module apc128bits(in, out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_a ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_b ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_cin ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_cout ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_d ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv1_m3_d ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv2_b ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv2_cin ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv2_cout ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv2_d ;
  wire _apc64_1_apc32_1_apc16_1_adder1_lv2_m3_d ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv1_a ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv1_b ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv1_cin ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv1_d ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv1_m3_d ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv2_cin ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv2_d ;
  wire _apc64_1_apc32_1_apc16_1_adder2_lv2_m3_d ;
  wire _apc64_1_apc32_1_apc16_1_half1_a ;
  wire _apc64_1_apc32_1_apc16_1_half1_cout ;
  wire _apc64_1_apc32_1_apc16_1_half1_s ;
  wire _apc64_1_apc32_1_apc16_1_half2_cout ;
  wire _apc64_1_apc32_1_apc16_1_half2_s ;
  wire _apc64_1_apc32_1_apc16_1_half3_cout ;
  wire _apc64_1_apc32_1_apc16_1_half3_s ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_a ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_b ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_cin ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_cout ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_d ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv1_m3_d ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv2_b ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv2_cin ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv2_cout ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv2_d ;
  wire _apc64_1_apc32_1_apc16_2_adder1_lv2_m3_d ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv1_a ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv1_b ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv1_cin ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv1_d ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv1_m3_d ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv2_cin ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv2_d ;
  wire _apc64_1_apc32_1_apc16_2_adder2_lv2_m3_d ;
  wire _apc64_1_apc32_1_apc16_2_half1_a ;
  wire _apc64_1_apc32_1_apc16_2_half1_cout ;
  wire _apc64_1_apc32_1_apc16_2_half1_s ;
  wire _apc64_1_apc32_1_apc16_2_half2_cout ;
  wire _apc64_1_apc32_1_apc16_2_half2_s ;
  wire _apc64_1_apc32_1_apc16_2_half3_cout ;
  wire _apc64_1_apc32_1_apc16_2_half3_s ;
  wire _apc64_1_apc32_1_out_0_;
  wire _apc64_1_apc32_1_out_1_;
  wire _apc64_1_apc32_1_out_2_;
  wire _apc64_1_apc32_1_out_3_;
  wire _apc64_1_apc32_1_out_4_;
  wire _apc64_1_apc32_1_out_5_;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_a ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_b ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_cin ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_cout ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_d ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv1_m3_d ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv2_b ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv2_cin ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv2_cout ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv2_d ;
  wire _apc64_1_apc32_2_apc16_1_adder1_lv2_m3_d ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv1_a ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv1_b ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv1_cin ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv1_d ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv1_m3_d ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv2_cin ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv2_d ;
  wire _apc64_1_apc32_2_apc16_1_adder2_lv2_m3_d ;
  wire _apc64_1_apc32_2_apc16_1_half1_a ;
  wire _apc64_1_apc32_2_apc16_1_half1_cout ;
  wire _apc64_1_apc32_2_apc16_1_half1_s ;
  wire _apc64_1_apc32_2_apc16_1_half2_cout ;
  wire _apc64_1_apc32_2_apc16_1_half2_s ;
  wire _apc64_1_apc32_2_apc16_1_half3_cout ;
  wire _apc64_1_apc32_2_apc16_1_half3_s ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_a ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_b ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_cin ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_cout ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_d ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv1_m3_d ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv2_b ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv2_cin ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv2_cout ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv2_d ;
  wire _apc64_1_apc32_2_apc16_2_adder1_lv2_m3_d ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv1_a ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv1_b ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv1_cin ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv1_d ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv1_m3_d ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv2_cin ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv2_d ;
  wire _apc64_1_apc32_2_apc16_2_adder2_lv2_m3_d ;
  wire _apc64_1_apc32_2_apc16_2_half1_a ;
  wire _apc64_1_apc32_2_apc16_2_half1_cout ;
  wire _apc64_1_apc32_2_apc16_2_half1_s ;
  wire _apc64_1_apc32_2_apc16_2_half2_cout ;
  wire _apc64_1_apc32_2_apc16_2_half2_s ;
  wire _apc64_1_apc32_2_apc16_2_half3_cout ;
  wire _apc64_1_apc32_2_apc16_2_half3_s ;
  wire _apc64_1_apc32_2_out_0_;
  wire _apc64_1_apc32_2_out_1_;
  wire _apc64_1_apc32_2_out_2_;
  wire _apc64_1_apc32_2_out_3_;
  wire _apc64_1_apc32_2_out_4_;
  wire _apc64_1_apc32_2_out_5_;
  wire _apc64_1_out_0_;
  wire _apc64_1_out_1_;
  wire _apc64_1_out_2_;
  wire _apc64_1_out_3_;
  wire _apc64_1_out_4_;
  wire _apc64_1_out_5_;
  wire _apc64_1_out_6_;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_a ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_b ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_cin ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_cout ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_d ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv1_m3_d ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv2_b ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv2_cin ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv2_cout ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv2_d ;
  wire _apc64_2_apc32_1_apc16_1_adder1_lv2_m3_d ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv1_a ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv1_b ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv1_cin ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv1_d ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv1_m3_d ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv2_cin ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv2_d ;
  wire _apc64_2_apc32_1_apc16_1_adder2_lv2_m3_d ;
  wire _apc64_2_apc32_1_apc16_1_half1_a ;
  wire _apc64_2_apc32_1_apc16_1_half1_cout ;
  wire _apc64_2_apc32_1_apc16_1_half1_s ;
  wire _apc64_2_apc32_1_apc16_1_half2_cout ;
  wire _apc64_2_apc32_1_apc16_1_half2_s ;
  wire _apc64_2_apc32_1_apc16_1_half3_cout ;
  wire _apc64_2_apc32_1_apc16_1_half3_s ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_a ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_b ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_cin ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_cout ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_d ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv1_m3_d ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv2_b ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv2_cin ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv2_cout ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv2_d ;
  wire _apc64_2_apc32_1_apc16_2_adder1_lv2_m3_d ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv1_a ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv1_b ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv1_cin ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv1_d ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv1_m3_d ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv2_cin ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv2_d ;
  wire _apc64_2_apc32_1_apc16_2_adder2_lv2_m3_d ;
  wire _apc64_2_apc32_1_apc16_2_half1_a ;
  wire _apc64_2_apc32_1_apc16_2_half1_cout ;
  wire _apc64_2_apc32_1_apc16_2_half1_s ;
  wire _apc64_2_apc32_1_apc16_2_half2_cout ;
  wire _apc64_2_apc32_1_apc16_2_half2_s ;
  wire _apc64_2_apc32_1_apc16_2_half3_cout ;
  wire _apc64_2_apc32_1_apc16_2_half3_s ;
  wire _apc64_2_apc32_1_out_0_;
  wire _apc64_2_apc32_1_out_1_;
  wire _apc64_2_apc32_1_out_2_;
  wire _apc64_2_apc32_1_out_3_;
  wire _apc64_2_apc32_1_out_4_;
  wire _apc64_2_apc32_1_out_5_;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_a ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_b ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_cin ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_cout ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_d ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv1_m3_d ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv2_b ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv2_cin ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv2_cout ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv2_d ;
  wire _apc64_2_apc32_2_apc16_1_adder1_lv2_m3_d ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv1_a ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv1_b ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv1_cin ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv1_d ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv1_m3_d ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv2_cin ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv2_d ;
  wire _apc64_2_apc32_2_apc16_1_adder2_lv2_m3_d ;
  wire _apc64_2_apc32_2_apc16_1_half1_a ;
  wire _apc64_2_apc32_2_apc16_1_half1_cout ;
  wire _apc64_2_apc32_2_apc16_1_half1_s ;
  wire _apc64_2_apc32_2_apc16_1_half2_cout ;
  wire _apc64_2_apc32_2_apc16_1_half2_s ;
  wire _apc64_2_apc32_2_apc16_1_half3_cout ;
  wire _apc64_2_apc32_2_apc16_1_half3_s ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_a ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_b ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_cin ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_cout ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_d ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv1_m3_d ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv2_b ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv2_cin ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv2_cout ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv2_d ;
  wire _apc64_2_apc32_2_apc16_2_adder1_lv2_m3_d ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv1_a ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv1_b ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv1_cin ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv1_d ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv1_m3_d ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv2_cin ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv2_d ;
  wire _apc64_2_apc32_2_apc16_2_adder2_lv2_m3_d ;
  wire _apc64_2_apc32_2_apc16_2_half1_a ;
  wire _apc64_2_apc32_2_apc16_2_half1_cout ;
  wire _apc64_2_apc32_2_apc16_2_half1_s ;
  wire _apc64_2_apc32_2_apc16_2_half2_cout ;
  wire _apc64_2_apc32_2_apc16_2_half2_s ;
  wire _apc64_2_apc32_2_apc16_2_half3_cout ;
  wire _apc64_2_apc32_2_apc16_2_half3_s ;
  wire _apc64_2_apc32_2_out_0_;
  wire _apc64_2_apc32_2_out_1_;
  wire _apc64_2_apc32_2_out_2_;
  wire _apc64_2_apc32_2_out_3_;
  wire _apc64_2_apc32_2_out_4_;
  wire _apc64_2_apc32_2_out_5_;
  wire _apc64_2_out_0_;
  wire _apc64_2_out_1_;
  wire _apc64_2_out_2_;
  wire _apc64_2_out_3_;
  wire _apc64_2_out_4_;
  wire _apc64_2_out_5_;
  wire _apc64_2_out_6_;
  input in_0_;
  input in_1_;
  input in_2_;
  input in_3_;
  input in_4_;
  input in_5_;
  input in_6_;
  input in_7_;
  input in_8_;
  input in_9_;
  input in_10_;
  input in_11_;
  input in_12_;
  input in_13_;
  input in_14_;
  input in_15_;
  input in_16_;
  input in_17_;
  input in_18_;
  input in_19_;
  input in_20_;
  input in_21_;
  input in_22_;
  input in_23_;
  input in_24_;
  input in_25_;
  input in_26_;
  input in_27_;
  input in_28_;
  input in_29_;
  input in_30_;
  input in_31_;
  input in_32_;
  input in_33_;
  input in_34_;
  input in_35_;
  input in_36_;
  input in_37_;
  input in_38_;
  input in_39_;
  input in_40_;
  input in_41_;
  input in_42_;
  input in_43_;
  input in_44_;
  input in_45_;
  input in_46_;
  input in_47_;
  input in_48_;
  input in_49_;
  input in_50_;
  input in_51_;
  input in_52_;
  input in_53_;
  input in_54_;
  input in_55_;
  input in_56_;
  input in_57_;
  input in_58_;
  input in_59_;
  input in_60_;
  input in_61_;
  input in_62_;
  input in_63_;
  input in_64_;
  input in_65_;
  input in_66_;
  input in_67_;
  input in_68_;
  input in_69_;
  input in_70_;
  input in_71_;
  input in_72_;
  input in_73_;
  input in_74_;
  input in_75_;
  input in_76_;
  input in_77_;
  input in_78_;
  input in_79_;
  input in_80_;
  input in_81_;
  input in_82_;
  input in_83_;
  input in_84_;
  input in_85_;
  input in_86_;
  input in_87_;
  input in_88_;
  input in_89_;
  input in_90_;
  input in_91_;
  input in_92_;
  input in_93_;
  input in_94_;
  input in_95_;
  input in_96_;
  input in_97_;
  input in_98_;
  input in_99_;
  input in_100_;
  input in_101_;
  input in_102_;
  input in_103_;
  input in_104_;
  input in_105_;
  input in_106_;
  input in_107_;
  input in_108_;
  input in_109_;
  input in_110_;
  input in_111_;
  input in_112_;
  input in_113_;
  input in_114_;
  input in_115_;
  input in_116_;
  input in_117_;
  input in_118_;
  input in_119_;
  input in_120_;
  input in_121_;
  input in_122_;
  input in_123_;
  input in_124_;
  input in_125_;
  input in_126_;
  input in_127_;
  output out_0_;
  output out_1_;
  output out_2_;
  output out_3_;
  output out_4_;
  output out_5_;
  output out_6_;
  output out_7_;
  or_ii _223_ (
    .a(_apc64_2_out_0_),
    .b(_apc64_1_out_0_),
    .c(_000_)
  );
  or_ii _224_ (
    .a(_apc64_2_out_1_),
    .b(_apc64_1_out_1_),
    .c(_001_)
  );
  and_ii _225_ (
    .a(_apc64_2_out_1_),
    .b(_apc64_1_out_1_),
    .c(_002_)
  );
  and_bi _226_ (
    .a(_001_),
    .b(_002_),
    .c(_003_)
  );
  or_bi _227_ (
    .a(_000_),
    .b(_003_),
    .c(_004_)
  );
  and_bi _228_ (
    .a(_000_),
    .b(_003_),
    .c(_005_)
  );
  and_bi _229_ (
    .a(_004_),
    .b(_005_),
    .c(out_1_)
  );
  maj_bii _230_ (
    .a(_000_),
    .b(_apc64_2_out_1_),
    .c(_apc64_1_out_1_),
    .d(_006_)
  );
  or_ii _231_ (
    .a(_apc64_2_out_2_),
    .b(_apc64_1_out_2_),
    .c(_007_)
  );
  and_ii _232_ (
    .a(_apc64_2_out_2_),
    .b(_apc64_1_out_2_),
    .c(_008_)
  );
  and_bi _233_ (
    .a(_007_),
    .b(_008_),
    .c(_009_)
  );
  or_bi _234_ (
    .a(_006_),
    .b(_009_),
    .c(_010_)
  );
  and_bi _235_ (
    .a(_006_),
    .b(_009_),
    .c(_011_)
  );
  and_bi _236_ (
    .a(_010_),
    .b(_011_),
    .c(out_2_)
  );
  maj_bii _237_ (
    .a(_006_),
    .b(_apc64_2_out_2_),
    .c(_apc64_1_out_2_),
    .d(_012_)
  );
  or_ii _238_ (
    .a(_apc64_2_out_3_),
    .b(_apc64_1_out_3_),
    .c(_013_)
  );
  and_ii _239_ (
    .a(_apc64_2_out_3_),
    .b(_apc64_1_out_3_),
    .c(_014_)
  );
  and_bi _240_ (
    .a(_013_),
    .b(_014_),
    .c(_015_)
  );
  or_bi _241_ (
    .a(_012_),
    .b(_015_),
    .c(_016_)
  );
  and_bi _242_ (
    .a(_012_),
    .b(_015_),
    .c(_017_)
  );
  and_bi _243_ (
    .a(_016_),
    .b(_017_),
    .c(out_3_)
  );
  maj_bii _244_ (
    .a(_012_),
    .b(_apc64_2_out_3_),
    .c(_apc64_1_out_3_),
    .d(_018_)
  );
  or_ii _245_ (
    .a(_apc64_2_out_4_),
    .b(_apc64_1_out_4_),
    .c(_019_)
  );
  and_ii _246_ (
    .a(_apc64_2_out_4_),
    .b(_apc64_1_out_4_),
    .c(_020_)
  );
  and_bi _247_ (
    .a(_019_),
    .b(_020_),
    .c(_021_)
  );
  or_bi _248_ (
    .a(_018_),
    .b(_021_),
    .c(_022_)
  );
  and_bi _249_ (
    .a(_018_),
    .b(_021_),
    .c(_023_)
  );
  and_bi _250_ (
    .a(_022_),
    .b(_023_),
    .c(out_4_)
  );
  maj_bii _251_ (
    .a(_018_),
    .b(_apc64_2_out_4_),
    .c(_apc64_1_out_4_),
    .d(_024_)
  );
  or_ii _252_ (
    .a(_apc64_2_out_5_),
    .b(_apc64_1_out_5_),
    .c(_025_)
  );
  and_ii _253_ (
    .a(_apc64_2_out_5_),
    .b(_apc64_1_out_5_),
    .c(_026_)
  );
  and_bi _254_ (
    .a(_025_),
    .b(_026_),
    .c(_027_)
  );
  or_bi _255_ (
    .a(_024_),
    .b(_027_),
    .c(_028_)
  );
  and_bi _256_ (
    .a(_024_),
    .b(_027_),
    .c(_029_)
  );
  and_bi _257_ (
    .a(_028_),
    .b(_029_),
    .c(out_5_)
  );
  maj_bii _258_ (
    .a(_024_),
    .b(_apc64_2_out_5_),
    .c(_apc64_1_out_5_),
    .d(_030_)
  );
  or_ii _259_ (
    .a(_apc64_2_out_6_),
    .b(_apc64_1_out_6_),
    .c(_031_)
  );
  and_ii _260_ (
    .a(_apc64_2_out_6_),
    .b(_apc64_1_out_6_),
    .c(_032_)
  );
  and_bi _261_ (
    .a(_031_),
    .b(_032_),
    .c(_033_)
  );
  or_bi _262_ (
    .a(_030_),
    .b(_033_),
    .c(_034_)
  );
  and_bi _263_ (
    .a(_030_),
    .b(_033_),
    .c(_035_)
  );
  and_bi _264_ (
    .a(_034_),
    .b(_035_),
    .c(out_6_)
  );
  maj_bbi _265_ (
    .a(_apc64_2_out_6_),
    .b(_apc64_1_out_6_),
    .c(_030_),
    .d(out_7_)
  );
  and_ii _266_ (
    .a(_apc64_2_out_0_),
    .b(_apc64_1_out_0_),
    .c(_036_)
  );
  and_bi _267_ (
    .a(_000_),
    .b(_036_),
    .c(out_0_)
  );
  or_ii _268_ (
    .a(_apc64_1_apc32_2_out_0_),
    .b(_apc64_1_apc32_1_out_0_),
    .c(_037_)
  );
  or_ii _269_ (
    .a(_apc64_1_apc32_2_out_1_),
    .b(_apc64_1_apc32_1_out_1_),
    .c(_038_)
  );
  and_ii _270_ (
    .a(_apc64_1_apc32_2_out_1_),
    .b(_apc64_1_apc32_1_out_1_),
    .c(_039_)
  );
  and_bi _271_ (
    .a(_038_),
    .b(_039_),
    .c(_040_)
  );
  or_bi _272_ (
    .a(_037_),
    .b(_040_),
    .c(_041_)
  );
  and_bi _273_ (
    .a(_037_),
    .b(_040_),
    .c(_042_)
  );
  and_bi _274_ (
    .a(_041_),
    .b(_042_),
    .c(_apc64_1_out_1_)
  );
  maj_bii _275_ (
    .a(_037_),
    .b(_apc64_1_apc32_2_out_1_),
    .c(_apc64_1_apc32_1_out_1_),
    .d(_043_)
  );
  or_ii _276_ (
    .a(_apc64_1_apc32_2_out_2_),
    .b(_apc64_1_apc32_1_out_2_),
    .c(_044_)
  );
  and_ii _277_ (
    .a(_apc64_1_apc32_2_out_2_),
    .b(_apc64_1_apc32_1_out_2_),
    .c(_045_)
  );
  and_bi _278_ (
    .a(_044_),
    .b(_045_),
    .c(_046_)
  );
  or_bi _279_ (
    .a(_043_),
    .b(_046_),
    .c(_047_)
  );
  and_bi _280_ (
    .a(_043_),
    .b(_046_),
    .c(_048_)
  );
  and_bi _281_ (
    .a(_047_),
    .b(_048_),
    .c(_apc64_1_out_2_)
  );
  maj_bii _282_ (
    .a(_043_),
    .b(_apc64_1_apc32_2_out_2_),
    .c(_apc64_1_apc32_1_out_2_),
    .d(_049_)
  );
  or_ii _283_ (
    .a(_apc64_1_apc32_2_out_3_),
    .b(_apc64_1_apc32_1_out_3_),
    .c(_050_)
  );
  and_ii _284_ (
    .a(_apc64_1_apc32_2_out_3_),
    .b(_apc64_1_apc32_1_out_3_),
    .c(_051_)
  );
  and_bi _285_ (
    .a(_050_),
    .b(_051_),
    .c(_052_)
  );
  or_bi _286_ (
    .a(_049_),
    .b(_052_),
    .c(_053_)
  );
  and_bi _287_ (
    .a(_049_),
    .b(_052_),
    .c(_054_)
  );
  and_bi _288_ (
    .a(_053_),
    .b(_054_),
    .c(_apc64_1_out_3_)
  );
  maj_bii _289_ (
    .a(_049_),
    .b(_apc64_1_apc32_2_out_3_),
    .c(_apc64_1_apc32_1_out_3_),
    .d(_055_)
  );
  or_ii _290_ (
    .a(_apc64_1_apc32_2_out_4_),
    .b(_apc64_1_apc32_1_out_4_),
    .c(_056_)
  );
  and_ii _291_ (
    .a(_apc64_1_apc32_2_out_4_),
    .b(_apc64_1_apc32_1_out_4_),
    .c(_057_)
  );
  and_bi _292_ (
    .a(_056_),
    .b(_057_),
    .c(_058_)
  );
  or_bi _293_ (
    .a(_055_),
    .b(_058_),
    .c(_059_)
  );
  and_bi _294_ (
    .a(_055_),
    .b(_058_),
    .c(_060_)
  );
  and_bi _295_ (
    .a(_059_),
    .b(_060_),
    .c(_apc64_1_out_4_)
  );
  maj_bii _296_ (
    .a(_055_),
    .b(_apc64_1_apc32_2_out_4_),
    .c(_apc64_1_apc32_1_out_4_),
    .d(_061_)
  );
  or_ii _297_ (
    .a(_apc64_1_apc32_2_out_5_),
    .b(_apc64_1_apc32_1_out_5_),
    .c(_062_)
  );
  and_ii _298_ (
    .a(_apc64_1_apc32_2_out_5_),
    .b(_apc64_1_apc32_1_out_5_),
    .c(_063_)
  );
  and_bi _299_ (
    .a(_062_),
    .b(_063_),
    .c(_064_)
  );
  or_bi _300_ (
    .a(_061_),
    .b(_064_),
    .c(_065_)
  );
  and_bi _301_ (
    .a(_061_),
    .b(_064_),
    .c(_066_)
  );
  and_bi _302_ (
    .a(_065_),
    .b(_066_),
    .c(_apc64_1_out_5_)
  );
  and_ii _303_ (
    .a(_apc64_1_apc32_2_out_0_),
    .b(_apc64_1_apc32_1_out_0_),
    .c(_067_)
  );
  and_bi _304_ (
    .a(_037_),
    .b(_067_),
    .c(_apc64_1_out_0_)
  );
  maj_bbi _305_ (
    .a(_apc64_1_apc32_2_out_5_),
    .b(_apc64_1_apc32_1_out_5_),
    .c(_061_),
    .d(_apc64_1_out_6_)
  );
  or_ii _306_ (
    .a(1'b0),
    .b(1'b0),
    .c(_068_)
  );
  or_ii _307_ (
    .a(_apc64_1_apc32_1_apc16_2_half1_s ),
    .b(_apc64_1_apc32_1_apc16_1_half1_s ),
    .c(_069_)
  );
  and_ii _308_ (
    .a(_apc64_1_apc32_1_apc16_2_half1_s ),
    .b(_apc64_1_apc32_1_apc16_1_half1_s ),
    .c(_070_)
  );
  and_bi _309_ (
    .a(_069_),
    .b(_070_),
    .c(_071_)
  );
  or_bi _310_ (
    .a(_068_),
    .b(_071_),
    .c(_072_)
  );
  and_bi _311_ (
    .a(_068_),
    .b(_071_),
    .c(_073_)
  );
  and_bi _312_ (
    .a(_072_),
    .b(_073_),
    .c(_apc64_1_apc32_1_out_1_)
  );
  maj_bii _313_ (
    .a(_068_),
    .b(_apc64_1_apc32_1_apc16_2_half1_s ),
    .c(_apc64_1_apc32_1_apc16_1_half1_s ),
    .d(_074_)
  );
  or_ii _314_ (
    .a(_apc64_1_apc32_1_apc16_2_half2_s ),
    .b(_apc64_1_apc32_1_apc16_1_half2_s ),
    .c(_075_)
  );
  and_ii _315_ (
    .a(_apc64_1_apc32_1_apc16_2_half2_s ),
    .b(_apc64_1_apc32_1_apc16_1_half2_s ),
    .c(_076_)
  );
  and_bi _316_ (
    .a(_075_),
    .b(_076_),
    .c(_077_)
  );
  or_bi _317_ (
    .a(_074_),
    .b(_077_),
    .c(_078_)
  );
  and_bi _318_ (
    .a(_074_),
    .b(_077_),
    .c(_079_)
  );
  and_bi _319_ (
    .a(_078_),
    .b(_079_),
    .c(_apc64_1_apc32_1_out_2_)
  );
  maj_bii _320_ (
    .a(_074_),
    .b(_apc64_1_apc32_1_apc16_2_half2_s ),
    .c(_apc64_1_apc32_1_apc16_1_half2_s ),
    .d(_080_)
  );
  or_ii _321_ (
    .a(_apc64_1_apc32_1_apc16_2_half3_s ),
    .b(_apc64_1_apc32_1_apc16_1_half3_s ),
    .c(_081_)
  );
  and_ii _322_ (
    .a(_apc64_1_apc32_1_apc16_2_half3_s ),
    .b(_apc64_1_apc32_1_apc16_1_half3_s ),
    .c(_082_)
  );
  and_bi _323_ (
    .a(_081_),
    .b(_082_),
    .c(_083_)
  );
  or_bi _324_ (
    .a(_080_),
    .b(_083_),
    .c(_084_)
  );
  and_bi _325_ (
    .a(_080_),
    .b(_083_),
    .c(_085_)
  );
  and_bi _326_ (
    .a(_084_),
    .b(_085_),
    .c(_apc64_1_apc32_1_out_3_)
  );
  maj_bii _327_ (
    .a(_080_),
    .b(_apc64_1_apc32_1_apc16_2_half3_s ),
    .c(_apc64_1_apc32_1_apc16_1_half3_s ),
    .d(_086_)
  );
  or_ii _328_ (
    .a(_apc64_1_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_1_apc16_1_half3_cout ),
    .c(_087_)
  );
  and_ii _329_ (
    .a(_apc64_1_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_1_apc16_1_half3_cout ),
    .c(_088_)
  );
  and_bi _330_ (
    .a(_087_),
    .b(_088_),
    .c(_089_)
  );
  or_bi _331_ (
    .a(_086_),
    .b(_089_),
    .c(_090_)
  );
  and_bi _332_ (
    .a(_086_),
    .b(_089_),
    .c(_091_)
  );
  and_bi _333_ (
    .a(_090_),
    .b(_091_),
    .c(_apc64_1_apc32_1_out_4_)
  );
  and_ii _334_ (
    .a(1'b0),
    .b(1'b0),
    .c(_092_)
  );
  and_bi _335_ (
    .a(_068_),
    .b(_092_),
    .c(_apc64_1_apc32_1_out_0_)
  );
  maj_bbi _336_ (
    .a(_apc64_1_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_1_apc16_1_half3_cout ),
    .c(_086_),
    .d(_apc64_1_apc32_1_out_5_)
  );
  or_bb _337_ (
    .a(in_113_),
    .b(in_112_),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_a )
  );
  and_bb _338_ (
    .a(in_115_),
    .b(in_114_),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_b )
  );
  or_bb _339_ (
    .a(in_117_),
    .b(in_116_),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_cin )
  );
  and_bb _340_ (
    .a(in_119_),
    .b(in_118_),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv1_a )
  );
  or_bb _341_ (
    .a(in_121_),
    .b(in_120_),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv1_b )
  );
  and_bb _342_ (
    .a(in_123_),
    .b(in_122_),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv1_cin )
  );
  or_bb _343_ (
    .a(in_125_),
    .b(in_124_),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv2_cin )
  );
  and_bb _344_ (
    .a(in_127_),
    .b(in_126_),
    .c(_apc64_1_apc32_1_apc16_1_half1_a )
  );
  maj_bbb _345_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv1_cin ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv1_b ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_a ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _346_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv1_b ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv1_a ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_cin ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv1_d )
  );
  maj_bbi _347_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv1_d ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv1_cin ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _348_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv2_cin ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_b ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _349_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv2_b ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv1_cout ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv2_d )
  );
  maj_bbi _350_ (
    .a(_apc64_1_apc32_1_apc16_1_adder1_lv2_d ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_cin ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv2_cout ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _351_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv1_cin ),
    .b(_apc64_1_apc32_1_apc16_1_adder2_lv1_b ),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv1_a ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv2_b )
  );
  maj_bbi _352_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv1_b ),
    .b(_apc64_1_apc32_1_apc16_1_adder2_lv1_a ),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv1_cin ),
    .d(_apc64_1_apc32_1_apc16_1_adder2_lv1_d )
  );
  maj_bbi _353_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv1_d ),
    .b(_apc64_1_apc32_1_apc16_1_adder2_lv1_cin ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv2_b ),
    .d(_apc64_1_apc32_1_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _354_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv2_cin ),
    .b(_apc64_1_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .d(_apc64_1_apc32_1_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _355_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .c(_apc64_1_apc32_1_apc16_1_adder2_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_1_adder2_lv2_d )
  );
  maj_bbi _356_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv2_d ),
    .b(_apc64_1_apc32_1_apc16_1_adder2_lv2_cin ),
    .c(_apc64_1_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _357_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_1_apc16_1_half1_a ),
    .c(_apc64_1_apc32_1_apc16_1_half1_cout )
  );
  or_bb _358_ (
    .a(_apc64_1_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_1_apc16_1_half1_a ),
    .c(_093_)
  );
  and_bi _359_ (
    .a(_093_),
    .b(_apc64_1_apc32_1_apc16_1_half1_cout ),
    .c(_apc64_1_apc32_1_apc16_1_half1_s )
  );
  and_bb _360_ (
    .a(_apc64_1_apc32_1_apc16_1_half1_cout ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_apc64_1_apc32_1_apc16_1_half2_cout )
  );
  or_bb _361_ (
    .a(_apc64_1_apc32_1_apc16_1_half1_cout ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_094_)
  );
  and_bi _362_ (
    .a(_094_),
    .b(_apc64_1_apc32_1_apc16_1_half2_cout ),
    .c(_apc64_1_apc32_1_apc16_1_half2_s )
  );
  and_bb _363_ (
    .a(_apc64_1_apc32_1_apc16_1_half2_cout ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_apc64_1_apc32_1_apc16_1_half3_cout )
  );
  or_bb _364_ (
    .a(_apc64_1_apc32_1_apc16_1_half2_cout ),
    .b(_apc64_1_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_095_)
  );
  and_bi _365_ (
    .a(_095_),
    .b(_apc64_1_apc32_1_apc16_1_half3_cout ),
    .c(_apc64_1_apc32_1_apc16_1_half3_s )
  );
  or_bb _366_ (
    .a(in_97_),
    .b(in_96_),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_a )
  );
  and_bb _367_ (
    .a(in_99_),
    .b(in_98_),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_b )
  );
  or_bb _368_ (
    .a(in_101_),
    .b(in_100_),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_cin )
  );
  and_bb _369_ (
    .a(in_103_),
    .b(in_102_),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv1_a )
  );
  or_bb _370_ (
    .a(in_105_),
    .b(in_104_),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv1_b )
  );
  and_bb _371_ (
    .a(in_107_),
    .b(in_106_),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv1_cin )
  );
  or_bb _372_ (
    .a(in_109_),
    .b(in_108_),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv2_cin )
  );
  and_bb _373_ (
    .a(in_111_),
    .b(in_110_),
    .c(_apc64_1_apc32_1_apc16_2_half1_a )
  );
  maj_bbb _374_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv1_cin ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv1_b ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_a ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _375_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv1_b ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv1_a ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_cin ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv1_d )
  );
  maj_bbi _376_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv1_d ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv1_cin ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _377_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv2_cin ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_b ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _378_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv2_b ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv1_cout ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv2_d )
  );
  maj_bbi _379_ (
    .a(_apc64_1_apc32_1_apc16_2_adder1_lv2_d ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_cin ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv2_cout ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _380_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv1_cin ),
    .b(_apc64_1_apc32_1_apc16_2_adder2_lv1_b ),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv1_a ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv2_b )
  );
  maj_bbi _381_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv1_b ),
    .b(_apc64_1_apc32_1_apc16_2_adder2_lv1_a ),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv1_cin ),
    .d(_apc64_1_apc32_1_apc16_2_adder2_lv1_d )
  );
  maj_bbi _382_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv1_d ),
    .b(_apc64_1_apc32_1_apc16_2_adder2_lv1_cin ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv2_b ),
    .d(_apc64_1_apc32_1_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _383_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv2_cin ),
    .b(_apc64_1_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .d(_apc64_1_apc32_1_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _384_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .c(_apc64_1_apc32_1_apc16_2_adder2_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_2_adder2_lv2_d )
  );
  maj_bbi _385_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv2_d ),
    .b(_apc64_1_apc32_1_apc16_2_adder2_lv2_cin ),
    .c(_apc64_1_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc64_1_apc32_1_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _386_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_1_apc16_2_half1_a ),
    .c(_apc64_1_apc32_1_apc16_2_half1_cout )
  );
  or_bb _387_ (
    .a(_apc64_1_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_1_apc16_2_half1_a ),
    .c(_096_)
  );
  and_bi _388_ (
    .a(_096_),
    .b(_apc64_1_apc32_1_apc16_2_half1_cout ),
    .c(_apc64_1_apc32_1_apc16_2_half1_s )
  );
  and_bb _389_ (
    .a(_apc64_1_apc32_1_apc16_2_half1_cout ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_apc64_1_apc32_1_apc16_2_half2_cout )
  );
  or_bb _390_ (
    .a(_apc64_1_apc32_1_apc16_2_half1_cout ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_097_)
  );
  and_bi _391_ (
    .a(_097_),
    .b(_apc64_1_apc32_1_apc16_2_half2_cout ),
    .c(_apc64_1_apc32_1_apc16_2_half2_s )
  );
  and_bb _392_ (
    .a(_apc64_1_apc32_1_apc16_2_half2_cout ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_apc64_1_apc32_1_apc16_2_half3_cout )
  );
  or_bb _393_ (
    .a(_apc64_1_apc32_1_apc16_2_half2_cout ),
    .b(_apc64_1_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_098_)
  );
  and_bi _394_ (
    .a(_098_),
    .b(_apc64_1_apc32_1_apc16_2_half3_cout ),
    .c(_apc64_1_apc32_1_apc16_2_half3_s )
  );
  or_ii _395_ (
    .a(1'b0),
    .b(1'b0),
    .c(_099_)
  );
  or_ii _396_ (
    .a(_apc64_1_apc32_2_apc16_2_half1_s ),
    .b(_apc64_1_apc32_2_apc16_1_half1_s ),
    .c(_100_)
  );
  and_ii _397_ (
    .a(_apc64_1_apc32_2_apc16_2_half1_s ),
    .b(_apc64_1_apc32_2_apc16_1_half1_s ),
    .c(_101_)
  );
  and_bi _398_ (
    .a(_100_),
    .b(_101_),
    .c(_102_)
  );
  or_bi _399_ (
    .a(_099_),
    .b(_102_),
    .c(_103_)
  );
  and_bi _400_ (
    .a(_099_),
    .b(_102_),
    .c(_104_)
  );
  and_bi _401_ (
    .a(_103_),
    .b(_104_),
    .c(_apc64_1_apc32_2_out_1_)
  );
  maj_bii _402_ (
    .a(_099_),
    .b(_apc64_1_apc32_2_apc16_2_half1_s ),
    .c(_apc64_1_apc32_2_apc16_1_half1_s ),
    .d(_105_)
  );
  or_ii _403_ (
    .a(_apc64_1_apc32_2_apc16_2_half2_s ),
    .b(_apc64_1_apc32_2_apc16_1_half2_s ),
    .c(_106_)
  );
  and_ii _404_ (
    .a(_apc64_1_apc32_2_apc16_2_half2_s ),
    .b(_apc64_1_apc32_2_apc16_1_half2_s ),
    .c(_107_)
  );
  and_bi _405_ (
    .a(_106_),
    .b(_107_),
    .c(_108_)
  );
  or_bi _406_ (
    .a(_105_),
    .b(_108_),
    .c(_109_)
  );
  and_bi _407_ (
    .a(_105_),
    .b(_108_),
    .c(_110_)
  );
  and_bi _408_ (
    .a(_109_),
    .b(_110_),
    .c(_apc64_1_apc32_2_out_2_)
  );
  maj_bii _409_ (
    .a(_105_),
    .b(_apc64_1_apc32_2_apc16_2_half2_s ),
    .c(_apc64_1_apc32_2_apc16_1_half2_s ),
    .d(_111_)
  );
  or_ii _410_ (
    .a(_apc64_1_apc32_2_apc16_2_half3_s ),
    .b(_apc64_1_apc32_2_apc16_1_half3_s ),
    .c(_112_)
  );
  and_ii _411_ (
    .a(_apc64_1_apc32_2_apc16_2_half3_s ),
    .b(_apc64_1_apc32_2_apc16_1_half3_s ),
    .c(_113_)
  );
  and_bi _412_ (
    .a(_112_),
    .b(_113_),
    .c(_114_)
  );
  or_bi _413_ (
    .a(_111_),
    .b(_114_),
    .c(_115_)
  );
  and_bi _414_ (
    .a(_111_),
    .b(_114_),
    .c(_116_)
  );
  and_bi _415_ (
    .a(_115_),
    .b(_116_),
    .c(_apc64_1_apc32_2_out_3_)
  );
  maj_bii _416_ (
    .a(_111_),
    .b(_apc64_1_apc32_2_apc16_2_half3_s ),
    .c(_apc64_1_apc32_2_apc16_1_half3_s ),
    .d(_117_)
  );
  or_ii _417_ (
    .a(_apc64_1_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_2_apc16_1_half3_cout ),
    .c(_118_)
  );
  and_ii _418_ (
    .a(_apc64_1_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_2_apc16_1_half3_cout ),
    .c(_119_)
  );
  and_bi _419_ (
    .a(_118_),
    .b(_119_),
    .c(_120_)
  );
  or_bi _420_ (
    .a(_117_),
    .b(_120_),
    .c(_121_)
  );
  and_bi _421_ (
    .a(_117_),
    .b(_120_),
    .c(_122_)
  );
  and_bi _422_ (
    .a(_121_),
    .b(_122_),
    .c(_apc64_1_apc32_2_out_4_)
  );
  and_ii _423_ (
    .a(1'b0),
    .b(1'b0),
    .c(_123_)
  );
  and_bi _424_ (
    .a(_099_),
    .b(_123_),
    .c(_apc64_1_apc32_2_out_0_)
  );
  maj_bbi _425_ (
    .a(_apc64_1_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_1_apc32_2_apc16_1_half3_cout ),
    .c(_117_),
    .d(_apc64_1_apc32_2_out_5_)
  );
  or_bb _426_ (
    .a(in_81_),
    .b(in_80_),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_a )
  );
  and_bb _427_ (
    .a(in_83_),
    .b(in_82_),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_b )
  );
  or_bb _428_ (
    .a(in_85_),
    .b(in_84_),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_cin )
  );
  and_bb _429_ (
    .a(in_87_),
    .b(in_86_),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv1_a )
  );
  or_bb _430_ (
    .a(in_89_),
    .b(in_88_),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv1_b )
  );
  and_bb _431_ (
    .a(in_91_),
    .b(in_90_),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv1_cin )
  );
  or_bb _432_ (
    .a(in_93_),
    .b(in_92_),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv2_cin )
  );
  and_bb _433_ (
    .a(in_95_),
    .b(in_94_),
    .c(_apc64_1_apc32_2_apc16_1_half1_a )
  );
  maj_bbb _434_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv1_cin ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv1_b ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_a ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _435_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv1_b ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv1_a ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_cin ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv1_d )
  );
  maj_bbi _436_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv1_d ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv1_cin ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _437_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv2_cin ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_b ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _438_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv2_b ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv1_cout ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv2_d )
  );
  maj_bbi _439_ (
    .a(_apc64_1_apc32_2_apc16_1_adder1_lv2_d ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_cin ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv2_cout ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _440_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv1_cin ),
    .b(_apc64_1_apc32_2_apc16_1_adder2_lv1_b ),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv1_a ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv2_b )
  );
  maj_bbi _441_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv1_b ),
    .b(_apc64_1_apc32_2_apc16_1_adder2_lv1_a ),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv1_cin ),
    .d(_apc64_1_apc32_2_apc16_1_adder2_lv1_d )
  );
  maj_bbi _442_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv1_d ),
    .b(_apc64_1_apc32_2_apc16_1_adder2_lv1_cin ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv2_b ),
    .d(_apc64_1_apc32_2_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _443_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv2_cin ),
    .b(_apc64_1_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .d(_apc64_1_apc32_2_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _444_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .c(_apc64_1_apc32_2_apc16_1_adder2_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_1_adder2_lv2_d )
  );
  maj_bbi _445_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv2_d ),
    .b(_apc64_1_apc32_2_apc16_1_adder2_lv2_cin ),
    .c(_apc64_1_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _446_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_2_apc16_1_half1_a ),
    .c(_apc64_1_apc32_2_apc16_1_half1_cout )
  );
  or_bb _447_ (
    .a(_apc64_1_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_2_apc16_1_half1_a ),
    .c(_124_)
  );
  and_bi _448_ (
    .a(_124_),
    .b(_apc64_1_apc32_2_apc16_1_half1_cout ),
    .c(_apc64_1_apc32_2_apc16_1_half1_s )
  );
  and_bb _449_ (
    .a(_apc64_1_apc32_2_apc16_1_half1_cout ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_apc64_1_apc32_2_apc16_1_half2_cout )
  );
  or_bb _450_ (
    .a(_apc64_1_apc32_2_apc16_1_half1_cout ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_125_)
  );
  and_bi _451_ (
    .a(_125_),
    .b(_apc64_1_apc32_2_apc16_1_half2_cout ),
    .c(_apc64_1_apc32_2_apc16_1_half2_s )
  );
  and_bb _452_ (
    .a(_apc64_1_apc32_2_apc16_1_half2_cout ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_apc64_1_apc32_2_apc16_1_half3_cout )
  );
  or_bb _453_ (
    .a(_apc64_1_apc32_2_apc16_1_half2_cout ),
    .b(_apc64_1_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_126_)
  );
  and_bi _454_ (
    .a(_126_),
    .b(_apc64_1_apc32_2_apc16_1_half3_cout ),
    .c(_apc64_1_apc32_2_apc16_1_half3_s )
  );
  or_bb _455_ (
    .a(in_65_),
    .b(in_64_),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_a )
  );
  and_bb _456_ (
    .a(in_67_),
    .b(in_66_),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_b )
  );
  or_bb _457_ (
    .a(in_69_),
    .b(in_68_),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_cin )
  );
  and_bb _458_ (
    .a(in_71_),
    .b(in_70_),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv1_a )
  );
  or_bb _459_ (
    .a(in_73_),
    .b(in_72_),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv1_b )
  );
  and_bb _460_ (
    .a(in_75_),
    .b(in_74_),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv1_cin )
  );
  or_bb _461_ (
    .a(in_77_),
    .b(in_76_),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv2_cin )
  );
  and_bb _462_ (
    .a(in_79_),
    .b(in_78_),
    .c(_apc64_1_apc32_2_apc16_2_half1_a )
  );
  maj_bbb _463_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv1_cin ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv1_b ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_a ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _464_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv1_b ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv1_a ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_cin ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv1_d )
  );
  maj_bbi _465_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv1_d ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv1_cin ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _466_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv2_cin ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_b ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _467_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv2_b ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv1_cout ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv2_d )
  );
  maj_bbi _468_ (
    .a(_apc64_1_apc32_2_apc16_2_adder1_lv2_d ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_cin ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv2_cout ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _469_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv1_cin ),
    .b(_apc64_1_apc32_2_apc16_2_adder2_lv1_b ),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv1_a ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv2_b )
  );
  maj_bbi _470_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv1_b ),
    .b(_apc64_1_apc32_2_apc16_2_adder2_lv1_a ),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv1_cin ),
    .d(_apc64_1_apc32_2_apc16_2_adder2_lv1_d )
  );
  maj_bbi _471_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv1_d ),
    .b(_apc64_1_apc32_2_apc16_2_adder2_lv1_cin ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv2_b ),
    .d(_apc64_1_apc32_2_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _472_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv2_cin ),
    .b(_apc64_1_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .d(_apc64_1_apc32_2_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _473_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .c(_apc64_1_apc32_2_apc16_2_adder2_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_2_adder2_lv2_d )
  );
  maj_bbi _474_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv2_d ),
    .b(_apc64_1_apc32_2_apc16_2_adder2_lv2_cin ),
    .c(_apc64_1_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc64_1_apc32_2_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _475_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_2_apc16_2_half1_a ),
    .c(_apc64_1_apc32_2_apc16_2_half1_cout )
  );
  or_bb _476_ (
    .a(_apc64_1_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_1_apc32_2_apc16_2_half1_a ),
    .c(_127_)
  );
  and_bi _477_ (
    .a(_127_),
    .b(_apc64_1_apc32_2_apc16_2_half1_cout ),
    .c(_apc64_1_apc32_2_apc16_2_half1_s )
  );
  and_bb _478_ (
    .a(_apc64_1_apc32_2_apc16_2_half1_cout ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_apc64_1_apc32_2_apc16_2_half2_cout )
  );
  or_bb _479_ (
    .a(_apc64_1_apc32_2_apc16_2_half1_cout ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_128_)
  );
  and_bi _480_ (
    .a(_128_),
    .b(_apc64_1_apc32_2_apc16_2_half2_cout ),
    .c(_apc64_1_apc32_2_apc16_2_half2_s )
  );
  and_bb _481_ (
    .a(_apc64_1_apc32_2_apc16_2_half2_cout ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_apc64_1_apc32_2_apc16_2_half3_cout )
  );
  or_bb _482_ (
    .a(_apc64_1_apc32_2_apc16_2_half2_cout ),
    .b(_apc64_1_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_129_)
  );
  and_bi _483_ (
    .a(_129_),
    .b(_apc64_1_apc32_2_apc16_2_half3_cout ),
    .c(_apc64_1_apc32_2_apc16_2_half3_s )
  );
  or_ii _484_ (
    .a(_apc64_2_apc32_2_out_0_),
    .b(_apc64_2_apc32_1_out_0_),
    .c(_130_)
  );
  or_ii _485_ (
    .a(_apc64_2_apc32_2_out_1_),
    .b(_apc64_2_apc32_1_out_1_),
    .c(_131_)
  );
  and_ii _486_ (
    .a(_apc64_2_apc32_2_out_1_),
    .b(_apc64_2_apc32_1_out_1_),
    .c(_132_)
  );
  and_bi _487_ (
    .a(_131_),
    .b(_132_),
    .c(_133_)
  );
  or_bi _488_ (
    .a(_130_),
    .b(_133_),
    .c(_134_)
  );
  and_bi _489_ (
    .a(_130_),
    .b(_133_),
    .c(_135_)
  );
  and_bi _490_ (
    .a(_134_),
    .b(_135_),
    .c(_apc64_2_out_1_)
  );
  maj_bii _491_ (
    .a(_130_),
    .b(_apc64_2_apc32_2_out_1_),
    .c(_apc64_2_apc32_1_out_1_),
    .d(_136_)
  );
  or_ii _492_ (
    .a(_apc64_2_apc32_2_out_2_),
    .b(_apc64_2_apc32_1_out_2_),
    .c(_137_)
  );
  and_ii _493_ (
    .a(_apc64_2_apc32_2_out_2_),
    .b(_apc64_2_apc32_1_out_2_),
    .c(_138_)
  );
  and_bi _494_ (
    .a(_137_),
    .b(_138_),
    .c(_139_)
  );
  or_bi _495_ (
    .a(_136_),
    .b(_139_),
    .c(_140_)
  );
  and_bi _496_ (
    .a(_136_),
    .b(_139_),
    .c(_141_)
  );
  and_bi _497_ (
    .a(_140_),
    .b(_141_),
    .c(_apc64_2_out_2_)
  );
  maj_bii _498_ (
    .a(_136_),
    .b(_apc64_2_apc32_2_out_2_),
    .c(_apc64_2_apc32_1_out_2_),
    .d(_142_)
  );
  or_ii _499_ (
    .a(_apc64_2_apc32_2_out_3_),
    .b(_apc64_2_apc32_1_out_3_),
    .c(_143_)
  );
  and_ii _500_ (
    .a(_apc64_2_apc32_2_out_3_),
    .b(_apc64_2_apc32_1_out_3_),
    .c(_144_)
  );
  and_bi _501_ (
    .a(_143_),
    .b(_144_),
    .c(_145_)
  );
  or_bi _502_ (
    .a(_142_),
    .b(_145_),
    .c(_146_)
  );
  and_bi _503_ (
    .a(_142_),
    .b(_145_),
    .c(_147_)
  );
  and_bi _504_ (
    .a(_146_),
    .b(_147_),
    .c(_apc64_2_out_3_)
  );
  maj_bii _505_ (
    .a(_142_),
    .b(_apc64_2_apc32_2_out_3_),
    .c(_apc64_2_apc32_1_out_3_),
    .d(_148_)
  );
  or_ii _506_ (
    .a(_apc64_2_apc32_2_out_4_),
    .b(_apc64_2_apc32_1_out_4_),
    .c(_149_)
  );
  and_ii _507_ (
    .a(_apc64_2_apc32_2_out_4_),
    .b(_apc64_2_apc32_1_out_4_),
    .c(_150_)
  );
  and_bi _508_ (
    .a(_149_),
    .b(_150_),
    .c(_151_)
  );
  or_bi _509_ (
    .a(_148_),
    .b(_151_),
    .c(_152_)
  );
  and_bi _510_ (
    .a(_148_),
    .b(_151_),
    .c(_153_)
  );
  and_bi _511_ (
    .a(_152_),
    .b(_153_),
    .c(_apc64_2_out_4_)
  );
  maj_bii _512_ (
    .a(_148_),
    .b(_apc64_2_apc32_2_out_4_),
    .c(_apc64_2_apc32_1_out_4_),
    .d(_154_)
  );
  or_ii _513_ (
    .a(_apc64_2_apc32_2_out_5_),
    .b(_apc64_2_apc32_1_out_5_),
    .c(_155_)
  );
  and_ii _514_ (
    .a(_apc64_2_apc32_2_out_5_),
    .b(_apc64_2_apc32_1_out_5_),
    .c(_156_)
  );
  and_bi _515_ (
    .a(_155_),
    .b(_156_),
    .c(_157_)
  );
  or_bi _516_ (
    .a(_154_),
    .b(_157_),
    .c(_158_)
  );
  and_bi _517_ (
    .a(_154_),
    .b(_157_),
    .c(_159_)
  );
  and_bi _518_ (
    .a(_158_),
    .b(_159_),
    .c(_apc64_2_out_5_)
  );
  and_ii _519_ (
    .a(_apc64_2_apc32_2_out_0_),
    .b(_apc64_2_apc32_1_out_0_),
    .c(_160_)
  );
  and_bi _520_ (
    .a(_130_),
    .b(_160_),
    .c(_apc64_2_out_0_)
  );
  maj_bbi _521_ (
    .a(_apc64_2_apc32_2_out_5_),
    .b(_apc64_2_apc32_1_out_5_),
    .c(_154_),
    .d(_apc64_2_out_6_)
  );
  or_ii _522_ (
    .a(1'b0),
    .b(1'b0),
    .c(_161_)
  );
  or_ii _523_ (
    .a(_apc64_2_apc32_1_apc16_2_half1_s ),
    .b(_apc64_2_apc32_1_apc16_1_half1_s ),
    .c(_162_)
  );
  and_ii _524_ (
    .a(_apc64_2_apc32_1_apc16_2_half1_s ),
    .b(_apc64_2_apc32_1_apc16_1_half1_s ),
    .c(_163_)
  );
  and_bi _525_ (
    .a(_162_),
    .b(_163_),
    .c(_164_)
  );
  or_bi _526_ (
    .a(_161_),
    .b(_164_),
    .c(_165_)
  );
  and_bi _527_ (
    .a(_161_),
    .b(_164_),
    .c(_166_)
  );
  and_bi _528_ (
    .a(_165_),
    .b(_166_),
    .c(_apc64_2_apc32_1_out_1_)
  );
  maj_bii _529_ (
    .a(_161_),
    .b(_apc64_2_apc32_1_apc16_2_half1_s ),
    .c(_apc64_2_apc32_1_apc16_1_half1_s ),
    .d(_167_)
  );
  or_ii _530_ (
    .a(_apc64_2_apc32_1_apc16_2_half2_s ),
    .b(_apc64_2_apc32_1_apc16_1_half2_s ),
    .c(_168_)
  );
  and_ii _531_ (
    .a(_apc64_2_apc32_1_apc16_2_half2_s ),
    .b(_apc64_2_apc32_1_apc16_1_half2_s ),
    .c(_169_)
  );
  and_bi _532_ (
    .a(_168_),
    .b(_169_),
    .c(_170_)
  );
  or_bi _533_ (
    .a(_167_),
    .b(_170_),
    .c(_171_)
  );
  and_bi _534_ (
    .a(_167_),
    .b(_170_),
    .c(_172_)
  );
  and_bi _535_ (
    .a(_171_),
    .b(_172_),
    .c(_apc64_2_apc32_1_out_2_)
  );
  maj_bii _536_ (
    .a(_167_),
    .b(_apc64_2_apc32_1_apc16_2_half2_s ),
    .c(_apc64_2_apc32_1_apc16_1_half2_s ),
    .d(_173_)
  );
  or_ii _537_ (
    .a(_apc64_2_apc32_1_apc16_2_half3_s ),
    .b(_apc64_2_apc32_1_apc16_1_half3_s ),
    .c(_174_)
  );
  and_ii _538_ (
    .a(_apc64_2_apc32_1_apc16_2_half3_s ),
    .b(_apc64_2_apc32_1_apc16_1_half3_s ),
    .c(_175_)
  );
  and_bi _539_ (
    .a(_174_),
    .b(_175_),
    .c(_176_)
  );
  or_bi _540_ (
    .a(_173_),
    .b(_176_),
    .c(_177_)
  );
  and_bi _541_ (
    .a(_173_),
    .b(_176_),
    .c(_178_)
  );
  and_bi _542_ (
    .a(_177_),
    .b(_178_),
    .c(_apc64_2_apc32_1_out_3_)
  );
  maj_bii _543_ (
    .a(_173_),
    .b(_apc64_2_apc32_1_apc16_2_half3_s ),
    .c(_apc64_2_apc32_1_apc16_1_half3_s ),
    .d(_179_)
  );
  or_ii _544_ (
    .a(_apc64_2_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_1_apc16_1_half3_cout ),
    .c(_180_)
  );
  and_ii _545_ (
    .a(_apc64_2_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_1_apc16_1_half3_cout ),
    .c(_181_)
  );
  and_bi _546_ (
    .a(_180_),
    .b(_181_),
    .c(_182_)
  );
  or_bi _547_ (
    .a(_179_),
    .b(_182_),
    .c(_183_)
  );
  and_bi _548_ (
    .a(_179_),
    .b(_182_),
    .c(_184_)
  );
  and_bi _549_ (
    .a(_183_),
    .b(_184_),
    .c(_apc64_2_apc32_1_out_4_)
  );
  and_ii _550_ (
    .a(1'b0),
    .b(1'b0),
    .c(_185_)
  );
  and_bi _551_ (
    .a(_161_),
    .b(_185_),
    .c(_apc64_2_apc32_1_out_0_)
  );
  maj_bbi _552_ (
    .a(_apc64_2_apc32_1_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_1_apc16_1_half3_cout ),
    .c(_179_),
    .d(_apc64_2_apc32_1_out_5_)
  );
  or_bb _553_ (
    .a(in_49_),
    .b(in_48_),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_a )
  );
  and_bb _554_ (
    .a(in_51_),
    .b(in_50_),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_b )
  );
  or_bb _555_ (
    .a(in_53_),
    .b(in_52_),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_cin )
  );
  and_bb _556_ (
    .a(in_55_),
    .b(in_54_),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv1_a )
  );
  or_bb _557_ (
    .a(in_57_),
    .b(in_56_),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv1_b )
  );
  and_bb _558_ (
    .a(in_59_),
    .b(in_58_),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv1_cin )
  );
  or_bb _559_ (
    .a(in_61_),
    .b(in_60_),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv2_cin )
  );
  and_bb _560_ (
    .a(in_63_),
    .b(in_62_),
    .c(_apc64_2_apc32_1_apc16_1_half1_a )
  );
  maj_bbb _561_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv1_cin ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv1_b ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_a ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _562_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv1_b ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv1_a ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_cin ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv1_d )
  );
  maj_bbi _563_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv1_d ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv1_cin ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _564_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv2_cin ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_b ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _565_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv2_b ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv1_cout ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv2_d )
  );
  maj_bbi _566_ (
    .a(_apc64_2_apc32_1_apc16_1_adder1_lv2_d ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_cin ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv2_cout ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _567_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv1_cin ),
    .b(_apc64_2_apc32_1_apc16_1_adder2_lv1_b ),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv1_a ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv2_b )
  );
  maj_bbi _568_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv1_b ),
    .b(_apc64_2_apc32_1_apc16_1_adder2_lv1_a ),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv1_cin ),
    .d(_apc64_2_apc32_1_apc16_1_adder2_lv1_d )
  );
  maj_bbi _569_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv1_d ),
    .b(_apc64_2_apc32_1_apc16_1_adder2_lv1_cin ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv2_b ),
    .d(_apc64_2_apc32_1_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _570_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv2_cin ),
    .b(_apc64_2_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .d(_apc64_2_apc32_1_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _571_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .c(_apc64_2_apc32_1_apc16_1_adder2_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_1_adder2_lv2_d )
  );
  maj_bbi _572_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv2_d ),
    .b(_apc64_2_apc32_1_apc16_1_adder2_lv2_cin ),
    .c(_apc64_2_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _573_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_1_apc16_1_half1_a ),
    .c(_apc64_2_apc32_1_apc16_1_half1_cout )
  );
  or_bb _574_ (
    .a(_apc64_2_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_1_apc16_1_half1_a ),
    .c(_186_)
  );
  and_bi _575_ (
    .a(_186_),
    .b(_apc64_2_apc32_1_apc16_1_half1_cout ),
    .c(_apc64_2_apc32_1_apc16_1_half1_s )
  );
  and_bb _576_ (
    .a(_apc64_2_apc32_1_apc16_1_half1_cout ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_apc64_2_apc32_1_apc16_1_half2_cout )
  );
  or_bb _577_ (
    .a(_apc64_2_apc32_1_apc16_1_half1_cout ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_187_)
  );
  and_bi _578_ (
    .a(_187_),
    .b(_apc64_2_apc32_1_apc16_1_half2_cout ),
    .c(_apc64_2_apc32_1_apc16_1_half2_s )
  );
  and_bb _579_ (
    .a(_apc64_2_apc32_1_apc16_1_half2_cout ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_apc64_2_apc32_1_apc16_1_half3_cout )
  );
  or_bb _580_ (
    .a(_apc64_2_apc32_1_apc16_1_half2_cout ),
    .b(_apc64_2_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_188_)
  );
  and_bi _581_ (
    .a(_188_),
    .b(_apc64_2_apc32_1_apc16_1_half3_cout ),
    .c(_apc64_2_apc32_1_apc16_1_half3_s )
  );
  or_bb _582_ (
    .a(in_33_),
    .b(in_32_),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_a )
  );
  and_bb _583_ (
    .a(in_35_),
    .b(in_34_),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_b )
  );
  or_bb _584_ (
    .a(in_37_),
    .b(in_36_),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_cin )
  );
  and_bb _585_ (
    .a(in_39_),
    .b(in_38_),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv1_a )
  );
  or_bb _586_ (
    .a(in_41_),
    .b(in_40_),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv1_b )
  );
  and_bb _587_ (
    .a(in_43_),
    .b(in_42_),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv1_cin )
  );
  or_bb _588_ (
    .a(in_45_),
    .b(in_44_),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv2_cin )
  );
  and_bb _589_ (
    .a(in_47_),
    .b(in_46_),
    .c(_apc64_2_apc32_1_apc16_2_half1_a )
  );
  maj_bbb _590_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv1_cin ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv1_b ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_a ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _591_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv1_b ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv1_a ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_cin ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv1_d )
  );
  maj_bbi _592_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv1_d ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv1_cin ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _593_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv2_cin ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_b ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _594_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv2_b ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv1_cout ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv2_d )
  );
  maj_bbi _595_ (
    .a(_apc64_2_apc32_1_apc16_2_adder1_lv2_d ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_cin ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv2_cout ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _596_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv1_cin ),
    .b(_apc64_2_apc32_1_apc16_2_adder2_lv1_b ),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv1_a ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv2_b )
  );
  maj_bbi _597_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv1_b ),
    .b(_apc64_2_apc32_1_apc16_2_adder2_lv1_a ),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv1_cin ),
    .d(_apc64_2_apc32_1_apc16_2_adder2_lv1_d )
  );
  maj_bbi _598_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv1_d ),
    .b(_apc64_2_apc32_1_apc16_2_adder2_lv1_cin ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv2_b ),
    .d(_apc64_2_apc32_1_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _599_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv2_cin ),
    .b(_apc64_2_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .d(_apc64_2_apc32_1_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _600_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .c(_apc64_2_apc32_1_apc16_2_adder2_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_2_adder2_lv2_d )
  );
  maj_bbi _601_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv2_d ),
    .b(_apc64_2_apc32_1_apc16_2_adder2_lv2_cin ),
    .c(_apc64_2_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc64_2_apc32_1_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _602_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_1_apc16_2_half1_a ),
    .c(_apc64_2_apc32_1_apc16_2_half1_cout )
  );
  or_bb _603_ (
    .a(_apc64_2_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_1_apc16_2_half1_a ),
    .c(_189_)
  );
  and_bi _604_ (
    .a(_189_),
    .b(_apc64_2_apc32_1_apc16_2_half1_cout ),
    .c(_apc64_2_apc32_1_apc16_2_half1_s )
  );
  and_bb _605_ (
    .a(_apc64_2_apc32_1_apc16_2_half1_cout ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_apc64_2_apc32_1_apc16_2_half2_cout )
  );
  or_bb _606_ (
    .a(_apc64_2_apc32_1_apc16_2_half1_cout ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_190_)
  );
  and_bi _607_ (
    .a(_190_),
    .b(_apc64_2_apc32_1_apc16_2_half2_cout ),
    .c(_apc64_2_apc32_1_apc16_2_half2_s )
  );
  and_bb _608_ (
    .a(_apc64_2_apc32_1_apc16_2_half2_cout ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_apc64_2_apc32_1_apc16_2_half3_cout )
  );
  or_bb _609_ (
    .a(_apc64_2_apc32_1_apc16_2_half2_cout ),
    .b(_apc64_2_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_191_)
  );
  and_bi _610_ (
    .a(_191_),
    .b(_apc64_2_apc32_1_apc16_2_half3_cout ),
    .c(_apc64_2_apc32_1_apc16_2_half3_s )
  );
  or_ii _611_ (
    .a(1'b0),
    .b(1'b0),
    .c(_192_)
  );
  or_ii _612_ (
    .a(_apc64_2_apc32_2_apc16_2_half1_s ),
    .b(_apc64_2_apc32_2_apc16_1_half1_s ),
    .c(_193_)
  );
  and_ii _613_ (
    .a(_apc64_2_apc32_2_apc16_2_half1_s ),
    .b(_apc64_2_apc32_2_apc16_1_half1_s ),
    .c(_194_)
  );
  and_bi _614_ (
    .a(_193_),
    .b(_194_),
    .c(_195_)
  );
  or_bi _615_ (
    .a(_192_),
    .b(_195_),
    .c(_196_)
  );
  and_bi _616_ (
    .a(_192_),
    .b(_195_),
    .c(_197_)
  );
  and_bi _617_ (
    .a(_196_),
    .b(_197_),
    .c(_apc64_2_apc32_2_out_1_)
  );
  maj_bii _618_ (
    .a(_192_),
    .b(_apc64_2_apc32_2_apc16_2_half1_s ),
    .c(_apc64_2_apc32_2_apc16_1_half1_s ),
    .d(_198_)
  );
  or_ii _619_ (
    .a(_apc64_2_apc32_2_apc16_2_half2_s ),
    .b(_apc64_2_apc32_2_apc16_1_half2_s ),
    .c(_199_)
  );
  and_ii _620_ (
    .a(_apc64_2_apc32_2_apc16_2_half2_s ),
    .b(_apc64_2_apc32_2_apc16_1_half2_s ),
    .c(_200_)
  );
  and_bi _621_ (
    .a(_199_),
    .b(_200_),
    .c(_201_)
  );
  or_bi _622_ (
    .a(_198_),
    .b(_201_),
    .c(_202_)
  );
  and_bi _623_ (
    .a(_198_),
    .b(_201_),
    .c(_203_)
  );
  and_bi _624_ (
    .a(_202_),
    .b(_203_),
    .c(_apc64_2_apc32_2_out_2_)
  );
  maj_bii _625_ (
    .a(_198_),
    .b(_apc64_2_apc32_2_apc16_2_half2_s ),
    .c(_apc64_2_apc32_2_apc16_1_half2_s ),
    .d(_204_)
  );
  or_ii _626_ (
    .a(_apc64_2_apc32_2_apc16_2_half3_s ),
    .b(_apc64_2_apc32_2_apc16_1_half3_s ),
    .c(_205_)
  );
  and_ii _627_ (
    .a(_apc64_2_apc32_2_apc16_2_half3_s ),
    .b(_apc64_2_apc32_2_apc16_1_half3_s ),
    .c(_206_)
  );
  and_bi _628_ (
    .a(_205_),
    .b(_206_),
    .c(_207_)
  );
  or_bi _629_ (
    .a(_204_),
    .b(_207_),
    .c(_208_)
  );
  and_bi _630_ (
    .a(_204_),
    .b(_207_),
    .c(_209_)
  );
  and_bi _631_ (
    .a(_208_),
    .b(_209_),
    .c(_apc64_2_apc32_2_out_3_)
  );
  maj_bii _632_ (
    .a(_204_),
    .b(_apc64_2_apc32_2_apc16_2_half3_s ),
    .c(_apc64_2_apc32_2_apc16_1_half3_s ),
    .d(_210_)
  );
  or_ii _633_ (
    .a(_apc64_2_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_2_apc16_1_half3_cout ),
    .c(_211_)
  );
  and_ii _634_ (
    .a(_apc64_2_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_2_apc16_1_half3_cout ),
    .c(_212_)
  );
  and_bi _635_ (
    .a(_211_),
    .b(_212_),
    .c(_213_)
  );
  or_bi _636_ (
    .a(_210_),
    .b(_213_),
    .c(_214_)
  );
  and_bi _637_ (
    .a(_210_),
    .b(_213_),
    .c(_215_)
  );
  and_bi _638_ (
    .a(_214_),
    .b(_215_),
    .c(_apc64_2_apc32_2_out_4_)
  );
  and_ii _639_ (
    .a(1'b0),
    .b(1'b0),
    .c(_216_)
  );
  and_bi _640_ (
    .a(_192_),
    .b(_216_),
    .c(_apc64_2_apc32_2_out_0_)
  );
  maj_bbi _641_ (
    .a(_apc64_2_apc32_2_apc16_2_half3_cout ),
    .b(_apc64_2_apc32_2_apc16_1_half3_cout ),
    .c(_210_),
    .d(_apc64_2_apc32_2_out_5_)
  );
  or_bb _642_ (
    .a(in_17_),
    .b(in_16_),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_a )
  );
  and_bb _643_ (
    .a(in_19_),
    .b(in_18_),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_b )
  );
  or_bb _644_ (
    .a(in_21_),
    .b(in_20_),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_cin )
  );
  and_bb _645_ (
    .a(in_23_),
    .b(in_22_),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv1_a )
  );
  or_bb _646_ (
    .a(in_25_),
    .b(in_24_),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv1_b )
  );
  and_bb _647_ (
    .a(in_27_),
    .b(in_26_),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv1_cin )
  );
  or_bb _648_ (
    .a(in_29_),
    .b(in_28_),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv2_cin )
  );
  and_bb _649_ (
    .a(in_31_),
    .b(in_30_),
    .c(_apc64_2_apc32_2_apc16_1_half1_a )
  );
  maj_bbb _650_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv1_cin ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv1_b ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_a ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _651_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv1_b ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv1_a ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_cin ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv1_d )
  );
  maj_bbi _652_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv1_d ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv1_cin ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _653_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv2_cin ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_b ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _654_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv2_b ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv1_cout ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv2_d )
  );
  maj_bbi _655_ (
    .a(_apc64_2_apc32_2_apc16_1_adder1_lv2_d ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_cin ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv2_cout ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _656_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv1_cin ),
    .b(_apc64_2_apc32_2_apc16_1_adder2_lv1_b ),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv1_a ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv2_b )
  );
  maj_bbi _657_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv1_b ),
    .b(_apc64_2_apc32_2_apc16_1_adder2_lv1_a ),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv1_cin ),
    .d(_apc64_2_apc32_2_apc16_1_adder2_lv1_d )
  );
  maj_bbi _658_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv1_d ),
    .b(_apc64_2_apc32_2_apc16_1_adder2_lv1_cin ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv2_b ),
    .d(_apc64_2_apc32_2_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _659_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv2_cin ),
    .b(_apc64_2_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .d(_apc64_2_apc32_2_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _660_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .c(_apc64_2_apc32_2_apc16_1_adder2_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_1_adder2_lv2_d )
  );
  maj_bbi _661_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv2_d ),
    .b(_apc64_2_apc32_2_apc16_1_adder2_lv2_cin ),
    .c(_apc64_2_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _662_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_2_apc16_1_half1_a ),
    .c(_apc64_2_apc32_2_apc16_1_half1_cout )
  );
  or_bb _663_ (
    .a(_apc64_2_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_2_apc16_1_half1_a ),
    .c(_217_)
  );
  and_bi _664_ (
    .a(_217_),
    .b(_apc64_2_apc32_2_apc16_1_half1_cout ),
    .c(_apc64_2_apc32_2_apc16_1_half1_s )
  );
  and_bb _665_ (
    .a(_apc64_2_apc32_2_apc16_1_half1_cout ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_apc64_2_apc32_2_apc16_1_half2_cout )
  );
  or_bb _666_ (
    .a(_apc64_2_apc32_2_apc16_1_half1_cout ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_218_)
  );
  and_bi _667_ (
    .a(_218_),
    .b(_apc64_2_apc32_2_apc16_1_half2_cout ),
    .c(_apc64_2_apc32_2_apc16_1_half2_s )
  );
  and_bb _668_ (
    .a(_apc64_2_apc32_2_apc16_1_half2_cout ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_apc64_2_apc32_2_apc16_1_half3_cout )
  );
  or_bb _669_ (
    .a(_apc64_2_apc32_2_apc16_1_half2_cout ),
    .b(_apc64_2_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_219_)
  );
  and_bi _670_ (
    .a(_219_),
    .b(_apc64_2_apc32_2_apc16_1_half3_cout ),
    .c(_apc64_2_apc32_2_apc16_1_half3_s )
  );
  or_bb _671_ (
    .a(in_1_),
    .b(in_0_),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_a )
  );
  and_bb _672_ (
    .a(in_3_),
    .b(in_2_),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_b )
  );
  or_bb _673_ (
    .a(in_5_),
    .b(in_4_),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_cin )
  );
  and_bb _674_ (
    .a(in_7_),
    .b(in_6_),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv1_a )
  );
  or_bb _675_ (
    .a(in_9_),
    .b(in_8_),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv1_b )
  );
  and_bb _676_ (
    .a(in_11_),
    .b(in_10_),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv1_cin )
  );
  or_bb _677_ (
    .a(in_13_),
    .b(in_12_),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv2_cin )
  );
  and_bb _678_ (
    .a(in_15_),
    .b(in_14_),
    .c(_apc64_2_apc32_2_apc16_2_half1_a )
  );
  maj_bbb _679_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv1_cin ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv1_b ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_a ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _680_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv1_b ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv1_a ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_cin ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv1_d )
  );
  maj_bbi _681_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv1_d ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv1_cin ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _682_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv2_cin ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_b ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _683_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv2_b ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv1_cout ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv2_d )
  );
  maj_bbi _684_ (
    .a(_apc64_2_apc32_2_apc16_2_adder1_lv2_d ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_cin ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv2_cout ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _685_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv1_cin ),
    .b(_apc64_2_apc32_2_apc16_2_adder2_lv1_b ),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv1_a ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv2_b )
  );
  maj_bbi _686_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv1_b ),
    .b(_apc64_2_apc32_2_apc16_2_adder2_lv1_a ),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv1_cin ),
    .d(_apc64_2_apc32_2_apc16_2_adder2_lv1_d )
  );
  maj_bbi _687_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv1_d ),
    .b(_apc64_2_apc32_2_apc16_2_adder2_lv1_cin ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv2_b ),
    .d(_apc64_2_apc32_2_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _688_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv2_cin ),
    .b(_apc64_2_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .d(_apc64_2_apc32_2_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _689_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .c(_apc64_2_apc32_2_apc16_2_adder2_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_2_adder2_lv2_d )
  );
  maj_bbi _690_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv2_d ),
    .b(_apc64_2_apc32_2_apc16_2_adder2_lv2_cin ),
    .c(_apc64_2_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc64_2_apc32_2_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _691_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_2_apc16_2_half1_a ),
    .c(_apc64_2_apc32_2_apc16_2_half1_cout )
  );
  or_bb _692_ (
    .a(_apc64_2_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc64_2_apc32_2_apc16_2_half1_a ),
    .c(_220_)
  );
  and_bi _693_ (
    .a(_220_),
    .b(_apc64_2_apc32_2_apc16_2_half1_cout ),
    .c(_apc64_2_apc32_2_apc16_2_half1_s )
  );
  and_bb _694_ (
    .a(_apc64_2_apc32_2_apc16_2_half1_cout ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_apc64_2_apc32_2_apc16_2_half2_cout )
  );
  or_bb _695_ (
    .a(_apc64_2_apc32_2_apc16_2_half1_cout ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_221_)
  );
  and_bi _696_ (
    .a(_221_),
    .b(_apc64_2_apc32_2_apc16_2_half2_cout ),
    .c(_apc64_2_apc32_2_apc16_2_half2_s )
  );
  and_bb _697_ (
    .a(_apc64_2_apc32_2_apc16_2_half2_cout ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_apc64_2_apc32_2_apc16_2_half3_cout )
  );
  or_bb _698_ (
    .a(_apc64_2_apc32_2_apc16_2_half2_cout ),
    .b(_apc64_2_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_222_)
  );
  and_bi _699_ (
    .a(_222_),
    .b(_apc64_2_apc32_2_apc16_2_half3_cout ),
    .c(_apc64_2_apc32_2_apc16_2_half3_s )
  );
endmodule
