module c6288(N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528, N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288);
	wire new_net_1720;
	wire new_net_20316;
	wire new_net_2272;
	wire new_net_5105;
	wire new_net_5250;
	wire new_net_9846;
	wire new_net_8109;
	wire new_net_19832;
	wire new_net_20464;
	wire _1106_;
	wire new_net_1867;
	wire new_net_12198;
	wire new_net_12434;
	wire new_net_13769;
	wire new_net_12885;
	wire new_net_14016;
	wire new_net_17696;
	wire new_net_16857;
	wire new_net_4638;
	wire new_net_4;
	wire new_net_2278;
	wire new_net_4927;
	wire new_net_5787;
	wire new_net_8445;
	wire new_net_18146;
	wire new_net_798;
	wire new_net_14479;
	wire new_net_3567;
	wire _1107_;
	wire new_net_2162;
	wire new_net_3667;
	wire new_net_7681;
	wire new_net_9849;
	wire new_net_4111;
	wire new_net_21313;
	wire new_net_18782;
	wire new_net_12;
	wire new_net_103;
	wire new_net_3458;
	wire new_net_5790;
	wire new_net_9848;
	wire new_net_7848;
	wire new_net_9288;
	wire new_net_19285;
	wire _1108_;
	wire new_net_3672;
	wire new_net_4106;
	wire new_net_15283;
	wire new_net_17778;
	wire new_net_20739;
	wire new_net_1647;
	wire new_net_3454;
	wire new_net_7115;
	wire new_net_8916;
	wire new_net_16228;
	wire new_net_11134;
	wire new_net_15970;
	wire new_net_7851;
	wire new_net_9291;
	wire new_net_21286;
	wire new_net_17949;
	wire new_net_105;
	wire _1109_;
	wire new_net_7321;
	wire new_net_10612;
	wire new_net_4640;
	wire new_net_19458;
	wire new_net_19833;
	wire new_net_20465;
	wire new_net_16064;
	wire new_net_1636;
	wire new_net_7114;
	wire new_net_12199;
	wire new_net_12435;
	wire new_net_13770;
	wire new_net_17281;
	wire new_net_12886;
	wire new_net_14017;
	wire new_net_17697;
	wire new_net_16858;
	wire _1110_;
	wire new_net_11;
	wire new_net_695;
	wire new_net_2799;
	wire new_net_8908;
	wire new_net_18144;
	wire new_net_20905;
	wire new_net_14;
	wire new_net_8904;
	wire new_net_9295;
	wire new_net_16466;
	wire new_net_21314;
	wire _1111_;
	wire new_net_3826;
	wire new_net_7312;
	wire new_net_14819;
	wire new_net_19500;
	wire new_net_21320;
	wire new_net_2034;
	wire new_net_19034;
	wire new_net_4107;
	wire new_net_7539;
	wire new_net_8914;
	wire new_net_9406;
	wire new_net_20740;
	wire _1112_;
	wire new_net_4637;
	wire new_net_4851;
	wire new_net_8909;
	wire new_net_15282;
	wire new_net_17777;
	wire new_net_7678;
	wire new_net_11135;
	wire new_net_16458;
	wire new_net_9173;
	wire new_net_697;
	wire new_net_4928;
	wire new_net_7195;
	wire new_net_7849;
	wire new_net_7865;
	wire new_net_19834;
	wire new_net_20466;
	wire new_net_100;
	wire new_net_696;
	wire _1113_;
	wire new_net_7536;
	wire new_net_7543;
	wire new_net_8907;
	wire new_net_12200;
	wire new_net_12436;
	wire new_net_13771;
	wire new_net_1644;
	wire _1582_;
	wire new_net_7311;
	wire new_net_17279;
	wire new_net_16227;
	wire new_net_9411;
	wire new_net_15969;
	wire new_net_20354;
	wire new_net_3537;
	wire new_net_13548;
	wire _1114_;
	wire new_net_6;
	wire new_net_688;
	wire new_net_16455;
	wire new_net_18138;
	wire new_net_21315;
	wire new_net_17309;
	wire new_net_19099;
	wire new_net_18564;
	wire new_net_9178;
	wire new_net_2644;
	wire new_net_104;
	wire new_net_5256;
	wire new_net_10300;
	wire new_net_19237;
	wire new_net_19053;
	wire _1115_;
	wire new_net_7541;
	wire new_net_7112;
	wire new_net_9852;
	wire new_net_8104;
	wire new_net_7852;
	wire new_net_10113;
	wire new_net_20353;
	wire new_net_20741;
	wire new_net_21188;
	wire new_net_6282;
	wire new_net_2277;
	wire new_net_4105;
	wire new_net_4859;
	wire new_net_5107;
	wire new_net_15281;
	wire new_net_5258;
	wire new_net_11136;
	wire new_net_9845;
	wire new_net_2525;
	wire _1116_;
	wire new_net_5970;
	wire new_net_7871;
	wire new_net_19242;
	wire new_net_13132;
	wire new_net_19835;
	wire new_net_20467;
	wire new_net_5685;
	wire new_net_1864;
	wire new_net_2276;
	wire new_net_4061;
	wire new_net_7117;
	wire new_net_14617;
	wire new_net_12201;
	wire new_net_12437;
	wire new_net_13772;
	wire new_net_8918;
	wire new_net_12888;
	wire new_net_19511;
	wire _1117_;
	wire new_net_2643;
	wire new_net_5793;
	wire new_net_8917;
	wire new_net_16226;
	wire new_net_15968;
	wire new_net_10114;
	wire new_net_691;
	wire new_net_4108;
	wire new_net_5792;
	wire new_net_8671;
	wire new_net_17776;
	wire new_net_10607;
	wire new_net_9294;
	wire new_net_16465;
	wire new_net_19286;
	wire new_net_20352;
	wire _1118_;
	wire new_net_2159;
	wire new_net_9179;
	wire new_net_7676;
	wire new_net_4065;
	wire new_net_18143;
	wire new_net_19287;
	wire new_net_19451;
	wire new_net_17759;
	wire new_net_3828;
	wire new_net_4066;
	wire new_net_4068;
	wire new_net_7868;
	wire new_net_9176;
	wire new_net_8164;
	wire new_net_10609;
	wire new_net_8113;
	wire new_net_10299;
	wire new_net_20742;
	wire _1119_;
	wire new_net_3459;
	wire new_net_3671;
	wire new_net_7194;
	wire new_net_9175;
	wire new_net_17278;
	wire new_net_17775;
	wire new_net_11137;
	wire new_net_18153;
	wire new_net_3824;
	wire new_net_7320;
	wire new_net_9405;
	wire new_net_9287;
	wire new_net_19288;
	wire new_net_19836;
	wire new_net_20468;
	wire new_net_12711;
	wire new_net_17700;
	wire _1120_;
	wire new_net_4860;
	wire new_net_14618;
	wire new_net_12048;
	wire new_net_13773;
	wire new_net_12202;
	wire new_net_12438;
	wire new_net_7679;
	wire _0133_;
	wire new_net_16225;
	wire new_net_2275;
	wire new_net_1639;
	wire new_net_1872;
	wire new_net_4063;
	wire new_net_4104;
	wire new_net_7113;
	wire new_net_9404;
	wire new_net_10611;
	wire new_net_8912;
	wire new_net_13641;
	wire _1121_;
	wire new_net_5791;
	wire new_net_9734;
	wire new_net_16459;
	wire new_net_7866;
	wire new_net_7530;
	wire new_net_8451;
	wire new_net_21317;
	wire new_net_18601;
	wire new_net_2797;
	wire new_net_3918;
	wire new_net_7850;
	wire new_net_9739;
	wire new_net_10295;
	wire new_net_19061;
	wire new_net_19203;
	wire _1122_;
	wire new_net_1634;
	wire new_net_1869;
	wire new_net_2641;
	wire new_net_4852;
	wire new_net_20743;
	wire new_net_21190;
	wire new_net_7;
	wire new_net_4853;
	wire new_net_17277;
	wire new_net_11138;
	wire new_net_17173;
	wire _1123_;
	wire new_net_7684;
	wire new_net_10605;
	wire new_net_9412;
	wire new_net_19457;
	wire new_net_19837;
	wire new_net_20469;
	wire new_net_5794;
	wire new_net_9292;
	wire new_net_12049;
	wire new_net_12712;
	wire new_net_3668;
	wire new_net_4109;
	wire new_net_14619;
	wire new_net_12203;
	wire new_net_12439;
	wire new_net_13774;
	wire new_net_5789;
	wire _1124_;
	wire new_net_1637;
	wire new_net_1866;
	wire new_net_15278;
	wire new_net_16224;
	wire new_net_15966;
	wire new_net_16464;
	wire new_net_1640;
	wire new_net_3457;
	wire new_net_3827;
	wire new_net_7314;
	wire new_net_9174;
	wire new_net_9851;
	wire new_net_18142;
	wire new_net_21318;
	wire new_net_7847;
	wire new_net_8452;
	wire _1125_;
	wire new_net_7317;
	wire new_net_10298;
	wire new_net_692;
	wire new_net_2161;
	wire new_net_7853;
	wire new_net_8910;
	wire new_net_9403;
	wire new_net_19491;
	wire new_net_20345;
	wire new_net_20744;
	wire new_net_21191;
	wire new_net_20227;
	wire new_net_101;
	wire _1126_;
	wire new_net_2639;
	wire new_net_4062;
	wire new_net_4929;
	wire new_net_3670;
	wire new_net_11139;
	wire new_net_17950;
	wire new_net_10;
	wire new_net_2279;
	wire new_net_3456;
	wire new_net_4636;
	wire new_net_9733;
	wire new_net_7109;
	wire new_net_9853;
	wire new_net_18135;
	wire new_net_19838;
	wire new_net_20470;
	wire _1127_;
	wire new_net_2798;
	wire new_net_5254;
	wire new_net_17478;
	wire new_net_5796;
	wire new_net_16863;
	wire new_net_12891;
	wire new_net_9290;
	wire new_net_12204;
	wire new_net_12440;
	wire new_net_7111;
	wire new_net_7537;
	wire new_net_8163;
	wire new_net_10301;
	wire new_net_8906;
	wire new_net_17772;
	wire new_net_16223;
	wire new_net_9407;
	wire new_net_15965;
	wire new_net_19498;
	wire _1128_;
	wire new_net_2642;
	wire new_net_3663;
	wire new_net_5795;
	wire new_net_8673;
	wire new_net_7542;
	wire new_net_12056;
	wire new_net_18141;
	wire new_net_18853;
	wire new_net_20351;
	wire new_net_3665;
	wire new_net_7193;
	wire new_net_21321;
	wire new_net_19035;
	wire _1129_;
	wire new_net_16456;
	wire new_net_2160;
	wire new_net_4067;
	wire new_net_9844;
	wire new_net_19492;
	wire new_net_20745;
	wire new_net_21192;
	wire new_net_19510;
	wire new_net_8;
	wire new_net_3460;
	wire new_net_7192;
	wire new_net_9738;
	wire new_net_15277;
	wire new_net_7313;
	wire new_net_11140;
	wire new_net_9409;
	wire new_net_18140;
	wire _1130_;
	wire new_net_7190;
	wire new_net_4926;
	wire new_net_4858;
	wire new_net_9850;
	wire new_net_19839;
	wire new_net_20471;
	wire new_net_16722;
	wire new_net_693;
	wire new_net_9296;
	wire new_net_12051;
	wire new_net_7191;
	wire new_net_14621;
	wire new_net_12205;
	wire new_net_12441;
	wire new_net_12892;
	wire new_net_17275;
	wire new_net_5563;
	wire _1131_;
	wire new_net_4110;
	wire new_net_4855;
	wire new_net_9735;
	wire new_net_15964;
	wire new_net_12050;
	wire new_net_17271;
	wire new_net_16222;
	wire new_net_4243;
	wire new_net_8112;
	wire new_net_13;
	wire new_net_3666;
	wire new_net_4633;
	wire new_net_4930;
	wire new_net_5106;
	wire new_net_16463;
	wire new_net_7677;
	wire new_net_5251;
	wire new_net_9181;
	wire new_net_19100;
	wire _1132_;
	wire new_net_4639;
	wire new_net_19243;
	wire new_net_18565;
	wire new_net_19054;
	wire new_net_10294;
	wire new_net_19497;
	wire new_net_20350;
	wire new_net_20746;
	wire new_net_21193;
	wire _1133_;
	wire new_net_1638;
	wire new_net_1868;
	wire new_net_2157;
	wire new_net_7873;
	wire new_net_15276;
	wire new_net_3825;
	wire new_net_11141;
	wire new_net_9847;
	wire new_net_17479;
	wire new_net_1643;
	wire new_net_3664;
	wire new_net_3829;
	wire new_net_8672;
	wire new_net_9732;
	wire new_net_10608;
	wire new_net_19244;
	wire new_net_19289;
	wire new_net_19840;
	wire new_net_20472;
	wire _0063_;
	wire new_net_16723;
	wire _1134_;
	wire new_net_2273;
	wire new_net_8450;
	wire new_net_12052;
	wire new_net_12715;
	wire new_net_14622;
	wire new_net_12206;
	wire new_net_12442;
	wire new_net_13777;
	wire new_net_15963;
	wire new_net_2795;
	wire new_net_5257;
	wire new_net_9289;
	wire new_net_9731;
	wire new_net_16221;
	wire new_net_20344;
	wire new_net_8111;
	wire new_net_2155;
	wire _1135_;
	wire new_net_694;
	wire new_net_5786;
	wire new_net_8453;
	wire new_net_7322;
	wire new_net_18139;
	wire new_net_19290;
	wire new_net_19456;
	wire new_net_4931;
	wire new_net_19638;
	wire new_net_1648;
	wire _1136_;
	wire new_net_3;
	wire new_net_10302;
	wire new_net_7680;
	wire new_net_19245;
	wire new_net_19496;
	wire new_net_20349;
	wire new_net_20747;
	wire new_net_21194;
	wire new_net_1870;
	wire new_net_1;
	wire new_net_4635;
	wire new_net_11142;
	wire new_net_9410;
	wire new_net_18154;
	wire _1137_;
	wire new_net_1646;
	wire new_net_1865;
	wire new_net_7854;
	wire new_net_9180;
	wire new_net_7116;
	wire new_net_19841;
	wire new_net_20473;
	wire new_net_7538;
	wire new_net_9177;
	wire new_net_16724;
	wire new_net_12053;
	wire new_net_12716;
	wire new_net_14623;
	wire new_net_12207;
	wire new_net_12443;
	wire new_net_13778;
	wire new_net_15275;
	wire _1138_;
	wire new_net_1645;
	wire new_net_2156;
	wire new_net_15962;
	wire new_net_16460;
	wire new_net_7683;
	wire new_net_16220;
	wire new_net_3946;
	wire new_net_8106;
	wire new_net_9297;
	wire new_net_16462;
	wire new_net_438;
	wire new_net_19455;
	wire new_net_21322;
	wire _1139_;
	wire new_net_10112;
	wire new_net_3669;
	wire new_net_8161;
	wire new_net_7319;
	wire new_net_18602;
	wire new_net_20370;
	wire new_net_19062;
	wire new_net_5;
	wire new_net_5969;
	wire new_net_20748;
	wire new_net_21195;
	wire new_net_19204;
	wire new_net_2;
	wire new_net_689;
	wire new_net_2282;
	wire _1140_;
	wire new_net_1642;
	wire new_net_2163;
	wire new_net_10610;
	wire new_net_11143;
	wire new_net_14275;
	wire new_net_4923;
	wire new_net_698;
	wire new_net_8905;
	wire new_net_19842;
	wire new_net_20474;
	wire new_net_18854;
	wire new_net_16844;
	wire new_net_17481;
	wire _1141_;
	wire new_net_1635;
	wire new_net_16725;
	wire new_net_12054;
	wire new_net_12717;
	wire new_net_16457;
	wire new_net_7869;
	wire new_net_14624;
	wire new_net_2281;
	wire new_net_4634;
	wire new_net_5253;
	wire new_net_15961;
	wire new_net_7189;
	wire new_net_7540;
	wire new_net_15273;
	wire new_net_16219;
	wire new_net_18137;
	wire new_net_1663;
	wire new_net_14481;
	wire new_net_4857;
	wire _1142_;
	wire new_net_8110;
	wire new_net_4064;
	wire new_net_8447;
	wire new_net_9298;
	wire new_net_10293;
	wire new_net_9736;
	wire new_net_5252;
	wire new_net_7110;
	wire new_net_102;
	wire new_net_2158;
	wire new_net_3830;
	wire new_net_8107;
	wire new_net_9293;
	wire new_net_10297;
	wire new_net_7196;
	wire new_net_16250;
	wire new_net_4854;
	wire new_net_9408;
	wire _1143_;
	wire new_net_2796;
	wire new_net_5564;
	wire new_net_15959;
	wire new_net_4112;
	wire new_net_7845;
	wire new_net_8449;
	wire new_net_16217;
	wire new_net_2274;
	wire new_net_4856;
	wire new_net_5968;
	wire new_net_10296;
	wire new_net_7864;
	wire new_net_8911;
	wire new_net_11144;
	wire new_net_19453;
	wire _1144_;
	wire new_net_8915;
	wire new_net_19494;
	wire new_net_19843;
	wire new_net_20347;
	wire new_net_20475;
	wire new_net_17951;
	wire new_net_20008;
	wire new_net_16845;
	wire new_net_17482;
	wire new_net_2640;
	wire new_net_7870;
	wire new_net_16726;
	wire new_net_12055;
	wire new_net_12718;
	wire new_net_14625;
	wire new_net_8913;
	wire new_net_12209;
	wire _1145_;
	wire new_net_1641;
	wire new_net_15960;
	wire new_net_10111;
	wire new_net_9737;
	wire new_net_8921;
	wire new_net_10613;
	wire new_net_16218;
	wire new_net_16461;
	wire new_net_17270;
	wire new_net_17767;
	wire new_net_21324;
	wire new_net_18852;
	wire new_net_690;
	wire _1146_;
	wire new_net_1871;
	wire new_net_3823;
	wire new_net_5249;
	wire new_net_19493;
	wire new_net_20346;
	wire new_net_12166;
	wire new_net_19036;
	wire new_net_2280;
	wire new_net_9;
	wire new_net_4924;
	wire new_net_5785;
	wire new_net_7846;
	wire new_net_8162;
	wire new_net_15272;
	wire new_net_8920;
	wire new_net_20750;
	wire new_net_21197;
	wire _1147_;
	wire new_net_7118;
	wire new_net_11145;
	wire new_net_5394;
	wire new_net_1365;
	wire new_net_1606;
	wire new_net_3865;
	wire new_net_9905;
	wire new_net_5870;
	wire new_net_9391;
	wire new_net_6945;
	wire new_net_14757;
	wire new_net_21462;
	wire _1589_;
	wire _1232_;
	wire _1064_;
	wire new_net_1406;
	wire new_net_12778;
	wire new_net_11880;
	wire new_net_12479;
	wire new_net_16372;
	wire new_net_10009;
	wire new_net_10710;
	wire new_net_14685;
	wire new_net_10147;
	wire new_net_19101;
	wire _1233_;
	wire new_net_1326;
	wire _1065_;
	wire new_net_1438;
	wire new_net_6407;
	wire new_net_10709;
	wire new_net_3860;
	wire new_net_9385;
	wire new_net_14756;
	wire new_net_8795;
	wire new_net_18566;
	wire new_net_3007;
	wire new_net_6411;
	wire new_net_19646;
	wire new_net_20906;
	wire new_net_6284;
	wire _1234_;
	wire new_net_1940;
	wire new_net_4602;
	wire new_net_5321;
	wire _1066_;
	wire new_net_5521;
	wire new_net_8280;
	wire new_net_1364;
	wire new_net_19527;
	wire new_net_20833;
	wire new_net_10850;
	wire new_net_227;
	wire new_net_1428;
	wire new_net_12480;
	wire new_net_10957;
	wire new_net_8802;
	wire new_net_5748;
	wire new_net_8299;
	wire new_net_5688;
	wire _1235_;
	wire _1067_;
	wire new_net_10703;
	wire new_net_10141;
	wire new_net_11724;
	wire new_net_3438;
	wire new_net_11881;
	wire new_net_12478;
	wire new_net_13004;
	wire new_net_9937;
	wire new_net_14158;
	wire new_net_16373;
	wire new_net_12779;
	wire new_net_13463;
	wire new_net_10144;
	wire _1236_;
	wire new_net_228;
	wire _1068_;
	wire new_net_1437;
	wire new_net_9075;
	wire new_net_6787;
	wire new_net_15666;
	wire new_net_8797;
	wire new_net_8302;
	wire new_net_20832;
	wire _1237_;
	wire _1069_;
	wire new_net_9073;
	wire new_net_9902;
	wire new_net_6409;
	wire new_net_15674;
	wire new_net_5747;
	wire new_net_18300;
	wire new_net_20824;
	wire new_net_621;
	wire new_net_5871;
	wire new_net_6939;
	wire new_net_19528;
	wire new_net_20907;
	wire new_net_18155;
	wire new_net_10851;
	wire _1238_;
	wire new_net_3001;
	wire _1070_;
	wire new_net_6402;
	wire new_net_9021;
	wire new_net_10958;
	wire new_net_14758;
	wire new_net_5517;
	wire new_net_6935;
	wire new_net_9386;
	wire new_net_10707;
	wire new_net_15663;
	wire new_net_19272;
	wire _1239_;
	wire new_net_224;
	wire new_net_11882;
	wire new_net_12477;
	wire new_net_13005;
	wire new_net_14159;
	wire new_net_16374;
	wire new_net_12780;
	wire new_net_6780;
	wire new_net_13464;
	wire new_net_225;
	wire new_net_1409;
	wire new_net_5319;
	wire new_net_13810;
	wire new_net_18603;
	wire new_net_8301;
	wire new_net_5400;
	wire new_net_1601;
	wire _1240_;
	wire new_net_2284;
	wire _1072_;
	wire new_net_15673;
	wire new_net_18299;
	wire new_net_20371;
	wire new_net_19063;
	wire new_net_9272;
	wire new_net_10525;
	wire new_net_2289;
	wire new_net_3005;
	wire new_net_1608;
	wire new_net_8801;
	wire new_net_19205;
	wire new_net_1357;
	wire new_net_1433;
	wire new_net_1605;
	wire _1241_;
	wire new_net_2286;
	wire new_net_6403;
	wire new_net_9019;
	wire _1073_;
	wire new_net_8803;
	wire new_net_19529;
	wire new_net_1408;
	wire new_net_2290;
	wire new_net_5671;
	wire new_net_10852;
	wire new_net_10959;
	wire new_net_5875;
	wire new_net_14759;
	wire _1074_;
	wire new_net_1354;
	wire new_net_1602;
	wire _1242_;
	wire new_net_231;
	wire new_net_6423;
	wire new_net_6779;
	wire new_net_19319;
	wire new_net_1607;
	wire new_net_1435;
	wire new_net_9072;
	wire new_net_11883;
	wire new_net_12476;
	wire new_net_13006;
	wire new_net_14160;
	wire new_net_16375;
	wire new_net_12781;
	wire new_net_13465;
	wire new_net_793;
	wire new_net_14482;
	wire new_net_6537;
	wire _1075_;
	wire _1243_;
	wire new_net_229;
	wire new_net_10528;
	wire new_net_5515;
	wire new_net_3323;
	wire new_net_5668;
	wire new_net_5756;
	wire new_net_9017;
	wire _1076_;
	wire new_net_4597;
	wire new_net_3862;
	wire _1244_;
	wire new_net_8284;
	wire new_net_1603;
	wire new_net_2997;
	wire new_net_9074;
	wire new_net_6784;
	wire new_net_8281;
	wire new_net_19530;
	wire new_net_20909;
	wire _1077_;
	wire _1245_;
	wire new_net_5397;
	wire new_net_10853;
	wire new_net_9933;
	wire new_net_10960;
	wire new_net_15671;
	wire new_net_14760;
	wire new_net_17952;
	wire new_net_18297;
	wire new_net_2303;
	wire new_net_6546;
	wire new_net_8304;
	wire new_net_1411;
	wire new_net_2285;
	wire new_net_9079;
	wire new_net_9934;
	wire new_net_5669;
	wire new_net_9388;
	wire new_net_6944;
	wire new_net_19316;
	wire new_net_1361;
	wire _1078_;
	wire _1246_;
	wire new_net_1325;
	wire new_net_2287;
	wire new_net_16376;
	wire new_net_9903;
	wire new_net_11884;
	wire new_net_12475;
	wire new_net_13007;
	wire new_net_13675;
	wire new_net_1436;
	wire new_net_6642;
	wire new_net_9078;
	wire new_net_10015;
	wire new_net_5869;
	wire new_net_18851;
	wire new_net_18319;
	wire _1079_;
	wire new_net_1412;
	wire new_net_10711;
	wire new_net_1943;
	wire _1247_;
	wire new_net_8800;
	wire new_net_20831;
	wire new_net_21323;
	wire new_net_19037;
	wire new_net_1434;
	wire new_net_1356;
	wire new_net_10706;
	wire new_net_6785;
	wire new_net_15672;
	wire new_net_10138;
	wire new_net_8287;
	wire new_net_18298;
	wire new_net_19693;
	wire _1248_;
	wire new_net_232;
	wire new_net_3000;
	wire new_net_5398;
	wire new_net_9938;
	wire new_net_10011;
	wire _1080_;
	wire new_net_6936;
	wire new_net_19531;
	wire new_net_20910;
	wire new_net_8285;
	wire new_net_6539;
	wire new_net_2293;
	wire new_net_10854;
	wire new_net_9910;
	wire new_net_9020;
	wire new_net_10013;
	wire new_net_10961;
	wire new_net_14761;
	wire new_net_19273;
	wire new_net_6540;
	wire _1249_;
	wire new_net_1611;
	wire _1081_;
	wire new_net_9906;
	wire new_net_9932;
	wire new_net_12262;
	wire new_net_14690;
	wire new_net_2283;
	wire new_net_5757;
	wire new_net_6545;
	wire new_net_6938;
	wire new_net_11885;
	wire new_net_12474;
	wire new_net_13008;
	wire new_net_14162;
	wire _1250_;
	wire new_net_235;
	wire new_net_1942;
	wire new_net_3003;
	wire new_net_4600;
	wire new_net_6410;
	wire new_net_9936;
	wire new_net_10017;
	wire _1082_;
	wire new_net_6943;
	wire new_net_19102;
	wire new_net_234;
	wire new_net_5317;
	wire new_net_5672;
	wire new_net_18567;
	wire new_net_8290;
	wire _1251_;
	wire new_net_1328;
	wire new_net_1432;
	wire _1083_;
	wire new_net_1358;
	wire new_net_5867;
	wire new_net_19532;
	wire new_net_20830;
	wire new_net_20911;
	wire _1252_;
	wire new_net_3006;
	wire _1084_;
	wire new_net_1430;
	wire new_net_10855;
	wire new_net_9081;
	wire new_net_10962;
	wire new_net_14762;
	wire _0070_;
	wire new_net_3002;
	wire new_net_1414;
	wire new_net_10016;
	wire new_net_9382;
	wire new_net_13322;
	wire new_net_12263;
	wire new_net_14691;
	wire _1253_;
	wire _1085_;
	wire new_net_1609;
	wire new_net_3863;
	wire new_net_5750;
	wire new_net_10526;
	wire new_net_11886;
	wire new_net_12473;
	wire new_net_8288;
	wire new_net_9076;
	wire new_net_9935;
	wire new_net_6942;
	wire new_net_10140;
	wire _1254_;
	wire new_net_230;
	wire new_net_2291;
	wire new_net_5665;
	wire new_net_16986;
	wire _1086_;
	wire new_net_5516;
	wire new_net_19208;
	wire new_net_20828;
	wire new_net_8289;
	wire new_net_1429;
	wire new_net_4599;
	wire new_net_5514;
	wire new_net_9930;
	wire new_net_10142;
	wire new_net_4909;
	wire _1255_;
	wire _1087_;
	wire new_net_1610;
	wire new_net_6640;
	wire new_net_10524;
	wire new_net_9907;
	wire new_net_19533;
	wire new_net_19647;
	wire new_net_20829;
	wire new_net_18156;
	wire new_net_10527;
	wire new_net_10856;
	wire new_net_10014;
	wire new_net_10963;
	wire new_net_14763;
	wire new_net_19209;
	wire _1256_;
	wire new_net_1405;
	wire new_net_5754;
	wire new_net_9080;
	wire new_net_4598;
	wire new_net_9016;
	wire new_net_3859;
	wire new_net_5873;
	wire new_net_6783;
	wire new_net_9390;
	wire new_net_10145;
	wire new_net_15232;
	wire new_net_16248;
	wire new_net_12264;
	wire new_net_14692;
	wire new_net_5520;
	wire new_net_11887;
	wire new_net_13010;
	wire new_net_10705;
	wire new_net_14164;
	wire _1257_;
	wire new_net_3004;
	wire _1089_;
	wire new_net_5395;
	wire new_net_6641;
	wire new_net_14620;
	wire new_net_10704;
	wire new_net_5868;
	wire new_net_18290;
	wire new_net_1407;
	wire new_net_1604;
	wire new_net_5518;
	wire new_net_9270;
	wire new_net_18604;
	wire new_net_20372;
	wire new_net_19064;
	wire new_net_8799;
	wire new_net_1403;
	wire _1258_;
	wire _1090_;
	wire new_net_9071;
	wire new_net_10713;
	wire new_net_19206;
	wire new_net_1329;
	wire new_net_9273;
	wire new_net_10708;
	wire new_net_15670;
	wire new_net_18296;
	wire new_net_19534;
	wire new_net_19648;
	wire new_net_20913;
	wire new_net_14764;
	wire _1091_;
	wire _1259_;
	wire new_net_6422;
	wire new_net_10857;
	wire new_net_10964;
	wire new_net_19210;
	wire new_net_21105;
	wire new_net_10139;
	wire new_net_8282;
	wire new_net_226;
	wire new_net_1363;
	wire new_net_10532;
	wire new_net_18289;
	wire new_net_15233;
	wire new_net_16249;
	wire new_net_12265;
	wire new_net_14693;
	wire _1092_;
	wire _1260_;
	wire new_net_3440;
	wire new_net_11888;
	wire new_net_13011;
	wire new_net_9939;
	wire new_net_1367;
	wire new_net_5755;
	wire new_net_6401;
	wire new_net_15664;
	wire _1093_;
	wire new_net_4910;
	wire _1261_;
	wire new_net_1327;
	wire new_net_1941;
	wire new_net_9268;
	wire new_net_3857;
	wire new_net_5874;
	wire new_net_12364;
	wire new_net_3864;
	wire new_net_6542;
	wire new_net_6408;
	wire new_net_20228;
	wire new_net_1366;
	wire _1262_;
	wire _1094_;
	wire new_net_5322;
	wire new_net_19535;
	wire new_net_20914;
	wire new_net_14765;
	wire new_net_10858;
	wire new_net_1330;
	wire new_net_1353;
	wire new_net_1410;
	wire new_net_10965;
	wire new_net_5320;
	wire new_net_10531;
	wire new_net_19211;
	wire new_net_1360;
	wire _1095_;
	wire _1263_;
	wire new_net_8300;
	wire new_net_9387;
	wire new_net_6786;
	wire new_net_18292;
	wire new_net_20827;
	wire new_net_14166;
	wire new_net_15234;
	wire new_net_1331;
	wire new_net_3439;
	wire new_net_5749;
	wire new_net_8283;
	wire new_net_12266;
	wire new_net_12787;
	wire new_net_16381;
	wire new_net_11889;
	wire new_net_6940;
	wire _1096_;
	wire new_net_1427;
	wire new_net_2288;
	wire _1264_;
	wire new_net_12472;
	wire new_net_6405;
	wire new_net_9018;
	wire new_net_5666;
	wire new_net_18850;
	wire new_net_15668;
	wire new_net_5519;
	wire new_net_8303;
	wire new_net_9392;
	wire new_net_18294;
	wire new_net_20662;
	wire new_net_18536;
	wire new_net_17401;
	wire new_net_10137;
	wire _1265_;
	wire new_net_2292;
	wire new_net_1355;
	wire _1097_;
	wire new_net_6406;
	wire new_net_10712;
	wire new_net_19038;
	wire new_net_20444;
	wire new_net_1332;
	wire new_net_8796;
	wire new_net_19536;
	wire new_net_20915;
	wire new_net_6778;
	wire new_net_10143;
	wire new_net_14766;
	wire _1266_;
	wire new_net_1333;
	wire _1098_;
	wire new_net_6544;
	wire new_net_6639;
	wire new_net_10859;
	wire new_net_10966;
	wire new_net_1939;
	wire new_net_2996;
	wire new_net_5318;
	wire _1596_;
	wire new_net_13472;
	wire new_net_15235;
	wire new_net_16251;
	wire _1267_;
	wire new_net_1404;
	wire _1099_;
	wire new_net_12267;
	wire new_net_14695;
	wire new_net_5752;
	wire new_net_5393;
	wire new_net_6781;
	wire new_net_1362;
	wire new_net_3861;
	wire new_net_8804;
	wire new_net_9077;
	wire new_net_15665;
	wire new_net_9908;
	wire new_net_20826;
	wire new_net_3991;
	wire new_net_17313;
	wire new_net_9269;
	wire _1100_;
	wire _1268_;
	wire new_net_3008;
	wire new_net_10529;
	wire new_net_1352;
	wire new_net_3327;
	wire new_net_18568;
	wire new_net_10530;
	wire new_net_6638;
	wire new_net_20404;
	wire new_net_10148;
	wire _1269_;
	wire new_net_1359;
	wire new_net_1413;
	wire new_net_1431;
	wire _1101_;
	wire new_net_19537;
	wire new_net_20916;
	wire new_net_14767;
	wire new_net_10860;
	wire new_net_10967;
	wire new_net_19321;
	wire new_net_9389;
	wire _1102_;
	wire new_net_6941;
	wire _1270_;
	wire new_net_2998;
	wire new_net_5753;
	wire new_net_5399;
	wire new_net_9931;
	wire new_net_19322;
	wire new_net_13473;
	wire new_net_15236;
	wire new_net_16252;
	wire new_net_2294;
	wire new_net_233;
	wire new_net_12268;
	wire new_net_14696;
	wire new_net_9271;
	wire new_net_11891;
	wire new_net_13014;
	wire _1271_;
	wire new_net_1324;
	wire new_net_2999;
	wire _1103_;
	wire new_net_5751;
	wire new_net_5396;
	wire new_net_10010;
	wire new_net_19315;
	wire new_net_20825;
	wire new_net_17874;
	wire new_net_9384;
	wire new_net_3324;
	wire new_net_5667;
	wire new_net_9909;
	wire new_net_15667;
	wire _1272_;
	wire _1104_;
	wire new_net_8286;
	wire new_net_18293;
	wire new_net_19274;
	wire new_net_6782;
	wire new_net_8798;
	wire new_net_9275;
	wire new_net_9904;
	wire new_net_17610;
	wire new_net_19538;
	wire new_net_20917;
	wire new_net_18157;
	wire new_net_1376;
	wire new_net_10968;
	wire _1273_;
	wire _1105_;
	wire new_net_3858;
	wire new_net_6937;
	wire new_net_6543;
	wire new_net_10861;
	wire new_net_769;
	wire new_net_2212;
	wire new_net_2859;
	wire new_net_13911;
	wire new_net_3767;
	wire new_net_7838;
	wire new_net_8434;
	wire new_net_5190;
	wire new_net_18949;
	wire new_net_20583;
	wire new_net_20229;
	wire new_net_9762;
	wire new_net_13687;
	wire new_net_13392;
	wire new_net_15722;
	wire _1484_;
	wire new_net_565;
	wire new_net_17365;
	wire new_net_15178;
	wire new_net_17388;
	wire new_net_14849;
	wire new_net_5290;
	wire new_net_5962;
	wire new_net_8015;
	wire new_net_759;
	wire new_net_2208;
	wire new_net_4317;
	wire new_net_8181;
	wire new_net_7008;
	wire new_net_8499;
	wire new_net_8945;
	wire new_net_18605;
	wire new_net_20373;
	wire new_net_19065;
	wire _1485_;
	wire new_net_2219;
	wire new_net_7808;
	wire new_net_6527;
	wire new_net_6831;
	wire new_net_19207;
	wire new_net_9606;
	wire new_net_768;
	wire new_net_1184;
	wire new_net_2179;
	wire new_net_3766;
	wire new_net_7809;
	wire _1486_;
	wire new_net_576;
	wire new_net_7257;
	wire new_net_20715;
	wire new_net_17957;
	wire new_net_21057;
	wire new_net_21106;
	wire new_net_1693;
	wire new_net_11495;
	wire new_net_11401;
	wire new_net_14322;
	wire new_net_19234;
	wire new_net_20811;
	wire new_net_5957;
	wire _1487_;
	wire new_net_1691;
	wire new_net_2858;
	wire new_net_7810;
	wire new_net_2213;
	wire new_net_6533;
	wire new_net_10742;
	wire new_net_20584;
	wire new_net_21361;
	wire new_net_13688;
	wire new_net_16904;
	wire new_net_13393;
	wire new_net_2216;
	wire new_net_3761;
	wire new_net_8184;
	wire new_net_17366;
	wire new_net_15723;
	wire new_net_9840;
	wire new_net_14170;
	wire _1488_;
	wire new_net_8178;
	wire new_net_4041;
	wire new_net_6530;
	wire new_net_5294;
	wire new_net_5437;
	wire new_net_8021;
	wire new_net_8428;
	wire new_net_20042;
	wire _1489_;
	wire new_net_8435;
	wire new_net_6740;
	wire new_net_18441;
	wire new_net_18960;
	wire new_net_19233;
	wire new_net_20040;
	wire new_net_566;
	wire new_net_1173;
	wire new_net_2184;
	wire new_net_8180;
	wire new_net_13910;
	wire new_net_20716;
	wire new_net_13912;
	wire new_net_2884;
	wire _1490_;
	wire new_net_3109;
	wire new_net_11496;
	wire new_net_11402;
	wire new_net_4036;
	wire new_net_2454;
	wire new_net_6159;
	wire new_net_19292;
	wire new_net_1692;
	wire new_net_2214;
	wire new_net_4037;
	wire new_net_6150;
	wire new_net_20585;
	wire new_net_13157;
	wire new_net_13689;
	wire new_net_13394;
	wire new_net_15724;
	wire new_net_2217;
	wire new_net_2853;
	wire _1491_;
	wire new_net_17367;
	wire new_net_15180;
	wire new_net_17390;
	wire new_net_18849;
	wire new_net_17774;
	wire new_net_2387;
	wire new_net_2882;
	wire new_net_7010;
	wire new_net_10735;
	wire new_net_18431;
	wire new_net_20043;
	wire new_net_18537;
	wire new_net_19039;
	wire _1492_;
	wire new_net_4039;
	wire new_net_6160;
	wire new_net_18440;
	wire new_net_20445;
	wire new_net_2182;
	wire new_net_2857;
	wire new_net_4900;
	wire new_net_6297;
	wire new_net_21369;
	wire new_net_20933;
	wire new_net_5958;
	wire new_net_8176;
	wire new_net_766;
	wire new_net_1181;
	wire _1493_;
	wire new_net_7262;
	wire new_net_2209;
	wire new_net_4184;
	wire new_net_7839;
	wire new_net_18959;
	wire new_net_3764;
	wire new_net_13913;
	wire new_net_11403;
	wire new_net_11497;
	wire new_net_16069;
	wire new_net_6154;
	wire new_net_18161;
	wire new_net_20813;
	wire new_net_2885;
	wire _1494_;
	wire new_net_3111;
	wire new_net_4320;
	wire new_net_16739;
	wire new_net_20586;
	wire new_net_14172;
	wire new_net_13158;
	wire new_net_15725;
	wire new_net_13395;
	wire new_net_17391;
	wire new_net_13690;
	wire new_net_16906;
	wire new_net_8430;
	wire new_net_15181;
	wire new_net_14324;
	wire new_net_20007;
	wire new_net_5966;
	wire new_net_2382;
	wire new_net_2185;
	wire _1495_;
	wire new_net_7806;
	wire new_net_9760;
	wire new_net_8183;
	wire new_net_4322;
	wire new_net_6532;
	wire new_net_20044;
	wire new_net_18569;
	wire new_net_5287;
	wire new_net_5439;
	wire new_net_15912;
	wire new_net_18242;
	wire new_net_20405;
	wire new_net_9611;
	wire new_net_2183;
	wire _1496_;
	wire new_net_3765;
	wire new_net_7259;
	wire new_net_19231;
	wire new_net_20045;
	wire new_net_5964;
	wire new_net_2177;
	wire new_net_1699;
	wire new_net_7261;
	wire new_net_9838;
	wire new_net_7004;
	wire new_net_6743;
	wire new_net_19232;
	wire new_net_20718;
	wire _1497_;
	wire new_net_1694;
	wire new_net_4182;
	wire new_net_6157;
	wire new_net_11498;
	wire new_net_13914;
	wire new_net_6293;
	wire new_net_8431;
	wire new_net_11404;
	wire _0077_;
	wire new_net_6826;
	wire new_net_764;
	wire new_net_2880;
	wire new_net_5189;
	wire new_net_7005;
	wire new_net_6153;
	wire new_net_18430;
	wire new_net_20587;
	wire new_net_13159;
	wire new_net_9604;
	wire new_net_13691;
	wire _1498_;
	wire new_net_15726;
	wire new_net_17369;
	wire new_net_15182;
	wire new_net_17392;
	wire new_net_17803;
	wire new_net_14853;
	wire new_net_17875;
	wire new_net_6830;
	wire new_net_9761;
	wire new_net_1695;
	wire _1499_;
	wire new_net_2383;
	wire new_net_3113;
	wire new_net_3762;
	wire new_net_4183;
	wire new_net_9843;
	wire new_net_6151;
	wire new_net_18439;
	wire new_net_9834;
	wire new_net_6824;
	wire new_net_2851;
	wire new_net_2174;
	wire new_net_4898;
	wire new_net_8179;
	wire new_net_18158;
	wire _1500_;
	wire new_net_2180;
	wire new_net_7258;
	wire new_net_20047;
	wire new_net_20719;
	wire new_net_4894;
	wire new_net_13396;
	wire new_net_7814;
	wire new_net_11499;
	wire new_net_13915;
	wire new_net_11405;
	wire new_net_14213;
	wire new_net_20815;
	wire new_net_21366;
	wire _1501_;
	wire new_net_5293;
	wire new_net_7807;
	wire new_net_18957;
	wire new_net_20588;
	wire new_net_17393;
	wire new_net_12486;
	wire new_net_13066;
	wire new_net_14174;
	wire new_net_13160;
	wire new_net_13692;
	wire new_net_2380;
	wire new_net_758;
	wire new_net_1178;
	wire new_net_3110;
	wire _1502_;
	wire new_net_5191;
	wire new_net_9832;
	wire new_net_18606;
	wire new_net_20160;
	wire new_net_19066;
	wire new_net_757;
	wire new_net_7813;
	wire new_net_18438;
	wire new_net_4318;
	wire new_net_5632;
	wire new_net_9610;
	wire _1503_;
	wire new_net_2181;
	wire new_net_2854;
	wire new_net_8022;
	wire new_net_7805;
	wire new_net_4323;
	wire new_net_1701;
	wire new_net_4034;
	wire new_net_9609;
	wire new_net_4178;
	wire new_net_6298;
	wire new_net_7836;
	wire new_net_20048;
	wire new_net_20720;
	wire new_net_21367;
	wire new_net_17958;
	wire new_net_21058;
	wire new_net_117;
	wire new_net_1988;
	wire new_net_20231;
	wire new_net_21107;
	wire new_net_6528;
	wire _1504_;
	wire new_net_9763;
	wire new_net_8016;
	wire new_net_7263;
	wire new_net_9839;
	wire new_net_11500;
	wire new_net_13916;
	wire new_net_11406;
	wire new_net_4038;
	wire new_net_6529;
	wire new_net_10734;
	wire new_net_1177;
	wire new_net_14437;
	wire new_net_20589;
	wire new_net_18276;
	wire new_net_10741;
	wire new_net_12487;
	wire new_net_13067;
	wire new_net_14175;
	wire new_net_13161;
	wire _1505_;
	wire new_net_567;
	wire new_net_1176;
	wire new_net_9608;
	wire new_net_13693;
	wire new_net_14485;
	wire new_net_4319;
	wire new_net_4897;
	wire new_net_5963;
	wire new_net_9614;
	wire new_net_6299;
	wire new_net_18433;
	wire new_net_6536;
	wire new_net_10732;
	wire _1506_;
	wire new_net_2455;
	wire new_net_5960;
	wire new_net_8182;
	wire new_net_7843;
	wire new_net_19228;
	wire new_net_10738;
	wire new_net_1700;
	wire new_net_2452;
	wire new_net_5965;
	wire new_net_6828;
	wire _1507_;
	wire new_net_2883;
	wire new_net_5292;
	wire new_net_9841;
	wire new_net_7837;
	wire new_net_20721;
	wire new_net_17954;
	wire new_net_19260;
	wire new_net_1174;
	wire new_net_5192;
	wire new_net_11501;
	wire new_net_13917;
	wire new_net_11407;
	wire new_net_18436;
	wire new_net_20046;
	wire new_net_20817;
	wire _1508_;
	wire new_net_1180;
	wire new_net_2385;
	wire new_net_9836;
	wire new_net_20590;
	wire new_net_14328;
	wire new_net_14916;
	wire new_net_16910;
	wire new_net_12488;
	wire new_net_13068;
	wire new_net_14176;
	wire new_net_13162;
	wire new_net_2176;
	wire new_net_2852;
	wire new_net_1183;
	wire new_net_13436;
	wire new_net_18848;
	wire _1509_;
	wire new_net_575;
	wire new_net_2881;
	wire new_net_13775;
	wire new_net_17773;
	wire new_net_18955;
	wire new_net_19293;
	wire new_net_18538;
	wire new_net_765;
	wire new_net_1179;
	wire new_net_9612;
	wire new_net_9842;
	wire new_net_17403;
	wire new_net_20395;
	wire new_net_19040;
	wire new_net_20446;
	wire _1510_;
	wire new_net_5291;
	wire new_net_3284;
	wire new_net_6294;
	wire new_net_8429;
	wire new_net_14343;
	wire new_net_18437;
	wire new_net_10740;
	wire new_net_4180;
	wire new_net_6156;
	wire new_net_6291;
	wire new_net_8175;
	wire new_net_19294;
	wire new_net_20722;
	wire new_net_19415;
	wire new_net_6825;
	wire _1511_;
	wire new_net_568;
	wire new_net_2389;
	wire new_net_11502;
	wire new_net_13918;
	wire new_net_11408;
	wire new_net_20818;
	wire new_net_20611;
	wire _1603_;
	wire new_net_6534;
	wire new_net_2877;
	wire new_net_4895;
	wire new_net_5438;
	wire new_net_7256;
	wire new_net_18432;
	wire new_net_20591;
	wire new_net_14329;
	wire new_net_14917;
	wire new_net_16911;
	wire new_net_2451;
	wire new_net_6155;
	wire new_net_12489;
	wire new_net_13069;
	wire new_net_14177;
	wire new_net_8947;
	wire new_net_13163;
	wire new_net_6741;
	wire new_net_10737;
	wire new_net_2175;
	wire new_net_4896;
	wire new_net_6292;
	wire new_net_18570;
	wire _1513_;
	wire new_net_1696;
	wire new_net_5967;
	wire new_net_7006;
	wire new_net_9605;
	wire new_net_18954;
	wire new_net_15913;
	wire new_net_18243;
	wire new_net_6827;
	wire new_net_4185;
	wire new_net_5286;
	wire new_net_6295;
	wire new_net_15950;
	wire _1514_;
	wire new_net_8018;
	wire new_net_7844;
	wire new_net_20723;
	wire new_net_21365;
	wire new_net_570;
	wire new_net_2879;
	wire new_net_11503;
	wire new_net_13919;
	wire new_net_11409;
	wire new_net_19295;
	wire new_net_20049;
	wire new_net_20819;
	wire _1515_;
	wire new_net_5961;
	wire new_net_8020;
	wire new_net_7260;
	wire new_net_4179;
	wire new_net_8177;
	wire new_net_7842;
	wire new_net_20592;
	wire new_net_7003;
	wire new_net_14330;
	wire new_net_14918;
	wire new_net_16912;
	wire new_net_12490;
	wire new_net_13070;
	wire new_net_4316;
	wire new_net_5193;
	wire new_net_13164;
	wire new_net_13696;
	wire new_net_17876;
	wire new_net_12347;
	wire _1516_;
	wire new_net_5631;
	wire new_net_6152;
	wire new_net_2215;
	wire new_net_21359;
	wire new_net_16989;
	wire new_net_2386;
	wire new_net_2218;
	wire new_net_4315;
	wire new_net_5288;
	wire new_net_6829;
	wire new_net_19722;
	wire new_net_6535;
	wire _1517_;
	wire new_net_762;
	wire new_net_9837;
	wire new_net_18953;
	wire new_net_2453;
	wire new_net_6161;
	wire new_net_7009;
	wire new_net_20724;
	wire new_net_1369;
	wire new_net_11410;
	wire new_net_14178;
	wire _1518_;
	wire new_net_573;
	wire new_net_2887;
	wire new_net_2855;
	wire new_net_4177;
	wire new_net_11504;
	wire new_net_13920;
	wire new_net_19229;
	wire new_net_574;
	wire new_net_763;
	wire new_net_2211;
	wire new_net_4181;
	wire new_net_20593;
	wire new_net_14859;
	wire new_net_14331;
	wire new_net_14919;
	wire new_net_16913;
	wire new_net_12491;
	wire new_net_13071;
	wire _1519_;
	wire new_net_760;
	wire new_net_13165;
	wire new_net_5289;
	wire new_net_1182;
	wire new_net_761;
	wire new_net_18607;
	wire _1520_;
	wire new_net_1698;
	wire new_net_2178;
	wire new_net_7264;
	wire new_net_21363;
	wire new_net_2384;
	wire new_net_4321;
	wire new_net_7841;
	wire _1521_;
	wire new_net_1697;
	wire new_net_2388;
	wire new_net_2886;
	wire new_net_18435;
	wire new_net_18952;
	wire new_net_20725;
	wire new_net_17959;
	wire new_net_21059;
	wire new_net_6739;
	wire new_net_571;
	wire new_net_2856;
	wire new_net_3112;
	wire new_net_16765;
	wire new_net_11505;
	wire new_net_20821;
	wire new_net_21108;
	wire new_net_5188;
	wire new_net_10733;
	wire _1522_;
	wire new_net_20594;
	wire new_net_14860;
	wire new_net_14332;
	wire new_net_14920;
	wire new_net_16914;
	wire new_net_12492;
	wire new_net_13072;
	wire new_net_14179;
	wire new_net_2876;
	wire new_net_572;
	wire new_net_13166;
	wire new_net_5194;
	wire _1523_;
	wire new_net_4040;
	wire new_net_4314;
	wire new_net_4899;
	wire new_net_9613;
	wire new_net_8019;
	wire new_net_13921;
	wire new_net_12367;
	wire new_net_6742;
	wire new_net_767;
	wire new_net_2860;
	wire new_net_7811;
	wire new_net_4176;
	wire new_net_18608;
	wire new_net_11411;
	wire new_net_5187;
	wire _1524_;
	wire new_net_2381;
	wire new_net_20050;
	wire new_net_16778;
	wire new_net_8433;
	wire new_net_8946;
	wire new_net_20051;
	wire new_net_20726;
	wire new_net_17955;
	wire new_net_9833;
	wire new_net_11506;
	wire new_net_6296;
	wire _1525_;
	wire new_net_1175;
	wire new_net_5959;
	wire new_net_9607;
	wire new_net_8017;
	wire new_net_18951;
	wire new_net_19296;
	wire new_net_13437;
	wire new_net_889;
	wire new_net_4190;
	wire new_net_20559;
	wire new_net_12062;
	wire new_net_18847;
	wire new_net_13776;
	wire new_net_8211;
	wire new_net_13887;
	wire new_net_14896;
	wire new_net_15853;
	wire new_net_17460;
	wire new_net_292;
	wire _0098_;
	wire _1148_;
	wire new_net_11832;
	wire new_net_16018;
	wire new_net_18539;
	wire new_net_17404;
	wire new_net_10379;
	wire new_net_897;
	wire new_net_2744;
	wire new_net_7384;
	wire new_net_19041;
	wire new_net_19723;
	wire new_net_20037;
	wire new_net_20835;
	wire new_net_1955;
	wire _0099_;
	wire _1149_;
	wire new_net_3136;
	wire new_net_8720;
	wire new_net_19827;
	wire new_net_21248;
	wire new_net_3138;
	wire new_net_7273;
	wire new_net_5369;
	wire _0100_;
	wire _1150_;
	wire new_net_893;
	wire _0476_;
	wire new_net_9912;
	wire new_net_20631;
	wire new_net_21011;
	wire new_net_11193;
	wire new_net_10383;
	wire new_net_1949;
	wire new_net_3149;
	wire new_net_10862;
	wire new_net_8490;
	wire new_net_5372;
	wire _1151_;
	wire _0101_;
	wire new_net_8275;
	wire new_net_20560;
	wire new_net_18349;
	wire new_net_17316;
	wire new_net_13888;
	wire new_net_14366;
	wire new_net_15854;
	wire new_net_17461;
	wire new_net_4103;
	wire new_net_5096;
	wire new_net_11833;
	wire new_net_16019;
	wire new_net_7390;
	wire new_net_13052;
	wire new_net_19506;
	wire new_net_18571;
	wire new_net_21015;
	wire new_net_14801;
	wire new_net_895;
	wire _0102_;
	wire _1152_;
	wire new_net_8276;
	wire new_net_19724;
	wire new_net_15914;
	wire new_net_18244;
	wire new_net_11610;
	wire new_net_10377;
	wire new_net_2743;
	wire new_net_9987;
	wire new_net_10466;
	wire new_net_1944;
	wire _0103_;
	wire _1153_;
	wire new_net_8273;
	wire new_net_899;
	wire new_net_4982;
	wire new_net_7391;
	wire new_net_19161;
	wire new_net_20632;
	wire new_net_21012;
	wire _0084_;
	wire new_net_11194;
	wire _0104_;
	wire _1154_;
	wire new_net_10863;
	wire new_net_14365;
	wire new_net_14895;
	wire new_net_1945;
	wire new_net_3878;
	wire new_net_5095;
	wire new_net_7275;
	wire new_net_20561;
	wire new_net_21237;
	wire new_net_12666;
	wire new_net_17048;
	wire new_net_17877;
	wire new_net_15736;
	wire new_net_13889;
	wire new_net_4098;
	wire new_net_15855;
	wire new_net_17462;
	wire _1155_;
	wire _0105_;
	wire new_net_11834;
	wire new_net_16020;
	wire new_net_9992;
	wire new_net_16990;
	wire new_net_19554;
	wire new_net_896;
	wire new_net_8712;
	wire new_net_19171;
	wire new_net_19725;
	wire new_net_898;
	wire _1156_;
	wire _0106_;
	wire new_net_4096;
	wire new_net_9084;
	wire new_net_7381;
	wire new_net_19326;
	wire new_net_14800;
	wire new_net_3127;
	wire new_net_3139;
	wire new_net_4867;
	wire new_net_10376;
	wire new_net_9082;
	wire _1157_;
	wire new_net_5371;
	wire new_net_900;
	wire _0107_;
	wire new_net_3134;
	wire new_net_7382;
	wire new_net_1953;
	wire new_net_20633;
	wire new_net_21013;
	wire new_net_11195;
	wire new_net_297;
	wire new_net_4100;
	wire new_net_8270;
	wire new_net_10864;
	wire new_net_19328;
	wire _1158_;
	wire _0108_;
	wire new_net_14894;
	wire new_net_4716;
	wire new_net_5891;
	wire new_net_20562;
	wire new_net_15737;
	wire new_net_8212;
	wire new_net_11611;
	wire new_net_13890;
	wire new_net_5168;
	wire new_net_14364;
	wire new_net_15856;
	wire new_net_17463;
	wire new_net_11835;
	wire new_net_4379;
	wire new_net_3143;
	wire new_net_8207;
	wire _1159_;
	wire _0109_;
	wire new_net_3128;
	wire new_net_7122;
	wire new_net_8487;
	wire new_net_19726;
	wire new_net_21238;
	wire new_net_1516;
	wire new_net_4097;
	wire new_net_8213;
	wire new_net_19170;
	wire new_net_21246;
	wire new_net_14922;
	wire new_net_18228;
	wire _1160_;
	wire _0110_;
	wire new_net_1950;
	wire new_net_4862;
	wire new_net_7488;
	wire new_net_17960;
	wire new_net_21060;
	wire new_net_16766;
	wire new_net_21109;
	wire new_net_890;
	wire new_net_1954;
	wire new_net_4099;
	wire new_net_4195;
	wire new_net_7120;
	wire new_net_16417;
	wire new_net_19327;
	wire new_net_20634;
	wire new_net_21014;
	wire new_net_8206;
	wire new_net_11196;
	wire new_net_1514;
	wire _1161_;
	wire _0111_;
	wire new_net_4980;
	wire new_net_10865;
	wire new_net_1511;
	wire new_net_3132;
	wire new_net_14893;
	wire new_net_20563;
	wire new_net_15738;
	wire new_net_8715;
	wire new_net_16683;
	wire new_net_11612;
	wire new_net_13891;
	wire _1162_;
	wire _0112_;
	wire new_net_12269;
	wire new_net_13055;
	wire new_net_14363;
	wire new_net_3425;
	wire new_net_19079;
	wire new_net_12368;
	wire new_net_805;
	wire new_net_8718;
	wire new_net_5370;
	wire new_net_1520;
	wire new_net_290;
	wire new_net_4095;
	wire new_net_14799;
	wire new_net_14362;
	wire new_net_19727;
	wire new_net_12247;
	wire new_net_3142;
	wire _1163_;
	wire _0113_;
	wire new_net_3133;
	wire new_net_3875;
	wire new_net_4861;
	wire new_net_7123;
	wire new_net_15565;
	wire new_net_17110;
	wire new_net_1947;
	wire new_net_1512;
	wire new_net_4191;
	wire new_net_8208;
	wire new_net_8488;
	wire new_net_19169;
	wire new_net_17956;
	wire new_net_8205;
	wire new_net_1515;
	wire _1164_;
	wire _0114_;
	wire new_net_3130;
	wire new_net_4987;
	wire new_net_7383;
	wire new_net_5097;
	wire new_net_19251;
	wire new_net_20635;
	wire new_net_11197;
	wire new_net_291;
	wire new_net_10381;
	wire new_net_10866;
	wire new_net_21244;
	wire new_net_16550;
	wire new_net_1948;
	wire _1165_;
	wire _0115_;
	wire new_net_3129;
	wire new_net_14892;
	wire new_net_20564;
	wire new_net_13438;
	wire new_net_12063;
	wire new_net_3976;
	wire new_net_2716;
	wire new_net_18846;
	wire new_net_13244;
	wire new_net_15739;
	wire new_net_11613;
	wire new_net_13892;
	wire new_net_3872;
	wire new_net_4102;
	wire new_net_15858;
	wire new_net_17465;
	wire new_net_17771;
	wire new_net_11837;
	wire new_net_17368;
	wire new_net_18540;
	wire new_net_8491;
	wire new_net_10464;
	wire new_net_14798;
	wire _1166_;
	wire _0116_;
	wire new_net_11644;
	wire new_net_9993;
	wire new_net_19728;
	wire new_net_17405;
	wire new_net_19042;
	wire new_net_345;
	wire new_net_5266;
	wire new_net_10373;
	wire new_net_7279;
	wire new_net_19687;
	wire new_net_19503;
	wire _0117_;
	wire _1167_;
	wire new_net_7126;
	wire new_net_21245;
	wire new_net_852;
	wire new_net_3876;
	wire new_net_19168;
	wire new_net_20636;
	wire new_net_21016;
	wire new_net_16072;
	wire new_net_11198;
	wire new_net_10867;
	wire new_net_14361;
	wire _0118_;
	wire _1168_;
	wire new_net_4983;
	wire new_net_4540;
	wire new_net_8489;
	wire new_net_14891;
	wire new_net_3144;
	wire new_net_4194;
	wire new_net_5630;
	wire new_net_7486;
	wire new_net_9918;
	wire new_net_20565;
	wire new_net_18350;
	wire new_net_16024;
	wire new_net_12109;
	wire new_net_13245;
	wire new_net_5166;
	wire new_net_13893;
	wire new_net_8209;
	wire new_net_11614;
	wire new_net_14527;
	wire _0119_;
	wire _1169_;
	wire new_net_17317;
	wire new_net_14797;
	wire new_net_4186;
	wire new_net_10382;
	wire new_net_19729;
	wire new_net_10944;
	wire new_net_15915;
	wire new_net_18245;
	wire _0120_;
	wire _1170_;
	wire new_net_8714;
	wire new_net_9914;
	wire new_net_894;
	wire new_net_3877;
	wire new_net_4193;
	wire new_net_9996;
	wire new_net_8719;
	wire new_net_19324;
	wire new_net_13140;
	wire _0121_;
	wire _1171_;
	wire new_net_4189;
	wire new_net_1518;
	wire new_net_20637;
	wire new_net_21017;
	wire new_net_10868;
	wire new_net_11199;
	wire new_net_14360;
	wire new_net_13056;
	wire new_net_19167;
	wire new_net_3146;
	wire new_net_5165;
	wire new_net_10462;
	wire new_net_1946;
	wire _1172_;
	wire _0122_;
	wire new_net_14890;
	wire new_net_20566;
	wire new_net_21239;
	wire new_net_706;
	wire new_net_17878;
	wire new_net_16686;
	wire new_net_7124;
	wire new_net_12110;
	wire new_net_7487;
	wire new_net_13246;
	wire new_net_10460;
	wire new_net_15741;
	wire new_net_11615;
	wire new_net_13894;
	wire new_net_2742;
	wire new_net_18489;
	wire new_net_16991;
	wire new_net_15179;
	wire new_net_8711;
	wire new_net_7274;
	wire new_net_14796;
	wire new_net_901;
	wire _0123_;
	wire _1173_;
	wire new_net_7128;
	wire new_net_7315;
	wire new_net_17389;
	wire new_net_19730;
	wire new_net_20432;
	wire new_net_17124;
	wire new_net_892;
	wire new_net_5628;
	wire new_net_8269;
	wire new_net_5744;
	wire new_net_10468;
	wire _0124_;
	wire _1174_;
	wire new_net_9990;
	wire new_net_19325;
	wire new_net_20638;
	wire new_net_20934;
	wire new_net_21018;
	wire new_net_4864;
	wire new_net_10869;
	wire _1175_;
	wire new_net_1952;
	wire _0125_;
	wire new_net_11200;
	wire new_net_20791;
	wire new_net_9916;
	wire new_net_294;
	wire new_net_14889;
	wire new_net_19166;
	wire new_net_19828;
	wire new_net_20567;
	wire new_net_8710;
	wire new_net_12111;
	wire new_net_14529;
	wire new_net_16687;
	wire new_net_13247;
	wire new_net_10467;
	wire new_net_15742;
	wire new_net_11616;
	wire new_net_13895;
	wire new_net_289;
	wire new_net_10592;
	wire new_net_7129;
	wire new_net_14795;
	wire new_net_1519;
	wire new_net_4868;
	wire new_net_10205;
	wire new_net_19731;
	wire new_net_20377;
	wire new_net_7276;
	wire new_net_10463;
	wire _1177_;
	wire _0127_;
	wire new_net_4192;
	wire new_net_14923;
	wire new_net_10461;
	wire new_net_17961;
	wire new_net_21061;
	wire new_net_7125;
	wire _1178_;
	wire _0128_;
	wire new_net_4986;
	wire new_net_3131;
	wire new_net_9989;
	wire new_net_20639;
	wire new_net_20935;
	wire new_net_21019;
	wire new_net_21110;
	wire new_net_10870;
	wire new_net_293;
	wire new_net_3137;
	wire new_net_11201;
	wire new_net_3873;
	wire new_net_4869;
	wire new_net_7271;
	wire _1179_;
	wire _0129_;
	wire new_net_296;
	wire new_net_3140;
	wire new_net_8210;
	wire new_net_10378;
	wire new_net_14888;
	wire new_net_18274;
	wire new_net_12112;
	wire new_net_14530;
	wire new_net_16688;
	wire new_net_13248;
	wire new_net_15743;
	wire new_net_11617;
	wire new_net_13896;
	wire new_net_14358;
	wire new_net_15862;
	wire new_net_17469;
	wire new_net_19080;
	wire new_net_9991;
	wire new_net_5098;
	wire new_net_8271;
	wire new_net_8485;
	wire new_net_5627;
	wire new_net_2745;
	wire _1180_;
	wire _0130_;
	wire new_net_14794;
	wire new_net_14357;
	wire new_net_12248;
	wire new_net_7388;
	wire new_net_7119;
	wire new_net_9919;
	wire new_net_8717;
	wire new_net_9915;
	wire _1181_;
	wire _0131_;
	wire new_net_3148;
	wire new_net_17111;
	wire new_net_4979;
	wire new_net_7387;
	wire new_net_10374;
	wire new_net_19162;
	wire new_net_20640;
	wire new_net_20936;
	wire new_net_21020;
	wire new_net_10871;
	wire new_net_3141;
	wire new_net_1513;
	wire _1182_;
	wire _0132_;
	wire new_net_11202;
	wire new_net_19253;
	wire new_net_16551;
	wire new_net_10459;
	wire new_net_9913;
	wire new_net_10375;
	wire new_net_14887;
	wire new_net_19830;
	wire new_net_20569;
	wire new_net_18845;
	wire new_net_9995;
	wire new_net_13059;
	wire new_net_8274;
	wire new_net_12113;
	wire new_net_14531;
	wire new_net_16689;
	wire new_net_8484;
	wire new_net_13249;
	wire new_net_15744;
	wire _1183_;
	wire new_net_17770;
	wire new_net_2231;
	wire new_net_18541;
	wire new_net_10465;
	wire new_net_14793;
	wire new_net_10380;
	wire new_net_14885;
	wire new_net_19164;
	wire new_net_19733;
	wire new_net_8841;
	wire new_net_11645;
	wire new_net_17406;
	wire new_net_12173;
	wire new_net_19043;
	wire new_net_9988;
	wire _0134_;
	wire _1184_;
	wire new_net_21241;
	wire new_net_17464;
	wire new_net_8713;
	wire new_net_4101;
	wire new_net_4187;
	wire new_net_7386;
	wire new_net_20568;
	wire _0135_;
	wire new_net_7392;
	wire new_net_8272;
	wire new_net_295;
	wire _1185_;
	wire new_net_16105;
	wire new_net_20038;
	wire new_net_20641;
	wire new_net_20937;
	wire new_net_21021;
	wire _0483_;
	wire new_net_20614;
	wire new_net_7277;
	wire new_net_10872;
	wire new_net_10458;
	wire new_net_902;
	wire new_net_5167;
	wire new_net_11203;
	wire new_net_14356;
	wire new_net_3126;
	wire new_net_7127;
	wire new_net_7278;
	wire new_net_5629;
	wire _1186_;
	wire _0136_;
	wire new_net_14886;
	wire new_net_19323;
	wire new_net_19831;
	wire new_net_20570;
	wire new_net_13060;
	wire new_net_12114;
	wire new_net_14532;
	wire new_net_16690;
	wire new_net_13250;
	wire new_net_15745;
	wire new_net_888;
	wire new_net_7272;
	wire new_net_11619;
	wire new_net_13898;
	wire new_net_9911;
	wire new_net_3145;
	wire new_net_1517;
	wire _1187_;
	wire _0137_;
	wire new_net_14792;
	wire new_net_4188;
	wire new_net_19734;
	wire new_net_15916;
	wire new_net_18246;
	wire new_net_14355;
	wire new_net_19163;
	wire new_net_17257;
	wire new_net_16859;
	wire new_net_2719;
	wire new_net_4865;
	wire new_net_8486;
	wire new_net_3147;
	wire _0138_;
	wire new_net_1951;
	wire _1188_;
	wire new_net_8204;
	wire new_net_9083;
	wire new_net_3135;
	wire new_net_20039;
	wire new_net_20642;
	wire new_net_20938;
	wire new_net_21022;
	wire new_net_9986;
	wire new_net_4863;
	wire new_net_10873;
	wire new_net_891;
	wire _0139_;
	wire _1189_;
	wire new_net_14791;
	wire new_net_11204;
	wire new_net_4985;
	wire new_net_21240;
	wire new_net_4125;
	wire new_net_9325;
	wire new_net_12745;
	wire new_net_16229;
	wire new_net_17879;
	wire new_net_12350;
	wire new_net_10190;
	wire new_net_1839;
	wire new_net_14710;
	wire new_net_7974;
	wire new_net_6237;
	wire new_net_20524;
	wire new_net_18490;
	wire new_net_16992;
	wire new_net_14533;
	wire new_net_13569;
	wire new_net_13215;
	wire new_net_13390;
	wire new_net_15521;
	wire new_net_17412;
	wire new_net_9668;
	wire new_net_1076;
	wire new_net_10354;
	wire new_net_15095;
	wire new_net_20433;
	wire new_net_17125;
	wire new_net_10546;
	wire new_net_9664;
	wire new_net_970;
	wire new_net_2191;
	wire new_net_4990;
	wire new_net_5345;
	wire new_net_20505;
	wire new_net_14217;
	wire _1779_;
	wire new_net_14709;
	wire new_net_20530;
	wire new_net_579;
	wire new_net_1841;
	wire new_net_2809;
	wire new_net_7306;
	wire new_net_8310;
	wire new_net_2095;
	wire _1780_;
	wire new_net_13650;
	wire new_net_20320;
	wire new_net_7567;
	wire new_net_13391;
	wire new_net_14556;
	wire new_net_1299;
	wire new_net_2091;
	wire new_net_11507;
	wire new_net_11519;
	wire new_net_10353;
	wire new_net_5890;
	wire new_net_7371;
	wire new_net_16445;
	wire _1781_;
	wire new_net_620;
	wire new_net_1039;
	wire new_net_2800;
	wire new_net_7976;
	wire new_net_20525;
	wire new_net_10690;
	wire new_net_13133;
	wire new_net_13216;
	wire new_net_14534;
	wire new_net_16575;
	wire new_net_16740;
	wire new_net_12000;
	wire new_net_13389;
	wire new_net_13570;
	wire new_net_14554;
	wire _1782_;
	wire new_net_10196;
	wire new_net_1834;
	wire new_net_622;
	wire new_net_288;
	wire new_net_14924;
	wire new_net_19275;
	wire new_net_16454;
	wire new_net_2102;
	wire new_net_2812;
	wire new_net_4969;
	wire new_net_5136;
	wire new_net_16834;
	wire new_net_20355;
	wire new_net_17962;
	wire new_net_21062;
	wire new_net_5529;
	wire new_net_10361;
	wire _1783_;
	wire new_net_16768;
	wire new_net_7318;
	wire new_net_1842;
	wire new_net_21111;
	wire new_net_2801;
	wire new_net_1844;
	wire new_net_5943;
	wire new_net_10065;
	wire new_net_5889;
	wire _1784_;
	wire new_net_11508;
	wire new_net_14711;
	wire new_net_11520;
	wire new_net_287;
	wire new_net_17922;
	wire new_net_10359;
	wire new_net_1843;
	wire new_net_578;
	wire new_net_2194;
	wire new_net_4988;
	wire new_net_8307;
	wire new_net_20526;
	wire new_net_12271;
	wire new_net_19081;
	wire new_net_9214;
	wire new_net_12370;
	wire new_net_15310;
	wire new_net_17154;
	wire _1785_;
	wire new_net_13134;
	wire new_net_5531;
	wire new_net_10199;
	wire new_net_13217;
	wire new_net_14535;
	wire new_net_16576;
	wire new_net_16741;
	wire new_net_12249;
	wire new_net_968;
	wire new_net_4332;
	wire new_net_6241;
	wire new_net_10171;
	wire new_net_1465;
	wire new_net_15567;
	wire _1786_;
	wire new_net_4995;
	wire new_net_5104;
	wire new_net_282;
	wire new_net_971;
	wire new_net_6236;
	wire new_net_124;
	wire new_net_580;
	wire new_net_2097;
	wire new_net_2190;
	wire new_net_9665;
	wire new_net_8309;
	wire new_net_18351;
	wire _1787_;
	wire new_net_4991;
	wire new_net_1072;
	wire new_net_8305;
	wire new_net_20859;
	wire new_net_13682;
	wire new_net_585;
	wire new_net_967;
	wire new_net_11509;
	wire new_net_12840;
	wire new_net_14712;
	wire new_net_11521;
	wire new_net_18844;
	wire _1788_;
	wire new_net_10547;
	wire new_net_1074;
	wire new_net_4903;
	wire new_net_20527;
	wire new_net_17370;
	wire new_net_12208;
	wire new_net_13779;
	wire new_net_17769;
	wire new_net_18542;
	wire new_net_15311;
	wire new_net_17155;
	wire new_net_13135;
	wire new_net_7336;
	wire new_net_13218;
	wire new_net_14536;
	wire new_net_16577;
	wire new_net_16742;
	wire new_net_1295;
	wire new_net_5350;
	wire new_net_11646;
	wire new_net_17407;
	wire _1789_;
	wire new_net_16443;
	wire new_net_14347;
	wire new_net_8308;
	wire new_net_8576;
	wire new_net_10200;
	wire new_net_16453;
	wire new_net_16106;
	wire new_net_5137;
	wire _1790_;
	wire new_net_4992;
	wire new_net_10193;
	wire new_net_588;
	wire new_net_4531;
	wire new_net_16074;
	wire new_net_10180;
	wire new_net_1290;
	wire new_net_5524;
	wire new_net_16744;
	wire new_net_13204;
	wire _1791_;
	wire new_net_6679;
	wire new_net_11510;
	wire new_net_14713;
	wire new_net_11522;
	wire new_net_10470;
	wire new_net_7565;
	wire new_net_2098;
	wire new_net_6676;
	wire new_net_20528;
	wire new_net_12308;
	wire new_net_4331;
	wire new_net_15312;
	wire new_net_17156;
	wire _1792_;
	wire new_net_13136;
	wire new_net_7335;
	wire new_net_13219;
	wire new_net_14537;
	wire new_net_16578;
	wire new_net_16743;
	wire new_net_18620;
	wire new_net_11618;
	wire new_net_10268;
	wire new_net_15917;
	wire new_net_18247;
	wire new_net_6683;
	wire new_net_2195;
	wire new_net_7307;
	wire new_net_9889;
	wire new_net_15954;
	wire new_net_16860;
	wire new_net_4337;
	wire new_net_6677;
	wire new_net_5525;
	wire new_net_10358;
	wire new_net_5346;
	wire _1793_;
	wire new_net_11944;
	wire new_net_13142;
	wire new_net_625;
	wire new_net_1038;
	wire new_net_4904;
	wire new_net_10181;
	wire new_net_5103;
	wire new_net_10360;
	wire _1794_;
	wire new_net_628;
	wire new_net_1035;
	wire new_net_2803;
	wire new_net_586;
	wire new_net_16447;
	wire new_net_13329;
	wire new_net_7975;
	wire new_net_5140;
	wire new_net_6234;
	wire new_net_10198;
	wire new_net_2186;
	wire new_net_2805;
	wire new_net_123;
	wire new_net_1835;
	wire new_net_5886;
	wire new_net_9667;
	wire new_net_12744;
	wire new_net_15307;
	wire new_net_1296;
	wire new_net_6233;
	wire new_net_10170;
	wire new_net_17051;
	wire new_net_5354;
	wire _1795_;
	wire new_net_4534;
	wire new_net_16230;
	wire new_net_12351;
	wire new_net_17880;
	wire new_net_18491;
	wire new_net_6955;
	wire new_net_7763;
	wire new_net_16993;
	wire new_net_15100;
	wire new_net_15526;
	wire new_net_17606;
	wire new_net_15313;
	wire new_net_17157;
	wire new_net_13137;
	wire new_net_8573;
	wire new_net_13220;
	wire new_net_14538;
	wire new_net_16579;
	wire new_net_10545;
	wire _1796_;
	wire new_net_2187;
	wire new_net_7308;
	wire new_net_4920;
	wire new_net_1030;
	wire new_net_4339;
	wire new_net_5349;
	wire new_net_16452;
	wire new_net_7460;
	wire new_net_14218;
	wire new_net_16021;
	wire new_net_6678;
	wire _1797_;
	wire new_net_1028;
	wire new_net_18005;
	wire new_net_10351;
	wire new_net_4338;
	wire new_net_8575;
	wire new_net_2810;
	wire _1798_;
	wire new_net_10201;
	wire new_net_9662;
	wire new_net_11512;
	wire new_net_14715;
	wire new_net_11524;
	wire new_net_127;
	wire new_net_286;
	wire new_net_1040;
	wire new_net_1085;
	wire new_net_10197;
	wire _0770_;
	wire new_net_15101;
	wire new_net_15527;
	wire new_net_17607;
	wire new_net_14549;
	wire new_net_15314;
	wire new_net_17158;
	wire _1799_;
	wire new_net_4996;
	wire new_net_13138;
	wire new_net_10544;
	wire new_net_20379;
	wire new_net_5530;
	wire new_net_1075;
	wire new_net_1845;
	wire new_net_2804;
	wire new_net_2092;
	wire new_net_4901;
	wire new_net_4968;
	wire new_net_9959;
	wire new_net_14925;
	wire _1800_;
	wire new_net_2193;
	wire new_net_129;
	wire new_net_18225;
	wire new_net_16835;
	wire new_net_17963;
	wire new_net_21063;
	wire new_net_112;
	wire new_net_583;
	wire new_net_623;
	wire new_net_2093;
	wire new_net_4333;
	wire new_net_16769;
	wire new_net_21112;
	wire new_net_1027;
	wire new_net_5139;
	wire new_net_6240;
	wire _1801_;
	wire new_net_587;
	wire new_net_122;
	wire new_net_3298;
	wire new_net_18866;
	wire new_net_5938;
	wire new_net_11525;
	wire new_net_2811;
	wire new_net_4840;
	wire new_net_9658;
	wire new_net_11513;
	wire new_net_14716;
	wire new_net_17923;
	wire new_net_2189;
	wire new_net_4334;
	wire new_net_10177;
	wire _1802_;
	wire new_net_10548;
	wire new_net_130;
	wire new_net_973;
	wire new_net_16444;
	wire new_net_19082;
	wire new_net_12868;
	wire new_net_15173;
	wire new_net_17419;
	wire new_net_15102;
	wire new_net_15528;
	wire new_net_17608;
	wire new_net_15315;
	wire new_net_17159;
	wire new_net_13139;
	wire new_net_1837;
	wire new_net_12371;
	wire new_net_12250;
	wire _1803_;
	wire new_net_5522;
	wire new_net_131;
	wire new_net_1297;
	wire new_net_2100;
	wire new_net_9661;
	wire new_net_10689;
	wire new_net_16451;
	wire new_net_15323;
	wire new_net_16782;
	wire new_net_17113;
	wire new_net_2196;
	wire _1804_;
	wire new_net_10688;
	wire new_net_581;
	wire new_net_974;
	wire new_net_16448;
	wire new_net_8313;
	wire new_net_2814;
	wire new_net_619;
	wire new_net_1083;
	wire new_net_9114;
	wire new_net_13683;
	wire new_net_11526;
	wire new_net_6239;
	wire new_net_10174;
	wire _1805_;
	wire new_net_5527;
	wire new_net_7303;
	wire new_net_11514;
	wire new_net_14717;
	wire new_net_16542;
	wire new_net_18616;
	wire new_net_12066;
	wire new_net_18843;
	wire new_net_2813;
	wire new_net_2802;
	wire new_net_4533;
	wire new_net_5352;
	wire new_net_20531;
	wire new_net_17371;
	wire new_net_13780;
	wire new_net_17768;
	wire new_net_18543;
	wire new_net_4532;
	wire new_net_12869;
	wire new_net_15174;
	wire new_net_17420;
	wire new_net_15103;
	wire new_net_15529;
	wire new_net_17609;
	wire new_net_15316;
	wire new_net_17160;
	wire _1806_;
	wire new_net_11647;
	wire new_net_17408;
	wire new_net_339;
	wire new_net_1041;
	wire new_net_6232;
	wire new_net_6315;
	wire new_net_14837;
	wire new_net_15877;
	wire new_net_14348;
	wire new_net_626;
	wire _1807_;
	wire new_net_5523;
	wire new_net_10541;
	wire new_net_1840;
	wire new_net_17466;
	wire new_net_4340;
	wire new_net_10175;
	wire new_net_618;
	wire new_net_3448;
	wire new_net_5526;
	wire new_net_7338;
	wire new_net_10542;
	wire new_net_7309;
	wire new_net_16107;
	wire _0490_;
	wire new_net_16075;
	wire new_net_2831;
	wire new_net_6238;
	wire _1808_;
	wire new_net_6680;
	wire new_net_584;
	wire new_net_1301;
	wire new_net_7337;
	wire new_net_16745;
	wire new_net_11527;
	wire new_net_14718;
	wire new_net_8312;
	wire new_net_10192;
	wire new_net_4993;
	wire new_net_6682;
	wire new_net_7301;
	wire new_net_11515;
	wire new_net_10178;
	wire new_net_13205;
	wire new_net_15701;
	wire new_net_2096;
	wire new_net_1836;
	wire _1809_;
	wire new_net_8574;
	wire new_net_20532;
	wire new_net_18352;
	wire new_net_12870;
	wire new_net_15530;
	wire new_net_16583;
	wire new_net_17161;
	wire new_net_13141;
	wire new_net_17421;
	wire new_net_14542;
	wire new_net_15317;
	wire new_net_13224;
	wire new_net_7566;
	wire new_net_18621;
	wire new_net_15918;
	wire new_net_18248;
	wire new_net_4902;
	wire new_net_6231;
	wire new_net_4989;
	wire _1810_;
	wire new_net_1031;
	wire new_net_128;
	wire new_net_284;
	wire new_net_5528;
	wire new_net_10352;
	wire new_net_5351;
	wire new_net_15955;
	wire new_net_16861;
	wire new_net_283;
	wire new_net_624;
	wire new_net_972;
	wire new_net_2808;
	wire new_net_4335;
	wire new_net_16450;
	wire new_net_4535;
	wire _1811_;
	wire new_net_2192;
	wire new_net_11945;
	wire new_net_8577;
	wire new_net_18304;
	wire new_net_5237;
	wire new_net_285;
	wire new_net_9666;
	wire new_net_13330;
	wire new_net_11516;
	wire new_net_14719;
	wire new_net_1846;
	wire new_net_11528;
	wire new_net_4994;
	wire _1812_;
	wire new_net_1082;
	wire new_net_8569;
	wire new_net_2099;
	wire new_net_16979;
	wire new_net_9328;
	wire new_net_12743;
	wire new_net_6876;
	wire new_net_17809;
	wire new_net_2188;
	wire new_net_1293;
	wire new_net_5347;
	wire new_net_20533;
	wire new_net_9757;
	wire new_net_17052;
	wire new_net_17881;
	wire new_net_18492;
	wire new_net_16994;
	wire new_net_8306;
	wire new_net_12847;
	wire new_net_12871;
	wire new_net_15176;
	wire new_net_14545;
	wire new_net_15105;
	wire new_net_15531;
	wire new_net_17611;
	wire new_net_10173;
	wire new_net_15318;
	wire new_net_1033;
	wire new_net_1084;
	wire new_net_2101;
	wire new_net_19697;
	wire new_net_15049;
	wire new_net_19717;
	wire new_net_5735;
	wire new_net_2466;
	wire new_net_6261;
	wire new_net_5138;
	wire new_net_6235;
	wire _1814_;
	wire new_net_627;
	wire new_net_5348;
	wire new_net_2094;
	wire new_net_582;
	wire new_net_16022;
	wire new_net_1298;
	wire new_net_10357;
	wire new_net_9660;
	wire new_net_18052;
	wire new_net_18006;
	wire new_net_10543;
	wire new_net_1300;
	wire _1815_;
	wire new_net_16116;
	wire new_net_1034;
	wire new_net_10194;
	wire new_net_11529;
	wire new_net_11517;
	wire new_net_10179;
	wire new_net_1029;
	wire new_net_975;
	wire new_net_4967;
	wire new_net_5353;
	wire new_net_14720;
	wire new_net_5133;
	wire _1816_;
	wire new_net_20534;
	wire new_net_12848;
	wire new_net_12872;
	wire new_net_15177;
	wire new_net_17423;
	wire new_net_15106;
	wire new_net_15532;
	wire new_net_17612;
	wire new_net_15319;
	wire new_net_17163;
	wire new_net_13143;
	wire new_net_15832;
	wire new_net_125;
	wire new_net_1294;
	wire _1817_;
	wire new_net_1079;
	wire new_net_969;
	wire new_net_9663;
	wire new_net_19698;
	wire new_net_1725;
	wire new_net_14926;
	wire new_net_10172;
	wire new_net_1292;
	wire new_net_4537;
	wire new_net_5134;
	wire new_net_16449;
	wire new_net_9752;
	wire new_net_16836;
	wire new_net_17964;
	wire new_net_21064;
	wire new_net_8311;
	wire new_net_616;
	wire new_net_2807;
	wire _1818_;
	wire new_net_4839;
	wire new_net_10362;
	wire new_net_10191;
	wire new_net_7302;
	wire new_net_16446;
	wire new_net_16770;
	wire new_net_21113;
	wire new_net_5238;
	wire new_net_8571;
	wire new_net_2806;
	wire new_net_1081;
	wire new_net_1291;
	wire new_net_6681;
	wire new_net_10687;
	wire new_net_10356;
	wire new_net_13581;
	wire new_net_14649;
	wire new_net_13664;
	wire new_net_5885;
	wire new_net_11518;
	wire new_net_11530;
	wire new_net_1032;
	wire new_net_4336;
	wire new_net_1080;
	wire _1819_;
	wire new_net_8572;
	wire new_net_18867;
	wire new_net_17924;
	wire _0630_;
	wire new_net_19083;
	wire new_net_12289;
	wire new_net_12372;
	wire new_net_10388;
	wire new_net_417;
	wire new_net_1891;
	wire new_net_2067;
	wire new_net_4437;
	wire new_net_20396;
	wire new_net_12251;
	wire new_net_8220;
	wire new_net_12660;
	wire new_net_12281;
	wire new_net_16134;
	wire new_net_13699;
	wire new_net_7205;
	wire new_net_15604;
	wire new_net_17483;
	wire new_net_17732;
	wire new_net_163;
	wire new_net_15888;
	wire new_net_1886;
	wire new_net_8155;
	wire new_net_16783;
	wire new_net_19747;
	wire new_net_19783;
	wire new_net_14239;
	wire new_net_18309;
	wire new_net_171;
	wire new_net_3755;
	wire new_net_4492;
	wire new_net_3683;
	wire new_net_10776;
	wire new_net_19363;
	wire new_net_3789;
	wire new_net_8867;
	wire new_net_21443;
	wire new_net_4387;
	wire new_net_20861;
	wire new_net_13684;
	wire new_net_10484;
	wire new_net_5277;
	wire new_net_2747;
	wire new_net_5308;
	wire new_net_20100;
	wire new_net_20727;
	wire new_net_16543;
	wire new_net_12067;
	wire new_net_8051;
	wire new_net_11321;
	wire new_net_555;
	wire new_net_1703;
	wire new_net_8152;
	wire new_net_10922;
	wire new_net_14061;
	wire new_net_17372;
	wire new_net_2230;
	wire new_net_18544;
	wire new_net_8061;
	wire new_net_9101;
	wire new_net_6487;
	wire new_net_6491;
	wire new_net_711;
	wire new_net_2065;
	wire new_net_12623;
	wire new_net_5316;
	wire new_net_11648;
	wire new_net_17409;
	wire new_net_15545;
	wire new_net_17544;
	wire new_net_16325;
	wire new_net_12661;
	wire new_net_17484;
	wire new_net_16610;
	wire new_net_17733;
	wire new_net_12282;
	wire new_net_16135;
	wire new_net_13700;
	wire new_net_15605;
	wire new_net_14349;
	wire new_net_17734;
	wire new_net_17467;
	wire new_net_10487;
	wire new_net_15889;
	wire new_net_9100;
	wire new_net_1240;
	wire new_net_95;
	wire new_net_2752;
	wire new_net_418;
	wire new_net_10693;
	wire new_net_169;
	wire new_net_19748;
	wire new_net_90;
	wire new_net_4439;
	wire new_net_7202;
	wire new_net_16108;
	wire new_net_12622;
	wire new_net_19364;
	wire new_net_1045;
	wire new_net_16076;
	wire new_net_3787;
	wire new_net_6496;
	wire new_net_420;
	wire new_net_6399;
	wire new_net_21444;
	wire new_net_16395;
	wire new_net_13276;
	wire new_net_16746;
	wire new_net_8555;
	wire new_net_6144;
	wire new_net_18996;
	wire new_net_20101;
	wire new_net_20728;
	wire new_net_12652;
	wire new_net_13290;
	wire new_net_15702;
	wire new_net_10477;
	wire new_net_10700;
	wire new_net_10774;
	wire new_net_11322;
	wire new_net_173;
	wire new_net_1892;
	wire new_net_3759;
	wire new_net_3774;
	wire new_net_19149;
	wire new_net_20397;
	wire new_net_18353;
	wire new_net_13840;
	wire new_net_8553;
	wire new_net_1890;
	wire new_net_1232;
	wire new_net_3790;
	wire new_net_4490;
	wire new_net_18622;
	wire new_net_15919;
	wire new_net_18249;
	wire new_net_13606;
	wire new_net_12662;
	wire new_net_4432;
	wire new_net_12283;
	wire new_net_16136;
	wire new_net_13701;
	wire new_net_17545;
	wire new_net_15305;
	wire new_net_15606;
	wire new_net_17485;
	wire new_net_4042;
	wire new_net_21370;
	wire new_net_16862;
	wire new_net_2720;
	wire new_net_10767;
	wire new_net_8055;
	wire new_net_8222;
	wire new_net_15890;
	wire new_net_556;
	wire new_net_700;
	wire new_net_1708;
	wire new_net_19006;
	wire new_net_19140;
	wire new_net_19749;
	wire new_net_11946;
	wire new_net_5278;
	wire new_net_8561;
	wire new_net_19365;
	wire new_net_10775;
	wire new_net_3791;
	wire new_net_10923;
	wire new_net_21445;
	wire new_net_13331;
	wire new_net_7199;
	wire new_net_165;
	wire new_net_1238;
	wire new_net_20102;
	wire new_net_20729;
	wire new_net_17810;
	wire new_net_8863;
	wire new_net_9862;
	wire new_net_707;
	wire new_net_3788;
	wire new_net_6397;
	wire new_net_11323;
	wire new_net_20398;
	wire new_net_17882;
	wire new_net_18493;
	wire new_net_16995;
	wire new_net_21360;
	wire new_net_8556;
	wire new_net_1707;
	wire new_net_419;
	wire new_net_4491;
	wire new_net_121;
	wire new_net_5282;
	wire new_net_8647;
	wire new_net_15183;
	wire new_net_19559;
	wire new_net_9825;
	wire new_net_20436;
	wire new_net_13607;
	wire new_net_17735;
	wire new_net_12663;
	wire new_net_13702;
	wire new_net_12284;
	wire new_net_17546;
	wire new_net_16327;
	wire new_net_16612;
	wire new_net_5280;
	wire new_net_15050;
	wire new_net_20212;
	wire new_net_2462;
	wire new_net_4431;
	wire new_net_3771;
	wire new_net_6485;
	wire new_net_19750;
	wire new_net_19786;
	wire new_net_14220;
	wire new_net_18088;
	wire new_net_16023;
	wire new_net_8862;
	wire new_net_10481;
	wire new_net_558;
	wire new_net_3758;
	wire new_net_3768;
	wire new_net_5313;
	wire new_net_19005;
	wire new_net_19366;
	wire new_net_18053;
	wire new_net_18007;
	wire new_net_16117;
	wire new_net_712;
	wire new_net_2751;
	wire new_net_168;
	wire new_net_414;
	wire new_net_560;
	wire new_net_3786;
	wire new_net_6495;
	wire new_net_5315;
	wire new_net_21446;
	wire new_net_6053;
	wire new_net_8562;
	wire new_net_4436;
	wire new_net_6493;
	wire new_net_12620;
	wire new_net_20103;
	wire new_net_20730;
	wire new_net_13509;
	wire new_net_9859;
	wire new_net_8218;
	wire new_net_11324;
	wire new_net_15607;
	wire new_net_10924;
	wire new_net_19148;
	wire new_net_20399;
	wire new_net_4380;
	wire new_net_9673;
	wire new_net_422;
	wire new_net_2755;
	wire new_net_15833;
	wire new_net_3688;
	wire new_net_9858;
	wire new_net_13608;
	wire new_net_4434;
	wire new_net_12285;
	wire new_net_16138;
	wire new_net_13703;
	wire new_net_175;
	wire new_net_89;
	wire new_net_17129;
	wire new_net_14927;
	wire new_net_8147;
	wire new_net_14058;
	wire new_net_8056;
	wire new_net_8219;
	wire new_net_564;
	wire new_net_167;
	wire new_net_3446;
	wire new_net_3756;
	wire new_net_4488;
	wire new_net_6141;
	wire new_net_16837;
	wire new_net_17965;
	wire new_net_21065;
	wire new_net_3776;
	wire new_net_3685;
	wire new_net_92;
	wire new_net_164;
	wire new_net_2749;
	wire new_net_19367;
	wire new_net_20326;
	wire new_net_16771;
	wire new_net_21114;
	wire new_net_4455;
	wire new_net_8059;
	wire new_net_1230;
	wire new_net_4433;
	wire new_net_10694;
	wire new_net_19004;
	wire new_net_21447;
	wire new_net_13582;
	wire new_net_14650;
	wire new_net_18868;
	wire new_net_10480;
	wire new_net_4429;
	wire new_net_9098;
	wire new_net_703;
	wire new_net_2068;
	wire new_net_20104;
	wire new_net_20731;
	wire new_net_17925;
	wire new_net_8153;
	wire new_net_10925;
	wire new_net_9863;
	wire new_net_12664;
	wire new_net_9097;
	wire new_net_11325;
	wire new_net_705;
	wire new_net_1233;
	wire new_net_6139;
	wire new_net_20400;
	wire new_net_19084;
	wire new_net_8149;
	wire new_net_7206;
	wire new_net_708;
	wire new_net_557;
	wire new_net_1704;
	wire new_net_19147;
	wire new_net_12373;
	wire new_net_15239;
	wire new_net_12252;
	wire new_net_14056;
	wire new_net_16329;
	wire new_net_16614;
	wire new_net_17548;
	wire new_net_10701;
	wire new_net_13609;
	wire new_net_12286;
	wire new_net_16139;
	wire new_net_13704;
	wire new_net_15892;
	wire new_net_8868;
	wire new_net_10486;
	wire new_net_9671;
	wire new_net_1889;
	wire new_net_17579;
	wire new_net_6142;
	wire new_net_19752;
	wire new_net_19788;
	wire new_net_15325;
	wire new_net_16784;
	wire new_net_17115;
	wire new_net_14240;
	wire new_net_10698;
	wire new_net_1237;
	wire new_net_415;
	wire new_net_561;
	wire new_net_1702;
	wire new_net_3785;
	wire new_net_19368;
	wire new_net_4164;
	wire new_net_4417;
	wire new_net_6841;
	wire new_net_6393;
	wire new_net_10479;
	wire new_net_2754;
	wire new_net_7200;
	wire new_net_12619;
	wire new_net_21448;
	wire new_net_16555;
	wire new_net_13685;
	wire new_net_10691;
	wire new_net_10773;
	wire new_net_8214;
	wire new_net_10390;
	wire new_net_152;
	wire new_net_3681;
	wire new_net_19003;
	wire new_net_20105;
	wire new_net_20732;
	wire new_net_16544;
	wire new_net_5312;
	wire new_net_10926;
	wire new_net_1888;
	wire new_net_11326;
	wire new_net_20401;
	wire new_net_569;
	wire new_net_17373;
	wire new_net_8154;
	wire new_net_10699;
	wire new_net_8050;
	wire new_net_9676;
	wire new_net_1706;
	wire new_net_18545;
	wire new_net_8847;
	wire new_net_11649;
	wire new_net_17410;
	wire new_net_18303;
	wire new_net_15546;
	wire new_net_3773;
	wire new_net_14055;
	wire new_net_16330;
	wire new_net_16615;
	wire new_net_10692;
	wire new_net_10772;
	wire new_net_13610;
	wire new_net_12665;
	wire new_net_12287;
	wire new_net_16140;
	wire new_net_344;
	wire new_net_15879;
	wire new_net_14350;
	wire new_net_10483;
	wire new_net_8558;
	wire new_net_3760;
	wire new_net_4438;
	wire new_net_4487;
	wire new_net_5285;
	wire new_net_12618;
	wire new_net_19753;
	wire new_net_14359;
	wire new_net_17468;
	wire new_net_10697;
	wire new_net_3684;
	wire new_net_3792;
	wire new_net_19369;
	wire new_net_16109;
	wire _0497_;
	wire new_net_16077;
	wire new_net_9854;
	wire new_net_2750;
	wire new_net_99;
	wire new_net_166;
	wire new_net_21449;
	wire new_net_13277;
	wire new_net_16747;
	wire new_net_172;
	wire new_net_1709;
	wire new_net_20106;
	wire new_net_20733;
	wire new_net_13207;
	wire new_net_18819;
	wire new_net_7826;
	wire new_net_12653;
	wire new_net_8151;
	wire new_net_10927;
	wire new_net_11327;
	wire new_net_18531;
	wire new_net_19002;
	wire new_net_19139;
	wire new_net_20402;
	wire new_net_18354;
	wire new_net_13841;
	wire new_net_12311;
	wire new_net_12612;
	wire new_net_4113;
	wire new_net_8052;
	wire new_net_10386;
	wire new_net_5284;
	wire new_net_18623;
	wire new_net_6147;
	wire new_net_12617;
	wire new_net_16095;
	wire new_net_17550;
	wire new_net_6398;
	wire new_net_14054;
	wire new_net_16331;
	wire new_net_16616;
	wire new_net_8869;
	wire new_net_13611;
	wire new_net_15920;
	wire new_net_10270;
	wire new_net_18250;
	wire new_net_15957;
	wire new_net_10768;
	wire new_net_416;
	wire new_net_2069;
	wire new_net_6497;
	wire new_net_19145;
	wire new_net_19754;
	wire new_net_19790;
	wire new_net_10619;
	wire new_net_10503;
	wire new_net_8864;
	wire new_net_9860;
	wire new_net_8060;
	wire new_net_2066;
	wire new_net_174;
	wire new_net_704;
	wire new_net_18997;
	wire new_net_19370;
	wire new_net_11947;
	wire new_net_8866;
	wire new_net_21450;
	wire new_net_14450;
	wire new_net_13332;
	wire new_net_9857;
	wire new_net_9670;
	wire new_net_559;
	wire new_net_20107;
	wire new_net_20734;
	wire new_net_16981;
	wire new_net_17811;
	wire new_net_6396;
	wire new_net_10928;
	wire new_net_10485;
	wire new_net_12288;
	wire new_net_7201;
	wire new_net_11328;
	wire new_net_20403;
	wire new_net_16233;
	wire new_net_17883;
	wire new_net_18494;
	wire new_net_16996;
	wire new_net_2746;
	wire new_net_19001;
	wire new_net_126;
	wire new_net_15184;
	wire new_net_17394;
	wire new_net_19784;
	wire new_net_19560;
	wire new_net_8646;
	wire new_net_12616;
	wire new_net_16096;
	wire new_net_17551;
	wire new_net_14053;
	wire new_net_16332;
	wire new_net_16617;
	wire new_net_13612;
	wire new_net_8057;
	wire new_net_12667;
	wire new_net_15051;
	wire new_net_20209;
	wire new_net_7824;
	wire new_net_6391;
	wire new_net_9669;
	wire new_net_19755;
	wire new_net_19791;
	wire new_net_13073;
	wire new_net_14221;
	wire new_net_18089;
	wire new_net_5310;
	wire new_net_8150;
	wire new_net_10482;
	wire new_net_1883;
	wire new_net_702;
	wire new_net_19144;
	wire new_net_19371;
	wire new_net_18054;
	wire new_net_19481;
	wire new_net_6148;
	wire new_net_10771;
	wire new_net_563;
	wire new_net_5279;
	wire new_net_18008;
	wire new_net_21451;
	wire new_net_16118;
	wire new_net_554;
	wire new_net_3775;
	wire new_net_8554;
	wire new_net_9672;
	wire new_net_20108;
	wire new_net_20735;
	wire new_net_13510;
	wire new_net_5888;
	wire new_net_10929;
	wire new_net_10696;
	wire new_net_10770;
	wire new_net_10389;
	wire new_net_1885;
	wire new_net_2064;
	wire new_net_98;
	wire new_net_709;
	wire new_net_11329;
	wire new_net_12851;
	wire new_net_1255;
	wire new_net_5314;
	wire new_net_9861;
	wire new_net_562;
	wire new_net_9674;
	wire new_net_6484;
	wire new_net_10585;
	wire new_net_3914;
	wire new_net_15612;
	wire new_net_17492;
	wire new_net_17741;
	wire new_net_17552;
	wire new_net_14052;
	wire new_net_16333;
	wire new_net_16618;
	wire new_net_13613;
	wire new_net_8054;
	wire new_net_12668;
	wire new_net_17130;
	wire new_net_15893;
	wire new_net_14928;
	wire new_net_4486;
	wire new_net_8861;
	wire new_net_94;
	wire new_net_2756;
	wire new_net_4115;
	wire new_net_19756;
	wire new_net_19792;
	wire new_net_16838;
	wire new_net_9099;
	wire new_net_1705;
	wire new_net_5281;
	wire new_net_7197;
	wire new_net_17966;
	wire new_net_19372;
	wire new_net_21066;
	wire new_net_16772;
	wire new_net_21115;
	wire new_net_10231;
	wire new_net_8645;
	wire new_net_9096;
	wire new_net_10385;
	wire new_net_176;
	wire new_net_4676;
	wire new_net_5283;
	wire new_net_19143;
	wire new_net_21452;
	wire new_net_13583;
	wire new_net_14651;
	wire new_net_8643;
	wire new_net_12615;
	wire new_net_1231;
	wire new_net_3754;
	wire new_net_10088;
	wire new_net_18869;
	wire new_net_20109;
	wire new_net_20736;
	wire new_net_17926;
	wire new_net_8644;
	wire new_net_16097;
	wire new_net_5309;
	wire new_net_6395;
	wire new_net_10930;
	wire new_net_8058;
	wire new_net_1235;
	wire new_net_421;
	wire new_net_4440;
	wire new_net_8560;
	wire new_net_18584;
	wire new_net_19085;
	wire new_net_6149;
	wire new_net_8642;
	wire new_net_9856;
	wire new_net_8223;
	wire new_net_701;
	wire new_net_155;
	wire new_net_6249;
	wire new_net_12253;
	wire new_net_15613;
	wire new_net_17493;
	wire new_net_17742;
	wire new_net_17553;
	wire new_net_14051;
	wire new_net_16334;
	wire new_net_16619;
	wire new_net_13614;
	wire new_net_12669;
	wire new_net_12290;
	wire new_net_423;
	wire new_net_699;
	wire new_net_18999;
	wire new_net_19757;
	wire new_net_19793;
	wire new_net_17580;
	wire new_net_15326;
	wire new_net_16785;
	wire new_net_17116;
	wire new_net_14241;
	wire new_net_6488;
	wire new_net_6140;
	wire new_net_5311;
	wire new_net_9865;
	wire new_net_10695;
	wire new_net_1236;
	wire new_net_3769;
	wire new_net_19373;
	wire new_net_12614;
	wire new_net_8870;
	wire new_net_9855;
	wire new_net_6392;
	wire new_net_6489;
	wire new_net_10702;
	wire new_net_21453;
	wire new_net_19142;
	wire new_net_20110;
	wire new_net_20737;
	wire new_net_20863;
	wire new_net_13686;
	wire new_net_2082;
	wire new_net_16545;
	wire new_net_20792;
	wire new_net_10931;
	wire new_net_10769;
	wire new_net_8053;
	wire new_net_6146;
	wire new_net_11331;
	wire new_net_20406;
	wire new_net_21368;
	wire new_net_17374;
	wire new_net_6494;
	wire new_net_10766;
	wire new_net_8216;
	wire new_net_97;
	wire new_net_14744;
	wire new_net_7786;
	wire new_net_18546;
	wire new_net_1158;
	wire new_net_11650;
	wire new_net_17411;
	wire new_net_15614;
	wire new_net_17494;
	wire new_net_17743;
	wire new_net_16098;
	wire new_net_17554;
	wire new_net_16335;
	wire new_net_16620;
	wire new_net_13615;
	wire new_net_12670;
	wire new_net_12291;
	wire new_net_14840;
	wire new_net_15880;
	wire new_net_14351;
	wire new_net_3770;
	wire new_net_19758;
	wire new_net_19794;
	wire new_net_6486;
	wire new_net_17736;
	wire new_net_6390;
	wire new_net_93;
	wire new_net_1234;
	wire new_net_18998;
	wire new_net_19374;
	wire new_net_5087;
	wire new_net_16110;
	wire new_net_8648;
	wire new_net_4114;
	wire new_net_8217;
	wire new_net_91;
	wire new_net_710;
	wire new_net_21454;
	wire new_net_13278;
	wire new_net_7203;
	wire new_net_6490;
	wire new_net_8865;
	wire new_net_9864;
	wire new_net_8221;
	wire new_net_16748;
	wire new_net_3686;
	wire new_net_4430;
	wire new_net_10384;
	wire new_net_20111;
	wire new_net_20273;
	wire new_net_12080;
	wire new_net_13602;
	wire new_net_13208;
	wire new_net_18820;
	wire new_net_7198;
	wire new_net_11332;
	wire new_net_12613;
	wire new_net_10932;
	wire new_net_424;
	wire new_net_9095;
	wire new_net_11416;
	wire new_net_12654;
	wire new_net_19141;
	wire new_net_20407;
	wire new_net_18355;
	wire new_net_13842;
	wire new_net_4155;
	wire new_net_12312;
	wire new_net_18624;
	wire new_net_14004;
	wire new_net_15332;
	wire new_net_15921;
	wire new_net_18251;
	wire new_net_17755;
	wire new_net_6707;
	wire new_net_5862;
	wire new_net_1522;
	wire new_net_2707;
	wire new_net_5743;
	wire new_net_8496;
	wire new_net_15369;
	wire new_net_1380;
	wire new_net_15958;
	wire new_net_16864;
	wire new_net_5182;
	wire new_net_13934;
	wire new_net_14311;
	wire new_net_15449;
	wire new_net_16774;
	wire new_net_17105;
	wire new_net_11939;
	wire new_net_13274;
	wire new_net_16668;
	wire new_net_11668;
	wire new_net_12541;
	wire new_net_7625;
	wire new_net_3893;
	wire new_net_8014;
	wire new_net_11948;
	wire new_net_14451;
	wire _1191_;
	wire new_net_934;
	wire new_net_1521;
	wire new_net_6353;
	wire new_net_6369;
	wire new_net_10183;
	wire new_net_11962;
	wire new_net_5746;
	wire new_net_16982;
	wire new_net_17812;
	wire new_net_4675;
	wire new_net_9491;
	wire _1192_;
	wire new_net_1021;
	wire new_net_2497;
	wire new_net_6042;
	wire new_net_6376;
	wire new_net_19262;
	wire new_net_20691;
	wire new_net_20930;
	wire new_net_17055;
	wire new_net_17884;
	wire new_net_18495;
	wire new_net_7762;
	wire new_net_16997;
	wire new_net_10793;
	wire new_net_10040;
	wire new_net_12992;
	wire new_net_10945;
	wire new_net_5861;
	wire new_net_7324;
	wire new_net_13556;
	wire new_net_1527;
	wire new_net_10093;
	wire new_net_12409;
	wire new_net_15185;
	wire new_net_17395;
	wire new_net_5216;
	wire new_net_5737;
	wire new_net_10041;
	wire _1193_;
	wire new_net_1665;
	wire new_net_2822;
	wire new_net_4751;
	wire new_net_15052;
	wire new_net_6260;
	wire new_net_13935;
	wire new_net_14312;
	wire new_net_15450;
	wire new_net_16775;
	wire new_net_17106;
	wire new_net_17092;
	wire new_net_11940;
	wire new_net_9489;
	wire new_net_13275;
	wire new_net_11669;
	wire new_net_20510;
	wire new_net_13074;
	wire new_net_14222;
	wire new_net_15402;
	wire new_net_18090;
	wire new_net_16025;
	wire new_net_5739;
	wire new_net_2714;
	wire new_net_17754;
	wire new_net_4454;
	wire new_net_9495;
	wire new_net_3532;
	wire new_net_6339;
	wire new_net_16469;
	wire _1194_;
	wire new_net_5499;
	wire new_net_18055;
	wire new_net_18009;
	wire new_net_16478;
	wire new_net_1526;
	wire new_net_2818;
	wire new_net_6375;
	wire new_net_19263;
	wire new_net_6243;
	wire new_net_9213;
	wire new_net_12707;
	wire new_net_11217;
	wire new_net_6706;
	wire new_net_6520;
	wire new_net_6334;
	wire _1195_;
	wire new_net_2817;
	wire new_net_5582;
	wire new_net_6050;
	wire new_net_3654;
	wire new_net_13511;
	wire new_net_5887;
	wire new_net_7305;
	wire new_net_939;
	wire new_net_3534;
	wire new_net_4750;
	wire new_net_20692;
	wire new_net_20931;
	wire new_net_6041;
	wire new_net_10794;
	wire new_net_4458;
	wire new_net_10946;
	wire new_net_16669;
	wire new_net_6341;
	wire new_net_2826;
	wire _1196_;
	wire new_net_1659;
	wire new_net_3535;
	wire new_net_12257;
	wire new_net_15835;
	wire new_net_15011;
	wire new_net_17091;
	wire new_net_2499;
	wire new_net_10099;
	wire new_net_4308;
	wire new_net_15894;
	wire new_net_14929;
	wire new_net_19279;
	wire new_net_12164;
	wire new_net_12406;
	wire new_net_14699;
	wire new_net_13936;
	wire new_net_14313;
	wire new_net_15451;
	wire new_net_16776;
	wire new_net_17107;
	wire new_net_16467;
	wire new_net_11941;
	wire new_net_19974;
	wire new_net_7471;
	wire new_net_16839;
	wire new_net_6587;
	wire new_net_17967;
	wire new_net_21067;
	wire new_net_5585;
	wire new_net_6047;
	wire new_net_17753;
	wire new_net_8984;
	wire new_net_4677;
	wire new_net_2824;
	wire new_net_12594;
	wire new_net_11511;
	wire new_net_16773;
	wire new_net_21116;
	wire new_net_10230;
	wire new_net_1023;
	wire _1198_;
	wire new_net_6344;
	wire new_net_16470;
	wire new_net_8502;
	wire new_net_10098;
	wire new_net_13584;
	wire new_net_14652;
	wire new_net_10079;
	wire new_net_18870;
	wire new_net_1907;
	wire new_net_3891;
	wire new_net_3993;
	wire new_net_5181;
	wire new_net_6343;
	wire new_net_6371;
	wire new_net_10097;
	wire new_net_17927;
	wire new_net_18585;
	wire new_net_3292;
	wire new_net_4680;
	wire _1199_;
	wire new_net_10094;
	wire new_net_20693;
	wire new_net_20932;
	wire new_net_15265;
	wire new_net_19086;
	wire new_net_11218;
	wire new_net_10947;
	wire new_net_3400;
	wire new_net_3889;
	wire new_net_4456;
	wire new_net_20434;
	wire new_net_12254;
	wire new_net_15010;
	wire new_net_6712;
	wire _1200_;
	wire new_net_17090;
	wire new_net_8505;
	wire new_net_6290;
	wire new_net_5255;
	wire new_net_5583;
	wire new_net_12165;
	wire new_net_12405;
	wire new_net_14700;
	wire new_net_13937;
	wire new_net_14314;
	wire new_net_15452;
	wire new_net_16777;
	wire new_net_17108;
	wire new_net_11942;
	wire new_net_17581;
	wire new_net_15327;
	wire new_net_14242;
	wire new_net_17752;
	wire new_net_1020;
	wire new_net_2493;
	wire _1201_;
	wire new_net_4753;
	wire new_net_18049;
	wire new_net_20834;
	wire new_net_16609;
	wire new_net_4601;
	wire new_net_9493;
	wire new_net_938;
	wire new_net_1024;
	wire new_net_1524;
	wire new_net_6046;
	wire new_net_16477;
	wire new_net_10095;
	wire new_net_14468;
	wire new_net_11182;
	wire new_net_16557;
	wire new_net_8007;
	wire new_net_5180;
	wire new_net_5741;
	wire new_net_10795;
	wire new_net_6519;
	wire new_net_9492;
	wire _1202_;
	wire new_net_2819;
	wire new_net_6335;
	wire new_net_4756;
	wire new_net_2080;
	wire new_net_16546;
	wire new_net_5579;
	wire new_net_5745;
	wire new_net_6714;
	wire new_net_3994;
	wire new_net_5864;
	wire new_net_20694;
	wire _1190_;
	wire new_net_12386;
	wire new_net_15782;
	wire new_net_18383;
	wire new_net_17375;
	wire new_net_14745;
	wire new_net_5186;
	wire new_net_11219;
	wire new_net_10948;
	wire new_net_2703;
	wire _1203_;
	wire new_net_20435;
	wire new_net_18547;
	wire new_net_9963;
	wire new_net_11651;
	wire new_net_15009;
	wire new_net_6708;
	wire new_net_7481;
	wire new_net_932;
	wire new_net_2702;
	wire new_net_17089;
	wire new_net_8506;
	wire new_net_14841;
	wire new_net_15881;
	wire new_net_14352;
	wire new_net_12404;
	wire new_net_13551;
	wire new_net_8009;
	wire new_net_13938;
	wire new_net_17109;
	wire new_net_14315;
	wire new_net_15453;
	wire new_net_13513;
	wire new_net_8816;
	wire new_net_11943;
	wire new_net_15608;
	wire new_net_17737;
	wire new_net_17470;
	wire new_net_17751;
	wire new_net_9571;
	wire new_net_1525;
	wire new_net_2494;
	wire new_net_6336;
	wire new_net_6374;
	wire _0504_;
	wire new_net_10186;
	wire new_net_2705;
	wire new_net_10827;
	wire new_net_1657;
	wire _1205_;
	wire new_net_1022;
	wire new_net_1911;
	wire new_net_2491;
	wire new_net_13279;
	wire new_net_16749;
	wire new_net_8978;
	wire new_net_2815;
	wire new_net_4673;
	wire new_net_4755;
	wire new_net_12081;
	wire new_net_13601;
	wire new_net_13209;
	wire new_net_2104;
	wire new_net_18821;
	wire new_net_15705;
	wire new_net_12655;
	wire new_net_13293;
	wire _1206_;
	wire new_net_2712;
	wire new_net_3896;
	wire new_net_20695;
	wire new_net_10146;
	wire new_net_18356;
	wire new_net_13843;
	wire new_net_11220;
	wire new_net_10796;
	wire new_net_10949;
	wire new_net_1915;
	wire new_net_2492;
	wire new_net_2715;
	wire new_net_5184;
	wire new_net_5740;
	wire new_net_12313;
	wire new_net_19264;
	wire new_net_18625;
	wire new_net_14005;
	wire new_net_10089;
	wire new_net_15008;
	wire _1207_;
	wire new_net_1529;
	wire new_net_2496;
	wire new_net_2821;
	wire new_net_17088;
	wire new_net_15333;
	wire new_net_15922;
	wire new_net_18252;
	wire new_net_6272;
	wire new_net_15370;
	wire new_net_12391;
	wire new_net_13808;
	wire new_net_10185;
	wire new_net_12167;
	wire new_net_12403;
	wire new_net_14702;
	wire new_net_13939;
	wire new_net_14316;
	wire new_net_15454;
	wire new_net_16779;
	wire new_net_16865;
	wire new_net_5183;
	wire new_net_17750;
	wire new_net_8985;
	wire new_net_4674;
	wire new_net_17567;
	wire _1208_;
	wire new_net_1016;
	wire new_net_3538;
	wire new_net_16471;
	wire new_net_11949;
	wire new_net_6890;
	wire new_net_3290;
	wire new_net_7478;
	wire new_net_16476;
	wire new_net_14452;
	wire new_net_20164;
	wire new_net_8980;
	wire _1209_;
	wire new_net_4154;
	wire new_net_16983;
	wire new_net_17813;
	wire new_net_8497;
	wire new_net_6373;
	wire new_net_1660;
	wire new_net_2825;
	wire new_net_2708;
	wire new_net_8817;
	wire new_net_20696;
	wire new_net_16235;
	wire new_net_8079;
	wire new_net_17056;
	wire new_net_17885;
	wire new_net_8778;
	wire new_net_18496;
	wire new_net_10797;
	wire new_net_936;
	wire new_net_11221;
	wire new_net_10950;
	wire new_net_3989;
	wire _1210_;
	wire new_net_20437;
	wire new_net_15186;
	wire new_net_17396;
	wire new_net_17087;
	wire new_net_8986;
	wire new_net_5742;
	wire new_net_15485;
	wire new_net_15053;
	wire new_net_16780;
	wire new_net_12392;
	wire new_net_15788;
	wire new_net_16673;
	wire new_net_12168;
	wire new_net_12402;
	wire new_net_13940;
	wire new_net_15455;
	wire new_net_14317;
	wire new_net_13809;
	wire new_net_8617;
	wire new_net_5813;
	wire new_net_13075;
	wire new_net_14223;
	wire new_net_8503;
	wire new_net_10092;
	wire new_net_15007;
	wire new_net_17749;
	wire new_net_3992;
	wire new_net_18091;
	wire new_net_16026;
	wire new_net_18056;
	wire _1212_;
	wire new_net_1661;
	wire new_net_3894;
	wire new_net_11820;
	wire new_net_18010;
	wire new_net_16120;
	wire new_net_12708;
	wire new_net_18612;
	wire new_net_8012;
	wire new_net_5736;
	wire new_net_7485;
	wire new_net_13512;
	wire new_net_7304;
	wire new_net_3892;
	wire new_net_3988;
	wire new_net_5865;
	wire new_net_16468;
	wire new_net_5738;
	wire new_net_1913;
	wire _1213_;
	wire new_net_9488;
	wire new_net_20697;
	wire new_net_12853;
	wire new_net_12139;
	wire new_net_11222;
	wire new_net_10798;
	wire new_net_1912;
	wire new_net_1015;
	wire new_net_5860;
	wire new_net_10951;
	wire new_net_20438;
	wire new_net_12258;
	wire new_net_15836;
	wire new_net_6337;
	wire new_net_17086;
	wire new_net_6704;
	wire new_net_8979;
	wire new_net_4453;
	wire new_net_4679;
	wire new_net_1914;
	wire _1214_;
	wire new_net_6563;
	wire new_net_17132;
	wire new_net_15895;
	wire new_net_17112;
	wire new_net_11675;
	wire new_net_13516;
	wire new_net_5500;
	wire new_net_12393;
	wire new_net_12401;
	wire new_net_16781;
	wire new_net_6045;
	wire new_net_12169;
	wire new_net_13941;
	wire new_net_14930;
	wire new_net_4752;
	wire new_net_17748;
	wire new_net_8976;
	wire new_net_4452;
	wire new_net_2820;
	wire _1215_;
	wire new_net_2500;
	wire new_net_16840;
	wire new_net_17968;
	wire new_net_21068;
	wire new_net_12595;
	wire new_net_16475;
	wire new_net_1531;
	wire new_net_2706;
	wire new_net_5673;
	wire new_net_13585;
	wire new_net_14653;
	wire new_net_8982;
	wire new_net_6044;
	wire new_net_10182;
	wire _1216_;
	wire new_net_6523;
	wire new_net_6562;
	wire new_net_13668;
	wire new_net_18871;
	wire new_net_17928;
	wire new_net_18269;
	wire new_net_10042;
	wire new_net_1523;
	wire new_net_3288;
	wire new_net_3397;
	wire new_net_6372;
	wire new_net_6524;
	wire new_net_20698;
	wire new_net_18586;
	wire new_net_19479;
	wire new_net_15266;
	wire new_net_19087;
	wire new_net_3539;
	wire new_net_11223;
	wire new_net_10799;
	wire new_net_6705;
	wire _1217_;
	wire new_net_1656;
	wire new_net_10952;
	wire new_net_20439;
	wire new_net_6250;
	wire new_net_15242;
	wire new_net_12255;
	wire new_net_17085;
	wire new_net_15006;
	wire new_net_4757;
	wire new_net_5858;
	wire new_net_6518;
	wire new_net_15096;
	wire new_net_10328;
	wire new_net_11676;
	wire new_net_13517;
	wire new_net_13547;
	wire new_net_16472;
	wire new_net_12394;
	wire new_net_13811;
	wire new_net_15790;
	wire new_net_12170;
	wire new_net_12400;
	wire new_net_14705;
	wire new_net_17582;
	wire new_net_15328;
	wire new_net_14243;
	wire new_net_8501;
	wire new_net_5586;
	wire new_net_17747;
	wire new_net_2489;
	wire new_net_4451;
	wire new_net_7827;
	wire new_net_7477;
	wire new_net_13094;
	wire new_net_18076;
	wire new_net_21141;
	wire new_net_20163;
	wire new_net_6368;
	wire _1219_;
	wire new_net_6525;
	wire new_net_7479;
	wire new_net_19265;
	wire new_net_6404;
	wire new_net_14469;
	wire new_net_8006;
	wire new_net_1910;
	wire new_net_3533;
	wire new_net_5581;
	wire new_net_6561;
	wire new_net_11183;
	wire new_net_16558;
	wire new_net_20865;
	wire new_net_16547;
	wire _1220_;
	wire new_net_10187;
	wire new_net_5185;
	wire new_net_10038;
	wire new_net_20699;
	wire new_net_12387;
	wire new_net_15783;
	wire new_net_18384;
	wire new_net_17376;
	wire new_net_18434;
	wire new_net_11224;
	wire new_net_10800;
	wire new_net_4831;
	wire new_net_7325;
	wire new_net_10044;
	wire new_net_10953;
	wire new_net_20440;
	wire new_net_14746;
	wire new_net_11652;
	wire new_net_3895;
	wire new_net_17084;
	wire new_net_5584;
	wire new_net_15005;
	wire new_net_6710;
	wire new_net_2823;
	wire _1221_;
	wire new_net_1655;
	wire new_net_3536;
	wire new_net_9570;
	wire new_net_14865;
	wire new_net_15549;
	wire new_net_5605;
	wire new_net_16891;
	wire new_net_15882;
	wire new_net_14353;
	wire new_net_13283;
	wire new_net_12395;
	wire new_net_13812;
	wire new_net_12171;
	wire new_net_12399;
	wire new_net_13546;
	wire new_net_14706;
	wire new_net_13943;
	wire new_net_17114;
	wire new_net_14320;
	wire new_net_15609;
	wire new_net_17738;
	wire new_net_17471;
	wire new_net_7217;
	wire new_net_9494;
	wire new_net_6342;
	wire new_net_8818;
	wire new_net_5179;
	wire new_net_6711;
	wire _1222_;
	wire new_net_17746;
	wire new_net_16474;
	wire new_net_6040;
	wire new_net_6713;
	wire _1223_;
	wire new_net_13280;
	wire new_net_10195;
	wire new_net_16750;
	wire new_net_12082;
	wire new_net_13600;
	wire new_net_13210;
	wire new_net_2711;
	wire new_net_8010;
	wire new_net_20700;
	wire new_net_18822;
	wire new_net_12656;
	wire new_net_13294;
	wire new_net_15706;
	wire new_net_18307;
	wire new_net_18357;
	wire new_net_6526;
	wire new_net_7534;
	wire new_net_10954;
	wire new_net_15791;
	wire new_net_6377;
	wire new_net_11225;
	wire new_net_10801;
	wire _1224_;
	wire new_net_20441;
	wire new_net_13844;
	wire new_net_12314;
	wire new_net_18626;
	wire new_net_5859;
	wire new_net_6340;
	wire new_net_15004;
	wire new_net_17083;
	wire new_net_8983;
	wire new_net_2488;
	wire new_net_4832;
	wire new_net_14006;
	wire new_net_15334;
	wire new_net_15301;
	wire new_net_15371;
	wire new_net_6564;
	wire new_net_13284;
	wire new_net_16677;
	wire new_net_5857;
	wire new_net_11678;
	wire new_net_13519;
	wire new_net_13545;
	wire new_net_12396;
	wire new_net_13813;
	wire new_net_12172;
	wire new_net_16866;
	wire new_net_15983;
	wire new_net_17745;
	wire new_net_3890;
	wire new_net_6370;
	wire new_net_17568;
	wire new_net_11950;
	wire new_net_6788;
	wire new_net_17744;
	wire _1226_;
	wire new_net_1909;
	wire new_net_2498;
	wire new_net_14453;
	wire new_net_8500;
	wire new_net_935;
	wire new_net_16984;
	wire new_net_8011;
	wire new_net_10189;
	wire new_net_937;
	wire _1227_;
	wire new_net_6871;
	wire new_net_2501;
	wire new_net_2827;
	wire new_net_20701;
	wire new_net_17814;
	wire new_net_16236;
	wire new_net_10955;
	wire new_net_17081;
	wire new_net_15002;
	wire new_net_11226;
	wire new_net_10802;
	wire new_net_1019;
	wire new_net_4678;
	wire new_net_20442;
	wire new_net_1044;
	wire new_net_18497;
	wire new_net_15187;
	wire new_net_17397;
	wire new_net_7482;
	wire new_net_5866;
	wire new_net_6338;
	wire new_net_17082;
	wire new_net_6039;
	wire new_net_8815;
	wire new_net_15003;
	wire new_net_1662;
	wire _1228_;
	wire new_net_14873;
	wire new_net_17625;
	wire new_net_15486;
	wire new_net_15054;
	wire new_net_19714;
	wire new_net_13285;
	wire new_net_16678;
	wire new_net_5863;
	wire new_net_11679;
	wire new_net_13520;
	wire new_net_10090;
	wire new_net_12397;
	wire new_net_13814;
	wire new_net_15792;
	wire new_net_8013;
	wire new_net_13076;
	wire new_net_14224;
	wire new_net_3990;
	wire new_net_4754;
	wire new_net_10091;
	wire new_net_6043;
	wire new_net_2710;
	wire _1229_;
	wire new_net_933;
	wire new_net_1530;
	wire new_net_18092;
	wire new_net_16027;
	wire new_net_14180;
	wire new_net_18057;
	wire new_net_16473;
	wire new_net_8498;
	wire new_net_11821;
	wire new_net_18011;
	wire new_net_16121;
	wire new_net_5788;
	wire new_net_12709;
	wire new_net_6521;
	wire _1230_;
	wire new_net_4450;
	wire new_net_6709;
	wire new_net_10043;
	wire new_net_9490;
	wire new_net_8008;
	wire new_net_7483;
	wire new_net_20702;
	wire new_net_17898;
	wire new_net_12854;
	wire new_net_12140;
	wire new_net_10956;
	wire new_net_11227;
	wire new_net_10803;
	wire new_net_1025;
	wire new_net_2713;
	wire _0791_;
	wire _1231_;
	wire new_net_1658;
	wire new_net_19126;
	wire new_net_20443;
	wire new_net_12259;
	wire new_net_15837;
	wire new_net_17133;
	wire new_net_15896;
	wire new_net_14931;
	wire new_net_6599;
	wire new_net_9415;
	wire new_net_10219;
	wire new_net_10534;
	wire new_net_7549;
	wire new_net_2928;
	wire new_net_785;
	wire new_net_2632;
	wire new_net_6281;
	wire new_net_19976;
	wire new_net_16841;
	wire new_net_17708;
	wire new_net_9416;
	wire new_net_16396;
	wire new_net_16727;
	wire new_net_10214;
	wire new_net_13474;
	wire new_net_13993;
	wire new_net_17637;
	wire new_net_15060;
	wire new_net_16078;
	wire new_net_12596;
	wire new_net_20041;
	wire new_net_3315;
	wire new_net_20196;
	wire new_net_4448;
	wire new_net_3279;
	wire new_net_14402;
	wire new_net_14654;
	wire new_net_9565;
	wire new_net_8480;
	wire new_net_10218;
	wire new_net_6701;
	wire _0981_;
	wire _0141_;
	wire _0561_;
	wire new_net_18872;
	wire new_net_21349;
	wire new_net_17929;
	wire new_net_9249;
	wire new_net_2920;
	wire new_net_18587;
	wire new_net_7215;
	wire new_net_19088;
	wire new_net_10215;
	wire new_net_197;
	wire _0142_;
	wire _0562_;
	wire new_net_15142;
	wire _0982_;
	wire new_net_6070;
	wire new_net_2911;
	wire new_net_20918;
	wire new_net_9750;
	wire new_net_15243;
	wire new_net_12256;
	wire new_net_10980;
	wire new_net_4282;
	wire new_net_782;
	wire new_net_12610;
	wire new_net_19280;
	wire new_net_19575;
	wire new_net_15097;
	wire new_net_788;
	wire new_net_9112;
	wire new_net_4279;
	wire _0143_;
	wire _0563_;
	wire _0983_;
	wire new_net_20453;
	wire new_net_15329;
	wire new_net_6389;
	wire new_net_13120;
	wire new_net_6169;
	wire new_net_14244;
	wire new_net_16397;
	wire new_net_16728;
	wire new_net_9253;
	wire new_net_13676;
	wire new_net_13475;
	wire new_net_17804;
	wire new_net_12270;
	wire new_net_12957;
	wire new_net_15061;
	wire new_net_13982;
	wire new_net_7835;
	wire new_net_10023;
	wire new_net_13093;
	wire new_net_18077;
	wire new_net_21142;
	wire new_net_16611;
	wire new_net_9413;
	wire new_net_3719;
	wire _0984_;
	wire _0144_;
	wire _0564_;
	wire new_net_2549;
	wire new_net_20197;
	wire new_net_14470;
	wire new_net_9251;
	wire new_net_10536;
	wire new_net_5656;
	wire new_net_2565;
	wire new_net_16559;
	wire new_net_20866;
	wire new_net_21350;
	wire new_net_18360;
	wire new_net_16548;
	wire _0985_;
	wire new_net_192;
	wire _0145_;
	wire _0565_;
	wire new_net_2635;
	wire _1197_;
	wire new_net_12388;
	wire new_net_15784;
	wire new_net_18385;
	wire new_net_3707;
	wire new_net_20919;
	wire new_net_14747;
	wire new_net_8848;
	wire new_net_11653;
	wire new_net_12611;
	wire new_net_5304;
	wire new_net_5950;
	wire new_net_9250;
	wire new_net_13994;
	wire new_net_10981;
	wire new_net_10561;
	wire new_net_2553;
	wire new_net_190;
	wire _0566_;
	wire new_net_14866;
	wire new_net_15550;
	wire new_net_17226;
	wire new_net_16892;
	wire new_net_14843;
	wire new_net_15883;
	wire new_net_14354;
	wire new_net_12607;
	wire new_net_9414;
	wire new_net_20454;
	wire new_net_15610;
	wire new_net_17739;
	wire new_net_10150;
	wire new_net_11858;
	wire new_net_16080;
	wire new_net_16398;
	wire new_net_16729;
	wire new_net_17639;
	wire new_net_17131;
	wire new_net_13677;
	wire new_net_13476;
	wire new_net_17805;
	wire new_net_4594;
	wire new_net_8108;
	wire _0511_;
	wire new_net_10790;
	wire new_net_5954;
	wire new_net_2560;
	wire new_net_2628;
	wire new_net_2912;
	wire new_net_20198;
	wire new_net_862;
	wire new_net_10726;
	wire new_net_13374;
	wire new_net_11523;
	wire new_net_13281;
	wire new_net_5953;
	wire new_net_9255;
	wire new_net_10216;
	wire _0148_;
	wire _0568_;
	wire _0988_;
	wire new_net_21351;
	wire new_net_20276;
	wire new_net_12083;
	wire new_net_13599;
	wire new_net_13211;
	wire new_net_11442;
	wire new_net_8477;
	wire new_net_18823;
	wire new_net_7442;
	wire new_net_10557;
	wire new_net_2551;
	wire new_net_13295;
	wire new_net_5046;
	wire new_net_18358;
	wire new_net_9117;
	wire new_net_9252;
	wire new_net_6686;
	wire new_net_6797;
	wire _0569_;
	wire new_net_787;
	wire _0149_;
	wire _0989_;
	wire new_net_188;
	wire new_net_12315;
	wire new_net_19879;
	wire new_net_10886;
	wire new_net_18627;
	wire new_net_6596;
	wire new_net_10982;
	wire new_net_6798;
	wire new_net_6289;
	wire new_net_7209;
	wire new_net_10560;
	wire new_net_791;
	wire new_net_4284;
	wire new_net_5661;
	wire new_net_8314;
	wire new_net_14007;
	wire new_net_147;
	wire new_net_15372;
	wire new_net_3319;
	wire new_net_3710;
	wire new_net_2634;
	wire _0570_;
	wire _0990_;
	wire _0150_;
	wire new_net_7545;
	wire new_net_20455;
	wire new_net_16867;
	wire new_net_20529;
	wire new_net_15984;
	wire new_net_7310;
	wire new_net_11859;
	wire new_net_16399;
	wire new_net_16730;
	wire new_net_13678;
	wire new_net_13477;
	wire new_net_17806;
	wire new_net_12272;
	wire new_net_12959;
	wire new_net_13995;
	wire new_net_15063;
	wire new_net_3834;
	wire new_net_4384;
	wire new_net_12609;
	wire new_net_3706;
	wire new_net_5306;
	wire new_net_3721;
	wire new_net_10558;
	wire _0571_;
	wire _0991_;
	wire _0151_;
	wire new_net_20199;
	wire new_net_14454;
	wire new_net_8622;
	wire new_net_3430;
	wire new_net_21352;
	wire new_net_16985;
	wire new_net_6280;
	wire new_net_7207;
	wire new_net_789;
	wire _0572_;
	wire _0992_;
	wire _0152_;
	wire new_net_6702;
	wire new_net_16237;
	wire new_net_10539;
	wire new_net_2918;
	wire new_net_196;
	wire new_net_4596;
	wire new_net_6700;
	wire new_net_18498;
	wire new_net_20921;
	wire new_net_12408;
	wire new_net_14697;
	wire new_net_15188;
	wire new_net_17398;
	wire new_net_5305;
	wire new_net_10983;
	wire new_net_4590;
	wire _0993_;
	wire _0573_;
	wire new_net_2919;
	wire _0153_;
	wire new_net_756;
	wire new_net_19578;
	wire new_net_15487;
	wire new_net_15055;
	wire new_net_20215;
	wire new_net_3422;
	wire new_net_3708;
	wire new_net_6605;
	wire new_net_20456;
	wire new_net_9684;
	wire new_net_13077;
	wire new_net_14225;
	wire new_net_15419;
	wire new_net_17641;
	wire new_net_11860;
	wire new_net_16400;
	wire new_net_16731;
	wire new_net_13679;
	wire new_net_13478;
	wire new_net_17807;
	wire new_net_11856;
	wire new_net_12960;
	wire new_net_18093;
	wire new_net_16028;
	wire new_net_14181;
	wire new_net_18058;
	wire new_net_6600;
	wire new_net_10222;
	wire new_net_4592;
	wire new_net_8049;
	wire new_net_3411;
	wire new_net_20200;
	wire new_net_11822;
	wire new_net_18012;
	wire new_net_12710;
	wire new_net_6601;
	wire new_net_3408;
	wire new_net_4281;
	wire new_net_191;
	wire _0575_;
	wire _0995_;
	wire _0155_;
	wire new_net_19281;
	wire new_net_21353;
	wire new_net_3314;
	wire new_net_6819;
	wire new_net_11987;
	wire new_net_13514;
	wire new_net_9417;
	wire new_net_10789;
	wire new_net_2916;
	wire new_net_17899;
	wire new_net_12855;
	wire new_net_12141;
	wire new_net_7439;
	wire new_net_4309;
	wire _0156_;
	wire new_net_2559;
	wire new_net_2638;
	wire _0576_;
	wire _0996_;
	wire new_net_20922;
	wire new_net_12260;
	wire new_net_12608;
	wire new_net_16081;
	wire new_net_7446;
	wire new_net_9118;
	wire new_net_10984;
	wire new_net_2550;
	wire new_net_19282;
	wire new_net_19579;
	wire new_net_15426;
	wire new_net_17134;
	wire new_net_15897;
	wire new_net_5658;
	wire new_net_7551;
	wire _0157_;
	wire new_net_7444;
	wire new_net_10781;
	wire new_net_781;
	wire _0577_;
	wire _0997_;
	wire new_net_14932;
	wire new_net_20457;
	wire new_net_15420;
	wire new_net_17642;
	wire new_net_11861;
	wire new_net_16401;
	wire new_net_16732;
	wire new_net_15065;
	wire new_net_13680;
	wire new_net_13479;
	wire new_net_17808;
	wire new_net_12961;
	wire new_net_16842;
	wire new_net_6703;
	wire new_net_7437;
	wire new_net_6796;
	wire _0998_;
	wire _0158_;
	wire _0578_;
	wire new_net_10005;
	wire new_net_20201;
	wire new_net_4457;
	wire new_net_8395;
	wire new_net_14403;
	wire new_net_14655;
	wire new_net_8838;
	wire new_net_19125;
	wire new_net_4285;
	wire new_net_6286;
	wire new_net_10004;
	wire new_net_21354;
	wire new_net_13670;
	wire new_net_18873;
	wire new_net_17930;
	wire new_net_7550;
	wire new_net_10223;
	wire _0579_;
	wire _0999_;
	wire _0159_;
	wire new_net_2633;
	wire new_net_6288;
	wire new_net_18588;
	wire new_net_8693;
	wire new_net_19089;
	wire new_net_12606;
	wire new_net_10221;
	wire new_net_4283;
	wire new_net_8046;
	wire new_net_10008;
	wire new_net_10562;
	wire new_net_20923;
	wire new_net_15143;
	wire new_net_9591;
	wire new_net_2913;
	wire new_net_10985;
	wire new_net_4286;
	wire new_net_4595;
	wire new_net_193;
	wire _0580_;
	wire _1000_;
	wire _0160_;
	wire new_net_2557;
	wire new_net_3720;
	wire new_net_15098;
	wire new_net_10788;
	wire new_net_12273;
	wire new_net_2914;
	wire new_net_1473;
	wire new_net_7210;
	wire new_net_19283;
	wire new_net_20458;
	wire new_net_15330;
	wire new_net_15421;
	wire new_net_11862;
	wire new_net_16082;
	wire new_net_9421;
	wire new_net_16402;
	wire new_net_16733;
	wire new_net_3711;
	wire new_net_5951;
	wire new_net_13681;
	wire new_net_6457;
	wire new_net_13092;
	wire new_net_18078;
	wire new_net_21143;
	wire new_net_7547;
	wire new_net_10217;
	wire new_net_199;
	wire new_net_5176;
	wire new_net_20202;
	wire new_net_7438;
	wire new_net_9113;
	wire _1002_;
	wire _0162_;
	wire _0582_;
	wire new_net_13227;
	wire new_net_21355;
	wire new_net_16560;
	wire new_net_18361;
	wire new_net_16549;
	wire new_net_20796;
	wire new_net_7208;
	wire new_net_5663;
	wire new_net_2925;
	wire new_net_189;
	wire new_net_20348;
	wire new_net_12389;
	wire new_net_15785;
	wire new_net_18386;
	wire new_net_5175;
	wire new_net_6602;
	wire new_net_9419;
	wire _0163_;
	wire _0583_;
	wire _1003_;
	wire new_net_20924;
	wire new_net_14748;
	wire new_net_13815;
	wire new_net_11654;
	wire new_net_17643;
	wire new_net_10415;
	wire new_net_10986;
	wire new_net_4591;
	wire new_net_2563;
	wire new_net_198;
	wire new_net_4312;
	wire new_net_19581;
	wire new_net_6541;
	wire new_net_14867;
	wire new_net_16893;
	wire new_net_14844;
	wire new_net_15884;
	wire new_net_12604;
	wire new_net_10782;
	wire _1004_;
	wire new_net_790;
	wire new_net_2556;
	wire _0164_;
	wire _0584_;
	wire new_net_20459;
	wire new_net_15611;
	wire new_net_17740;
	wire new_net_13988;
	wire new_net_15516;
	wire new_net_17136;
	wire new_net_17715;
	wire new_net_15422;
	wire new_net_11863;
	wire new_net_16083;
	wire new_net_9424;
	wire new_net_16403;
	wire new_net_16734;
	wire new_net_783;
	wire _0165_;
	wire _0585_;
	wire _1005_;
	wire new_net_20203;
	wire new_net_13375;
	wire new_net_9120;
	wire new_net_12274;
	wire new_net_5659;
	wire new_net_5955;
	wire new_net_13282;
	wire new_net_12084;
	wire new_net_13598;
	wire new_net_13212;
	wire new_net_11443;
	wire new_net_7552;
	wire new_net_9422;
	wire new_net_9256;
	wire new_net_6688;
	wire new_net_4593;
	wire _0586_;
	wire _1006_;
	wire _0166_;
	wire new_net_18824;
	wire new_net_12658;
	wire new_net_13296;
	wire new_net_15708;
	wire new_net_18359;
	wire new_net_20925;
	wire new_net_4032;
	wire new_net_13846;
	wire new_net_8740;
	wire new_net_18628;
	wire new_net_4313;
	wire new_net_3709;
	wire new_net_9254;
	wire new_net_10987;
	wire new_net_10535;
	wire new_net_8047;
	wire new_net_2562;
	wire _0587_;
	wire _1007_;
	wire _0167_;
	wire new_net_14008;
	wire new_net_15336;
	wire new_net_15373;
	wire new_net_12605;
	wire new_net_9119;
	wire new_net_2564;
	wire new_net_20460;
	wire new_net_4035;
	wire new_net_16868;
	wire new_net_15985;
	wire new_net_4307;
	wire new_net_13989;
	wire new_net_15517;
	wire new_net_17137;
	wire new_net_17716;
	wire new_net_17644;
	wire new_net_11864;
	wire new_net_16084;
	wire new_net_9423;
	wire new_net_16404;
	wire new_net_17570;
	wire new_net_19344;
	wire new_net_10414;
	wire new_net_12602;
	wire new_net_784;
	wire new_net_3316;
	wire new_net_20204;
	wire _0797_;
	wire new_net_14455;
	wire new_net_8623;
	wire new_net_6285;
	wire new_net_6598;
	wire new_net_7443;
	wire new_net_12275;
	wire _0169_;
	wire _0589_;
	wire _1009_;
	wire new_net_8832;
	wire new_net_12603;
	wire new_net_9420;
	wire new_net_9116;
	wire new_net_6799;
	wire new_net_11274;
	wire new_net_15299;
	wire new_net_16238;
	wire new_net_5946;
	wire new_net_10533;
	wire _0590_;
	wire _0170_;
	wire _1010_;
	wire new_net_194;
	wire new_net_20926;
	wire new_net_18499;
	wire new_net_12407;
	wire new_net_14698;
	wire new_net_15189;
	wire new_net_17399;
	wire new_net_15423;
	wire new_net_10988;
	wire new_net_13482;
	wire new_net_2636;
	wire new_net_19583;
	wire new_net_14875;
	wire new_net_17627;
	wire new_net_15488;
	wire new_net_15056;
	wire new_net_10783;
	wire new_net_5952;
	wire new_net_6687;
	wire new_net_2555;
	wire _0591_;
	wire _1011_;
	wire _0171_;
	wire new_net_20461;
	wire new_net_7461;
	wire new_net_14226;
	wire new_net_7418;
	wire new_net_12965;
	wire new_net_14001;
	wire new_net_15069;
	wire new_net_13990;
	wire new_net_15518;
	wire new_net_17138;
	wire new_net_17717;
	wire new_net_17645;
	wire new_net_11865;
	wire new_net_10413;
	wire new_net_11857;
	wire new_net_18094;
	wire new_net_16029;
	wire new_net_14182;
	wire new_net_18059;
	wire new_net_10564;
	wire new_net_5662;
	wire _0592_;
	wire _1012_;
	wire _0172_;
	wire new_net_20205;
	wire new_net_11823;
	wire new_net_18013;
	wire new_net_10007;
	wire new_net_12276;
	wire new_net_7416;
	wire new_net_12101;
	wire new_net_6055;
	wire new_net_11988;
	wire new_net_3722;
	wire new_net_6279;
	wire new_net_10785;
	wire new_net_13515;
	wire new_net_10540;
	wire new_net_2924;
	wire _0593_;
	wire _1013_;
	wire _0173_;
	wire new_net_21356;
	wire new_net_12211;
	wire new_net_17900;
	wire new_net_12856;
	wire new_net_11465;
	wire new_net_5664;
	wire new_net_9418;
	wire new_net_10786;
	wire new_net_5948;
	wire new_net_12142;
	wire new_net_2631;
	wire new_net_20927;
	wire _0798_;
	wire new_net_12261;
	wire new_net_6287;
	wire new_net_10784;
	wire new_net_10989;
	wire _1014_;
	wire new_net_410;
	wire _0594_;
	wire new_net_2558;
	wire _0174_;
	wire new_net_19584;
	wire new_net_15839;
	wire new_net_15427;
	wire new_net_17135;
	wire new_net_7204;
	wire new_net_15898;
	wire new_net_6597;
	wire new_net_10787;
	wire new_net_6800;
	wire new_net_792;
	wire new_net_2922;
	wire new_net_4311;
	wire new_net_20462;
	wire new_net_19978;
	wire new_net_12966;
	wire new_net_14002;
	wire new_net_15070;
	wire new_net_13991;
	wire new_net_15519;
	wire new_net_17139;
	wire new_net_15424;
	wire new_net_17646;
	wire _0175_;
	wire new_net_11866;
	wire new_net_16843;
	wire new_net_12598;
	wire new_net_7417;
	wire new_net_10538;
	wire new_net_7445;
	wire new_net_9115;
	wire new_net_10220;
	wire new_net_20206;
	wire new_net_4449;
	wire new_net_14404;
	wire new_net_14656;
	wire new_net_13587;
	wire new_net_12277;
	wire new_net_4277;
	wire new_net_2629;
	wire _0596_;
	wire _1016_;
	wire _0176_;
	wire new_net_3705;
	wire new_net_13671;
	wire new_net_18874;
	wire new_net_10559;
	wire new_net_21357;
	wire new_net_17931;
	wire new_net_18589;
	wire new_net_5177;
	wire _0177_;
	wire new_net_2915;
	wire _0597_;
	wire _1017_;
	wire new_net_19284;
	wire new_net_7709;
	wire new_net_20928;
	wire new_net_12279;
	wire new_net_19090;
	wire new_net_15144;
	wire new_net_12600;
	wire new_net_10990;
	wire new_net_19585;
	wire new_net_5464;
	wire new_net_15245;
	wire new_net_15099;
	wire new_net_2926;
	wire _0598_;
	wire _1018_;
	wire _0178_;
	wire new_net_18100;
	wire new_net_20463;
	wire new_net_10326;
	wire new_net_17584;
	wire new_net_15331;
	wire new_net_12967;
	wire new_net_14003;
	wire new_net_15071;
	wire new_net_13992;
	wire new_net_15520;
	wire new_net_15425;
	wire new_net_17647;
	wire new_net_17719;
	wire new_net_11867;
	wire new_net_16087;
	wire new_net_13122;
	wire new_net_14246;
	wire new_net_13091;
	wire new_net_18079;
	wire new_net_21144;
	wire new_net_2917;
	wire new_net_10780;
	wire _1019_;
	wire _0179_;
	wire _0599_;
	wire new_net_2552;
	wire new_net_20207;
	wire new_net_16613;
	wire new_net_14472;
	wire new_net_12278;
	wire new_net_12601;
	wire new_net_4310;
	wire new_net_13228;
	wire new_net_16561;
	wire new_net_20868;
	wire new_net_18362;
	wire new_net_10003;
	wire new_net_6603;
	wire new_net_2927;
	wire _0600_;
	wire _1020_;
	wire _0180_;
	wire new_net_20797;
	wire new_net_21358;
	wire new_net_15786;
	wire new_net_12390;
	wire new_net_12280;
	wire _1204_;
	wire new_net_2566;
	wire new_net_195;
	wire new_net_5660;
	wire new_net_10006;
	wire new_net_18387;
	wire new_net_20929;
	wire new_net_13863;
	wire new_net_18738;
	wire new_net_14749;
	wire new_net_13816;
	wire new_net_7546;
	wire new_net_7441;
	wire new_net_10991;
	wire _0601_;
	wire _1021_;
	wire _0181_;
	wire new_net_19586;
	wire new_net_11655;
	wire new_net_6538;
	wire new_net_14868;
	wire new_net_16894;
	wire _1652_;
	wire new_net_1938;
	wire new_net_3027;
	wire new_net_7246;
	wire new_net_6012;
	wire new_net_10568;
	wire new_net_19844;
	wire new_net_20571;
	wire new_net_262;
	wire new_net_2546;
	wire new_net_11632;
	wire new_net_12221;
	wire new_net_12316;
	wire new_net_17057;
	wire new_net_12174;
	wire new_net_17400;
	wire new_net_14981;
	wire new_net_15320;
	wire new_net_5382;
	wire new_net_7621;
	wire new_net_9246;
	wire new_net_6522;
	wire new_net_6737;
	wire new_net_2966;
	wire new_net_18825;
	wire new_net_260;
	wire new_net_1501;
	wire new_net_1668;
	wire new_net_3738;
	wire new_net_5549;
	wire new_net_6812;
	wire new_net_21431;
	wire new_net_20738;
	wire new_net_18629;
	wire new_net_2542;
	wire new_net_1276;
	wire new_net_1671;
	wire new_net_6820;
	wire new_net_19539;
	wire new_net_19551;
	wire new_net_261;
	wire new_net_1289;
	wire new_net_1652;
	wire new_net_3026;
	wire new_net_7619;
	wire new_net_9172;
	wire new_net_10969;
	wire new_net_10569;
	wire new_net_19721;
	wire new_net_2537;
	wire new_net_3019;
	wire new_net_6014;
	wire new_net_9722;
	wire new_net_19845;
	wire new_net_20572;
	wire new_net_20556;
	wire new_net_258;
	wire new_net_5545;
	wire new_net_11633;
	wire new_net_12175;
	wire new_net_12222;
	wire new_net_17058;
	wire new_net_12317;
	wire new_net_14264;
	wire new_net_14982;
	wire new_net_15321;
	wire new_net_3224;
	wire new_net_7372;
	wire new_net_21078;
	wire new_net_2600;
	wire new_net_263;
	wire new_net_6838;
	wire new_net_8344;
	wire new_net_3740;
	wire new_net_7376;
	wire new_net_21432;
	wire new_net_1048;
	wire new_net_18500;
	wire new_net_1678;
	wire new_net_994;
	wire new_net_1508;
	wire new_net_5546;
	wire new_net_9593;
	wire new_net_7623;
	wire new_net_19540;
	wire new_net_6816;
	wire new_net_3812;
	wire new_net_8346;
	wire new_net_10970;
	wire new_net_3742;
	wire new_net_4257;
	wire new_net_19846;
	wire new_net_20573;
	wire new_net_21079;
	wire new_net_18095;
	wire new_net_18060;
	wire new_net_1672;
	wire new_net_11989;
	wire new_net_11634;
	wire new_net_12223;
	wire new_net_12318;
	wire new_net_17059;
	wire new_net_8349;
	wire new_net_12176;
	wire new_net_17402;
	wire new_net_15322;
	wire new_net_18014;
	wire new_net_6011;
	wire new_net_6818;
	wire new_net_9164;
	wire new_net_20018;
	wire new_net_1503;
	wire new_net_2965;
	wire new_net_3225;
	wire new_net_8362;
	wire new_net_9166;
	wire new_net_17901;
	wire new_net_1504;
	wire new_net_3226;
	wire new_net_5548;
	wire new_net_10566;
	wire new_net_9169;
	wire new_net_10229;
	wire new_net_19627;
	wire new_net_21433;
	wire new_net_18305;
	wire new_net_1277;
	wire new_net_2543;
	wire new_net_1677;
	wire new_net_3020;
	wire new_net_1506;
	wire new_net_9716;
	wire new_net_19541;
	wire new_net_1675;
	wire new_net_3029;
	wire new_net_10971;
	wire new_net_7374;
	wire new_net_265;
	wire new_net_7243;
	wire new_net_8347;
	wire new_net_19847;
	wire new_net_20574;
	wire new_net_21076;
	wire new_net_1509;
	wire new_net_2541;
	wire new_net_11990;
	wire new_net_13030;
	wire new_net_8345;
	wire new_net_12177;
	wire new_net_13265;
	wire new_net_16754;
	wire new_net_12224;
	wire new_net_17060;
	wire new_net_383;
	wire new_net_3018;
	wire new_net_6811;
	wire new_net_9805;
	wire new_net_18875;
	wire new_net_20823;
	wire new_net_17932;
	wire new_net_2964;
	wire new_net_4507;
	wire new_net_5035;
	wire new_net_7375;
	wire new_net_19720;
	wire new_net_18590;
	wire new_net_2972;
	wire new_net_6009;
	wire new_net_21434;
	wire new_net_150;
	wire new_net_1931;
	wire new_net_10572;
	wire new_net_19306;
	wire new_net_19542;
	wire new_net_18101;
	wire new_net_268;
	wire new_net_1930;
	wire new_net_2547;
	wire new_net_9717;
	wire new_net_14983;
	wire new_net_3806;
	wire new_net_4510;
	wire new_net_10972;
	wire new_net_3379;
	wire new_net_7377;
	wire new_net_1935;
	wire new_net_3744;
	wire new_net_5378;
	wire new_net_19848;
	wire new_net_20575;
	wire new_net_21077;
	wire new_net_18080;
	wire new_net_21145;
	wire new_net_11695;
	wire new_net_13266;
	wire new_net_17061;
	wire new_net_5034;
	wire new_net_12320;
	wire new_net_14267;
	wire new_net_11991;
	wire new_net_15324;
	wire new_net_17593;
	wire new_net_11636;
	wire new_net_251;
	wire new_net_1502;
	wire new_net_9721;
	wire new_net_4511;
	wire new_net_5033;
	wire new_net_8367;
	wire new_net_6814;
	wire new_net_21075;
	wire new_net_20869;
	wire new_net_18363;
	wire new_net_20798;
	wire new_net_7241;
	wire new_net_9145;
	wire new_net_19712;
	wire new_net_15787;
	wire new_net_18388;
	wire new_net_264;
	wire new_net_1280;
	wire new_net_6836;
	wire new_net_21435;
	wire new_net_18739;
	wire new_net_995;
	wire new_net_10571;
	wire new_net_3227;
	wire new_net_4512;
	wire new_net_8366;
	wire new_net_9170;
	wire new_net_19543;
	wire new_net_19719;
	wire new_net_20010;
	wire new_net_16895;
	wire new_net_2963;
	wire new_net_3025;
	wire new_net_6005;
	wire new_net_10973;
	wire new_net_7380;
	wire new_net_1288;
	wire new_net_4258;
	wire new_net_6837;
	wire new_net_19849;
	wire new_net_20576;
	wire new_net_1674;
	wire new_net_3809;
	wire new_net_7379;
	wire new_net_9247;
	wire new_net_11696;
	wire new_net_13267;
	wire new_net_9715;
	wire new_net_11992;
	wire new_net_11637;
	wire new_net_12226;
	wire new_net_3017;
	wire new_net_5542;
	wire new_net_19302;
	wire new_net_21074;
	wire new_net_20218;
	wire new_net_18826;
	wire new_net_1654;
	wire new_net_2548;
	wire new_net_1281;
	wire new_net_2973;
	wire new_net_6815;
	wire new_net_20009;
	wire new_net_21436;
	wire new_net_18630;
	wire new_net_2968;
	wire new_net_8369;
	wire new_net_9167;
	wire new_net_19544;
	wire new_net_19718;
	wire new_net_2247;
	wire new_net_2545;
	wire new_net_2969;
	wire new_net_9713;
	wire new_net_8342;
	wire new_net_7624;
	wire new_net_10974;
	wire new_net_20013;
	wire new_net_989;
	wire new_net_7627;
	wire new_net_19711;
	wire new_net_19850;
	wire new_net_20577;
	wire new_net_20600;
	wire new_net_2439;
	wire new_net_267;
	wire new_net_3808;
	wire new_net_11697;
	wire new_net_13268;
	wire new_net_6821;
	wire new_net_11993;
	wire new_net_11638;
	wire new_net_12227;
	wire new_net_12322;
	wire new_net_17063;
	wire new_net_1507;
	wire new_net_9719;
	wire new_net_20017;
	wire new_net_1284;
	wire new_net_2971;
	wire new_net_8340;
	wire new_net_7620;
	wire new_net_12790;
	wire new_net_16240;
	wire _0000_;
	wire new_net_1650;
	wire new_net_21437;
	wire new_net_1279;
	wire new_net_2962;
	wire new_net_3745;
	wire new_net_5782;
	wire new_net_7240;
	wire new_net_19545;
	wire new_net_748;
	wire new_net_10975;
	wire new_net_16757;
	wire new_net_1673;
	wire new_net_1278;
	wire new_net_4506;
	wire new_net_6007;
	wire new_net_19716;
	wire new_net_1933;
	wire new_net_3739;
	wire new_net_5781;
	wire new_net_19851;
	wire new_net_20578;
	wire new_net_18096;
	wire new_net_8364;
	wire _0001_;
	wire new_net_1653;
	wire new_net_3811;
	wire new_net_9248;
	wire new_net_11698;
	wire new_net_13269;
	wire new_net_11994;
	wire new_net_11639;
	wire new_net_12228;
	wire new_net_18061;
	wire new_net_18015;
	wire new_net_992;
	wire new_net_6822;
	wire new_net_5784;
	wire new_net_12713;
	wire new_net_8361;
	wire new_net_1669;
	wire new_net_3022;
	wire new_net_4508;
	wire new_net_5543;
	wire new_net_5783;
	wire new_net_9144;
	wire new_net_9595;
	wire new_net_17902;
	wire new_net_1666;
	wire new_net_21438;
	wire new_net_15249;
	wire new_net_9165;
	wire new_net_3030;
	wire _0002_;
	wire new_net_6004;
	wire new_net_19546;
	wire new_net_20011;
	wire new_net_8370;
	wire new_net_10976;
	wire new_net_993;
	wire new_net_1283;
	wire new_net_3311;
	wire new_net_3023;
	wire new_net_2538;
	wire new_net_3443;
	wire new_net_19303;
	wire new_net_19852;
	wire new_net_20579;
	wire new_net_21071;
	wire new_net_259;
	wire new_net_8360;
	wire new_net_16758;
	wire new_net_11699;
	wire new_net_13270;
	wire new_net_11995;
	wire new_net_11640;
	wire new_net_12229;
	wire new_net_12324;
	wire new_net_17065;
	wire new_net_378;
	wire _0003_;
	wire new_net_996;
	wire new_net_1667;
	wire new_net_2540;
	wire new_net_18876;
	wire new_net_1239;
	wire new_net_255;
	wire new_net_10227;
	wire new_net_2539;
	wire new_net_7622;
	wire new_net_17933;
	wire new_net_18591;
	wire new_net_1932;
	wire new_net_5377;
	wire new_net_19304;
	wire new_net_21439;
	wire new_net_158;
	wire new_net_3021;
	wire new_net_254;
	wire new_net_5384;
	wire new_net_4504;
	wire new_net_19305;
	wire new_net_19547;
	wire _0004_;
	wire new_net_253;
	wire new_net_2970;
	wire new_net_9171;
	wire new_net_18102;
	wire new_net_1929;
	wire new_net_3028;
	wire new_net_7378;
	wire new_net_9594;
	wire new_net_19853;
	wire new_net_20580;
	wire new_net_21072;
	wire new_net_19649;
	wire new_net_20361;
	wire new_net_18081;
	wire new_net_21146;
	wire new_net_13036;
	wire new_net_14272;
	wire new_net_17598;
	wire new_net_2544;
	wire new_net_1275;
	wire new_net_4259;
	wire new_net_9142;
	wire new_net_16759;
	wire new_net_11700;
	wire new_net_13271;
	wire new_net_257;
	wire new_net_8341;
	wire new_net_21070;
	wire new_net_20870;
	wire new_net_18364;
	wire _0005_;
	wire new_net_256;
	wire new_net_1285;
	wire new_net_2967;
	wire new_net_5380;
	wire new_net_6010;
	wire new_net_9720;
	wire new_net_10567;
	wire new_net_988;
	wire new_net_1676;
	wire new_net_3312;
	wire new_net_10977;
	wire new_net_5547;
	wire _1211_;
	wire new_net_18389;
	wire new_net_20016;
	wire new_net_21440;
	wire new_net_18740;
	wire new_net_1651;
	wire new_net_4503;
	wire new_net_5037;
	wire new_net_8348;
	wire new_net_19548;
	wire new_net_6839;
	wire _0006_;
	wire new_net_998;
	wire new_net_8368;
	wire new_net_3024;
	wire new_net_5780;
	wire new_net_19715;
	wire new_net_16896;
	wire new_net_1937;
	wire new_net_3810;
	wire new_net_19854;
	wire new_net_20581;
	wire _1659_;
	wire new_net_3588;
	wire new_net_7626;
	wire new_net_13037;
	wire new_net_14273;
	wire new_net_17599;
	wire new_net_1936;
	wire _0007_;
	wire new_net_1287;
	wire new_net_16760;
	wire new_net_11701;
	wire new_net_13272;
	wire new_net_1649;
	wire new_net_252;
	wire new_net_1286;
	wire new_net_1510;
	wire new_net_10224;
	wire new_net_5541;
	wire new_net_7239;
	wire new_net_6013;
	wire _0008_;
	wire new_net_990;
	wire new_net_1670;
	wire new_net_10228;
	wire new_net_3741;
	wire new_net_10570;
	wire new_net_8343;
	wire new_net_18827;
	wire new_net_1282;
	wire new_net_5381;
	wire new_net_6813;
	wire new_net_21441;
	wire new_net_4256;
	wire _0009_;
	wire new_net_997;
	wire new_net_3310;
	wire new_net_9714;
	wire new_net_5779;
	wire new_net_9143;
	wire new_net_5379;
	wire new_net_15219;
	wire new_net_18631;
	wire new_net_19877;
	wire new_net_10226;
	wire new_net_10978;
	wire new_net_20015;
	wire new_net_21364;
	wire _0010_;
	wire new_net_999;
	wire new_net_1505;
	wire new_net_5038;
	wire new_net_8359;
	wire new_net_19855;
	wire new_net_20582;
	wire new_net_3406;
	wire new_net_13038;
	wire new_net_14274;
	wire new_net_17600;
	wire new_net_266;
	wire new_net_4509;
	wire new_net_8365;
	wire new_net_10225;
	wire new_net_16761;
	wire new_net_11702;
	wire new_net_13273;
	wire _0011_;
	wire new_net_991;
	wire new_net_7373;
	wire new_net_9245;
	wire new_net_7242;
	wire new_net_21069;
	wire new_net_6817;
	wire new_net_3807;
	wire _0012_;
	wire new_net_1934;
	wire new_net_5544;
	wire new_net_3743;
	wire new_net_19713;
	wire new_net_21442;
	wire new_net_14701;
	wire new_net_5383;
	wire new_net_10233;
	wire new_net_19550;
	wire _0013_;
	wire new_net_4505;
	wire new_net_8363;
	wire new_net_10232;
	wire new_net_10979;
	wire new_net_9718;
	wire new_net_15491;
	wire new_net_7244;
	wire new_net_20014;
	wire new_net_2923;
	wire new_net_18097;
	wire new_net_18062;
	wire new_net_3231;
	wire new_net_7501;
	wire new_net_6983;
	wire new_net_18016;
	wire new_net_12714;
	wire new_net_9439;
	wire new_net_14944;
	wire new_net_15438;
	wire new_net_15615;
	wire new_net_955;
	wire new_net_7504;
	wire new_net_16099;
	wire new_net_12624;
	wire new_net_14074;
	wire new_net_16111;
	wire new_net_3010;
	wire new_net_7529;
	wire new_net_7672;
	wire new_net_13518;
	wire new_net_9003;
	wire new_net_19771;
	wire new_net_19878;
	wire new_net_17903;
	wire new_net_7154;
	wire new_net_10449;
	wire new_net_5359;
	wire new_net_15261;
	wire new_net_2007;
	wire new_net_2062;
	wire new_net_4960;
	wire new_net_7666;
	wire new_net_480;
	wire new_net_8277;
	wire new_net_3881;
	wire new_net_9094;
	wire new_net_5607;
	wire new_net_15224;
	wire new_net_20999;
	wire new_net_946;
	wire new_net_3617;
	wire new_net_4966;
	wire new_net_7153;
	wire new_net_10992;
	wire new_net_5357;
	wire new_net_5611;
	wire new_net_16193;
	wire new_net_19150;
	wire new_net_3518;
	wire new_net_7156;
	wire new_net_2055;
	wire new_net_10642;
	wire new_net_8999;
	wire new_net_13590;
	wire new_net_15616;
	wire new_net_3522;
	wire new_net_3616;
	wire new_net_4498;
	wire new_net_4977;
	wire new_net_5355;
	wire new_net_16100;
	wire new_net_12625;
	wire new_net_14075;
	wire new_net_16112;
	wire new_net_18877;
	wire new_net_8691;
	wire new_net_15262;
	wire new_net_15223;
	wire new_net_19772;
	wire new_net_18592;
	wire new_net_21325;
	wire new_net_2675;
	wire new_net_4891;
	wire new_net_5854;
	wire new_net_7668;
	wire new_net_9444;
	wire new_net_9087;
	wire new_net_10633;
	wire new_net_6452;
	wire new_net_4964;
	wire new_net_19127;
	wire new_net_21000;
	wire new_net_18103;
	wire new_net_15439;
	wire new_net_7505;
	wire new_net_8787;
	wire new_net_10451;
	wire new_net_10993;
	wire new_net_3230;
	wire new_net_6873;
	wire new_net_18082;
	wire new_net_21147;
	wire new_net_14943;
	wire new_net_19160;
	wire new_net_15428;
	wire new_net_2058;
	wire new_net_2672;
	wire new_net_15617;
	wire new_net_16101;
	wire new_net_477;
	wire new_net_12626;
	wire new_net_14076;
	wire new_net_13300;
	wire new_net_16552;
	wire new_net_10120;
	wire new_net_18365;
	wire new_net_2053;
	wire new_net_3233;
	wire new_net_8786;
	wire new_net_8689;
	wire new_net_15263;
	wire new_net_16192;
	wire new_net_19137;
	wire new_net_19773;
	wire new_net_15789;
	wire new_net_18390;
	wire new_net_3464;
	wire new_net_483;
	wire new_net_5174;
	wire new_net_5092;
	wire new_net_7395;
	wire new_net_18741;
	wire new_net_2678;
	wire new_net_953;
	wire new_net_6875;
	wire new_net_2060;
	wire new_net_3622;
	wire new_net_5094;
	wire new_net_5856;
	wire new_net_6450;
	wire new_net_6990;
	wire new_net_21001;
	wire new_net_950;
	wire new_net_3715;
	wire new_net_4611;
	wire new_net_5851;
	wire new_net_10994;
	wire new_net_16113;
	wire new_net_6993;
	wire new_net_15222;
	wire new_net_14942;
	wire new_net_10637;
	wire new_net_7399;
	wire new_net_9004;
	wire new_net_15429;
	wire new_net_943;
	wire new_net_15440;
	wire new_net_15618;
	wire new_net_16102;
	wire new_net_12627;
	wire new_net_14077;
	wire new_net_13301;
	wire new_net_16553;
	wire new_net_14417;
	wire new_net_3467;
	wire new_net_2061;
	wire new_net_4978;
	wire new_net_3234;
	wire new_net_6872;
	wire new_net_6982;
	wire new_net_16191;
	wire new_net_19774;
	wire new_net_19876;
	wire new_net_18828;
	wire new_net_2681;
	wire new_net_478;
	wire new_net_4607;
	wire new_net_5849;
	wire new_net_9442;
	wire new_net_7507;
	wire new_net_9086;
	wire new_net_6989;
	wire new_net_8696;
	wire new_net_19136;
	wire new_net_4501;
	wire new_net_7509;
	wire new_net_9090;
	wire new_net_6933;
	wire new_net_6449;
	wire new_net_6994;
	wire new_net_6986;
	wire new_net_19474;
	wire new_net_3519;
	wire new_net_3619;
	wire new_net_3883;
	wire new_net_8686;
	wire new_net_19880;
	wire new_net_21002;
	wire new_net_4605;
	wire new_net_10995;
	wire new_net_5356;
	wire new_net_15264;
	wire new_net_15221;
	wire new_net_3009;
	wire new_net_951;
	wire new_net_3462;
	wire new_net_14941;
	wire new_net_7151;
	wire new_net_8005;
	wire new_net_7671;
	wire new_net_19159;
	wire new_net_12296;
	wire new_net_15430;
	wire new_net_15441;
	wire new_net_15619;
	wire new_net_16103;
	wire new_net_12628;
	wire new_net_14078;
	wire new_net_16114;
	wire new_net_16554;
	wire new_net_12770;
	wire new_net_2612;
	wire new_net_16190;
	wire new_net_3013;
	wire new_net_4499;
	wire new_net_5503;
	wire new_net_19775;
	wire new_net_15688;
	wire new_net_3712;
	wire new_net_7528;
	wire new_net_8998;
	wire new_net_8788;
	wire new_net_3880;
	wire new_net_6870;
	wire new_net_6985;
	wire new_net_3884;
	wire new_net_4889;
	wire new_net_6453;
	wire new_net_19135;
	wire new_net_2676;
	wire new_net_485;
	wire new_net_949;
	wire new_net_4497;
	wire new_net_8783;
	wire new_net_3236;
	wire new_net_8687;
	wire new_net_19152;
	wire new_net_21003;
	wire new_net_3465;
	wire new_net_7603;
	wire new_net_10996;
	wire new_net_6934;
	wire new_net_13302;
	wire new_net_13081;
	wire new_net_10640;
	wire new_net_18098;
	wire new_net_14940;
	wire new_net_5088;
	wire new_net_4575;
	wire new_net_12297;
	wire new_net_15220;
	wire new_net_2680;
	wire new_net_15431;
	wire new_net_15442;
	wire new_net_15620;
	wire new_net_16104;
	wire new_net_12629;
	wire new_net_14079;
	wire new_net_16115;
	wire new_net_16189;
	wire new_net_3516;
	wire new_net_3882;
	wire new_net_7148;
	wire new_net_3387;
	wire new_net_6988;
	wire new_net_14438;
	wire new_net_7667;
	wire new_net_19776;
	wire new_net_19881;
	wire new_net_17904;
	wire new_net_4577;
	wire new_net_4892;
	wire new_net_10638;
	wire new_net_8690;
	wire new_net_17355;
	wire new_net_3011;
	wire new_net_7502;
	wire new_net_5848;
	wire new_net_10634;
	wire new_net_4962;
	wire new_net_401;
	wire new_net_19221;
	wire new_net_20714;
	wire new_net_20299;
	wire new_net_6987;
	wire new_net_2682;
	wire new_net_2054;
	wire new_net_4500;
	wire new_net_5850;
	wire new_net_7503;
	wire new_net_8785;
	wire new_net_19134;
	wire new_net_21004;
	wire new_net_19982;
	wire new_net_5847;
	wire new_net_6877;
	wire new_net_10997;
	wire new_net_3435;
	wire _1512_;
	wire new_net_3885;
	wire new_net_4888;
	wire new_net_5846;
	wire new_net_14939;
	wire new_net_7606;
	wire new_net_8688;
	wire new_net_7394;
	wire new_net_19158;
	wire new_net_19882;
	wire _0350_;
	wire new_net_17981;
	wire new_net_12630;
	wire new_net_12298;
	wire new_net_16556;
	wire new_net_15432;
	wire new_net_3524;
	wire new_net_9005;
	wire new_net_13456;
	wire new_net_15443;
	wire new_net_14080;
	wire new_net_12772;
	wire new_net_6431;
	wire new_net_14408;
	wire new_net_16188;
	wire new_net_2059;
	wire new_net_3469;
	wire new_net_3623;
	wire new_net_5086;
	wire new_net_7147;
	wire new_net_10450;
	wire new_net_6997;
	wire new_net_7398;
	wire new_net_15267;
	wire new_net_18593;
	wire new_net_7402;
	wire new_net_2057;
	wire new_net_7526;
	wire new_net_3887;
	wire new_net_14825;
	wire new_net_15651;
	wire new_net_9091;
	wire _1358_;
	wire new_net_3228;
	wire new_net_12980;
	wire new_net_3468;
	wire new_net_4612;
	wire new_net_9000;
	wire new_net_9092;
	wire new_net_6454;
	wire new_net_19153;
	wire new_net_8695;
	wire new_net_4496;
	wire new_net_4608;
	wire new_net_5090;
	wire new_net_8792;
	wire new_net_9089;
	wire new_net_6995;
	wire new_net_21005;
	wire new_net_18104;
	wire new_net_7674;
	wire new_net_6979;
	wire new_net_4574;
	wire new_net_5852;
	wire new_net_6446;
	wire new_net_10453;
	wire new_net_10998;
	wire new_net_19133;
	wire new_net_18083;
	wire new_net_21148;
	wire new_net_942;
	wire new_net_3463;
	wire new_net_3520;
	wire new_net_9438;
	wire new_net_14938;
	wire new_net_4887;
	wire new_net_19883;
	wire new_net_12335;
	wire new_net_15270;
	wire new_net_12299;
	wire new_net_15218;
	wire new_net_2063;
	wire new_net_3466;
	wire new_net_4981;
	wire new_net_15433;
	wire new_net_15444;
	wire new_net_15622;
	wire new_net_1829;
	wire new_net_7396;
	wire new_net_6980;
	wire new_net_3620;
	wire new_net_5362;
	wire new_net_16187;
	wire new_net_15268;
	wire new_net_18366;
	wire new_net_19778;
	wire new_net_19884;
	wire new_net_3240;
	wire new_net_4609;
	wire new_net_4965;
	wire _1218_;
	wire new_net_18391;
	wire new_net_18742;
	wire new_net_7393;
	wire new_net_4606;
	wire new_net_9446;
	wire new_net_3014;
	wire new_net_947;
	wire new_net_3618;
	wire new_net_9441;
	wire new_net_8278;
	wire new_net_9085;
	wire new_net_21006;
	wire new_net_484;
	wire new_net_3879;
	wire new_net_5610;
	wire new_net_10999;
	wire new_net_2673;
	wire new_net_954;
	wire new_net_14937;
	wire new_net_7500;
	wire new_net_8784;
	wire new_net_19132;
	wire new_net_19157;
	wire new_net_8570;
	wire new_net_5606;
	wire new_net_12336;
	wire new_net_17041;
	wire new_net_4573;
	wire new_net_12300;
	wire new_net_15217;
	wire new_net_15445;
	wire new_net_15623;
	wire new_net_15434;
	wire new_net_7506;
	wire new_net_3238;
	wire new_net_3621;
	wire new_net_16186;
	wire new_net_10447;
	wire new_net_13593;
	wire new_net_19779;
	wire new_net_18829;
	wire new_net_7397;
	wire new_net_9006;
	wire new_net_6456;
	wire new_net_5612;
	wire new_net_487;
	wire new_net_5172;
	wire new_net_9093;
	wire new_net_6445;
	wire new_net_7670;
	wire new_net_948;
	wire new_net_3239;
	wire new_net_3461;
	wire new_net_8002;
	wire new_net_4576;
	wire new_net_10635;
	wire new_net_19154;
	wire new_net_21007;
	wire new_net_9436;
	wire new_net_11000;
	wire new_net_3012;
	wire new_net_476;
	wire new_net_6868;
	wire new_net_5358;
	wire new_net_8004;
	wire new_net_15269;
	wire new_net_8791;
	wire new_net_2674;
	wire new_net_7527;
	wire new_net_14936;
	wire new_net_19610;
	wire new_net_12775;
	wire new_net_13459;
	wire new_net_12337;
	wire new_net_17042;
	wire new_net_7149;
	wire new_net_14083;
	wire new_net_12301;
	wire new_net_16119;
	wire new_net_15446;
	wire new_net_15624;
	wire new_net_4572;
	wire new_net_482;
	wire new_net_16185;
	wire new_net_4493;
	wire new_net_7499;
	wire new_net_3229;
	wire new_net_19780;
	wire new_net_7150;
	wire new_net_8794;
	wire new_net_9447;
	wire new_net_18655;
	wire new_net_19185;
	wire new_net_6455;
	wire new_net_6992;
	wire new_net_10636;
	wire new_net_3716;
	wire new_net_14703;
	wire new_net_4502;
	wire new_net_5609;
	wire new_net_7401;
	wire new_net_2677;
	wire new_net_3237;
	wire new_net_4963;
	wire new_net_5091;
	wire new_net_7155;
	wire new_net_5360;
	wire new_net_19128;
	wire new_net_21008;
	wire new_net_7669;
	wire new_net_4571;
	wire new_net_9002;
	wire new_net_5173;
	wire new_net_5093;
	wire new_net_9088;
	wire new_net_11001;
	wire new_net_425;
	wire new_net_18099;
	wire new_net_7403;
	wire new_net_15271;
	wire new_net_479;
	wire new_net_5089;
	wire new_net_5502;
	wire new_net_14935;
	wire new_net_7508;
	wire new_net_19156;
	wire new_net_6998;
	wire new_net_10639;
	wire new_net_12776;
	wire new_net_13460;
	wire new_net_8694;
	wire new_net_12338;
	wire new_net_17043;
	wire new_net_12302;
	wire new_net_15215;
	wire new_net_15436;
	wire new_net_7400;
	wire new_net_3517;
	wire new_net_16184;
	wire new_net_9001;
	wire new_net_9443;
	wire new_net_14933;
	wire new_net_4495;
	wire new_net_10452;
	wire new_net_19130;
	wire new_net_19781;
	wire new_net_17905;
	wire new_net_6448;
	wire new_net_481;
	wire new_net_952;
	wire new_net_4893;
	wire new_net_4959;
	wire new_net_486;
	wire new_net_3713;
	wire new_net_3886;
	wire new_net_4610;
	wire new_net_8692;
	wire new_net_16182;
	wire new_net_3523;
	wire new_net_9440;
	wire new_net_4494;
	wire new_net_21009;
	wire new_net_17140;
	wire new_net_3016;
	wire new_net_944;
	wire new_net_5853;
	wire new_net_7152;
	wire new_net_11002;
	wire new_net_6451;
	wire new_net_4961;
	wire new_net_941;
	wire new_net_3015;
	wire new_net_14934;
	wire new_net_8279;
	wire new_net_10454;
	wire new_net_17979;
	wire new_net_17982;
	wire new_net_12777;
	wire new_net_13461;
	wire new_net_945;
	wire new_net_3714;
	wire new_net_12339;
	wire new_net_17044;
	wire new_net_12303;
	wire new_net_15214;
	wire new_net_15437;
	wire new_net_5171;
	wire new_net_16183;
	wire new_net_9437;
	wire new_net_19782;
	wire new_net_19875;
	wire new_net_18594;
	wire new_net_5855;
	wire new_net_6874;
	wire new_net_3521;
	wire new_net_3888;
	wire new_net_4890;
	wire new_net_5361;
	wire new_net_5501;
	wire new_net_6981;
	wire new_net_9445;
	wire new_net_10448;
	wire new_net_19777;
	wire new_net_21327;
	wire new_net_12887;
	wire new_net_3235;
	wire new_net_6984;
	wire new_net_2056;
	wire new_net_2679;
	wire new_net_5504;
	wire new_net_15213;
	wire new_net_15104;
	wire new_net_10456;
	wire new_net_21010;
	wire new_net_18105;
	wire new_net_3530;
	wire new_net_6447;
	wire new_net_6869;
	wire new_net_10643;
	wire new_net_8790;
	wire new_net_11003;
	wire new_net_19267;
	wire new_net_19886;
	wire new_net_6380;
	wire new_net_18084;
	wire new_net_21149;
	wire new_net_18887;
	wire new_net_21296;
	wire new_net_2952;
	wire new_net_7420;
	wire new_net_4420;
	wire new_net_20547;
	wire new_net_18367;
	wire new_net_12553;
	wire new_net_12731;
	wire new_net_15048;
	wire new_net_11894;
	wire new_net_17351;
	wire _0392_;
	wire new_net_3039;
	wire new_net_2951;
	wire new_net_10262;
	wire new_net_16514;
	wire new_net_21362;
	wire new_net_12225;
	wire new_net_5940;
	wire new_net_3897;
	wire new_net_4383;
	wire new_net_4905;
	wire new_net_6137;
	wire new_net_10208;
	wire new_net_18392;
	wire new_net_18443;
	wire new_net_18743;
	wire new_net_10478;
	wire _0393_;
	wire new_net_3040;
	wire new_net_3724;
	wire new_net_5443;
	wire new_net_7937;
	wire new_net_21337;
	wire new_net_10471;
	wire new_net_9201;
	wire new_net_8261;
	wire new_net_11892;
	wire new_net_20210;
	wire new_net_16899;
	wire new_net_10475;
	wire _0394_;
	wire new_net_5776;
	wire new_net_20088;
	wire new_net_17495;
	wire new_net_10666;
	wire new_net_11588;
	wire new_net_11436;
	wire new_net_17246;
	wire new_net_11240;
	wire new_net_11460;
	wire new_net_11893;
	wire new_net_19623;
	wire new_net_20871;
	wire new_net_496;
	wire _0395_;
	wire new_net_2297;
	wire new_net_17352;
	wire new_net_8843;
	wire new_net_4819;
	wire new_net_3042;
	wire new_net_20548;
	wire new_net_13592;
	wire new_net_12022;
	wire new_net_14639;
	wire new_net_12732;
	wire new_net_13652;
	wire new_net_14439;
	wire new_net_16515;
	wire new_net_1152;
	wire new_net_4427;
	wire new_net_12910;
	wire new_net_13724;
	wire new_net_18830;
	wire new_net_10472;
	wire _0396_;
	wire new_net_3728;
	wire new_net_10261;
	wire new_net_17350;
	wire new_net_17245;
	wire new_net_4424;
	wire new_net_19874;
	wire new_net_20211;
	wire new_net_10060;
	wire new_net_6128;
	wire new_net_21338;
	wire new_net_15216;
	wire new_net_16643;
	wire _0397_;
	wire new_net_3223;
	wire new_net_4080;
	wire new_net_4378;
	wire new_net_8903;
	wire new_net_9210;
	wire new_net_18452;
	wire new_net_10203;
	wire new_net_3213;
	wire new_net_3725;
	wire new_net_7422;
	wire new_net_19873;
	wire new_net_20089;
	wire new_net_10061;
	wire new_net_497;
	wire _0398_;
	wire new_net_2960;
	wire new_net_11589;
	wire new_net_7089;
	wire new_net_11437;
	wire new_net_14157;
	wire new_net_11241;
	wire new_net_11461;
	wire new_net_19212;
	wire new_net_16633;
	wire new_net_498;
	wire new_net_2953;
	wire new_net_3036;
	wire new_net_1256;
	wire new_net_5391;
	wire new_net_20549;
	wire new_net_17569;
	wire new_net_3647;
	wire new_net_10210;
	wire new_net_12023;
	wire new_net_16871;
	wire _0399_;
	wire new_net_3218;
	wire new_net_12733;
	wire new_net_13653;
	wire new_net_14440;
	wire new_net_17886;
	wire new_net_3222;
	wire new_net_7936;
	wire new_net_17349;
	wire new_net_17244;
	wire new_net_18656;
	wire new_net_19186;
	wire new_net_14704;
	wire new_net_16642;
	wire new_net_12671;
	wire _0400_;
	wire new_net_3309;
	wire new_net_4382;
	wire new_net_5440;
	wire new_net_17243;
	wire new_net_18451;
	wire new_net_19872;
	wire new_net_21339;
	wire new_net_5945;
	wire new_net_492;
	wire new_net_2302;
	wire new_net_5447;
	wire new_net_15494;
	wire new_net_21405;
	wire new_net_10204;
	wire _0401_;
	wire new_net_1248;
	wire new_net_2299;
	wire new_net_4381;
	wire new_net_20090;
	wire new_net_14640;
	wire new_net_3038;
	wire new_net_4821;
	wire new_net_5385;
	wire new_net_11590;
	wire new_net_9207;
	wire new_net_11438;
	wire new_net_11242;
	wire new_net_11462;
	wire new_net_6138;
	wire new_net_10063;
	wire _0402_;
	wire new_net_1262;
	wire new_net_5446;
	wire new_net_8260;
	wire new_net_16574;
	wire new_net_18444;
	wire new_net_20550;
	wire new_net_3363;
	wire new_net_12024;
	wire new_net_1150;
	wire new_net_1250;
	wire new_net_3219;
	wire new_net_12734;
	wire new_net_13654;
	wire new_net_14441;
	wire new_net_16517;
	wire new_net_12912;
	wire new_net_16516;
	wire new_net_17906;
	wire new_net_17589;
	wire new_net_4419;
	wire new_net_10209;
	wire _0403_;
	wire new_net_17348;
	wire new_net_6131;
	wire new_net_17357;
	wire new_net_19119;
	wire new_net_12672;
	wire new_net_4073;
	wire new_net_4081;
	wire new_net_4822;
	wire new_net_5141;
	wire new_net_5387;
	wire new_net_20213;
	wire new_net_21340;
	wire new_net_18888;
	wire new_net_10057;
	wire _0404_;
	wire new_net_10720;
	wire new_net_10058;
	wire new_net_3033;
	wire new_net_3217;
	wire new_net_3650;
	wire new_net_5144;
	wire new_net_10715;
	wire new_net_7934;
	wire new_net_20091;
	wire new_net_1528;
	wire new_net_18050;
	wire new_net_16640;
	wire _0405_;
	wire new_net_3453;
	wire new_net_5148;
	wire new_net_11591;
	wire new_net_10716;
	wire new_net_11439;
	wire new_net_11243;
	wire new_net_4521;
	wire new_net_11463;
	wire new_net_17983;
	wire new_net_6134;
	wire new_net_3898;
	wire new_net_4069;
	wire new_net_8844;
	wire new_net_9203;
	wire new_net_20551;
	wire new_net_21396;
	wire new_net_12557;
	wire new_net_16873;
	wire new_net_17571;
	wire new_net_5774;
	wire new_net_12025;
	wire new_net_14641;
	wire _0406_;
	wire new_net_1257;
	wire new_net_2955;
	wire new_net_3649;
	wire new_net_18595;
	wire new_net_10066;
	wire new_net_493;
	wire new_net_1155;
	wire new_net_3318;
	wire new_net_17347;
	wire new_net_5143;
	wire new_net_21397;
	wire _1365_;
	wire new_net_12673;
	wire _0407_;
	wire new_net_1261;
	wire new_net_1157;
	wire new_net_8846;
	wire new_net_8262;
	wire new_net_21341;
	wire new_net_6135;
	wire new_net_16641;
	wire new_net_5772;
	wire new_net_10067;
	wire new_net_4815;
	wire new_net_5444;
	wire new_net_8842;
	wire new_net_9204;
	wire new_net_19227;
	wire new_net_18106;
	wire _0408_;
	wire new_net_4818;
	wire new_net_20092;
	wire new_net_19650;
	wire new_net_2957;
	wire new_net_5150;
	wire new_net_5390;
	wire new_net_6136;
	wire new_net_10259;
	wire new_net_11592;
	wire new_net_11440;
	wire new_net_11244;
	wire new_net_11464;
	wire new_net_17583;
	wire new_net_18085;
	wire new_net_21150;
	wire new_net_18886;
	wire _0409_;
	wire new_net_20552;
	wire new_net_21223;
	wire new_net_12558;
	wire new_net_16874;
	wire new_net_17572;
	wire new_net_12026;
	wire new_net_14642;
	wire new_net_12736;
	wire new_net_13656;
	wire new_net_14443;
	wire new_net_16519;
	wire new_net_12914;
	wire new_net_18368;
	wire _0410_;
	wire new_net_1247;
	wire new_net_5942;
	wire new_net_17346;
	wire new_net_7978;
	wire new_net_17242;
	wire new_net_18445;
	wire new_net_17062;
	wire _1225_;
	wire new_net_18393;
	wire new_net_18744;
	wire new_net_19268;
	wire new_net_2295;
	wire new_net_4817;
	wire new_net_12674;
	wire new_net_8258;
	wire new_net_19257;
	wire new_net_19871;
	wire new_net_21342;
	wire _0411_;
	wire new_net_489;
	wire new_net_3644;
	wire new_net_9964;
	wire new_net_7090;
	wire new_net_19258;
	wire new_net_3082;
	wire new_net_1249;
	wire new_net_2304;
	wire new_net_4071;
	wire new_net_5771;
	wire new_net_5389;
	wire new_net_20093;
	wire new_net_20216;
	wire new_net_21403;
	wire _1673_;
	wire _0412_;
	wire new_net_488;
	wire new_net_2961;
	wire new_net_3646;
	wire new_net_10476;
	wire new_net_10264;
	wire new_net_11593;
	wire new_net_9208;
	wire new_net_11441;
	wire new_net_7935;
	wire new_net_16632;
	wire new_net_1259;
	wire new_net_4077;
	wire new_net_10265;
	wire new_net_10718;
	wire new_net_20553;
	wire new_net_12559;
	wire new_net_16875;
	wire new_net_17573;
	wire _0413_;
	wire new_net_1251;
	wire new_net_3643;
	wire new_net_12027;
	wire new_net_14643;
	wire new_net_12737;
	wire new_net_13657;
	wire new_net_1160;
	wire new_net_3903;
	wire new_net_17345;
	wire new_net_17241;
	wire new_net_3317;
	wire new_net_494;
	wire _0414_;
	wire new_net_4377;
	wire new_net_12675;
	wire new_net_20214;
	wire new_net_21343;
	wire new_net_1252;
	wire new_net_4070;
	wire new_net_4076;
	wire new_net_8839;
	wire new_net_3034;
	wire _0415_;
	wire new_net_2296;
	wire new_net_7087;
	wire new_net_19870;
	wire new_net_20094;
	wire new_net_20217;
	wire new_net_11246;
	wire new_net_11466;
	wire new_net_11898;
	wire new_net_10207;
	wire new_net_3640;
	wire new_net_5142;
	wire new_net_5941;
	wire new_net_11594;
	wire new_net_9209;
	wire new_net_7982;
	wire new_net_6132;
	wire _0416_;
	wire new_net_5770;
	wire new_net_5939;
	wire new_net_7981;
	wire new_net_20554;
	wire new_net_7930;
	wire new_net_16886;
	wire new_net_17585;
	wire new_net_6130;
	wire new_net_12560;
	wire new_net_16876;
	wire new_net_17574;
	wire new_net_3652;
	wire new_net_1154;
	wire new_net_2956;
	wire new_net_19885;
	wire new_net_17887;
	wire _0417_;
	wire new_net_5392;
	wire new_net_7088;
	wire new_net_17344;
	wire new_net_17240;
	wire new_net_18657;
	wire new_net_19187;
	wire new_net_18051;
	wire new_net_10056;
	wire new_net_12676;
	wire new_net_10263;
	wire new_net_19868;
	wire new_net_21344;
	wire new_net_21401;
	wire new_net_4421;
	wire _0418_;
	wire new_net_9961;
	wire new_net_4816;
	wire new_net_21382;
	wire new_net_16639;
	wire new_net_5777;
	wire new_net_18449;
	wire new_net_19869;
	wire new_net_20095;
	wire new_net_2910;
	wire new_net_7931;
	wire new_net_11247;
	wire new_net_11467;
	wire new_net_5436;
	wire _0419_;
	wire new_net_3221;
	wire new_net_11595;
	wire new_net_8845;
	wire new_net_10721;
	wire new_net_7980;
	wire new_net_14509;
	wire new_net_3729;
	wire new_net_5149;
	wire new_net_18442;
	wire new_net_20555;
	wire new_net_12095;
	wire new_net_16887;
	wire new_net_17586;
	wire new_net_12561;
	wire new_net_17575;
	wire _0420_;
	wire new_net_5435;
	wire new_net_16638;
	wire new_net_5778;
	wire new_net_5936;
	wire new_net_12029;
	wire new_net_2959;
	wire new_net_1258;
	wire new_net_5445;
	wire new_net_6129;
	wire new_net_16634;
	wire new_net_12218;
	wire new_net_17343;
	wire new_net_17239;
	wire new_net_17907;
	wire new_net_18989;
	wire new_net_15254;
	wire new_net_17358;
	wire _0421_;
	wire new_net_3035;
	wire new_net_12677;
	wire new_net_8901;
	wire new_net_21345;
	wire new_net_3305;
	wire new_net_4428;
	wire new_net_4820;
	wire new_net_6400;
	wire _0422_;
	wire new_net_10202;
	wire new_net_10719;
	wire new_net_20096;
	wire new_net_11444;
	wire new_net_11248;
	wire new_net_11468;
	wire new_net_5773;
	wire new_net_3900;
	wire new_net_11596;
	wire new_net_10717;
	wire new_net_19226;
	wire new_net_20879;
	wire new_net_21399;
	wire new_net_17984;
	wire new_net_11899;
	wire new_net_2298;
	wire _0423_;
	wire new_net_1153;
	wire new_net_3032;
	wire new_net_3726;
	wire new_net_4423;
	wire new_net_5441;
	wire new_net_5161;
	wire new_net_19259;
	wire new_net_15057;
	wire new_net_15365;
	wire new_net_17681;
	wire new_net_16888;
	wire new_net_17587;
	wire new_net_12562;
	wire new_net_17576;
	wire new_net_495;
	wire new_net_3306;
	wire new_net_5162;
	wire new_net_17238;
	wire new_net_8263;
	wire _0424_;
	wire new_net_1156;
	wire new_net_3648;
	wire new_net_3901;
	wire new_net_4074;
	wire new_net_5448;
	wire new_net_17342;
	wire new_net_21329;
	wire new_net_14828;
	wire new_net_15654;
	wire new_net_12889;
	wire new_net_7929;
	wire new_net_6133;
	wire new_net_3220;
	wire new_net_16637;
	wire new_net_12678;
	wire new_net_10474;
	wire new_net_18447;
	wire new_net_19261;
	wire new_net_21346;
	wire new_net_7938;
	wire _0425_;
	wire new_net_3727;
	wire new_net_3899;
	wire new_net_4426;
	wire new_net_4376;
	wire new_net_10260;
	wire new_net_21400;
	wire new_net_18107;
	wire new_net_491;
	wire new_net_20097;
	wire new_net_3529;
	wire new_net_11445;
	wire new_net_11249;
	wire new_net_11469;
	wire new_net_11900;
	wire new_net_16877;
	wire _0426_;
	wire new_net_3639;
	wire new_net_5775;
	wire new_net_11597;
	wire new_net_4078;
	wire new_net_19651;
	wire new_net_18086;
	wire new_net_21151;
	wire new_net_11901;
	wire new_net_3037;
	wire new_net_4422;
	wire new_net_5147;
	wire new_net_19867;
	wire new_net_20557;
	wire new_net_18885;
	wire new_net_1741;
	wire new_net_15058;
	wire new_net_15366;
	wire new_net_17682;
	wire new_net_16889;
	wire new_net_17588;
	wire new_net_13661;
	wire new_net_12563;
	wire new_net_17577;
	wire _0427_;
	wire new_net_3031;
	wire new_net_18369;
	wire new_net_2301;
	wire new_net_5146;
	wire new_net_5937;
	wire new_net_10469;
	wire new_net_17237;
	wire new_net_10258;
	wire new_net_18394;
	wire new_net_18745;
	wire new_net_12679;
	wire new_net_3041;
	wire _0428_;
	wire new_net_10714;
	wire new_net_3651;
	wire new_net_3642;
	wire new_net_17236;
	wire new_net_1260;
	wire new_net_5442;
	wire new_net_5388;
	wire new_net_3723;
	wire new_net_5164;
	wire _0429_;
	wire new_net_9962;
	wire new_net_1151;
	wire new_net_4079;
	wire new_net_20098;
	wire new_net_20208;
	wire new_net_7086;
	wire new_net_11446;
	wire new_net_8259;
	wire new_net_11250;
	wire new_net_11470;
	wire new_net_6127;
	wire new_net_2958;
	wire new_net_4425;
	wire new_net_10064;
	wire new_net_11598;
	wire new_net_2954;
	wire _0430_;
	wire new_net_2300;
	wire new_net_490;
	wire new_net_4072;
	wire new_net_1159;
	wire new_net_4082;
	wire new_net_20558;
	wire new_net_21395;
	wire new_net_864;
	wire new_net_15059;
	wire new_net_15367;
	wire new_net_17683;
	wire new_net_16525;
	wire new_net_16890;
	wire new_net_17578;
	wire new_net_5944;
	wire new_net_11902;
	wire new_net_12564;
	wire new_net_16878;
	wire new_net_7933;
	wire _0431_;
	wire new_net_1254;
	wire new_net_3645;
	wire new_net_16635;
	wire new_net_10059;
	wire new_net_17341;
	wire new_net_19224;
	wire new_net_19346;
	wire new_net_5386;
	wire new_net_1253;
	wire new_net_12680;
	wire new_net_10473;
	wire new_net_20219;
	wire new_net_21348;
	wire new_net_12353;
	wire new_net_17698;
	wire new_net_8840;
	wire new_net_9206;
	wire _0432_;
	wire new_net_3215;
	wire new_net_3641;
	wire new_net_3902;
	wire new_net_16636;
	wire new_net_10062;
	wire new_net_18446;
	wire new_net_7979;
	wire new_net_7932;
	wire new_net_5163;
	wire new_net_19225;
	wire new_net_20099;
	wire new_net_4083;
	wire new_net_11447;
	wire new_net_11251;
	wire new_net_11599;
	wire _0433_;
	wire new_net_3904;
	wire new_net_11471;
	wire new_net_10266;
	wire new_net_10206;
	wire new_net_12920;
	wire new_net_17779;
	wire new_net_18889;
	wire new_net_6126;
	wire new_net_8239;
	wire new_net_3104;
	wire new_net_4658;
	wire new_net_5003;
	wire new_net_14781;
	wire new_net_20774;
	wire new_net_21385;
	wire new_net_1309;
	wire new_net_12796;
	wire new_net_15692;
	wire new_net_17888;
	wire new_net_5512;
	wire new_net_17282;
	wire new_net_15130;
	wire new_net_15947;
	wire new_net_14251;
	wire new_net_17519;
	wire _0518_;
	wire new_net_1087;
	wire _0182_;
	wire new_net_631;
	wire new_net_18658;
	wire new_net_19188;
	wire new_net_12178;
	wire new_net_5734;
	wire new_net_4295;
	wire new_net_4800;
	wire new_net_20773;
	wire new_net_14883;
	wire new_net_17635;
	wire new_net_3525;
	wire new_net_6015;
	wire _0183_;
	wire _0519_;
	wire new_net_8413;
	wire new_net_14780;
	wire new_net_19628;
	wire new_net_20764;
	wire new_net_6023;
	wire new_net_1393;
	wire new_net_8534;
	wire new_net_10034;
	wire new_net_4663;
	wire new_net_7266;
	wire _0184_;
	wire _0520_;
	wire new_net_3509;
	wire new_net_5000;
	wire new_net_18229;
	wire new_net_14510;
	wire new_net_16205;
	wire new_net_6120;
	wire new_net_11285;
	wire new_net_17269;
	wire new_net_3510;
	wire new_net_4662;
	wire new_net_10839;
	wire new_net_10036;
	wire new_net_11064;
	wire new_net_20799;
	wire new_net_2878;
	wire new_net_13694;
	wire new_net_2446;
	wire new_net_5728;
	wire new_net_9866;
	wire new_net_6760;
	wire new_net_8972;
	wire _0521_;
	wire _0185_;
	wire new_net_3107;
	wire new_net_3508;
	wire new_net_3850;
	wire new_net_14442;
	wire new_net_16518;
	wire new_net_11996;
	wire new_net_17908;
	wire new_net_15948;
	wire new_net_17283;
	wire new_net_7944;
	wire new_net_17520;
	wire new_net_14252;
	wire new_net_1396;
	wire new_net_1091;
	wire new_net_12530;
	wire new_net_15131;
	wire new_net_15995;
	wire new_net_15255;
	wire new_net_17359;
	wire new_net_5509;
	wire new_net_3747;
	wire _0522_;
	wire _0186_;
	wire new_net_17268;
	wire new_net_4772;
	wire new_net_408;
	wire new_net_20300;
	wire new_net_3515;
	wire new_net_4296;
	wire new_net_4799;
	wire new_net_7960;
	wire new_net_16312;
	wire new_net_15435;
	wire new_net_19629;
	wire _0523_;
	wire _0187_;
	wire new_net_8538;
	wire new_net_4249;
	wire new_net_9629;
	wire new_net_19184;
	wire new_net_19621;
	wire new_net_642;
	wire new_net_4824;
	wire new_net_5727;
	wire new_net_6121;
	wire new_net_17985;
	wire new_net_14782;
	wire new_net_5732;
	wire new_net_11286;
	wire new_net_638;
	wire _0188_;
	wire _0524_;
	wire new_net_10840;
	wire new_net_4828;
	wire new_net_11065;
	wire new_net_16304;
	wire new_net_2697;
	wire new_net_1851;
	wire new_net_4305;
	wire new_net_8612;
	wire new_net_17284;
	wire new_net_15132;
	wire new_net_15949;
	wire _0189_;
	wire _0525_;
	wire new_net_14253;
	wire new_net_17521;
	wire new_net_12531;
	wire new_net_14111;
	wire new_net_4255;
	wire new_net_12984;
	wire new_net_14829;
	wire new_net_15655;
	wire _1372_;
	wire new_net_300;
	wire new_net_18679;
	wire new_net_12890;
	wire new_net_16204;
	wire new_net_17267;
	wire new_net_636;
	wire new_net_3750;
	wire new_net_4770;
	wire new_net_7269;
	wire new_net_19173;
	wire new_net_1856;
	wire _0190_;
	wire _0526_;
	wire new_net_7736;
	wire new_net_10028;
	wire new_net_8416;
	wire new_net_19630;
	wire new_net_18108;
	wire new_net_8532;
	wire new_net_19620;
	wire new_net_21393;
	wire new_net_6019;
	wire new_net_5730;
	wire new_net_639;
	wire _0527_;
	wire _0191_;
	wire new_net_1088;
	wire new_net_18227;
	wire new_net_19183;
	wire new_net_18087;
	wire new_net_19652;
	wire new_net_21152;
	wire new_net_10841;
	wire new_net_641;
	wire new_net_4778;
	wire new_net_6123;
	wire new_net_11287;
	wire new_net_14583;
	wire new_net_11066;
	wire new_net_14783;
	wire new_net_18884;
	wire new_net_20801;
	wire new_net_1833;
	wire new_net_9636;
	wire new_net_8238;
	wire new_net_9875;
	wire _0528_;
	wire _0192_;
	wire new_net_6758;
	wire new_net_19619;
	wire new_net_21186;
	wire new_net_18370;
	wire new_net_1754;
	wire new_net_15133;
	wire new_net_15997;
	wire new_net_17285;
	wire new_net_9868;
	wire new_net_14112;
	wire new_net_1852;
	wire new_net_3105;
	wire new_net_4253;
	wire new_net_14254;
	wire new_net_13182;
	wire new_net_17064;
	wire new_net_18746;
	wire new_net_16203;
	wire new_net_6119;
	wire new_net_17266;
	wire _0529_;
	wire _0193_;
	wire new_net_8611;
	wire new_net_16301;
	wire new_net_4997;
	wire new_net_9010;
	wire new_net_20772;
	wire new_net_1855;
	wire new_net_1400;
	wire new_net_4303;
	wire new_net_7265;
	wire new_net_8240;
	wire new_net_16311;
	wire new_net_8533;
	wire new_net_8606;
	wire new_net_10031;
	wire new_net_19631;
	wire new_net_6025;
	wire _0194_;
	wire _0530_;
	wire new_net_3102;
	wire new_net_9193;
	wire new_net_9625;
	wire _1680_;
	wire new_net_640;
	wire new_net_4664;
	wire new_net_4829;
	wire new_net_10037;
	wire new_net_19618;
	wire new_net_17934;
	wire new_net_7948;
	wire new_net_11288;
	wire _0195_;
	wire _0531_;
	wire new_net_10842;
	wire new_net_8607;
	wire new_net_11067;
	wire new_net_16305;
	wire new_net_870;
	wire new_net_19182;
	wire new_net_1398;
	wire new_net_4661;
	wire new_net_21185;
	wire new_net_5883;
	wire new_net_13183;
	wire new_net_17286;
	wire new_net_15134;
	wire new_net_15951;
	wire _0196_;
	wire new_net_637;
	wire _0532_;
	wire new_net_14255;
	wire new_net_17523;
	wire new_net_14113;
	wire _0560_;
	wire new_net_12375;
	wire new_net_12921;
	wire new_net_7738;
	wire new_net_17265;
	wire new_net_3093;
	wire new_net_4776;
	wire new_net_16202;
	wire new_net_9061;
	wire new_net_18226;
	wire new_net_12354;
	wire new_net_17699;
	wire new_net_10030;
	wire new_net_4803;
	wire new_net_9199;
	wire _0197_;
	wire _0533_;
	wire new_net_3094;
	wire new_net_8242;
	wire new_net_3906;
	wire new_net_9633;
	wire new_net_19632;
	wire new_net_14784;
	wire new_net_629;
	wire new_net_7962;
	wire new_net_20771;
	wire new_net_5506;
	wire new_net_1096;
	wire _0198_;
	wire _0534_;
	wire new_net_18985;
	wire new_net_4251;
	wire new_net_8613;
	wire new_net_11289;
	wire new_net_11068;
	wire new_net_9195;
	wire new_net_20803;
	wire new_net_3232;
	wire new_net_16940;
	wire _0535_;
	wire _0199_;
	wire new_net_18890;
	wire new_net_15752;
	wire new_net_19181;
	wire new_net_21184;
	wire new_net_21384;
	wire new_net_12797;
	wire new_net_15693;
	wire new_net_13184;
	wire new_net_17287;
	wire new_net_1093;
	wire new_net_3910;
	wire new_net_5170;
	wire new_net_15135;
	wire new_net_15952;
	wire new_net_14256;
	wire new_net_17524;
	wire new_net_12534;
	wire new_net_17889;
	wire new_net_18659;
	wire new_net_19189;
	wire new_net_4801;
	wire new_net_6021;
	wire new_net_16201;
	wire new_net_1401;
	wire _0536_;
	wire _0200_;
	wire new_net_8902;
	wire new_net_8235;
	wire new_net_17264;
	wire new_net_12179;
	wire new_net_12398;
	wire new_net_14707;
	wire new_net_14884;
	wire new_net_17636;
	wire new_net_6024;
	wire new_net_1092;
	wire new_net_3100;
	wire new_net_4297;
	wire new_net_4798;
	wire new_net_16310;
	wire new_net_18224;
	wire new_net_19611;
	wire new_net_19633;
	wire new_net_1089;
	wire _0537_;
	wire _0201_;
	wire new_net_1847;
	wire new_net_9874;
	wire new_net_8536;
	wire new_net_10843;
	wire new_net_4659;
	wire new_net_4773;
	wire new_net_20770;
	wire new_net_2921;
	wire new_net_634;
	wire new_net_3106;
	wire new_net_3909;
	wire new_net_4306;
	wire new_net_7959;
	wire new_net_21391;
	wire new_net_14511;
	wire new_net_14785;
	wire _0538_;
	wire _0202_;
	wire new_net_3748;
	wire new_net_11290;
	wire new_net_11069;
	wire new_net_20804;
	wire new_net_13695;
	wire new_net_1392;
	wire new_net_3753;
	wire new_net_4825;
	wire new_net_5511;
	wire new_net_8236;
	wire new_net_21183;
	wire new_net_11997;
	wire new_net_13185;
	wire new_net_17288;
	wire _0539_;
	wire _0203_;
	wire new_net_15136;
	wire new_net_15953;
	wire new_net_14257;
	wire new_net_17525;
	wire new_net_12535;
	wire new_net_14115;
	wire new_net_17909;
	wire new_net_17360;
	wire new_net_9200;
	wire new_net_16200;
	wire new_net_1391;
	wire new_net_4300;
	wire new_net_9872;
	wire new_net_17263;
	wire new_net_10035;
	wire new_net_18223;
	wire new_net_4771;
	wire new_net_1850;
	wire new_net_1086;
	wire _0204_;
	wire _0540_;
	wire new_net_9869;
	wire new_net_3328;
	wire new_net_6759;
	wire new_net_8604;
	wire new_net_19634;
	wire new_net_20301;
	wire new_net_4777;
	wire new_net_3442;
	wire new_net_8541;
	wire new_net_18048;
	wire new_net_4660;
	wire _0205_;
	wire _0541_;
	wire new_net_7951;
	wire new_net_7734;
	wire new_net_8975;
	wire new_net_4826;
	wire new_net_16306;
	wire new_net_19617;
	wire new_net_17986;
	wire new_net_9198;
	wire new_net_14786;
	wire new_net_1848;
	wire new_net_3099;
	wire new_net_4250;
	wire new_net_4299;
	wire new_net_9867;
	wire new_net_11291;
	wire new_net_7731;
	wire new_net_10844;
	wire new_net_2690;
	wire new_net_9630;
	wire new_net_8415;
	wire _0542_;
	wire new_net_5507;
	wire new_net_1854;
	wire _0206_;
	wire new_net_6756;
	wire new_net_7953;
	wire new_net_21182;
	wire new_net_9012;
	wire new_net_11757;
	wire new_net_12809;
	wire new_net_13186;
	wire new_net_17289;
	wire new_net_1402;
	wire new_net_3752;
	wire new_net_4301;
	wire new_net_4999;
	wire new_net_6125;
	wire new_net_14830;
	wire new_net_15656;
	wire new_net_18680;
	wire new_net_16199;
	wire _0543_;
	wire _0207_;
	wire new_net_3848;
	wire new_net_7946;
	wire new_net_17262;
	wire new_net_10032;
	wire new_net_19179;
	wire new_net_17620;
	wire new_net_3746;
	wire new_net_16309;
	wire new_net_19635;
	wire new_net_21389;
	wire new_net_18109;
	wire new_net_3097;
	wire new_net_9058;
	wire new_net_633;
	wire _0544_;
	wire _0208_;
	wire new_net_4830;
	wire new_net_18222;
	wire new_net_9007;
	wire new_net_9635;
	wire new_net_1853;
	wire new_net_1397;
	wire new_net_3512;
	wire new_net_6757;
	wire new_net_7954;
	wire new_net_18218;
	wire new_net_19653;
	wire new_net_3096;
	wire new_net_5002;
	wire new_net_9631;
	wire new_net_3849;
	wire new_net_14787;
	wire _0209_;
	wire _0545_;
	wire new_net_5733;
	wire new_net_8237;
	wire new_net_9873;
	wire new_net_18883;
	wire new_net_14498;
	wire new_net_9008;
	wire new_net_6018;
	wire new_net_7735;
	wire new_net_8531;
	wire new_net_10033;
	wire new_net_19616;
	wire new_net_21181;
	wire new_net_18371;
	wire new_net_4779;
	wire new_net_11758;
	wire new_net_12810;
	wire new_net_13187;
	wire _0210_;
	wire _0546_;
	wire new_net_3447;
	wire new_net_5505;
	wire new_net_17290;
	wire new_net_15138;
	wire new_net_15205;
	wire new_net_9192;
	wire new_net_1090;
	wire new_net_3514;
	wire new_net_4774;
	wire new_net_7268;
	wire new_net_16198;
	wire new_net_5726;
	wire new_net_9876;
	wire new_net_17261;
	wire new_net_5169;
	wire new_net_18747;
	wire new_net_21045;
	wire new_net_9009;
	wire new_net_1094;
	wire _0211_;
	wire _0547_;
	wire new_net_19178;
	wire new_net_19636;
	wire new_net_7270;
	wire new_net_8610;
	wire new_net_9014;
	wire new_net_17522;
	wire new_net_2738;
	wire new_net_643;
	wire _0548_;
	wire _0212_;
	wire new_net_3749;
	wire new_net_9870;
	wire new_net_19614;
	wire new_net_21153;
	wire new_net_17935;
	wire new_net_4248;
	wire new_net_11072;
	wire new_net_8414;
	wire new_net_14788;
	wire new_net_632;
	wire new_net_3908;
	wire new_net_11293;
	wire new_net_7957;
	wire new_net_10846;
	wire new_net_20807;
	wire new_net_9627;
	wire new_net_4806;
	wire _0549_;
	wire _0213_;
	wire new_net_3751;
	wire new_net_7945;
	wire new_net_19615;
	wire new_net_21180;
	wire new_net_21383;
	wire new_net_18407;
	wire new_net_16003;
	wire new_net_11759;
	wire new_net_12811;
	wire new_net_13188;
	wire new_net_3101;
	wire new_net_4302;
	wire new_net_17291;
	wire new_net_15139;
	wire new_net_15956;
	wire new_net_14260;
	wire new_net_12922;
	wire new_net_12376;
	wire new_net_3108;
	wire new_net_5001;
	wire new_net_4797;
	wire _0550_;
	wire _0214_;
	wire new_net_16197;
	wire new_net_17260;
	wire new_net_12355;
	wire new_net_16308;
	wire new_net_1095;
	wire new_net_1394;
	wire new_net_3281;
	wire new_net_4254;
	wire new_net_7950;
	wire new_net_6755;
	wire new_net_18221;
	wire new_net_19637;
	wire new_net_9596;
	wire new_net_16303;
	wire _0551_;
	wire new_net_630;
	wire _0215_;
	wire new_net_7733;
	wire new_net_19177;
	wire new_net_21388;
	wire new_net_7943;
	wire new_net_14195;
	wire new_net_14161;
	wire new_net_9628;
	wire new_net_14789;
	wire _0552_;
	wire _0216_;
	wire new_net_6017;
	wire new_net_7267;
	wire new_net_8243;
	wire new_net_11294;
	wire new_net_8537;
	wire new_net_10847;
	wire new_net_5729;
	wire new_net_7955;
	wire new_net_8241;
	wire new_net_18220;
	wire new_net_21179;
	wire new_net_18891;
	wire new_net_19241;
	wire new_net_15694;
	wire new_net_16004;
	wire new_net_9632;
	wire new_net_11760;
	wire new_net_12812;
	wire new_net_13189;
	wire new_net_1849;
	wire _0553_;
	wire _0217_;
	wire new_net_4298;
	wire new_net_17292;
	wire new_net_17890;
	wire new_net_18660;
	wire new_net_19190;
	wire new_net_8605;
	wire new_net_9194;
	wire new_net_3511;
	wire new_net_4775;
	wire new_net_4802;
	wire new_net_4998;
	wire new_net_16196;
	wire new_net_17259;
	wire new_net_7961;
	wire new_net_21177;
	wire new_net_12180;
	wire new_net_14708;
	wire new_net_5004;
	wire new_net_9196;
	wire new_net_1399;
	wire _0554_;
	wire _0218_;
	wire new_net_4304;
	wire new_net_5513;
	wire new_net_6020;
	wire new_net_17258;
	wire new_net_7737;
	wire new_net_11073;
	wire new_net_6016;
	wire new_net_7949;
	wire new_net_8535;
	wire new_net_20765;
	wire new_net_3171;
	wire new_net_16006;
	wire new_net_17436;
	wire new_net_4827;
	wire new_net_3098;
	wire new_net_9011;
	wire new_net_9062;
	wire _0219_;
	wire _0555_;
	wire new_net_16194;
	wire new_net_18219;
	wire new_net_19176;
	wire new_net_14790;
	wire new_net_4804;
	wire new_net_5510;
	wire new_net_6022;
	wire new_net_5731;
	wire new_net_7947;
	wire new_net_11295;
	wire new_net_10848;
	wire new_net_20809;
	wire new_net_20812;
	wire new_net_1857;
	wire new_net_3095;
	wire new_net_9063;
	wire new_net_9197;
	wire _0556_;
	wire _0220_;
	wire new_net_3907;
	wire new_net_21178;
	wire new_net_16484;
	wire new_net_14444;
	wire new_net_16520;
	wire new_net_11998;
	wire new_net_12540;
	wire new_net_14120;
	wire new_net_16005;
	wire new_net_11761;
	wire new_net_12813;
	wire new_net_13190;
	wire new_net_3905;
	wire new_net_4769;
	wire new_net_17293;
	wire new_net_15141;
	wire new_net_713;
	wire new_net_9370;
	wire new_net_15257;
	wire new_net_17361;
	wire new_net_4252;
	wire new_net_3513;
	wire new_net_8412;
	wire _0221_;
	wire _0557_;
	wire new_net_16195;
	wire new_net_6124;
	wire new_net_19613;
	wire new_net_21301;
	wire new_net_17648;
	wire new_net_16307;
	wire new_net_1097;
	wire new_net_1395;
	wire new_net_4823;
	wire new_net_19639;
	wire new_net_20302;
	wire new_net_18145;
	wire new_net_10029;
	wire _0222_;
	wire new_net_635;
	wire _0558_;
	wire new_net_8973;
	wire new_net_18047;
	wire new_net_3282;
	wire new_net_5508;
	wire new_net_9871;
	wire new_net_14133;
	wire new_net_17976;
	wire new_net_4329;
	wire new_net_8539;
	wire new_net_10849;
	wire new_net_8609;
	wire new_net_11074;
	wire new_net_4805;
	wire _0559_;
	wire _0223_;
	wire new_net_6122;
	wire new_net_11296;
	wire new_net_17987;
	wire new_net_17069;
	wire new_net_12831;
	wire new_net_12123;
	wire new_net_5083;
	wire new_net_10489;
	wire new_net_2337;
	wire new_net_3153;
	wire new_net_3344;
	wire new_net_3391;
	wire new_net_10235;
	wire new_net_20595;
	wire new_net_12986;
	wire new_net_14831;
	wire new_net_15657;
	wire _1379_;
	wire new_net_18681;
	wire new_net_7346;
	wire new_net_11796;
	wire new_net_6104;
	wire new_net_11951;
	wire new_net_12126;
	wire new_net_5845;
	wire new_net_12648;
	wire new_net_13286;
	wire new_net_15698;
	wire new_net_16963;
	wire new_net_17621;
	wire new_net_12125;
	wire new_net_3562;
	wire new_net_9351;
	wire new_net_10244;
	wire new_net_19795;
	wire new_net_19819;
	wire new_net_18110;
	wire new_net_2049;
	wire new_net_7651;
	wire _0351_;
	wire _0771_;
	wire new_net_3553;
	wire new_net_4146;
	wire new_net_7730;
	wire new_net_9343;
	wire new_net_19654;
	wire new_net_6604;
	wire new_net_7030;
	wire new_net_6365;
	wire _0352_;
	wire _0772_;
	wire new_net_19515;
	wire new_net_20124;
	wire new_net_20987;
	wire new_net_13562;
	wire new_net_14585;
	wire new_net_14499;
	wire new_net_5079;
	wire new_net_5837;
	wire new_net_10495;
	wire new_net_2200;
	wire new_net_8328;
	wire new_net_10439;
	wire new_net_13980;
	wire new_net_11075;
	wire new_net_11472;
	wire new_net_10234;
	wire new_net_17018;
	wire new_net_7340;
	wire _0353_;
	wire _0773_;
	wire new_net_9347;
	wire new_net_18454;
	wire new_net_20596;
	wire new_net_4075;
	wire new_net_12230;
	wire new_net_17066;
	wire new_net_2579;
	wire new_net_6902;
	wire new_net_15206;
	wire new_net_1900;
	wire new_net_13873;
	wire new_net_18748;
	wire new_net_11797;
	wire new_net_16964;
	wire new_net_11952;
	wire new_net_12649;
	wire new_net_13287;
	wire new_net_15699;
	wire new_net_11621;
	wire new_net_17295;
	wire new_net_9563;
	wire new_net_15014;
	wire new_net_20487;
	wire new_net_21046;
	wire new_net_13826;
	wire new_net_5051;
	wire new_net_5081;
	wire new_net_10496;
	wire _0354_;
	wire _0774_;
	wire new_net_2330;
	wire new_net_4148;
	wire new_net_3555;
	wire new_net_19796;
	wire new_net_19820;
	wire new_net_10245;
	wire new_net_14229;
	wire new_net_5801;
	wire new_net_12124;
	wire new_net_6358;
	wire new_net_21187;
	wire _1687_;
	wire new_net_2741;
	wire new_net_21154;
	wire new_net_7726;
	wire new_net_10236;
	wire new_net_14228;
	wire new_net_5043;
	wire new_net_2202;
	wire _0775_;
	wire _0355_;
	wire new_net_9158;
	wire new_net_3554;
	wire new_net_18312;
	wire new_net_12993;
	wire new_net_2487;
	wire new_net_17936;
	wire new_net_19516;
	wire new_net_20125;
	wire new_net_20988;
	wire new_net_11112;
	wire new_net_11390;
	wire new_net_5805;
	wire new_net_12122;
	wire _0356_;
	wire _0776_;
	wire new_net_13462;
	wire new_net_9567;
	wire new_net_5407;
	wire new_net_11076;
	wire new_net_10105;
	wire new_net_14424;
	wire new_net_18408;
	wire new_net_2197;
	wire new_net_3564;
	wire new_net_7655;
	wire new_net_7828;
	wire new_net_20597;
	wire _0567_;
	wire new_net_12377;
	wire new_net_12923;
	wire new_net_11798;
	wire new_net_11953;
	wire new_net_15700;
	wire new_net_9500;
	wire new_net_16965;
	wire _0357_;
	wire new_net_1098;
	wire new_net_12650;
	wire new_net_13288;
	wire _0777_;
	wire new_net_12356;
	wire new_net_17701;
	wire new_net_7029;
	wire new_net_9159;
	wire new_net_9435;
	wire new_net_13979;
	wire new_net_19797;
	wire new_net_19821;
	wire new_net_14230;
	wire new_net_13616;
	wire _0358_;
	wire new_net_6367;
	wire _0778_;
	wire new_net_18311;
	wire new_net_18463;
	wire new_net_19213;
	wire new_net_20447;
	wire new_net_7723;
	wire new_net_7347;
	wire new_net_2201;
	wire new_net_3418;
	wire new_net_10440;
	wire new_net_20451;
	wire new_net_2440;
	wire new_net_9342;
	wire _0779_;
	wire _0359_;
	wire new_net_2043;
	wire new_net_13173;
	wire new_net_10494;
	wire new_net_3159;
	wire new_net_19517;
	wire new_net_20126;
	wire new_net_20989;
	wire new_net_11113;
	wire new_net_11391;
	wire new_net_7362;
	wire new_net_12121;
	wire new_net_646;
	wire new_net_2042;
	wire new_net_17782;
	wire new_net_10442;
	wire new_net_9564;
	wire new_net_5404;
	wire new_net_18892;
	wire new_net_1310;
	wire new_net_15695;
	wire new_net_10238;
	wire new_net_10070;
	wire _0780_;
	wire _0360_;
	wire new_net_6357;
	wire new_net_18301;
	wire new_net_20598;
	wire new_net_17891;
	wire new_net_12444;
	wire new_net_9920;
	wire new_net_13833;
	wire new_net_18661;
	wire new_net_19191;
	wire new_net_10242;
	wire new_net_7366;
	wire new_net_10074;
	wire new_net_11799;
	wire new_net_11954;
	wire new_net_7024;
	wire new_net_649;
	wire new_net_5843;
	wire new_net_12651;
	wire new_net_13289;
	wire new_net_12181;
	wire new_net_7532;
	wire new_net_645;
	wire new_net_7341;
	wire new_net_10076;
	wire new_net_7022;
	wire new_net_9499;
	wire _0361_;
	wire new_net_7656;
	wire _0781_;
	wire new_net_2338;
	wire new_net_14231;
	wire new_net_13617;
	wire new_net_7657;
	wire new_net_16007;
	wire new_net_17437;
	wire new_net_3565;
	wire new_net_5044;
	wire _0362_;
	wire new_net_10492;
	wire _0782_;
	wire new_net_14613;
	wire new_net_648;
	wire new_net_2199;
	wire new_net_5406;
	wire new_net_6106;
	wire new_net_9156;
	wire new_net_19518;
	wire new_net_20127;
	wire new_net_20990;
	wire new_net_21255;
	wire new_net_13697;
	wire new_net_11078;
	wire new_net_11475;
	wire new_net_10241;
	wire new_net_11114;
	wire new_net_11392;
	wire new_net_5798;
	wire _0783_;
	wire _0363_;
	wire new_net_2047;
	wire new_net_14492;
	wire new_net_14445;
	wire new_net_16521;
	wire new_net_7369;
	wire new_net_3155;
	wire new_net_5844;
	wire new_net_6107;
	wire new_net_8325;
	wire new_net_1993;
	wire new_net_20599;
	wire new_net_15258;
	wire new_net_17362;
	wire new_net_15017;
	wire new_net_15489;
	wire new_net_9344;
	wire new_net_5802;
	wire new_net_11800;
	wire new_net_11955;
	wire _0784_;
	wire _0364_;
	wire new_net_2048;
	wire new_net_6361;
	wire new_net_12956;
	wire _0980_;
	wire new_net_13897;
	wire new_net_17649;
	wire new_net_404;
	wire new_net_9346;
	wire new_net_2206;
	wire new_net_3151;
	wire new_net_7825;
	wire new_net_13977;
	wire new_net_18456;
	wire new_net_19799;
	wire new_net_19823;
	wire new_net_15137;
	wire new_net_20303;
	wire new_net_14232;
	wire new_net_3345;
	wire new_net_13618;
	wire _0785_;
	wire _0365_;
	wire new_net_1101;
	wire new_net_2052;
	wire new_net_3152;
	wire new_net_9566;
	wire new_net_18046;
	wire new_net_9502;
	wire new_net_9162;
	wire new_net_18310;
	wire new_net_18462;
	wire new_net_14134;
	wire new_net_17975;
	wire new_net_17988;
	wire new_net_3416;
	wire new_net_5401;
	wire _0366_;
	wire new_net_1104;
	wire new_net_9505;
	wire _0786_;
	wire new_net_3157;
	wire new_net_4147;
	wire new_net_19519;
	wire new_net_20128;
	wire new_net_11079;
	wire new_net_11476;
	wire new_net_11115;
	wire new_net_11393;
	wire new_net_2331;
	wire new_net_7026;
	wire new_net_6360;
	wire new_net_18776;
	wire new_net_20374;
	wire new_net_17070;
	wire new_net_2198;
	wire new_net_7728;
	wire new_net_5807;
	wire _0367_;
	wire new_net_1110;
	wire _0787_;
	wire new_net_12832;
	wire new_net_5050;
	wire new_net_9497;
	wire new_net_12119;
	wire new_net_21333;
	wire new_net_12987;
	wire new_net_14832;
	wire new_net_15658;
	wire new_net_312;
	wire new_net_15018;
	wire new_net_15490;
	wire new_net_13291;
	wire new_net_15703;
	wire new_net_16968;
	wire new_net_11801;
	wire new_net_11956;
	wire new_net_3156;
	wire new_net_5408;
	wire new_net_5840;
	wire new_net_12893;
	wire new_net_18682;
	wire new_net_7725;
	wire new_net_9350;
	wire new_net_5803;
	wire _0788_;
	wire _0368_;
	wire new_net_12120;
	wire new_net_15356;
	wire new_net_13976;
	wire new_net_19800;
	wire new_net_19824;
	wire new_net_18111;
	wire new_net_10493;
	wire new_net_7729;
	wire new_net_14233;
	wire new_net_652;
	wire new_net_2038;
	wire new_net_3160;
	wire new_net_5080;
	wire new_net_13619;
	wire new_net_5842;
	wire new_net_5709;
	wire new_net_9349;
	wire _0369_;
	wire _0789_;
	wire new_net_8326;
	wire new_net_19655;
	wire new_net_15994;
	wire new_net_5048;
	wire new_net_5804;
	wire new_net_7368;
	wire new_net_19266;
	wire new_net_19520;
	wire new_net_20129;
	wire new_net_20992;
	wire new_net_21257;
	wire new_net_13561;
	wire new_net_14586;
	wire new_net_14500;
	wire new_net_11116;
	wire new_net_11394;
	wire new_net_10497;
	wire new_net_6105;
	wire new_net_9430;
	wire new_net_11080;
	wire _0370_;
	wire _0790_;
	wire new_net_11477;
	wire new_net_20375;
	wire new_net_12118;
	wire new_net_9431;
	wire new_net_5084;
	wire new_net_7345;
	wire new_net_17019;
	wire new_net_10446;
	wire new_net_20601;
	wire new_net_3150;
	wire new_net_11620;
	wire new_net_12231;
	wire new_net_17067;
	wire new_net_11802;
	wire new_net_3548;
	wire new_net_15019;
	wire new_net_13292;
	wire new_net_15704;
	wire new_net_16969;
	wire new_net_11957;
	wire new_net_17300;
	wire _0371_;
	wire new_net_9523;
	wire new_net_13874;
	wire new_net_18749;
	wire new_net_21047;
	wire new_net_13975;
	wire new_net_5797;
	wire new_net_6359;
	wire new_net_10437;
	wire new_net_19801;
	wire new_net_19825;
	wire new_net_3550;
	wire new_net_7360;
	wire new_net_10069;
	wire _0372_;
	wire _0792_;
	wire new_net_15923;
	wire new_net_13620;
	wire new_net_18206;
	wire new_net_20449;
	wire new_net_15447;
	wire new_net_9568;
	wire new_net_3556;
	wire new_net_21155;
	wire new_net_12994;
	wire new_net_17937;
	wire new_net_651;
	wire new_net_5800;
	wire new_net_3563;
	wire new_net_2204;
	wire _0373_;
	wire _0793_;
	wire new_net_19521;
	wire new_net_20130;
	wire new_net_20993;
	wire new_net_21258;
	wire new_net_18450;
	wire new_net_11081;
	wire new_net_11478;
	wire new_net_11117;
	wire new_net_11395;
	wire new_net_14234;
	wire new_net_4149;
	wire new_net_4230;
	wire new_net_10438;
	wire new_net_20376;
	wire new_net_14425;
	wire _1449_;
	wire new_net_3557;
	wire new_net_10071;
	wire new_net_2205;
	wire _0374_;
	wire new_net_12117;
	wire _0794_;
	wire new_net_9161;
	wire new_net_18455;
	wire new_net_20602;
	wire new_net_12924;
	wire new_net_15020;
	wire new_net_15492;
	wire new_net_17301;
	wire new_net_7344;
	wire new_net_11803;
	wire new_net_9433;
	wire new_net_11958;
	wire new_net_1099;
	wire new_net_2335;
	wire new_net_3560;
	wire new_net_8974;
	wire new_net_12357;
	wire new_net_13974;
	wire new_net_3419;
	wire new_net_3551;
	wire new_net_7342;
	wire new_net_17702;
	wire new_net_7829;
	wire new_net_2332;
	wire _0375_;
	wire new_net_5085;
	wire _0795_;
	wire new_net_13621;
	wire new_net_3561;
	wire new_net_7361;
	wire new_net_7724;
	wire new_net_10240;
	wire new_net_20448;
	wire new_net_9341;
	wire new_net_7370;
	wire new_net_1103;
	wire _0796_;
	wire _0376_;
	wire new_net_5045;
	wire new_net_7027;
	wire new_net_10498;
	wire new_net_19448;
	wire new_net_14163;
	wire new_net_9348;
	wire new_net_1109;
	wire new_net_7364;
	wire new_net_7722;
	wire new_net_9503;
	wire new_net_18308;
	wire new_net_18460;
	wire new_net_19522;
	wire new_net_20131;
	wire new_net_20994;
	wire new_net_13174;
	wire new_net_2561;
	wire new_net_11082;
	wire new_net_11479;
	wire new_net_5235;
	wire new_net_7727;
	wire new_net_11118;
	wire new_net_11396;
	wire new_net_7365;
	wire _0377_;
	wire new_net_1106;
	wire new_net_2203;
	wire new_net_2614;
	wire new_net_16943;
	wire new_net_17783;
	wire new_net_18893;
	wire new_net_11292;
	wire new_net_18501;
	wire new_net_15696;
	wire new_net_12800;
	wire new_net_9559;
	wire new_net_9501;
	wire new_net_5799;
	wire new_net_5052;
	wire new_net_7028;
	wire new_net_12116;
	wire new_net_20603;
	wire new_net_17892;
	wire new_net_12445;
	wire new_net_18662;
	wire new_net_19192;
	wire new_net_16971;
	wire new_net_15021;
	wire new_net_15493;
	wire new_net_7531;
	wire new_net_7363;
	wire new_net_11804;
	wire _0378_;
	wire new_net_1102;
	wire new_net_11959;
	wire new_net_7023;
	wire new_net_12182;
	wire new_net_13973;
	wire new_net_1107;
	wire new_net_7339;
	wire new_net_9163;
	wire new_net_10441;
	wire new_net_18453;
	wire new_net_19803;
	wire new_net_3549;
	wire new_net_14235;
	wire _0379_;
	wire new_net_3558;
	wire new_net_6109;
	wire new_net_13622;
	wire new_net_7658;
	wire _0799_;
	wire new_net_16008;
	wire new_net_17438;
	wire new_net_2039;
	wire new_net_2336;
	wire new_net_5049;
	wire new_net_10243;
	wire _0800_;
	wire _0380_;
	wire new_net_2040;
	wire new_net_16691;
	wire new_net_19523;
	wire new_net_20132;
	wire new_net_20995;
	wire new_net_21260;
	wire new_net_14514;
	wire new_net_18958;
	wire new_net_20814;
	wire new_net_16580;
	wire new_net_13698;
	wire new_net_9434;
	wire new_net_11083;
	wire new_net_11480;
	wire new_net_2207;
	wire new_net_9498;
	wire new_net_11119;
	wire new_net_11397;
	wire new_net_20378;
	wire new_net_14446;
	wire new_net_16522;
	wire new_net_12115;
	wire new_net_10072;
	wire new_net_7343;
	wire new_net_3347;
	wire _0801_;
	wire _0381_;
	wire new_net_10444;
	wire new_net_8876;
	wire new_net_20604;
	wire new_net_17363;
	wire new_net_15707;
	wire new_net_9569;
	wire new_net_16972;
	wire new_net_14238;
	wire new_net_11960;
	wire new_net_10073;
	wire new_net_9429;
	wire new_net_12657;
	wire new_net_15022;
	wire new_net_11805;
	wire new_net_21303;
	wire new_net_17650;
	wire new_net_13972;
	wire _0802_;
	wire new_net_2334;
	wire _0382_;
	wire new_net_5047;
	wire new_net_7025;
	wire new_net_19804;
	wire new_net_20304;
	wire new_net_14236;
	wire new_net_13623;
	wire new_net_10488;
	wire new_net_18306;
	wire new_net_18458;
	wire new_net_9157;
	wire new_net_10443;
	wire new_net_5236;
	wire _0803_;
	wire _0383_;
	wire new_net_1105;
	wire new_net_8977;
	wire new_net_18045;
	wire new_net_11929;
	wire new_net_14135;
	wire new_net_8327;
	wire new_net_2050;
	wire new_net_3158;
	wire new_net_9496;
	wire new_net_5082;
	wire new_net_19524;
	wire new_net_20133;
	wire new_net_20996;
	wire new_net_17989;
	wire new_net_21261;
	wire new_net_12782;
	wire new_net_11084;
	wire new_net_11481;
	wire new_net_11120;
	wire new_net_11398;
	wire new_net_10075;
	wire new_net_650;
	wire _0804_;
	wire _0384_;
	wire new_net_5078;
	wire new_net_12688;
	wire new_net_13480;
	wire new_net_2044;
	wire new_net_20605;
	wire new_net_17071;
	wire new_net_12833;
	wire new_net_12988;
	wire new_net_14833;
	wire new_net_15659;
	wire _1386_;
	wire new_net_11630;
	wire new_net_17304;
	wire new_net_9560;
	wire new_net_5405;
	wire new_net_15023;
	wire new_net_15495;
	wire new_net_11806;
	wire _0805_;
	wire _0385_;
	wire new_net_11961;
	wire new_net_18683;
	wire new_net_12894;
	wire new_net_15344;
	wire new_net_18650;
	wire new_net_13971;
	wire new_net_4231;
	wire new_net_5403;
	wire new_net_9504;
	wire new_net_18302;
	wire new_net_19269;
	wire new_net_19805;
	wire new_net_15357;
	wire new_net_4227;
	wire new_net_14237;
	wire new_net_3390;
	wire new_net_7348;
	wire _0806_;
	wire _0386_;
	wire new_net_13624;
	wire new_net_20476;
	wire new_net_9345;
	wire new_net_2041;
	wire new_net_5402;
	wire new_net_12471;
	wire new_net_19829;
	wire new_net_16431;
	wire new_net_19656;
	wire new_net_13969;
	wire _0807_;
	wire _0387_;
	wire new_net_6108;
	wire new_net_10457;
	wire new_net_2045;
	wire new_net_19270;
	wire new_net_19525;
	wire new_net_7440;
	wire new_net_20134;
	wire new_net_14587;
	wire new_net_18881;
	wire new_net_11085;
	wire new_net_11482;
	wire new_net_11399;
	wire new_net_2333;
	wire new_net_1100;
	wire new_net_9432;
	wire new_net_13626;
	wire new_net_16973;
	wire new_net_20380;
	wire _0808_;
	wire new_net_10068;
	wire _0388_;
	wire new_net_6364;
	wire new_net_7653;
	wire new_net_20606;
	wire new_net_1684;
	wire new_net_17020;
	wire new_net_1757;
	wire new_net_12232;
	wire new_net_17068;
	wire new_net_12659;
	wire new_net_13297;
	wire new_net_11631;
	wire new_net_17305;
	wire new_net_15024;
	wire new_net_15496;
	wire new_net_1111;
	wire new_net_5839;
	wire new_net_11807;
	wire new_net_15709;
	wire new_net_15208;
	wire new_net_21048;
	wire new_net_6356;
	wire new_net_13970;
	wire _0389_;
	wire new_net_1108;
	wire _0809_;
	wire new_net_3343;
	wire new_net_3559;
	wire new_net_19806;
	wire new_net_7830;
	wire new_net_2046;
	wire new_net_644;
	wire new_net_3394;
	wire new_net_7367;
	wire new_net_13625;
	wire new_net_15924;
	wire new_net_18207;
	wire new_net_15448;
	wire new_net_7654;
	wire new_net_10491;
	wire new_net_4151;
	wire new_net_9561;
	wire new_net_3552;
	wire new_net_4226;
	wire new_net_10239;
	wire new_net_11121;
	wire _0390_;
	wire _0810_;
	wire new_net_21156;
	wire new_net_12995;
	wire new_net_17938;
	wire new_net_7659;
	wire new_net_7419;
	wire new_net_9352;
	wire new_net_10237;
	wire new_net_3427;
	wire new_net_4145;
	wire new_net_4228;
	wire new_net_19526;
	wire new_net_20135;
	wire new_net_20998;
	wire new_net_6363;
	wire new_net_10445;
	wire new_net_9562;
	wire new_net_11086;
	wire new_net_11400;
	wire _0391_;
	wire _0811_;
	wire new_net_5806;
	wire new_net_19271;
	wire new_net_20381;
	wire _0574_;
	wire new_net_12161;
	wire new_net_12379;
	wire new_net_12925;
	wire new_net_7970;
	wire new_net_6897;
	wire new_net_2514;
	wire new_net_1383;
	wire new_net_1832;
	wire new_net_12358;
	wire new_net_3763;
	wire new_net_17703;
	wire new_net_16253;
	wire new_net_7770;
	wire new_net_17531;
	wire new_net_16420;
	wire new_net_14391;
	wire new_net_17318;
	wire new_net_12245;
	wire new_net_12352;
	wire new_net_15025;
	wire new_net_13639;
	wire new_net_3115;
	wire new_net_19938;
	wire new_net_6559;
	wire new_net_210;
	wire new_net_3265;
	wire new_net_7409;
	wire new_net_18619;
	wire new_net_8517;
	wire new_net_8030;
	wire _1569_;
	wire new_net_14198;
	wire new_net_1825;
	wire _1359_;
	wire new_net_212;
	wire new_net_1390;
	wire new_net_10279;
	wire new_net_6511;
	wire new_net_21247;
	wire new_net_5832;
	wire new_net_7819;
	wire new_net_6555;
	wire new_net_7473;
	wire new_net_2515;
	wire new_net_5927;
	wire _0986_;
	wire new_net_19746;
	wire new_net_13175;
	wire new_net_21467;
	wire new_net_2554;
	wire _1570_;
	wire _1360_;
	wire new_net_311;
	wire new_net_21264;
	wire new_net_2625;
	wire new_net_16944;
	wire new_net_18894;
	wire new_net_15756;
	wire new_net_18502;
	wire new_net_12801;
	wire new_net_15697;
	wire new_net_15687;
	wire new_net_8031;
	wire new_net_11087;
	wire new_net_11297;
	wire new_net_4395;
	wire new_net_7064;
	wire new_net_7968;
	wire new_net_9225;
	wire new_net_10804;
	wire new_net_9981;
	wire new_net_17893;
	wire new_net_17333;
	wire new_net_13835;
	wire new_net_18663;
	wire new_net_19193;
	wire new_net_3917;
	wire new_net_3936;
	wire _1571_;
	wire _1361_;
	wire new_net_200;
	wire new_net_666;
	wire new_net_18618;
	wire new_net_12183;
	wire new_net_12057;
	wire new_net_12791;
	wire new_net_14392;
	wire new_net_16587;
	wire new_net_12981;
	wire new_net_14826;
	wire new_net_15652;
	wire new_net_16254;
	wire new_net_16987;
	wire new_net_12246;
	wire new_net_21378;
	wire new_net_3928;
	wire new_net_2779;
	wire _1362_;
	wire new_net_1388;
	wire _1572_;
	wire new_net_16009;
	wire new_net_17439;
	wire new_net_18632;
	wire new_net_310;
	wire new_net_2775;
	wire new_net_9223;
	wire new_net_8789;
	wire new_net_19340;
	wire new_net_19736;
	wire new_net_14611;
	wire new_net_16715;
	wire new_net_19450;
	wire new_net_5456;
	wire new_net_7582;
	wire new_net_8520;
	wire _1363_;
	wire new_net_818;
	wire new_net_1384;
	wire new_net_2772;
	wire _1573_;
	wire new_net_3264;
	wire new_net_9226;
	wire new_net_21468;
	wire new_net_16581;
	wire new_net_9977;
	wire new_net_8518;
	wire new_net_2124;
	wire new_net_2520;
	wire new_net_21265;
	wire new_net_14447;
	wire new_net_16523;
	wire _1364_;
	wire _1574_;
	wire new_net_3915;
	wire new_net_11088;
	wire new_net_11298;
	wire new_net_10805;
	wire new_net_16421;
	wire new_net_12447;
	wire new_net_15260;
	wire new_net_17364;
	wire new_net_823;
	wire new_net_1824;
	wire new_net_7435;
	wire new_net_19341;
	wire new_net_12958;
	wire _0987_;
	wire new_net_17651;
	wire new_net_12011;
	wire new_net_13229;
	wire new_net_12058;
	wire new_net_12792;
	wire new_net_6956;
	wire new_net_12982;
	wire new_net_14827;
	wire new_net_15653;
	wire new_net_16255;
	wire new_net_16988;
	wire new_net_20305;
	wire new_net_16903;
	wire new_net_17256;
	wire new_net_3272;
	wire new_net_6558;
	wire new_net_14308;
	wire new_net_16847;
	wire new_net_18044;
	wire new_net_7963;
	wire new_net_6551;
	wire _1366_;
	wire new_net_213;
	wire _1576_;
	wire new_net_3267;
	wire new_net_6510;
	wire new_net_11930;
	wire new_net_14136;
	wire new_net_16662;
	wire new_net_305;
	wire new_net_1828;
	wire new_net_6517;
	wire new_net_6560;
	wire new_net_7818;
	wire new_net_17990;
	wire new_net_21469;
	wire new_net_3392;
	wire new_net_12103;
	wire new_net_14521;
	wire new_net_12783;
	wire new_net_6948;
	wire new_net_6556;
	wire _1367_;
	wire new_net_206;
	wire new_net_309;
	wire _1577_;
	wire new_net_2122;
	wire new_net_21266;
	wire new_net_13481;
	wire new_net_9983;
	wire new_net_2524;
	wire new_net_6954;
	wire new_net_11089;
	wire new_net_11299;
	wire new_net_10806;
	wire new_net_12834;
	wire new_net_21335;
	wire new_net_12989;
	wire new_net_14834;
	wire new_net_15660;
	wire _1368_;
	wire _1578_;
	wire new_net_3938;
	wire new_net_15166;
	wire new_net_9835;
	wire new_net_18684;
	wire new_net_12895;
	wire new_net_1348;
	wire new_net_12012;
	wire new_net_13230;
	wire new_net_13642;
	wire new_net_12059;
	wire new_net_12793;
	wire new_net_14394;
	wire new_net_15689;
	wire new_net_16589;
	wire new_net_7772;
	wire new_net_12983;
	wire new_net_15358;
	wire new_net_7967;
	wire new_net_17255;
	wire _1369_;
	wire new_net_202;
	wire new_net_2777;
	wire _1579_;
	wire new_net_3338;
	wire new_net_6145;
	wire new_net_16088;
	wire new_net_17543;
	wire new_net_11890;
	wire new_net_12470;
	wire new_net_5829;
	wire new_net_7964;
	wire new_net_2125;
	wire new_net_7065;
	wire new_net_19737;
	wire new_net_16432;
	wire new_net_19657;
	wire new_net_15996;
	wire _1370_;
	wire new_net_822;
	wire new_net_3271;
	wire new_net_6208;
	wire _1580_;
	wire new_net_6514;
	wire new_net_21470;
	wire new_net_13559;
	wire new_net_14588;
	wire new_net_18880;
	wire new_net_9976;
	wire new_net_8525;
	wire new_net_2771;
	wire new_net_3273;
	wire new_net_3944;
	wire new_net_7476;
	wire new_net_9221;
	wire new_net_21267;
	wire new_net_8521;
	wire new_net_9890;
	wire _1581_;
	wire _1371_;
	wire new_net_14307;
	wire new_net_11090;
	wire new_net_11300;
	wire new_net_10807;
	wire new_net_11622;
	wire new_net_6899;
	wire new_net_8027;
	wire new_net_2118;
	wire new_net_211;
	wire new_net_18617;
	wire new_net_15209;
	wire new_net_21049;
	wire new_net_11824;
	wire new_net_12013;
	wire new_net_13231;
	wire new_net_13643;
	wire new_net_5836;
	wire new_net_8526;
	wire new_net_12060;
	wire new_net_12794;
	wire new_net_14395;
	wire new_net_15690;
	wire new_net_15509;
	wire new_net_6894;
	wire new_net_9727;
	wire new_net_17254;
	wire new_net_19339;
	wire new_net_19744;
	wire new_net_15925;
	wire new_net_18208;
	wire new_net_14258;
	wire new_net_17526;
	wire new_net_17503;
	wire new_net_5834;
	wire new_net_8522;
	wire new_net_6953;
	wire _1583_;
	wire _1373_;
	wire new_net_1826;
	wire new_net_21157;
	wire new_net_12996;
	wire new_net_17939;
	wire new_net_6509;
	wire new_net_8137;
	wire new_net_5827;
	wire new_net_2129;
	wire new_net_817;
	wire new_net_4399;
	wire new_net_21471;
	wire new_net_5932;
	wire new_net_7771;
	wire _1584_;
	wire new_net_2526;
	wire _1374_;
	wire new_net_308;
	wire new_net_7475;
	wire new_net_21268;
	wire new_net_18410;
	wire new_net_14306;
	wire new_net_8026;
	wire new_net_5826;
	wire new_net_9729;
	wire new_net_11091;
	wire new_net_11301;
	wire new_net_9227;
	wire new_net_10808;
	wire new_net_19743;
	wire new_net_5608;
	wire new_net_17033;
	wire new_net_12160;
	wire new_net_9979;
	wire new_net_4957;
	wire _1585_;
	wire _1375_;
	wire new_net_209;
	wire new_net_2776;
	wire new_net_9723;
	wire new_net_7406;
	wire new_net_21297;
	wire new_net_12359;
	wire new_net_11825;
	wire new_net_12014;
	wire new_net_13232;
	wire new_net_13644;
	wire new_net_7973;
	wire new_net_12061;
	wire new_net_12795;
	wire new_net_15691;
	wire new_net_7773;
	wire new_net_12985;
	wire new_net_17704;
	wire new_net_17144;
	wire new_net_9975;
	wire new_net_7972;
	wire new_net_6896;
	wire new_net_7768;
	wire _1586_;
	wire new_net_2126;
	wire _1376_;
	wire new_net_204;
	wire new_net_4657;
	wire new_net_17253;
	wire new_net_5831;
	wire new_net_2121;
	wire new_net_3920;
	wire new_net_14165;
	wire new_net_7822;
	wire _1587_;
	wire _1377_;
	wire new_net_4397;
	wire new_net_4953;
	wire new_net_21472;
	wire new_net_13176;
	wire new_net_11750;
	wire new_net_8134;
	wire new_net_7821;
	wire new_net_669;
	wire new_net_3587;
	wire new_net_4958;
	wire new_net_18642;
	wire new_net_21269;
	wire new_net_14380;
	wire new_net_16945;
	wire new_net_17785;
	wire new_net_18895;
	wire new_net_15757;
	wire new_net_18503;
	wire new_net_9978;
	wire new_net_14396;
	wire new_net_16591;
	wire new_net_4954;
	wire _1588_;
	wire _1378_;
	wire new_net_2778;
	wire new_net_4394;
	wire new_net_11092;
	wire new_net_11302;
	wire new_net_17894;
	wire new_net_17334;
	wire new_net_820;
	wire new_net_7769;
	wire new_net_7965;
	wire new_net_13836;
	wire new_net_18614;
	wire new_net_18664;
	wire new_net_19194;
	wire new_net_19741;
	wire new_net_12184;
	wire new_net_14305;
	wire new_net_16425;
	wire new_net_17513;
	wire new_net_8135;
	wire new_net_11826;
	wire new_net_5935;
	wire new_net_9980;
	wire new_net_12015;
	wire new_net_13233;
	wire new_net_13645;
	wire new_net_7767;
	wire new_net_8029;
	wire new_net_214;
	wire new_net_17252;
	wire new_net_7470;
	wire new_net_17486;
	wire new_net_18615;
	wire new_net_4984;
	wire new_net_16010;
	wire new_net_17440;
	wire new_net_7405;
	wire _1380_;
	wire new_net_1389;
	wire _1590_;
	wire new_net_2120;
	wire new_net_17993;
	wire new_net_16716;
	wire new_net_19447;
	wire new_net_3916;
	wire new_net_4392;
	wire new_net_4956;
	wire new_net_21473;
	wire new_net_14516;
	wire new_net_20816;
	wire new_net_16670;
	wire new_net_16582;
	wire _1381_;
	wire new_net_824;
	wire _1591_;
	wire new_net_19735;
	wire new_net_21270;
	wire new_net_10490;
	wire new_net_14448;
	wire new_net_16524;
	wire new_net_7404;
	wire new_net_10810;
	wire new_net_9984;
	wire new_net_215;
	wire new_net_1386;
	wire new_net_7474;
	wire new_net_11093;
	wire new_net_11303;
	wire new_net_20793;
	wire new_net_12448;
	wire _1382_;
	wire new_net_208;
	wire new_net_825;
	wire _1592_;
	wire new_net_9892;
	wire new_net_17652;
	wire new_net_7407;
	wire new_net_14304;
	wire new_net_16426;
	wire new_net_17514;
	wire new_net_6515;
	wire new_net_11827;
	wire new_net_12016;
	wire new_net_13234;
	wire new_net_13646;
	wire new_net_8519;
	wire new_net_15140;
	wire new_net_20306;
	wire new_net_21189;
	wire new_net_14303;
	wire new_net_9982;
	wire new_net_4396;
	wire new_net_5828;
	wire _1383_;
	wire _1593_;
	wire new_net_3268;
	wire new_net_3942;
	wire new_net_8351;
	wire new_net_17251;
	wire new_net_7069;
	wire new_net_16848;
	wire new_net_6893;
	wire new_net_7817;
	wire new_net_2128;
	wire new_net_672;
	wire new_net_3589;
	wire new_net_5833;
	wire new_net_8981;
	wire new_net_18043;
	wire new_net_879;
	wire new_net_11931;
	wire new_net_14137;
	wire _1384_;
	wire new_net_2768;
	wire _1594_;
	wire new_net_3940;
	wire new_net_18855;
	wire new_net_21474;
	wire new_net_17991;
	wire new_net_12104;
	wire new_net_14522;
	wire new_net_12784;
	wire new_net_7411;
	wire new_net_6951;
	wire new_net_1827;
	wire new_net_2769;
	wire new_net_671;
	wire new_net_2516;
	wire new_net_3926;
	wire new_net_21271;
	wire new_net_12690;
	wire new_net_10811;
	wire new_net_6516;
	wire new_net_8028;
	wire _1385_;
	wire new_net_676;
	wire _1595_;
	wire new_net_6557;
	wire new_net_11094;
	wire new_net_11304;
	wire new_net_20794;
	wire new_net_17073;
	wire new_net_12990;
	wire new_net_14835;
	wire new_net_15661;
	wire new_net_7414;
	wire new_net_9228;
	wire new_net_7765;
	wire new_net_7816;
	wire new_net_2774;
	wire new_net_2513;
	wire new_net_3934;
	wire new_net_7066;
	wire new_net_18609;
	wire new_net_15167;
	wire new_net_17413;
	wire new_net_18685;
	wire new_net_18956;
	wire new_net_12896;
	wire new_net_15346;
	wire new_net_16427;
	wire new_net_17515;
	wire new_net_11828;
	wire new_net_12017;
	wire new_net_13235;
	wire new_net_13647;
	wire new_net_8516;
	wire new_net_12064;
	wire new_net_12798;
	wire new_net_14398;
	wire new_net_15359;
	wire new_net_207;
	wire new_net_670;
	wire new_net_1381;
	wire new_net_8202;
	wire new_net_2119;
	wire new_net_3590;
	wire new_net_5835;
	wire new_net_6553;
	wire new_net_17250;
	wire new_net_14333;
	wire new_net_16089;
	wire new_net_3270;
	wire new_net_7766;
	wire _1387_;
	wire new_net_2773;
	wire _1597_;
	wire new_net_16433;
	wire new_net_2132;
	wire new_net_3922;
	wire new_net_6552;
	wire new_net_18613;
	wire new_net_21475;
	wire new_net_20885;
	wire new_net_13558;
	wire new_net_14589;
	wire new_net_18879;
	wire new_net_7063;
	wire new_net_7410;
	wire new_net_9222;
	wire new_net_6947;
	wire _1598_;
	wire new_net_2130;
	wire _1388_;
	wire new_net_21272;
	wire new_net_1739;
	wire new_net_9659;
	wire new_net_11095;
	wire new_net_11305;
	wire new_net_7412;
	wire new_net_10812;
	wire new_net_4393;
	wire new_net_1830;
	wire new_net_9725;
	wire new_net_20795;
	wire new_net_11623;
	wire new_net_3269;
	wire new_net_4398;
	wire new_net_6898;
	wire _1599_;
	wire _1389_;
	wire new_net_665;
	wire new_net_19740;
	wire new_net_15210;
	wire new_net_17720;
	wire new_net_21050;
	wire new_net_15932;
	wire new_net_17540;
	wire new_net_16428;
	wire new_net_17516;
	wire new_net_11829;
	wire new_net_12018;
	wire new_net_13236;
	wire new_net_13648;
	wire new_net_12065;
	wire new_net_12799;
	wire new_net_15510;
	wire new_net_17709;
	wire new_net_7472;
	wire new_net_8136;
	wire _1600_;
	wire _1390_;
	wire new_net_302;
	wire new_net_17249;
	wire new_net_19338;
	wire new_net_15926;
	wire new_net_18209;
	wire new_net_6761;
	wire new_net_14259;
	wire new_net_17527;
	wire new_net_9220;
	wire new_net_14302;
	wire new_net_677;
	wire new_net_5830;
	wire _1394_;
	wire new_net_301;
	wire new_net_10052;
	wire new_net_19658;
	wire new_net_9168;
	wire new_net_9985;
	wire _1601_;
	wire _1391_;
	wire new_net_303;
	wire new_net_4955;
	wire new_net_12997;
	wire new_net_17940;
	wire new_net_21476;
	wire new_net_7562;
	wire new_net_4952;
	wire new_net_2517;
	wire new_net_1382;
	wire new_net_21273;
	wire new_net_8437;
	wire new_net_13466;
	wire new_net_11096;
	wire new_net_11306;
	wire new_net_10813;
	wire new_net_6513;
	wire new_net_5930;
	wire new_net_8032;
	wire _1602_;
	wire _1392_;
	wire new_net_12360;
	wire new_net_18411;
	wire new_net_17034;
	wire new_net_19138;
	wire _0581_;
	wire new_net_3266;
	wire new_net_7434;
	wire new_net_2519;
	wire new_net_2131;
	wire new_net_203;
	wire new_net_306;
	wire new_net_3930;
	wire new_net_12159;
	wire new_net_12381;
	wire new_net_12927;
	wire new_net_20751;
	wire new_net_13649;
	wire new_net_15933;
	wire new_net_17541;
	wire new_net_16429;
	wire new_net_17517;
	wire new_net_11830;
	wire new_net_16595;
	wire new_net_5931;
	wire new_net_12019;
	wire new_net_13237;
	wire new_net_17705;
	wire new_net_15461;
	wire new_net_17145;
	wire new_net_5933;
	wire new_net_3924;
	wire new_net_5825;
	wire new_net_17248;
	wire new_net_19739;
	wire new_net_8025;
	wire new_net_7408;
	wire new_net_17247;
	wire new_net_8133;
	wire new_net_14301;
	wire new_net_7815;
	wire new_net_7966;
	wire new_net_4950;
	wire new_net_6949;
	wire _1604_;
	wire new_net_2127;
	wire new_net_299;
	wire new_net_3274;
	wire new_net_21477;
	wire new_net_11666;
	wire new_net_13177;
	wire new_net_11751;
	wire _1605_;
	wire _1395_;
	wire new_net_819;
	wire new_net_3585;
	wire new_net_15967;
	wire new_net_21274;
	wire new_net_14381;
	wire new_net_16946;
	wire new_net_17786;
	wire new_net_18896;
	wire new_net_11097;
	wire new_net_11307;
	wire new_net_10814;
	wire new_net_7969;
	wire new_net_1831;
	wire new_net_3932;
	wire new_net_6950;
	wire new_net_9893;
	wire new_net_18504;
	wire new_net_18611;
	wire new_net_17895;
	wire _1396_;
	wire new_net_674;
	wire _1606_;
	wire new_net_19337;
	wire new_net_13837;
	wire new_net_18665;
	wire new_net_19195;
	wire new_net_12185;
	wire new_net_15036;
	wire new_net_15934;
	wire new_net_17542;
	wire new_net_14299;
	wire new_net_16430;
	wire new_net_17518;
	wire new_net_11831;
	wire new_net_5929;
	wire new_net_12020;
	wire new_net_13238;
	wire new_net_9724;
	wire new_net_8523;
	wire _1397_;
	wire new_net_826;
	wire _1607_;
	wire new_net_3586;
	wire new_net_4951;
	wire new_net_18610;
	wire new_net_19738;
	wire new_net_17487;
	wire new_net_16011;
	wire new_net_17441;
	wire new_net_14300;
	wire new_net_6512;
	wire new_net_7433;
	wire new_net_2521;
	wire new_net_8024;
	wire new_net_17994;
	wire new_net_8793;
	wire new_net_16717;
	wire new_net_9730;
	wire _1398_;
	wire new_net_298;
	wire new_net_1385;
	wire _1608_;
	wire new_net_6952;
	wire new_net_14517;
	wire new_net_16671;
	wire new_net_304;
	wire new_net_673;
	wire new_net_6957;
	wire new_net_19336;
	wire new_net_21275;
	wire new_net_18372;
	wire new_net_12755;
	wire new_net_9891;
	wire new_net_10815;
	wire new_net_11098;
	wire _1399_;
	wire new_net_821;
	wire _1609_;
	wire new_net_1387;
	wire new_net_11256;
	wire new_net_14449;
	wire new_net_7764;
	wire _1071_;
	wire new_net_2003;
	wire new_net_12449;
	wire new_net_19732;
	wire _0994_;
	wire new_net_18667;
	wire new_net_17653;
	wire new_net_10083;
	wire new_net_839;
	wire new_net_3531;
	wire new_net_20619;
	wire new_net_5716;
	wire new_net_20307;
	wire new_net_16905;
	wire new_net_15391;
	wire new_net_17660;
	wire new_net_14192;
	wire new_net_13039;
	wire new_net_16030;
	wire new_net_16313;
	wire new_net_13663;
	wire new_net_8479;
	wire new_net_12754;
	wire _1274_;
	wire new_net_16849;
	wire new_net_9260;
	wire new_net_1337;
	wire new_net_2763;
	wire new_net_2105;
	wire new_net_4812;
	wire new_net_6350;
	wire new_net_9898;
	wire new_net_18042;
	wire new_net_20232;
	wire new_net_11932;
	wire new_net_14138;
	wire new_net_17971;
	wire new_net_18856;
	wire new_net_5335;
	wire new_net_8436;
	wire new_net_10084;
	wire _1275_;
	wire new_net_17992;
	wire new_net_12105;
	wire new_net_14523;
	wire new_net_12785;
	wire new_net_10272;
	wire new_net_10654;
	wire new_net_9475;
	wire new_net_6809;
	wire new_net_21419;
	wire new_net_12691;
	wire new_net_11914;
	wire new_net_8481;
	wire new_net_1563;
	wire new_net_2767;
	wire _1276_;
	wire new_net_20112;
	wire new_net_20975;
	wire new_net_17074;
	wire new_net_12836;
	wire new_net_307;
	wire new_net_12991;
	wire new_net_14836;
	wire new_net_15662;
	wire new_net_11377;
	wire new_net_10898;
	wire new_net_8482;
	wire new_net_1571;
	wire new_net_2005;
	wire new_net_5558;
	wire new_net_12433;
	wire new_net_1838;
	wire new_net_15168;
	wire new_net_17414;
	wire new_net_18686;
	wire new_net_15347;
	wire new_net_6580;
	wire _1277_;
	wire new_net_2103;
	wire new_net_20620;
	wire new_net_15360;
	wire new_net_17448;
	wire new_net_12431;
	wire new_net_15392;
	wire new_net_8264;
	wire new_net_14193;
	wire new_net_13040;
	wire new_net_15084;
	wire new_net_16314;
	wire new_net_9541;
	wire new_net_8882;
	wire new_net_8543;
	wire new_net_14334;
	wire new_net_16090;
	wire new_net_10520;
	wire new_net_14039;
	wire new_net_14743;
	wire new_net_9709;
	wire new_net_9258;
	wire new_net_8476;
	wire _1278_;
	wire new_net_844;
	wire new_net_20233;
	wire new_net_7492;
	wire new_net_16434;
	wire new_net_15998;
	wire new_net_6808;
	wire new_net_8547;
	wire new_net_8442;
	wire new_net_9263;
	wire new_net_19684;
	wire new_net_19502;
	wire new_net_20886;
	wire new_net_13557;
	wire new_net_14590;
	wire new_net_18878;
	wire new_net_9540;
	wire new_net_10280;
	wire _1279_;
	wire new_net_14503;
	wire new_net_21420;
	wire new_net_11913;
	wire new_net_4463;
	wire new_net_6802;
	wire new_net_19686;
	wire new_net_20113;
	wire new_net_20976;
	wire new_net_3154;
	wire new_net_11624;
	wire new_net_10400;
	wire new_net_11484;
	wire new_net_11378;
	wire new_net_10656;
	wire new_net_10899;
	wire new_net_10087;
	wire _1280_;
	wire new_net_2113;
	wire new_net_2581;
	wire new_net_15211;
	wire new_net_17721;
	wire new_net_5619;
	wire new_net_21051;
	wire new_net_10663;
	wire new_net_10086;
	wire new_net_3570;
	wire new_net_4814;
	wire new_net_5604;
	wire new_net_8090;
	wire new_net_9803;
	wire new_net_20621;
	wire new_net_17710;
	wire new_net_15511;
	wire new_net_13817;
	wire new_net_15085;
	wire new_net_15393;
	wire new_net_17662;
	wire new_net_14194;
	wire new_net_5330;
	wire new_net_13041;
	wire new_net_16032;
	wire new_net_16315;
	wire new_net_13665;
	wire new_net_15927;
	wire new_net_18210;
	wire new_net_17528;
	wire new_net_10736;
	wire new_net_12481;
	wire new_net_14169;
	wire new_net_14038;
	wire new_net_6574;
	wire new_net_10277;
	wire new_net_8548;
	wire new_net_8440;
	wire new_net_1567;
	wire new_net_2765;
	wire new_net_4210;
	wire new_net_4326;
	wire new_net_4462;
	wire new_net_19659;
	wire new_net_21159;
	wire new_net_4484;
	wire new_net_12998;
	wire new_net_2490;
	wire new_net_10281;
	wire new_net_4464;
	wire new_net_8618;
	wire new_net_3293;
	wire _1282_;
	wire new_net_13627;
	wire new_net_4205;
	wire new_net_17941;
	wire new_net_9538;
	wire new_net_10274;
	wire new_net_4327;
	wire new_net_5653;
	wire new_net_21421;
	wire new_net_17862;
	wire new_net_13467;
	wire new_net_21375;
	wire new_net_13743;
	wire new_net_11912;
	wire new_net_8721;
	wire new_net_9894;
	wire _1463_;
	wire _1283_;
	wire new_net_1368;
	wire new_net_18412;
	wire new_net_20114;
	wire new_net_20977;
	wire new_net_17035;
	wire new_net_11485;
	wire new_net_10900;
	wire new_net_11379;
	wire new_net_3452;
	wire new_net_5556;
	wire new_net_12158;
	wire new_net_19692;
	wire new_net_12382;
	wire new_net_12928;
	wire new_net_21299;
	wire new_net_841;
	wire new_net_5428;
	wire new_net_5651;
	wire new_net_1569;
	wire new_net_8085;
	wire new_net_1336;
	wire new_net_8614;
	wire new_net_10080;
	wire _1284_;
	wire new_net_2108;
	wire new_net_17706;
	wire new_net_15462;
	wire new_net_17146;
	wire new_net_13818;
	wire new_net_15086;
	wire new_net_15394;
	wire new_net_13666;
	wire new_net_12757;
	wire new_net_17663;
	wire new_net_12429;
	wire new_net_13042;
	wire new_net_16033;
	wire new_net_16316;
	wire new_net_14741;
	wire new_net_5649;
	wire new_net_14037;
	wire new_net_1570;
	wire new_net_5597;
	wire new_net_6354;
	wire _1285_;
	wire new_net_2009;
	wire new_net_4209;
	wire new_net_19317;
	wire new_net_14201;
	wire new_net_16324;
	wire new_net_14167;
	wire new_net_10519;
	wire new_net_9542;
	wire new_net_6355;
	wire new_net_9261;
	wire new_net_13628;
	wire new_net_19124;
	wire new_net_11665;
	wire new_net_14598;
	wire new_net_13178;
	wire new_net_9013;
	wire new_net_11752;
	wire new_net_5654;
	wire new_net_4810;
	wire _1286_;
	wire new_net_1340;
	wire new_net_9477;
	wire new_net_21422;
	wire new_net_8411;
	wire new_net_14382;
	wire new_net_16947;
	wire new_net_17787;
	wire new_net_18897;
	wire new_net_18505;
	wire new_net_4207;
	wire new_net_8266;
	wire new_net_10271;
	wire new_net_4881;
	wire new_net_6346;
	wire new_net_11911;
	wire new_net_9259;
	wire new_net_1338;
	wire new_net_1378;
	wire new_net_2112;
	wire new_net_7812;
	wire new_net_17896;
	wire new_net_5550;
	wire new_net_11486;
	wire new_net_11380;
	wire new_net_10275;
	wire new_net_10901;
	wire _1287_;
	wire new_net_838;
	wire new_net_13838;
	wire new_net_18666;
	wire new_net_19196;
	wire new_net_2013;
	wire new_net_9470;
	wire new_net_19116;
	wire new_net_12143;
	wire new_net_12428;
	wire new_net_15087;
	wire new_net_13819;
	wire new_net_15395;
	wire new_net_14196;
	wire new_net_13667;
	wire new_net_5600;
	wire new_net_13043;
	wire new_net_17664;
	wire new_net_17488;
	wire new_net_16012;
	wire new_net_17442;
	wire new_net_10082;
	wire new_net_8722;
	wire new_net_14740;
	wire new_net_10522;
	wire new_net_14036;
	wire new_net_10658;
	wire new_net_8083;
	wire new_net_2759;
	wire new_net_4208;
	wire new_net_6345;
	wire new_net_17995;
	wire new_net_16718;
	wire _1289_;
	wire new_net_13629;
	wire new_net_5332;
	wire new_net_8267;
	wire new_net_4883;
	wire new_net_2758;
	wire new_net_14518;
	wire new_net_13262;
	wire new_net_16672;
	wire new_net_16584;
	wire new_net_8880;
	wire new_net_6584;
	wire new_net_9473;
	wire new_net_1370;
	wire new_net_2111;
	wire new_net_4460;
	wire new_net_8439;
	wire new_net_19123;
	wire new_net_19685;
	wire new_net_21423;
	wire new_net_18373;
	wire new_net_12756;
	wire new_net_5841;
	wire new_net_848;
	wire new_net_8086;
	wire new_net_6578;
	wire new_net_8621;
	wire new_net_9704;
	wire new_net_9539;
	wire new_net_11910;
	wire new_net_5331;
	wire new_net_2106;
	wire _1290_;
	wire new_net_3838;
	wire new_net_12450;
	wire new_net_16317;
	wire new_net_11487;
	wire new_net_11381;
	wire new_net_10902;
	wire new_net_4880;
	wire new_net_5652;
	wire new_net_9257;
	wire new_net_18726;
	wire new_net_9675;
	wire new_net_7612;
	wire new_net_6577;
	wire new_net_4325;
	wire _1291_;
	wire new_net_17654;
	wire new_net_18668;
	wire new_net_3333;
	wire new_net_13820;
	wire new_net_12144;
	wire new_net_12427;
	wire new_net_9895;
	wire new_net_15088;
	wire new_net_15396;
	wire new_net_17665;
	wire new_net_14197;
	wire new_net_13044;
	wire new_net_16035;
	wire new_net_7074;
	wire new_net_16850;
	wire new_net_14035;
	wire new_net_14739;
	wire _1292_;
	wire new_net_1334;
	wire new_net_20237;
	wire new_net_21406;
	wire new_net_18041;
	wire new_net_883;
	wire new_net_11933;
	wire new_net_14139;
	wire new_net_17970;
	wire new_net_8723;
	wire new_net_10662;
	wire new_net_8620;
	wire new_net_8877;
	wire new_net_4808;
	wire new_net_9267;
	wire new_net_13630;
	wire new_net_18857;
	wire new_net_12106;
	wire new_net_14524;
	wire new_net_12786;
	wire new_net_4324;
	wire new_net_6349;
	wire _1293_;
	wire new_net_1371;
	wire new_net_9266;
	wire new_net_21424;
	wire new_net_7741;
	wire new_net_12692;
	wire new_net_13483;
	wire new_net_9899;
	wire new_net_10399;
	wire new_net_8624;
	wire new_net_11909;
	wire new_net_1561;
	wire new_net_2762;
	wire new_net_3528;
	wire new_net_3569;
	wire new_net_19122;
	wire new_net_20117;
	wire new_net_17075;
	wire new_net_12837;
	wire new_net_11488;
	wire new_net_11382;
	wire new_net_4328;
	wire new_net_5323;
	wire new_net_10903;
	wire _1294_;
	wire new_net_5336;
	wire new_net_6461;
	wire new_net_2107;
	wire new_net_19691;
	wire new_net_20749;
	wire new_net_15169;
	wire new_net_17415;
	wire new_net_18687;
	wire new_net_15348;
	wire new_net_1346;
	wire new_net_9544;
	wire new_net_1373;
	wire new_net_4885;
	wire new_net_8542;
	wire new_net_15013;
	wire new_net_7421;
	wire new_net_15361;
	wire new_net_4212;
	wire new_net_13669;
	wire new_net_12760;
	wire new_net_16036;
	wire new_net_13821;
	wire new_net_15089;
	wire new_net_6805;
	wire new_net_12145;
	wire new_net_12426;
	wire new_net_15397;
	wire new_net_5213;
	wire new_net_14335;
	wire new_net_7130;
	wire new_net_14034;
	wire new_net_14738;
	wire new_net_10398;
	wire new_net_2011;
	wire new_net_3571;
	wire new_net_6351;
	wire new_net_16091;
	wire new_net_20238;
	wire new_net_16435;
	wire new_net_13631;
	wire new_net_4811;
	wire new_net_5551;
	wire new_net_10273;
	wire new_net_10660;
	wire _1296_;
	wire new_net_18017;
	wire new_net_21081;
	wire new_net_15999;
	wire new_net_10455;
	wire new_net_14591;
	wire new_net_6803;
	wire new_net_4467;
	wire new_net_5337;
	wire new_net_5427;
	wire new_net_5598;
	wire new_net_21425;
	wire new_net_14504;
	wire new_net_8483;
	wire new_net_6348;
	wire new_net_11908;
	wire _1297_;
	wire new_net_1379;
	wire new_net_8444;
	wire new_net_20118;
	wire new_net_20625;
	wire new_net_20981;
	wire new_net_1923;
	wire new_net_12432;
	wire new_net_11625;
	wire new_net_6575;
	wire new_net_11489;
	wire new_net_11383;
	wire new_net_8552;
	wire new_net_10904;
	wire new_net_1375;
	wire new_net_19121;
	wire new_net_19690;
	wire new_net_14686;
	wire new_net_19318;
	wire new_net_15212;
	wire new_net_17722;
	wire new_net_21052;
	wire new_net_4211;
	wire new_net_8084;
	wire new_net_8724;
	wire new_net_4809;
	wire new_net_6576;
	wire new_net_10657;
	wire _1298_;
	wire new_net_9262;
	wire new_net_15512;
	wire new_net_17711;
	wire new_net_18178;
	wire new_net_8478;
	wire new_net_12761;
	wire new_net_12146;
	wire new_net_12425;
	wire new_net_8091;
	wire new_net_13822;
	wire new_net_15090;
	wire new_net_15398;
	wire new_net_17667;
	wire new_net_14199;
	wire new_net_15928;
	wire new_net_18211;
	wire new_net_14261;
	wire new_net_17529;
	wire new_net_12482;
	wire new_net_9897;
	wire new_net_14033;
	wire new_net_14737;
	wire new_net_5552;
	wire new_net_10396;
	wire new_net_9708;
	wire new_net_9546;
	wire new_net_4466;
	wire new_net_5599;
	wire new_net_6347;
	wire new_net_17506;
	wire new_net_19660;
	wire new_net_21160;
	wire new_net_13632;
	wire new_net_1377;
	wire new_net_5603;
	wire new_net_19115;
	wire new_net_12999;
	wire new_net_17942;
	wire new_net_19866;
	wire new_net_3566;
	wire new_net_8082;
	wire new_net_6804;
	wire new_net_9707;
	wire _1300_;
	wire new_net_1568;
	wire new_net_2008;
	wire new_net_21426;
	wire new_net_17863;
	wire new_net_13468;
	wire new_net_9901;
	wire new_net_8088;
	wire new_net_11907;
	wire new_net_20119;
	wire new_net_20626;
	wire new_net_20982;
	wire new_net_18413;
	wire new_net_17036;
	wire _0588_;
	wire new_net_9468;
	wire new_net_5655;
	wire new_net_8092;
	wire new_net_6806;
	wire new_net_11490;
	wire new_net_11384;
	wire new_net_10278;
	wire _1301_;
	wire new_net_2109;
	wire new_net_4459;
	wire new_net_12157;
	wire new_net_12383;
	wire new_net_12929;
	wire new_net_8089;
	wire new_net_10397;
	wire new_net_1565;
	wire new_net_19120;
	wire new_net_17707;
	wire new_net_15463;
	wire new_net_17147;
	wire new_net_12762;
	wire new_net_4214;
	wire new_net_12147;
	wire new_net_12424;
	wire new_net_13823;
	wire new_net_15091;
	wire new_net_15399;
	wire new_net_17668;
	wire new_net_14200;
	wire _1302_;
	wire new_net_14032;
	wire new_net_9710;
	wire new_net_10276;
	wire new_net_3527;
	wire new_net_8549;
	wire new_net_8878;
	wire new_net_19682;
	wire new_net_20240;
	wire new_net_14202;
	wire new_net_3772;
	wire new_net_13633;
	wire new_net_4206;
	wire _1303_;
	wire new_net_8616;
	wire new_net_3793;
	wire new_net_9940;
	wire new_net_14168;
	wire new_net_11664;
	wire new_net_5495;
	wire new_net_14599;
	wire new_net_14736;
	wire new_net_8265;
	wire new_net_9712;
	wire new_net_843;
	wire new_net_3568;
	wire new_net_4461;
	wire new_net_11753;
	wire new_net_21427;
	wire new_net_8405;
	wire new_net_14383;
	wire new_net_16948;
	wire new_net_17788;
	wire new_net_18898;
	wire new_net_9472;
	wire new_net_6579;
	wire new_net_9545;
	wire _1304_;
	wire new_net_1335;
	wire new_net_11906;
	wire new_net_20120;
	wire new_net_20627;
	wire new_net_20983;
	wire new_net_18506;
	wire new_net_14683;
	wire new_net_17897;
	wire new_net_11491;
	wire new_net_11385;
	wire new_net_846;
	wire new_net_8441;
	wire new_net_10906;
	wire new_net_17336;
	wire new_net_18448;
	wire _1305_;
	wire new_net_4330;
	wire new_net_10905;
	wire new_net_15533;
	wire new_net_13672;
	wire new_net_12763;
	wire new_net_13638;
	wire new_net_12148;
	wire new_net_12423;
	wire new_net_10523;
	wire new_net_13824;
	wire new_net_15092;
	wire new_net_15400;
	wire new_net_17669;
	wire new_net_20482;
	wire new_net_17638;
	wire new_net_17489;
	wire new_net_17443;
	wire new_net_16013;
	wire new_net_10077;
	wire new_net_9474;
	wire new_net_5650;
	wire new_net_14031;
	wire new_net_2006;
	wire _1306_;
	wire new_net_845;
	wire new_net_6352;
	wire new_net_8546;
	wire new_net_20241;
	wire new_net_17996;
	wire new_net_19348;
	wire new_net_16719;
	wire new_net_13634;
	wire new_net_2010;
	wire new_net_5327;
	wire new_net_14519;
	wire new_net_13263;
	wire new_net_9896;
	wire new_net_2014;
	wire _1307_;
	wire new_net_1372;
	wire new_net_2110;
	wire new_net_5326;
	wire new_net_21428;
	wire new_net_16585;
	wire new_net_18374;
	wire new_net_9705;
	wire new_net_2764;
	wire new_net_8550;
	wire new_net_8619;
	wire new_net_11905;
	wire new_net_20121;
	wire new_net_20628;
	wire new_net_20984;
	wire new_net_4807;
	wire new_net_11492;
	wire new_net_11386;
	wire _1308_;
	wire new_net_4465;
	wire new_net_4879;
	wire new_net_8544;
	wire new_net_10907;
	wire new_net_12451;
	wire new_net_18727;
	wire new_net_12962;
	wire _1001_;
	wire new_net_8087;
	wire new_net_3526;
	wire new_net_3574;
	wire new_net_18669;
	wire new_net_17655;
	wire new_net_19501;
	wire new_net_6554;
	wire new_net_13673;
	wire new_net_12764;
	wire new_net_13637;
	wire new_net_12149;
	wire new_net_12422;
	wire new_net_13825;
	wire new_net_15093;
	wire new_net_6582;
	wire new_net_15401;
	wire new_net_17670;
	wire new_net_16907;
	wire new_net_16851;
	wire new_net_10521;
	wire new_net_14030;
	wire new_net_14735;
	wire new_net_840;
	wire new_net_1339;
	wire new_net_6583;
	wire new_net_6807;
	wire new_net_19118;
	wire new_net_20242;
	wire new_net_14140;
	wire new_net_11934;
	wire new_net_13635;
	wire _1310_;
	wire new_net_18858;
	wire new_net_12107;
	wire new_net_7121;
	wire new_net_8475;
	wire new_net_9706;
	wire new_net_4813;
	wire new_net_6462;
	wire new_net_14525;
	wire new_net_8875;
	wire new_net_19688;
	wire new_net_21429;
	wire new_net_12693;
	wire _1311_;
	wire new_net_5553;
	wire new_net_1374;
	wire new_net_5602;
	wire new_net_11904;
	wire new_net_20122;
	wire new_net_20629;
	wire new_net_20985;
	wire new_net_13484;
	wire new_net_17076;
	wire new_net_8438;
	wire new_net_9265;
	wire new_net_9467;
	wire new_net_11493;
	wire new_net_11387;
	wire new_net_6581;
	wire new_net_10661;
	wire new_net_10908;
	wire new_net_17799;
	wire new_net_19689;
	wire new_net_15170;
	wire new_net_17416;
	wire new_net_18688;
	wire new_net_18950;
	wire _1312_;
	wire new_net_3794;
	wire new_net_5329;
	wire new_net_10655;
	wire new_net_15349;
	wire new_net_18647;
	wire new_net_15362;
	wire new_net_8545;
	wire new_net_8615;
	wire new_net_13050;
	wire new_net_16041;
	wire new_net_16323;
	wire new_net_13674;
	wire new_net_9469;
	wire new_net_12765;
	wire new_net_12150;
	wire new_net_8081;
	wire new_net_17450;
	wire new_net_14336;
	wire new_net_9900;
	wire new_net_14029;
	wire new_net_14734;
	wire _1313_;
	wire new_net_1562;
	wire new_net_19683;
	wire new_net_20243;
	wire new_net_16092;
	wire new_net_17547;
	wire new_net_21117;
	wire new_net_16436;
	wire new_net_13636;
	wire new_net_1566;
	wire new_net_9537;
	wire new_net_10078;
	wire new_net_10659;
	wire new_net_19117;
	wire new_net_18018;
	wire new_net_21082;
	wire new_net_16000;
	wire new_net_16302;
	wire new_net_5601;
	wire new_net_8883;
	wire new_net_6460;
	wire new_net_10085;
	wire _1314_;
	wire new_net_2760;
	wire new_net_21430;
	wire new_net_14505;
	wire new_net_8881;
	wire new_net_11903;
	wire new_net_10081;
	wire new_net_9471;
	wire new_net_1564;
	wire new_net_2012;
	wire new_net_2766;
	wire new_net_5555;
	wire new_net_20123;
	wire new_net_20630;
	wire new_net_15710;
	wire new_net_4882;
	wire new_net_8551;
	wire new_net_10909;
	wire new_net_14028;
	wire new_net_14733;
	wire new_net_5557;
	wire new_net_6810;
	wire new_net_11494;
	wire new_net_11388;
	wire _1315_;
	wire new_net_11626;
	wire new_net_14687;
	wire new_net_17723;
	wire new_net_21053;
	wire new_net_15513;
	wire new_net_17712;
	wire new_net_7510;
	wire new_net_10282;
	wire new_net_6963;
	wire new_net_15929;
	wire new_net_18212;
	wire new_net_14262;
	wire new_net_17530;
	wire new_net_12483;
	wire new_net_14171;
	wire new_net_16384;
	wire new_net_13333;
	wire new_net_14673;
	wire new_net_14768;
	wire new_net_17791;
	wire new_net_3958;
	wire new_net_15072;
	wire new_net_15237;
	wire new_net_6276;
	wire new_net_15368;
	wire new_net_19661;
	wire new_net_21161;
	wire new_net_9822;
	wire new_net_9024;
	wire new_net_20256;
	wire new_net_2495;
	wire new_net_13000;
	wire new_net_17943;
	wire new_net_11976;
	wire new_net_7138;
	wire new_net_2031;
	wire new_net_10286;
	wire new_net_10765;
	wire new_net_5270;
	wire new_net_1053;
	wire new_net_1543;
	wire new_net_4050;
	wire new_net_21224;
	wire new_net_17864;
	wire new_net_13469;
	wire new_net_21374;
	wire new_net_6209;
	wire new_net_3635;
	wire new_net_4203;
	wire new_net_6964;
	wire new_net_13744;
	wire _1470_;
	wire new_net_18414;
	wire new_net_17037;
	wire new_net_14108;
	wire new_net_1748;
	wire new_net_6774;
	wire new_net_2036;
	wire new_net_10289;
	wire new_net_8700;
	wire new_net_2530;
	wire new_net_6438;
	wire new_net_20667;
	wire new_net_12156;
	wire new_net_18633;
	wire new_net_12384;
	wire new_net_12361;
	wire new_net_11004;
	wire new_net_9816;
	wire new_net_11543;
	wire new_net_10755;
	wire new_net_3634;
	wire new_net_509;
	wire new_net_1535;
	wire new_net_2026;
	wire new_net_19563;
	wire new_net_20883;
	wire new_net_15464;
	wire new_net_5231;
	wire new_net_17148;
	wire new_net_10285;
	wire new_net_7185;
	wire new_net_5269;
	wire new_net_4972;
	wire new_net_1538;
	wire new_net_14087;
	wire new_net_16409;
	wire new_net_16385;
	wire new_net_10166;
	wire new_net_13334;
	wire new_net_14674;
	wire new_net_14769;
	wire new_net_17792;
	wire new_net_15073;
	wire new_net_15238;
	wire new_net_10664;
	wire new_net_14203;
	wire new_net_16326;
	wire new_net_5822;
	wire new_net_5725;
	wire new_net_6274;
	wire new_net_4976;
	wire new_net_3637;
	wire new_net_20257;
	wire new_net_11663;
	wire new_net_14600;
	wire new_net_11754;
	wire new_net_8702;
	wire new_net_10764;
	wire new_net_1311;
	wire new_net_14384;
	wire new_net_16949;
	wire new_net_17789;
	wire new_net_18899;
	wire new_net_4048;
	wire new_net_6959;
	wire new_net_18507;
	wire new_net_14684;
	wire new_net_510;
	wire new_net_3638;
	wire new_net_20668;
	wire new_net_20752;
	wire new_net_21404;
	wire new_net_17337;
	wire new_net_6439;
	wire new_net_11005;
	wire new_net_14107;
	wire new_net_6776;
	wire new_net_11544;
	wire new_net_10305;
	wire new_net_1055;
	wire new_net_10828;
	wire new_net_19564;
	wire new_net_20884;
	wire new_net_15534;
	wire new_net_7141;
	wire new_net_5821;
	wire new_net_3656;
	wire new_net_4046;
	wire new_net_4202;
	wire new_net_5720;
	wire new_net_17490;
	wire new_net_4003;
	wire new_net_5624;
	wire new_net_16014;
	wire new_net_17444;
	wire new_net_14088;
	wire new_net_16410;
	wire new_net_16386;
	wire new_net_13335;
	wire new_net_14675;
	wire new_net_10290;
	wire new_net_14770;
	wire new_net_17793;
	wire new_net_7183;
	wire new_net_15074;
	wire new_net_7611;
	wire new_net_17997;
	wire new_net_6823;
	wire new_net_16720;
	wire new_net_19452;
	wire new_net_10163;
	wire new_net_4197;
	wire new_net_1542;
	wire new_net_3658;
	wire new_net_6210;
	wire new_net_20258;
	wire new_net_13252;
	wire new_net_16697;
	wire new_net_10331;
	wire new_net_14520;
	wire new_net_20820;
	wire new_net_13264;
	wire new_net_16674;
	wire new_net_6965;
	wire new_net_5433;
	wire new_net_6770;
	wire new_net_2529;
	wire new_net_18375;
	wire new_net_11473;
	wire new_net_12758;
	wire new_net_500;
	wire new_net_5717;
	wire new_net_6212;
	wire new_net_1996;
	wire new_net_6968;
	wire new_net_7758;
	wire new_net_10287;
	wire new_net_5714;
	wire new_net_501;
	wire new_net_12452;
	wire new_net_20669;
	wire new_net_20753;
	wire new_net_18728;
	wire new_net_21309;
	wire new_net_12963;
	wire new_net_11006;
	wire new_net_14106;
	wire new_net_11545;
	wire new_net_8703;
	wire new_net_10303;
	wire new_net_5723;
	wire new_net_6269;
	wire new_net_6216;
	wire new_net_17656;
	wire new_net_10829;
	wire new_net_18670;
	wire new_net_2622;
	wire new_net_7512;
	wire new_net_10307;
	wire new_net_6211;
	wire new_net_15308;
	wire new_net_19694;
	wire new_net_16908;
	wire new_net_18136;
	wire new_net_19246;
	wire new_net_7067;
	wire new_net_16852;
	wire new_net_14089;
	wire new_net_16411;
	wire new_net_16387;
	wire new_net_10167;
	wire new_net_13336;
	wire new_net_14676;
	wire new_net_14771;
	wire new_net_17794;
	wire new_net_15075;
	wire new_net_15240;
	wire new_net_7143;
	wire new_net_11935;
	wire new_net_14141;
	wire new_net_10304;
	wire new_net_10756;
	wire new_net_499;
	wire new_net_10431;
	wire new_net_20259;
	wire new_net_9274;
	wire new_net_18859;
	wire new_net_18291;
	wire new_net_12108;
	wire new_net_14526;
	wire new_net_12788;
	wire new_net_9031;
	wire new_net_7513;
	wire new_net_10763;
	wire new_net_3441;
	wire new_net_1054;
	wire new_net_3633;
	wire new_net_9677;
	wire new_net_11969;
	wire new_net_12694;
	wire new_net_11330;
	wire new_net_5057;
	wire new_net_10436;
	wire new_net_5824;
	wire new_net_17184;
	wire new_net_17077;
	wire new_net_6775;
	wire new_net_8697;
	wire new_net_10754;
	wire new_net_5054;
	wire new_net_5715;
	wire new_net_20670;
	wire new_net_20754;
	wire new_net_15171;
	wire new_net_17417;
	wire new_net_20411;
	wire new_net_18689;
	wire new_net_6219;
	wire new_net_10830;
	wire new_net_4051;
	wire new_net_11007;
	wire new_net_15350;
	wire new_net_11546;
	wire new_net_4198;
	wire new_net_7181;
	wire new_net_1313;
	wire new_net_2531;
	wire new_net_18646;
	wire new_net_15015;
	wire new_net_15363;
	wire new_net_6275;
	wire new_net_17451;
	wire new_net_14337;
	wire new_net_16412;
	wire new_net_14105;
	wire new_net_16388;
	wire new_net_13337;
	wire new_net_14677;
	wire new_net_14772;
	wire new_net_17795;
	wire new_net_15076;
	wire new_net_15241;
	wire new_net_6143;
	wire _0140_;
	wire new_net_16093;
	wire new_net_21118;
	wire new_net_16437;
	wire new_net_4975;
	wire new_net_9025;
	wire new_net_8701;
	wire new_net_502;
	wire new_net_1532;
	wire new_net_20260;
	wire new_net_18019;
	wire new_net_21083;
	wire new_net_16001;
	wire new_net_1743;
	wire new_net_14506;
	wire new_net_6333;
	wire new_net_6960;
	wire new_net_7755;
	wire new_net_7514;
	wire new_net_15711;
	wire new_net_12430;
	wire new_net_11627;
	wire new_net_4973;
	wire new_net_10161;
	wire new_net_1303;
	wire new_net_1537;
	wire new_net_20671;
	wire new_net_20755;
	wire new_net_14688;
	wire new_net_17724;
	wire new_net_10429;
	wire new_net_10831;
	wire new_net_14090;
	wire new_net_11008;
	wire new_net_4199;
	wire new_net_5460;
	wire new_net_8704;
	wire new_net_19567;
	wire new_net_20887;
	wire new_net_21054;
	wire new_net_7548;
	wire new_net_15514;
	wire new_net_17713;
	wire new_net_7142;
	wire new_net_7759;
	wire new_net_1305;
	wire new_net_15930;
	wire new_net_18213;
	wire new_net_16413;
	wire new_net_9029;
	wire new_net_14104;
	wire new_net_16389;
	wire new_net_7753;
	wire new_net_13338;
	wire new_net_14678;
	wire new_net_14773;
	wire new_net_17796;
	wire new_net_10757;
	wire new_net_12484;
	wire new_net_19662;
	wire new_net_21162;
	wire new_net_14103;
	wire new_net_1051;
	wire new_net_5273;
	wire new_net_20261;
	wire new_net_9572;
	wire new_net_13001;
	wire new_net_17944;
	wire new_net_6768;
	wire new_net_10762;
	wire new_net_3813;
	wire new_net_5058;
	wire new_net_11977;
	wire new_net_9917;
	wire new_net_17865;
	wire new_net_13470;
	wire new_net_15669;
	wire new_net_10283;
	wire new_net_5724;
	wire new_net_18415;
	wire new_net_17038;
	wire _0595_;
	wire new_net_10291;
	wire new_net_10309;
	wire new_net_2035;
	wire new_net_1540;
	wire new_net_5056;
	wire new_net_5434;
	wire new_net_6213;
	wire new_net_20672;
	wire new_net_20756;
	wire new_net_12155;
	wire new_net_12385;
	wire new_net_12931;
	wire new_net_5272;
	wire new_net_11009;
	wire new_net_10832;
	wire new_net_6771;
	wire new_net_1306;
	wire new_net_19568;
	wire new_net_20888;
	wire new_net_10435;
	wire new_net_6772;
	wire new_net_7184;
	wire new_net_17149;
	wire new_net_1042;
	wire new_net_5465;
	wire new_net_5036;
	wire new_net_5274;
	wire new_net_15374;
	wire new_net_15905;
	wire new_net_14091;
	wire new_net_16414;
	wire new_net_16390;
	wire new_net_13339;
	wire new_net_14679;
	wire new_net_14774;
	wire new_net_17797;
	wire new_net_6268;
	wire new_net_9022;
	wire new_net_7756;
	wire new_net_7515;
	wire new_net_7186;
	wire new_net_1747;
	wire new_net_6217;
	wire new_net_20262;
	wire new_net_11587;
	wire new_net_11662;
	wire new_net_14601;
	wire new_net_10430;
	wire new_net_11547;
	wire new_net_5934;
	wire new_net_11755;
	wire new_net_14385;
	wire new_net_16950;
	wire new_net_17790;
	wire new_net_18900;
	wire new_net_11548;
	wire new_net_3814;
	wire new_net_18508;
	wire new_net_7007;
	wire new_net_6961;
	wire new_net_10758;
	wire new_net_1533;
	wire new_net_507;
	wire new_net_3655;
	wire new_net_20673;
	wire new_net_20757;
	wire new_net_17338;
	wire new_net_10833;
	wire new_net_11010;
	wire new_net_14102;
	wire new_net_5819;
	wire new_net_1746;
	wire new_net_2027;
	wire new_net_1308;
	wire new_net_19569;
	wire new_net_20889;
	wire new_net_15535;
	wire new_net_6214;
	wire new_net_9817;
	wire new_net_4201;
	wire new_net_8698;
	wire new_net_1534;
	wire new_net_1737;
	wire new_net_1312;
	wire new_net_17640;
	wire new_net_17491;
	wire new_net_15375;
	wire new_net_15906;
	wire new_net_14092;
	wire new_net_16415;
	wire new_net_16391;
	wire new_net_13340;
	wire new_net_14680;
	wire new_net_14775;
	wire new_net_17798;
	wire new_net_15244;
	wire new_net_9015;
	wire new_net_14086;
	wire new_net_17998;
	wire new_net_18473;
	wire new_net_14605;
	wire new_net_6277;
	wire new_net_10432;
	wire new_net_10306;
	wire new_net_8705;
	wire new_net_16721;
	wire new_net_5466;
	wire new_net_1307;
	wire new_net_20263;
	wire new_net_13253;
	wire new_net_16698;
	wire new_net_9819;
	wire new_net_10761;
	wire new_net_4196;
	wire new_net_5820;
	wire new_net_16675;
	wire new_net_11474;
	wire new_net_5060;
	wire new_net_10165;
	wire new_net_3653;
	wire new_net_4043;
	wire new_net_12759;
	wire new_net_5838;
	wire new_net_6773;
	wire new_net_2527;
	wire new_net_508;
	wire new_net_5275;
	wire new_net_6215;
	wire new_net_20674;
	wire new_net_20758;
	wire new_net_12453;
	wire new_net_18729;
	wire new_net_19151;
	wire new_net_12964;
	wire _1008_;
	wire new_net_10834;
	wire new_net_11011;
	wire new_net_14101;
	wire new_net_10160;
	wire new_net_9820;
	wire new_net_15079;
	wire new_net_19570;
	wire new_net_20890;
	wire new_net_18671;
	wire new_net_17657;
	wire new_net_1541;
	wire new_net_6278;
	wire new_net_15309;
	wire new_net_19695;
	wire new_net_16909;
	wire new_net_5718;
	wire new_net_6270;
	wire new_net_15376;
	wire new_net_15907;
	wire new_net_14093;
	wire new_net_16416;
	wire new_net_16392;
	wire new_net_7752;
	wire new_net_13341;
	wire new_net_14681;
	wire new_net_7140;
	wire new_net_20264;
	wire new_net_885;
	wire new_net_11936;
	wire new_net_9160;
	wire new_net_18860;
	wire new_net_8879;
	wire new_net_9821;
	wire new_net_4866;
	wire new_net_12789;
	wire new_net_11970;
	wire new_net_7182;
	wire new_net_6966;
	wire new_net_10759;
	wire new_net_2028;
	wire new_net_504;
	wire new_net_3661;
	wire new_net_5462;
	wire new_net_17078;
	wire new_net_5722;
	wire new_net_3660;
	wire new_net_1046;
	wire new_net_20675;
	wire new_net_20759;
	wire new_net_10739;
	wire new_net_17801;
	wire new_net_15012;
	wire new_net_15172;
	wire new_net_17418;
	wire new_net_18690;
	wire new_net_7187;
	wire new_net_10168;
	wire new_net_10835;
	wire new_net_7760;
	wire new_net_11549;
	wire new_net_11012;
	wire new_net_7139;
	wire new_net_1302;
	wire new_net_1047;
	wire new_net_5459;
	wire new_net_15351;
	wire new_net_15016;
	wire new_net_14570;
	wire new_net_15364;
	wire new_net_6218;
	wire new_net_1043;
	wire new_net_21222;
	wire new_net_17452;
	wire new_net_15080;
	wire new_net_15377;
	wire new_net_15908;
	wire new_net_13342;
	wire new_net_14094;
	wire new_net_16393;
	wire new_net_14100;
	wire new_net_14682;
	wire new_net_15246;
	wire new_net_17800;
	wire new_net_21243;
	wire new_net_16094;
	wire new_net_17549;
	wire new_net_21119;
	wire new_net_16438;
	wire new_net_7188;
	wire new_net_3659;
	wire new_net_10288;
	wire new_net_1049;
	wire new_net_20265;
	wire new_net_18020;
	wire new_net_21084;
	wire new_net_16002;
	wire new_net_19499;
	wire new_net_10760;
	wire new_net_10433;
	wire new_net_10162;
	wire new_net_1742;
	wire new_net_4049;
	wire new_net_6273;
	wire new_net_7761;
	wire new_net_7165;
	wire new_net_13497;
	wire new_net_14507;
	wire new_net_1017;
	wire new_net_6038;
	wire new_net_6267;
	wire new_net_6769;
	wire new_net_7511;
	wire new_net_1052;
	wire new_net_1740;
	wire new_net_15712;
	wire new_net_11389;
	wire new_net_11245;
	wire new_net_1536;
	wire new_net_20676;
	wire new_net_20760;
	wire new_net_11628;
	wire new_net_14689;
	wire new_net_4200;
	wire new_net_6271;
	wire new_net_10836;
	wire new_net_11013;
	wire new_net_6777;
	wire new_net_7754;
	wire new_net_11550;
	wire new_net_505;
	wire new_net_19572;
	wire new_net_17725;
	wire new_net_21055;
	wire new_net_15515;
	wire new_net_17714;
	wire new_net_10312;
	wire new_net_6962;
	wire new_net_9030;
	wire new_net_2983;
	wire new_net_15931;
	wire new_net_18214;
	wire new_net_15081;
	wire new_net_15247;
	wire new_net_15378;
	wire new_net_15909;
	wire new_net_14095;
	wire new_net_16418;
	wire new_net_14099;
	wire new_net_16394;
	wire new_net_6767;
	wire new_net_13343;
	wire new_net_12485;
	wire new_net_14173;
	wire new_net_19291;
	wire new_net_19663;
	wire new_net_21163;
	wire new_net_2532;
	wire new_net_3662;
	wire new_net_5271;
	wire new_net_5721;
	wire new_net_20266;
	wire new_net_13002;
	wire new_net_17945;
	wire new_net_4366;
	wire new_net_5719;
	wire new_net_4047;
	wire new_net_9023;
	wire new_net_3636;
	wire new_net_11978;
	wire new_net_8443;
	wire new_net_17866;
	wire new_net_10164;
	wire new_net_9814;
	wire new_net_1744;
	wire new_net_2033;
	wire new_net_7757;
	wire new_net_9026;
	wire new_net_13471;
	wire new_net_10292;
	wire new_net_5537;
	wire new_net_15190;
	wire new_net_16158;
	wire new_net_13742;
	wire _1477_;
	wire new_net_18416;
	wire new_net_5463;
	wire new_net_10310;
	wire new_net_9818;
	wire new_net_17039;
	wire new_net_1050;
	wire new_net_20677;
	wire new_net_20761;
	wire new_net_12154;
	wire new_net_11551;
	wire new_net_7180;
	wire new_net_10308;
	wire new_net_10837;
	wire new_net_11014;
	wire new_net_1738;
	wire new_net_4044;
	wire new_net_4974;
	wire new_net_5059;
	wire new_net_19573;
	wire new_net_10284;
	wire new_net_8699;
	wire new_net_4045;
	wire new_net_6437;
	wire new_net_14097;
	wire new_net_1745;
	wire new_net_1304;
	wire new_net_15466;
	wire new_net_17150;
	wire new_net_14779;
	wire new_net_17802;
	wire new_net_15082;
	wire new_net_15248;
	wire new_net_15379;
	wire new_net_15910;
	wire new_net_10428;
	wire new_net_6958;
	wire new_net_14096;
	wire new_net_16419;
	wire new_net_7516;
	wire new_net_20267;
	wire new_net_16328;
	wire new_net_21242;
	wire new_net_5982;
	wire new_net_7922;
	wire new_net_14602;
	wire new_net_675;
	wire new_net_11756;
	wire new_net_14386;
	wire new_net_3657;
	wire new_net_7750;
	wire new_net_18509;
	wire new_net_10096;
	wire new_net_10169;
	wire new_net_5276;
	wire new_net_5461;
	wire new_net_9027;
	wire new_net_9815;
	wire new_net_20678;
	wire new_net_20762;
	wire new_net_12968;
	wire new_net_17339;
	wire new_net_11552;
	wire new_net_10838;
	wire new_net_9028;
	wire new_net_11015;
	wire new_net_19574;
	wire new_net_20894;
	wire new_net_8900;
	wire _1088_;
	wire new_net_74;
	wire new_net_5031;
	wire new_net_8893;
	wire new_net_10247;
	wire new_net_13923;
	wire new_net_7466;
	wire new_net_17999;
	wire _0644_;
	wire _1022_;
	wire new_net_8988;
	wire new_net_17353;
	wire new_net_12410;
	wire new_net_16786;
	wire new_net_11975;
	wire new_net_13757;
	wire new_net_14121;
	wire new_net_14216;
	wire new_net_1014;
	wire new_net_20822;
	wire new_net_1315;
	wire new_net_6572;
	wire new_net_10252;
	wire new_net_8937;
	wire new_net_16676;
	wire new_net_21372;
	wire new_net_18795;
	wire _1023_;
	wire _0645_;
	wire new_net_77;
	wire new_net_8894;
	wire new_net_5027;
	wire new_net_8952;
	wire new_net_4163;
	wire new_net_8172;
	wire new_net_19375;
	wire new_net_8812;
	wire new_net_7468;
	wire new_net_8949;
	wire new_net_8167;
	wire new_net_9056;
	wire new_net_9357;
	wire _0146_;
	wire new_net_18938;
	wire new_net_18730;
	wire _1024_;
	wire _0646_;
	wire new_net_8810;
	wire new_net_20775;
	wire new_net_18672;
	wire new_net_4411;
	wire new_net_7462;
	wire new_net_13956;
	wire new_net_11333;
	wire new_net_19587;
	wire new_net_20420;
	wire new_net_19696;
	wire _1025_;
	wire new_net_278;
	wire _0647_;
	wire new_net_15817;
	wire new_net_4711;
	wire new_net_8934;
	wire new_net_8171;
	wire new_net_9582;
	wire new_net_9878;
	wire new_net_15250;
	wire new_net_5130;
	wire new_net_5708;
	wire new_net_13310;
	wire new_net_15628;
	wire new_net_12411;
	wire new_net_15581;
	wire new_net_17354;
	wire new_net_14344;
	wire new_net_14122;
	wire new_net_18861;
	wire new_net_14528;
	wire new_net_1314;
	wire _0648_;
	wire _1026_;
	wire new_net_3913;
	wire new_net_8993;
	wire new_net_19215;
	wire new_net_20477;
	wire new_net_1775;
	wire new_net_4416;
	wire new_net_5124;
	wire new_net_7686;
	wire new_net_9050;
	wire new_net_9880;
	wire new_net_15828;
	wire new_net_18134;
	wire new_net_19376;
	wire new_net_17079;
	wire _0649_;
	wire _1027_;
	wire new_net_9879;
	wire new_net_8943;
	wire new_net_4346;
	wire new_net_4414;
	wire new_net_13922;
	wire new_net_9049;
	wire new_net_8762;
	wire new_net_10404;
	wire new_net_7628;
	wire new_net_19216;
	wire new_net_20776;
	wire _0650_;
	wire _1028_;
	wire new_net_5642;
	wire new_net_9573;
	wire new_net_13924;
	wire new_net_11334;
	wire new_net_8936;
	wire new_net_19588;
	wire new_net_20421;
	wire new_net_21380;
	wire new_net_1774;
	wire new_net_5128;
	wire new_net_7638;
	wire _0147_;
	wire new_net_21120;
	wire _0651_;
	wire _1029_;
	wire new_net_9578;
	wire new_net_12412;
	wire new_net_13759;
	wire new_net_15251;
	wire new_net_15582;
	wire new_net_8811;
	wire new_net_14345;
	wire new_net_15819;
	wire new_net_18021;
	wire new_net_21085;
	wire new_net_271;
	wire new_net_9358;
	wire new_net_9365;
	wire new_net_13955;
	wire new_net_10410;
	wire new_net_18947;
	wire new_net_20891;
	wire new_net_21371;
	wire _0652_;
	wire _1030_;
	wire new_net_6565;
	wire new_net_8809;
	wire new_net_18133;
	wire new_net_19377;
	wire new_net_4713;
	wire new_net_7132;
	wire new_net_9051;
	wire new_net_9583;
	wire new_net_11629;
	wire new_net_21381;
	wire _0653_;
	wire _1031_;
	wire new_net_6834;
	wire new_net_8806;
	wire new_net_15820;
	wire new_net_5127;
	wire new_net_7136;
	wire new_net_7634;
	wire new_net_20479;
	wire new_net_21056;
	wire new_net_3361;
	wire new_net_5129;
	wire new_net_9364;
	wire new_net_13925;
	wire new_net_11335;
	wire new_net_8770;
	wire new_net_19589;
	wire new_net_20422;
	wire new_net_5055;
	wire new_net_18215;
	wire _0654_;
	wire _1032_;
	wire new_net_279;
	wire new_net_9048;
	wire _1778_;
	wire new_net_7637;
	wire new_net_19664;
	wire new_net_21164;
	wire new_net_3673;
	wire new_net_12413;
	wire new_net_13760;
	wire new_net_15252;
	wire new_net_17356;
	wire new_net_15583;
	wire new_net_14346;
	wire new_net_16789;
	wire new_net_14124;
	wire new_net_14219;
	wire _0655_;
	wire _1033_;
	wire new_net_5647;
	wire new_net_13954;
	wire new_net_8814;
	wire new_net_20356;
	wire new_net_17867;
	wire new_net_3437;
	wire new_net_9354;
	wire new_net_10257;
	wire new_net_15827;
	wire new_net_8766;
	wire new_net_18131;
	wire new_net_18946;
	wire new_net_19378;
	wire new_net_18980;
	wire new_net_18417;
	wire new_net_17040;
	wire new_net_270;
	wire new_net_1777;
	wire _0656_;
	wire _1034_;
	wire new_net_1320;
	wire new_net_8896;
	wire new_net_3679;
	wire new_net_1780;
	wire new_net_2929;
	wire new_net_68;
	wire new_net_5368;
	wire new_net_9359;
	wire new_net_7012;
	wire new_net_8950;
	wire new_net_6842;
	wire new_net_8944;
	wire _0657_;
	wire _1035_;
	wire new_net_9883;
	wire new_net_8159;
	wire new_net_13926;
	wire new_net_6569;
	wire new_net_8813;
	wire new_net_11336;
	wire new_net_5132;
	wire new_net_7463;
	wire new_net_1316;
	wire new_net_4412;
	wire new_net_8989;
	wire new_net_21373;
	wire new_net_11979;
	wire new_net_13313;
	wire new_net_15631;
	wire _0658_;
	wire _1036_;
	wire new_net_4342;
	wire new_net_5125;
	wire new_net_12414;
	wire new_net_13761;
	wire new_net_15253;
	wire new_net_4489;
	wire new_net_1322;
	wire new_net_6835;
	wire new_net_13953;
	wire new_net_10246;
	wire new_net_5131;
	wire new_net_7135;
	wire _1037_;
	wire _0659_;
	wire new_net_1318;
	wire new_net_9356;
	wire new_net_8897;
	wire new_net_10253;
	wire new_net_19379;
	wire new_net_18510;
	wire new_net_10254;
	wire new_net_8173;
	wire new_net_18945;
	wire new_net_20991;
	wire _1281_;
	wire _0660_;
	wire _1038_;
	wire new_net_5030;
	wire new_net_4413;
	wire new_net_18126;
	wire new_net_4407;
	wire new_net_7631;
	wire new_net_13927;
	wire new_net_6571;
	wire new_net_19591;
	wire new_net_20424;
	wire _0661_;
	wire _1039_;
	wire new_net_1317;
	wire new_net_5032;
	wire new_net_8808;
	wire new_net_8764;
	wire new_net_18132;
	wire new_net_205;
	wire new_net_18000;
	wire new_net_277;
	wire new_net_2933;
	wire new_net_4344;
	wire new_net_5562;
	wire new_net_7630;
	wire new_net_11980;
	wire new_net_13314;
	wire new_net_15632;
	wire new_net_12415;
	wire new_net_13762;
	wire _0662_;
	wire _1040_;
	wire new_net_5561;
	wire new_net_13952;
	wire new_net_3912;
	wire new_net_12021;
	wire new_net_14638;
	wire new_net_8174;
	wire new_net_18796;
	wire new_net_18377;
	wire new_net_14742;
	wire new_net_5643;
	wire new_net_6832;
	wire new_net_8948;
	wire new_net_9367;
	wire new_net_15826;
	wire new_net_10401;
	wire new_net_19380;
	wire new_net_18295;
	wire _0663_;
	wire _1041_;
	wire new_net_2936;
	wire new_net_8939;
	wire new_net_18731;
	wire _1015_;
	wire new_net_269;
	wire new_net_8899;
	wire new_net_10250;
	wire new_net_10409;
	wire new_net_8165;
	wire new_net_18944;
	wire new_net_21379;
	wire new_net_18673;
	wire _0664_;
	wire _1042_;
	wire new_net_1776;
	wire new_net_13928;
	wire new_net_7464;
	wire new_net_18129;
	wire new_net_19256;
	wire new_net_19592;
	wire new_net_20425;
	wire new_net_21196;
	wire new_net_1779;
	wire new_net_3678;
	wire new_net_9887;
	wire new_net_16854;
	wire new_net_14456;
	wire _0665_;
	wire _1043_;
	wire new_net_4410;
	wire new_net_11981;
	wire new_net_13315;
	wire new_net_15633;
	wire new_net_9055;
	wire new_net_12416;
	wire new_net_13763;
	wire new_net_18862;
	wire new_net_6566;
	wire new_net_8995;
	wire new_net_13951;
	wire new_net_8955;
	wire new_net_8771;
	wire _0666_;
	wire _1044_;
	wire new_net_5644;
	wire new_net_8987;
	wire new_net_9366;
	wire new_net_4161;
	wire new_net_8941;
	wire new_net_19381;
	wire new_net_1319;
	wire new_net_2935;
	wire new_net_4165;
	wire new_net_9363;
	wire new_net_11337;
	wire new_net_10403;
	wire new_net_3677;
	wire new_net_4343;
	wire _0667_;
	wire new_net_71;
	wire _1045_;
	wire new_net_275;
	wire new_net_2931;
	wire new_net_9581;
	wire new_net_8892;
	wire new_net_9369;
	wire new_net_20450;
	wire new_net_2937;
	wire new_net_13929;
	wire new_net_18943;
	wire new_net_19593;
	wire new_net_20426;
	wire _0668_;
	wire new_net_72;
	wire _1046_;
	wire new_net_3364;
	wire new_net_9576;
	wire new_net_10255;
	wire new_net_5126;
	wire new_net_18130;
	wire new_net_3757;
	wire new_net_21121;
	wire new_net_14457;
	wire new_net_5029;
	wire new_net_5646;
	wire new_net_5710;
	wire new_net_11982;
	wire new_net_13316;
	wire new_net_15634;
	wire new_net_12417;
	wire new_net_13764;
	wire new_net_15256;
	wire new_net_18022;
	wire new_net_21086;
	wire new_net_8170;
	wire _0669_;
	wire _1047_;
	wire new_net_13950;
	wire new_net_7467;
	wire new_net_8938;
	wire new_net_20892;
	wire new_net_273;
	wire new_net_9888;
	wire new_net_15825;
	wire new_net_8768;
	wire new_net_10407;
	wire new_net_19382;
	wire new_net_21377;
	wire _0670_;
	wire _1048_;
	wire new_net_272;
	wire new_net_8160;
	wire new_net_15818;
	wire new_net_20360;
	wire new_net_19172;
	wire new_net_274;
	wire new_net_6881;
	wire new_net_7685;
	wire new_net_8996;
	wire new_net_8935;
	wire new_net_19217;
	wire new_net_20777;
	wire _0671_;
	wire _1049_;
	wire new_net_8990;
	wire new_net_13930;
	wire new_net_11338;
	wire new_net_18128;
	wire new_net_19218;
	wire new_net_19594;
	wire new_net_20427;
	wire new_net_18216;
	wire new_net_7636;
	wire new_net_9368;
	wire new_net_9580;
	wire new_net_10408;
	wire new_net_18942;
	wire new_net_20357;
	wire new_net_4223;
	wire new_net_19665;
	wire _0672_;
	wire _1050_;
	wire new_net_3675;
	wire new_net_4345;
	wire new_net_14458;
	wire new_net_11983;
	wire new_net_13317;
	wire new_net_15635;
	wire new_net_5648;
	wire new_net_7687;
	wire new_net_4160;
	wire new_net_4348;
	wire new_net_13949;
	wire new_net_6568;
	wire new_net_6843;
	wire new_net_19219;
	wire new_net_19254;
	wire new_net_20181;
	wire new_net_4167;
	wire _0673_;
	wire _1051_;
	wire new_net_76;
	wire new_net_5367;
	wire new_net_9361;
	wire new_net_5713;
	wire new_net_17868;
	wire new_net_19383;
	wire new_net_3676;
	wire new_net_8156;
	wire new_net_7469;
	wire new_net_8954;
	wire _0674_;
	wire _1052_;
	wire new_net_67;
	wire new_net_10248;
	wire new_net_8958;
	wire new_net_19255;
	wire new_net_20778;
	wire new_net_4833;
	wire new_net_280;
	wire new_net_1321;
	wire new_net_4715;
	wire new_net_9886;
	wire new_net_10249;
	wire new_net_13931;
	wire new_net_11339;
	wire new_net_5712;
	wire new_net_18127;
	wire new_net_19595;
	wire new_net_8933;
	wire _1053_;
	wire _0675_;
	wire new_net_6567;
	wire new_net_7011;
	wire new_net_7133;
	wire new_net_7465;
	wire new_net_8767;
	wire new_net_14459;
	wire new_net_11984;
	wire new_net_13318;
	wire new_net_15636;
	wire new_net_9574;
	wire new_net_9881;
	wire new_net_12419;
	wire new_net_13766;
	wire new_net_4409;
	wire _1054_;
	wire new_net_281;
	wire new_net_1782;
	wire _0676_;
	wire new_net_8168;
	wire new_net_9362;
	wire new_net_13948;
	wire new_net_15822;
	wire new_net_668;
	wire new_net_18636;
	wire new_net_6840;
	wire new_net_2932;
	wire new_net_4712;
	wire new_net_9885;
	wire new_net_8994;
	wire new_net_10256;
	wire new_net_15824;
	wire new_net_19384;
	wire new_net_19335;
	wire new_net_18511;
	wire new_net_8769;
	wire _0677_;
	wire _1055_;
	wire new_net_3360;
	wire new_net_9575;
	wire new_net_8991;
	wire new_net_21376;
	wire new_net_2930;
	wire new_net_7137;
	wire new_net_8807;
	wire new_net_18937;
	wire new_net_20779;
	wire new_net_4714;
	wire new_net_10405;
	wire _0678_;
	wire _1056_;
	wire new_net_3674;
	wire new_net_10251;
	wire new_net_13932;
	wire new_net_11340;
	wire new_net_19596;
	wire new_net_15538;
	wire new_net_5641;
	wire new_net_6833;
	wire new_net_8805;
	wire new_net_9882;
	wire new_net_201;
	wire new_net_18001;
	wire _0679_;
	wire _1057_;
	wire new_net_14460;
	wire new_net_15259;
	wire new_net_7629;
	wire new_net_11985;
	wire new_net_13319;
	wire new_net_15637;
	wire new_net_12420;
	wire new_net_13767;
	wire new_net_8940;
	wire new_net_1323;
	wire new_net_4418;
	wire new_net_13947;
	wire new_net_6573;
	wire new_net_18125;
	wire new_net_18940;
	wire new_net_18797;
	wire new_net_18378;
	wire new_net_2934;
	wire _1058_;
	wire new_net_1778;
	wire _0680_;
	wire new_net_4341;
	wire new_net_8997;
	wire new_net_8763;
	wire new_net_8898;
	wire new_net_9353;
	wire new_net_3349;
	wire new_net_9054;
	wire new_net_75;
	wire new_net_5028;
	wire new_net_5645;
	wire new_net_13946;
	wire _0681_;
	wire _1059_;
	wire new_net_3911;
	wire new_net_8942;
	wire new_net_7635;
	wire new_net_9355;
	wire new_net_8992;
	wire new_net_18732;
	wire new_net_20780;
	wire new_net_18674;
	wire new_net_73;
	wire new_net_1781;
	wire new_net_4408;
	wire new_net_8169;
	wire new_net_7688;
	wire new_net_9360;
	wire new_net_8158;
	wire new_net_11341;
	wire new_net_18865;
	wire new_net_19597;
	wire _0682_;
	wire _1060_;
	wire new_net_8765;
	wire new_net_9052;
	wire new_net_9579;
	wire new_net_20540;
	wire new_net_21402;
	wire new_net_14132;
	wire new_net_14227;
	wire new_net_70;
	wire new_net_4166;
	wire new_net_4347;
	wire new_net_8166;
	wire new_net_14461;
	wire new_net_11986;
	wire new_net_13320;
	wire new_net_15638;
	wire new_net_18863;
	wire new_net_69;
	wire _0683_;
	wire _1061_;
	wire new_net_13933;
	wire new_net_4162;
	wire new_net_8956;
	wire new_net_9057;
	wire new_net_10402;
	wire new_net_15823;
	wire new_net_18939;
	wire new_net_19386;
	wire new_net_20358;
	wire new_net_18172;
	wire new_net_5711;
	wire new_net_7134;
	wire _0684_;
	wire _1062_;
	wire new_net_276;
	wire new_net_4415;
	wire new_net_9053;
	wire new_net_9577;
	wire new_net_7131;
	wire new_net_10411;
	wire new_net_9884;
	wire new_net_15175;
	wire new_net_20781;
	wire _1063_;
	wire _0685_;
	wire new_net_8895;
	wire new_net_7633;
	wire new_net_9877;
	wire new_net_8157;
	wire new_net_11342;
	wire new_net_18123;
	wire new_net_19598;
	wire new_net_20431;
	wire _0154_;
	wire new_net_21122;
	wire new_net_1959;
	wire new_net_2137;
	wire new_net_3505;
	wire new_net_7164;
	wire new_net_7900;
	wire new_net_19983;
	wire new_net_20031;
	wire new_net_18023;
	wire new_net_21087;
	wire new_net_16822;
	wire _1526_;
	wire _1820_;
	wire new_net_11844;
	wire new_net_12458;
	wire new_net_16762;
	wire new_net_3485;
	wire new_net_4877;
	wire new_net_12636;
	wire new_net_13415;
	wire new_net_20893;
	wire new_net_1130;
	wire new_net_7354;
	wire new_net_7904;
	wire new_net_8116;
	wire new_net_9483;
	wire new_net_19552;
	wire new_net_20655;
	wire new_net_13758;
	wire _1527_;
	wire new_net_1964;
	wire _1821_;
	wire new_net_3486;
	wire new_net_7882;
	wire new_net_2503;
	wire new_net_18948;
	wire new_net_20665;
	wire new_net_21201;
	wire new_net_1482;
	wire new_net_1129;
	wire new_net_4736;
	wire new_net_19576;
	wire _1528_;
	wire new_net_1478;
	wire new_net_2143;
	wire _1822_;
	wire new_net_6613;
	wire new_net_8780;
	wire new_net_3307;
	wire new_net_3356;
	wire new_net_20666;
	wire new_net_18217;
	wire new_net_1628;
	wire new_net_2357;
	wire new_net_5071;
	wire new_net_11040;
	wire new_net_11565;
	wire new_net_7283;
	wire new_net_9305;
	wire new_net_11122;
	wire new_net_19666;
	wire _1823_;
	wire new_net_2394;
	wire _1529_;
	wire new_net_10338;
	wire new_net_6056;
	wire new_net_7159;
	wire new_net_19984;
	wire new_net_20032;
	wire new_net_15557;
	wire new_net_16823;
	wire new_net_2400;
	wire new_net_3184;
	wire new_net_4481;
	wire new_net_6325;
	wire new_net_11845;
	wire new_net_12459;
	wire new_net_16763;
	wire new_net_12637;
	wire new_net_17869;
	wire new_net_15806;
	wire _1824_;
	wire _1530_;
	wire new_net_3189;
	wire new_net_6612;
	wire new_net_15816;
	wire new_net_2392;
	wire new_net_3491;
	wire new_net_9134;
	wire new_net_9481;
	wire new_net_19131;
	wire _1825_;
	wire new_net_1627;
	wire _1531_;
	wire new_net_1961;
	wire new_net_9480;
	wire new_net_4871;
	wire new_net_6054;
	wire new_net_10048;
	wire new_net_9587;
	wire new_net_21200;
	wire new_net_19454;
	wire new_net_2509;
	wire new_net_1444;
	wire new_net_1481;
	wire new_net_1630;
	wire new_net_2141;
	wire new_net_4728;
	wire new_net_4872;
	wire new_net_6052;
	wire _1826_;
	wire _1532_;
	wire new_net_7356;
	wire new_net_3186;
	wire new_net_11041;
	wire new_net_13003;
	wire new_net_6058;
	wire new_net_11566;
	wire new_net_11123;
	wire new_net_4443;
	wire new_net_1446;
	wire new_net_2140;
	wire new_net_3358;
	wire new_net_8114;
	wire new_net_10330;
	wire new_net_9592;
	wire new_net_19985;
	wire new_net_20033;
	wire new_net_15558;
	wire _1827_;
	wire new_net_2355;
	wire _1533_;
	wire new_net_16824;
	wire new_net_11846;
	wire new_net_12460;
	wire new_net_16764;
	wire new_net_12638;
	wire new_net_13417;
	wire new_net_18395;
	wire new_net_2504;
	wire new_net_2138;
	wire new_net_19334;
	wire new_net_18512;
	wire _1828_;
	wire new_net_2362;
	wire _1534_;
	wire new_net_6048;
	wire new_net_21199;
	wire _1288_;
	wire new_net_2390;
	wire new_net_2512;
	wire new_net_4733;
	wire new_net_6606;
	wire new_net_20182;
	wire _1829_;
	wire _1535_;
	wire new_net_3487;
	wire new_net_3423;
	wire new_net_15539;
	wire new_net_1486;
	wire new_net_3188;
	wire new_net_6331;
	wire new_net_11567;
	wire new_net_9588;
	wire new_net_9482;
	wire new_net_11124;
	wire new_net_11042;
	wire new_net_11918;
	wire new_net_19553;
	wire new_net_18002;
	wire new_net_7357;
	wire _1830_;
	wire _1536_;
	wire new_net_5062;
	wire new_net_10050;
	wire new_net_10599;
	wire new_net_7907;
	wire new_net_19986;
	wire new_net_20034;
	wire new_net_20664;
	wire new_net_19461;
	wire new_net_14501;
	wire new_net_15559;
	wire new_net_2358;
	wire new_net_1133;
	wire new_net_1242;
	wire new_net_1479;
	wire new_net_4734;
	wire new_net_16825;
	wire new_net_11847;
	wire new_net_14512;
	wire new_net_18798;
	wire new_net_18379;
	wire new_net_15810;
	wire _1831_;
	wire new_net_1245;
	wire _1537_;
	wire new_net_9140;
	wire new_net_1443;
	wire new_net_3339;
	wire new_net_10046;
	wire new_net_3855;
	wire new_net_7899;
	wire new_net_15815;
	wire new_net_1441;
	wire new_net_1453;
	wire new_net_3196;
	wire new_net_8122;
	wire new_net_13958;
	wire new_net_16266;
	wire new_net_18733;
	wire _1538_;
	wire new_net_1447;
	wire _1832_;
	wire new_net_1626;
	wire new_net_7351;
	wire new_net_6332;
	wire new_net_3489;
	wire new_net_10600;
	wire new_net_7281;
	wire new_net_8777;
	wire new_net_18675;
	wire new_net_1957;
	wire new_net_2136;
	wire new_net_1241;
	wire new_net_9135;
	wire new_net_6327;
	wire new_net_10051;
	wire new_net_7161;
	wire new_net_11125;
	wire _1539_;
	wire _1833_;
	wire new_net_3191;
	wire new_net_5068;
	wire new_net_6323;
	wire new_net_6607;
	wire new_net_11043;
	wire new_net_11568;
	wire new_net_8779;
	wire new_net_1460;
	wire new_net_1632;
	wire new_net_4480;
	wire new_net_7350;
	wire new_net_7160;
	wire new_net_7291;
	wire new_net_9299;
	wire new_net_19987;
	wire new_net_20035;
	wire new_net_18864;
	wire new_net_15869;
	wire new_net_15560;
	wire _1540_;
	wire _1834_;
	wire new_net_16826;
	wire new_net_11848;
	wire new_net_12462;
	wire new_net_12640;
	wire new_net_13419;
	wire new_net_14513;
	wire new_net_6608;
	wire new_net_1137;
	wire new_net_3185;
	wire new_net_5067;
	wire new_net_7901;
	wire new_net_7879;
	wire new_net_20663;
	wire new_net_18471;
	wire new_net_7902;
	wire _1541_;
	wire new_net_1477;
	wire _1835_;
	wire new_net_9132;
	wire new_net_6324;
	wire new_net_1026;
	wire new_net_17422;
	wire new_net_2139;
	wire new_net_1485;
	wire new_net_3502;
	wire new_net_6610;
	wire new_net_10595;
	wire new_net_1345;
	wire _1542_;
	wire new_net_1965;
	wire new_net_2144;
	wire new_net_2365;
	wire new_net_1631;
	wire new_net_8120;
	wire _1836_;
	wire new_net_1132;
	wire new_net_10598;
	wire new_net_3854;
	wire new_net_11126;
	wire new_net_1960;
	wire new_net_2361;
	wire new_net_3490;
	wire new_net_5066;
	wire new_net_11044;
	wire new_net_14502;
	wire new_net_11569;
	wire new_net_19555;
	wire _1543_;
	wire _1837_;
	wire new_net_2393;
	wire new_net_15807;
	wire new_net_8117;
	wire new_net_3354;
	wire new_net_7286;
	wire new_net_9308;
	wire new_net_19988;
	wire new_net_20036;
	wire new_net_21123;
	wire new_net_18024;
	wire new_net_21088;
	wire new_net_15870;
	wire new_net_17760;
	wire new_net_6057;
	wire new_net_14631;
	wire new_net_15561;
	wire new_net_16827;
	wire new_net_11849;
	wire new_net_12463;
	wire new_net_16767;
	wire new_net_12641;
	wire new_net_1963;
	wire _1544_;
	wire new_net_1440;
	wire new_net_1489;
	wire new_net_1244;
	wire new_net_7355;
	wire new_net_2396;
	wire new_net_4731;
	wire new_net_13651;
	wire new_net_1135;
	wire _0875_;
	wire new_net_1448;
	wire new_net_2510;
	wire new_net_3383;
	wire new_net_3504;
	wire new_net_4873;
	wire new_net_15814;
	wire new_net_8123;
	wire new_net_6330;
	wire new_net_9300;
	wire _1545_;
	wire new_net_1958;
	wire new_net_1459;
	wire new_net_2399;
	wire new_net_4482;
	wire new_net_4876;
	wire new_net_10596;
	wire new_net_9303;
	wire new_net_21094;
	wire new_net_19577;
	wire new_net_17718;
	wire new_net_3187;
	wire new_net_6615;
	wire new_net_9484;
	wire new_net_10336;
	wire new_net_7883;
	wire new_net_20661;
	wire _1546_;
	wire new_net_11570;
	wire new_net_11127;
	wire new_net_11045;
	wire new_net_10337;
	wire new_net_9141;
	wire new_net_19556;
	wire new_net_19449;
	wire new_net_2356;
	wire new_net_1476;
	wire new_net_8118;
	wire new_net_10601;
	wire new_net_19667;
	wire new_net_19989;
	wire new_net_12820;
	wire new_net_15871;
	wire new_net_16828;
	wire new_net_14515;
	wire _1547_;
	wire new_net_3190;
	wire new_net_13421;
	wire new_net_15562;
	wire new_net_12642;
	wire new_net_17761;
	wire new_net_7167;
	wire new_net_2395;
	wire new_net_3852;
	wire new_net_8119;
	wire new_net_17870;
	wire new_net_7158;
	wire new_net_7282;
	wire new_net_8782;
	wire _1548_;
	wire new_net_1450;
	wire new_net_5064;
	wire new_net_9133;
	wire new_net_9487;
	wire new_net_20660;
	wire new_net_9306;
	wire new_net_1454;
	wire new_net_1480;
	wire new_net_1136;
	wire new_net_10332;
	wire new_net_20656;
	wire new_net_19495;
	wire new_net_9586;
	wire new_net_2398;
	wire _1549_;
	wire new_net_15805;
	wire new_net_9139;
	wire new_net_7880;
	wire new_net_11128;
	wire new_net_2511;
	wire new_net_3195;
	wire new_net_11046;
	wire new_net_11571;
	wire new_net_19557;
	wire new_net_1243;
	wire new_net_1461;
	wire new_net_2507;
	wire _1550_;
	wire new_net_19990;
	wire new_net_12821;
	wire new_net_14820;
	wire new_net_15872;
	wire new_net_17762;
	wire new_net_1624;
	wire new_net_2142;
	wire new_net_3352;
	wire new_net_15563;
	wire new_net_7352;
	wire new_net_16829;
	wire new_net_18396;
	wire _1551_;
	wire new_net_9589;
	wire _0819_;
	wire new_net_3501;
	wire new_net_6614;
	wire new_net_7280;
	wire new_net_15813;
	wire new_net_12319;
	wire _1552_;
	wire new_net_15808;
	wire new_net_7353;
	wire new_net_8121;
	wire new_net_6326;
	wire new_net_3506;
	wire new_net_18714;
	wire new_net_1456;
	wire new_net_1967;
	wire new_net_9590;
	wire new_net_6322;
	wire new_net_10339;
	wire _1553_;
	wire new_net_11129;
	wire new_net_11047;
	wire new_net_11572;
	wire new_net_19558;
	wire new_net_18003;
	wire new_net_7157;
	wire new_net_8781;
	wire new_net_2364;
	wire new_net_4874;
	wire new_net_9585;
	wire new_net_10047;
	wire new_net_19991;
	wire new_net_12822;
	wire new_net_14821;
	wire _1554_;
	wire new_net_4730;
	wire new_net_15873;
	wire new_net_17763;
	wire new_net_15564;
	wire new_net_16830;
	wire new_net_11852;
	wire new_net_12466;
	wire new_net_1599;
	wire new_net_18799;
	wire new_net_1488;
	wire new_net_1969;
	wire new_net_3488;
	wire new_net_3507;
	wire new_net_4875;
	wire new_net_10045;
	wire new_net_18380;
	wire new_net_3455;
	wire new_net_7288;
	wire _1555_;
	wire new_net_1484;
	wire new_net_5061;
	wire new_net_6051;
	wire new_net_7885;
	wire new_net_13959;
	wire new_net_16267;
	wire new_net_3335;
	wire new_net_5301;
	wire new_net_10604;
	wire new_net_18734;
	wire new_net_18676;
	wire new_net_18634;
	wire new_net_7166;
	wire _1556_;
	wire new_net_1462;
	wire new_net_9138;
	wire new_net_4479;
	wire new_net_10335;
	wire new_net_11573;
	wire new_net_1966;
	wire new_net_1131;
	wire new_net_2505;
	wire new_net_11130;
	wire new_net_7349;
	wire new_net_8115;
	wire new_net_6616;
	wire new_net_9486;
	wire new_net_11048;
	wire _1557_;
	wire new_net_7886;
	wire new_net_19992;
	wire new_net_13720;
	wire new_net_7284;
	wire new_net_12823;
	wire new_net_14822;
	wire new_net_1449;
	wire new_net_1956;
	wire new_net_1452;
	wire new_net_7903;
	wire new_net_15874;
	wire new_net_17764;
	wire new_net_5949;
	wire new_net_3682;
	wire new_net_3856;
	wire _1558_;
	wire new_net_9584;
	wire new_net_3197;
	wire new_net_4729;
	wire new_net_10333;
	wire new_net_18171;
	wire new_net_1457;
	wire new_net_15812;
	wire new_net_20659;
	wire new_net_3405;
	wire new_net_7162;
	wire _1559_;
	wire new_net_1445;
	wire new_net_6611;
	wire new_net_10049;
	wire new_net_7285;
	wire new_net_9307;
	wire new_net_1487;
	wire new_net_1968;
	wire new_net_2502;
	wire new_net_9137;
	wire new_net_6329;
	wire new_net_10334;
	wire new_net_903;
	wire new_net_11574;
	wire new_net_7163;
	wire new_net_7290;
	wire _1560_;
	wire new_net_1134;
	wire new_net_2506;
	wire new_net_7905;
	wire new_net_11131;
	wire new_net_15809;
	wire new_net_4737;
	wire new_net_20332;
	wire _0161_;
	wire new_net_7289;
	wire new_net_1629;
	wire new_net_3199;
	wire new_net_19993;
	wire new_net_21124;
	wire new_net_18025;
	wire new_net_21089;
	wire new_net_13721;
	wire new_net_12824;
	wire new_net_14823;
	wire _1561_;
	wire new_net_1455;
	wire new_net_2359;
	wire new_net_15875;
	wire new_net_17765;
	wire new_net_15566;
	wire new_net_5063;
	wire new_net_18901;
	wire new_net_9304;
	wire new_net_2397;
	wire new_net_3193;
	wire new_net_9131;
	wire new_net_2075;
	wire new_net_15717;
	wire new_net_3853;
	wire _1562_;
	wire new_net_1483;
	wire new_net_1962;
	wire new_net_9301;
	wire new_net_1633;
	wire new_net_2391;
	wire new_net_4483;
	wire new_net_1127;
	wire new_net_1442;
	wire new_net_4485;
	wire new_net_9309;
	wire new_net_7359;
	wire new_net_14694;
	wire new_net_6328;
	wire new_net_7884;
	wire new_net_10597;
	wire _1563_;
	wire new_net_1439;
	wire new_net_3353;
	wire new_net_20657;
	wire new_net_3540;
	wire new_net_11575;
	wire new_net_3484;
	wire new_net_3851;
	wire new_net_4732;
	wire new_net_11132;
	wire new_net_11050;
	wire new_net_19561;
	wire new_net_1128;
	wire new_net_1625;
	wire _1564_;
	wire new_net_2133;
	wire new_net_9130;
	wire new_net_9478;
	wire new_net_3198;
	wire new_net_19994;
	wire new_net_4218;
	wire new_net_19668;
	wire new_net_13544;
	wire new_net_14508;
	wire new_net_14637;
	wire new_net_13722;
	wire new_net_1458;
	wire new_net_2508;
	wire new_net_12825;
	wire new_net_14824;
	wire new_net_15876;
	wire new_net_17766;
	wire _1565_;
	wire new_net_3192;
	wire new_net_17871;
	wire new_net_6049;
	wire new_net_7878;
	wire new_net_4735;
	wire new_net_4878;
	wire new_net_15811;
	wire new_net_8919;
	wire new_net_2360;
	wire _1566_;
	wire new_net_5065;
	wire new_net_4870;
	wire new_net_20658;
	wire new_net_1451;
	wire new_net_2363;
	wire new_net_2135;
	wire new_net_1246;
	wire new_net_7287;
	wire new_net_9302;
	wire new_net_17661;
	wire new_net_7881;
	wire new_net_11576;
	wire _1567_;
	wire new_net_2134;
	wire new_net_11133;
	wire new_net_4738;
	wire new_net_11051;
	wire new_net_19562;
	wire new_net_21198;
	wire new_net_9329;
	wire new_net_9801;
	wire new_net_50;
	wire new_net_1818;
	wire new_net_5595;
	wire new_net_7096;
	wire new_net_19887;
	wire new_net_667;
	wire new_net_18397;
	wire new_net_4133;
	wire new_net_11785;
	wire new_net_12233;
	wire _0602_;
	wire new_net_1814;
	wire new_net_2308;
	wire new_net_12304;
	wire new_net_13781;
	wire new_net_8888;
	wire new_net_15829;
	wire new_net_39;
	wire new_net_2307;
	wire new_net_9191;
	wire new_net_19699;
	wire new_net_20622;
	wire new_net_18715;
	wire _0603_;
	wire new_net_5430;
	wire new_net_6725;
	wire _1295_;
	wire new_net_2896;
	wire new_net_2791;
	wire new_net_3998;
	wire new_net_8855;
	wire new_net_15592;
	wire new_net_4121;
	wire new_net_9957;
	wire new_net_15541;
	wire _0604_;
	wire new_net_3995;
	wire new_net_4782;
	wire new_net_5616;
	wire new_net_6718;
	wire new_net_7098;
	wire new_net_20052;
	wire new_net_20703;
	wire new_net_19129;
	wire new_net_18004;
	wire new_net_12753;
	wire new_net_2895;
	wire new_net_5620;
	wire new_net_11577;
	wire new_net_11424;
	wire new_net_11170;
	wire new_net_10933;
	wire new_net_13095;
	wire new_net_20478;
	wire new_net_20895;
	wire _0605_;
	wire new_net_2315;
	wire new_net_19888;
	wire new_net_1590;
	wire new_net_18800;
	wire new_net_18381;
	wire new_net_14378;
	wire new_net_5613;
	wire new_net_12234;
	wire new_net_12305;
	wire new_net_13782;
	wire new_net_15593;
	wire new_net_15830;
	wire new_net_14838;
	wire new_net_15878;
	wire new_net_17165;
	wire _0606_;
	wire new_net_2482;
	wire new_net_591;
	wire new_net_2306;
	wire new_net_19700;
	wire new_net_13960;
	wire new_net_16268;
	wire new_net_9323;
	wire new_net_1822;
	wire new_net_4129;
	wire new_net_4781;
	wire new_net_18735;
	wire new_net_18677;
	wire _0607_;
	wire new_net_1812;
	wire new_net_3426;
	wire new_net_4120;
	wire new_net_5429;
	wire new_net_8889;
	wire new_net_15594;
	wire new_net_6548;
	wire new_net_9683;
	wire new_net_20486;
	wire new_net_9321;
	wire new_net_2782;
	wire new_net_2404;
	wire new_net_3999;
	wire new_net_19220;
	wire new_net_20053;
	wire new_net_20704;
	wire new_net_7780;
	wire new_net_3372;
	wire new_net_11786;
	wire _0608_;
	wire new_net_2479;
	wire new_net_11578;
	wire new_net_11425;
	wire new_net_11171;
	wire new_net_10934;
	wire new_net_20896;
	wire new_net_19320;
	wire new_net_7774;
	wire new_net_14377;
	wire new_net_51;
	wire new_net_5705;
	wire new_net_6547;
	wire new_net_19889;
	wire new_net_12751;
	wire _0609_;
	wire new_net_43;
	wire new_net_2485;
	wire new_net_12235;
	wire new_net_12306;
	wire new_net_13783;
	wire new_net_15595;
	wire new_net_15831;
	wire new_net_14839;
	wire new_net_59;
	wire new_net_12752;
	wire new_net_5594;
	wire new_net_19701;
	wire new_net_20485;
	wire _0610_;
	wire new_net_832;
	wire new_net_9800;
	wire new_net_6720;
	wire new_net_603;
	wire new_net_2783;
	wire new_net_2310;
	wire new_net_2406;
	wire new_net_8884;
	wire new_net_5702;
	wire new_net_913;
	wire new_net_10419;
	wire new_net_2892;
	wire _0611_;
	wire new_net_7094;
	wire new_net_20054;
	wire new_net_20705;
	wire new_net_9950;
	wire new_net_2403;
	wire new_net_4152;
	wire new_net_5295;
	wire new_net_9799;
	wire new_net_11579;
	wire new_net_11426;
	wire new_net_11172;
	wire new_net_10935;
	wire new_net_20897;
	wire new_net_21125;
	wire new_net_18026;
	wire new_net_21090;
	wire new_net_14376;
	wire _0612_;
	wire new_net_1214;
	wire new_net_2481;
	wire new_net_2781;
	wire new_net_8891;
	wire new_net_6550;
	wire new_net_18807;
	wire new_net_19223;
	wire new_net_19890;
	wire new_net_2647;
	wire new_net_18902;
	wire new_net_11787;
	wire new_net_12750;
	wire new_net_1209;
	wire new_net_2409;
	wire new_net_3697;
	wire new_net_12236;
	wire new_net_4153;
	wire new_net_12307;
	wire new_net_13784;
	wire new_net_5614;
	wire _0882_;
	wire _0613_;
	wire new_net_2949;
	wire new_net_2415;
	wire new_net_3996;
	wire new_net_5591;
	wire new_net_19702;
	wire new_net_18525;
	wire new_net_5639;
	wire new_net_9958;
	wire new_net_45;
	wire new_net_597;
	wire new_net_4126;
	wire new_net_5621;
	wire new_net_5635;
	wire _0614_;
	wire new_net_3690;
	wire new_net_4130;
	wire new_net_7097;
	wire new_net_835;
	wire new_net_2483;
	wire new_net_3429;
	wire new_net_5432;
	wire new_net_6715;
	wire new_net_5053;
	wire new_net_20055;
	wire new_net_20706;
	wire new_net_6684;
	wire new_net_10936;
	wire new_net_10417;
	wire _0615_;
	wire new_net_3694;
	wire new_net_5808;
	wire new_net_11427;
	wire new_net_11173;
	wire new_net_20898;
	wire new_net_19669;
	wire new_net_14375;
	wire new_net_3695;
	wire new_net_4132;
	wire new_net_19891;
	wire new_net_16565;
	wire new_net_5633;
	wire new_net_13090;
	wire new_net_14208;
	wire new_net_7777;
	wire new_net_11788;
	wire new_net_12749;
	wire new_net_594;
	wire _0616_;
	wire new_net_4786;
	wire new_net_12237;
	wire new_net_17872;
	wire new_net_46;
	wire new_net_1813;
	wire new_net_2305;
	wire new_net_6726;
	wire new_net_15596;
	wire new_net_19703;
	wire new_net_7091;
	wire _0617_;
	wire new_net_4128;
	wire new_net_6670;
	wire new_net_11580;
	wire new_net_5615;
	wire new_net_6721;
	wire new_net_9185;
	wire _0618_;
	wire new_net_589;
	wire new_net_1823;
	wire new_net_4156;
	wire new_net_20056;
	wire new_net_20707;
	wire new_net_10937;
	wire new_net_593;
	wire new_net_1207;
	wire new_net_8885;
	wire new_net_11428;
	wire new_net_11174;
	wire new_net_20899;
	wire _0619_;
	wire new_net_1820;
	wire new_net_41;
	wire new_net_1217;
	wire new_net_2938;
	wire new_net_14374;
	wire new_net_8854;
	wire new_net_15597;
	wire new_net_19892;
	wire new_net_13089;
	wire new_net_14209;
	wire new_net_7775;
	wire new_net_5818;
	wire new_net_11789;
	wire new_net_12748;
	wire new_net_12238;
	wire new_net_12309;
	wire new_net_15834;
	wire new_net_14842;
	wire new_net_18398;
	wire new_net_10421;
	wire _0620_;
	wire new_net_2891;
	wire new_net_3693;
	wire new_net_5590;
	wire new_net_13723;
	wire new_net_15601;
	wire new_net_19704;
	wire new_net_20484;
	wire new_net_12321;
	wire new_net_7095;
	wire new_net_10022;
	wire new_net_602;
	wire new_net_833;
	wire new_net_2888;
	wire new_net_1216;
	wire new_net_2784;
	wire new_net_5815;
	wire new_net_8886;
	wire new_net_18716;
	wire new_net_20623;
	wire new_net_9190;
	wire new_net_2402;
	wire _0621_;
	wire new_net_2480;
	wire new_net_3689;
	wire new_net_5704;
	wire new_net_21394;
	wire new_net_5636;
	wire new_net_7092;
	wire new_net_10426;
	wire new_net_1815;
	wire new_net_1213;
	wire new_net_4122;
	wire new_net_20057;
	wire new_net_20708;
	wire new_net_13078;
	wire new_net_10938;
	wire new_net_1212;
	wire new_net_2786;
	wire new_net_2939;
	wire _0622_;
	wire new_net_11581;
	wire new_net_13786;
	wire new_net_11429;
	wire new_net_11175;
	wire new_net_10024;
	wire new_net_10424;
	wire new_net_1208;
	wire new_net_592;
	wire new_net_2313;
	wire new_net_4124;
	wire new_net_14373;
	wire new_net_9804;
	wire new_net_19893;
	wire new_net_13088;
	wire new_net_14210;
	wire new_net_9182;
	wire new_net_2947;
	wire _0623_;
	wire new_net_11790;
	wire new_net_12747;
	wire new_net_9802;
	wire new_net_12239;
	wire new_net_12310;
	wire new_net_12074;
	wire new_net_18382;
	wire new_net_18801;
	wire _1299_;
	wire new_net_9678;
	wire new_net_9183;
	wire new_net_2411;
	wire new_net_3698;
	wire new_net_4118;
	wire new_net_16137;
	wire new_net_19705;
	wire new_net_13961;
	wire new_net_16269;
	wire new_net_10425;
	wire _0624_;
	wire new_net_4119;
	wire new_net_6727;
	wire new_net_18736;
	wire new_net_1057;
	wire new_net_18678;
	wire new_net_1215;
	wire new_net_15598;
	wire new_net_20483;
	wire new_net_2701;
	wire new_net_9187;
	wire new_net_9960;
	wire _0625_;
	wire new_net_837;
	wire new_net_5814;
	wire new_net_9798;
	wire new_net_20058;
	wire new_net_20709;
	wire new_net_9679;
	wire new_net_14338;
	wire new_net_10020;
	wire new_net_10939;
	wire new_net_11582;
	wire new_net_8857;
	wire new_net_11430;
	wire new_net_11176;
	wire new_net_20901;
	wire new_net_10019;
	wire new_net_9952;
	wire _0626_;
	wire new_net_601;
	wire new_net_836;
	wire new_net_14372;
	wire new_net_5593;
	wire new_net_8887;
	wire new_net_19894;
	wire new_net_4116;
	wire new_net_13079;
	wire new_net_1817;
	wire new_net_13087;
	wire new_net_7779;
	wire new_net_44;
	wire new_net_14211;
	wire new_net_11791;
	wire new_net_12746;
	wire new_net_12240;
	wire _0627_;
	wire new_net_8860;
	wire new_net_9951;
	wire new_net_19706;
	wire new_net_20481;
	wire new_net_2790;
	wire new_net_4157;
	wire new_net_8856;
	wire new_net_10423;
	wire new_net_15599;
	wire new_net_19222;
	wire new_net_1018;
	wire new_net_20149;
	wire _0628_;
	wire new_net_49;
	wire new_net_2484;
	wire new_net_2943;
	wire new_net_600;
	wire new_net_831;
	wire new_net_7778;
	wire new_net_9953;
	wire new_net_3369;
	wire new_net_6724;
	wire new_net_10018;
	wire new_net_2941;
	wire new_net_2793;
	wire new_net_2408;
	wire new_net_8859;
	wire new_net_20059;
	wire new_net_20710;
	wire _0168_;
	wire new_net_10940;
	wire _0629_;
	wire new_net_1816;
	wire new_net_2412;
	wire new_net_11583;
	wire new_net_6728;
	wire new_net_11431;
	wire new_net_11177;
	wire new_net_20902;
	wire new_net_21126;
	wire new_net_18027;
	wire new_net_21091;
	wire new_net_2940;
	wire new_net_2898;
	wire new_net_4785;
	wire new_net_6668;
	wire new_net_9324;
	wire new_net_14371;
	wire new_net_10420;
	wire new_net_19895;
	wire new_net_18808;
	wire new_net_18903;
	wire new_net_4001;
	wire new_net_14845;
	wire new_net_15885;
	wire new_net_17172;
	wire new_net_13080;
	wire new_net_14339;
	wire new_net_7093;
	wire new_net_13086;
	wire new_net_14212;
	wire new_net_830;
	wire new_net_9327;
	wire new_net_19707;
	wire new_net_18526;
	wire new_net_2897;
	wire _0631_;
	wire new_net_4131;
	wire new_net_8858;
	wire new_net_19580;
	wire new_net_2894;
	wire new_net_2785;
	wire new_net_2950;
	wire new_net_5638;
	wire new_net_8849;
	wire new_net_10025;
	wire _0632_;
	wire new_net_1210;
	wire new_net_4123;
	wire new_net_4159;
	wire new_net_4787;
	wire new_net_5817;
	wire new_net_9184;
	wire new_net_20060;
	wire new_net_20711;
	wire new_net_11178;
	wire new_net_2945;
	wire new_net_2312;
	wire new_net_1206;
	wire new_net_3421;
	wire new_net_3692;
	wire new_net_11432;
	wire new_net_5596;
	wire new_net_11584;
	wire new_net_10941;
	wire new_net_9681;
	wire _0633_;
	wire new_net_2893;
	wire new_net_14370;
	wire new_net_15600;
	wire new_net_5587;
	wire new_net_19896;
	wire new_net_5706;
	wire new_net_14846;
	wire new_net_15886;
	wire new_net_9680;
	wire new_net_14340;
	wire new_net_13085;
	wire new_net_2309;
	wire new_net_52;
	wire new_net_8850;
	wire new_net_15838;
	wire new_net_17873;
	wire new_net_16165;
	wire new_net_3997;
	wire new_net_5634;
	wire new_net_598;
	wire new_net_2311;
	wire new_net_2948;
	wire _0634_;
	wire new_net_42;
	wire new_net_9955;
	wire new_net_4127;
	wire new_net_6669;
	wire new_net_7776;
	wire new_net_9186;
	wire new_net_10418;
	wire new_net_6719;
	wire new_net_5296;
	wire new_net_590;
	wire _0635_;
	wire new_net_2942;
	wire new_net_5431;
	wire new_net_20061;
	wire new_net_20712;
	wire new_net_11179;
	wire new_net_10942;
	wire _0636_;
	wire new_net_2788;
	wire new_net_9956;
	wire new_net_9322;
	wire new_net_11585;
	wire new_net_11433;
	wire new_net_20480;
	wire new_net_20904;
	wire new_net_6549;
	wire new_net_9682;
	wire new_net_2414;
	wire new_net_595;
	wire new_net_14369;
	wire new_net_5618;
	wire new_net_19897;
	wire new_net_4783;
	wire new_net_14847;
	wire new_net_17174;
	wire new_net_13082;
	wire new_net_14341;
	wire new_net_13084;
	wire new_net_14214;
	wire new_net_834;
	wire new_net_2405;
	wire _0637_;
	wire new_net_18399;
	wire new_net_2401;
	wire new_net_2899;
	wire new_net_2789;
	wire new_net_10021;
	wire new_net_19709;
	wire new_net_5812;
	wire new_net_596;
	wire _0638_;
	wire new_net_2946;
	wire new_net_10027;
	wire new_net_8851;
	wire new_net_15602;
	wire new_net_21398;
	wire new_net_20624;
	wire new_net_20997;
	wire new_net_18717;
	wire new_net_2794;
	wire new_net_3367;
	wire new_net_5592;
	wire new_net_5707;
	wire new_net_4117;
	wire new_net_47;
	wire _0639_;
	wire new_net_828;
	wire new_net_10416;
	wire new_net_4158;
	wire new_net_20062;
	wire new_net_20713;
	wire new_net_3691;
	wire new_net_11434;
	wire new_net_11180;
	wire new_net_2787;
	wire new_net_48;
	wire new_net_829;
	wire new_net_2410;
	wire new_net_5640;
	wire new_net_10943;
	wire new_net_11586;
	wire new_net_1071;
	wire new_net_6722;
	wire new_net_8853;
	wire new_net_15603;
	wire new_net_6716;
	wire new_net_40;
	wire new_net_1211;
	wire _0640_;
	wire new_net_1819;
	wire new_net_2889;
	wire new_net_7781;
	wire new_net_15840;
	wire new_net_14848;
	wire new_net_17175;
	wire new_net_13083;
	wire new_net_14342;
	wire new_net_5589;
	wire new_net_5809;
	wire new_net_14215;
	wire new_net_11795;
	wire new_net_12244;
	wire new_net_18802;
	wire new_net_8890;
	wire new_net_5811;
	wire _0641_;
	wire new_net_3696;
	wire new_net_10422;
	wire new_net_19710;
	wire new_net_13962;
	wire new_net_5617;
	wire new_net_5703;
	wire new_net_2486;
	wire new_net_38;
	wire new_net_1821;
	wire new_net_2413;
	wire new_net_10026;
	wire new_net_9954;
	wire new_net_18737;
	wire new_net_6717;
	wire new_net_5810;
	wire _0642_;
	wire new_net_3450;
	wire new_net_9326;
	wire new_net_14367;
	wire new_net_2704;
	wire new_net_15887;
	wire new_net_2478;
	wire new_net_2944;
	wire new_net_2314;
	wire new_net_2890;
	wire new_net_3424;
	wire new_net_4780;
	wire new_net_5637;
	wire new_net_9188;
	wire new_net_5135;
	wire new_net_5588;
	wire new_net_6723;
	wire new_net_11435;
	wire new_net_4784;
	wire new_net_11181;
	wire new_net_15891;
	wire new_net_5816;
	wire _0643_;
	wire new_net_599;
	wire new_net_2407;
	wire _0014_;
	wire new_net_24;
	wire new_net_5477;
	wire new_net_19856;
	wire new_net_19995;
	wire new_net_7971;
	wire new_net_17117;
	wire new_net_17613;
	wire new_net_8386;
	wire new_net_10502;
	wire new_net_2242;
	wire _1694_;
	wire new_net_12588;
	wire new_net_13369;
	wire new_net_11738;
	wire new_net_16146;
	wire new_net_3046;
	wire new_net_3614;
	wire new_net_4142;
	wire new_net_5040;
	wire new_net_7044;
	wire new_net_19460;
	wire new_net_20075;
	wire new_net_20280;
	wire new_net_16787;
	wire new_net_2236;
	wire _1695_;
	wire new_net_18;
	wire new_net_7424;
	wire new_net_316;
	wire new_net_2264;
	wire new_net_3610;
	wire new_net_4473;
	wire new_net_4666;
	wire new_net_20327;
	wire _1696_;
	wire new_net_2258;
	wire new_net_7748;
	wire new_net_20322;
	wire new_net_20963;
	wire new_net_21035;
	wire new_net_21276;
	wire new_net_21288;
	wire new_net_19155;
	wire new_net_21127;
	wire new_net_18028;
	wire new_net_21092;
	wire new_net_11146;
	wire new_net_12552;
	wire new_net_4139;
	wire new_net_4654;
	wire new_net_5041;
	wire new_net_18809;
	wire new_net_18904;
	wire new_net_3202;
	wire new_net_3733;
	wire new_net_7221;
	wire _1697_;
	wire new_net_317;
	wire new_net_2261;
	wire new_net_3615;
	wire new_net_6627;
	wire new_net_19857;
	wire new_net_19996;
	wire new_net_13655;
	wire new_net_17843;
	wire new_net_15720;
	wire _0889_;
	wire new_net_17118;
	wire new_net_16692;
	wire new_net_17614;
	wire new_net_16;
	wire new_net_3048;
	wire new_net_4669;
	wire new_net_12589;
	wire new_net_13370;
	wire new_net_17816;
	wire new_net_11739;
	wire new_net_18527;
	wire _1698_;
	wire new_net_19;
	wire new_net_2369;
	wire new_net_19309;
	wire new_net_19470;
	wire new_net_20281;
	wire new_net_8382;
	wire new_net_318;
	wire new_net_3211;
	wire new_net_3546;
	wire new_net_2982;
	wire _1699_;
	wire new_net_4056;
	wire new_net_4136;
	wire new_net_9136;
	wire new_net_8773;
	wire new_net_15686;
	wire new_net_19307;
	wire new_net_4471;
	wire new_net_8772;
	wire new_net_7050;
	wire new_net_9283;
	wire new_net_16351;
	wire new_net_20073;
	wire new_net_20325;
	wire new_net_20964;
	wire new_net_21036;
	wire new_net_21277;
	wire new_net_8640;
	wire new_net_11147;
	wire _1700_;
	wire new_net_8391;
	wire new_net_12551;
	wire new_net_7300;
	wire new_net_8638;
	wire new_net_7431;
	wire new_net_19468;
	wire new_net_19858;
	wire new_net_19997;
	wire new_net_20074;
	wire new_net_8215;
	wire new_net_21392;
	wire new_net_15198;
	wire new_net_16166;
	wire new_net_17119;
	wire new_net_17615;
	wire new_net_7222;
	wire _1701_;
	wire new_net_321;
	wire new_net_2241;
	wire new_net_16693;
	wire new_net_4134;
	wire new_net_12590;
	wire new_net_13371;
	wire new_net_2373;
	wire new_net_3735;
	wire new_net_4053;
	wire new_net_4472;
	wire new_net_7052;
	wire new_net_8383;
	wire new_net_19314;
	wire new_net_19469;
	wire new_net_20282;
	wire _1702_;
	wire new_net_5482;
	wire new_net_15685;
	wire new_net_8641;
	wire new_net_21;
	wire new_net_2234;
	wire new_net_3730;
	wire new_net_4665;
	wire new_net_5483;
	wire new_net_5995;
	wire new_net_6629;
	wire new_net_7051;
	wire new_net_3044;
	wire _1703_;
	wire new_net_17;
	wire new_net_314;
	wire new_net_20965;
	wire new_net_21037;
	wire new_net_21278;
	wire new_net_21290;
	wire new_net_11148;
	wire new_net_2378;
	wire new_net_2684;
	wire new_net_4476;
	wire new_net_10055;
	wire new_net_20321;
	wire new_net_5928;
	wire new_net_4469;
	wire _1704_;
	wire new_net_4650;
	wire new_net_19859;
	wire new_net_11999;
	wire new_net_14555;
	wire new_net_19998;
	wire new_net_15727;
	wire new_net_18400;
	wire _0833_;
	wire new_net_19329;
	wire new_net_17120;
	wire new_net_17616;
	wire new_net_7229;
	wire new_net_3050;
	wire new_net_5485;
	wire new_net_12550;
	wire new_net_12591;
	wire new_net_16694;
	wire new_net_6630;
	wire new_net_13725;
	wire new_net_12323;
	wire new_net_15676;
	wire new_net_3210;
	wire new_net_7228;
	wire _1705_;
	wire new_net_3870;
	wire new_net_20283;
	wire new_net_18718;
	wire new_net_7046;
	wire _1706_;
	wire new_net_4052;
	wire new_net_7749;
	wire new_net_10053;
	wire new_net_5039;
	wire new_net_20966;
	wire new_net_21038;
	wire new_net_21279;
	wire new_net_21291;
	wire new_net_4655;
	wire new_net_5480;
	wire new_net_15683;
	wire new_net_3208;
	wire new_net_11149;
	wire _1707_;
	wire new_net_4055;
	wire new_net_3612;
	wire new_net_1000;
	wire new_net_13372;
	wire new_net_20847;
	wire new_net_12028;
	wire new_net_14644;
	wire new_net_3866;
	wire new_net_4059;
	wire new_net_7042;
	wire new_net_8387;
	wire new_net_19312;
	wire new_net_19860;
	wire new_net_19999;
	wire new_net_18803;
	wire new_net_16150;
	wire new_net_17819;
	wire new_net_17121;
	wire new_net_17617;
	wire _1708_;
	wire new_net_25;
	wire new_net_4057;
	wire new_net_4137;
	wire new_net_12592;
	wire new_net_16695;
	wire new_net_13963;
	wire new_net_16271;
	wire new_net_4058;
	wire new_net_10499;
	wire new_net_20072;
	wire new_net_20284;
	wire _1709_;
	wire new_net_15;
	wire new_net_7428;
	wire new_net_5999;
	wire new_net_9277;
	wire new_net_3294;
	wire new_net_15684;
	wire new_net_6001;
	wire new_net_12549;
	wire new_net_19467;
	wire new_net_20328;
	wire new_net_7751;
	wire _1710_;
	wire new_net_4140;
	wire new_net_20967;
	wire new_net_21039;
	wire new_net_21280;
	wire new_net_21292;
	wire new_net_11150;
	wire new_net_4144;
	wire new_net_19310;
	wire new_net_13298;
	wire new_net_5947;
	wire new_net_3687;
	wire new_net_4648;
	wire new_net_3049;
	wire _1711_;
	wire new_net_2271;
	wire new_net_7224;
	wire new_net_7048;
	wire new_net_19861;
	wire new_net_20000;
	wire new_net_20323;
	wire new_net_16151;
	wire new_net_17820;
	wire new_net_17122;
	wire new_net_17618;
	wire new_net_12593;
	wire new_net_13373;
	wire new_net_16696;
	wire new_net_11743;
	wire new_net_21158;
	wire new_net_3206;
	wire _1712_;
	wire new_net_22;
	wire new_net_3868;
	wire new_net_7423;
	wire new_net_3611;
	wire new_net_2257;
	wire new_net_4672;
	wire new_net_20285;
	wire new_net_2368;
	wire new_net_322;
	wire new_net_4649;
	wire new_net_12548;
	wire new_net_16788;
	wire new_net_3203;
	wire new_net_3052;
	wire new_net_7225;
	wire new_net_7425;
	wire _1713_;
	wire new_net_20071;
	wire new_net_313;
	wire new_net_5484;
	wire new_net_20968;
	wire new_net_21040;
	wire new_net_21281;
	wire new_net_21293;
	wire new_net_21128;
	wire new_net_11151;
	wire _1714_;
	wire new_net_4141;
	wire new_net_4670;
	wire new_net_12546;
	wire new_net_5996;
	wire new_net_19466;
	wire new_net_20324;
	wire new_net_18810;
	wire new_net_16955;
	wire new_net_18905;
	wire new_net_19862;
	wire new_net_20001;
	wire new_net_15642;
	wire new_net_11744;
	wire new_net_16152;
	wire new_net_17821;
	wire new_net_3734;
	wire new_net_17123;
	wire new_net_17619;
	wire _1715_;
	wire new_net_2366;
	wire new_net_3201;
	wire new_net_7430;
	wire new_net_2473;
	wire new_net_15721;
	wire new_net_320;
	wire new_net_6003;
	wire new_net_10501;
	wire new_net_20286;
	wire new_net_18528;
	wire new_net_19582;
	wire new_net_7049;
	wire new_net_9278;
	wire new_net_3732;
	wire _1716_;
	wire new_net_5998;
	wire new_net_2266;
	wire new_net_3207;
	wire new_net_3737;
	wire new_net_4054;
	wire new_net_4667;
	wire new_net_10506;
	wire new_net_12547;
	wire new_net_19459;
	wire new_net_20070;
	wire _1717_;
	wire new_net_2262;
	wire new_net_3047;
	wire new_net_20969;
	wire new_net_21282;
	wire new_net_21294;
	wire new_net_11152;
	wire new_net_3043;
	wire new_net_3867;
	wire new_net_19313;
	wire new_net_19465;
	wire new_net_7043;
	wire new_net_9280;
	wire new_net_15678;
	wire new_net_3204;
	wire _1718_;
	wire new_net_7429;
	wire new_net_3609;
	wire new_net_19863;
	wire new_net_20002;
	wire new_net_20069;
	wire new_net_6628;
	wire new_net_7053;
	wire new_net_9276;
	wire new_net_11745;
	wire new_net_16153;
	wire new_net_17822;
	wire new_net_2260;
	wire new_net_3051;
	wire new_net_4468;
	wire new_net_8636;
	wire new_net_16167;
	wire _1719_;
	wire new_net_3212;
	wire new_net_8389;
	wire new_net_19464;
	wire new_net_20287;
	wire new_net_2263;
	wire new_net_20;
	wire new_net_2243;
	wire new_net_4143;
	wire new_net_10500;
	wire new_net_940;
	wire _1720_;
	wire new_net_2687;
	wire new_net_2377;
	wire new_net_13009;
	wire new_net_15682;
	wire new_net_2259;
	wire new_net_3736;
	wire new_net_7294;
	wire new_net_20068;
	wire new_net_20970;
	wire new_net_21283;
	wire new_net_21295;
	wire new_net_16735;
	wire _1721_;
	wire new_net_11153;
	wire new_net_3503;
	wire new_net_13533;
	wire new_net_14626;
	wire new_net_9285;
	wire new_net_15675;
	wire new_net_319;
	wire new_net_8775;
	wire new_net_19463;
	wire new_net_19864;
	wire new_net_20003;
	wire new_net_13397;
	wire new_net_15728;
	wire new_net_18401;
	wire new_net_13376;
	wire new_net_16699;
	wire new_net_9281;
	wire new_net_11746;
	wire new_net_4653;
	wire new_net_15681;
	wire new_net_16154;
	wire new_net_17823;
	wire new_net_2370;
	wire _1722_;
	wire new_net_13726;
	wire new_net_2367;
	wire new_net_3053;
	wire new_net_7223;
	wire new_net_12977;
	wire new_net_12545;
	wire new_net_7292;
	wire new_net_20288;
	wire new_net_21347;
	wire new_net_18719;
	wire _1309_;
	wire new_net_2371;
	wire _1723_;
	wire new_net_10505;
	wire new_net_7295;
	wire new_net_20065;
	wire new_net_5022;
	wire new_net_2372;
	wire new_net_4478;
	wire new_net_12544;
	wire new_net_19311;
	wire new_net_2235;
	wire _1724_;
	wire new_net_2268;
	wire new_net_4138;
	wire new_net_20971;
	wire new_net_21284;
	wire new_net_2244;
	wire new_net_315;
	wire new_net_3613;
	wire new_net_3731;
	wire new_net_11154;
	wire new_net_4094;
	wire new_net_20848;
	wire new_net_14645;
	wire new_net_4475;
	wire _1725_;
	wire new_net_4135;
	wire new_net_19308;
	wire new_net_19865;
	wire new_net_20004;
	wire new_net_17838;
	wire new_net_18804;
	wire new_net_13377;
	wire new_net_16700;
	wire new_net_11747;
	wire new_net_16155;
	wire new_net_17824;
	wire new_net_5481;
	wire new_net_17126;
	wire new_net_17622;
	wire new_net_12597;
	wire new_net_21042;
	wire new_net_10371;
	wire new_net_16272;
	wire new_net_13964;
	wire new_net_2237;
	wire _1726_;
	wire new_net_20289;
	wire new_net_7045;
	wire new_net_15680;
	wire new_net_2238;
	wire new_net_4060;
	wire new_net_5478;
	wire new_net_664;
	wire new_net_10507;
	wire new_net_8774;
	wire new_net_2239;
	wire _1727_;
	wire new_net_3209;
	wire new_net_4477;
	wire new_net_4668;
	wire new_net_7427;
	wire new_net_20972;
	wire new_net_21285;
	wire new_net_3200;
	wire new_net_3045;
	wire _1728_;
	wire new_net_8637;
	wire new_net_11155;
	wire new_net_12543;
	wire new_net_7298;
	wire new_net_13299;
	wire new_net_15677;
	wire new_net_7297;
	wire new_net_20005;
	wire new_net_20329;
	wire _0021_;
	wire new_net_17825;
	wire new_net_13378;
	wire new_net_16701;
	wire new_net_9279;
	wire new_net_11748;
	wire new_net_16156;
	wire _1729_;
	wire new_net_17127;
	wire new_net_17623;
	wire new_net_8388;
	wire new_net_5997;
	wire new_net_8390;
	wire new_net_2379;
	wire new_net_3871;
	wire new_net_20290;
	wire new_net_8385;
	wire _1730_;
	wire new_net_4470;
	wire new_net_7047;
	wire new_net_10504;
	wire new_net_20331;
	wire new_net_19964;
	wire new_net_7299;
	wire new_net_3608;
	wire new_net_10054;
	wire _1731_;
	wire new_net_2265;
	wire new_net_2685;
	wire new_net_4603;
	wire new_net_20067;
	wire new_net_20330;
	wire new_net_20973;
	wire new_net_9282;
	wire new_net_2267;
	wire new_net_2688;
	wire new_net_3869;
	wire new_net_5479;
	wire new_net_8639;
	wire new_net_11156;
	wire new_net_7226;
	wire new_net_18811;
	wire _1732_;
	wire new_net_23;
	wire new_net_2270;
	wire new_net_2374;
	wire new_net_19462;
	wire new_net_20006;
	wire new_net_18906;
	wire new_net_12599;
	wire new_net_16702;
	wire new_net_11749;
	wire new_net_16157;
	wire new_net_17826;
	wire new_net_26;
	wire new_net_8776;
	wire new_net_17128;
	wire new_net_17624;
	wire new_net_12542;
	wire new_net_17845;
	wire new_net_13765;
	wire new_net_6000;
	wire new_net_13379;
	wire new_net_4651;
	wire _1733_;
	wire new_net_5042;
	wire new_net_7230;
	wire new_net_8392;
	wire new_net_20291;
	wire new_net_18529;
	wire new_net_19165;
	wire new_net_7062;
	wire new_net_7296;
	wire new_net_6002;
	wire new_net_9286;
	wire new_net_2240;
	wire new_net_2376;
	wire new_net_4652;
	wire new_net_4671;
	wire new_net_15026;
	wire new_net_7293;
	wire new_net_9284;
	wire new_net_15679;
	wire _1734_;
	wire new_net_323;
	wire new_net_2375;
	wire new_net_4474;
	wire new_net_7426;
	wire new_net_20064;
	wire new_net_2686;
	wire new_net_7432;
	wire new_net_8384;
	wire new_net_20974;
	wire new_net_21287;
	wire new_net_16644;
	wire new_net_5328;
	wire _1735_;
	wire new_net_3054;
	wire new_net_2683;
	wire new_net_3205;
	wire new_net_11157;
	wire new_net_4604;
	wire new_net_7227;
	wire new_net_20066;
	wire new_net_2316;
	wire new_net_11792;
	wire new_net_15770;
	wire _1316_;
	wire new_net_18277;
	wire new_net_16168;
	wire new_net_12493;
	wire new_net_3470;
	wire new_net_10128;
	wire new_net_3974;
	wire new_net_12495;
	wire new_net_13015;
	wire new_net_13167;
	wire new_net_12683;
	wire new_net_16974;
	wire _1442_;
	wire new_net_12446;
	wire new_net_13839;
	wire new_net_17377;
	wire new_net_21041;
	wire new_net_4386;
	wire new_net_19599;
	wire new_net_4834;
	wire new_net_18234;
	wire new_net_4726;
	wire _1443_;
	wire new_net_956;
	wire new_net_17666;
	wire new_net_5011;
	wire new_net_19483;
	wire new_net_9231;
	wire new_net_858;
	wire new_net_4720;
	wire new_net_4935;
	wire new_net_13023;
	wire new_net_16736;
	wire new_net_9647;
	wire _1444_;
	wire new_net_856;
	wire new_net_962;
	wire new_net_13534;
	wire new_net_14627;
	wire new_net_8253;
	wire new_net_12494;
	wire new_net_16503;
	wire new_net_4722;
	wire new_net_4934;
	wire new_net_11205;
	wire new_net_15390;
	wire new_net_12001;
	wire new_net_13571;
	wire new_net_14553;
	wire new_net_577;
	wire new_net_13398;
	wire new_net_15729;
	wire new_net_18402;
	wire _0840_;
	wire new_net_5922;
	wire _1445_;
	wire new_net_5018;
	wire new_net_17225;
	wire new_net_13727;
	wire new_net_12325;
	wire new_net_12978;
	wire new_net_16361;
	wire new_net_13016;
	wire new_net_13168;
	wire new_net_12684;
	wire new_net_16975;
	wire new_net_1558;
	wire new_net_2568;
	wire new_net_4938;
	wire new_net_5012;
	wire new_net_9233;
	wire new_net_18720;
	wire new_net_3475;
	wire new_net_8246;
	wire _1446_;
	wire new_net_1550;
	wire new_net_8139;
	wire new_net_5017;
	wire new_net_20137;
	wire new_net_9107;
	wire new_net_961;
	wire new_net_17224;
	wire new_net_19484;
	wire new_net_19608;
	wire new_net_17472;
	wire new_net_11925;
	wire new_net_16631;
	wire _1447_;
	wire new_net_2577;
	wire new_net_9479;
	wire new_net_1078;
	wire new_net_5920;
	wire new_net_19609;
	wire new_net_20872;
	wire new_net_20849;
	wire new_net_12030;
	wire new_net_14646;
	wire new_net_4724;
	wire new_net_3257;
	wire new_net_6654;
	wire _1448_;
	wire new_net_6187;
	wire new_net_3083;
	wire new_net_11206;
	wire new_net_12078;
	wire new_net_4747;
	wire new_net_18805;
	wire new_net_9398;
	wire new_net_9110;
	wire new_net_1713;
	wire new_net_2574;
	wire new_net_6196;
	wire new_net_8144;
	wire new_net_8660;
	wire new_net_16141;
	wire new_net_13965;
	wire new_net_16273;
	wire new_net_9395;
	wire new_net_16362;
	wire new_net_17227;
	wire new_net_9232;
	wire new_net_13017;
	wire new_net_13169;
	wire new_net_5919;
	wire new_net_12685;
	wire new_net_16504;
	wire new_net_16976;
	wire new_net_15413;
	wire new_net_20138;
	wire new_net_14318;
	wire new_net_2709;
	wire new_net_9393;
	wire new_net_16630;
	wire new_net_3256;
	wire _1450_;
	wire new_net_8140;
	wire new_net_2571;
	wire new_net_4940;
	wire new_net_3086;
	wire new_net_19485;
	wire new_net_8131;
	wire new_net_1721;
	wire new_net_8143;
	wire new_net_7385;
	wire new_net_9109;
	wire new_net_9652;
	wire _1451_;
	wire new_net_1716;
	wire new_net_8146;
	wire new_net_9230;
	wire new_net_10126;
	wire new_net_786;
	wire new_net_16629;
	wire new_net_8127;
	wire new_net_964;
	wire new_net_2995;
	wire new_net_1548;
	wire new_net_3091;
	wire new_net_4939;
	wire new_net_11207;
	wire new_net_18409;
	wire new_net_9394;
	wire new_net_6659;
	wire new_net_8653;
	wire new_net_2575;
	wire _1452_;
	wire new_net_5016;
	wire new_net_5375;
	wire new_net_15386;
	wire new_net_15536;
	wire new_net_16363;
	wire new_net_13018;
	wire new_net_16977;
	wire new_net_6658;
	wire new_net_8729;
	wire new_net_13170;
	wire new_net_8132;
	wire new_net_12686;
	wire new_net_8456;
	wire new_net_15943;
	wire new_net_12496;
	wire new_net_2572;
	wire new_net_2988;
	wire _1453_;
	wire new_net_20139;
	wire new_net_16790;
	wire new_net_4388;
	wire new_net_8129;
	wire new_net_8252;
	wire new_net_3261;
	wire new_net_7085;
	wire new_net_8125;
	wire _1454_;
	wire new_net_855;
	wire new_net_7083;
	wire new_net_5559;
	wire new_net_7986;
	wire new_net_18812;
	wire new_net_11208;
	wire new_net_4390;
	wire new_net_8732;
	wire new_net_957;
	wire _1455_;
	wire new_net_1553;
	wire new_net_6193;
	wire new_net_18907;
	wire new_net_3214;
	wire new_net_13658;
	wire new_net_9103;
	wire new_net_1557;
	wire new_net_2986;
	wire new_net_4723;
	wire new_net_10132;
	wire new_net_19607;
	wire new_net_17846;
	wire new_net_18941;
	wire new_net_15385;
	wire new_net_15537;
	wire new_net_16506;
	wire new_net_13019;
	wire new_net_13171;
	wire new_net_16978;
	wire _1456_;
	wire new_net_860;
	wire new_net_12687;
	wire new_net_17231;
	wire new_net_18530;
	wire new_net_8466;
	wire new_net_10127;
	wire new_net_854;
	wire new_net_960;
	wire new_net_12497;
	wire new_net_20140;
	wire new_net_15027;
	wire new_net_3368;
	wire new_net_4721;
	wire new_net_1717;
	wire new_net_1546;
	wire _1457_;
	wire new_net_6192;
	wire new_net_13027;
	wire new_net_21165;
	wire _1813_;
	wire new_net_8726;
	wire new_net_1545;
	wire new_net_8130;
	wire new_net_13097;
	wire new_net_16645;
	wire new_net_8251;
	wire new_net_2578;
	wire new_net_2994;
	wire _1458_;
	wire new_net_11687;
	wire new_net_16570;
	wire new_net_11209;
	wire new_net_8248;
	wire new_net_4385;
	wire new_net_966;
	wire new_net_2993;
	wire new_net_3259;
	wire new_net_8652;
	wire new_net_11793;
	wire new_net_20362;
	wire new_net_6991;
	wire new_net_12766;
	wire new_net_13450;
	wire new_net_18278;
	wire new_net_17229;
	wire new_net_16624;
	wire new_net_1714;
	wire new_net_2992;
	wire _1459_;
	wire new_net_8142;
	wire new_net_19600;
	wire new_net_15200;
	wire new_net_16169;
	wire new_net_15384;
	wire new_net_16365;
	wire new_net_9655;
	wire new_net_13020;
	wire new_net_13172;
	wire new_net_16507;
	wire new_net_3362;
	wire new_net_3476;
	wire new_net_6660;
	wire new_net_8128;
	wire new_net_3085;
	wire new_net_16623;
	wire new_net_3252;
	wire new_net_6655;
	wire new_net_8727;
	wire new_net_958;
	wire _1460_;
	wire new_net_19606;
	wire new_net_20141;
	wire new_net_7245;
	wire new_net_14984;
	wire new_net_5373;
	wire new_net_9229;
	wire new_net_12499;
	wire new_net_959;
	wire new_net_14123;
	wire new_net_3084;
	wire new_net_17228;
	wire new_net_8730;
	wire _1461_;
	wire new_net_859;
	wire new_net_6185;
	wire new_net_13024;
	wire new_net_16737;
	wire new_net_5925;
	wire new_net_7082;
	wire new_net_8141;
	wire new_net_13535;
	wire new_net_14628;
	wire new_net_9653;
	wire new_net_8250;
	wire _1462_;
	wire new_net_1719;
	wire new_net_849;
	wire new_net_3260;
	wire new_net_11210;
	wire new_net_20363;
	wire new_net_12002;
	wire new_net_13572;
	wire new_net_14552;
	wire new_net_13399;
	wire new_net_15730;
	wire new_net_18403;
	wire new_net_12500;
	wire new_net_17230;
	wire new_net_8725;
	wire new_net_2990;
	wire new_net_5013;
	wire new_net_5560;
	wire new_net_17294;
	wire new_net_13728;
	wire new_net_12326;
	wire new_net_16980;
	wire new_net_3088;
	wire new_net_17233;
	wire new_net_17726;
	wire new_net_12689;
	wire new_net_16366;
	wire new_net_9399;
	wire new_net_13021;
	wire new_net_16897;
	wire new_net_13845;
	wire new_net_12979;
	wire new_net_18968;
	wire new_net_18721;
	wire new_net_9046;
	wire new_net_2573;
	wire new_net_3472;
	wire new_net_4719;
	wire new_net_19605;
	wire new_net_20142;
	wire new_net_10427;
	wire new_net_3348;
	wire new_net_9104;
	wire new_net_12498;
	wire new_net_4389;
	wire _1464_;
	wire new_net_8650;
	wire new_net_17473;
	wire new_net_11926;
	wire new_net_1551;
	wire new_net_1718;
	wire new_net_2991;
	wire new_net_3081;
	wire new_net_7985;
	wire new_net_8657;
	wire new_net_3366;
	wire new_net_9650;
	wire _1465_;
	wire new_net_5916;
	wire new_net_10125;
	wire new_net_19604;
	wire new_net_16530;
	wire new_net_20873;
	wire new_net_20850;
	wire new_net_14647;
	wire new_net_12031;
	wire new_net_11211;
	wire new_net_16627;
	wire new_net_963;
	wire new_net_6657;
	wire new_net_8655;
	wire new_net_17383;
	wire new_net_20364;
	wire new_net_4748;
	wire new_net_18806;
	wire new_net_8254;
	wire new_net_4725;
	wire new_net_12501;
	wire new_net_16621;
	wire _1466_;
	wire new_net_1547;
	wire new_net_4391;
	wire new_net_10387;
	wire new_net_16142;
	wire new_net_17727;
	wire new_net_15540;
	wire new_net_16898;
	wire new_net_17232;
	wire new_net_16367;
	wire new_net_13022;
	wire new_net_16628;
	wire new_net_13966;
	wire new_net_2987;
	wire new_net_3471;
	wire new_net_14850;
	wire new_net_9402;
	wire _1467_;
	wire new_net_861;
	wire new_net_2570;
	wire new_net_20143;
	wire new_net_1544;
	wire new_net_3255;
	wire new_net_5921;
	wire new_net_19603;
	wire new_net_14319;
	wire _1468_;
	wire new_net_3254;
	wire new_net_2569;
	wire new_net_10129;
	wire new_net_1552;
	wire new_net_3087;
	wire new_net_5015;
	wire new_net_10131;
	wire new_net_19486;
	wire new_net_5956;
	wire new_net_5014;
	wire new_net_5374;
	wire new_net_11212;
	wire new_net_3970;
	wire _1469_;
	wire new_net_8126;
	wire new_net_20365;
	wire new_net_13711;
	wire new_net_8651;
	wire new_net_9397;
	wire new_net_12502;
	wire new_net_2989;
	wire new_net_3351;
	wire new_net_12454;
	wire new_net_13847;
	wire new_net_17384;
	wire new_net_9041;
	wire new_net_16510;
	wire new_net_5019;
	wire new_net_15382;
	wire new_net_17728;
	wire new_net_9400;
	wire new_net_16368;
	wire new_net_15383;
	wire new_net_7084;
	wire new_net_20144;
	wire new_net_15944;
	wire new_net_16791;
	wire new_net_10123;
	wire new_net_3092;
	wire new_net_9108;
	wire _1471_;
	wire new_net_5918;
	wire new_net_6195;
	wire new_net_4936;
	wire new_net_9044;
	wire new_net_3473;
	wire new_net_9396;
	wire new_net_3972;
	wire new_net_1711;
	wire new_net_965;
	wire new_net_3080;
	wire new_net_5923;
	wire new_net_9043;
	wire _1472_;
	wire new_net_6662;
	wire new_net_19487;
	wire new_net_14539;
	wire new_net_18813;
	wire new_net_8658;
	wire new_net_11213;
	wire new_net_9105;
	wire new_net_5917;
	wire new_net_7984;
	wire new_net_8138;
	wire new_net_8245;
	wire new_net_8728;
	wire new_net_20366;
	wire new_net_18908;
	wire new_net_13659;
	wire new_net_9102;
	wire new_net_12503;
	wire _1473_;
	wire new_net_17847;
	wire new_net_2471;
	wire new_net_7987;
	wire new_net_10124;
	wire new_net_12455;
	wire new_net_13848;
	wire new_net_17385;
	wire new_net_17729;
	wire new_net_15381;
	wire new_net_15542;
	wire new_net_16900;
	wire new_net_16369;
	wire new_net_7060;
	wire new_net_8124;
	wire _1474_;
	wire new_net_20145;
	wire new_net_15028;
	wire new_net_8649;
	wire new_net_9106;
	wire new_net_9651;
	wire new_net_850;
	wire new_net_18064;
	wire new_net_13028;
	wire _1475_;
	wire new_net_3262;
	wire new_net_21166;
	wire new_net_13098;
	wire new_net_16646;
	wire new_net_4933;
	wire new_net_1555;
	wire new_net_3253;
	wire new_net_19488;
	wire new_net_16571;
	wire new_net_10130;
	wire new_net_11214;
	wire new_net_17234;
	wire _1476_;
	wire new_net_20367;
	wire new_net_11794;
	wire new_net_12767;
	wire new_net_13451;
	wire new_net_9657;
	wire new_net_1556;
	wire new_net_5376;
	wire _1323_;
	wire new_net_15772;
	wire new_net_18279;
	wire new_net_12456;
	wire new_net_13849;
	wire new_net_17386;
	wire new_net_17730;
	wire new_net_15380;
	wire new_net_15543;
	wire new_net_16901;
	wire new_net_16370;
	wire new_net_1715;
	wire new_net_2567;
	wire new_net_1226;
	wire new_net_21043;
	wire new_net_7988;
	wire new_net_853;
	wire new_net_20146;
	wire new_net_14985;
	wire new_net_8145;
	wire new_net_3350;
	wire new_net_9042;
	wire new_net_8249;
	wire _1478_;
	wire new_net_4718;
	wire new_net_9654;
	wire new_net_11836;
	wire new_net_8247;
	wire new_net_3477;
	wire new_net_4717;
	wire new_net_7983;
	wire new_net_13012;
	wire new_net_13025;
	wire new_net_8654;
	wire _1479_;
	wire new_net_1549;
	wire new_net_1710;
	wire new_net_9656;
	wire new_net_16626;
	wire new_net_19489;
	wire new_net_19601;
	wire new_net_16738;
	wire new_net_6190;
	wire new_net_11215;
	wire new_net_3090;
	wire new_net_4937;
	wire new_net_9648;
	wire new_net_14629;
	wire new_net_13536;
	wire new_net_20368;
	wire new_net_12003;
	wire new_net_13573;
	wire new_net_14551;
	wire new_net_8023;
	wire new_net_13400;
	wire new_net_15731;
	wire new_net_18404;
	wire new_net_17235;
	wire new_net_9401;
	wire _1480_;
	wire new_net_1560;
	wire new_net_5924;
	wire new_net_19602;
	wire new_net_17027;
	wire _0847_;
	wire new_net_13729;
	wire new_net_12327;
	wire new_net_12457;
	wire new_net_13850;
	wire new_net_17387;
	wire new_net_17731;
	wire new_net_15544;
	wire new_net_16902;
	wire new_net_16371;
	wire new_net_2576;
	wire new_net_3263;
	wire new_net_13026;
	wire new_net_18722;
	wire new_net_3089;
	wire _1481_;
	wire new_net_16622;
	wire new_net_6656;
	wire new_net_20147;
	wire new_net_6973;
	wire new_net_857;
	wire new_net_6661;
	wire new_net_17532;
	wire new_net_21390;
	wire new_net_17474;
	wire new_net_1712;
	wire _1482_;
	wire new_net_851;
	wire new_net_1559;
	wire new_net_12504;
	wire new_net_2816;
	wire new_net_6189;
	wire new_net_4932;
	wire new_net_8656;
	wire new_net_1077;
	wire new_net_3474;
	wire new_net_19490;
	wire new_net_20874;
	wire new_net_6194;
	wire new_net_11216;
	wire new_net_8244;
	wire _1483_;
	wire new_net_9649;
	wire new_net_20369;
	wire new_net_20851;
	wire new_net_12032;
	wire new_net_14648;
	wire new_net_19751;
	wire new_net_16143;
	wire new_net_12932;
	wire new_net_16275;
	wire new_net_13967;
	wire new_net_1751;
	wire new_net_4524;
	wire new_net_19759;
	wire new_net_19947;
	wire new_net_20523;
	wire new_net_21249;
	wire new_net_14851;
	wire new_net_16277;
	wire new_net_17010;
	wire new_net_9929;
	wire new_net_13827;
	wire new_net_16846;
	wire _0812_;
	wire new_net_4844;
	wire new_net_10728;
	wire new_net_13251;
	wire new_net_16597;
	wire new_net_8064;
	wire new_net_1013;
	wire new_net_4556;
	wire new_net_4846;
	wire new_net_19807;
	wire new_net_21250;
	wire new_net_14062;
	wire _0813_;
	wire new_net_4578;
	wire new_net_10510;
	wire new_net_11714;
	wire new_net_9827;
	wire new_net_7070;
	wire new_net_868;
	wire new_net_1750;
	wire new_net_1469;
	wire new_net_4523;
	wire new_net_7061;
	wire new_net_15643;
	wire new_net_5215;
	wire new_net_1145;
	wire new_net_1467;
	wire _0814_;
	wire new_net_4697;
	wire new_net_14557;
	wire new_net_4848;
	wire new_net_20076;
	wire new_net_13712;
	wire new_net_12102;
	wire new_net_17141;
	wire new_net_4522;
	wire new_net_4581;
	wire new_net_18654;
	wire new_net_20408;
	wire new_net_3251;
	wire new_net_15639;
	wire _0815_;
	wire new_net_1753;
	wire new_net_10722;
	wire new_net_19948;
	wire new_net_18464;
	wire new_net_15945;
	wire new_net_11712;
	wire new_net_12100;
	wire new_net_13498;
	wire new_net_16492;
	wire new_net_16278;
	wire new_net_17011;
	wire new_net_13828;
	wire new_net_8066;
	wire new_net_9831;
	wire new_net_4842;
	wire new_net_16792;
	wire new_net_5554;
	wire _0816_;
	wire new_net_865;
	wire new_net_14426;
	wire new_net_18644;
	wire new_net_19770;
	wire new_net_19808;
	wire new_net_15650;
	wire new_net_14427;
	wire new_net_20514;
	wire new_net_9826;
	wire new_net_3122;
	wire new_net_4843;
	wire _0817_;
	wire new_net_4727;
	wire new_net_14098;
	wire new_net_14540;
	wire new_net_18814;
	wire new_net_8070;
	wire new_net_1142;
	wire new_net_3117;
	wire new_net_8333;
	wire new_net_20077;
	wire new_net_16959;
	wire new_net_18909;
	wire new_net_13660;
	wire new_net_8069;
	wire _0818_;
	wire new_net_4085;
	wire new_net_20409;
	wire new_net_6946;
	wire new_net_20423;
	wire new_net_17848;
	wire new_net_2470;
	wire new_net_13768;
	wire new_net_19785;
	wire new_net_9970;
	wire new_net_1148;
	wire new_net_4701;
	wire new_net_19949;
	wire new_net_14368;
	wire new_net_15062;
	wire new_net_11711;
	wire new_net_12099;
	wire new_net_13499;
	wire new_net_16493;
	wire new_net_16279;
	wire new_net_17012;
	wire new_net_9971;
	wire new_net_13829;
	wire new_net_17142;
	wire new_net_1472;
	wire new_net_15029;
	wire new_net_14909;
	wire new_net_18159;
	wire new_net_9969;
	wire new_net_3121;
	wire new_net_4703;
	wire new_net_7075;
	wire new_net_19809;
	wire new_net_18065;
	wire new_net_6008;
	wire new_net_13029;
	wire new_net_21167;
	wire _0820_;
	wire new_net_869;
	wire new_net_4589;
	wire new_net_10515;
	wire new_net_14428;
	wire new_net_18653;
	wire new_net_19769;
	wire new_net_13099;
	wire new_net_16647;
	wire new_net_4765;
	wire new_net_16356;
	wire new_net_7791;
	wire new_net_20522;
	wire new_net_647;
	wire new_net_11689;
	wire new_net_16572;
	wire new_net_9926;
	wire _0821_;
	wire new_net_8337;
	wire new_net_1006;
	wire new_net_20078;
	wire new_net_12768;
	wire new_net_13452;
	wire new_net_20410;
	wire new_net_15773;
	wire new_net_18280;
	wire new_net_20717;
	wire _0822_;
	wire new_net_10513;
	wire new_net_19950;
	wire new_net_20512;
	wire new_net_21044;
	wire new_net_10727;
	wire new_net_16600;
	wire new_net_16706;
	wire new_net_11710;
	wire new_net_13500;
	wire new_net_16494;
	wire new_net_16280;
	wire new_net_17013;
	wire new_net_13830;
	wire new_net_17143;
	wire new_net_14986;
	wire new_net_5218;
	wire _0823_;
	wire new_net_3124;
	wire new_net_4529;
	wire new_net_8334;
	wire new_net_19810;
	wire new_net_14125;
	wire new_net_13013;
	wire new_net_14429;
	wire new_net_8068;
	wire new_net_6763;
	wire new_net_2443;
	wire new_net_19768;
	wire new_net_20452;
	wire new_net_16625;
	wire new_net_12631;
	wire new_net_14081;
	wire new_net_1756;
	wire _0824_;
	wire new_net_4702;
	wire new_net_8293;
	wire new_net_13537;
	wire new_net_14630;
	wire new_net_1139;
	wire new_net_18652;
	wire new_net_19333;
	wire new_net_20079;
	wire new_net_12004;
	wire new_net_13574;
	wire new_net_14550;
	wire new_net_13401;
	wire new_net_15732;
	wire new_net_18405;
	wire new_net_10731;
	wire new_net_13254;
	wire new_net_7793;
	wire new_net_9973;
	wire new_net_727;
	wire new_net_872;
	wire _0825_;
	wire new_net_4588;
	wire new_net_4699;
	wire new_net_19767;
	wire new_net_17296;
	wire new_net_13730;
	wire new_net_1749;
	wire new_net_1005;
	wire new_net_4554;
	wire new_net_19951;
	wire new_net_8099;
	wire new_net_18723;
	wire new_net_16601;
	wire new_net_16707;
	wire new_net_11709;
	wire new_net_13501;
	wire new_net_16495;
	wire new_net_16281;
	wire new_net_17014;
	wire new_net_9966;
	wire new_net_13831;
	wire _0826_;
	wire new_net_7783;
	wire new_net_9967;
	wire new_net_10517;
	wire new_net_19811;
	wire new_net_17533;
	wire new_net_17475;
	wire new_net_10723;
	wire new_net_14430;
	wire new_net_8600;
	wire new_net_5219;
	wire _0827_;
	wire new_net_2448;
	wire new_net_10509;
	wire new_net_16751;
	wire new_net_18029;
	wire new_net_21080;
	wire new_net_10729;
	wire new_net_15649;
	wire new_net_7789;
	wire new_net_9924;
	wire new_net_1003;
	wire new_net_5221;
	wire new_net_19766;
	wire new_net_11730;
	wire new_net_16532;
	wire new_net_20875;
	wire new_net_7785;
	wire new_net_8062;
	wire _0828_;
	wire new_net_1144;
	wire new_net_1471;
	wire new_net_3118;
	wire new_net_4528;
	wire new_net_18651;
	wire new_net_19332;
	wire new_net_20080;
	wire new_net_9972;
	wire new_net_4558;
	wire new_net_20412;
	wire new_net_20520;
	wire new_net_12328;
	wire new_net_18325;
	wire new_net_16144;
	wire new_net_4435;
	wire new_net_15648;
	wire new_net_9921;
	wire _0829_;
	wire new_net_10512;
	wire new_net_19952;
	wire new_net_13968;
	wire new_net_16276;
	wire new_net_13255;
	wire new_net_16602;
	wire new_net_16708;
	wire new_net_11708;
	wire new_net_12097;
	wire new_net_13502;
	wire new_net_16282;
	wire new_net_17015;
	wire new_net_13832;
	wire new_net_16496;
	wire new_net_14852;
	wire new_net_12098;
	wire _0830_;
	wire new_net_19812;
	wire new_net_20519;
	wire new_net_16879;
	wire new_net_14321;
	wire new_net_14063;
	wire new_net_14431;
	wire new_net_8063;
	wire new_net_1007;
	wire new_net_10724;
	wire _0831_;
	wire new_net_4583;
	wire new_net_6764;
	wire new_net_3283;
	wire new_net_8003;
	wire new_net_8596;
	wire new_net_2441;
	wire new_net_1009;
	wire new_net_4557;
	wire new_net_20081;
	wire new_net_14558;
	wire _0035_;
	wire new_net_13713;
	wire _0832_;
	wire new_net_18649;
	wire new_net_20413;
	wire new_net_13879;
	wire new_net_9928;
	wire new_net_2445;
	wire new_net_1012;
	wire new_net_19953;
	wire new_net_20518;
	wire new_net_18513;
	wire new_net_4696;
	wire new_net_13256;
	wire new_net_16603;
	wire new_net_16709;
	wire new_net_11707;
	wire new_net_12096;
	wire new_net_13503;
	wire new_net_16497;
	wire new_net_16283;
	wire new_net_17016;
	wire new_net_15946;
	wire new_net_16793;
	wire new_net_15647;
	wire new_net_19813;
	wire new_net_4585;
	wire new_net_14432;
	wire new_net_5222;
	wire _0834_;
	wire new_net_3125;
	wire new_net_17507;
	wire new_net_19331;
	wire new_net_8339;
	wire new_net_9927;
	wire new_net_3114;
	wire new_net_14541;
	wire new_net_18815;
	wire new_net_10135;
	wire _0835_;
	wire new_net_5214;
	wire new_net_6766;
	wire new_net_7072;
	wire new_net_20082;
	wire new_net_11777;
	wire new_net_18910;
	wire new_net_3216;
	wire new_net_15640;
	wire new_net_8598;
	wire new_net_9823;
	wire new_net_1001;
	wire new_net_4580;
	wire new_net_20414;
	wire new_net_17849;
	wire new_net_4549;
	wire new_net_1138;
	wire new_net_1470;
	wire _0836_;
	wire new_net_730;
	wire new_net_19954;
	wire new_net_18532;
	wire new_net_16498;
	wire new_net_13257;
	wire new_net_16604;
	wire new_net_11706;
	wire new_net_16284;
	wire new_net_17017;
	wire new_net_13834;
	wire new_net_1464;
	wire new_net_4579;
	wire new_net_13504;
	wire new_net_15899;
	wire new_net_15030;
	wire new_net_14910;
	wire _0837_;
	wire new_net_18160;
	wire new_net_19814;
	wire new_net_725;
	wire new_net_18066;
	wire new_net_14433;
	wire new_net_8336;
	wire new_net_9925;
	wire new_net_21168;
	wire new_net_13100;
	wire new_net_8335;
	wire new_net_9830;
	wire new_net_2450;
	wire _0838_;
	wire new_net_4526;
	wire new_net_19670;
	wire new_net_19765;
	wire new_net_11690;
	wire new_net_16573;
	wire new_net_15645;
	wire new_net_8601;
	wire new_net_20083;
	wire new_net_12769;
	wire new_net_13453;
	wire new_net_4698;
	wire new_net_7792;
	wire _0839_;
	wire new_net_726;
	wire new_net_5114;
	wire new_net_14997;
	wire new_net_16853;
	wire new_net_19760;
	wire new_net_20415;
	wire _1330_;
	wire new_net_15774;
	wire new_net_18281;
	wire new_net_728;
	wire new_net_863;
	wire new_net_19955;
	wire new_net_4536;
	wire new_net_7073;
	wire new_net_4586;
	wire new_net_13258;
	wire new_net_16605;
	wire new_net_16711;
	wire new_net_11705;
	wire new_net_12094;
	wire new_net_13505;
	wire new_net_16499;
	wire new_net_16285;
	wire new_net_14987;
	wire new_net_7782;
	wire new_net_1468;
	wire new_net_4527;
	wire new_net_4584;
	wire new_net_8071;
	wire new_net_19815;
	wire new_net_14126;
	wire new_net_10518;
	wire new_net_14434;
	wire new_net_15646;
	wire new_net_1002;
	wire _0841_;
	wire new_net_3116;
	wire new_net_11838;
	wire new_net_9828;
	wire new_net_19330;
	wire new_net_8751;
	wire new_net_21235;
	wire new_net_10725;
	wire new_net_1755;
	wire new_net_1011;
	wire new_net_3123;
	wire new_net_4587;
	wire new_net_12632;
	wire new_net_14082;
	wire new_net_8625;
	wire new_net_9974;
	wire _0842_;
	wire new_net_2442;
	wire new_net_4850;
	wire new_net_6765;
	wire new_net_20084;
	wire new_net_13538;
	wire new_net_12005;
	wire new_net_13575;
	wire new_net_13402;
	wire new_net_15733;
	wire new_net_18406;
	wire new_net_1147;
	wire new_net_1474;
	wire new_net_2449;
	wire new_net_9829;
	wire new_net_10133;
	wire new_net_18648;
	wire new_net_19764;
	wire new_net_20416;
	wire new_net_17297;
	wire new_net_13731;
	wire new_net_4530;
	wire new_net_2444;
	wire _0843_;
	wire new_net_8067;
	wire new_net_19956;
	wire new_net_20517;
	wire new_net_21251;
	wire new_net_18724;
	wire new_net_16606;
	wire new_net_16286;
	wire new_net_7071;
	wire new_net_10508;
	wire new_net_13506;
	wire new_net_13259;
	wire new_net_16500;
	wire new_net_11704;
	wire new_net_12093;
	wire new_net_16712;
	wire new_net_6978;
	wire new_net_7077;
	wire new_net_8330;
	wire new_net_8602;
	wire _0844_;
	wire new_net_19816;
	wire new_net_17534;
	wire new_net_17476;
	wire new_net_8338;
	wire new_net_10511;
	wire new_net_14435;
	wire new_net_3377;
	wire new_net_10603;
	wire new_net_16752;
	wire new_net_7076;
	wire new_net_8563;
	wire new_net_9923;
	wire new_net_1475;
	wire _0845_;
	wire new_net_3119;
	wire new_net_18030;
	wire new_net_19762;
	wire new_net_1073;
	wire new_net_16533;
	wire new_net_20876;
	wire new_net_10516;
	wire new_net_15644;
	wire new_net_8566;
	wire new_net_8595;
	wire new_net_873;
	wire new_net_5220;
	wire new_net_20085;
	wire new_net_5670;
	wire _0846_;
	wire new_net_9824;
	wire new_net_19763;
	wire new_net_20417;
	wire _0686_;
	wire new_net_12329;
	wire new_net_18326;
	wire new_net_16145;
	wire new_net_4847;
	wire new_net_1752;
	wire new_net_1141;
	wire new_net_9968;
	wire new_net_19957;
	wire new_net_12934;
	wire new_net_7692;
	wire new_net_16855;
	wire new_net_13260;
	wire new_net_16607;
	wire new_net_16713;
	wire new_net_11703;
	wire new_net_12092;
	wire new_net_13507;
	wire new_net_15641;
	wire new_net_16501;
	wire new_net_16287;
	wire new_net_9623;
	wire new_net_16927;
	wire new_net_4841;
	wire new_net_4849;
	wire new_net_8565;
	wire new_net_1010;
	wire new_net_4525;
	wire new_net_4700;
	wire new_net_7788;
	wire new_net_19817;
	wire new_net_20516;
	wire new_net_16880;
	wire new_net_14064;
	wire new_net_10730;
	wire new_net_10136;
	wire new_net_7790;
	wire new_net_1008;
	wire _0848_;
	wire new_net_14436;
	wire new_net_7389;
	wire new_net_1463;
	wire new_net_8065;
	wire new_net_8599;
	wire new_net_14661;
	wire new_net_18913;
	wire new_net_9060;
	wire new_net_4582;
	wire new_net_4555;
	wire new_net_1149;
	wire _0849_;
	wire new_net_13303;
	wire new_net_18643;
	wire new_net_20086;
	wire new_net_14559;
	wire new_net_8564;
	wire new_net_1004;
	wire new_net_5217;
	wire new_net_20418;
	wire new_net_13714;
	wire new_net_8331;
	wire new_net_1466;
	wire new_net_866;
	wire _0850_;
	wire new_net_4084;
	wire new_net_7787;
	wire new_net_16170;
	wire new_net_18548;
	wire new_net_19958;
	wire new_net_18514;
	wire new_net_17151;
	wire new_net_16856;
	wire new_net_10514;
	wire new_net_13261;
	wire new_net_16608;
	wire new_net_16714;
	wire new_net_13508;
	wire new_net_16502;
	wire new_net_16288;
	wire new_net_17021;
	wire new_net_16794;
	wire new_net_6762;
	wire new_net_8568;
	wire _0851_;
	wire new_net_19818;
	wire new_net_20515;
	wire new_net_1143;
	wire new_net_4551;
	wire new_net_8597;
	wire new_net_9922;
	wire new_net_18645;
	wire new_net_14310;
	wire new_net_17508;
	wire new_net_7068;
	wire new_net_8332;
	wire new_net_867;
	wire _0852_;
	wire new_net_7784;
	wire new_net_8329;
	wire new_net_2447;
	wire new_net_729;
	wire new_net_3120;
	wire new_net_4559;
	wire new_net_9965;
	wire new_net_18816;
	wire new_net_20087;
	wire new_net_11778;
	wire new_net_18911;
	wire new_net_4550;
	wire new_net_8567;
	wire new_net_871;
	wire _0853_;
	wire new_net_19761;
	wire new_net_20419;
	wire new_net_21252;
	wire new_net_13662;
	wire new_net_10665;
	wire new_net_19787;
	wire new_net_15064;
	wire new_net_8557;
	wire new_net_18533;
	wire new_net_14969;
	wire new_net_405;
	wire new_net_458;
	wire new_net_811;
	wire new_net_5115;
	wire new_net_15900;
	wire new_net_15031;
	wire new_net_14911;
	wire new_net_14592;
	wire new_net_13403;
	wire new_net_4793;
	wire new_net_17200;
	wire new_net_14462;
	wire new_net_9239;
	wire new_net_17684;
	wire new_net_15118;
	wire new_net_12954;
	wire _0224_;
	wire new_net_18067;
	wire new_net_13031;
	wire new_net_6006;
	wire new_net_7742;
	wire new_net_3579;
	wire new_net_20292;
	wire new_net_21169;
	wire new_net_12576;
	wire new_net_13101;
	wire new_net_16649;
	wire new_net_18461;
	wire new_net_16358;
	wire new_net_19671;
	wire new_net_8825;
	wire new_net_1491;
	wire new_net_5123;
	wire new_net_5497;
	wire new_net_13045;
	wire new_net_6791;
	wire _0687_;
	wire _0225_;
	wire _0897_;
	wire new_net_813;
	wire new_net_5325;
	wire new_net_8716;
	wire new_net_11964;
	wire new_net_403;
	wire new_net_812;
	wire new_net_3582;
	wire new_net_6911;
	wire new_net_13406;
	wire new_net_21214;
	wire new_net_13454;
	wire new_net_9241;
	wire new_net_7920;
	wire _0688_;
	wire _0898_;
	wire _0226_;
	wire new_net_6093;
	wire new_net_19020;
	wire new_net_15775;
	wire new_net_18282;
	wire new_net_21387;
	wire new_net_9238;
	wire new_net_11016;
	wire new_net_7718;
	wire new_net_11963;
	wire new_net_2609;
	wire new_net_3580;
	wire new_net_4272;
	wire new_net_12955;
	wire new_net_11600;
	wire new_net_10134;
	wire new_net_8871;
	wire new_net_4276;
	wire new_net_7715;
	wire new_net_11965;
	wire _0227_;
	wire _0689_;
	wire _0899_;
	wire new_net_3346;
	wire new_net_3584;
	wire new_net_14988;
	wire new_net_7334;
	wire new_net_18237;
	wire new_net_17201;
	wire new_net_14276;
	wire new_net_14958;
	wire new_net_14593;
	wire new_net_17104;
	wire new_net_14463;
	wire new_net_13404;
	wire new_net_1727;
	wire new_net_4270;
	wire new_net_6101;
	wire new_net_19928;
	wire new_net_14127;
	wire new_net_17671;
	wire new_net_11839;
	wire new_net_9242;
	wire new_net_5344;
	wire _0228_;
	wire new_net_2611;
	wire _0690_;
	wire new_net_1732;
	wire _0900_;
	wire new_net_8826;
	wire new_net_20293;
	wire new_net_20343;
	wire new_net_9148;
	wire new_net_6793;
	wire new_net_4646;
	wire new_net_5116;
	wire new_net_12633;
	wire new_net_11538;
	wire new_net_21302;
	wire new_net_7921;
	wire _0229_;
	wire _0691_;
	wire new_net_14632;
	wire new_net_13539;
	wire _0901_;
	wire new_net_810;
	wire new_net_3607;
	wire new_net_13344;
	wire new_net_18984;
	wire new_net_11670;
	wire new_net_12006;
	wire new_net_13576;
	wire new_net_14548;
	wire new_net_9948;
	wire new_net_88;
	wire new_net_3340;
	wire new_net_4791;
	wire new_net_17298;
	wire new_net_4767;
	wire new_net_13732;
	wire new_net_11017;
	wire new_net_5120;
	wire new_net_7745;
	wire _0692_;
	wire _0902_;
	wire _0230_;
	wire new_net_11601;
	wire new_net_8094;
	wire new_net_18725;
	wire new_net_11966;
	wire new_net_3578;
	wire new_net_9150;
	wire new_net_17103;
	wire new_net_17202;
	wire new_net_17686;
	wire new_net_14277;
	wire new_net_14959;
	wire new_net_9941;
	wire new_net_14464;
	wire new_net_14594;
	wire new_net_6789;
	wire new_net_13405;
	wire _0693_;
	wire new_net_17535;
	wire new_net_13061;
	wire new_net_17477;
	wire new_net_3606;
	wire new_net_3950;
	wire new_net_6096;
	wire new_net_20294;
	wire new_net_9485;
	wire new_net_16753;
	wire new_net_18031;
	wire new_net_7942;
	wire new_net_9240;
	wire new_net_5496;
	wire new_net_7923;
	wire _0232_;
	wire _0694_;
	wire _0904_;
	wire new_net_456;
	wire new_net_2601;
	wire new_net_6855;
	wire new_net_11728;
	wire new_net_16534;
	wire new_net_20877;
	wire new_net_5333;
	wire new_net_9155;
	wire new_net_7720;
	wire new_net_7928;
	wire new_net_3295;
	wire new_net_20342;
	wire new_net_20854;
	wire new_net_21216;
	wire new_net_13239;
	wire new_net_12953;
	wire _0233_;
	wire _0695_;
	wire new_net_412;
	wire _0905_;
	wire new_net_18983;
	wire new_net_12330;
	wire new_net_18327;
	wire new_net_7941;
	wire new_net_11018;
	wire new_net_7926;
	wire new_net_7740;
	wire new_net_459;
	wire new_net_2608;
	wire new_net_4792;
	wire new_net_7169;
	wire new_net_12935;
	wire new_net_11602;
	wire new_net_7522;
	wire new_net_11967;
	wire new_net_460;
	wire new_net_1724;
	wire _0696_;
	wire _0906_;
	wire _0234_;
	wire new_net_1492;
	wire new_net_17102;
	wire new_net_14854;
	wire new_net_16928;
	wire new_net_17203;
	wire new_net_14465;
	wire new_net_17687;
	wire new_net_15121;
	wire new_net_14278;
	wire new_net_14960;
	wire new_net_7743;
	wire new_net_14595;
	wire new_net_1731;
	wire new_net_4788;
	wire new_net_16881;
	wire new_net_14065;
	wire new_net_8593;
	wire new_net_6912;
	wire new_net_7001;
	wire new_net_5338;
	wire _0697_;
	wire _0907_;
	wire _0235_;
	wire new_net_6856;
	wire new_net_20295;
	wire new_net_10012;
	wire new_net_7721;
	wire new_net_1497;
	wire new_net_5339;
	wire new_net_6861;
	wire new_net_21304;
	wire new_net_14662;
	wire new_net_18914;
	wire new_net_13304;
	wire new_net_8872;
	wire new_net_8820;
	wire new_net_7924;
	wire new_net_449;
	wire _0698_;
	wire _0908_;
	wire _0236_;
	wire new_net_20341;
	wire new_net_21217;
	wire new_net_1811;
	wire new_net_14560;
	wire _0042_;
	wire new_net_13715;
	wire new_net_6103;
	wire new_net_6794;
	wire new_net_84;
	wire new_net_3583;
	wire new_net_18477;
	wire new_net_18549;
	wire new_net_11603;
	wire new_net_7939;
	wire new_net_8822;
	wire new_net_11019;
	wire _0237_;
	wire _0909_;
	wire new_net_454;
	wire _0699_;
	wire new_net_13881;
	wire new_net_18982;
	wire new_net_18515;
	wire new_net_85;
	wire new_net_4004;
	wire new_net_17101;
	wire new_net_20340;
	wire new_net_16795;
	wire new_net_15122;
	wire new_net_17204;
	wire new_net_17688;
	wire new_net_14279;
	wire new_net_14961;
	wire new_net_7716;
	wire new_net_14466;
	wire new_net_14596;
	wire _0238_;
	wire _0910_;
	wire new_net_10211;
	wire new_net_7168;
	wire new_net_7927;
	wire new_net_6853;
	wire new_net_20296;
	wire new_net_14309;
	wire new_net_17509;
	wire new_net_7518;
	wire new_net_5118;
	wire _0701_;
	wire _0911_;
	wire _0239_;
	wire new_net_81;
	wire new_net_7744;
	wire new_net_21305;
	wire new_net_14543;
	wire new_net_18817;
	wire new_net_87;
	wire new_net_406;
	wire new_net_21218;
	wire new_net_11779;
	wire new_net_2656;
	wire new_net_18912;
	wire new_net_9244;
	wire _0702_;
	wire _0912_;
	wire _0240_;
	wire new_net_455;
	wire new_net_2604;
	wire new_net_19300;
	wire new_net_20339;
	wire new_net_18964;
	wire new_net_11604;
	wire new_net_8594;
	wire new_net_8819;
	wire new_net_11020;
	wire new_net_413;
	wire new_net_807;
	wire new_net_2605;
	wire new_net_6858;
	wire new_net_12292;
	wire new_net_8559;
	wire new_net_18534;
	wire new_net_8874;
	wire _0703_;
	wire _0913_;
	wire _0241_;
	wire new_net_6795;
	wire new_net_13735;
	wire new_net_17100;
	wire new_net_18981;
	wire new_net_15901;
	wire new_net_2770;
	wire new_net_15032;
	wire new_net_15123;
	wire new_net_17205;
	wire new_net_17689;
	wire new_net_14280;
	wire new_net_14962;
	wire new_net_14467;
	wire new_net_14597;
	wire new_net_4031;
	wire new_net_6097;
	wire new_net_14912;
	wire new_net_18068;
	wire new_net_4029;
	wire new_net_6098;
	wire new_net_10212;
	wire _0704_;
	wire new_net_16869;
	wire _0914_;
	wire _0242_;
	wire new_net_20297;
	wire new_net_13032;
	wire new_net_21170;
	wire new_net_12577;
	wire new_net_13102;
	wire new_net_16650;
	wire new_net_16359;
	wire new_net_78;
	wire new_net_1729;
	wire new_net_4271;
	wire new_net_4796;
	wire new_net_11968;
	wire new_net_21306;
	wire new_net_19672;
	wire new_net_13046;
	wire new_net_13738;
	wire new_net_6094;
	wire new_net_7525;
	wire new_net_7719;
	wire _0705_;
	wire _0915_;
	wire _0243_;
	wire new_net_3602;
	wire new_net_21219;
	wire new_net_13407;
	wire new_net_20063;
	wire new_net_5926;
	wire new_net_6996;
	wire new_net_12771;
	wire new_net_13455;
	wire new_net_8591;
	wire new_net_4790;
	wire new_net_9152;
	wire new_net_1494;
	wire new_net_452;
	wire new_net_19021;
	wire _1337_;
	wire new_net_15776;
	wire new_net_18283;
	wire new_net_3576;
	wire new_net_11605;
	wire new_net_4794;
	wire new_net_8827;
	wire new_net_11021;
	wire new_net_5117;
	wire _0706_;
	wire _0916_;
	wire _0244_;
	wire new_net_3297;
	wire new_net_17099;
	wire new_net_8824;
	wire new_net_1499;
	wire new_net_4008;
	wire new_net_6792;
	wire new_net_14989;
	wire new_net_7037;
	wire new_net_12948;
	wire new_net_17690;
	wire new_net_15124;
	wire new_net_7940;
	wire new_net_8590;
	wire new_net_17206;
	wire new_net_4795;
	wire new_net_14281;
	wire new_net_14963;
	wire new_net_7925;
	wire new_net_14128;
	wire new_net_1490;
	wire new_net_4027;
	wire new_net_6910;
	wire new_net_20298;
	wire new_net_11840;
	wire new_net_8821;
	wire _0708_;
	wire _0246_;
	wire _0918_;
	wire new_net_82;
	wire new_net_4006;
	wire new_net_21307;
	wire new_net_12634;
	wire new_net_14084;
	wire new_net_10110;
	wire new_net_6860;
	wire new_net_86;
	wire new_net_6790;
	wire new_net_21220;
	wire new_net_11740;
	wire new_net_13540;
	wire new_net_14633;
	wire new_net_11671;
	wire new_net_12007;
	wire new_net_13577;
	wire new_net_14547;
	wire new_net_3954;
	wire _0709_;
	wire _0919_;
	wire _0247_;
	wire new_net_808;
	wire new_net_4005;
	wire new_net_17030;
	wire new_net_4213;
	wire new_net_17299;
	wire new_net_3313;
	wire new_net_13733;
	wire new_net_13740;
	wire new_net_11606;
	wire new_net_11022;
	wire new_net_1495;
	wire new_net_3581;
	wire new_net_5121;
	wire new_net_18974;
	wire new_net_9045;
	wire new_net_17098;
	wire new_net_9149;
	wire new_net_9243;
	wire new_net_9946;
	wire _0248_;
	wire _0710_;
	wire _0920_;
	wire new_net_79;
	wire new_net_4275;
	wire new_net_10563;
	wire new_net_12947;
	wire new_net_7519;
	wire new_net_15125;
	wire new_net_17207;
	wire new_net_17691;
	wire new_net_14282;
	wire new_net_14964;
	wire new_net_1500;
	wire new_net_2603;
	wire new_net_3449;
	wire new_net_17536;
	wire new_net_13062;
	wire new_net_3575;
	wire new_net_4641;
	wire new_net_4028;
	wire new_net_7524;
	wire _0249_;
	wire _0711_;
	wire _0921_;
	wire new_net_2610;
	wire new_net_4007;
	wire new_net_18979;
	wire new_net_21308;
	wire new_net_18032;
	wire new_net_2828;
	wire new_net_9697;
	wire new_net_11727;
	wire new_net_16535;
	wire new_net_20878;
	wire _0922_;
	wire new_net_7171;
	wire new_net_9947;
	wire _0250_;
	wire new_net_13309;
	wire new_net_15627;
	wire _0712_;
	wire new_net_2607;
	wire new_net_21221;
	wire new_net_13240;
	wire new_net_5872;
	wire new_net_9154;
	wire new_net_407;
	wire new_net_6859;
	wire new_net_20338;
	wire new_net_12952;
	wire new_net_10628;
	wire new_net_12331;
	wire new_net_18328;
	wire new_net_10537;
	wire new_net_13737;
	wire new_net_11607;
	wire new_net_11023;
	wire new_net_1735;
	wire _0713_;
	wire _0923_;
	wire _0251_;
	wire new_net_12936;
	wire new_net_10845;
	wire new_net_7906;
	wire new_net_17097;
	wire new_net_8823;
	wire new_net_83;
	wire new_net_6102;
	wire new_net_6999;
	wire new_net_14855;
	wire new_net_16929;
	wire new_net_11971;
	wire new_net_13411;
	wire new_net_12946;
	wire new_net_6095;
	wire new_net_15126;
	wire new_net_17208;
	wire new_net_17692;
	wire new_net_14283;
	wire new_net_14965;
	wire new_net_9151;
	wire new_net_16882;
	wire new_net_14066;
	wire new_net_6854;
	wire new_net_7517;
	wire new_net_9942;
	wire new_net_1730;
	wire new_net_450;
	wire new_net_4033;
	wire new_net_5341;
	wire new_net_9146;
	wire _0925_;
	wire new_net_453;
	wire new_net_806;
	wire new_net_1722;
	wire _0253_;
	wire _0715_;
	wire new_net_1496;
	wire new_net_18978;
	wire new_net_14663;
	wire new_net_18915;
	wire new_net_6092;
	wire new_net_7170;
	wire new_net_9236;
	wire new_net_3956;
	wire new_net_4273;
	wire new_net_13305;
	wire new_net_14561;
	wire _0926_;
	wire new_net_1728;
	wire new_net_2613;
	wire _0254_;
	wire _0716_;
	wire new_net_1498;
	wire new_net_13716;
	wire new_net_18478;
	wire new_net_13741;
	wire new_net_11608;
	wire new_net_9944;
	wire new_net_11024;
	wire new_net_2602;
	wire new_net_3952;
	wire new_net_4645;
	wire new_net_16172;
	wire new_net_18550;
	wire new_net_18516;
	wire new_net_6857;
	wire new_net_17096;
	wire new_net_4026;
	wire new_net_9147;
	wire new_net_9945;
	wire _0927_;
	wire _0255_;
	wire _0717_;
	wire new_net_20337;
	wire new_net_16796;
	wire new_net_11972;
	wire new_net_13412;
	wire new_net_12945;
	wire new_net_15127;
	wire new_net_17209;
	wire new_net_17693;
	wire new_net_14284;
	wire new_net_14966;
	wire new_net_815;
	wire new_net_14471;
	wire new_net_9949;
	wire new_net_2606;
	wire _0718_;
	wire _0928_;
	wire _0256_;
	wire new_net_5119;
	wire new_net_3275;
	wire new_net_16422;
	wire new_net_17510;
	wire new_net_9943;
	wire new_net_3605;
	wire new_net_4789;
	wire new_net_6099;
	wire new_net_21310;
	wire new_net_16703;
	wire new_net_3194;
	wire new_net_4030;
	wire _0257_;
	wire new_net_1723;
	wire _0719_;
	wire _0929_;
	wire new_net_7717;
	wire new_net_18977;
	wire new_net_20334;
	wire new_net_14544;
	wire new_net_18818;
	wire new_net_11780;
	wire new_net_13978;
	wire new_net_4642;
	wire new_net_20335;
	wire new_net_9476;
	wire new_net_11609;
	wire _0258_;
	wire _0930_;
	wire _0720_;
	wire _0896_;
	wire new_net_3577;
	wire new_net_4002;
	wire new_net_11025;
	wire new_net_8659;
	wire new_net_19789;
	wire new_net_12293;
	wire new_net_15066;
	wire new_net_18535;
	wire new_net_7746;
	wire new_net_17095;
	wire new_net_7523;
	wire new_net_457;
	wire new_net_809;
	wire new_net_1726;
	wire new_net_3601;
	wire new_net_6913;
	wire new_net_20336;
	wire new_net_14971;
	wire new_net_20943;
	wire _1340_;
	wire new_net_15902;
	wire new_net_15033;
	wire new_net_11973;
	wire new_net_17694;
	wire new_net_12944;
	wire new_net_6100;
	wire new_net_15128;
	wire new_net_411;
	wire new_net_17210;
	wire new_net_14285;
	wire new_net_14967;
	wire new_net_13413;
	wire new_net_14913;
	wire new_net_18162;
	wire new_net_16915;
	wire new_net_18069;
	wire new_net_4647;
	wire new_net_7919;
	wire new_net_11895;
	wire new_net_12554;
	wire new_net_16870;
	wire new_net_13033;
	wire new_net_21171;
	wire new_net_5567;
	wire new_net_6667;
	wire new_net_12578;
	wire new_net_13103;
	wire new_net_3604;
	wire new_net_4274;
	wire new_net_409;
	wire _0722_;
	wire _0932_;
	wire _0260_;
	wire new_net_451;
	wire new_net_1734;
	wire new_net_21311;
	wire new_net_19673;
	wire new_net_13047;
	wire new_net_18963;
	wire new_net_7000;
	wire new_net_6862;
	wire new_net_8589;
	wire new_net_1493;
	wire new_net_80;
	wire new_net_4643;
	wire new_net_5122;
	wire new_net_9373;
	wire new_net_13408;
	wire _0723_;
	wire _0933_;
	wire _0261_;
	wire new_net_814;
	wire new_net_1733;
	wire new_net_9237;
	wire new_net_18976;
	wire new_net_19022;
	wire new_net_15777;
	wire new_net_18284;
	wire new_net_21386;
	wire new_net_17093;
	wire new_net_7520;
	wire new_net_3603;
	wire new_net_11026;
	wire new_net_14862;
	wire new_net_14776;
	wire new_net_13736;
	wire new_net_17094;
	wire _0724_;
	wire _0934_;
	wire _0262_;
	wire new_net_14990;
	wire new_net_7002;
	wire new_net_14473;
	wire new_net_14603;
	wire new_net_13414;
	wire new_net_13739;
	wire new_net_15129;
	wire new_net_17211;
	wire new_net_17695;
	wire new_net_14286;
	wire new_net_14968;
	wire new_net_14129;
	wire new_net_5498;
	wire new_net_1736;
	wire new_net_7739;
	wire new_net_11974;
	wire new_net_4644;
	wire new_net_7521;
	wire new_net_8873;
	wire new_net_9153;
	wire _0725_;
	wire _0935_;
	wire new_net_11841;
	wire new_net_15971;
	wire new_net_8748;
	wire new_net_7747;
	wire new_net_18973;
	wire new_net_21312;
	wire new_net_12635;
	wire new_net_14085;
	wire new_net_11540;
	wire _0726_;
	wire _0936_;
	wire _0264_;
	wire new_net_5342;
	wire new_net_11741;
	wire new_net_13541;
	wire new_net_14634;
	wire new_net_11672;
	wire new_net_402;
	wire new_net_20333;
	wire new_net_13578;
	wire new_net_12008;
	wire new_net_14546;
	wire new_net_17031;
	wire new_net_11027;
	wire new_net_3948;
	wire _0937_;
	wire _0727_;
	wire _0265_;
	wire new_net_18975;
	wire new_net_13734;
	wire new_net_2424;
	wire new_net_10565;
	wire new_net_15473;
	wire new_net_9638;
	wire new_net_7888;
	wire new_net_10685;
	wire new_net_2233;
	wire new_net_6029;
	wire new_net_6110;
	wire new_net_19935;
	wire new_net_17537;
	wire new_net_6531;
	wire new_net_13063;
	wire new_net_13357;
	wire new_net_14486;
	wire new_net_16479;
	wire new_net_16951;
	wire new_net_12873;
	wire new_net_14802;
	wire new_net_17022;
	wire new_net_17435;
	wire new_net_13875;
	wire new_net_17330;
	wire new_net_16755;
	wire new_net_18033;
	wire new_net_9646;
	wire new_net_1682;
	wire new_net_389;
	wire new_net_1218;
	wire new_net_1344;
	wire new_net_1862;
	wire new_net_5994;
	wire new_net_20268;
	wire new_net_12729;
	wire new_net_13191;
	wire new_net_13448;
	wire new_net_11726;
	wire new_net_16536;
	wire new_net_10682;
	wire new_net_394;
	wire new_net_6266;
	wire new_net_2757;
	wire new_net_3960;
	wire new_net_6031;
	wire new_net_747;
	wire _0057_;
	wire new_net_19351;
	wire new_net_19399;
	wire new_net_20856;
	wire new_net_13241;
	wire new_net_9383;
	wire new_net_10318;
	wire new_net_6696;
	wire new_net_34;
	wire new_net_397;
	wire new_net_12951;
	wire new_net_12332;
	wire new_net_18329;
	wire new_net_5232;
	wire new_net_10329;
	wire _0058_;
	wire new_net_1681;
	wire new_net_12937;
	wire _1342_;
	wire new_net_10681;
	wire new_net_16216;
	wire new_net_3342;
	wire new_net_4018;
	wire new_net_2232;
	wire new_net_1229;
	wire new_net_1037;
	wire new_net_14856;
	wire new_net_16930;
	wire new_net_8580;
	wire new_net_6699;
	wire new_net_13756;
	wire new_net_5991;
	wire new_net_1863;
	wire new_net_2222;
	wire new_net_2650;
	wire _0059_;
	wire new_net_1924;
	wire new_net_19936;
	wire new_net_16883;
	wire _1736_;
	wire new_net_14067;
	wire new_net_13358;
	wire new_net_14487;
	wire new_net_16480;
	wire new_net_16952;
	wire new_net_12874;
	wire new_net_14803;
	wire new_net_17023;
	wire new_net_13876;
	wire new_net_17331;
	wire new_net_15345;
	wire new_net_19904;
	wire new_net_5906;
	wire new_net_6914;
	wire new_net_5155;
	wire _0060_;
	wire new_net_20269;
	wire new_net_14664;
	wire new_net_18916;
	wire new_net_9059;
	wire new_net_9463;
	wire new_net_7890;
	wire new_net_6698;
	wire new_net_6113;
	wire new_net_1224;
	wire new_net_1685;
	wire new_net_4569;
	wire new_net_13306;
	wire new_net_19352;
	wire new_net_19400;
	wire new_net_7872;
	wire new_net_14562;
	wire _0049_;
	wire new_net_16147;
	wire _0061_;
	wire new_net_13717;
	wire new_net_18479;
	wire new_net_9645;
	wire new_net_13755;
	wire new_net_2224;
	wire new_net_2648;
	wire new_net_6036;
	wire new_net_16173;
	wire new_net_18551;
	wire new_net_13883;
	wire new_net_18517;
	wire new_net_6690;
	wire new_net_10686;
	wire new_net_3249;
	wire new_net_6917;
	wire new_net_4565;
	wire new_net_6262;
	wire _0062_;
	wire new_net_16797;
	wire new_net_6466;
	wire new_net_10316;
	wire new_net_17434;
	wire new_net_6922;
	wire new_net_2653;
	wire new_net_3244;
	wire new_net_19937;
	wire new_net_13359;
	wire new_net_14488;
	wire new_net_16481;
	wire new_net_16953;
	wire new_net_12875;
	wire new_net_14804;
	wire new_net_17024;
	wire new_net_13877;
	wire new_net_17332;
	wire new_net_4567;
	wire new_net_16423;
	wire new_net_17511;
	wire new_net_13155;
	wire new_net_21093;
	wire new_net_6467;
	wire new_net_13754;
	wire new_net_16215;
	wire new_net_4570;
	wire new_net_5153;
	wire new_net_9619;
	wire new_net_35;
	wire new_net_3248;
	wire new_net_20270;
	wire new_net_16704;
	wire new_net_5687;
	wire new_net_4092;
	wire new_net_4168;
	wire new_net_6114;
	wire _0064_;
	wire new_net_3278;
	wire new_net_19353;
	wire new_net_19401;
	wire new_net_19642;
	wire new_net_11781;
	wire new_net_752;
	wire new_net_5157;
	wire new_net_6116;
	wire new_net_15734;
	wire new_net_20428;
	wire new_net_5233;
	wire _0065_;
	wire new_net_746;
	wire new_net_3393;
	wire new_net_6032;
	wire new_net_12294;
	wire new_net_15067;
	wire new_net_5683;
	wire new_net_7892;
	wire new_net_1922;
	wire new_net_1351;
	wire new_net_3388;
	wire new_net_4016;
	wire new_net_14972;
	wire new_net_15903;
	wire new_net_15034;
	wire new_net_6037;
	wire new_net_17433;
	wire new_net_4015;
	wire new_net_6919;
	wire new_net_3386;
	wire new_net_32;
	wire new_net_2220;
	wire _0066_;
	wire new_net_17152;
	wire new_net_14914;
	wire new_net_18163;
	wire new_net_16916;
	wire new_net_7316;
	wire new_net_18070;
	wire new_net_15986;
	wire new_net_16918;
	wire new_net_13360;
	wire new_net_14489;
	wire new_net_16482;
	wire new_net_16954;
	wire new_net_12876;
	wire new_net_14805;
	wire new_net_17025;
	wire new_net_13878;
	wire new_net_11896;
	wire new_net_12555;
	wire new_net_13034;
	wire new_net_21172;
	wire new_net_12579;
	wire new_net_16652;
	wire new_net_13104;
	wire new_net_4174;
	wire new_net_7898;
	wire new_net_16214;
	wire new_net_4561;
	wire new_net_5701;
	wire new_net_5993;
	wire _0067_;
	wire new_net_3401;
	wire new_net_20271;
	wire new_net_19674;
	wire new_net_13048;
	wire new_net_13604;
	wire new_net_9637;
	wire new_net_4014;
	wire new_net_1342;
	wire new_net_1859;
	wire new_net_31;
	wire new_net_384;
	wire new_net_750;
	wire new_net_1220;
	wire new_net_3398;
	wire new_net_19354;
	wire new_net_9376;
	wire new_net_13409;
	wire new_net_12773;
	wire new_net_13457;
	wire new_net_9234;
	wire new_net_7894;
	wire new_net_8587;
	wire new_net_1222;
	wire new_net_386;
	wire new_net_1860;
	wire _0068_;
	wire new_net_19023;
	wire _1344_;
	wire new_net_15778;
	wire new_net_18285;
	wire new_net_10319;
	wire new_net_6694;
	wire new_net_10683;
	wire new_net_749;
	wire new_net_5908;
	wire new_net_6111;
	wire new_net_14777;
	wire new_net_10321;
	wire new_net_6027;
	wire new_net_1919;
	wire _0069_;
	wire new_net_5154;
	wire new_net_1223;
	wire new_net_13449;
	wire new_net_17432;
	wire new_net_1861;
	wire new_net_10324;
	wire new_net_19939;
	wire new_net_1585;
	wire new_net_14130;
	wire new_net_15987;
	wire new_net_16919;
	wire new_net_13361;
	wire new_net_16931;
	wire new_net_14490;
	wire new_net_16483;
	wire new_net_12877;
	wire new_net_14806;
	wire new_net_17026;
	wire new_net_15465;
	wire new_net_11842;
	wire new_net_15972;
	wire new_net_21415;
	wire new_net_16213;
	wire new_net_5699;
	wire new_net_751;
	wire new_net_399;
	wire new_net_3395;
	wire new_net_20272;
	wire new_net_7436;
	wire new_net_7990;
	wire new_net_6697;
	wire new_net_3250;
	wire new_net_6921;
	wire new_net_6112;
	wire new_net_13753;
	wire new_net_1228;
	wire _0071_;
	wire new_net_396;
	wire new_net_5156;
	wire new_net_11742;
	wire new_net_13542;
	wire new_net_14635;
	wire new_net_11673;
	wire new_net_12009;
	wire new_net_13579;
	wire new_net_7991;
	wire new_net_9460;
	wire new_net_8586;
	wire new_net_10317;
	wire new_net_5689;
	wire new_net_17032;
	wire new_net_10816;
	wire new_net_4221;
	wire new_net_385;
	wire _0072_;
	wire new_net_9047;
	wire new_net_1679;
	wire new_net_755;
	wire new_net_1225;
	wire new_net_2221;
	wire new_net_3341;
	wire new_net_4175;
	wire new_net_5160;
	wire new_net_5989;
	wire new_net_10323;
	wire new_net_20920;
	wire new_net_15474;
	wire new_net_4224;
	wire new_net_5684;
	wire new_net_13749;
	wire new_net_17431;
	wire new_net_393;
	wire _0073_;
	wire new_net_6265;
	wire new_net_19940;
	wire new_net_17538;
	wire new_net_3417;
	wire new_net_15988;
	wire new_net_16920;
	wire new_net_16956;
	wire new_net_13362;
	wire new_net_6468;
	wire new_net_14491;
	wire new_net_12878;
	wire new_net_13752;
	wire new_net_14807;
	wire new_net_13880;
	wire new_net_13064;
	wire new_net_4225;
	wire new_net_9464;
	wire new_net_4172;
	wire new_net_8584;
	wire new_net_16212;
	wire new_net_390;
	wire new_net_6916;
	wire new_net_1683;
	wire _0074_;
	wire new_net_16756;
	wire new_net_18034;
	wire new_net_12728;
	wire new_net_13192;
	wire new_net_16537;
	wire new_net_20880;
	wire new_net_9616;
	wire new_net_6473;
	wire new_net_2225;
	wire new_net_1686;
	wire new_net_30;
	wire new_net_388;
	wire new_net_19356;
	wire new_net_19404;
	wire new_net_19645;
	wire new_net_13311;
	wire new_net_15629;
	wire new_net_20857;
	wire new_net_13242;
	wire new_net_5700;
	wire new_net_9641;
	wire new_net_13751;
	wire _0075_;
	wire new_net_2652;
	wire new_net_3243;
	wire new_net_4012;
	wire new_net_19708;
	wire _0700_;
	wire new_net_12950;
	wire new_net_18762;
	wire new_net_12333;
	wire new_net_18330;
	wire new_net_9644;
	wire new_net_4173;
	wire new_net_12938;
	wire new_net_7690;
	wire new_net_17335;
	wire new_net_5681;
	wire new_net_9622;
	wire new_net_6030;
	wire new_net_1219;
	wire new_net_1341;
	wire _0076_;
	wire new_net_1690;
	wire new_net_14857;
	wire new_net_9620;
	wire new_net_17430;
	wire new_net_7896;
	wire new_net_29;
	wire new_net_3246;
	wire new_net_4568;
	wire new_net_19941;
	wire new_net_16884;
	wire new_net_5158;
	wire new_net_5698;
	wire new_net_17028;
	wire new_net_13363;
	wire new_net_6026;
	wire new_net_15989;
	wire new_net_16485;
	wire new_net_15467;
	wire new_net_16957;
	wire new_net_16921;
	wire new_net_14068;
	wire new_net_9621;
	wire new_net_6692;
	wire new_net_16211;
	wire new_net_398;
	wire new_net_745;
	wire new_net_3964;
	wire new_net_6115;
	wire new_net_20274;
	wire new_net_14665;
	wire new_net_18917;
	wire new_net_8579;
	wire new_net_2229;
	wire new_net_1689;
	wire _0078_;
	wire new_net_19357;
	wire new_net_19405;
	wire new_net_13307;
	wire new_net_7867;
	wire new_net_1802;
	wire new_net_6750;
	wire new_net_14563;
	wire new_net_7897;
	wire new_net_10320;
	wire new_net_10684;
	wire new_net_2655;
	wire new_net_391;
	wire new_net_3242;
	wire new_net_4017;
	wire new_net_16148;
	wire new_net_13718;
	wire new_net_18480;
	wire new_net_6465;
	wire new_net_28;
	wire _0079_;
	wire new_net_16174;
	wire new_net_18552;
	wire new_net_13884;
	wire new_net_5657;
	wire new_net_15083;
	wire new_net_18518;
	wire new_net_5145;
	wire new_net_5914;
	wire new_net_6470;
	wire new_net_8588;
	wire new_net_1916;
	wire new_net_3968;
	wire new_net_6117;
	wire new_net_5983;
	wire new_net_10327;
	wire new_net_5913;
	wire new_net_7887;
	wire new_net_17429;
	wire new_net_37;
	wire new_net_2649;
	wire _0080_;
	wire new_net_1350;
	wire new_net_19942;
	wire new_net_15468;
	wire new_net_16934;
	wire new_net_15990;
	wire new_net_16922;
	wire new_net_13364;
	wire new_net_14493;
	wire new_net_16486;
	wire new_net_16958;
	wire new_net_12880;
	wire new_net_13882;
	wire new_net_3103;
	wire new_net_6967;
	wire new_net_16424;
	wire new_net_17512;
	wire new_net_13156;
	wire new_net_6263;
	wire new_net_10322;
	wire new_net_4169;
	wire new_net_6469;
	wire new_net_16210;
	wire _0081_;
	wire new_net_753;
	wire new_net_4013;
	wire new_net_20275;
	wire new_net_4552;
	wire new_net_16705;
	wire new_net_36;
	wire new_net_4219;
	wire new_net_5987;
	wire new_net_19358;
	wire new_net_19406;
	wire new_net_3357;
	wire new_net_11077;
	wire new_net_11782;
	wire new_net_9465;
	wire new_net_5911;
	wire new_net_387;
	wire _0082_;
	wire new_net_1349;
	wire new_net_6118;
	wire new_net_15735;
	wire new_net_20429;
	wire new_net_7895;
	wire new_net_13750;
	wire new_net_14808;
	wire new_net_6920;
	wire new_net_1925;
	wire _0903_;
	wire new_net_12295;
	wire new_net_15068;
	wire new_net_4562;
	wire new_net_9615;
	wire new_net_4217;
	wire new_net_5915;
	wire new_net_17029;
	wire new_net_1343;
	wire new_net_2226;
	wire _0083_;
	wire new_net_3402;
	wire new_net_17953;
	wire new_net_14973;
	wire new_net_7057;
	wire new_net_15904;
	wire new_net_15035;
	wire new_net_9642;
	wire new_net_17428;
	wire new_net_4215;
	wire new_net_19943;
	wire new_net_10176;
	wire new_net_17153;
	wire new_net_5108;
	wire new_net_14915;
	wire new_net_18164;
	wire new_net_10602;
	wire new_net_16917;
	wire new_net_18071;
	wire new_net_15352;
	wire new_net_15469;
	wire new_net_16935;
	wire new_net_15991;
	wire new_net_16923;
	wire new_net_9461;
	wire new_net_13365;
	wire new_net_14494;
	wire new_net_16487;
	wire new_net_12881;
	wire new_net_11897;
	wire new_net_12556;
	wire new_net_16872;
	wire new_net_13035;
	wire new_net_21173;
	wire new_net_12580;
	wire new_net_9624;
	wire new_net_8582;
	wire new_net_16209;
	wire new_net_1761;
	wire new_net_13105;
	wire new_net_16653;
	wire new_net_1918;
	wire new_net_2228;
	wire new_net_3280;
	wire new_net_6918;
	wire new_net_18783;
	wire new_net_19675;
	wire new_net_5324;
	wire new_net_13049;
	wire new_net_1884;
	wire new_net_8585;
	wire new_net_13605;
	wire new_net_1917;
	wire new_net_27;
	wire new_net_2223;
	wire _0085_;
	wire new_net_3403;
	wire new_net_19359;
	wire new_net_19407;
	wire new_net_13410;
	wire new_net_1680;
	wire new_net_4566;
	wire new_net_12774;
	wire new_net_13458;
	wire new_net_19024;
	wire new_net_15779;
	wire new_net_18286;
	wire new_net_5152;
	wire new_net_10325;
	wire new_net_6028;
	wire _0086_;
	wire new_net_14778;
	wire new_net_13748;
	wire new_net_1687;
	wire new_net_4563;
	wire new_net_5151;
	wire new_net_4220;
	wire new_net_9462;
	wire new_net_5909;
	wire new_net_6464;
	wire new_net_17427;
	wire new_net_1927;
	wire _0087_;
	wire new_net_4204;
	wire new_net_19944;
	wire new_net_16360;
	wire new_net_14131;
	wire new_net_15353;
	wire new_net_15470;
	wire new_net_16936;
	wire new_net_7989;
	wire new_net_15992;
	wire new_net_16924;
	wire new_net_13366;
	wire new_net_14495;
	wire new_net_16488;
	wire new_net_16960;
	wire new_net_4000;
	wire new_net_16079;
	wire new_net_11843;
	wire new_net_15973;
	wire new_net_4560;
	wire new_net_5988;
	wire new_net_3404;
	wire new_net_9466;
	wire new_net_9639;
	wire new_net_6471;
	wire new_net_7889;
	wire new_net_16208;
	wire _0088_;
	wire new_net_20277;
	wire new_net_8472;
	wire _1348_;
	wire new_net_1926;
	wire new_net_1227;
	wire new_net_4564;
	wire new_net_19360;
	wire new_net_19408;
	wire new_net_13543;
	wire new_net_14636;
	wire new_net_9640;
	wire new_net_6472;
	wire new_net_6693;
	wire new_net_16207;
	wire new_net_11674;
	wire new_net_2651;
	wire _0089_;
	wire new_net_3247;
	wire new_net_13580;
	wire new_net_11111;
	wire new_net_19822;
	wire new_net_5990;
	wire new_net_6463;
	wire new_net_7893;
	wire new_net_10314;
	wire new_net_6695;
	wire new_net_13745;
	wire new_net_2645;
	wire new_net_744;
	wire new_net_3277;
	wire new_net_5234;
	wire new_net_10817;
	wire new_net_17302;
	wire new_net_18459;
	wire new_net_5697;
	wire new_net_9618;
	wire new_net_3966;
	wire new_net_10679;
	wire _0090_;
	wire new_net_33;
	wire new_net_392;
	wire new_net_18253;
	wire new_net_9235;
	wire new_net_5682;
	wire new_net_5912;
	wire new_net_8578;
	wire new_net_13746;
	wire new_net_17426;
	wire new_net_395;
	wire new_net_3389;
	wire new_net_19945;
	wire new_net_15475;
	wire new_net_17539;
	wire new_net_15354;
	wire new_net_15471;
	wire new_net_16937;
	wire new_net_16925;
	wire _0091_;
	wire new_net_13367;
	wire new_net_4171;
	wire new_net_14496;
	wire new_net_16489;
	wire new_net_16961;
	wire new_net_13065;
	wire new_net_17480;
	wire new_net_6915;
	wire new_net_5992;
	wire new_net_7891;
	wire new_net_17424;
	wire new_net_4170;
	wire new_net_4656;
	wire new_net_5907;
	wire new_net_20278;
	wire new_net_18035;
	wire new_net_12727;
	wire new_net_13193;
	wire new_net_6264;
	wire new_net_9617;
	wire new_net_5686;
	wire _0092_;
	wire new_net_19361;
	wire new_net_19409;
	wire new_net_20881;
	wire new_net_13312;
	wire new_net_15630;
	wire new_net_20858;
	wire new_net_13243;
	wire new_net_10680;
	wire new_net_2654;
	wire new_net_3245;
	wire new_net_9458;
	wire new_net_16998;
	wire new_net_13851;
	wire new_net_12949;
	wire new_net_18763;
	wire new_net_5985;
	wire new_net_5905;
	wire new_net_10315;
	wire new_net_12334;
	wire new_net_16206;
	wire _0093_;
	wire new_net_18331;
	wire new_net_12939;
	wire new_net_7992;
	wire new_net_15993;
	wire new_net_8581;
	wire new_net_1928;
	wire new_net_3241;
	wire new_net_7977;
	wire new_net_14858;
	wire new_net_6034;
	wire new_net_9643;
	wire new_net_5910;
	wire new_net_8583;
	wire new_net_6691;
	wire new_net_13747;
	wire new_net_17425;
	wire _0094_;
	wire new_net_19946;
	wire new_net_5986;
	wire new_net_16932;
	wire new_net_16885;
	wire new_net_13886;
	wire new_net_17340;
	wire new_net_15355;
	wire new_net_15472;
	wire new_net_16938;
	wire new_net_16926;
	wire new_net_13368;
	wire new_net_14497;
	wire new_net_16490;
	wire new_net_16962;
	wire _1743_;
	wire new_net_14069;
	wire new_net_4710;
	wire new_net_4216;
	wire new_net_400;
	wire new_net_1858;
	wire new_net_1921;
	wire _0095_;
	wire new_net_20279;
	wire new_net_6394;
	wire new_net_14666;
	wire new_net_18918;
	wire new_net_2646;
	wire new_net_754;
	wire new_net_5984;
	wire new_net_9459;
	wire new_net_19362;
	wire new_net_19410;
	wire new_net_13308;
	wire new_net_1798;
	wire new_net_6035;
	wire new_net_10313;
	wire _0096_;
	wire new_net_1347;
	wire new_net_1920;
	wire new_net_16149;
	wire new_net_13719;
	wire new_net_18481;
	wire new_net_4093;
	wire new_net_470;
	wire new_net_6077;
	wire new_net_8760;
	wire new_net_16175;
	wire new_net_18553;
	wire new_net_13885;
	wire new_net_5159;
	wire new_net_4222;
	wire _0097_;
	wire new_net_2227;
	wire new_net_1688;
	wire new_net_3962;
	wire new_net_18519;
	wire _0434_;
	wire new_net_352;
	wire new_net_918;
	wire new_net_731;
	wire new_net_8745;
	wire new_net_5363;
	wire new_net_19959;
	wire new_net_21226;
	wire new_net_21095;
	wire new_net_351;
	wire _0728_;
	wire new_net_1195;
	wire new_net_1617;
	wire new_net_12127;
	wire new_net_12362;
	wire new_net_13957;
	wire new_net_16265;
	wire new_net_15911;
	wire new_net_14921;
	wire new_net_356;
	wire new_net_3177;
	wire new_net_8829;
	wire new_net_9377;
	wire new_net_219;
	wire new_net_1619;
	wire _0729_;
	wire new_net_926;
	wire new_net_19411;
	wire new_net_20311;
	wire new_net_21236;
	wire new_net_20430;
	wire new_net_10630;
	wire new_net_19482;
	wire new_net_21407;
	wire _0730_;
	wire new_net_359;
	wire new_net_20679;
	wire new_net_4240;
	wire new_net_11263;
	wire new_net_7495;
	wire new_net_9783;
	wire new_net_10874;
	wire new_net_11667;
	wire new_net_18165;
	wire new_net_18072;
	wire _0731_;
	wire new_net_223;
	wire new_net_354;
	wire new_net_8835;
	wire new_net_19960;
	wire new_net_20021;
	wire new_net_20319;
	wire new_net_21174;
	wire new_net_16654;
	wire new_net_924;
	wire new_net_5540;
	wire new_net_8228;
	wire new_net_12341;
	wire new_net_13852;
	wire new_net_15191;
	wire new_net_16159;
	wire new_net_16999;
	wire new_net_12128;
	wire new_net_12363;
	wire new_net_18784;
	wire new_net_19676;
	wire _0732_;
	wire new_net_3396;
	wire new_net_10625;
	wire new_net_8736;
	wire new_net_9528;
	wire new_net_20030;
	wire new_net_3399;
	wire new_net_5364;
	wire new_net_9535;
	wire new_net_19412;
	wire new_net_19025;
	wire _1351_;
	wire new_net_18287;
	wire _0733_;
	wire new_net_511;
	wire new_net_3173;
	wire new_net_3332;
	wire new_net_3494;
	wire new_net_7496;
	wire new_net_21408;
	wire new_net_738;
	wire new_net_3330;
	wire new_net_9790;
	wire new_net_8828;
	wire new_net_20029;
	wire new_net_20680;
	wire new_net_19624;
	wire new_net_1221;
	wire _0734_;
	wire new_net_2596;
	wire new_net_3182;
	wire new_net_3444;
	wire new_net_9686;
	wire new_net_11264;
	wire new_net_4971;
	wire new_net_10875;
	wire new_net_218;
	wire new_net_512;
	wire new_net_8749;
	wire new_net_8830;
	wire new_net_19961;
	wire new_net_21225;
	wire new_net_19898;
	wire _0735_;
	wire new_net_515;
	wire new_net_1613;
	wire new_net_357;
	wire new_net_12342;
	wire new_net_13853;
	wire new_net_15192;
	wire new_net_16160;
	wire new_net_17000;
	wire new_net_12129;
	wire new_net_9124;
	wire new_net_1621;
	wire new_net_3175;
	wire new_net_3498;
	wire new_net_9687;
	wire new_net_1140;
	wire _0736_;
	wire new_net_1186;
	wire new_net_3337;
	wire new_net_19413;
	wire new_net_20028;
	wire new_net_3500;
	wire new_net_8834;
	wire new_net_19471;
	wire new_net_17303;
	wire new_net_21409;
	wire new_net_17685;
	wire _0737_;
	wire new_net_1190;
	wire new_net_8231;
	wire new_net_4613;
	wire new_net_925;
	wire new_net_18254;
	wire new_net_20681;
	wire new_net_742;
	wire new_net_5365;
	wire new_net_10876;
	wire _0738_;
	wire new_net_5532;
	wire new_net_9782;
	wire new_net_19962;
	wire new_net_20313;
	wire new_net_13430;
	wire new_net_1192;
	wire new_net_2591;
	wire new_net_12343;
	wire new_net_13854;
	wire new_net_15193;
	wire new_net_16161;
	wire new_net_17001;
	wire new_net_12130;
	wire new_net_12365;
	wire new_net_18036;
	wire new_net_20882;
	wire new_net_919;
	wire _0739_;
	wire new_net_19276;
	wire new_net_5334;
	wire new_net_18831;
	wire new_net_3495;
	wire new_net_10269;
	wire new_net_10629;
	wire new_net_19414;
	wire new_net_19480;
	wire new_net_21234;
	wire _0707_;
	wire new_net_18764;
	wire new_net_18332;
	wire _0740_;
	wire new_net_217;
	wire new_net_3276;
	wire new_net_4233;
	wire new_net_9689;
	wire new_net_519;
	wire new_net_11265;
	wire new_net_5023;
	wire new_net_1616;
	wire new_net_21410;
	wire new_net_3174;
	wire new_net_9693;
	wire new_net_19277;
	wire new_net_20682;
	wire new_net_350;
	wire _0741_;
	wire new_net_9381;
	wire new_net_8227;
	wire new_net_7489;
	wire new_net_16933;
	wire new_net_8742;
	wire new_net_10877;
	wire new_net_522;
	wire new_net_2598;
	wire new_net_4260;
	wire new_net_9527;
	wire new_net_19963;
	wire _0742_;
	wire new_net_917;
	wire new_net_13431;
	wire new_net_7236;
	wire new_net_12344;
	wire new_net_13855;
	wire new_net_15194;
	wire new_net_16162;
	wire new_net_12131;
	wire new_net_12366;
	wire new_net_18919;
	wire new_net_931;
	wire new_net_2597;
	wire new_net_5533;
	wire new_net_8747;
	wire _0743_;
	wire new_net_1189;
	wire new_net_2592;
	wire new_net_3493;
	wire new_net_8833;
	wire new_net_9457;
	wire new_net_9529;
	wire new_net_8226;
	wire new_net_9692;
	wire new_net_11273;
	wire new_net_18482;
	wire new_net_1623;
	wire new_net_7493;
	wire new_net_21411;
	wire new_net_18554;
	wire new_net_18520;
	wire _0744_;
	wire new_net_216;
	wire new_net_1187;
	wire new_net_9532;
	wire new_net_7237;
	wire new_net_20683;
	wire new_net_1618;
	wire new_net_3703;
	wire new_net_9378;
	wire new_net_11266;
	wire new_net_8750;
	wire new_net_10878;
	wire new_net_19478;
	wire new_net_20309;
	wire new_net_21232;
	wire new_net_355;
	wire new_net_920;
	wire _0745_;
	wire new_net_2594;
	wire new_net_3700;
	wire new_net_9379;
	wire new_net_7231;
	wire new_net_9797;
	wire new_net_5024;
	wire new_net_10627;
	wire new_net_4232;
	wire new_net_5538;
	wire new_net_16270;
	wire new_net_13432;
	wire new_net_12345;
	wire new_net_13856;
	wire new_net_15195;
	wire new_net_16163;
	wire new_net_17003;
	wire new_net_9690;
	wire new_net_21096;
	wire new_net_8744;
	wire new_net_1614;
	wire _0746_;
	wire new_net_3161;
	wire new_net_3183;
	wire new_net_4235;
	wire new_net_20234;
	wire new_net_7491;
	wire new_net_8831;
	wire new_net_9372;
	wire new_net_19416;
	wire new_net_20027;
	wire new_net_1612;
	wire _0747_;
	wire new_net_5539;
	wire new_net_7498;
	wire new_net_10626;
	wire new_net_19477;
	wire new_net_21233;
	wire new_net_21412;
	wire new_net_4617;
	wire new_net_9795;
	wire new_net_20312;
	wire new_net_20684;
	wire new_net_10879;
	wire new_net_2593;
	wire _0748_;
	wire new_net_930;
	wire new_net_11267;
	wire new_net_20308;
	wire new_net_18166;
	wire new_net_19230;
	wire new_net_3702;
	wire new_net_7079;
	wire new_net_19965;
	wire new_net_18073;
	wire new_net_21175;
	wire new_net_14667;
	wire _0749_;
	wire new_net_3699;
	wire new_net_13433;
	wire new_net_12346;
	wire new_net_13857;
	wire new_net_15196;
	wire new_net_16164;
	wire new_net_17004;
	wire new_net_12133;
	wire new_net_18785;
	wire new_net_19677;
	wire new_net_353;
	wire new_net_928;
	wire new_net_8229;
	wire new_net_9536;
	wire _0750_;
	wire new_net_743;
	wire new_net_3168;
	wire new_net_9530;
	wire new_net_8233;
	wire new_net_4237;
	wire new_net_16586;
	wire new_net_19417;
	wire new_net_19026;
	wire new_net_18288;
	wire new_net_3163;
	wire new_net_8739;
	wire new_net_9531;
	wire new_net_21413;
	wire _0751_;
	wire new_net_514;
	wire new_net_7233;
	wire new_net_20026;
	wire new_net_20685;
	wire new_net_19625;
	wire new_net_922;
	wire new_net_10880;
	wire new_net_11268;
	wire new_net_18709;
	wire _0752_;
	wire new_net_741;
	wire new_net_3170;
	wire new_net_3180;
	wire new_net_11661;
	wire new_net_7078;
	wire new_net_19966;
	wire new_net_15975;
	wire new_net_358;
	wire new_net_3334;
	wire new_net_5025;
	wire new_net_15197;
	wire new_net_8737;
	wire new_net_14668;
	wire new_net_13434;
	wire new_net_8230;
	wire new_net_12134;
	wire new_net_12369;
	wire new_net_21230;
	wire _0753_;
	wire new_net_222;
	wire new_net_2599;
	wire new_net_3167;
	wire new_net_9792;
	wire new_net_8753;
	wire new_net_732;
	wire new_net_9788;
	wire new_net_19418;
	wire new_net_20024;
	wire new_net_20315;
	wire _0754_;
	wire new_net_2595;
	wire new_net_7080;
	wire new_net_7497;
	wire new_net_9775;
	wire new_net_21414;
	wire new_net_736;
	wire new_net_927;
	wire new_net_4234;
	wire new_net_10267;
	wire new_net_19278;
	wire new_net_20025;
	wire new_net_20686;
	wire new_net_18255;
	wire new_net_9778;
	wire new_net_929;
	wire _0755_;
	wire new_net_1185;
	wire new_net_10881;
	wire new_net_8232;
	wire new_net_9694;
	wire new_net_11269;
	wire new_net_3165;
	wire new_net_1620;
	wire new_net_9371;
	wire new_net_19967;
	wire new_net_7494;
	wire new_net_16439;
	wire _0756_;
	wire new_net_737;
	wire new_net_1622;
	wire new_net_3181;
	wire new_net_14669;
	wire new_net_13435;
	wire new_net_12348;
	wire new_net_13859;
	wire new_net_18037;
	wire new_net_21073;
	wire new_net_4239;
	wire new_net_5021;
	wire new_net_8741;
	wire new_net_9374;
	wire new_net_5535;
	wire new_net_2761;
	wire new_net_18832;
	wire _0757_;
	wire new_net_734;
	wire new_net_1188;
	wire new_net_5366;
	wire new_net_11660;
	wire new_net_3178;
	wire new_net_19419;
	wire new_net_10623;
	wire new_net_348;
	wire new_net_3336;
	wire new_net_3172;
	wire new_net_3701;
	wire new_net_8734;
	wire new_net_9793;
	wire new_net_18765;
	wire new_net_18333;
	wire new_net_19476;
	wire _0758_;
	wire new_net_3164;
	wire new_net_8735;
	wire new_net_8836;
	wire new_net_20687;
	wire new_net_21231;
	wire new_net_1193;
	wire new_net_11270;
	wire new_net_10882;
	wire new_net_8756;
	wire new_net_7238;
	wire new_net_19472;
	wire _0759_;
	wire new_net_4616;
	wire new_net_8837;
	wire new_net_10631;
	wire new_net_5534;
	wire new_net_8224;
	wire new_net_5020;
	wire new_net_19968;
	wire _1750_;
	wire new_net_20359;
	wire new_net_17007;
	wire new_net_12349;
	wire new_net_16440;
	wire new_net_220;
	wire new_net_518;
	wire new_net_16274;
	wire new_net_14154;
	wire new_net_14670;
	wire new_net_16015;
	wire new_net_17445;
	wire new_net_18920;
	wire _0760_;
	wire new_net_516;
	wire new_net_8743;
	wire new_net_735;
	wire new_net_4241;
	wire new_net_20314;
	wire new_net_740;
	wire new_net_5026;
	wire new_net_11659;
	wire new_net_9533;
	wire new_net_9685;
	wire new_net_19420;
	wire new_net_20020;
	wire new_net_20310;
	wire new_net_8746;
	wire new_net_9781;
	wire new_net_923;
	wire _0761_;
	wire new_net_3162;
	wire new_net_9534;
	wire new_net_18483;
	wire new_net_21416;
	wire new_net_18555;
	wire new_net_19798;
	wire new_net_521;
	wire new_net_8234;
	wire new_net_20688;
	wire new_net_842;
	wire new_net_18521;
	wire new_net_10883;
	wire new_net_9375;
	wire _0762_;
	wire new_net_8225;
	wire new_net_15199;
	wire new_net_4238;
	wire new_net_9789;
	wire new_net_11271;
	wire new_net_14957;
	wire new_net_19475;
	wire new_net_513;
	wire new_net_7081;
	wire new_net_19969;
	wire new_net_20023;
	wire _0441_;
	wire new_net_14155;
	wire new_net_16016;
	wire new_net_17446;
	wire new_net_1615;
	wire _0763_;
	wire new_net_921;
	wire new_net_16441;
	wire new_net_3499;
	wire new_net_14671;
	wire new_net_17008;
	wire new_net_21097;
	wire new_net_520;
	wire new_net_9780;
	wire new_net_5536;
	wire new_net_21227;
	wire _0764_;
	wire new_net_3166;
	wire new_net_11658;
	wire new_net_4236;
	wire new_net_19421;
	wire new_net_20235;
	wire new_net_21229;
	wire new_net_916;
	wire new_net_3385;
	wire new_net_8738;
	wire new_net_10632;
	wire new_net_19473;
	wire new_net_21417;
	wire _0765_;
	wire new_net_3176;
	wire new_net_9784;
	wire new_net_9787;
	wire new_net_20689;
	wire new_net_517;
	wire new_net_3169;
	wire new_net_4614;
	wire new_net_9777;
	wire new_net_10624;
	wire new_net_10884;
	wire new_net_7235;
	wire new_net_9691;
	wire new_net_9786;
	wire new_net_11272;
	wire new_net_18167;
	wire _0766_;
	wire new_net_3496;
	wire new_net_8752;
	wire new_net_9794;
	wire new_net_19970;
	wire new_net_20019;
	wire new_net_18074;
	wire new_net_21176;
	wire new_net_14156;
	wire new_net_16017;
	wire new_net_17447;
	wire new_net_3331;
	wire new_net_3704;
	wire new_net_7232;
	wire new_net_9779;
	wire new_net_16442;
	wire new_net_11656;
	wire new_net_14672;
	wire new_net_18786;
	wire new_net_19678;
	wire _0767_;
	wire new_net_739;
	wire new_net_3179;
	wire new_net_7490;
	wire new_net_18063;
	wire new_net_20022;
	wire new_net_3497;
	wire new_net_6801;
	wire new_net_8755;
	wire new_net_9796;
	wire new_net_11657;
	wire new_net_19422;
	wire new_net_17280;
	wire new_net_19027;
	wire new_net_221;
	wire new_net_733;
	wire _0768_;
	wire new_net_9380;
	wire new_net_21418;
	wire new_net_19640;
	wire new_net_1191;
	wire new_net_3492;
	wire new_net_8754;
	wire new_net_7234;
	wire new_net_9791;
	wire new_net_20690;
	wire new_net_19626;
	wire _0769_;
	wire new_net_349;
	wire new_net_10885;
	wire new_net_9688;
	wire new_net_21228;
	wire _0308_;
	wire new_net_611;
	wire new_net_2841;
	wire new_net_4759;
	wire new_net_10349;
	wire new_net_6091;
	wire new_net_8670;
	wire new_net_20159;
	wire new_net_20535;
	wire new_net_503;
	wire new_net_13203;
	wire new_net_2016;
	wire _0266_;
	wire _1400_;
	wire _1610_;
	wire new_net_16348;
	wire new_net_16526;
	wire new_net_11736;
	wire new_net_11773;
	wire new_net_12849;
	wire new_net_2269;
	wire new_net_606;
	wire new_net_5765;
	wire new_net_6885;
	wire new_net_11677;
	wire _0938_;
	wire new_net_18337;
	wire new_net_9811;
	wire _1401_;
	wire _1611_;
	wire new_net_2838;
	wire _0267_;
	wire new_net_3599;
	wire new_net_4693;
	wire new_net_7858;
	wire new_net_6088;
	wire new_net_2845;
	wire new_net_5260;
	wire new_net_5902;
	wire new_net_7863;
	wire new_net_18256;
	wire new_net_1554;
	wire new_net_3624;
	wire _1402_;
	wire _1612_;
	wire _0268_;
	wire new_net_1269;
	wire new_net_9812;
	wire new_net_20158;
	wire new_net_2123;
	wire new_net_10552;
	wire new_net_183;
	wire new_net_11737;
	wire new_net_8759;
	wire new_net_13909;
	wire new_net_11099;
	wire new_net_11365;
	wire new_net_17980;
	wire new_net_20394;
	wire _1403_;
	wire _1613_;
	wire new_net_2025;
	wire _0269_;
	wire new_net_604;
	wire new_net_9808;
	wire new_net_20536;
	wire new_net_18038;
	wire new_net_14874;
	wire new_net_4288;
	wire new_net_16171;
	wire new_net_7456;
	wire new_net_17626;
	wire new_net_12850;
	wire new_net_11735;
	wire new_net_11774;
	wire new_net_16527;
	wire new_net_16349;
	wire new_net_18833;
	wire _1404_;
	wire _1614_;
	wire _0270_;
	wire new_net_6081;
	wire new_net_5760;
	wire _0714_;
	wire new_net_19445;
	wire new_net_18766;
	wire new_net_18334;
	wire new_net_10555;
	wire _1405_;
	wire _1615_;
	wire new_net_683;
	wire _0271_;
	wire new_net_16667;
	wire new_net_1271;
	wire new_net_5261;
	wire new_net_20845;
	wire new_net_2849;
	wire new_net_325;
	wire new_net_608;
	wire new_net_3598;
	wire new_net_19345;
	wire _1406_;
	wire _1616_;
	wire new_net_2017;
	wire _0272_;
	wire new_net_2850;
	wire new_net_12034;
	wire new_net_8495;
	wire new_net_8757;
	wire new_net_11100;
	wire new_net_11366;
	wire new_net_3625;
	wire new_net_8492;
	wire new_net_20537;
	wire new_net_18921;
	wire _1407_;
	wire _1617_;
	wire new_net_680;
	wire new_net_2843;
	wire _0273_;
	wire new_net_7457;
	wire new_net_16350;
	wire new_net_11734;
	wire new_net_16528;
	wire new_net_11775;
	wire new_net_2024;
	wire new_net_2837;
	wire new_net_4768;
	wire new_net_9556;
	wire new_net_13908;
	wire new_net_18484;
	wire new_net_7995;
	wire _1408_;
	wire _1618_;
	wire _0274_;
	wire new_net_16666;
	wire new_net_6084;
	wire new_net_21023;
	wire new_net_18556;
	wire new_net_4289;
	wire new_net_4758;
	wire new_net_5268;
	wire new_net_18522;
	wire new_net_20844;
	wire new_net_18457;
	wire new_net_20908;
	wire new_net_2669;
	wire _1409_;
	wire _1619_;
	wire new_net_682;
	wire _0275_;
	wire new_net_4293;
	wire new_net_11101;
	wire new_net_3632;
	wire new_net_5899;
	wire new_net_11367;
	wire _0276_;
	wire _1410_;
	wire _1620_;
	wire new_net_3594;
	wire new_net_17978;
	wire new_net_20538;
	wire new_net_20843;
	wire new_net_21098;
	wire new_net_14876;
	wire new_net_4762;
	wire new_net_5901;
	wire new_net_11733;
	wire new_net_16529;
	wire new_net_11776;
	wire new_net_12035;
	wire new_net_13206;
	wire new_net_17628;
	wire new_net_12852;
	wire new_net_328;
	wire _1411_;
	wire _1621_;
	wire _0277_;
	wire new_net_13907;
	wire new_net_20236;
	wire new_net_18691;
	wire new_net_8000;
	wire new_net_8493;
	wire _0917_;
	wire _0278_;
	wire _1412_;
	wire new_net_3628;
	wire _1622_;
	wire new_net_6886;
	wire new_net_2018;
	wire new_net_185;
	wire new_net_13906;
	wire new_net_5262;
	wire new_net_609;
	wire new_net_2844;
	wire new_net_20157;
	wire new_net_20842;
	wire new_net_18168;
	wire new_net_11102;
	wire new_net_11368;
	wire _0279_;
	wire _1413_;
	wire _1623_;
	wire new_net_2840;
	wire new_net_16664;
	wire new_net_17977;
	wire new_net_18075;
	wire new_net_4761;
	wire new_net_7999;
	wire new_net_9806;
	wire new_net_7855;
	wire new_net_20539;
	wire new_net_18787;
	wire new_net_19679;
	wire new_net_5767;
	wire new_net_14877;
	wire new_net_17629;
	wire _0280_;
	wire _1414_;
	wire _1624_;
	wire new_net_9807;
	wire new_net_4763;
	wire new_net_16352;
	wire new_net_11732;
	wire new_net_1273;
	wire new_net_178;
	wire new_net_331;
	wire new_net_2021;
	wire new_net_9810;
	wire new_net_16659;
	wire new_net_8661;
	wire new_net_16588;
	wire new_net_14393;
	wire new_net_20787;
	wire new_net_19028;
	wire new_net_11308;
	wire _0281_;
	wire new_net_329;
	wire new_net_1268;
	wire _1415_;
	wire _1625_;
	wire new_net_9552;
	wire new_net_6086;
	wire new_net_10346;
	wire new_net_20836;
	wire new_net_19641;
	wire new_net_687;
	wire new_net_5764;
	wire new_net_6884;
	wire new_net_16665;
	wire _0282_;
	wire new_net_1424;
	wire _1626_;
	wire new_net_2023;
	wire new_net_4291;
	wire new_net_7856;
	wire _1416_;
	wire new_net_6087;
	wire new_net_20156;
	wire new_net_16364;
	wire new_net_11103;
	wire new_net_11369;
	wire new_net_3592;
	wire new_net_3629;
	wire new_net_5761;
	wire new_net_20151;
	wire new_net_612;
	wire _0283_;
	wire _1417_;
	wire _1627_;
	wire new_net_7996;
	wire new_net_6882;
	wire new_net_3365;
	wire new_net_16293;
	wire new_net_2015;
	wire new_net_2842;
	wire new_net_14878;
	wire new_net_17630;
	wire new_net_177;
	wire new_net_605;
	wire new_net_4691;
	wire new_net_5075;
	wire new_net_10556;
	wire new_net_16353;
	wire new_net_11731;
	wire new_net_16531;
	wire new_net_5265;
	wire _1418_;
	wire _1628_;
	wire new_net_186;
	wire new_net_8001;
	wire _0284_;
	wire new_net_3591;
	wire new_net_18418;
	wire new_net_18338;
	wire new_net_2350;
	wire new_net_19826;
	wire new_net_5072;
	wire new_net_8669;
	wire new_net_686;
	wire new_net_20153;
	wire new_net_5077;
	wire _1419_;
	wire _1629_;
	wire new_net_2846;
	wire new_net_332;
	wire new_net_1267;
	wire _0285_;
	wire new_net_7862;
	wire new_net_18257;
	wire new_net_10348;
	wire new_net_180;
	wire new_net_9549;
	wire new_net_9813;
	wire new_net_11104;
	wire new_net_11370;
	wire _1420_;
	wire _1630_;
	wire new_net_182;
	wire new_net_684;
	wire _0286_;
	wire new_net_1415;
	wire new_net_4766;
	wire new_net_5758;
	wire new_net_7857;
	wire new_net_20541;
	wire new_net_21253;
	wire new_net_18039;
	wire new_net_14750;
	wire new_net_16176;
	wire new_net_14879;
	wire new_net_17631;
	wire _1421_;
	wire _1631_;
	wire _0287_;
	wire new_net_7998;
	wire new_net_9551;
	wire new_net_16354;
	wire new_net_13905;
	wire new_net_3289;
	wire new_net_4294;
	wire new_net_5696;
	wire new_net_6089;
	wire new_net_16658;
	wire new_net_17974;
	wire new_net_18834;
	wire new_net_20148;
	wire new_net_17002;
	wire _1422_;
	wire _1632_;
	wire new_net_324;
	wire _0288_;
	wire new_net_5903;
	wire new_net_18767;
	wire new_net_18335;
	wire new_net_3627;
	wire new_net_20152;
	wire new_net_4912;
	wire new_net_8666;
	wire new_net_10342;
	wire _1423_;
	wire _1633_;
	wire _0289_;
	wire new_net_5263;
	wire new_net_5763;
	wire new_net_20841;
	wire new_net_685;
	wire new_net_1423;
	wire new_net_3631;
	wire new_net_4692;
	wire new_net_4911;
	wire new_net_11105;
	wire new_net_11371;
	wire new_net_9550;
	wire new_net_6883;
	wire new_net_7459;
	wire _1757_;
	wire new_net_6083;
	wire _1424_;
	wire _1634_;
	wire new_net_681;
	wire new_net_1274;
	wire new_net_10553;
	wire _0290_;
	wire new_net_1426;
	wire new_net_16656;
	wire new_net_20542;
	wire new_net_8664;
	wire new_net_14751;
	wire new_net_16177;
	wire new_net_1417;
	wire new_net_5073;
	wire new_net_6887;
	wire new_net_14880;
	wire new_net_17632;
	wire new_net_16355;
	wire new_net_11729;
	wire new_net_18922;
	wire new_net_5694;
	wire new_net_13904;
	wire _1425_;
	wire _1635_;
	wire _0291_;
	wire new_net_333;
	wire new_net_10550;
	wire new_net_6889;
	wire new_net_7859;
	wire new_net_4688;
	wire new_net_9555;
	wire new_net_11635;
	wire new_net_18485;
	wire new_net_18557;
	wire new_net_5074;
	wire _1426_;
	wire _1636_;
	wire new_net_181;
	wire new_net_2020;
	wire _0292_;
	wire new_net_1270;
	wire new_net_10549;
	wire new_net_4689;
	wire new_net_15580;
	wire new_net_18194;
	wire new_net_18523;
	wire new_net_614;
	wire new_net_678;
	wire new_net_5259;
	wire new_net_16663;
	wire new_net_5695;
	wire _1427_;
	wire _1637_;
	wire _0293_;
	wire new_net_5070;
	wire new_net_5762;
	wire new_net_11106;
	wire new_net_11372;
	wire new_net_9548;
	wire new_net_17973;
	wire new_net_1539;
	wire new_net_3286;
	wire new_net_5759;
	wire new_net_6090;
	wire new_net_6888;
	wire new_net_20543;
	wire new_net_20840;
	wire new_net_21099;
	wire new_net_16710;
	wire new_net_12857;
	wire new_net_14752;
	wire new_net_16178;
	wire _1428_;
	wire _1638_;
	wire new_net_2848;
	wire _0294_;
	wire new_net_14881;
	wire new_net_17633;
	wire new_net_9557;
	wire new_net_13903;
	wire new_net_2019;
	wire new_net_607;
	wire new_net_5264;
	wire new_net_19343;
	wire new_net_17910;
	wire new_net_19008;
	wire new_net_18692;
	wire new_net_4913;
	wire new_net_326;
	wire new_net_1263;
	wire new_net_1420;
	wire _1429_;
	wire _1639_;
	wire _0295_;
	wire new_net_15740;
	wire new_net_4292;
	wire new_net_8662;
	wire new_net_10345;
	wire new_net_1422;
	wire new_net_187;
	wire new_net_1264;
	wire new_net_3370;
	wire new_net_7993;
	wire new_net_8665;
	wire _1430_;
	wire _1640_;
	wire _0296_;
	wire new_net_5904;
	wire new_net_20155;
	wire new_net_20838;
	wire new_net_18169;
	wire new_net_8761;
	wire new_net_3285;
	wire new_net_11107;
	wire new_net_11373;
	wire new_net_4690;
	wire new_net_17972;
	wire new_net_4914;
	wire _1431_;
	wire _1641_;
	wire _0297_;
	wire new_net_4290;
	wire new_net_7997;
	wire new_net_16657;
	wire new_net_20544;
	wire new_net_20839;
	wire new_net_18788;
	wire new_net_19680;
	wire new_net_12858;
	wire new_net_8663;
	wire new_net_14753;
	wire new_net_16179;
	wire new_net_334;
	wire new_net_610;
	wire new_net_4760;
	wire new_net_14882;
	wire new_net_17634;
	wire new_net_16357;
	wire new_net_13902;
	wire _0298_;
	wire new_net_1266;
	wire _1432_;
	wire _1642_;
	wire new_net_5766;
	wire new_net_3600;
	wire new_net_15280;
	wire new_net_330;
	wire new_net_1418;
	wire new_net_16661;
	wire new_net_19029;
	wire new_net_327;
	wire _0299_;
	wire _1433_;
	wire _1643_;
	wire new_net_9553;
	wire new_net_615;
	wire new_net_3630;
	wire new_net_8494;
	wire new_net_4359;
	wire _0300_;
	wire _1434_;
	wire _1644_;
	wire new_net_11108;
	wire new_net_11374;
	wire new_net_10554;
	wire new_net_9558;
	wire new_net_4764;
	wire new_net_7458;
	wire new_net_2637;
	wire new_net_184;
	wire new_net_679;
	wire new_net_8667;
	wire new_net_20545;
	wire _0315_;
	wire new_net_11783;
	wire new_net_12042;
	wire new_net_13213;
	wire new_net_12859;
	wire _1435_;
	wire _1645_;
	wire new_net_179;
	wire _0301_;
	wire new_net_10341;
	wire new_net_14754;
	wire new_net_1146;
	wire new_net_2847;
	wire new_net_1425;
	wire new_net_3371;
	wire new_net_5076;
	wire new_net_13901;
	wire new_net_18419;
	wire _0945_;
	wire new_net_18339;
	wire new_net_4287;
	wire _1436_;
	wire _1646_;
	wire new_net_2022;
	wire new_net_8668;
	wire new_net_8758;
	wire new_net_10347;
	wire new_net_3626;
	wire new_net_7994;
	wire _0302_;
	wire new_net_1265;
	wire new_net_3595;
	wire new_net_4694;
	wire new_net_7455;
	wire new_net_20154;
	wire new_net_18703;
	wire new_net_18258;
	wire _1437_;
	wire _1647_;
	wire new_net_1419;
	wire new_net_13899;
	wire new_net_5267;
	wire _0303_;
	wire new_net_9547;
	wire new_net_3596;
	wire new_net_10340;
	wire new_net_10551;
	wire new_net_11109;
	wire new_net_11375;
	wire new_net_20150;
	wire _1438_;
	wire _1648_;
	wire new_net_5069;
	wire new_net_6085;
	wire new_net_1416;
	wire _0304_;
	wire new_net_4695;
	wire new_net_20546;
	wire new_net_18040;
	wire new_net_11784;
	wire new_net_12043;
	wire new_net_13214;
	wire new_net_12860;
	wire new_net_2839;
	wire new_net_3373;
	wire new_net_3593;
	wire new_net_10344;
	wire new_net_14755;
	wire new_net_16181;
	wire _1439_;
	wire _1649_;
	wire _0305_;
	wire new_net_5693;
	wire new_net_13900;
	wire new_net_17969;
	wire new_net_20837;
	wire new_net_18835;
	wire _0721_;
	wire new_net_19342;
	wire new_net_18768;
	wire new_net_19180;
	wire new_net_18336;
	wire new_net_5900;
	wire _1440_;
	wire _1650_;
	wire new_net_613;
	wire _0306_;
	wire new_net_3451;
	wire new_net_16660;
	wire new_net_7860;
	wire new_net_9809;
	wire new_net_1421;
	wire new_net_6082;
	wire new_net_9554;
	wire new_net_11110;
	wire new_net_1272;
	wire _1651_;
	wire _1441_;
	wire _0307_;
	wire new_net_3287;
	wire new_net_11376;
	wire new_net_10343;
	wire new_net_5769;
	wire new_net_18923;
	wire new_net_8075;
	wire new_net_238;
	wire new_net_987;
	wire new_net_2151;
	wire new_net_2906;
	wire new_net_10370;
	wire new_net_8316;
	wire new_net_5227;
	wire new_net_5623;
	wire new_net_6182;
	wire new_net_15746;
	wire new_net_3066;
	wire new_net_8077;
	wire new_net_12826;
	wire new_net_15284;
	wire new_net_17045;
	wire new_net_981;
	wire new_net_550;
	wire new_net_12374;
	wire new_net_15154;
	wire new_net_240;
	wire new_net_538;
	wire new_net_984;
	wire new_net_10154;
	wire new_net_10391;
	wire new_net_18486;
	wire new_net_6076;
	wire new_net_16180;
	wire new_net_18558;
	wire new_net_20978;
	wire new_net_18195;
	wire new_net_8190;
	wire new_net_979;
	wire new_net_1199;
	wire new_net_1787;
	wire new_net_1978;
	wire new_net_6252;
	wire new_net_10372;
	wire new_net_8473;
	wire new_net_6972;
	wire new_net_6174;
	wire new_net_18524;
	wire new_net_245;
	wire new_net_436;
	wire new_net_7058;
	wire new_net_8469;
	wire new_net_21202;
	wire new_net_21455;
	wire new_net_8678;
	wire new_net_5980;
	wire new_net_7212;
	wire new_net_10151;
	wire new_net_18181;
	wire new_net_20939;
	wire new_net_11762;
	wire new_net_243;
	wire new_net_980;
	wire new_net_4947;
	wire new_net_6179;
	wire new_net_8317;
	wire new_net_8420;
	wire new_net_11531;
	wire new_net_8470;
	wire new_net_15001;
	wire new_net_21100;
	wire new_net_8374;
	wire new_net_239;
	wire new_net_1200;
	wire new_net_1786;
	wire new_net_6248;
	wire new_net_8323;
	wire new_net_5224;
	wire new_net_6971;
	wire new_net_10392;
	wire new_net_1170;
	wire new_net_18925;
	wire new_net_8380;
	wire new_net_8427;
	wire new_net_8963;
	wire new_net_10580;
	wire new_net_15747;
	wire new_net_437;
	wire new_net_523;
	wire new_net_12827;
	wire new_net_15285;
	wire new_net_17046;
	wire new_net_17911;
	wire new_net_19009;
	wire new_net_18693;
	wire new_net_5979;
	wire new_net_426;
	wire new_net_535;
	wire new_net_1796;
	wire new_net_15000;
	wire new_net_6969;
	wire new_net_7711;
	wire new_net_18179;
	wire _0924_;
	wire new_net_8680;
	wire new_net_8966;
	wire new_net_541;
	wire new_net_3481;
	wire new_net_16300;
	wire new_net_3986;
	wire new_net_18180;
	wire new_net_21203;
	wire new_net_21456;
	wire new_net_8185;
	wire new_net_1970;
	wire new_net_8034;
	wire new_net_7697;
	wire new_net_5225;
	wire new_net_7707;
	wire new_net_20940;
	wire new_net_9032;
	wire new_net_543;
	wire new_net_2905;
	wire new_net_3055;
	wire new_net_11532;
	wire new_net_524;
	wire new_net_6970;
	wire new_net_11229;
	wire new_net_10887;
	wire new_net_20860;
	wire new_net_18789;
	wire new_net_19681;
	wire new_net_5489;
	wire new_net_9035;
	wire new_net_533;
	wire new_net_16132;
	wire new_net_7213;
	wire new_net_20800;
	wire new_net_8685;
	wire new_net_8964;
	wire new_net_11763;
	wire new_net_15748;
	wire new_net_545;
	wire new_net_2152;
	wire new_net_1789;
	wire new_net_12828;
	wire new_net_15286;
	wire new_net_17047;
	wire new_net_16590;
	wire new_net_15279;
	wire new_net_19030;
	wire new_net_3062;
	wire new_net_8320;
	wire new_net_8471;
	wire new_net_10158;
	wire new_net_14999;
	wire new_net_19643;
	wire new_net_2902;
	wire new_net_982;
	wire new_net_1797;
	wire new_net_3374;
	wire new_net_10368;
	wire new_net_5626;
	wire new_net_7713;
	wire new_net_10750;
	wire new_net_8961;
	wire new_net_2904;
	wire new_net_6244;
	wire new_net_21204;
	wire new_net_21457;
	wire new_net_18182;
	wire new_net_1582;
	wire new_net_16292;
	wire new_net_525;
	wire new_net_1788;
	wire new_net_3060;
	wire new_net_7216;
	wire new_net_20941;
	wire new_net_10888;
	wire new_net_534;
	wire new_net_3483;
	wire new_net_4267;
	wire new_net_8033;
	wire new_net_6247;
	wire new_net_11533;
	wire new_net_6223;
	wire new_net_6479;
	wire new_net_7013;
	wire new_net_8371;
	wire new_net_8422;
	wire new_net_10574;
	wire new_net_427;
	wire new_net_1198;
	wire new_net_7698;
	wire new_net_16131;
	wire new_net_10157;
	wire new_net_14183;
	wire new_net_15974;
	wire new_net_5487;
	wire new_net_8425;
	wire new_net_11764;
	wire new_net_15749;
	wire new_net_549;
	wire new_net_978;
	wire new_net_3071;
	wire new_net_12829;
	wire new_net_18420;
	wire new_net_18340;
	wire new_net_4945;
	wire new_net_435;
	wire new_net_1976;
	wire new_net_8072;
	wire new_net_10366;
	wire new_net_14998;
	wire new_net_6974;
	wire new_net_16299;
	wire new_net_8965;
	wire new_net_3375;
	wire new_net_7016;
	wire new_net_8322;
	wire new_net_6184;
	wire new_net_7219;
	wire new_net_18704;
	wire new_net_18259;
	wire new_net_428;
	wire new_net_10394;
	wire new_net_18176;
	wire new_net_21205;
	wire new_net_21458;
	wire new_net_5976;
	wire new_net_244;
	wire new_net_3067;
	wire new_net_3983;
	wire new_net_20942;
	wire new_net_10889;
	wire new_net_16290;
	wire new_net_8189;
	wire new_net_9219;
	wire new_net_11534;
	wire new_net_11231;
	wire new_net_20862;
	wire new_net_546;
	wire new_net_5494;
	wire new_net_16130;
	wire new_net_17049;
	wire new_net_10747;
	wire new_net_14184;
	wire new_net_15158;
	wire new_net_1973;
	wire new_net_11765;
	wire new_net_15750;
	wire new_net_8080;
	wire new_net_12830;
	wire new_net_12378;
	wire new_net_18836;
	wire new_net_9218;
	wire new_net_8186;
	wire new_net_1771;
	wire new_net_539;
	wire new_net_3072;
	wire new_net_7694;
	wire new_net_8464;
	wire new_net_10364;
	wire new_net_8381;
	wire new_net_6177;
	wire new_net_18769;
	wire new_net_4264;
	wire new_net_236;
	wire new_net_8423;
	wire new_net_3057;
	wire new_net_2149;
	wire new_net_2908;
	wire new_net_3980;
	wire new_net_4261;
	wire new_net_18175;
	wire new_net_21206;
	wire new_net_21459;
	wire new_net_10581;
	wire new_net_1794;
	wire new_net_542;
	wire new_net_3061;
	wire new_net_3480;
	wire new_net_4946;
	wire new_net_10363;
	wire new_net_7696;
	wire new_net_6977;
	wire new_net_10153;
	wire _1764_;
	wire new_net_10753;
	wire new_net_10890;
	wire new_net_8967;
	wire new_net_526;
	wire new_net_3376;
	wire new_net_4944;
	wire new_net_6246;
	wire new_net_11535;
	wire new_net_11232;
	wire new_net_6181;
	wire new_net_21215;
	wire new_net_3981;
	wire new_net_4262;
	wire new_net_16129;
	wire new_net_7019;
	wire new_net_10155;
	wire new_net_18924;
	wire new_net_14185;
	wire new_net_15976;
	wire new_net_8377;
	wire new_net_3056;
	wire new_net_5972;
	wire new_net_7214;
	wire new_net_11766;
	wire new_net_15751;
	wire new_net_17050;
	wire new_net_8035;
	wire new_net_10152;
	wire new_net_7689;
	wire new_net_14996;
	wire new_net_12909;
	wire new_net_18487;
	wire new_net_18559;
	wire new_net_19802;
	wire new_net_16298;
	wire new_net_1792;
	wire new_net_7693;
	wire new_net_6975;
	wire new_net_20979;
	wire new_net_18196;
	wire new_net_8426;
	wire new_net_529;
	wire new_net_4948;
	wire new_net_6891;
	wire new_net_21207;
	wire new_net_21460;
	wire new_net_7706;
	wire new_net_10744;
	wire new_net_3076;
	wire new_net_1205;
	wire new_net_7054;
	wire new_net_5228;
	wire new_net_18177;
	wire new_net_20944;
	wire _0455_;
	wire new_net_11536;
	wire new_net_10891;
	wire new_net_540;
	wire new_net_11233;
	wire new_net_5230;
	wire new_net_9034;
	wire new_net_10369;
	wire new_net_8373;
	wire new_net_20864;
	wire new_net_21101;
	wire new_net_247;
	wire new_net_5486;
	wire new_net_5974;
	wire new_net_16128;
	wire new_net_6976;
	wire new_net_18926;
	wire new_net_7220;
	wire new_net_15290;
	wire new_net_12380;
	wire new_net_11767;
	wire new_net_14186;
	wire new_net_1975;
	wire new_net_2147;
	wire new_net_527;
	wire new_net_15977;
	wire new_net_12926;
	wire new_net_20239;
	wire new_net_17912;
	wire new_net_19010;
	wire new_net_6176;
	wire new_net_8682;
	wire new_net_431;
	wire new_net_8191;
	wire new_net_14995;
	wire new_net_18694;
	wire _1176_;
	wire new_net_7714;
	wire new_net_10749;
	wire new_net_1793;
	wire new_net_1972;
	wire new_net_4266;
	wire new_net_8379;
	wire new_net_7014;
	wire new_net_20763;
	wire new_net_237;
	wire new_net_544;
	wire new_net_1770;
	wire new_net_3985;
	wire new_net_7691;
	wire new_net_7055;
	wire new_net_21208;
	wire new_net_21461;
	wire new_net_9033;
	wire new_net_7017;
	wire new_net_20945;
	wire new_net_21254;
	wire new_net_10892;
	wire new_net_249;
	wire new_net_1204;
	wire new_net_3070;
	wire new_net_5488;
	wire new_net_5971;
	wire new_net_6251;
	wire new_net_11537;
	wire new_net_7020;
	wire new_net_11234;
	wire new_net_18790;
	wire new_net_433;
	wire new_net_3078;
	wire new_net_10578;
	wire new_net_16127;
	wire new_net_6183;
	wire new_net_14187;
	wire new_net_15978;
	wire new_net_552;
	wire new_net_2907;
	wire new_net_3077;
	wire new_net_8676;
	wire new_net_3979;
	wire new_net_11768;
	wire new_net_15753;
	wire new_net_20769;
	wire new_net_16291;
	wire new_net_2909;
	wire new_net_250;
	wire new_net_17276;
	wire new_net_14994;
	wire new_net_19031;
	wire new_net_16297;
	wire new_net_5492;
	wire new_net_8679;
	wire new_net_18173;
	wire new_net_19644;
	wire new_net_10367;
	wire new_net_434;
	wire new_net_3068;
	wire new_net_4265;
	wire new_net_8372;
	wire new_net_3984;
	wire new_net_9216;
	wire new_net_8324;
	wire new_net_8474;
	wire new_net_21209;
	wire new_net_18183;
	wire new_net_1785;
	wire new_net_1202;
	wire new_net_3378;
	wire new_net_8424;
	wire new_net_7059;
	wire new_net_20946;
	wire new_net_11235;
	wire new_net_7211;
	wire new_net_10893;
	wire new_net_976;
	wire new_net_1197;
	wire new_net_551;
	wire new_net_2154;
	wire new_net_5973;
	wire new_net_10573;
	wire new_net_8074;
	wire new_net_548;
	wire new_net_3063;
	wire new_net_5493;
	wire new_net_10582;
	wire new_net_16126;
	wire new_net_17053;
	wire new_net_6175;
	wire new_net_10745;
	wire new_net_14188;
	wire new_net_15979;
	wire new_net_530;
	wire new_net_3075;
	wire new_net_8375;
	wire new_net_11769;
	wire new_net_15754;
	wire new_net_18421;
	wire _0952_;
	wire new_net_18341;
	wire new_net_10156;
	wire new_net_536;
	wire new_net_2145;
	wire new_net_6242;
	wire new_net_2347;
	wire new_net_9039;
	wire new_net_8319;
	wire new_net_14993;
	wire new_net_18174;
	wire new_net_18750;
	wire new_net_19067;
	wire new_net_18561;
	wire new_net_19007;
	wire new_net_10752;
	wire new_net_7705;
	wire new_net_8073;
	wire new_net_9215;
	wire new_net_19347;
	wire new_net_18705;
	wire new_net_18260;
	wire new_net_8078;
	wire new_net_18170;
	wire new_net_21210;
	wire new_net_21463;
	wire new_net_19565;
	wire new_net_2903;
	wire new_net_3322;
	wire new_net_8421;
	wire new_net_8684;
	wire new_net_9038;
	wire new_net_20947;
	wire new_net_11236;
	wire new_net_7708;
	wire new_net_10894;
	wire new_net_248;
	wire new_net_547;
	wire new_net_2148;
	wire new_net_9217;
	wire new_net_11539;
	wire new_net_8318;
	wire new_net_20867;
	wire new_net_19549;
	wire new_net_6180;
	wire new_net_10159;
	wire new_net_242;
	wire new_net_1784;
	wire new_net_3479;
	wire new_net_5981;
	wire new_net_8960;
	wire new_net_9212;
	wire new_net_16125;
	wire new_net_14189;
	wire new_net_15980;
	wire new_net_2153;
	wire new_net_3320;
	wire new_net_4941;
	wire new_net_11770;
	wire new_net_15755;
	wire new_net_12835;
	wire new_net_15293;
	wire new_net_17054;
	wire new_net_18837;
	wire new_net_17005;
	wire new_net_13858;
	wire new_net_16294;
	wire new_net_2150;
	wire new_net_3065;
	wire new_net_5490;
	wire new_net_3982;
	wire new_net_6245;
	wire new_net_7015;
	wire new_net_14992;
	wire new_net_19444;
	wire new_net_16256;
	wire new_net_18770;
	wire new_net_10743;
	wire new_net_16296;
	wire new_net_1791;
	wire new_net_0;
	wire new_net_3058;
	wire new_net_3073;
	wire new_net_5491;
	wire new_net_8419;
	wire new_net_7018;
	wire new_net_8315;
	wire new_net_5226;
	wire new_net_537;
	wire new_net_2900;
	wire new_net_4268;
	wire new_net_5978;
	wire new_net_21211;
	wire new_net_21464;
	wire new_net_1036;
	wire new_net_7544;
	wire new_net_531;
	wire new_net_3064;
	wire new_net_3079;
	wire new_net_7056;
	wire new_net_8378;
	wire new_net_10575;
	wire new_net_20948;
	wire new_net_11237;
	wire new_net_10393;
	wire new_net_432;
	wire new_net_3482;
	wire new_net_10751;
	wire new_net_10895;
	wire new_net_10577;
	wire new_net_8192;
	wire new_net_9036;
	wire new_net_7699;
	wire new_net_21129;
	wire new_net_7712;
	wire new_net_16124;
	wire new_net_19247;
	wire new_net_7021;
	wire new_net_17658;
	wire new_net_5223;
	wire new_net_553;
	wire new_net_429;
	wire new_net_986;
	wire new_net_14190;
	wire new_net_15981;
	wire new_net_12930;
	wire new_net_10579;
	wire new_net_10395;
	wire new_net_528;
	wire new_net_1974;
	wire new_net_4263;
	wire new_net_8376;
	wire new_net_8681;
	wire new_net_8188;
	wire new_net_18488;
	wire new_net_3069;
	wire new_net_1203;
	wire new_net_8677;
	wire new_net_9040;
	wire new_net_19349;
	wire new_net_20980;
	wire new_net_18197;
	wire new_net_20912;
	wire new_net_983;
	wire new_net_5625;
	wire new_net_8683;
	wire new_net_21212;
	wire new_net_21465;
	wire new_net_8468;
	wire new_net_246;
	wire new_net_1196;
	wire new_net_8418;
	wire new_net_1783;
	wire new_net_15621;
	wire new_net_20949;
	wire new_net_6892;
	wire new_net_11238;
	wire new_net_3074;
	wire new_net_532;
	wire new_net_10896;
	wire new_net_4269;
	wire new_net_12461;
	wire new_net_10365;
	wire new_net_11541;
	wire new_net_16122;
	wire new_net_21102;
	wire new_net_8321;
	wire new_net_5622;
	wire new_net_6178;
	wire new_net_1773;
	wire new_net_1790;
	wire new_net_3478;
	wire new_net_8193;
	wire new_net_16123;
	wire new_net_14991;
	wire new_net_17659;
	wire new_net_7218;
	wire new_net_7710;
	wire new_net_2901;
	wire new_net_3059;
	wire new_net_430;
	wire new_net_1772;
	wire new_net_10746;
	wire new_net_14191;
	wire new_net_17852;
	wire new_net_18927;
	wire new_net_17913;
	wire new_net_19011;
	wire new_net_8465;
	wire new_net_3978;
	wire new_net_18695;
	wire new_net_12132;
	wire _0931_;
	wire new_net_6173;
	wire new_net_241;
	wire new_net_1201;
	wire new_net_1979;
	wire new_net_16295;
	wire new_net_5975;
	wire new_net_10576;
	wire new_net_4942;
	wire new_net_19350;
	wire new_net_17319;
	wire new_net_14018;
	wire new_net_10149;
	wire new_net_2146;
	wire new_net_16289;
	wire new_net_5977;
	wire new_net_8417;
	wire new_net_8959;
	wire new_net_21213;
	wire new_net_21466;
	wire new_net_8467;
	wire new_net_977;
	wire new_net_1971;
	wire new_net_3977;
	wire new_net_9037;
	wire new_net_20950;
	wire new_net_11239;
	wire new_net_985;
	wire new_net_1795;
	wire new_net_1977;
	wire new_net_10897;
	wire new_net_8962;
	wire new_net_4943;
	wire new_net_8076;
	wire new_net_7695;
	wire new_net_11542;
	wire new_net_6844;
	wire new_net_18791;
	wire new_net_5302;
	wire new_net_170;
	wire new_net_20802;
	wire new_net_8460;
	wire new_net_10777;
	wire new_net_1762;
	wire new_net_1882;
	wire new_net_7559;
	wire new_net_20488;
	wire new_net_15935;
	wire new_net_5008;
	wire new_net_8510;
	wire new_net_17555;
	wire new_net_7099;
	wire new_net_14287;
	wire _0854_;
	wire new_net_2341;
	wire new_net_11927;
	wire new_net_13096;
	wire new_net_8197;
	wire new_net_135;
	wire new_net_18995;
	wire new_net_20184;
	wire new_net_20244;
	wire new_net_18112;
	wire new_net_6311;
	wire new_net_877;
	wire _0855_;
	wire new_net_6430;
	wire new_net_3781;
	wire new_net_18231;
	wire new_net_18184;
	wire new_net_6255;
	wire new_net_368;
	wire new_net_463;
	wire new_net_658;
	wire new_net_2343;
	wire new_net_18986;
	wire new_net_16085;
	wire new_net_9521;
	wire _0856_;
	wire new_net_2352;
	wire new_net_2533;
	wire new_net_7558;
	wire new_net_9699;
	wire new_net_7448;
	wire new_net_12565;
	wire new_net_20951;
	wire new_net_6222;
	wire new_net_13416;
	wire new_net_9522;
	wire new_net_11343;
	wire new_net_2865;
	wire new_net_878;
	wire new_net_2535;
	wire new_net_6459;
	wire new_net_13603;
	wire new_net_12210;
	wire new_net_6258;
	wire new_net_464;
	wire new_net_1768;
	wire _0857_;
	wire new_net_9698;
	wire new_net_3782;
	wire new_net_20489;
	wire new_net_12735;
	wire new_net_18422;
	wire new_net_19103;
	wire new_net_18342;
	wire new_net_12969;
	wire new_net_13864;
	wire new_net_5574;
	wire new_net_15047;
	wire new_net_15936;
	wire new_net_17556;
	wire new_net_1881;
	wire new_net_466;
	wire new_net_14288;
	wire new_net_11928;
	wire new_net_18751;
	wire new_net_19068;
	wire new_net_138;
	wire _0858_;
	wire new_net_363;
	wire new_net_9702;
	wire new_net_2339;
	wire new_net_14732;
	wire new_net_20185;
	wire new_net_20245;
	wire new_net_18706;
	wire new_net_18261;
	wire new_net_1765;
	wire new_net_2866;
	wire new_net_369;
	wire new_net_8931;
	wire _0326_;
	wire new_net_19566;
	wire new_net_15483;
	wire new_net_6256;
	wire new_net_2872;
	wire _0859_;
	wire new_net_8194;
	wire new_net_8509;
	wire new_net_10779;
	wire new_net_361;
	wire new_net_6733;
	wire new_net_7146;
	wire new_net_7553;
	wire new_net_20952;
	wire new_net_21024;
	wire new_net_11344;
	wire new_net_656;
	wire _0860_;
	wire new_net_360;
	wire new_net_2346;
	wire new_net_15046;
	wire new_net_139;
	wire new_net_3359;
	wire new_net_8923;
	wire new_net_20490;
	wire new_net_18838;
	wire new_net_15287;
	wire new_net_17006;
	wire new_net_12970;
	wire new_net_13865;
	wire new_net_14476;
	wire new_net_15937;
	wire new_net_17557;
	wire new_net_1766;
	wire _0861_;
	wire new_net_2353;
	wire new_net_14289;
	wire new_net_17308;
	wire new_net_4949;
	wire new_net_16257;
	wire new_net_18771;
	wire new_net_19174;
	wire new_net_10606;
	wire new_net_8454;
	wire new_net_10778;
	wire new_net_14731;
	wire new_net_20186;
	wire new_net_20246;
	wire new_net_8511;
	wire new_net_2861;
	wire _0862_;
	wire new_net_7447;
	wire new_net_18232;
	wire new_net_5467;
	wire _1771_;
	wire new_net_21130;
	wire new_net_4919;
	wire _0863_;
	wire new_net_461;
	wire new_net_655;
	wire new_net_20953;
	wire new_net_21025;
	wire new_net_8196;
	wire new_net_8515;
	wire new_net_11345;
	wire new_net_1769;
	wire new_net_474;
	wire new_net_3778;
	wire new_net_7105;
	wire new_net_19441;
	wire new_net_9740;
	wire new_net_6320;
	wire new_net_15045;
	wire new_net_8200;
	wire new_net_2344;
	wire new_net_140;
	wire new_net_2862;
	wire _0864_;
	wire new_net_3784;
	wire new_net_20491;
	wire new_net_12212;
	wire new_net_15713;
	wire new_net_12971;
	wire new_net_13866;
	wire new_net_15938;
	wire new_net_17558;
	wire new_net_1759;
	wire new_net_5573;
	wire new_net_6432;
	wire new_net_12911;
	wire new_net_14730;
	wire new_net_9525;
	wire new_net_6317;
	wire new_net_136;
	wire new_net_467;
	wire new_net_1760;
	wire _0865_;
	wire new_net_7556;
	wire new_net_20187;
	wire new_net_20247;
	wire new_net_15584;
	wire new_net_18198;
	wire new_net_8195;
	wire new_net_18994;
	wire _0866_;
	wire new_net_7102;
	wire new_net_19297;
	wire _0462_;
	wire new_net_370;
	wire new_net_20954;
	wire new_net_21026;
	wire new_net_20521;
	wire new_net_21103;
	wire new_net_9742;
	wire new_net_465;
	wire new_net_5575;
	wire new_net_6321;
	wire new_net_364;
	wire new_net_2348;
	wire _0867_;
	wire new_net_6259;
	wire new_net_11346;
	wire new_net_1763;
	wire new_net_9518;
	wire new_net_15044;
	wire new_net_20492;
	wire new_net_17853;
	wire new_net_18928;
	wire new_net_13493;
	wire new_net_17914;
	wire new_net_19012;
	wire new_net_12213;
	wire new_net_15714;
	wire new_net_17310;
	wire new_net_12972;
	wire new_net_13867;
	wire new_net_15939;
	wire new_net_2536;
	wire _0868_;
	wire new_net_653;
	wire new_net_16648;
	wire new_net_18572;
	wire new_net_18696;
	wire new_net_15155;
	wire new_net_16133;
	wire new_net_14729;
	wire new_net_6080;
	wire new_net_2534;
	wire new_net_365;
	wire new_net_473;
	wire new_net_3783;
	wire new_net_5680;
	wire new_net_20188;
	wire new_net_20248;
	wire new_net_17320;
	wire new_net_14019;
	wire new_net_2349;
	wire _0869_;
	wire new_net_874;
	wire new_net_7103;
	wire new_net_9701;
	wire new_net_18233;
	wire new_net_17162;
	wire new_net_876;
	wire new_net_2870;
	wire new_net_18230;
	wire new_net_18993;
	wire new_net_21256;
	wire new_net_2340;
	wire _0870_;
	wire new_net_6254;
	wire new_net_20955;
	wire new_net_21027;
	wire new_net_661;
	wire new_net_1764;
	wire new_net_5676;
	wire new_net_6429;
	wire new_net_7452;
	wire new_net_11347;
	wire new_net_8930;
	wire new_net_18376;
	wire new_net_18792;
	wire new_net_7453;
	wire new_net_15043;
	wire _0871_;
	wire new_net_8187;
	wire new_net_20493;
	wire new_net_14397;
	wire new_net_16592;
	wire new_net_12085;
	wire new_net_13597;
	wire new_net_9741;
	wire new_net_12214;
	wire new_net_15715;
	wire new_net_12973;
	wire new_net_13868;
	wire new_net_17311;
	wire new_net_15940;
	wire new_net_468;
	wire new_net_17274;
	wire new_net_14728;
	wire new_net_8459;
	wire new_net_654;
	wire new_net_1873;
	wire _0872_;
	wire new_net_6458;
	wire new_net_20189;
	wire new_net_20249;
	wire new_net_18113;
	wire new_net_1874;
	wire new_net_2351;
	wire new_net_8507;
	wire new_net_7107;
	wire new_net_6428;
	wire new_net_18235;
	wire new_net_18185;
	wire new_net_6738;
	wire new_net_657;
	wire new_net_887;
	wire _0873_;
	wire new_net_7958;
	wire new_net_12529;
	wire new_net_14109;
	wire new_net_16086;
	wire new_net_18992;
	wire new_net_20956;
	wire new_net_21028;
	wire _0329_;
	wire new_net_15982;
	wire new_net_6880;
	wire new_net_9519;
	wire _0874_;
	wire new_net_11348;
	wire new_net_6434;
	wire new_net_13586;
	wire new_net_9748;
	wire new_net_15042;
	wire new_net_20494;
	wire new_net_18423;
	wire new_net_19104;
	wire new_net_12086;
	wire new_net_13596;
	wire new_net_14480;
	wire new_net_3777;
	wire new_net_12215;
	wire new_net_15716;
	wire new_net_17312;
	wire new_net_12974;
	wire new_net_13869;
	wire new_net_15941;
	wire _0959_;
	wire new_net_15764;
	wire new_net_18343;
	wire new_net_18752;
	wire new_net_19069;
	wire new_net_14727;
	wire new_net_3329;
	wire new_net_6079;
	wire new_net_6314;
	wire new_net_6736;
	wire new_net_20190;
	wire new_net_20250;
	wire new_net_18707;
	wire new_net_18262;
	wire new_net_9520;
	wire new_net_1879;
	wire new_net_2869;
	wire _0876_;
	wire new_net_5009;
	wire new_net_7145;
	wire new_net_6071;
	wire new_net_9524;
	wire new_net_6318;
	wire new_net_8932;
	wire new_net_7557;
	wire new_net_2871;
	wire _0877_;
	wire new_net_367;
	wire new_net_5577;
	wire new_net_20957;
	wire new_net_21029;
	wire new_net_7415;
	wire new_net_8462;
	wire new_net_8198;
	wire new_net_11349;
	wire new_net_18991;
	wire _0878_;
	wire new_net_366;
	wire new_net_146;
	wire new_net_875;
	wire new_net_1877;
	wire new_net_2874;
	wire new_net_15041;
	wire new_net_7554;
	wire new_net_20495;
	wire new_net_18839;
	wire new_net_15288;
	wire new_net_12087;
	wire new_net_13595;
	wire new_net_16651;
	wire new_net_9749;
	wire new_net_12216;
	wire new_net_13860;
	wire new_net_12975;
	wire new_net_13870;
	wire new_net_884;
	wire new_net_15942;
	wire new_net_16258;
	wire new_net_6895;
	wire new_net_18772;
	wire new_net_14726;
	wire _0879_;
	wire new_net_8924;
	wire new_net_18238;
	wire new_net_19298;
	wire new_net_20191;
	wire new_net_20251;
	wire new_net_6074;
	wire new_net_4915;
	wire new_net_5578;
	wire new_net_9526;
	wire new_net_5678;
	wire new_net_13942;
	wire new_net_17559;
	wire new_net_5674;
	wire new_net_6735;
	wire new_net_472;
	wire new_net_1758;
	wire new_net_1876;
	wire _0880_;
	wire new_net_8457;
	wire new_net_5010;
	wire new_net_462;
	wire new_net_886;
	wire new_net_4916;
	wire new_net_8461;
	wire new_net_8926;
	wire new_net_19299;
	wire new_net_20958;
	wire new_net_21030;
	wire _0231_;
	wire new_net_21131;
	wire new_net_881;
	wire new_net_1875;
	wire _0881_;
	wire new_net_4922;
	wire new_net_11350;
	wire new_net_8929;
	wire new_net_20768;
	wire new_net_137;
	wire new_net_659;
	wire new_net_7564;
	wire new_net_8201;
	wire new_net_15040;
	wire new_net_18990;
	wire new_net_20496;
	wire new_net_11722;
	wire new_net_13588;
	wire new_net_14657;
	wire new_net_17314;
	wire new_net_12088;
	wire new_net_13594;
	wire new_net_12217;
	wire new_net_15718;
	wire new_net_12976;
	wire new_net_13871;
	wire new_net_14725;
	wire new_net_4917;
	wire new_net_5576;
	wire new_net_7106;
	wire new_net_20192;
	wire new_net_20252;
	wire new_net_15585;
	wire new_net_18199;
	wire new_net_847;
	wire new_net_6435;
	wire new_net_7555;
	wire _0883_;
	wire new_net_145;
	wire new_net_2868;
	wire new_net_6316;
	wire new_net_5005;
	wire new_net_18236;
	wire new_net_9700;
	wire new_net_6072;
	wire new_net_6436;
	wire new_net_7450;
	wire new_net_6073;
	wire new_net_2354;
	wire _0884_;
	wire new_net_5569;
	wire new_net_20959;
	wire new_net_21031;
	wire new_net_21104;
	wire new_net_6427;
	wire new_net_7563;
	wire new_net_11351;
	wire new_net_6879;
	wire new_net_1767;
	wire new_net_471;
	wire new_net_7104;
	wire new_net_6734;
	wire new_net_6878;
	wire _0885_;
	wire new_net_133;
	wire new_net_4921;
	wire new_net_8927;
	wire new_net_20497;
	wire new_net_17854;
	wire new_net_18929;
	wire new_net_20136;
	wire new_net_17915;
	wire new_net_19013;
	wire new_net_14483;
	wire new_net_11723;
	wire new_net_13589;
	wire new_net_14658;
	wire new_net_14142;
	wire new_net_16063;
	wire new_net_12089;
	wire new_net_13872;
	wire new_net_15719;
	wire new_net_17315;
	wire new_net_18573;
	wire new_net_18697;
	wire new_net_15156;
	wire new_net_5675;
	wire new_net_15039;
	wire new_net_14724;
	wire new_net_880;
	wire _0886_;
	wire new_net_2875;
	wire new_net_6257;
	wire new_net_20193;
	wire new_net_20253;
	wire new_net_17321;
	wire new_net_14020;
	wire new_net_9746;
	wire new_net_1880;
	wire new_net_2867;
	wire new_net_6313;
	wire new_net_8925;
	wire _0887_;
	wire new_net_5007;
	wire new_net_6078;
	wire new_net_8513;
	wire new_net_8928;
	wire new_net_18774;
	wire new_net_141;
	wire new_net_7454;
	wire new_net_8512;
	wire new_net_20960;
	wire new_net_21032;
	wire _0888_;
	wire new_net_132;
	wire new_net_663;
	wire new_net_6075;
	wire new_net_8458;
	wire new_net_11352;
	wire new_net_18793;
	wire new_net_1887;
	wire new_net_6730;
	wire new_net_9696;
	wire new_net_20498;
	wire new_net_16593;
	wire new_net_11937;
	wire new_net_13106;
	wire new_net_14143;
	wire new_net_9703;
	wire new_net_6732;
	wire new_net_12090;
	wire new_net_14484;
	wire new_net_14659;
	wire new_net_9744;
	wire new_net_12219;
	wire new_net_17273;
	wire new_net_20513;
	wire new_net_6433;
	wire new_net_7451;
	wire new_net_6731;
	wire new_net_882;
	wire new_net_2345;
	wire new_net_5677;
	wire new_net_14723;
	wire new_net_8922;
	wire new_net_18988;
	wire new_net_20194;
	wire new_net_5580;
	wire new_net_18114;
	wire new_net_2873;
	wire _0890_;
	wire new_net_5679;
	wire new_net_4918;
	wire new_net_8463;
	wire new_net_15857;
	wire new_net_18186;
	wire new_net_8199;
	wire new_net_142;
	wire new_net_469;
	wire new_net_6312;
	wire new_net_7561;
	wire new_net_14145;
	wire new_net_14110;
	wire new_net_3780;
	wire new_net_1878;
	wire new_net_2863;
	wire _0891_;
	wire new_net_8203;
	wire new_net_20961;
	wire new_net_21033;
	wire new_net_2630;
	wire new_net_7560;
	wire new_net_9747;
	wire new_net_134;
	wire new_net_362;
	wire new_net_13418;
	wire new_net_12639;
	wire new_net_5570;
	wire new_net_15037;
	wire new_net_11353;
	wire new_net_506;
	wire new_net_3779;
	wire new_net_9743;
	wire new_net_660;
	wire _0892_;
	wire new_net_12033;
	wire new_net_15038;
	wire new_net_8514;
	wire new_net_18241;
	wire new_net_19301;
	wire new_net_20499;
	wire new_net_18424;
	wire new_net_11938;
	wire new_net_13107;
	wire new_net_14144;
	wire new_net_16065;
	wire new_net_16655;
	wire new_net_11725;
	wire new_net_13591;
	wire new_net_14660;
	wire new_net_12091;
	wire new_net_12220;
	wire new_net_19105;
	wire new_net_15765;
	wire new_net_18344;
	wire new_net_18753;
	wire new_net_19070;
	wire new_net_12418;
	wire new_net_7144;
	wire new_net_7449;
	wire new_net_14722;
	wire new_net_143;
	wire new_net_2864;
	wire _0893_;
	wire new_net_18240;
	wire new_net_20195;
	wire new_net_20255;
	wire new_net_18708;
	wire new_net_18263;
	wire new_net_9745;
	wire new_net_144;
	wire new_net_3326;
	wire new_net_6319;
	wire new_net_6253;
	wire new_net_7101;
	wire new_net_18987;
	wire new_net_9726;
	wire new_net_4925;
	wire _0894_;
	wire new_net_5572;
	wire new_net_5006;
	wire new_net_7100;
	wire new_net_18239;
	wire new_net_475;
	wire new_net_662;
	wire new_net_7108;
	wire new_net_8508;
	wire new_net_20962;
	wire new_net_21034;
	wire new_net_16054;
	wire new_net_16031;
	wire new_net_9695;
	wire new_net_6729;
	wire new_net_14721;
	wire new_net_2342;
	wire _0895_;
	wire new_net_8455;
	wire new_net_3302;
	wire new_net_11354;
	wire new_net_16505;
	wire new_net_18840;
	wire new_net_15289;
	wire new_net_13861;
	wire new_net_14614;
	wire new_net_119;
	wire new_net_1118;
	wire new_net_2253;
	wire new_net_10116;
	wire new_net_19971;
	wire new_net_2032;
	wire new_net_16259;
	wire new_net_18773;
	wire new_net_3797;
	wire new_net_9332;
	wire new_net_11915;
	wire new_net_7797;
	wire new_net_13153;
	wire new_net_16066;
	wire new_net_13567;
	wire new_net_14581;
	wire new_net_16538;
	wire new_net_16939;
	wire new_net_2250;
	wire new_net_2736;
	wire new_net_6481;
	wire new_net_17560;
	wire _0015_;
	wire _0309_;
	wire _0435_;
	wire _1317_;
	wire _1653_;
	wire new_net_114;
	wire new_net_777;
	wire new_net_2248;
	wire new_net_12162;
	wire new_net_2975;
	wire new_net_9335;
	wire new_net_9451;
	wire new_net_7618;
	wire new_net_21132;
	wire new_net_9111;
	wire new_net_16405;
	wire new_net_3801;
	wire new_net_5113;
	wire new_net_7589;
	wire new_net_6653;
	wire _0016_;
	wire _0310_;
	wire _0436_;
	wire _1318_;
	wire _1654_;
	wire new_net_7615;
	wire new_net_13154;
	wire new_net_13568;
	wire new_net_17187;
	wire new_net_1987;
	wire new_net_2255;
	wire new_net_3301;
	wire new_net_4514;
	wire new_net_4709;
	wire new_net_7617;
	wire new_net_13388;
	wire new_net_10118;
	wire new_net_5110;
	wire new_net_7804;
	wire _0017_;
	wire _0311_;
	wire _0437_;
	wire _1319_;
	wire _1655_;
	wire new_net_159;
	wire new_net_19972;
	wire new_net_12913;
	wire new_net_11641;
	wire new_net_19044;
	wire new_net_11916;
	wire new_net_13152;
	wire new_net_13566;
	wire new_net_15108;
	wire new_net_16067;
	wire new_net_17780;
	wire new_net_15771;
	wire new_net_12933;
	wire new_net_16539;
	wire new_net_14970;
	wire new_net_15586;
	wire new_net_18200;
	wire new_net_15094;
	wire new_net_2737;
	wire new_net_5112;
	wire new_net_17186;
	wire _0018_;
	wire _0312_;
	wire new_net_2836;
	wire new_net_2251;
	wire _0438_;
	wire _1320_;
	wire _1656_;
	wire new_net_9339;
	wire new_net_7584;
	wire new_net_5203;
	wire new_net_2254;
	wire new_net_2116;
	wire new_net_2830;
	wire new_net_3802;
	wire new_net_3816;
	wire new_net_7610;
	wire new_net_21326;
	wire _0469_;
	wire _0439_;
	wire _0019_;
	wire _0313_;
	wire _1321_;
	wire _1657_;
	wire new_net_12464;
	wire new_net_149;
	wire new_net_11850;
	wire new_net_4618;
	wire new_net_20220;
	wire new_net_2984;
	wire new_net_3299;
	wire new_net_4623;
	wire new_net_5202;
	wire new_net_12682;
	wire new_net_6229;
	wire new_net_14582;
	wire new_net_5195;
	wire _0020_;
	wire _0314_;
	wire _0440_;
	wire _1322_;
	wire _1658_;
	wire new_net_161;
	wire new_net_9751;
	wire new_net_17855;
	wire new_net_18930;
	wire new_net_13495;
	wire new_net_17916;
	wire new_net_19014;
	wire new_net_9336;
	wire new_net_15306;
	wire new_net_9128;
	wire new_net_19973;
	wire new_net_18574;
	wire new_net_18698;
	wire new_net_15157;
	wire new_net_12135;
	wire new_net_9448;
	wire new_net_11917;
	wire new_net_6476;
	wire new_net_13151;
	wire new_net_16068;
	wire new_net_16231;
	wire new_net_13565;
	wire new_net_16540;
	wire new_net_16941;
	wire new_net_17781;
	wire new_net_17322;
	wire new_net_20767;
	wire new_net_14021;
	wire new_net_17198;
	wire new_net_2624;
	wire new_net_17185;
	wire new_net_18641;
	wire new_net_15456;
	wire new_net_1908;
	wire new_net_4516;
	wire new_net_6225;
	wire new_net_5893;
	wire _0022_;
	wire _0316_;
	wire _0442_;
	wire _1324_;
	wire _1660_;
	wire new_net_1122;
	wire new_net_5566;
	wire new_net_14290;
	wire new_net_4970;
	wire new_net_2977;
	wire new_net_116;
	wire new_net_151;
	wire new_net_13051;
	wire new_net_16377;
	wire new_net_5197;
	wire _0443_;
	wire _0023_;
	wire _0317_;
	wire _1661_;
	wire new_net_3258;
	wire _1325_;
	wire new_net_3817;
	wire new_net_18640;
	wire new_net_18794;
	wire new_net_11184;
	wire new_net_7613;
	wire new_net_11275;
	wire new_net_20805;
	wire new_net_14399;
	wire new_net_16594;
	wire new_net_1990;
	wire new_net_3800;
	wire new_net_2829;
	wire new_net_5200;
	wire _0444_;
	wire _0024_;
	wire _0318_;
	wire new_net_2619;
	wire _1326_;
	wire _1662_;
	wire new_net_12838;
	wire new_net_15274;
	wire new_net_17272;
	wire new_net_15476;
	wire new_net_17072;
	wire new_net_16541;
	wire new_net_15110;
	wire new_net_16942;
	wire new_net_13564;
	wire new_net_16232;
	wire new_net_15335;
	wire new_net_770;
	wire new_net_5565;
	wire new_net_9205;
	wire new_net_18115;
	wire _1663_;
	wire new_net_107;
	wire new_net_1983;
	wire new_net_4907;
	wire _0025_;
	wire _0319_;
	wire _0445_;
	wire new_net_2981;
	wire new_net_2249;
	wire _1327_;
	wire new_net_18187;
	wire new_net_120;
	wire new_net_2252;
	wire new_net_6224;
	wire new_net_9125;
	wire new_net_18639;
	wire new_net_21328;
	wire new_net_14146;
	wire new_net_10122;
	wire _0026_;
	wire _0320_;
	wire _0446_;
	wire _1328_;
	wire _1664_;
	wire new_net_110;
	wire new_net_1115;
	wire new_net_2114;
	wire new_net_5099;
	wire new_net_13146;
	wire _0336_;
	wire new_net_19440;
	wire new_net_19175;
	wire new_net_10119;
	wire new_net_7586;
	wire new_net_2115;
	wire new_net_3821;
	wire new_net_6226;
	wire new_net_19436;
	wire new_net_11276;
	wire _1665_;
	wire _0447_;
	wire _0027_;
	wire _0321_;
	wire new_net_2626;
	wire _1329_;
	wire new_net_20225;
	wire new_net_12738;
	wire new_net_18425;
	wire new_net_7590;
	wire new_net_7798;
	wire new_net_775;
	wire new_net_1986;
	wire new_net_15304;
	wire new_net_19106;
	wire new_net_19975;
	wire new_net_15766;
	wire _0966_;
	wire new_net_18345;
	wire new_net_13785;
	wire new_net_18754;
	wire new_net_19071;
	wire new_net_15477;
	wire _1666_;
	wire new_net_9334;
	wire new_net_11919;
	wire new_net_16070;
	wire new_net_13563;
	wire new_net_14584;
	wire _0448_;
	wire _0028_;
	wire _0322_;
	wire new_net_8048;
	wire new_net_2748;
	wire new_net_18264;
	wire new_net_6480;
	wire new_net_7583;
	wire new_net_157;
	wire new_net_776;
	wire new_net_2617;
	wire new_net_2245;
	wire new_net_3415;
	wire new_net_14612;
	wire new_net_17183;
	wire _1667_;
	wire new_net_10115;
	wire new_net_7585;
	wire new_net_779;
	wire _0449_;
	wire _0029_;
	wire _0323_;
	wire new_net_2834;
	wire _1331_;
	wire new_net_3818;
	wire new_net_16831;
	wire new_net_14263;
	wire new_net_2615;
	wire new_net_3798;
	wire new_net_5897;
	wire new_net_6474;
	wire new_net_9753;
	wire new_net_11185;
	wire new_net_16055;
	wire _1668_;
	wire new_net_774;
	wire _0450_;
	wire _0030_;
	wire _0324_;
	wire _1332_;
	wire new_net_1125;
	wire new_net_3822;
	wire new_net_19446;
	wire new_net_3717;
	wire new_net_11277;
	wire new_net_6227;
	wire new_net_772;
	wire new_net_2621;
	wire new_net_15111;
	wire new_net_20226;
	wire new_net_10641;
	wire new_net_18841;
	wire _1333_;
	wire _1669_;
	wire _0451_;
	wire _0031_;
	wire _0325_;
	wire new_net_160;
	wire new_net_15303;
	wire new_net_19442;
	wire new_net_13862;
	wire new_net_17009;
	wire new_net_2037;
	wire new_net_16260;
	wire new_net_14009;
	wire new_net_14974;
	wire new_net_15337;
	wire new_net_16234;
	wire new_net_15478;
	wire new_net_9338;
	wire new_net_11920;
	wire new_net_16071;
	wire new_net_13149;
	wire new_net_17784;
	wire new_net_7682;
	wire new_net_17182;
	wire new_net_4620;
	wire new_net_3804;
	wire new_net_6477;
	wire new_net_13150;
	wire new_net_17672;
	wire _1334_;
	wire _1670_;
	wire _0452_;
	wire _0032_;
	wire new_net_13944;
	wire new_net_17561;
	wire new_net_9450;
	wire new_net_2978;
	wire new_net_21330;
	wire new_net_3355;
	wire new_net_8951;
	wire new_net_9122;
	wire new_net_9455;
	wire new_net_10121;
	wire _0327_;
	wire _1335_;
	wire _1671_;
	wire new_net_773;
	wire new_net_1991;
	wire _0453_;
	wire _0033_;
	wire new_net_21133;
	wire new_net_16406;
	wire new_net_9453;
	wire new_net_115;
	wire new_net_2620;
	wire new_net_3420;
	wire new_net_11186;
	wire new_net_4622;
	wire new_net_11278;
	wire _1336_;
	wire _1672_;
	wire new_net_1116;
	wire _0454_;
	wire _0034_;
	wire _0328_;
	wire new_net_19439;
	wire new_net_13387;
	wire new_net_7607;
	wire new_net_9127;
	wire new_net_7581;
	wire new_net_15302;
	wire new_net_19977;
	wire new_net_2329;
	wire new_net_11642;
	wire new_net_19045;
	wire new_net_14010;
	wire new_net_14975;
	wire new_net_15112;
	wire new_net_15338;
	wire new_net_15479;
	wire new_net_4515;
	wire new_net_9452;
	wire new_net_11921;
	wire new_net_7587;
	wire new_net_13148;
	wire new_net_15587;
	wire new_net_18201;
	wire new_net_17181;
	wire new_net_6482;
	wire new_net_7588;
	wire new_net_3413;
	wire new_net_4513;
	wire new_net_14610;
	wire new_net_9189;
	wire _0036_;
	wire _0330_;
	wire _0456_;
	wire _1338_;
	wire _1674_;
	wire new_net_2522;
	wire new_net_18638;
	wire new_net_21331;
	wire new_net_15625;
	wire new_net_11851;
	wire new_net_12465;
	wire new_net_10039;
	wire new_net_10355;
	wire new_net_4625;
	wire _0037_;
	wire _0331_;
	wire _0457_;
	wire _1339_;
	wire _1675_;
	wire new_net_2740;
	wire new_net_6647;
	wire new_net_20652;
	wire new_net_12681;
	wire new_net_11187;
	wire new_net_11279;
	wire new_net_2733;
	wire new_net_5198;
	wire new_net_5898;
	wire new_net_17856;
	wire new_net_18931;
	wire new_net_17917;
	wire new_net_19015;
	wire new_net_2117;
	wire new_net_2979;
	wire new_net_3718;
	wire _1676_;
	wire new_net_1981;
	wire new_net_4706;
	wire new_net_7580;
	wire _0038_;
	wire _0332_;
	wire _0458_;
	wire new_net_4278;
	wire new_net_18575;
	wire new_net_18699;
	wire new_net_14011;
	wire new_net_14976;
	wire new_net_15113;
	wire new_net_15339;
	wire new_net_15480;
	wire new_net_11922;
	wire new_net_13147;
	wire new_net_16073;
	wire new_net_12136;
	wire new_net_13560;
	wire new_net_17323;
	wire new_net_20766;
	wire new_net_17180;
	wire _1677_;
	wire new_net_4518;
	wire new_net_14022;
	wire _0039_;
	wire _0333_;
	wire _0459_;
	wire new_net_14609;
	wire _1341_;
	wire new_net_18882;
	wire new_net_3803;
	wire new_net_19355;
	wire new_net_21332;
	wire new_net_15457;
	wire new_net_14291;
	wire new_net_18775;
	wire new_net_9121;
	wire _1678_;
	wire new_net_1980;
	wire new_net_2732;
	wire new_net_7799;
	wire new_net_2833;
	wire _0460_;
	wire _0040_;
	wire _0334_;
	wire new_net_10406;
	wire new_net_21259;
	wire new_net_16378;
	wire new_net_9333;
	wire new_net_18637;
	wire new_net_5303;
	wire new_net_11188;
	wire new_net_11280;
	wire new_net_4520;
	wire new_net_6475;
	wire _0041_;
	wire _0335_;
	wire _0461_;
	wire _1343_;
	wire _1679_;
	wire new_net_1117;
	wire new_net_6643;
	wire new_net_20806;
	wire new_net_14400;
	wire new_net_6228;
	wire new_net_3300;
	wire new_net_3410;
	wire new_net_15300;
	wire new_net_19979;
	wire new_net_12839;
	wire new_net_12153;
	wire new_net_12940;
	wire new_net_14012;
	wire new_net_14977;
	wire new_net_15114;
	wire new_net_15340;
	wire new_net_4619;
	wire new_net_15481;
	wire new_net_11923;
	wire new_net_6230;
	wire new_net_14901;
	wire new_net_18116;
	wire new_net_17179;
	wire new_net_4517;
	wire new_net_4704;
	wire new_net_9123;
	wire new_net_14608;
	wire new_net_17164;
	wire new_net_7803;
	wire new_net_2976;
	wire _0043_;
	wire _0337_;
	wire _0463_;
	wire _1345_;
	wire _1681_;
	wire new_net_111;
	wire new_net_15859;
	wire new_net_1119;
	wire new_net_18188;
	wire new_net_14147;
	wire new_net_20318;
	wire new_net_7614;
	wire new_net_2832;
	wire new_net_154;
	wire new_net_2246;
	wire new_net_5201;
	wire new_net_6650;
	wire new_net_9758;
	wire new_net_12532;
	wire _1682_;
	wire new_net_1985;
	wire new_net_9330;
	wire new_net_5109;
	wire new_net_7802;
	wire _0464_;
	wire _0044_;
	wire _0338_;
	wire _1346_;
	wire new_net_13420;
	wire new_net_13221;
	wire new_net_11189;
	wire new_net_11281;
	wire new_net_9337;
	wire new_net_1123;
	wire new_net_7794;
	wire new_net_16966;
	wire new_net_12739;
	wire new_net_18426;
	wire _1683_;
	wire new_net_106;
	wire new_net_2618;
	wire _0465_;
	wire _0045_;
	wire _0339_;
	wire _1347_;
	wire new_net_1124;
	wire new_net_19248;
	wire new_net_19980;
	wire new_net_19107;
	wire new_net_15767;
	wire new_net_18346;
	wire new_net_18755;
	wire new_net_19072;
	wire new_net_12152;
	wire new_net_12941;
	wire new_net_14013;
	wire new_net_14978;
	wire new_net_15115;
	wire new_net_15341;
	wire new_net_15482;
	wire new_net_9340;
	wire new_net_11924;
	wire new_net_13145;
	wire new_net_13705;
	wire new_net_19146;
	wire new_net_3815;
	wire new_net_5101;
	wire new_net_17178;
	wire _1684_;
	wire new_net_4519;
	wire _0046_;
	wire _0340_;
	wire _0466_;
	wire new_net_6221;
	wire new_net_14607;
	wire new_net_9449;
	wire new_net_2616;
	wire new_net_6644;
	wire new_net_19249;
	wire new_net_21298;
	wire new_net_21334;
	wire new_net_16832;
	wire new_net_17590;
	wire _1685_;
	wire new_net_4708;
	wire new_net_9454;
	wire _0047_;
	wire _0341_;
	wire new_net_2980;
	wire _0467_;
	wire _1349_;
	wire new_net_16056;
	wire new_net_4705;
	wire new_net_109;
	wire new_net_148;
	wire new_net_2623;
	wire new_net_2256;
	wire new_net_3799;
	wire new_net_4884;
	wire new_net_6646;
	wire new_net_9755;
	wire new_net_11190;
	wire new_net_11282;
	wire _1350_;
	wire _1686_;
	wire new_net_2734;
	wire _0468_;
	wire _0048_;
	wire _0342_;
	wire new_net_2627;
	wire new_net_18842;
	wire new_net_7608;
	wire new_net_9126;
	wire new_net_1989;
	wire new_net_4906;
	wire new_net_5204;
	wire new_net_6483;
	wire new_net_7801;
	wire new_net_19981;
	wire new_net_20230;
	wire new_net_1112;
	wire new_net_15291;
	wire new_net_7820;
	wire new_net_16261;
	wire new_net_15298;
	wire new_net_15780;
	wire new_net_16239;
	wire new_net_156;
	wire new_net_12151;
	wire new_net_12942;
	wire new_net_14014;
	wire new_net_14979;
	wire new_net_15116;
	wire new_net_15342;
	wire new_net_17177;
	wire new_net_1982;
	wire new_net_113;
	wire new_net_3304;
	wire new_net_7795;
	wire new_net_14606;
	wire new_net_20221;
	wire new_net_17673;
	wire new_net_13945;
	wire new_net_17562;
	wire new_net_3819;
	wire new_net_17176;
	wire _1352_;
	wire _1688_;
	wire new_net_108;
	wire new_net_1984;
	wire _0470_;
	wire _0050_;
	wire _0344_;
	wire new_net_7796;
	wire new_net_9456;
	wire new_net_4707;
	wire new_net_19250;
	wire new_net_19385;
	wire new_net_21134;
	wire new_net_8608;
	wire _1353_;
	wire _1689_;
	wire new_net_1121;
	wire _0471_;
	wire _0345_;
	wire new_net_2835;
	wire _0051_;
	wire new_net_14604;
	wire new_net_16407;
	wire new_net_7616;
	wire new_net_11191;
	wire new_net_11283;
	wire new_net_2974;
	wire new_net_3414;
	wire new_net_6220;
	wire new_net_13386;
	wire new_net_15296;
	wire new_net_4621;
	wire _0472_;
	wire _1354_;
	wire _1690_;
	wire new_net_1113;
	wire _0052_;
	wire _0346_;
	wire new_net_7800;
	wire new_net_18635;
	wire new_net_19091;
	wire new_net_12915;
	wire new_net_11643;
	wire new_net_15781;
	wire new_net_9759;
	wire new_net_15297;
	wire new_net_17080;
	wire new_net_12943;
	wire new_net_14015;
	wire new_net_14980;
	wire new_net_15117;
	wire new_net_15343;
	wire new_net_15484;
	wire new_net_19046;
	wire new_net_15588;
	wire new_net_18202;
	wire new_net_162;
	wire new_net_3820;
	wire _1355_;
	wire _1691_;
	wire new_net_118;
	wire new_net_2735;
	wire _0473_;
	wire _0347_;
	wire _0053_;
	wire new_net_3296;
	wire new_net_7609;
	wire new_net_9331;
	wire new_net_2985;
	wire new_net_4624;
	wire new_net_4908;
	wire new_net_5199;
	wire new_net_5892;
	wire new_net_19437;
	wire new_net_21300;
	wire new_net_21336;
	wire new_net_15626;
	wire new_net_9754;
	wire new_net_5100;
	wire new_net_10117;
	wire _1356_;
	wire _1692_;
	wire new_net_1120;
	wire _0474_;
	wire _0348_;
	wire new_net_5111;
	wire _0054_;
	wire new_net_9756;
	wire new_net_9129;
	wire new_net_153;
	wire new_net_1114;
	wire new_net_3805;
	wire new_net_5196;
	wire new_net_6648;
	wire new_net_5102;
	wire new_net_11284;
	wire new_net_2739;
	wire new_net_771;
	wire _1357_;
	wire _0475_;
	wire _1693_;
	wire new_net_11192;
	wire _0349_;
	wire _0055_;
	wire new_net_1167;
	wire new_net_17857;
	wire new_net_18932;
	wire new_net_2780;
	wire new_net_12241;
	wire new_net_17918;
	wire new_net_19016;
	wire new_net_18576;
	wire new_net_18700;
	wire new_net_15159;
	wire new_net_12137;
	wire new_net_7178;
	wire new_net_795;
	wire new_net_2460;
	wire new_net_9067;
	wire new_net_20500;
	wire new_net_20654;
	wire new_net_17324;
	wire new_net_6478;
	wire new_net_14023;
	wire new_net_12068;
	wire new_net_13485;
	wire new_net_14414;
	wire new_net_9767;
	wire new_net_15758;
	wire new_net_17839;
	wire new_net_15201;
	wire new_net_14897;
	wire new_net_14956;
	wire new_net_15841;
	wire new_net_10102;
	wire new_net_4687;
	wire new_net_6162;
	wire new_net_15458;
	wire new_net_14292;
	wire new_net_10412;
	wire new_net_4745;
	wire new_net_5248;
	wire new_net_7569;
	wire new_net_11483;
	wire new_net_2464;
	wire _0939_;
	wire new_net_2071;
	wire new_net_19387;
	wire new_net_13053;
	wire new_net_16379;
	wire new_net_9066;
	wire new_net_9772;
	wire new_net_6904;
	wire new_net_800;
	wire new_net_4682;
	wire new_net_4741;
	wire new_net_8396;
	wire new_net_7643;
	wire new_net_17827;
	wire new_net_8268;
	wire new_net_6905;
	wire new_net_5241;
	wire new_net_7833;
	wire new_net_7332;
	wire new_net_803;
	wire _0940_;
	wire new_net_11771;
	wire new_net_780;
	wire new_net_2528;
	wire new_net_8524;
	wire new_net_14401;
	wire new_net_16596;
	wire new_net_17828;
	wire new_net_11553;
	wire new_net_11252;
	wire new_net_11412;
	wire new_net_15508;
	wire new_net_6665;
	wire new_net_7639;
	wire new_net_13119;
	wire new_net_12730;
	wire new_net_5239;
	wire new_net_9770;
	wire new_net_7175;
	wire new_net_8102;
	wire _0941_;
	wire new_net_3837;
	wire new_net_14569;
	wire new_net_20501;
	wire new_net_14902;
	wire new_net_18117;
	wire new_net_12069;
	wire new_net_13486;
	wire new_net_14415;
	wire new_net_9769;
	wire new_net_15759;
	wire new_net_17840;
	wire new_net_15202;
	wire new_net_14898;
	wire new_net_15842;
	wire new_net_2169;
	wire new_net_15821;
	wire new_net_15860;
	wire new_net_18189;
	wire new_net_15507;
	wire _0942_;
	wire new_net_373;
	wire new_net_6168;
	wire new_net_20171;
	wire new_net_14148;
	wire new_net_12533;
	wire new_net_10586;
	wire new_net_1594;
	wire new_net_1901;
	wire new_net_5211;
	wire new_net_7605;
	wire new_net_19388;
	wire new_net_5894;
	wire _0343_;
	wire new_net_13144;
	wire new_net_19443;
	wire new_net_7326;
	wire _0943_;
	wire new_net_337;
	wire new_net_379;
	wire new_net_2468;
	wire new_net_7247;
	wire new_net_18972;
	wire new_net_20653;
	wire new_net_13222;
	wire new_net_7568;
	wire new_net_2172;
	wire new_net_5244;
	wire new_net_6171;
	wire new_net_6674;
	wire new_net_19513;
	wire new_net_16967;
	wire new_net_12740;
	wire new_net_18427;
	wire new_net_20254;
	wire new_net_11554;
	wire new_net_7173;
	wire new_net_11253;
	wire new_net_11413;
	wire new_net_16241;
	wire new_net_15225;
	wire _0944_;
	wire new_net_341;
	wire new_net_6420;
	wire new_net_7912;
	wire new_net_19108;
	wire new_net_15768;
	wire _0973_;
	wire new_net_18347;
	wire new_net_17378;
	wire new_net_18756;
	wire new_net_19073;
	wire new_net_12421;
	wire new_net_6903;
	wire new_net_7577;
	wire new_net_14955;
	wire new_net_3833;
	wire new_net_6663;
	wire new_net_20170;
	wire new_net_20502;
	wire new_net_13706;
	wire new_net_18710;
	wire new_net_13116;
	wire new_net_12070;
	wire new_net_13487;
	wire new_net_14416;
	wire new_net_9764;
	wire new_net_15760;
	wire new_net_15203;
	wire new_net_14899;
	wire new_net_15843;
	wire new_net_2164;
	wire new_net_9728;
	wire new_net_17222;
	wire new_net_17829;
	wire new_net_15506;
	wire new_net_2459;
	wire new_net_2076;
	wire new_net_19571;
	wire new_net_20645;
	wire new_net_7358;
	wire new_net_16833;
	wire new_net_19402;
	wire new_net_14265;
	wire new_net_17591;
	wire new_net_9070;
	wire new_net_6865;
	wire new_net_8096;
	wire new_net_2458;
	wire _0946_;
	wire new_net_5208;
	wire new_net_19389;
	wire new_net_16057;
	wire new_net_16034;
	wire new_net_8707;
	wire new_net_4837;
	wire new_net_6900;
	wire new_net_7918;
	wire new_net_16679;
	wire new_net_4364;
	wire new_net_6206;
	wire new_net_8098;
	wire new_net_1588;
	wire _0947_;
	wire new_net_16508;
	wire new_net_4684;
	wire new_net_18971;
	wire new_net_19512;
	wire new_net_11228;
	wire new_net_14571;
	wire new_net_11555;
	wire new_net_17841;
	wire new_net_11254;
	wire new_net_11414;
	wire new_net_1600;
	wire new_net_1899;
	wire new_net_382;
	wire new_net_6165;
	wire new_net_8097;
	wire new_net_15292;
	wire new_net_19438;
	wire new_net_16262;
	wire new_net_13447;
	wire new_net_6203;
	wire new_net_6866;
	wire new_net_14954;
	wire new_net_12861;
	wire new_net_347;
	wire _0948_;
	wire new_net_6172;
	wire new_net_6412;
	wire new_net_20503;
	wire new_net_7675;
	wire new_net_12726;
	wire new_net_13194;
	wire new_net_14405;
	wire new_net_7642;
	wire new_net_12071;
	wire new_net_13488;
	wire new_net_15761;
	wire new_net_17832;
	wire new_net_15204;
	wire new_net_14900;
	wire new_net_17674;
	wire new_net_15844;
	wire new_net_17563;
	wire new_net_7251;
	wire new_net_17830;
	wire new_net_8100;
	wire _0949_;
	wire new_net_2457;
	wire new_net_15505;
	wire new_net_19252;
	wire new_net_1898;
	wire new_net_4368;
	wire new_net_4836;
	wire new_net_5246;
	wire new_net_19390;
	wire new_net_20644;
	wire _0245_;
	wire new_net_21135;
	wire new_net_4375;
	wire new_net_9773;
	wire _0950_;
	wire new_net_2474;
	wire new_net_1587;
	wire new_net_20651;
	wire new_net_12698;
	wire new_net_7248;
	wire new_net_8101;
	wire new_net_4744;
	wire new_net_6666;
	wire new_net_13555;
	wire new_net_13385;
	wire new_net_19092;
	wire new_net_14572;
	wire new_net_11556;
	wire new_net_342;
	wire _0951_;
	wire new_net_1596;
	wire new_net_2171;
	wire new_net_12879;
	wire new_net_11255;
	wire new_net_11415;
	wire new_net_18970;
	wire new_net_12916;
	wire new_net_7704;
	wire new_net_7917;
	wire new_net_6205;
	wire new_net_2070;
	wire new_net_381;
	wire new_net_797;
	wire new_net_5207;
	wire new_net_14953;
	wire new_net_19047;
	wire new_net_20504;
	wire new_net_18124;
	wire new_net_20986;
	wire new_net_15589;
	wire new_net_18203;
	wire new_net_14418;
	wire new_net_13195;
	wire new_net_13489;
	wire new_net_12725;
	wire new_net_6204;
	wire new_net_12072;
	wire new_net_17833;
	wire new_net_15762;
	wire new_net_17842;
	wire new_net_14406;
	wire new_net_13981;
	wire new_net_346;
	wire new_net_372;
	wire new_net_4681;
	wire new_net_10108;
	wire new_net_15504;
	wire new_net_7640;
	wire new_net_2518;
	wire new_net_19745;
	wire new_net_20388;
	wire new_net_7874;
	wire new_net_16806;
	wire new_net_7911;
	wire new_net_13446;
	wire new_net_10103;
	wire new_net_1902;
	wire new_net_380;
	wire _0953_;
	wire new_net_19391;
	wire new_net_21289;
	wire new_net_11853;
	wire new_net_12467;
	wire new_net_7908;
	wire new_net_2168;
	wire new_net_2477;
	wire new_net_3831;
	wire new_net_10587;
	wire new_net_18961;
	wire new_net_11715;
	wire new_net_6207;
	wire new_net_6867;
	wire new_net_8093;
	wire _0954_;
	wire new_net_17858;
	wire new_net_18933;
	wire new_net_14573;
	wire new_net_7641;
	wire new_net_17831;
	wire new_net_11557;
	wire new_net_2074;
	wire new_net_2167;
	wire new_net_5571;
	wire new_net_6167;
	wire new_net_7330;
	wire new_net_12242;
	wire new_net_17919;
	wire new_net_19017;
	wire new_net_18577;
	wire new_net_18701;
	wire new_net_3835;
	wire new_net_4367;
	wire new_net_2465;
	wire _0955_;
	wire new_net_15160;
	wire new_net_5212;
	wire new_net_14952;
	wire new_net_18969;
	wire new_net_12138;
	wire new_net_20169;
	wire new_net_17325;
	wire new_net_12581;
	wire new_net_13113;
	wire new_net_7253;
	wire new_net_12724;
	wire new_net_13196;
	wire new_net_14407;
	wire new_net_12073;
	wire new_net_13490;
	wire new_net_14419;
	wire new_net_15763;
	wire new_net_14024;
	wire new_net_10106;
	wire new_net_6901;
	wire new_net_7832;
	wire new_net_2467;
	wire _0956_;
	wire new_net_5210;
	wire new_net_8257;
	wire new_net_7327;
	wire new_net_15503;
	wire new_net_15459;
	wire new_net_14293;
	wire new_net_7250;
	wire new_net_13445;
	wire new_net_6908;
	wire new_net_7573;
	wire new_net_376;
	wire new_net_4086;
	wire new_net_19392;
	wire new_net_19509;
	wire new_net_13054;
	wire new_net_16380;
	wire new_net_6675;
	wire new_net_7700;
	wire new_net_9065;
	wire new_net_9771;
	wire _0957_;
	wire new_net_5245;
	wire new_net_20643;
	wire new_net_8731;
	wire new_net_12802;
	wire new_net_19622;
	wire new_net_8402;
	wire new_net_336;
	wire new_net_6201;
	wire new_net_7331;
	wire new_net_13346;
	wire new_net_11772;
	wire new_net_20808;
	wire new_net_14574;
	wire new_net_2165;
	wire _0958_;
	wire new_net_2456;
	wire new_net_4685;
	wire new_net_11558;
	wire new_net_11417;
	wire new_net_20162;
	wire new_net_20852;
	wire new_net_14951;
	wire new_net_10584;
	wire new_net_2469;
	wire new_net_801;
	wire new_net_20506;
	wire new_net_19197;
	wire new_net_14245;
	wire new_net_12582;
	wire new_net_13112;
	wire new_net_15207;
	wire new_net_12723;
	wire new_net_9768;
	wire new_net_17844;
	wire new_net_14420;
	wire new_net_13197;
	wire new_net_13491;
	wire new_net_14903;
	wire new_net_18118;
	wire new_net_20650;
	wire new_net_17166;
	wire new_net_6570;
	wire new_net_10104;
	wire new_net_2077;
	wire new_net_6421;
	wire new_net_15502;
	wire new_net_20168;
	wire new_net_15861;
	wire new_net_18190;
	wire new_net_14149;
	wire new_net_7909;
	wire new_net_13444;
	wire new_net_802;
	wire _0960_;
	wire new_net_2078;
	wire new_net_19393;
	wire new_net_14114;
	wire new_net_9774;
	wire new_net_4372;
	wire new_net_6164;
	wire new_net_11257;
	wire new_net_12643;
	wire new_net_13422;
	wire new_net_13223;
	wire _0961_;
	wire new_net_4683;
	wire new_net_12036;
	wire new_net_12741;
	wire new_net_7535;
	wire new_net_18428;
	wire new_net_14575;
	wire new_net_7646;
	wire new_net_11559;
	wire new_net_1593;
	wire new_net_1904;
	wire new_net_799;
	wire new_net_4749;
	wire new_net_11418;
	wire new_net_20853;
	wire new_net_15226;
	wire new_net_16242;
	wire new_net_13797;
	wire new_net_19109;
	wire new_net_15769;
	wire new_net_18348;
	wire new_net_17379;
	wire new_net_13787;
	wire new_net_18757;
	wire new_net_6673;
	wire new_net_1591;
	wire _0962_;
	wire new_net_5209;
	wire new_net_14950;
	wire new_net_6163;
	wire new_net_19074;
	wire new_net_20166;
	wire new_net_20507;
	wire new_net_13707;
	wire new_net_6417;
	wire new_net_12583;
	wire new_net_13111;
	wire new_net_12722;
	wire new_net_13198;
	wire new_net_14409;
	wire new_net_6200;
	wire new_net_12075;
	wire new_net_13492;
	wire new_net_14421;
	wire new_net_18711;
	wire new_net_8394;
	wire new_net_4746;
	wire new_net_1592;
	wire new_net_1903;
	wire _0963_;
	wire new_net_15501;
	wire new_net_18967;
	wire new_net_20167;
	wire new_net_17223;
	wire new_net_17834;
	wire new_net_13443;
	wire new_net_7571;
	wire new_net_2170;
	wire new_net_375;
	wire new_net_7648;
	wire new_net_14266;
	wire new_net_17592;
	wire new_net_19394;
	wire new_net_19403;
	wire new_net_16058;
	wire new_net_19214;
	wire _0964_;
	wire new_net_7333;
	wire new_net_16680;
	wire new_net_13521;
	wire new_net_9765;
	wire new_net_7647;
	wire new_net_9064;
	wire new_net_6202;
	wire new_net_6419;
	wire new_net_10101;
	wire new_net_16509;
	wire new_net_6685;
	wire new_net_14576;
	wire new_net_11560;
	wire new_net_4742;
	wire new_net_343;
	wire new_net_371;
	wire new_net_1896;
	wire new_net_2166;
	wire _0965_;
	wire new_net_11258;
	wire new_net_11419;
	wire new_net_12814;
	wire new_net_14813;
	wire new_net_2030;
	wire new_net_16263;
	wire new_net_4686;
	wire new_net_6170;
	wire new_net_7575;
	wire new_net_14949;
	wire new_net_18962;
	wire new_net_20508;
	wire new_net_12862;
	wire new_net_2210;
	wire new_net_14070;
	wire new_net_14247;
	wire new_net_14422;
	wire new_net_12584;
	wire new_net_13110;
	wire new_net_4365;
	wire new_net_12721;
	wire new_net_13199;
	wire new_net_14410;
	wire new_net_12076;
	wire new_net_17675;
	wire new_net_6362;
	wire new_net_15845;
	wire new_net_1894;
	wire new_net_15500;
	wire new_net_17564;
	wire new_net_8953;
	wire new_net_7916;
	wire new_net_17835;
	wire new_net_7177;
	wire _0967_;
	wire new_net_1897;
	wire new_net_18966;
	wire new_net_19238;
	wire new_net_19395;
	wire new_net_20648;
	wire new_net_21136;
	wire new_net_7252;
	wire new_net_7702;
	wire new_net_6199;
	wire new_net_2072;
	wire new_net_4629;
	wire new_net_7831;
	wire new_net_19508;
	wire new_net_12506;
	wire new_net_12699;
	wire new_net_19435;
	wire new_net_7703;
	wire new_net_7910;
	wire new_net_13442;
	wire new_net_7644;
	wire new_net_7179;
	wire new_net_10591;
	wire new_net_1589;
	wire _0968_;
	wire new_net_13554;
	wire new_net_13384;
	wire new_net_5568;
	wire new_net_8393;
	wire new_net_14577;
	wire new_net_11561;
	wire new_net_374;
	wire new_net_11259;
	wire new_net_11420;
	wire new_net_20647;
	wire new_net_20855;
	wire new_net_19093;
	wire new_net_12917;
	wire new_net_6418;
	wire new_net_7915;
	wire new_net_10590;
	wire new_net_338;
	wire new_net_1598;
	wire new_net_1905;
	wire _0969_;
	wire new_net_14948;
	wire new_net_20509;
	wire new_net_12190;
	wire new_net_19048;
	wire new_net_15590;
	wire new_net_18204;
	wire new_net_14071;
	wire new_net_14248;
	wire new_net_12585;
	wire new_net_13109;
	wire new_net_12720;
	wire new_net_13200;
	wire new_net_14411;
	wire new_net_12077;
	wire new_net_13494;
	wire new_net_14423;
	wire new_net_4628;
	wire new_net_8709;
	wire _0970_;
	wire new_net_794;
	wire new_net_8103;
	wire new_net_10593;
	wire new_net_5247;
	wire new_net_7329;
	wire new_net_15499;
	wire new_net_7732;
	wire new_net_17836;
	wire new_net_2073;
	wire new_net_6664;
	wire new_net_6864;
	wire new_net_19396;
	wire new_net_6609;
	wire new_net_11854;
	wire new_net_12468;
	wire _0971_;
	wire new_net_6906;
	wire new_net_7574;
	wire new_net_7834;
	wire new_net_18965;
	wire new_net_19507;
	wire new_net_20165;
	wire new_net_20646;
	wire new_net_11716;
	wire new_net_7249;
	wire new_net_2472;
	wire new_net_796;
	wire new_net_1893;
	wire new_net_4627;
	wire new_net_4838;
	wire new_net_17859;
	wire new_net_18934;
	wire new_net_11260;
	wire new_net_11421;
	wire new_net_14578;
	wire new_net_11562;
	wire new_net_804;
	wire _0972_;
	wire new_net_4087;
	wire new_net_4630;
	wire new_net_18121;
	wire new_net_19504;
	wire new_net_2792;
	wire new_net_12243;
	wire new_net_17920;
	wire new_net_19018;
	wire new_net_18578;
	wire new_net_18702;
	wire new_net_5205;
	wire new_net_14947;
	wire new_net_4370;
	wire new_net_8400;
	wire new_net_10107;
	wire new_net_1895;
	wire new_net_340;
	wire new_net_6907;
	wire new_net_10588;
	wire new_net_3407;
	wire new_net_15161;
	wire new_net_17326;
	wire new_net_15851;
	wire new_net_14072;
	wire new_net_14249;
	wire new_net_6671;
	wire new_net_12586;
	wire new_net_13108;
	wire new_net_12719;
	wire new_net_13201;
	wire new_net_14412;
	wire new_net_7649;
	wire new_net_14025;
	wire new_net_18147;
	wire new_net_14945;
	wire new_net_15498;
	wire new_net_6414;
	wire new_net_6198;
	wire new_net_9069;
	wire new_net_3836;
	wire new_net_4740;
	wire new_net_6863;
	wire new_net_7176;
	wire new_net_15460;
	wire new_net_19235;
	wire new_net_14294;
	wire new_net_15497;
	wire new_net_4371;
	wire new_net_7913;
	wire new_net_13441;
	wire new_net_4739;
	wire new_net_17837;
	wire new_net_8708;
	wire new_net_2475;
	wire _0974_;
	wire new_net_7172;
	wire new_net_21262;
	wire new_net_9997;
	wire new_net_8706;
	wire new_net_4369;
	wire new_net_20161;
	wire new_net_8733;
	wire new_net_12803;
	wire new_net_5206;
	wire new_net_6413;
	wire new_net_4835;
	wire new_net_7645;
	wire new_net_7823;
	wire _0975_;
	wire new_net_377;
	wire new_net_2476;
	wire new_net_4374;
	wire new_net_7579;
	wire new_net_7328;
	wire new_net_11261;
	wire new_net_11422;
	wire new_net_8401;
	wire new_net_14579;
	wire new_net_9766;
	wire new_net_11563;
	wire new_net_1906;
	wire new_net_4373;
	wire new_net_4626;
	wire new_net_12841;
	wire new_net_14946;
	wire _0976_;
	wire new_net_6416;
	wire new_net_20511;
	wire new_net_19055;
	wire new_net_19198;
	wire new_net_15852;
	wire new_net_6166;
	wire new_net_14073;
	wire new_net_14250;
	wire new_net_12587;
	wire new_net_7255;
	wire new_net_13439;
	wire new_net_14413;
	wire new_net_12079;
	wire new_net_13496;
	wire new_net_14904;
	wire new_net_18119;
	wire new_net_17167;
	wire new_net_13202;
	wire new_net_14580;
	wire new_net_4743;
	wire new_net_10109;
	wire new_net_1595;
	wire _0977_;
	wire new_net_3832;
	wire new_net_8095;
	wire new_net_10583;
	wire new_net_18191;
	wire new_net_14150;
	wire new_net_8397;
	wire new_net_13440;
	wire new_net_10100;
	wire new_net_2463;
	wire new_net_1597;
	wire new_net_4631;
	wire new_net_6197;
	wire new_net_6909;
	wire new_net_10594;
	wire new_net_19239;
	wire new_net_7413;
	wire new_net_7604;
	wire new_net_11875;
	wire new_net_12571;
	wire new_net_8398;
	wire new_net_10213;
	wire _0978_;
	wire new_net_2173;
	wire new_net_335;
	wire new_net_7174;
	wire new_net_5243;
	wire new_net_19240;
	wire new_net_19505;
	wire new_net_12644;
	wire new_net_13423;
	wire new_net_1664;
	wire new_net_6672;
	wire new_net_7254;
	wire new_net_7701;
	wire new_net_8399;
	wire new_net_9068;
	wire new_net_4632;
	wire new_net_6415;
	wire new_net_10589;
	wire new_net_7576;
	wire new_net_14474;
	wire new_net_7861;
	wire new_net_12037;
	wire new_net_11262;
	wire new_net_11423;
	wire new_net_11564;
	wire new_net_2461;
	wire new_net_2079;
	wire _0979_;
	wire new_net_5242;
	wire new_net_18777;
	wire new_net_12742;
	wire new_net_18429;
	wire new_net_15227;
	wire new_net_16243;
	wire new_net_19110;
	wire new_net_17380;
	wire new_net_13788;
	wire new_net_18758;
	wire new_net_19075;
	wire new_net_13996;
	wire new_net_2753;
	wire new_net_13708;
	wire new_net_19000;
	wire new_net_15107;
	wire new_net_18712;
	wire new_net_1809;
	wire new_net_18316;
	wire new_net_18467;
	wire new_net_19911;
	wire new_net_20607;
	wire new_net_14323;
	wire new_net_15403;
	wire new_net_17212;
	wire new_net_14379;
	wire new_net_13345;
	wire new_net_16798;
	wire new_net_11868;
	wire new_net_17188;
	wire new_net_12907;
	wire new_net_4088;
	wire new_net_12695;
	wire new_net_8353;
	wire new_net_1810;
	wire new_net_6303;
	wire new_net_7600;
	wire new_net_18313;
	wire new_net_13118;
	wire new_net_16059;
	wire new_net_3795;
	wire new_net_7662;
	wire new_net_5298;
	wire new_net_6745;
	wire new_net_16318;
	wire _0477_;
	wire new_net_2089;
	wire new_net_19423;
	wire new_net_20649;
	wire new_net_16681;
	wire new_net_20900;
	wire new_net_9313;
	wire new_net_8634;
	wire new_net_1066;
	wire new_net_2324;
	wire new_net_6065;
	wire new_net_7663;
	wire new_net_11230;
	wire new_net_4354;
	wire new_net_6304;
	wire new_net_9312;
	wire new_net_12527;
	wire new_net_8408;
	wire _0478_;
	wire new_net_20782;
	wire new_net_15294;
	wire new_net_5896;
	wire new_net_12815;
	wire new_net_14814;
	wire new_net_16264;
	wire new_net_11309;
	wire new_net_9315;
	wire new_net_11448;
	wire new_net_7595;
	wire new_net_10910;
	wire new_net_8297;
	wire new_net_11052;
	wire new_net_1803;
	wire new_net_4545;
	wire new_net_5452;
	wire new_net_12863;
	wire new_net_4350;
	wire new_net_9318;
	wire new_net_10617;
	wire new_net_6589;
	wire new_net_6752;
	wire _0479_;
	wire new_net_6059;
	wire new_net_19912;
	wire new_net_20608;
	wire new_net_17676;
	wire new_net_15846;
	wire new_net_17565;
	wire new_net_15404;
	wire new_net_17189;
	wire new_net_9317;
	wire new_net_17213;
	wire new_net_16799;
	wire new_net_17496;
	wire new_net_11869;
	wire new_net_12566;
	wire new_net_6424;
	wire new_net_12696;
	wire new_net_9711;
	wire new_net_8626;
	wire new_net_5453;
	wire new_net_1800;
	wire new_net_6754;
	wire _0480_;
	wire new_net_443;
	wire _0252_;
	wire new_net_21137;
	wire new_net_20223;
	wire new_net_6631;
	wire new_net_8296;
	wire new_net_3543;
	wire new_net_4089;
	wire new_net_19424;
	wire new_net_12044;
	wire new_net_12700;
	wire new_net_20383;
	wire new_net_6300;
	wire new_net_14050;
	wire new_net_9320;
	wire new_net_7594;
	wire _0481_;
	wire new_net_18324;
	wire new_net_18476;
	wire new_net_20386;
	wire new_net_3987;
	wire new_net_13553;
	wire new_net_13383;
	wire new_net_12528;
	wire new_net_4543;
	wire new_net_6503;
	wire new_net_9603;
	wire new_net_19094;
	wire new_net_20783;
	wire new_net_14809;
	wire new_net_3597;
	wire new_net_19236;
	wire new_net_12918;
	wire new_net_11310;
	wire new_net_11449;
	wire new_net_10911;
	wire new_net_11053;
	wire _0482_;
	wire new_net_4553;
	wire new_net_12191;
	wire new_net_19049;
	wire new_net_15591;
	wire new_net_18205;
	wire new_net_9310;
	wire new_net_10614;
	wire new_net_57;
	wire new_net_2320;
	wire new_net_2726;
	wire new_net_19913;
	wire new_net_20609;
	wire new_net_13983;
	wire new_net_9626;
	wire new_net_15405;
	wire new_net_17190;
	wire new_net_17214;
	wire new_net_7599;
	wire new_net_16800;
	wire new_net_17497;
	wire new_net_11870;
	wire new_net_12567;
	wire new_net_12697;
	wire new_net_13347;
	wire new_net_6504;
	wire new_net_7602;
	wire new_net_6591;
	wire new_net_7591;
	wire new_net_55;
	wire new_net_4353;
	wire new_net_20384;
	wire new_net_14714;
	wire new_net_11855;
	wire new_net_12469;
	wire new_net_10001;
	wire new_net_6507;
	wire new_net_8630;
	wire new_net_5451;
	wire new_net_4091;
	wire new_net_5415;
	wire new_net_1799;
	wire _0484_;
	wire new_net_18323;
	wire new_net_18475;
	wire new_net_11717;
	wire new_net_8356;
	wire new_net_10618;
	wire new_net_20387;
	wire new_net_17860;
	wire new_net_18935;
	wire new_net_5454;
	wire new_net_9426;
	wire new_net_2723;
	wire _0485_;
	wire new_net_2318;
	wire new_net_20784;
	wire new_net_17921;
	wire new_net_19019;
	wire new_net_18579;
	wire new_net_11311;
	wire new_net_11450;
	wire new_net_10912;
	wire new_net_11054;
	wire new_net_6586;
	wire new_net_8969;
	wire new_net_15162;
	wire new_net_17327;
	wire _0486_;
	wire new_net_19914;
	wire new_net_20385;
	wire new_net_20610;
	wire new_net_17601;
	wire new_net_14026;
	wire new_net_18148;
	wire new_net_12904;
	wire new_net_15145;
	wire new_net_15406;
	wire new_net_17191;
	wire new_net_17215;
	wire new_net_6594;
	wire new_net_12526;
	wire new_net_16801;
	wire new_net_17498;
	wire new_net_11871;
	wire new_net_14295;
	wire new_net_6064;
	wire new_net_8530;
	wire new_net_14049;
	wire new_net_6500;
	wire _0487_;
	wire new_net_63;
	wire new_net_1068;
	wire new_net_21263;
	wire new_net_19397;
	wire new_net_14060;
	wire new_net_9994;
	wire new_net_16382;
	wire new_net_6426;
	wire new_net_439;
	wire new_net_4246;
	wire new_net_4544;
	wire new_net_6068;
	wire new_net_19426;
	wire new_net_12804;
	wire new_net_20222;
	wire new_net_6060;
	wire new_net_9319;
	wire new_net_6595;
	wire _0488_;
	wire new_net_1806;
	wire new_net_58;
	wire new_net_13348;
	wire new_net_20810;
	wire new_net_4247;
	wire new_net_5410;
	wire new_net_2081;
	wire new_net_20785;
	wire new_net_13803;
	wire new_net_18596;
	wire new_net_12842;
	wire new_net_19056;
	wire new_net_11312;
	wire new_net_11451;
	wire new_net_10913;
	wire new_net_12568;
	wire new_net_6632;
	wire new_net_11055;
	wire _0489_;
	wire new_net_61;
	wire new_net_2322;
	wire new_net_8971;
	wire new_net_9211;
	wire new_net_10000;
	wire new_net_7596;
	wire new_net_1808;
	wire new_net_2730;
	wire new_net_3308;
	wire new_net_4542;
	wire new_net_6749;
	wire new_net_19915;
	wire new_net_14905;
	wire new_net_18120;
	wire new_net_17168;
	wire new_net_12903;
	wire new_net_15146;
	wire new_net_15407;
	wire new_net_17192;
	wire new_net_17216;
	wire new_net_16802;
	wire new_net_17499;
	wire new_net_11872;
	wire new_net_5299;
	wire new_net_6635;
	wire new_net_15415;
	wire new_net_15863;
	wire new_net_18192;
	wire new_net_14151;
	wire new_net_20317;
	wire new_net_9601;
	wire new_net_14048;
	wire new_net_5411;
	wire new_net_18314;
	wire new_net_18468;
	wire new_net_9224;
	wire new_net_7956;
	wire new_net_12536;
	wire new_net_14116;
	wire new_net_11876;
	wire new_net_12572;
	wire new_net_20382;
	wire new_net_6067;
	wire new_net_2321;
	wire _0491_;
	wire new_net_19427;
	wire new_net_12645;
	wire new_net_13424;
	wire new_net_11691;
	wire new_net_7484;
	wire new_net_13225;
	wire new_net_6585;
	wire new_net_1804;
	wire new_net_18322;
	wire new_net_18474;
	wire new_net_14475;
	wire new_net_8105;
	wire new_net_12038;
	wire new_net_16970;
	wire new_net_18778;
	wire new_net_12525;
	wire new_net_9425;
	wire new_net_6633;
	wire _0492_;
	wire new_net_20786;
	wire new_net_15228;
	wire new_net_16244;
	wire new_net_13799;
	wire new_net_19111;
	wire new_net_17381;
	wire new_net_11313;
	wire new_net_11452;
	wire new_net_10914;
	wire new_net_11056;
	wire new_net_13789;
	wire new_net_18759;
	wire new_net_19076;
	wire new_net_13997;
	wire new_net_13709;
	wire new_net_3544;
	wire new_net_9311;
	wire new_net_6593;
	wire new_net_8298;
	wire _0493_;
	wire new_net_3321;
	wire new_net_19916;
	wire new_net_20612;
	wire new_net_18713;
	wire new_net_12902;
	wire new_net_15147;
	wire new_net_15408;
	wire new_net_17193;
	wire new_net_10622;
	wire new_net_17217;
	wire new_net_16803;
	wire new_net_17500;
	wire new_net_11873;
	wire new_net_12569;
	wire new_net_4351;
	wire new_net_14047;
	wire new_net_1063;
	wire _0494_;
	wire new_net_17594;
	wire new_net_14268;
	wire new_net_13117;
	wire new_net_16060;
	wire new_net_8527;
	wire new_net_9316;
	wire new_net_7597;
	wire new_net_1060;
	wire new_net_445;
	wire new_net_4546;
	wire new_net_19428;
	wire new_net_3680;
	wire new_net_4886;
	wire new_net_16037;
	wire new_net_16319;
	wire new_net_16682;
	wire new_net_6302;
	wire new_net_8357;
	wire new_net_8628;
	wire new_net_12523;
	wire new_net_1064;
	wire _0495_;
	wire new_net_16511;
	wire new_net_13179;
	wire new_net_4548;
	wire new_net_4355;
	wire new_net_6310;
	wire new_net_8358;
	wire new_net_9314;
	wire new_net_10616;
	wire new_net_5450;
	wire new_net_5409;
	wire new_net_1070;
	wire new_net_6753;
	wire new_net_15295;
	wire new_net_21316;
	wire new_net_12816;
	wire new_net_14815;
	wire new_net_9602;
	wire new_net_11314;
	wire new_net_11453;
	wire new_net_7601;
	wire new_net_10915;
	wire new_net_11057;
	wire new_net_64;
	wire new_net_1056;
	wire _0496_;
	wire new_net_446;
	wire new_net_12864;
	wire new_net_8970;
	wire new_net_6637;
	wire new_net_19917;
	wire new_net_20613;
	wire new_net_17677;
	wire new_net_4024;
	wire new_net_12901;
	wire new_net_15148;
	wire new_net_15409;
	wire new_net_17194;
	wire new_net_3547;
	wire new_net_17218;
	wire new_net_16804;
	wire new_net_17501;
	wire new_net_11874;
	wire new_net_12570;
	wire new_net_15847;
	wire new_net_17566;
	wire new_net_8957;
	wire new_net_14046;
	wire new_net_12524;
	wire new_net_9427;
	wire new_net_3409;
	wire new_net_3542;
	wire new_net_8410;
	wire new_net_12621;
	wire new_net_21138;
	wire new_net_6069;
	wire _0498_;
	wire new_net_2717;
	wire new_net_8295;
	wire _1568_;
	wire new_net_19429;
	wire new_net_12045;
	wire new_net_12701;
	wire new_net_778;
	wire new_net_9599;
	wire new_net_6505;
	wire new_net_7876;
	wire new_net_1807;
	wire new_net_5458;
	wire new_net_13552;
	wire new_net_13382;
	wire new_net_6066;
	wire new_net_7660;
	wire new_net_2728;
	wire _0499_;
	wire new_net_56;
	wire new_net_2323;
	wire new_net_5412;
	wire new_net_447;
	wire new_net_8407;
	wire new_net_20788;
	wire new_net_19095;
	wire new_net_12882;
	wire new_net_14810;
	wire new_net_3572;
	wire new_net_18560;
	wire new_net_12919;
	wire new_net_8968;
	wire new_net_11315;
	wire new_net_11454;
	wire new_net_6508;
	wire new_net_8629;
	wire new_net_12517;
	wire new_net_10916;
	wire new_net_2090;
	wire new_net_2718;
	wire new_net_3541;
	wire new_net_12192;
	wire new_net_19050;
	wire new_net_4356;
	wire new_net_6307;
	wire new_net_10615;
	wire new_net_1069;
	wire _0500_;
	wire new_net_3545;
	wire new_net_8294;
	wire new_net_6748;
	wire new_net_18465;
	wire new_net_19918;
	wire new_net_13984;
	wire new_net_6283;
	wire new_net_5229;
	wire new_net_14564;
	wire new_net_4539;
	wire new_net_12900;
	wire new_net_15410;
	wire new_net_17195;
	wire new_net_17219;
	wire new_net_15149;
	wire new_net_17502;
	wire new_net_8635;
	wire new_net_16805;
	wire new_net_14045;
	wire new_net_10620;
	wire _0501_;
	wire new_net_54;
	wire new_net_16809;
	wire new_net_10621;
	wire new_net_12522;
	wire new_net_2729;
	wire new_net_442;
	wire new_net_1058;
	wire new_net_5413;
	wire new_net_19430;
	wire new_net_11718;
	wire new_net_19199;
	wire new_net_3303;
	wire new_net_8403;
	wire new_net_6063;
	wire new_net_6506;
	wire new_net_2721;
	wire _0502_;
	wire new_net_66;
	wire new_net_1065;
	wire new_net_6634;
	wire new_net_3796;
	wire new_net_1161;
	wire new_net_17861;
	wire new_net_18936;
	wire new_net_2722;
	wire new_net_8631;
	wire new_net_18320;
	wire new_net_18472;
	wire new_net_20789;
	wire new_net_9776;
	wire new_net_18580;
	wire new_net_7664;
	wire new_net_11316;
	wire new_net_8350;
	wire new_net_11455;
	wire new_net_8632;
	wire new_net_10917;
	wire _0503_;
	wire new_net_62;
	wire new_net_11059;
	wire new_net_15163;
	wire new_net_19742;
	wire new_net_15865;
	wire new_net_15077;
	wire new_net_17328;
	wire new_net_1062;
	wire new_net_2325;
	wire new_net_19919;
	wire new_net_20390;
	wire new_net_20615;
	wire new_net_15522;
	wire new_net_17602;
	wire new_net_8432;
	wire new_net_14027;
	wire new_net_11049;
	wire new_net_18149;
	wire new_net_13353;
	wire new_net_14387;
	wire new_net_14565;
	wire new_net_9598;
	wire new_net_12899;
	wire new_net_15150;
	wire new_net_8529;
	wire new_net_15411;
	wire new_net_17196;
	wire new_net_17220;
	wire new_net_6061;
	wire new_net_14044;
	wire new_net_6590;
	wire new_net_14296;
	wire new_net_2087;
	wire new_net_441;
	wire new_net_6366;
	wire new_net_20389;
	wire new_net_14204;
	wire new_net_19398;
	wire new_net_14059;
	wire new_net_4541;
	wire new_net_12521;
	wire _0505_;
	wire new_net_19431;
	wire new_net_16383;
	wire new_net_6751;
	wire new_net_2086;
	wire new_net_2326;
	wire new_net_12805;
	wire new_net_13349;
	wire new_net_6649;
	wire new_net_65;
	wire new_net_1059;
	wire new_net_8355;
	wire new_net_1801;
	wire _0506_;
	wire new_net_17815;
	wire new_net_20790;
	wire new_net_13804;
	wire new_net_18597;
	wire new_net_12843;
	wire new_net_11060;
	wire new_net_11317;
	wire new_net_10918;
	wire new_net_8409;
	wire new_net_9600;
	wire new_net_11456;
	wire new_net_19057;
	wire new_net_8404;
	wire new_net_6306;
	wire _0507_;
	wire new_net_3325;
	wire new_net_18466;
	wire new_net_19920;
	wire new_net_20391;
	wire new_net_20616;
	wire new_net_14906;
	wire new_net_15389;
	wire new_net_17169;
	wire new_net_15151;
	wire new_net_17504;
	wire new_net_13354;
	wire new_net_14566;
	wire new_net_16807;
	wire new_net_15412;
	wire new_net_12898;
	wire new_net_17221;
	wire new_net_14388;
	wire new_net_17197;
	wire new_net_15416;
	wire new_net_6492;
	wire new_net_15864;
	wire new_net_18193;
	wire new_net_14152;
	wire new_net_14043;
	wire new_net_2085;
	wire new_net_4349;
	wire new_net_9999;
	wire new_net_6498;
	wire _0508_;
	wire new_net_2725;
	wire new_net_5414;
	wire new_net_12537;
	wire new_net_14117;
	wire new_net_9597;
	wire new_net_12520;
	wire new_net_2317;
	wire new_net_5449;
	wire new_net_11877;
	wire new_net_12573;
	wire new_net_8292;
	wire new_net_18318;
	wire new_net_18470;
	wire new_net_19432;
	wire new_net_12646;
	wire new_net_13425;
	wire new_net_11692;
	wire new_net_4538;
	wire new_net_6062;
	wire new_net_8352;
	wire new_net_6499;
	wire _0509_;
	wire new_net_7533;
	wire new_net_13226;
	wire new_net_12039;
	wire new_net_8354;
	wire new_net_448;
	wire new_net_5416;
	wire new_net_6309;
	wire new_net_6502;
	wire new_net_7875;
	wire new_net_7650;
	wire new_net_18779;
	wire new_net_15229;
	wire new_net_16245;
	wire new_net_13800;
	wire new_net_19112;
	wire new_net_11061;
	wire new_net_11318;
	wire new_net_11457;
	wire new_net_2327;
	wire new_net_816;
	wire _0510_;
	wire new_net_10919;
	wire new_net_17382;
	wire new_net_13790;
	wire new_net_18760;
	wire new_net_19077;
	wire new_net_13998;
	wire new_net_13710;
	wire new_net_6308;
	wire new_net_7661;
	wire new_net_2727;
	wire new_net_5457;
	wire new_net_19921;
	wire new_net_20617;
	wire new_net_15109;
	wire new_net_7952;
	wire new_net_8540;
	wire new_net_827;
	wire new_net_11058;
	wire new_net_5300;
	wire new_net_12705;
	wire new_net_6747;
	wire new_net_13355;
	wire new_net_14389;
	wire new_net_15152;
	wire new_net_17505;
	wire new_net_14567;
	wire new_net_12897;
	wire new_net_16808;
	wire new_net_14325;
	wire new_net_17946;
	wire new_net_14042;
	wire new_net_2088;
	wire new_net_18315;
	wire new_net_20392;
	wire new_net_14269;
	wire new_net_17595;
	wire new_net_16061;
	wire new_net_6425;
	wire new_net_8291;
	wire new_net_2731;
	wire new_net_7598;
	wire _0512_;
	wire new_net_1805;
	wire new_net_12519;
	wire new_net_19433;
	wire new_net_16038;
	wire new_net_16320;
	wire new_net_3874;
	wire new_net_6501;
	wire new_net_440;
	wire new_net_4090;
	wire new_net_7593;
	wire new_net_13427;
	wire new_net_16512;
	wire new_net_13180;
	wire new_net_8633;
	wire new_net_1061;
	wire new_net_2084;
	wire _0513_;
	wire new_net_6689;
	wire new_net_11062;
	wire new_net_6746;
	wire new_net_8406;
	wire new_net_10791;
	wire new_net_11319;
	wire new_net_11458;
	wire new_net_7877;
	wire new_net_60;
	wire new_net_2083;
	wire new_net_4352;
	wire new_net_12817;
	wire new_net_14816;
	wire new_net_12865;
	wire new_net_9998;
	wire _0514_;
	wire new_net_2724;
	wire new_net_9428;
	wire new_net_19922;
	wire new_net_20618;
	wire new_net_20846;
	wire new_net_17678;
	wire new_net_12706;
	wire new_net_6744;
	wire new_net_13356;
	wire new_net_14390;
	wire new_net_15153;
	wire new_net_6305;
	wire new_net_8528;
	wire new_net_15414;
	wire new_net_17199;
	wire new_net_14568;
	wire new_net_15848;
	wire new_net_4547;
	wire new_net_14041;
	wire new_net_6592;
	wire new_net_7592;
	wire new_net_8627;
	wire new_net_53;
	wire _0515_;
	wire new_net_5455;
	wire _0259_;
	wire new_net_21139;
	wire new_net_444;
	wire new_net_1067;
	wire new_net_5417;
	wire new_net_6636;
	wire new_net_19434;
	wire new_net_8446;
	wire new_net_12046;
	wire new_net_4244;
	wire new_net_12702;
	wire new_net_6301;
	wire new_net_10002;
	wire new_net_2328;
	wire _0516_;
	wire new_net_18317;
	wire new_net_18469;
	wire new_net_20393;
	wire new_net_7323;
	wire new_net_3412;
	wire new_net_4245;
	wire new_net_13381;
	wire new_net_17306;
	wire new_net_19096;
	wire new_net_12883;
	wire new_net_14811;
	wire new_net_3573;
	wire new_net_11063;
	wire new_net_10792;
	wire new_net_11320;
	wire new_net_14040;
	wire new_net_11459;
	wire new_net_6588;
	wire new_net_12518;
	wire new_net_2319;
	wire _0517_;
	wire new_net_10921;
	wire new_net_12193;
	wire new_net_19051;
	wire new_net_8852;
	wire new_net_13985;
	wire new_net_19612;
	wire new_net_4615;
	wire new_net_15569;
	wire new_net_4023;
	wire new_net_4446;
	wire new_net_18265;
	wire new_net_19899;
	wire new_net_19923;
	wire new_net_19425;
	wire new_net_16042;
	wire new_net_16336;
	wire new_net_11680;
	wire new_net_13321;
	wire new_net_13531;
	wire new_net_16562;
	wire new_net_17850;
	wire new_net_13792;
	wire new_net_12186;
	wire new_net_14861;
	wire new_net_2001;
	wire new_net_9513;
	wire new_net_19514;
	wire new_net_11719;
	wire new_net_20115;
	wire new_net_7632;
	wire new_net_2590;
	wire _1737_;
	wire new_net_2660;
	wire new_net_9264;
	wire new_net_10674;
	wire new_net_1580;
	wire new_net_724;
	wire new_net_3384;
	wire new_net_3847;
	wire new_net_4447;
	wire new_net_6191;
	wire new_net_18581;
	wire new_net_10669;
	wire new_net_6625;
	wire new_net_9510;
	wire new_net_1169;
	wire new_net_2428;
	wire _1738_;
	wire new_net_6378;
	wire new_net_15164;
	wire new_net_15866;
	wire new_net_17756;
	wire new_net_10311;
	wire new_net_15078;
	wire new_net_17329;
	wire new_net_11028;
	wire new_net_13532;
	wire new_net_11158;
	wire new_net_4011;
	wire new_net_722;
	wire new_net_907;
	wire new_net_1997;
	wire new_net_6388;
	wire new_net_6923;
	wire new_net_617;
	wire new_net_15523;
	wire new_net_17603;
	wire new_net_18150;
	wire new_net_2698;
	wire _1739_;
	wire new_net_719;
	wire new_net_6930;
	wire new_net_11808;
	wire new_net_19900;
	wire new_net_19924;
	wire new_net_20175;
	wire new_net_8256;
	wire new_net_12505;
	wire new_net_16810;
	wire new_net_14297;
	wire new_net_16043;
	wire new_net_6847;
	wire new_net_16337;
	wire new_net_11681;
	wire new_net_17851;
	wire new_net_16563;
	wire new_net_13793;
	wire new_net_13121;
	wire new_net_17449;
	wire new_net_12187;
	wire new_net_7570;
	wire new_net_14205;
	wire new_net_9543;
	wire new_net_5469;
	wire new_net_4445;
	wire new_net_1995;
	wire new_net_2588;
	wire _1740_;
	wire new_net_718;
	wire new_net_20174;
	wire new_net_12806;
	wire new_net_15804;
	wire new_net_10652;
	wire new_net_1166;
	wire new_net_1572;
	wire new_net_2431;
	wire new_net_4361;
	wire new_net_5421;
	wire new_net_11819;
	wire new_net_20176;
	wire new_net_13350;
	wire new_net_6652;
	wire new_net_11355;
	wire new_net_3843;
	wire new_net_2587;
	wire new_net_906;
	wire new_net_2429;
	wire _1741_;
	wire new_net_4441;
	wire new_net_20177;
	wire new_net_5823;
	wire new_net_13805;
	wire new_net_18598;
	wire new_net_12844;
	wire new_net_15568;
	wire new_net_6624;
	wire new_net_7039;
	wire new_net_8041;
	wire new_net_9517;
	wire new_net_19058;
	wire new_net_19200;
	wire new_net_9202;
	wire new_net_8040;
	wire new_net_3382;
	wire new_net_11029;
	wire new_net_5475;
	wire new_net_15570;
	wire new_net_11159;
	wire new_net_905;
	wire new_net_2432;
	wire _1742_;
	wire new_net_6924;
	wire new_net_19590;
	wire new_net_14907;
	wire new_net_15388;
	wire new_net_17170;
	wire new_net_6846;
	wire new_net_1168;
	wire new_net_1574;
	wire new_net_2659;
	wire new_net_19901;
	wire new_net_19925;
	wire new_net_5178;
	wire new_net_15417;
	wire new_net_96;
	wire new_net_5343;
	wire new_net_14153;
	wire new_net_10673;
	wire new_net_16044;
	wire new_net_16338;
	wire new_net_13323;
	wire new_net_16564;
	wire new_net_6441;
	wire new_net_12188;
	wire new_net_14863;
	wire new_net_15547;
	wire new_net_15797;
	wire new_net_5307;
	wire new_net_12538;
	wire new_net_14118;
	wire new_net_11878;
	wire new_net_12574;
	wire new_net_5876;
	wire new_net_15571;
	wire new_net_1999;
	wire new_net_2662;
	wire new_net_3844;
	wire new_net_4845;
	wire new_net_16598;
	wire new_net_12647;
	wire new_net_13426;
	wire new_net_11693;
	wire new_net_6384;
	wire new_net_11811;
	wire new_net_6850;
	wire new_net_5418;
	wire _1744_;
	wire new_net_714;
	wire new_net_1163;
	wire new_net_2420;
	wire new_net_14477;
	wire new_net_12040;
	wire new_net_8039;
	wire new_net_10678;
	wire new_net_2661;
	wire new_net_2423;
	wire new_net_2584;
	wire new_net_7652;
	wire new_net_18780;
	wire new_net_15230;
	wire new_net_16246;
	wire new_net_13801;
	wire new_net_19113;
	wire new_net_15119;
	wire new_net_5878;
	wire new_net_9507;
	wire new_net_4358;
	wire _1745_;
	wire new_net_13791;
	wire new_net_18761;
	wire new_net_19078;
	wire new_net_10748;
	wire new_net_13999;
	wire new_net_6929;
	wire new_net_13794;
	wire new_net_11356;
	wire new_net_11682;
	wire new_net_10677;
	wire new_net_11160;
	wire new_net_11030;
	wire new_net_10818;
	wire new_net_1576;
	wire new_net_1172;
	wire new_net_11070;
	wire new_net_6651;
	wire new_net_10671;
	wire new_net_13530;
	wire new_net_6619;
	wire _1746_;
	wire new_net_2438;
	wire new_net_2670;
	wire new_net_1584;
	wire new_net_19902;
	wire new_net_19926;
	wire new_net_14326;
	wire new_net_17947;
	wire new_net_6925;
	wire new_net_12508;
	wire new_net_15548;
	wire new_net_16045;
	wire new_net_16339;
	wire new_net_13123;
	wire new_net_13324;
	wire new_net_14864;
	wire new_net_16813;
	wire new_net_12189;
	wire new_net_14270;
	wire new_net_17596;
	wire new_net_13115;
	wire new_net_16062;
	wire new_net_8043;
	wire new_net_5882;
	wire _1747_;
	wire new_net_1998;
	wire new_net_1583;
	wire new_net_16039;
	wire new_net_16321;
	wire new_net_16684;
	wire new_net_11818;
	wire new_net_8045;
	wire new_net_6620;
	wire new_net_15803;
	wire new_net_1575;
	wire new_net_20903;
	wire new_net_13428;
	wire new_net_16513;
	wire new_net_13181;
	wire _1748_;
	wire new_net_720;
	wire new_net_5692;
	wire new_net_12818;
	wire new_net_14817;
	wire new_net_6443;
	wire new_net_5424;
	wire new_net_7032;
	wire new_net_18275;
	wire new_net_10188;
	wire new_net_19032;
	wire new_net_12866;
	wire new_net_5768;
	wire new_net_6932;
	wire new_net_10819;
	wire new_net_2436;
	wire new_net_11031;
	wire new_net_2585;
	wire new_net_11161;
	wire _1749_;
	wire new_net_717;
	wire new_net_5691;
	wire new_net_11357;
	wire new_net_17679;
	wire new_net_2426;
	wire new_net_5425;
	wire new_net_6387;
	wire new_net_9514;
	wire new_net_9515;
	wire new_net_15572;
	wire new_net_19903;
	wire new_net_19927;
	wire new_net_15849;
	wire new_net_6931;
	wire new_net_12509;
	wire new_net_13124;
	wire new_net_16814;
	wire new_net_16046;
	wire new_net_16340;
	wire new_net_11683;
	wire new_net_13325;
	wire new_net_16566;
	wire new_net_13795;
	wire new_net_21140;
	wire new_net_1573;
	wire new_net_2417;
	wire new_net_2589;
	wire new_net_3428;
	wire new_net_18268;
	wire _1575_;
	wire new_net_12908;
	wire new_net_8448;
	wire new_net_12047;
	wire new_net_4242;
	wire new_net_5297;
	wire new_net_12703;
	wire new_net_4442;
	wire new_net_10644;
	wire new_net_10667;
	wire new_net_15793;
	wire new_net_4400;
	wire new_net_13529;
	wire _1751_;
	wire new_net_2667;
	wire new_net_914;
	wire new_net_7041;
	wire new_net_20012;
	wire new_net_13550;
	wire new_net_13380;
	wire new_net_2694;
	wire new_net_4401;
	wire new_net_5472;
	wire new_net_6848;
	wire new_net_20178;
	wire new_net_17307;
	wire new_net_19097;
	wire new_net_12884;
	wire new_net_14812;
	wire new_net_18562;
	wire new_net_3434;
	wire _1752_;
	wire new_net_2699;
	wire new_net_9506;
	wire new_net_12194;
	wire new_net_11358;
	wire new_net_10820;
	wire new_net_11032;
	wire new_net_6444;
	wire new_net_11162;
	wire new_net_2437;
	wire new_net_4019;
	wire new_net_13986;
	wire _0263_;
	wire new_net_15573;
	wire new_net_6851;
	wire new_net_10649;
	wire new_net_2693;
	wire new_net_3846;
	wire new_net_1171;
	wire new_net_2418;
	wire new_net_2582;
	wire _1753_;
	wire new_net_716;
	wire new_net_10434;
	wire new_net_2523;
	wire new_net_17453;
	wire new_net_12510;
	wire new_net_13125;
	wire new_net_16047;
	wire new_net_16341;
	wire new_net_16815;
	wire new_net_11684;
	wire new_net_13326;
	wire new_net_16567;
	wire new_net_13796;
	wire new_net_6158;
	wire new_net_4025;
	wire new_net_7033;
	wire new_net_11812;
	wire new_net_8044;
	wire new_net_5880;
	wire new_net_2419;
	wire new_net_2435;
	wire _1754_;
	wire new_net_721;
	wire new_net_2664;
	wire new_net_11720;
	wire new_net_5690;
	wire new_net_15802;
	wire new_net_11817;
	wire new_net_6849;
	wire new_net_13528;
	wire new_net_909;
	wire new_net_2004;
	wire new_net_18273;
	wire new_net_20116;
	wire new_net_7578;
	wire new_net_7031;
	wire new_net_4403;
	wire _1755_;
	wire new_net_1994;
	wire new_net_6186;
	wire new_net_7673;
	wire new_net_18582;
	wire new_net_10670;
	wire new_net_3445;
	wire new_net_6622;
	wire new_net_12906;
	wire new_net_15165;
	wire new_net_15867;
	wire new_net_17757;
	wire new_net_4022;
	wire new_net_7034;
	wire new_net_11359;
	wire new_net_15577;
	wire new_net_10821;
	wire new_net_11033;
	wire new_net_11163;
	wire _1756_;
	wire new_net_10920;
	wire new_net_15524;
	wire new_net_17604;
	wire new_net_7840;
	wire new_net_18151;
	wire new_net_15574;
	wire new_net_5877;
	wire new_net_19905;
	wire new_net_19929;
	wire new_net_16811;
	wire new_net_17454;
	wire new_net_12511;
	wire new_net_13126;
	wire new_net_16816;
	wire new_net_16048;
	wire new_net_16342;
	wire new_net_11685;
	wire new_net_13327;
	wire new_net_16568;
	wire new_net_5470;
	wire new_net_14298;
	wire new_net_14206;
	wire new_net_6927;
	wire new_net_6440;
	wire new_net_1586;
	wire new_net_912;
	wire new_net_8148;
	wire _0126_;
	wire new_net_13057;
	wire new_net_9512;
	wire new_net_13527;
	wire new_net_6442;
	wire new_net_1577;
	wire _1758_;
	wire new_net_5468;
	wire new_net_20179;
	wire new_net_12807;
	wire new_net_1126;
	wire new_net_8674;
	wire new_net_14615;
	wire new_net_13351;
	wire new_net_5895;
	wire new_net_7040;
	wire new_net_910;
	wire new_net_3432;
	wire new_net_3842;
	wire new_net_17817;
	wire new_net_13806;
	wire new_net_18599;
	wire new_net_12845;
	wire new_net_6617;
	wire new_net_5476;
	wire new_net_908;
	wire _1759_;
	wire new_net_10350;
	wire new_net_19059;
	wire new_net_19201;
	wire new_net_11360;
	wire new_net_10822;
	wire new_net_11034;
	wire new_net_2433;
	wire new_net_3381;
	wire new_net_11164;
	wire new_net_15551;
	wire new_net_18271;
	wire new_net_7572;
	wire new_net_14908;
	wire new_net_18122;
	wire new_net_15387;
	wire new_net_17171;
	wire new_net_15798;
	wire _1760_;
	wire new_net_5474;
	wire new_net_5881;
	wire new_net_3436;
	wire new_net_19906;
	wire new_net_19930;
	wire new_net_15418;
	wire new_net_17455;
	wire new_net_12512;
	wire new_net_13127;
	wire new_net_16817;
	wire new_net_16049;
	wire new_net_16343;
	wire new_net_11686;
	wire new_net_13328;
	wire new_net_16569;
	wire new_net_13798;
	wire new_net_9634;
	wire new_net_16408;
	wire new_net_18321;
	wire new_net_12539;
	wire new_net_14119;
	wire new_net_9509;
	wire _1761_;
	wire new_net_2665;
	wire new_net_20173;
	wire new_net_11879;
	wire new_net_12575;
	wire _1393_;
	wire new_net_16599;
	wire new_net_15801;
	wire new_net_11816;
	wire new_net_10653;
	wire new_net_13526;
	wire new_net_2430;
	wire new_net_6623;
	wire new_net_11694;
	wire new_net_14478;
	wire new_net_12041;
	wire new_net_4362;
	wire new_net_15575;
	wire new_net_6621;
	wire new_net_5473;
	wire _1762_;
	wire new_net_723;
	wire new_net_18272;
	wire new_net_2051;
	wire new_net_18781;
	wire new_net_15231;
	wire new_net_16247;
	wire new_net_13802;
	wire new_net_19114;
	wire new_net_10646;
	wire new_net_2658;
	wire new_net_4010;
	wire new_net_4363;
	wire new_net_6382;
	wire new_net_15120;
	wire new_net_14000;
	wire new_net_5419;
	wire new_net_11165;
	wire new_net_4020;
	wire new_net_11361;
	wire new_net_10823;
	wire new_net_11035;
	wire _1763_;
	wire new_net_20180;
	wire new_net_20224;
	wire new_net_11071;
	wire new_net_15556;
	wire new_net_2666;
	wire new_net_3845;
	wire new_net_4360;
	wire new_net_6385;
	wire new_net_18267;
	wire new_net_19907;
	wire new_net_19931;
	wire new_net_14327;
	wire new_net_6033;
	wire new_net_17948;
	wire new_net_14869;
	wire new_net_15552;
	wire new_net_15794;
	wire new_net_17456;
	wire new_net_11809;
	wire new_net_12513;
	wire new_net_13128;
	wire new_net_16818;
	wire new_net_16050;
	wire new_net_16344;
	wire new_net_14271;
	wire new_net_17597;
	wire new_net_13114;
	wire new_net_6928;
	wire new_net_10651;
	wire new_net_2000;
	wire new_net_2695;
	wire new_net_16040;
	wire new_net_16322;
	wire new_net_15576;
	wire new_net_13525;
	wire new_net_5884;
	wire new_net_16685;
	wire _1765_;
	wire new_net_2692;
	wire new_net_13429;
	wire new_net_5340;
	wire new_net_9511;
	wire new_net_911;
	wire new_net_1165;
	wire new_net_3291;
	wire new_net_6645;
	wire new_net_15795;
	wire new_net_6381;
	wire new_net_6618;
	wire _1766_;
	wire new_net_2668;
	wire new_net_2700;
	wire new_net_1578;
	wire new_net_21319;
	wire new_net_12819;
	wire new_net_14818;
	wire new_net_2029;
	wire new_net_12163;
	wire new_net_19033;
	wire new_net_12867;
	wire new_net_11166;
	wire new_net_11362;
	wire new_net_15578;
	wire new_net_10824;
	wire new_net_6626;
	wire new_net_11036;
	wire new_net_2691;
	wire new_net_2416;
	wire new_net_2586;
	wire new_net_19052;
	wire new_net_17680;
	wire new_net_5422;
	wire _1767_;
	wire new_net_2689;
	wire new_net_3840;
	wire new_net_19908;
	wire new_net_19932;
	wire new_net_15850;
	wire new_net_14870;
	wire new_net_15553;
	wire new_net_17457;
	wire new_net_12514;
	wire new_net_13129;
	wire new_net_16819;
	wire new_net_10675;
	wire new_net_16051;
	wire new_net_16345;
	wire new_net_11688;
	wire new_net_9785;
	wire new_net_6379;
	wire new_net_3433;
	wire _1768_;
	wire new_net_2657;
	wire new_net_1581;
	wire new_net_2427;
	wire new_net_2434;
	wire new_net_2583;
	wire new_net_15800;
	wire new_net_11815;
	wire new_net_8036;
	wire new_net_10672;
	wire new_net_13524;
	wire new_net_1162;
	wire new_net_3431;
	wire new_net_12704;
	wire new_net_11713;
	wire new_net_16491;
	wire new_net_10184;
	wire new_net_7038;
	wire new_net_15796;
	wire _1769_;
	wire new_net_13549;
	wire new_net_20183;
	wire new_net_19098;
	wire new_net_8255;
	wire new_net_4229;
	wire new_net_6386;
	wire new_net_3841;
	wire new_net_18563;
	wire new_net_12195;
	wire new_net_11167;
	wire new_net_10825;
	wire new_net_6852;
	wire new_net_4405;
	wire new_net_11037;
	wire _1770_;
	wire new_net_2696;
	wire new_net_13987;
	wire new_net_5420;
	wire new_net_8037;
	wire new_net_1164;
	wire new_net_2580;
	wire new_net_3380;
	wire new_net_4404;
	wire new_net_19909;
	wire new_net_19933;
	wire new_net_12010;
	wire new_net_8603;
	wire new_net_12196;
	wire new_net_14871;
	wire new_net_15554;
	wire new_net_17458;
	wire new_net_12515;
	wire new_net_13130;
	wire new_net_16820;
	wire new_net_10648;
	wire new_net_16052;
	wire new_net_16346;
	wire _0056_;
	wire new_net_10645;
	wire new_net_4402;
	wire new_net_5879;
	wire new_net_7914;
	wire new_net_11721;
	wire new_net_5423;
	wire new_net_7035;
	wire new_net_11813;
	wire new_net_10650;
	wire new_net_13523;
	wire _1772_;
	wire new_net_4021;
	wire new_net_9508;
	wire new_net_11363;
	wire new_net_15579;
	wire new_net_915;
	wire new_net_20172;
	wire new_net_12340;
	wire new_net_6188;
	wire new_net_9516;
	wire new_net_11810;
	wire new_net_1579;
	wire new_net_2421;
	wire _1773_;
	wire new_net_4444;
	wire new_net_7665;
	wire new_net_18270;
	wire new_net_4280;
	wire new_net_18583;
	wire new_net_12905;
	wire new_net_10809;
	wire new_net_11168;
	wire new_net_10826;
	wire new_net_11038;
	wire new_net_2425;
	wire new_net_17758;
	wire new_net_2663;
	wire new_net_4406;
	wire new_net_15868;
	wire new_net_15525;
	wire new_net_17605;
	wire new_net_4009;
	wire new_net_4357;
	wire new_net_10647;
	wire new_net_2422;
	wire _1774_;
	wire new_net_3839;
	wire new_net_19910;
	wire new_net_19934;
	wire new_net_18152;
	wire new_net_12197;
	wire new_net_14872;
	wire new_net_15555;
	wire new_net_7036;
	wire new_net_17459;
	wire new_net_12516;
	wire new_net_13131;
	wire new_net_16821;
	wire new_net_16053;
	wire new_net_16347;
	wire new_net_6926;
	wire new_net_12507;
	wire new_net_16812;
	wire new_net_14207;
	wire new_net_8042;
	wire new_net_10676;
	wire _1775_;
	wire new_net_18266;
	wire new_net_8592;
	wire new_net_14057;
	wire new_net_13058;
	wire new_net_8675;
	wire new_net_15799;
	wire new_net_11814;
	wire new_net_13522;
	wire new_net_6845;
	wire new_net_13640;
	wire new_net_12808;
	wire new_net_14616;
	wire new_net_13352;
	wire new_net_6383;
	wire new_net_10668;
	wire new_net_5471;
	wire _1776_;
	wire new_net_715;
	wire new_net_2671;
	wire new_net_17818;
	wire new_net_13807;
	wire new_net_8504;
	wire new_net_1992;
	wire new_net_18600;
	wire new_net_5240;
	wire new_net_12846;
	wire new_net_7480;
	wire new_net_19060;
	wire new_net_11169;
	wire new_net_5426;
	wire new_net_11364;
	wire new_net_8038;
	wire new_net_11039;
	wire new_net_2002;
	wire new_net_904;
	wire _1777_;
	wire new_net_4150;
	wire new_net_19202;
	input N1;
	input N103;
	input N120;
	input N137;
	input N154;
	input N171;
	input N18;
	input N188;
	input N205;
	input N222;
	input N239;
	input N256;
	input N273;
	input N290;
	input N307;
	input N324;
	input N341;
	input N35;
	input N358;
	input N375;
	input N392;
	input N409;
	input N426;
	input N443;
	input N460;
	input N477;
	input N494;
	input N511;
	input N52;
	input N528;
	input N69;
	input N86;
	output N1581;
	output N1901;
	output N2223;
	output N2548;
	output N2877;
	output N3211;
	output N3552;
	output N3895;
	output N4241;
	output N4591;
	output N4946;
	output N5308;
	output N545;
	output N5672;
	output N5971;
	output N6123;
	output N6150;
	output N6160;
	output N6170;
	output N6180;
	output N6190;
	output N6200;
	output N6210;
	output N6220;
	output N6230;
	output N6240;
	output N6250;
	output N6260;
	output N6270;
	output N6280;
	output N6287;
	output N6288;

	and_bb _1838_ (
		.a(new_net_396),
		.b(new_net_2841),
		.c(_1458_)
	);

	and_bb _1839_ (
		.a(new_net_2551),
		.b(new_net_2907),
		.c(_1469_)
	);

	or_ii _1840_ (
		.a(new_net_3105),
		.b(new_net_3232),
		.c(_1480_)
	);

	and_bi _1841_ (
		.a(new_net_1020),
		.b(new_net_1425),
		.c(_1491_)
	);

	and_bb _1842_ (
		.a(new_net_2912),
		.b(new_net_3245),
		.c(_1502_)
	);

	or_ii _1843_ (
		.a(new_net_2552),
		.b(new_net_3093),
		.c(_1513_)
	);

	and_bi _1844_ (
		.a(new_net_2573),
		.b(new_net_488),
		.c(_1524_)
	);

	and_ii _1845_ (
		.a(new_net_3455),
		.b(new_net_254),
		.c(_1535_)
	);

	and_bb _1846_ (
		.a(new_net_2913),
		.b(new_net_2842),
		.c(new_net_0)
	);

	or_bi _1847_ (
		.a(new_net_2574),
		.b(new_net_1195),
		.c(_1556_)
	);

	or_bi _1848_ (
		.a(new_net_1908),
		.b(new_net_2754),
		.c(_1566_)
	);

	and_bb _1849_ (
		.a(new_net_36),
		.b(new_net_2833),
		.c(_1577_)
	);

	and_bi _1850_ (
		.a(new_net_1909),
		.b(new_net_2756),
		.c(_1588_)
	);

	or_bi _1851_ (
		.a(new_net_3456),
		.b(new_net_3193),
		.c(_1599_)
	);

	and_ii _1852_ (
		.a(new_net_2773),
		.b(new_net_2523),
		.c(_1610_)
	);

	and_bi _1853_ (
		.a(new_net_3194),
		.b(new_net_3123),
		.c(_1621_)
	);

	and_bb _1854_ (
		.a(new_net_2548),
		.b(new_net_49),
		.c(_1632_)
	);

	or_ii _1855_ (
		.a(new_net_741),
		.b(new_net_3094),
		.c(_1643_)
	);

	and_bi _1856_ (
		.a(new_net_489),
		.b(new_net_2880),
		.c(_1654_)
	);

	and_bb _1857_ (
		.a(new_net_737),
		.b(new_net_2917),
		.c(_1665_)
	);

	and_bi _1858_ (
		.a(new_net_1426),
		.b(new_net_2442),
		.c(_1676_)
	);

	and_ii _1859_ (
		.a(new_net_3457),
		.b(new_net_347),
		.c(_1686_)
	);

	or_bb _1860_ (
		.a(new_net_1269),
		.b(new_net_255),
		.c(_1697_)
	);

	or_ii _1861_ (
		.a(new_net_1270),
		.b(new_net_256),
		.c(_1708_)
	);

	or_ii _1862_ (
		.a(new_net_3458),
		.b(new_net_1706),
		.c(_1719_)
	);

	and_ii _1863_ (
		.a(new_net_2537),
		.b(new_net_836),
		.c(_1730_)
	);

	and_bb _1864_ (
		.a(new_net_2538),
		.b(new_net_837),
		.c(_1741_)
	);

	or_bb _1865_ (
		.a(new_net_3459),
		.b(new_net_3213),
		.c(_1752_)
	);

	or_bb _1866_ (
		.a(new_net_1586),
		.b(new_net_1886),
		.c(_1763_)
	);

	and_bb _1867_ (
		.a(new_net_1587),
		.b(new_net_1887),
		.c(_1774_)
	);

	or_bi _1868_ (
		.a(new_net_3460),
		.b(new_net_446),
		.c(_1785_)
	);

	and_ii _1869_ (
		.a(new_net_275),
		.b(new_net_620),
		.c(_1796_)
	);

	and_bb _1870_ (
		.a(new_net_276),
		.b(new_net_621),
		.c(_1806_)
	);

	or_bb _1871_ (
		.a(new_net_3461),
		.b(new_net_707),
		.c(new_net_3968)
	);

	and_bb _1872_ (
		.a(new_net_2843),
		.b(new_net_264),
		.c(_1827_)
	);

	and_bi _1873_ (
		.a(new_net_447),
		.b(new_net_708),
		.c(_0000_)
	);

	and_bb _1874_ (
		.a(new_net_2547),
		.b(new_net_403),
		.c(_0011_)
	);

	and_bi _1875_ (
		.a(new_net_1707),
		.b(new_net_3214),
		.c(_0022_)
	);

	and_bb _1876_ (
		.a(new_net_50),
		.b(new_net_3233),
		.c(_0033_)
	);

	or_ii _1877_ (
		.a(new_net_1405),
		.b(new_net_3100),
		.c(_0044_)
	);

	and_bi _1878_ (
		.a(new_net_2443),
		.b(new_net_888),
		.c(_0055_)
	);

	and_bb _1879_ (
		.a(new_net_1416),
		.b(new_net_2908),
		.c(_0066_)
	);

	and_bi _1880_ (
		.a(new_net_2881),
		.b(new_net_1632),
		.c(_0077_)
	);

	and_ii _1881_ (
		.a(new_net_3462),
		.b(new_net_1577),
		.c(_0088_)
	);

	or_bb _1882_ (
		.a(new_net_2819),
		.b(new_net_348),
		.c(_0099_)
	);

	or_ii _1883_ (
		.a(new_net_2820),
		.b(new_net_349),
		.c(_0110_)
	);

	or_ii _1884_ (
		.a(new_net_3463),
		.b(new_net_524),
		.c(_0121_)
	);

	and_ii _1885_ (
		.a(new_net_1499),
		.b(new_net_763),
		.c(_0132_)
	);

	and_bb _1886_ (
		.a(new_net_1500),
		.b(new_net_764),
		.c(_0143_)
	);

	or_bb _1887_ (
		.a(new_net_3464),
		.b(new_net_2905),
		.c(_0154_)
	);

	or_bb _1888_ (
		.a(new_net_1600),
		.b(new_net_3165),
		.c(_0165_)
	);

	or_ii _1889_ (
		.a(new_net_1601),
		.b(new_net_3166),
		.c(_0176_)
	);

	or_ii _1890_ (
		.a(new_net_3465),
		.b(new_net_460),
		.c(_0187_)
	);

	and_ii _1891_ (
		.a(new_net_88),
		.b(new_net_3226),
		.c(_0198_)
	);

	and_bb _1892_ (
		.a(new_net_89),
		.b(new_net_3227),
		.c(_0209_)
	);

	or_bb _1893_ (
		.a(new_net_3466),
		.b(new_net_2194),
		.c(_0219_)
	);

	or_bb _1894_ (
		.a(new_net_2949),
		.b(new_net_890),
		.c(_0230_)
	);

	and_bb _1895_ (
		.a(new_net_2832),
		.b(new_net_3177),
		.c(_0241_)
	);

	and_bb _1896_ (
		.a(new_net_2950),
		.b(new_net_891),
		.c(_0252_)
	);

	or_bi _1897_ (
		.a(new_net_3467),
		.b(new_net_2420),
		.c(_0263_)
	);

	and_ii _1898_ (
		.a(new_net_1485),
		.b(new_net_663),
		.c(_0274_)
	);

	and_bi _1899_ (
		.a(new_net_2421),
		.b(new_net_2985),
		.c(_0285_)
	);

	and_bb _1900_ (
		.a(new_net_2559),
		.b(new_net_3185),
		.c(_0296_)
	);

	and_bi _1901_ (
		.a(new_net_461),
		.b(new_net_2195),
		.c(_0307_)
	);

	and_bb _1902_ (
		.a(new_net_397),
		.b(new_net_3244),
		.c(_0318_)
	);

	and_bi _1903_ (
		.a(new_net_525),
		.b(new_net_2906),
		.c(_0328_)
	);

	and_bb _1904_ (
		.a(new_net_750),
		.b(new_net_42),
		.c(_0339_)
	);

	or_ii _1905_ (
		.a(new_net_1469),
		.b(new_net_3101),
		.c(_0350_)
	);

	and_bi _1906_ (
		.a(new_net_1633),
		.b(new_net_20),
		.c(_0361_)
	);

	and_bb _1907_ (
		.a(new_net_1473),
		.b(new_net_2909),
		.c(_0372_)
	);

	and_bi _1908_ (
		.a(new_net_889),
		.b(new_net_142),
		.c(_0383_)
	);

	and_ii _1909_ (
		.a(new_net_3468),
		.b(new_net_1232),
		.c(_0394_)
	);

	or_bb _1910_ (
		.a(new_net_1060),
		.b(new_net_1579),
		.c(_0405_)
	);

	or_ii _1911_ (
		.a(new_net_1061),
		.b(new_net_1578),
		.c(_0416_)
	);

	or_ii _1912_ (
		.a(new_net_3469),
		.b(new_net_3220),
		.c(_0427_)
	);

	and_ii _1913_ (
		.a(new_net_1310),
		.b(new_net_1028),
		.c(_0437_)
	);

	and_bb _1914_ (
		.a(new_net_1311),
		.b(new_net_1029),
		.c(_0448_)
	);

	or_bb _1915_ (
		.a(new_net_3470),
		.b(new_net_120),
		.c(_0459_)
	);

	or_bb _1916_ (
		.a(new_net_970),
		.b(new_net_2134),
		.c(_0470_)
	);

	or_ii _1917_ (
		.a(new_net_971),
		.b(new_net_2135),
		.c(_0481_)
	);

	or_ii _1918_ (
		.a(new_net_3471),
		.b(new_net_1340),
		.c(_0492_)
	);

	and_ii _1919_ (
		.a(new_net_1519),
		.b(new_net_287),
		.c(_0503_)
	);

	and_bb _1920_ (
		.a(new_net_1520),
		.b(new_net_288),
		.c(_0514_)
	);

	or_bb _1921_ (
		.a(new_net_3472),
		.b(new_net_356),
		.c(_0525_)
	);

	or_bb _1922_ (
		.a(new_net_2006),
		.b(new_net_2769),
		.c(_0535_)
	);

	or_ii _1923_ (
		.a(new_net_2007),
		.b(new_net_2770),
		.c(_0546_)
	);

	or_ii _1924_ (
		.a(new_net_3473),
		.b(new_net_795),
		.c(_0557_)
	);

	and_ii _1925_ (
		.a(new_net_3141),
		.b(new_net_2759),
		.c(_0568_)
	);

	and_bb _1926_ (
		.a(new_net_3142),
		.b(new_net_2760),
		.c(_0579_)
	);

	or_bb _1927_ (
		.a(new_net_3474),
		.b(new_net_1878),
		.c(_0590_)
	);

	or_bb _1928_ (
		.a(new_net_2761),
		.b(new_net_1770),
		.c(_0601_)
	);

	and_bb _1929_ (
		.a(new_net_1245),
		.b(new_net_2834),
		.c(_0612_)
	);

	and_bb _1930_ (
		.a(new_net_2762),
		.b(new_net_1771),
		.c(_0632_)
	);

	or_bi _1931_ (
		.a(new_net_3475),
		.b(new_net_301),
		.c(_0633_)
	);

	and_ii _1932_ (
		.a(new_net_1156),
		.b(new_net_1352),
		.c(_0644_)
	);

	and_bi _1933_ (
		.a(new_net_302),
		.b(new_net_30),
		.c(_0655_)
	);

	and_bb _1934_ (
		.a(new_net_2549),
		.b(new_net_1257),
		.c(_0666_)
	);

	and_bi _1935_ (
		.a(new_net_796),
		.b(new_net_1879),
		.c(_0677_)
	);

	and_bb _1936_ (
		.a(new_net_3192),
		.b(new_net_3234),
		.c(_0688_)
	);

	and_bi _1937_ (
		.a(new_net_1341),
		.b(new_net_357),
		.c(_0698_)
	);

	and_bb _1938_ (
		.a(new_net_738),
		.b(new_net_404),
		.c(_0709_)
	);

	and_bi _1939_ (
		.a(new_net_3221),
		.b(new_net_121),
		.c(_0720_)
	);

	and_bb _1940_ (
		.a(new_net_1419),
		.b(new_net_41),
		.c(_0731_)
	);

	or_ii _1941_ (
		.a(new_net_3077),
		.b(new_net_3102),
		.c(_0742_)
	);

	and_bi _1942_ (
		.a(new_net_143),
		.b(new_net_548),
		.c(_0753_)
	);

	and_bb _1943_ (
		.a(new_net_3089),
		.b(new_net_2910),
		.c(_0764_)
	);

	and_bi _1944_ (
		.a(new_net_21),
		.b(new_net_182),
		.c(_0774_)
	);

	and_ii _1945_ (
		.a(new_net_3476),
		.b(new_net_1295),
		.c(_0785_)
	);

	or_bb _1946_ (
		.a(new_net_602),
		.b(new_net_1234),
		.c(_0796_)
	);

	or_ii _1947_ (
		.a(new_net_603),
		.b(new_net_1233),
		.c(_0807_)
	);

	or_ii _1948_ (
		.a(new_net_3477),
		.b(new_net_2476),
		.c(_0818_)
	);

	and_ii _1949_ (
		.a(new_net_1780),
		.b(new_net_126),
		.c(_0828_)
	);

	and_bb _1950_ (
		.a(new_net_1781),
		.b(new_net_127),
		.c(_0839_)
	);

	or_bb _1951_ (
		.a(new_net_3478),
		.b(new_net_1038),
		.c(_0850_)
	);

	or_bb _1952_ (
		.a(new_net_3115),
		.b(new_net_2933),
		.c(_0861_)
	);

	or_ii _1953_ (
		.a(new_net_3116),
		.b(new_net_2934),
		.c(_0872_)
	);

	or_ii _1954_ (
		.a(new_net_3479),
		.b(new_net_1840),
		.c(_0882_)
	);

	and_ii _1955_ (
		.a(new_net_2669),
		.b(new_net_868),
		.c(_0893_)
	);

	and_bb _1956_ (
		.a(new_net_2670),
		.b(new_net_869),
		.c(_0904_)
	);

	or_bb _1957_ (
		.a(new_net_3480),
		.b(new_net_3143),
		.c(_0915_)
	);

	or_bb _1958_ (
		.a(new_net_757),
		.b(new_net_470),
		.c(_0925_)
	);

	or_ii _1959_ (
		.a(new_net_758),
		.b(new_net_471),
		.c(_0936_)
	);

	or_ii _1960_ (
		.a(new_net_3481),
		.b(new_net_345),
		.c(_0947_)
	);

	and_ii _1961_ (
		.a(new_net_138),
		.b(new_net_102),
		.c(_0958_)
	);

	and_bb _1962_ (
		.a(new_net_139),
		.b(new_net_103),
		.c(_0968_)
	);

	or_bb _1963_ (
		.a(new_net_3482),
		.b(new_net_358),
		.c(_0979_)
	);

	or_bb _1964_ (
		.a(new_net_3262),
		.b(new_net_2418),
		.c(_0989_)
	);

	or_ii _1965_ (
		.a(new_net_3263),
		.b(new_net_2419),
		.c(_1000_)
	);

	or_ii _1966_ (
		.a(new_net_3483),
		.b(new_net_2216),
		.c(_1010_)
	);

	and_ii _1967_ (
		.a(new_net_3041),
		.b(new_net_327),
		.c(_1013_)
	);

	and_bb _1968_ (
		.a(new_net_3042),
		.b(new_net_328),
		.c(_1014_)
	);

	or_bb _1969_ (
		.a(new_net_3484),
		.b(new_net_2855),
		.c(_1015_)
	);

	or_bb _1970_ (
		.a(new_net_787),
		.b(new_net_1439),
		.c(_1016_)
	);

	and_bb _1971_ (
		.a(new_net_1449),
		.b(new_net_2829),
		.c(_1017_)
	);

	and_bb _1972_ (
		.a(new_net_788),
		.b(new_net_1440),
		.c(_1018_)
	);

	or_bi _1973_ (
		.a(new_net_3485),
		.b(new_net_2995),
		.c(_1019_)
	);

	and_ii _1974_ (
		.a(new_net_1509),
		.b(new_net_1092),
		.c(_1020_)
	);

	and_bi _1975_ (
		.a(new_net_2996),
		.b(new_net_1672),
		.c(_1021_)
	);

	and_bb _1976_ (
		.a(new_net_2560),
		.b(new_net_1447),
		.c(_1022_)
	);

	and_bi _1977_ (
		.a(new_net_2217),
		.b(new_net_2856),
		.c(_1023_)
	);

	and_bb _1978_ (
		.a(new_net_1253),
		.b(new_net_3246),
		.c(_1024_)
	);

	and_bi _1979_ (
		.a(new_net_346),
		.b(new_net_359),
		.c(_1025_)
	);

	and_bb _1980_ (
		.a(new_net_751),
		.b(new_net_3183),
		.c(_1026_)
	);

	and_bi _1981_ (
		.a(new_net_1841),
		.b(new_net_3144),
		.c(_1027_)
	);

	and_bb _1982_ (
		.a(new_net_1414),
		.b(new_net_405),
		.c(_1028_)
	);

	and_bi _1983_ (
		.a(new_net_2477),
		.b(new_net_1039),
		.c(_1029_)
	);

	and_bb _1984_ (
		.a(new_net_1482),
		.b(new_net_43),
		.c(_1030_)
	);

	or_ii _1985_ (
		.a(new_net_2339),
		.b(new_net_3103),
		.c(_1031_)
	);

	and_bi _1986_ (
		.a(new_net_183),
		.b(new_net_335),
		.c(_1032_)
	);

	and_bb _1987_ (
		.a(new_net_2344),
		.b(new_net_2911),
		.c(_1033_)
	);

	and_bi _1988_ (
		.a(new_net_549),
		.b(new_net_422),
		.c(_1034_)
	);

	and_ii _1989_ (
		.a(new_net_3486),
		.b(new_net_2890),
		.c(_1035_)
	);

	or_bb _1990_ (
		.a(new_net_506),
		.b(new_net_1296),
		.c(_1036_)
	);

	or_ii _1991_ (
		.a(new_net_507),
		.b(new_net_1297),
		.c(_1037_)
	);

	or_ii _1992_ (
		.a(new_net_3487),
		.b(new_net_444),
		.c(_1038_)
	);

	and_ii _1993_ (
		.a(new_net_626),
		.b(new_net_303),
		.c(_1039_)
	);

	and_bb _1994_ (
		.a(new_net_627),
		.b(new_net_304),
		.c(_1040_)
	);

	or_bb _1995_ (
		.a(new_net_3488),
		.b(new_net_655),
		.c(_1041_)
	);

	or_bb _1996_ (
		.a(new_net_771),
		.b(new_net_2276),
		.c(_1042_)
	);

	or_ii _1997_ (
		.a(new_net_772),
		.b(new_net_2277),
		.c(_1043_)
	);

	or_ii _1998_ (
		.a(new_net_3489),
		.b(new_net_1590),
		.c(_1044_)
	);

	and_ii _1999_ (
		.a(new_net_1902),
		.b(new_net_2096),
		.c(_1045_)
	);

	and_bb _2000_ (
		.a(new_net_1903),
		.b(new_net_2097),
		.c(_1046_)
	);

	or_bb _2001_ (
		.a(new_net_3490),
		.b(new_net_2102),
		.c(_1047_)
	);

	or_bb _2002_ (
		.a(new_net_968),
		.b(new_net_1894),
		.c(_1048_)
	);

	or_ii _2003_ (
		.a(new_net_969),
		.b(new_net_1895),
		.c(_1049_)
	);

	or_ii _2004_ (
		.a(new_net_3491),
		.b(new_net_1000),
		.c(_1050_)
	);

	and_ii _2005_ (
		.a(new_net_3135),
		.b(new_net_168),
		.c(_1051_)
	);

	and_bb _2006_ (
		.a(new_net_3136),
		.b(new_net_169),
		.c(_1052_)
	);

	or_bb _2007_ (
		.a(new_net_3492),
		.b(new_net_1076),
		.c(_1053_)
	);

	or_bb _2008_ (
		.a(new_net_450),
		.b(new_net_1584),
		.c(_1054_)
	);

	or_ii _2009_ (
		.a(new_net_451),
		.b(new_net_1585),
		.c(_1055_)
	);

	or_ii _2010_ (
		.a(new_net_3493),
		.b(new_net_1184),
		.c(_1056_)
	);

	and_ii _2011_ (
		.a(new_net_1004),
		.b(new_net_96),
		.c(_1057_)
	);

	and_bb _2012_ (
		.a(new_net_1005),
		.b(new_net_97),
		.c(_1058_)
	);

	or_bb _2013_ (
		.a(new_net_3494),
		.b(new_net_1312),
		.c(_1059_)
	);

	or_bb _2014_ (
		.a(new_net_1596),
		.b(new_net_1158),
		.c(_1060_)
	);

	or_ii _2015_ (
		.a(new_net_1597),
		.b(new_net_1159),
		.c(_1061_)
	);

	or_ii _2016_ (
		.a(new_net_3495),
		.b(new_net_1403),
		.c(_1062_)
	);

	and_ii _2017_ (
		.a(new_net_2106),
		.b(new_net_998),
		.c(_1063_)
	);

	and_bb _2018_ (
		.a(new_net_2107),
		.b(new_net_999),
		.c(_1064_)
	);

	or_bb _2019_ (
		.a(new_net_3496),
		.b(new_net_2292),
		.c(_1065_)
	);

	or_bb _2020_ (
		.a(new_net_1650),
		.b(new_net_1830),
		.c(_1066_)
	);

	and_bb _2021_ (
		.a(new_net_1796),
		.b(new_net_2835),
		.c(_1067_)
	);

	and_bb _2022_ (
		.a(new_net_1651),
		.b(new_net_1831),
		.c(_1068_)
	);

	or_bi _2023_ (
		.a(new_net_3497),
		.b(new_net_1686),
		.c(_1069_)
	);

	and_ii _2024_ (
		.a(new_net_1752),
		.b(new_net_1702),
		.c(_1070_)
	);

	and_bi _2025_ (
		.a(new_net_1687),
		.b(new_net_1790),
		.c(_1071_)
	);

	and_bb _2026_ (
		.a(new_net_2550),
		.b(new_net_1810),
		.c(_1072_)
	);

	and_bi _2027_ (
		.a(new_net_1404),
		.b(new_net_2293),
		.c(_1073_)
	);

	and_bb _2028_ (
		.a(new_net_1454),
		.b(new_net_3235),
		.c(_1074_)
	);

	and_bi _2029_ (
		.a(new_net_1185),
		.b(new_net_1313),
		.c(_1075_)
	);

	and_bb _2030_ (
		.a(new_net_739),
		.b(new_net_1258),
		.c(_1076_)
	);

	and_bi _2031_ (
		.a(new_net_1001),
		.b(new_net_1077),
		.c(_1077_)
	);

	and_bb _2032_ (
		.a(new_net_1418),
		.b(new_net_3184),
		.c(_1078_)
	);

	and_bi _2033_ (
		.a(new_net_1591),
		.b(new_net_2103),
		.c(_1079_)
	);

	and_bb _2034_ (
		.a(new_net_1471),
		.b(new_net_406),
		.c(_1080_)
	);

	and_bi _2035_ (
		.a(new_net_445),
		.b(new_net_656),
		.c(_1081_)
	);

	and_bb _2036_ (
		.a(new_net_3091),
		.b(new_net_44),
		.c(_1082_)
	);

	or_ii _2037_ (
		.a(new_net_3095),
		.b(new_net_2400),
		.c(_1083_)
	);

	and_bi _2038_ (
		.a(new_net_423),
		.b(new_net_2206),
		.c(_1084_)
	);

	and_bb _2039_ (
		.a(new_net_2918),
		.b(new_net_2396),
		.c(_1085_)
	);

	and_bi _2040_ (
		.a(new_net_336),
		.b(new_net_2621),
		.c(_1086_)
	);

	and_ii _2041_ (
		.a(new_net_3498),
		.b(new_net_2363),
		.c(_1087_)
	);

	or_bb _2042_ (
		.a(new_net_2452),
		.b(new_net_2892),
		.c(_1088_)
	);

	or_ii _2043_ (
		.a(new_net_2453),
		.b(new_net_2891),
		.c(_1089_)
	);

	or_ii _2044_ (
		.a(new_net_3499),
		.b(new_net_3274),
		.c(_1090_)
	);

	and_ii _2045_ (
		.a(new_net_329),
		.b(new_net_1990),
		.c(_1091_)
	);

	and_bb _2046_ (
		.a(new_net_330),
		.b(new_net_1991),
		.c(_1092_)
	);

	or_bb _2047_ (
		.a(new_net_3500),
		.b(new_net_2649),
		.c(_1093_)
	);

	or_bb _2048_ (
		.a(new_net_932),
		.b(new_net_2230),
		.c(_1094_)
	);

	or_ii _2049_ (
		.a(new_net_933),
		.b(new_net_2231),
		.c(_1095_)
	);

	or_ii _2050_ (
		.a(new_net_3501),
		.b(new_net_1070),
		.c(_1096_)
	);

	and_ii _2051_ (
		.a(new_net_1495),
		.b(new_net_1656),
		.c(_1097_)
	);

	and_bb _2052_ (
		.a(new_net_1496),
		.b(new_net_1657),
		.c(_1098_)
	);

	or_bb _2053_ (
		.a(new_net_3502),
		.b(new_net_2849),
		.c(_1099_)
	);

	or_bb _2054_ (
		.a(new_net_2969),
		.b(new_net_1457),
		.c(_1100_)
	);

	or_ii _2055_ (
		.a(new_net_2970),
		.b(new_net_1458),
		.c(_1101_)
	);

	or_ii _2056_ (
		.a(new_net_3503),
		.b(new_net_2212),
		.c(_1102_)
	);

	and_ii _2057_ (
		.a(new_net_2625),
		.b(new_net_1261),
		.c(_1103_)
	);

	and_bb _2058_ (
		.a(new_net_2626),
		.b(new_net_1262),
		.c(_1104_)
	);

	or_bb _2059_ (
		.a(new_net_3504),
		.b(new_net_3147),
		.c(_1105_)
	);

	or_bb _2060_ (
		.a(new_net_3248),
		.b(new_net_2066),
		.c(_1106_)
	);

	or_ii _2061_ (
		.a(new_net_3249),
		.b(new_net_2067),
		.c(_1107_)
	);

	or_ii _2062_ (
		.a(new_net_3505),
		.b(new_net_32),
		.c(_1108_)
	);

	and_ii _2063_ (
		.a(new_net_2138),
		.b(new_net_2014),
		.c(_1109_)
	);

	and_bb _2064_ (
		.a(new_net_2139),
		.b(new_net_2015),
		.c(_1110_)
	);

	or_bb _2065_ (
		.a(new_net_3506),
		.b(new_net_2333),
		.c(_1111_)
	);

	or_bb _2066_ (
		.a(new_net_2742),
		.b(new_net_733),
		.c(_1112_)
	);

	or_ii _2067_ (
		.a(new_net_2743),
		.b(new_net_734),
		.c(_1113_)
	);

	or_ii _2068_ (
		.a(new_net_3507),
		.b(new_net_2951),
		.c(_1114_)
	);

	and_ii _2069_ (
		.a(new_net_112),
		.b(new_net_522),
		.c(_1115_)
	);

	and_bb _2070_ (
		.a(new_net_113),
		.b(new_net_523),
		.c(_1116_)
	);

	or_bb _2071_ (
		.a(new_net_3508),
		.b(new_net_289),
		.c(_1117_)
	);

	or_bb _2072_ (
		.a(new_net_424),
		.b(new_net_1922),
		.c(_1118_)
	);

	or_ii _2073_ (
		.a(new_net_425),
		.b(new_net_1923),
		.c(_1119_)
	);

	or_ii _2074_ (
		.a(new_net_3509),
		.b(new_net_464),
		.c(_1120_)
	);

	and_ii _2075_ (
		.a(new_net_1192),
		.b(new_net_1874),
		.c(_1121_)
	);

	and_bb _2076_ (
		.a(new_net_1193),
		.b(new_net_1875),
		.c(_1122_)
	);

	or_bb _2077_ (
		.a(new_net_3510),
		.b(new_net_1390),
		.c(_1123_)
	);

	or_bb _2078_ (
		.a(new_net_1748),
		.b(new_net_3270),
		.c(_1124_)
	);

	and_bb _2079_ (
		.a(new_net_209),
		.b(new_net_2830),
		.c(_1125_)
	);

	and_bb _2080_ (
		.a(new_net_1749),
		.b(new_net_3271),
		.c(_1126_)
	);

	or_bi _2081_ (
		.a(new_net_3511),
		.b(new_net_1934),
		.c(_1127_)
	);

	and_ii _2082_ (
		.a(new_net_856),
		.b(new_net_2146),
		.c(_1128_)
	);

	and_bi _2083_ (
		.a(new_net_1935),
		.b(new_net_876),
		.c(_1129_)
	);

	and_bb _2084_ (
		.a(new_net_2561),
		.b(new_net_206),
		.c(_1130_)
	);

	and_bi _2085_ (
		.a(new_net_465),
		.b(new_net_1391),
		.c(_1131_)
	);

	and_bb _2086_ (
		.a(new_net_1802),
		.b(new_net_3247),
		.c(_1132_)
	);

	and_bi _2087_ (
		.a(new_net_2952),
		.b(new_net_290),
		.c(_1133_)
	);

	and_bb _2088_ (
		.a(new_net_752),
		.b(new_net_1446),
		.c(_1134_)
	);

	and_bi _2089_ (
		.a(new_net_33),
		.b(new_net_2334),
		.c(_1135_)
	);

	and_bb _2090_ (
		.a(new_net_1415),
		.b(new_net_1259),
		.c(_1136_)
	);

	and_bi _2091_ (
		.a(new_net_2213),
		.b(new_net_3148),
		.c(_1137_)
	);

	and_bb _2092_ (
		.a(new_net_1483),
		.b(new_net_3186),
		.c(_1138_)
	);

	and_bi _2093_ (
		.a(new_net_1071),
		.b(new_net_2850),
		.c(_1139_)
	);

	and_bb _2094_ (
		.a(new_net_3087),
		.b(new_net_407),
		.c(_1140_)
	);

	and_bi _2095_ (
		.a(new_net_3275),
		.b(new_net_2650),
		.c(_1141_)
	);

	and_bb _2096_ (
		.a(new_net_2353),
		.b(new_net_45),
		.c(_1142_)
	);

	or_ii _2097_ (
		.a(new_net_3096),
		.b(new_net_384),
		.c(_1143_)
	);

	and_bi _2098_ (
		.a(new_net_2622),
		.b(new_net_1368),
		.c(_1144_)
	);

	and_bb _2099_ (
		.a(new_net_2919),
		.b(new_net_378),
		.c(_1145_)
	);

	and_bi _2100_ (
		.a(new_net_2207),
		.b(new_net_1467),
		.c(_1146_)
	);

	and_ii _2101_ (
		.a(new_net_3512),
		.b(new_net_1400),
		.c(_1147_)
	);

	or_bb _2102_ (
		.a(new_net_3205),
		.b(new_net_2365),
		.c(_1148_)
	);

	or_ii _2103_ (
		.a(new_net_3206),
		.b(new_net_2364),
		.c(_1149_)
	);

	or_ii _2104_ (
		.a(new_net_3513),
		.b(new_net_1900),
		.c(_1150_)
	);

	and_ii _2105_ (
		.a(new_net_2282),
		.b(new_net_2166),
		.c(_1151_)
	);

	and_bb _2106_ (
		.a(new_net_2283),
		.b(new_net_2167),
		.c(_1152_)
	);

	or_bb _2107_ (
		.a(new_net_3514),
		.b(new_net_2480),
		.c(_1153_)
	);

	or_bb _2108_ (
		.a(new_net_2897),
		.b(new_net_1318),
		.c(_1154_)
	);

	or_ii _2109_ (
		.a(new_net_2898),
		.b(new_net_1319),
		.c(_1155_)
	);

	or_ii _2110_ (
		.a(new_net_3515),
		.b(new_net_1786),
		.c(_1156_)
	);

	and_ii _2111_ (
		.a(new_net_1872),
		.b(new_net_1275),
		.c(_1157_)
	);

	and_bb _2112_ (
		.a(new_net_1873),
		.b(new_net_1276),
		.c(_1158_)
	);

	or_bb _2113_ (
		.a(new_net_3516),
		.b(new_net_448),
		.c(_1159_)
	);

	or_bb _2114_ (
		.a(new_net_1986),
		.b(new_net_1206),
		.c(_1160_)
	);

	or_ii _2115_ (
		.a(new_net_1987),
		.b(new_net_1207),
		.c(_1161_)
	);

	or_ii _2116_ (
		.a(new_net_3517),
		.b(new_net_1002),
		.c(_1162_)
	);

	and_ii _2117_ (
		.a(new_net_1358),
		.b(new_net_1178),
		.c(_1163_)
	);

	and_bb _2118_ (
		.a(new_net_1359),
		.b(new_net_1179),
		.c(_1164_)
	);

	or_bb _2119_ (
		.a(new_net_3518),
		.b(new_net_1594),
		.c(_1165_)
	);

	or_bb _2120_ (
		.a(new_net_2240),
		.b(new_net_1202),
		.c(_1166_)
	);

	or_ii _2121_ (
		.a(new_net_2241),
		.b(new_net_1203),
		.c(_1167_)
	);

	or_ii _2122_ (
		.a(new_net_3519),
		.b(new_net_2104),
		.c(_1168_)
	);

	and_ii _2123_ (
		.a(new_net_2357),
		.b(new_net_1110),
		.c(_1169_)
	);

	and_bb _2124_ (
		.a(new_net_2358),
		.b(new_net_1111),
		.c(_1170_)
	);

	or_bb _2125_ (
		.a(new_net_3520),
		.b(new_net_2412),
		.c(_1171_)
	);

	or_bb _2126_ (
		.a(new_net_2454),
		.b(new_net_1072),
		.c(_1172_)
	);

	or_ii _2127_ (
		.a(new_net_2455),
		.b(new_net_1073),
		.c(_1173_)
	);

	or_ii _2128_ (
		.a(new_net_3521),
		.b(new_net_2484),
		.c(_1174_)
	);

	and_ii _2129_ (
		.a(new_net_454),
		.b(new_net_681),
		.c(_1175_)
	);

	and_bb _2130_ (
		.a(new_net_455),
		.b(new_net_682),
		.c(_1176_)
	);

	or_bb _2131_ (
		.a(new_net_3522),
		.b(new_net_641),
		.c(_1177_)
	);

	or_bb _2132_ (
		.a(new_net_2716),
		.b(new_net_486),
		.c(_1178_)
	);

	or_ii _2133_ (
		.a(new_net_2717),
		.b(new_net_487),
		.c(_1179_)
	);

	or_ii _2134_ (
		.a(new_net_3523),
		.b(new_net_2757),
		.c(_1180_)
	);

	and_ii _2135_ (
		.a(new_net_1598),
		.b(new_net_293),
		.c(_1181_)
	);

	and_bb _2136_ (
		.a(new_net_1599),
		.b(new_net_294),
		.c(_1182_)
	);

	or_bb _2137_ (
		.a(new_net_3524),
		.b(new_net_2851),
		.c(_1183_)
	);

	or_bb _2138_ (
		.a(new_net_2126),
		.b(new_net_966),
		.c(_1184_)
	);

	or_ii _2139_ (
		.a(new_net_2127),
		.b(new_net_967),
		.c(_1185_)
	);

	or_ii _2140_ (
		.a(new_net_3525),
		.b(new_net_2315),
		.c(_1186_)
	);

	and_ii _2141_ (
		.a(new_net_2736),
		.b(new_net_938),
		.c(_1187_)
	);

	and_bb _2142_ (
		.a(new_net_2737),
		.b(new_net_939),
		.c(_1188_)
	);

	or_bb _2143_ (
		.a(new_net_3526),
		.b(new_net_2931),
		.c(_1189_)
	);

	or_bb _2144_ (
		.a(new_net_86),
		.b(new_net_2973),
		.c(_1190_)
	);

	and_bb _2145_ (
		.a(new_net_87),
		.b(new_net_2974),
		.c(_1191_)
	);

	or_bi _2146_ (
		.a(new_net_3527),
		.b(new_net_492),
		.c(_1192_)
	);

	and_ii _2147_ (
		.a(new_net_98),
		.b(new_net_814),
		.c(_1193_)
	);

	and_bb _2148_ (
		.a(new_net_99),
		.b(new_net_815),
		.c(_1194_)
	);

	or_bb _2149_ (
		.a(new_net_3528),
		.b(new_net_1036),
		.c(new_net_3956)
	);

	or_ii _2150_ (
		.a(new_net_3097),
		.b(new_net_2844),
		.c(_1195_)
	);

	and_bi _2151_ (
		.a(new_net_3529),
		.b(new_net_1021),
		.c(_1196_)
	);

	and_bi _2152_ (
		.a(new_net_2755),
		.b(new_net_3530),
		.c(new_net_3958)
	);

	and_bb _2153_ (
		.a(new_net_2774),
		.b(new_net_2524),
		.c(_1197_)
	);

	or_bb _2154_ (
		.a(new_net_3531),
		.b(new_net_3124),
		.c(new_net_3930)
	);

	and_bb _2155_ (
		.a(new_net_1510),
		.b(new_net_1093),
		.c(_1198_)
	);

	or_bb _2156_ (
		.a(new_net_3532),
		.b(new_net_1673),
		.c(new_net_3950)
	);

	and_bb _2157_ (
		.a(new_net_857),
		.b(new_net_2147),
		.c(_1199_)
	);

	or_bb _2158_ (
		.a(new_net_3533),
		.b(new_net_877),
		.c(new_net_3928)
	);

	and_bb _2159_ (
		.a(new_net_1753),
		.b(new_net_1703),
		.c(_1200_)
	);

	or_bb _2160_ (
		.a(new_net_3534),
		.b(new_net_1791),
		.c(new_net_3932)
	);

	and_bb _2161_ (
		.a(new_net_1157),
		.b(new_net_1353),
		.c(_1201_)
	);

	or_bb _2162_ (
		.a(new_net_3535),
		.b(new_net_31),
		.c(new_net_3954)
	);

	and_bb _2163_ (
		.a(new_net_1486),
		.b(new_net_664),
		.c(_1202_)
	);

	or_bb _2164_ (
		.a(new_net_3536),
		.b(new_net_2986),
		.c(new_net_3974)
	);

	and_bb _2165_ (
		.a(new_net_2605),
		.b(new_net_2836),
		.c(_1203_)
	);

	and_bi _2166_ (
		.a(new_net_493),
		.b(new_net_1037),
		.c(_1204_)
	);

	and_bb _2167_ (
		.a(new_net_2553),
		.b(new_net_259),
		.c(_1205_)
	);

	and_bi _2168_ (
		.a(new_net_2316),
		.b(new_net_2932),
		.c(_1206_)
	);

	and_bb _2169_ (
		.a(new_net_201),
		.b(new_net_3236),
		.c(_1207_)
	);

	and_bi _2170_ (
		.a(new_net_2758),
		.b(new_net_2852),
		.c(_1208_)
	);

	and_bb _2171_ (
		.a(new_net_742),
		.b(new_net_1797),
		.c(_1209_)
	);

	and_bi _2172_ (
		.a(new_net_2485),
		.b(new_net_642),
		.c(_1210_)
	);

	and_bb _2173_ (
		.a(new_net_1406),
		.b(new_net_1450),
		.c(_1211_)
	);

	and_bi _2174_ (
		.a(new_net_2105),
		.b(new_net_2413),
		.c(_1212_)
	);

	and_bb _2175_ (
		.a(new_net_1474),
		.b(new_net_1246),
		.c(_1213_)
	);

	and_bi _2176_ (
		.a(new_net_1003),
		.b(new_net_1595),
		.c(_1214_)
	);

	and_bb _2177_ (
		.a(new_net_3078),
		.b(new_net_3189),
		.c(_1215_)
	);

	and_bi _2178_ (
		.a(new_net_1787),
		.b(new_net_449),
		.c(_1216_)
	);

	and_bb _2179_ (
		.a(new_net_2343),
		.b(new_net_392),
		.c(_1217_)
	);

	and_bi _2180_ (
		.a(new_net_1901),
		.b(new_net_2481),
		.c(_1218_)
	);

	and_bb _2181_ (
		.a(new_net_37),
		.b(new_net_2401),
		.c(_1219_)
	);

	or_ii _2182_ (
		.a(new_net_2498),
		.b(new_net_3106),
		.c(_1220_)
	);

	and_bi _2183_ (
		.a(new_net_1468),
		.b(new_net_2987),
		.c(_1221_)
	);

	and_bb _2184_ (
		.a(new_net_2502),
		.b(new_net_2914),
		.c(_1222_)
	);

	and_bi _2185_ (
		.a(new_net_1369),
		.b(new_net_1174),
		.c(_1223_)
	);

	and_ii _2186_ (
		.a(new_net_3537),
		.b(new_net_3217),
		.c(_1224_)
	);

	or_bb _2187_ (
		.a(new_net_510),
		.b(new_net_1401),
		.c(_1225_)
	);

	or_ii _2188_ (
		.a(new_net_511),
		.b(new_net_1402),
		.c(_1226_)
	);

	or_ii _2189_ (
		.a(new_net_3538),
		.b(new_net_719),
		.c(_1227_)
	);

	and_ii _2190_ (
		.a(new_net_1374),
		.b(new_net_1082),
		.c(_1228_)
	);

	and_bb _2191_ (
		.a(new_net_1375),
		.b(new_net_1083),
		.c(_1229_)
	);

	or_bb _2192_ (
		.a(new_net_3539),
		.b(new_net_1230),
		.c(_1230_)
	);

	or_bb _2193_ (
		.a(new_net_1527),
		.b(new_net_1052),
		.c(_1231_)
	);

	or_ii _2194_ (
		.a(new_net_1528),
		.b(new_net_1053),
		.c(_1232_)
	);

	or_ii _2195_ (
		.a(new_net_3540),
		.b(new_net_1567),
		.c(_1233_)
	);

	and_ii _2196_ (
		.a(new_net_1652),
		.b(new_net_1016),
		.c(_1234_)
	);

	and_bb _2197_ (
		.a(new_net_1653),
		.b(new_net_1017),
		.c(_1235_)
	);

	or_bb _2198_ (
		.a(new_net_3541),
		.b(new_net_1678),
		.c(_1236_)
	);

	or_bb _2199_ (
		.a(new_net_1734),
		.b(new_net_2174),
		.c(_1237_)
	);

	or_ii _2200_ (
		.a(new_net_1735),
		.b(new_net_2175),
		.c(_1238_)
	);

	or_ii _2201_ (
		.a(new_net_3542),
		.b(new_net_1162),
		.c(_1239_)
	);

	and_ii _2202_ (
		.a(new_net_1842),
		.b(new_net_1964),
		.c(_1240_)
	);

	and_bb _2203_ (
		.a(new_net_1843),
		.b(new_net_1965),
		.c(_1241_)
	);

	or_bb _2204_ (
		.a(new_net_3543),
		.b(new_net_1716),
		.c(_1242_)
	);

	or_bb _2205_ (
		.a(new_net_1952),
		.b(new_net_1768),
		.c(_1243_)
	);

	or_ii _2206_ (
		.a(new_net_1953),
		.b(new_net_1769),
		.c(_1244_)
	);

	or_ii _2207_ (
		.a(new_net_3544),
		.b(new_net_2278),
		.c(_1245_)
	);

	and_ii _2208_ (
		.a(new_net_2693),
		.b(new_net_896),
		.c(_1246_)
	);

	and_bb _2209_ (
		.a(new_net_2694),
		.b(new_net_897),
		.c(_1247_)
	);

	or_bb _2210_ (
		.a(new_net_3545),
		.b(new_net_2895),
		.c(_1248_)
	);

	or_bb _2211_ (
		.a(new_net_2200),
		.b(new_net_872),
		.c(_1249_)
	);

	or_ii _2212_ (
		.a(new_net_2201),
		.b(new_net_873),
		.c(_1250_)
	);

	or_ii _2213_ (
		.a(new_net_3546),
		.b(new_net_2238),
		.c(_1251_)
	);

	and_ii _2214_ (
		.a(new_net_2309),
		.b(new_net_1212),
		.c(_1252_)
	);

	and_bb _2215_ (
		.a(new_net_2310),
		.b(new_net_1213),
		.c(_1253_)
	);

	or_bb _2216_ (
		.a(new_net_3547),
		.b(new_net_862),
		.c(_1254_)
	);

	or_bb _2217_ (
		.a(new_net_2430),
		.b(new_net_1034),
		.c(_1255_)
	);

	or_ii _2218_ (
		.a(new_net_2431),
		.b(new_net_1035),
		.c(_1256_)
	);

	or_ii _2219_ (
		.a(new_net_3548),
		.b(new_net_1356),
		.c(_1257_)
	);

	and_ii _2220_ (
		.a(new_net_2541),
		.b(new_net_894),
		.c(_1258_)
	);

	and_bb _2221_ (
		.a(new_net_2542),
		.b(new_net_895),
		.c(_1259_)
	);

	or_bb _2222_ (
		.a(new_net_3549),
		.b(new_net_1906),
		.c(_1260_)
	);

	or_bb _2223_ (
		.a(new_net_2288),
		.b(new_net_693),
		.c(_1261_)
	);

	or_ii _2224_ (
		.a(new_net_2289),
		.b(new_net_694),
		.c(_1262_)
	);

	or_ii _2225_ (
		.a(new_net_3550),
		.b(new_net_2714),
		.c(_1263_)
	);

	and_ii _2226_ (
		.a(new_net_2777),
		.b(new_net_496),
		.c(_1264_)
	);

	and_bb _2227_ (
		.a(new_net_2778),
		.b(new_net_497),
		.c(_1265_)
	);

	or_bb _2228_ (
		.a(new_net_3551),
		.b(new_net_3153),
		.c(_1266_)
	);

	or_bb _2229_ (
		.a(new_net_248),
		.b(new_net_299),
		.c(_1267_)
	);

	or_ii _2230_ (
		.a(new_net_249),
		.b(new_net_300),
		.c(_1268_)
	);

	or_ii _2231_ (
		.a(new_net_3552),
		.b(new_net_2965),
		.c(_1269_)
	);

	and_ii _2232_ (
		.a(new_net_864),
		.b(new_net_116),
		.c(_1270_)
	);

	and_bb _2233_ (
		.a(new_net_865),
		.b(new_net_117),
		.c(_1271_)
	);

	or_bb _2234_ (
		.a(new_net_3553),
		.b(new_net_3111),
		.c(_1272_)
	);

	or_bb _2235_ (
		.a(new_net_3175),
		.b(new_net_3211),
		.c(_1273_)
	);

	and_bb _2236_ (
		.a(new_net_3176),
		.b(new_net_3212),
		.c(_1274_)
	);

	or_bi _2237_ (
		.a(new_net_3554),
		.b(new_net_3230),
		.c(_1275_)
	);

	and_ii _2238_ (
		.a(new_net_72),
		.b(new_net_2981),
		.c(_1276_)
	);

	and_bb _2239_ (
		.a(new_net_73),
		.b(new_net_2982),
		.c(_1277_)
	);

	or_bb _2240_ (
		.a(new_net_3555),
		.b(new_net_2882),
		.c(new_net_3922)
	);

	and_bb _2241_ (
		.a(new_net_3011),
		.b(new_net_2837),
		.c(_1278_)
	);

	and_bi _2242_ (
		.a(new_net_3231),
		.b(new_net_2883),
		.c(_1279_)
	);

	and_bb _2243_ (
		.a(new_net_2554),
		.b(new_net_2608),
		.c(_1280_)
	);

	and_bi _2244_ (
		.a(new_net_2966),
		.b(new_net_3112),
		.c(_1281_)
	);

	and_bb _2245_ (
		.a(new_net_258),
		.b(new_net_3237),
		.c(_1282_)
	);

	and_bi _2246_ (
		.a(new_net_2715),
		.b(new_net_3154),
		.c(_1283_)
	);

	and_bb _2247_ (
		.a(new_net_743),
		.b(new_net_200),
		.c(_1284_)
	);

	and_bi _2248_ (
		.a(new_net_1357),
		.b(new_net_1907),
		.c(_1285_)
	);

	and_bb _2249_ (
		.a(new_net_1407),
		.b(new_net_1804),
		.c(_1286_)
	);

	and_bi _2250_ (
		.a(new_net_2239),
		.b(new_net_863),
		.c(_1287_)
	);

	and_bb _2251_ (
		.a(new_net_1475),
		.b(new_net_1441),
		.c(_1288_)
	);

	and_bi _2252_ (
		.a(new_net_2279),
		.b(new_net_2896),
		.c(_1289_)
	);

	and_bb _2253_ (
		.a(new_net_3079),
		.b(new_net_1254),
		.c(_1290_)
	);

	and_bi _2254_ (
		.a(new_net_1163),
		.b(new_net_1717),
		.c(_1291_)
	);

	and_bb _2255_ (
		.a(new_net_2345),
		.b(new_net_3178),
		.c(_1292_)
	);

	and_bi _2256_ (
		.a(new_net_1568),
		.b(new_net_1679),
		.c(_1293_)
	);

	and_bb _2257_ (
		.a(new_net_393),
		.b(new_net_2403),
		.c(_1294_)
	);

	and_bi _2258_ (
		.a(new_net_720),
		.b(new_net_1231),
		.c(_1295_)
	);

	and_bb _2259_ (
		.a(new_net_46),
		.b(new_net_376),
		.c(_1296_)
	);

	or_ii _2260_ (
		.a(new_net_1129),
		.b(new_net_3098),
		.c(_1297_)
	);

	and_bi _2261_ (
		.a(new_net_1175),
		.b(new_net_442),
		.c(_1298_)
	);

	and_bb _2262_ (
		.a(new_net_1117),
		.b(new_net_2921),
		.c(_1299_)
	);

	and_bi _2263_ (
		.a(new_net_2988),
		.b(new_net_962),
		.c(_1300_)
	);

	and_ii _2264_ (
		.a(new_net_3556),
		.b(new_net_630),
		.c(_1301_)
	);

	or_bb _2265_ (
		.a(new_net_1164),
		.b(new_net_3218),
		.c(_1302_)
	);

	or_ii _2266_ (
		.a(new_net_1165),
		.b(new_net_3219),
		.c(_1303_)
	);

	or_ii _2267_ (
		.a(new_net_3557),
		.b(new_net_1350),
		.c(_1304_)
	);

	and_ii _2268_ (
		.a(new_net_1718),
		.b(new_net_874),
		.c(_1305_)
	);

	and_bb _2269_ (
		.a(new_net_1719),
		.b(new_net_875),
		.c(_1306_)
	);

	or_bb _2270_ (
		.a(new_net_3558),
		.b(new_net_1898),
		.c(_1307_)
	);

	or_bb _2271_ (
		.a(new_net_2280),
		.b(new_net_854),
		.c(_1308_)
	);

	or_ii _2272_ (
		.a(new_net_2281),
		.b(new_net_855),
		.c(_1309_)
	);

	or_ii _2273_ (
		.a(new_net_3559),
		.b(new_net_1273),
		.c(_1310_)
	);

	and_ii _2274_ (
		.a(new_net_1346),
		.b(new_net_3129),
		.c(_1311_)
	);

	and_bb _2275_ (
		.a(new_net_1347),
		.b(new_net_3130),
		.c(_1312_)
	);

	or_bb _2276_ (
		.a(new_net_3560),
		.b(new_net_3133),
		.c(_1313_)
	);

	or_bb _2277_ (
		.a(new_net_244),
		.b(new_net_2888),
		.c(_1314_)
	);

	or_ii _2278_ (
		.a(new_net_245),
		.b(new_net_2889),
		.c(_1315_)
	);

	or_ii _2279_ (
		.a(new_net_3561),
		.b(new_net_1539),
		.c(_1316_)
	);

	and_ii _2280_ (
		.a(new_net_10),
		.b(new_net_699),
		.c(_1317_)
	);

	and_bb _2281_ (
		.a(new_net_11),
		.b(new_net_700),
		.c(_1318_)
	);

	or_bb _2282_ (
		.a(new_net_3562),
		.b(new_net_68),
		.c(_1319_)
	);

	or_bb _2283_ (
		.a(new_net_128),
		.b(new_net_2478),
		.c(_1320_)
	);

	or_ii _2284_ (
		.a(new_net_129),
		.b(new_net_2479),
		.c(_1321_)
	);

	or_ii _2285_ (
		.a(new_net_3563),
		.b(new_net_793),
		.c(_1322_)
	);

	and_ii _2286_ (
		.a(new_net_236),
		.b(new_net_2274),
		.c(_1323_)
	);

	and_bb _2287_ (
		.a(new_net_237),
		.b(new_net_2275),
		.c(_1324_)
	);

	or_bb _2288_ (
		.a(new_net_3564),
		.b(new_net_1298),
		.c(_1325_)
	);

	or_bb _2289_ (
		.a(new_net_337),
		.b(new_net_2092),
		.c(_1326_)
	);

	or_ii _2290_ (
		.a(new_net_338),
		.b(new_net_2093),
		.c(_1327_)
	);

	or_ii _2291_ (
		.a(new_net_3565),
		.b(new_net_1848),
		.c(_1328_)
	);

	and_ii _2292_ (
		.a(new_net_2246),
		.b(new_net_1892),
		.c(_1329_)
	);

	and_bb _2293_ (
		.a(new_net_2247),
		.b(new_net_1893),
		.c(_1330_)
	);

	or_bb _2294_ (
		.a(new_net_3566),
		.b(new_net_500),
		.c(_1331_)
	);

	or_bb _2295_ (
		.a(new_net_600),
		.b(new_net_504),
		.c(_1332_)
	);

	or_ii _2296_ (
		.a(new_net_601),
		.b(new_net_505),
		.c(_1333_)
	);

	or_ii _2297_ (
		.a(new_net_3567),
		.b(new_net_3063),
		.c(_1334_)
	);

	and_ii _2298_ (
		.a(new_net_697),
		.b(new_net_1580),
		.c(_1335_)
	);

	and_bb _2299_ (
		.a(new_net_698),
		.b(new_net_1581),
		.c(_1336_)
	);

	or_bb _2300_ (
		.a(new_net_3568),
		.b(new_net_765),
		.c(_1337_)
	);

	or_bb _2301_ (
		.a(new_net_801),
		.b(new_net_420),
		.c(_1338_)
	);

	or_ii _2302_ (
		.a(new_net_802),
		.b(new_net_421),
		.c(_1339_)
	);

	or_ii _2303_ (
		.a(new_net_3569),
		.b(new_net_870),
		.c(_1340_)
	);

	and_ii _2304_ (
		.a(new_net_1306),
		.b(new_net_366),
		.c(_1341_)
	);

	and_bb _2305_ (
		.a(new_net_1307),
		.b(new_net_367),
		.c(_1342_)
	);

	or_bb _2306_ (
		.a(new_net_3570),
		.b(new_net_1517),
		.c(_1343_)
	);

	or_bb _2307_ (
		.a(new_net_1856),
		.b(new_net_988),
		.c(_1344_)
	);

	or_ii _2308_ (
		.a(new_net_1857),
		.b(new_net_989),
		.c(_1345_)
	);

	or_ii _2309_ (
		.a(new_net_3571),
		.b(new_net_2030),
		.c(_1346_)
	);

	and_ii _2310_ (
		.a(new_net_2446),
		.b(new_net_842),
		.c(_1347_)
	);

	and_bb _2311_ (
		.a(new_net_2447),
		.b(new_net_843),
		.c(_1348_)
	);

	or_bb _2312_ (
		.a(new_net_3572),
		.b(new_net_2655),
		.c(_1349_)
	);

	or_bb _2313_ (
		.a(new_net_1214),
		.b(new_net_614),
		.c(_1350_)
	);

	or_ii _2314_ (
		.a(new_net_1215),
		.b(new_net_615),
		.c(_1351_)
	);

	or_ii _2315_ (
		.a(new_net_3573),
		.b(new_net_1281),
		.c(_1352_)
	);

	and_ii _2316_ (
		.a(new_net_354),
		.b(new_net_238),
		.c(_1353_)
	);

	and_bb _2317_ (
		.a(new_net_355),
		.b(new_net_239),
		.c(_1354_)
	);

	or_bb _2318_ (
		.a(new_net_3574),
		.b(new_net_1376),
		.c(_1355_)
	);

	or_bb _2319_ (
		.a(new_net_960),
		.b(new_net_226),
		.c(_1356_)
	);

	and_bb _2320_ (
		.a(new_net_961),
		.b(new_net_227),
		.c(_1357_)
	);

	or_bi _2321_ (
		.a(new_net_3575),
		.b(new_net_1535),
		.c(_1358_)
	);

	and_ii _2322_ (
		.a(new_net_1610),
		.b(new_net_172),
		.c(_1359_)
	);

	and_bb _2323_ (
		.a(new_net_1611),
		.b(new_net_173),
		.c(_1360_)
	);

	or_bb _2324_ (
		.a(new_net_3576),
		.b(new_net_2651),
		.c(new_net_3926)
	);

	and_bb _2325_ (
		.a(new_net_426),
		.b(new_net_2838),
		.c(_1361_)
	);

	and_bi _2326_ (
		.a(new_net_1536),
		.b(new_net_2652),
		.c(_1362_)
	);

	and_bb _2327_ (
		.a(new_net_2555),
		.b(new_net_3014),
		.c(_1363_)
	);

	and_bi _2328_ (
		.a(new_net_1282),
		.b(new_net_1377),
		.c(_1364_)
	);

	and_bb _2329_ (
		.a(new_net_2607),
		.b(new_net_3238),
		.c(_1365_)
	);

	and_bi _2330_ (
		.a(new_net_2031),
		.b(new_net_2656),
		.c(_1366_)
	);

	and_bb _2331_ (
		.a(new_net_744),
		.b(new_net_257),
		.c(_1367_)
	);

	and_bi _2332_ (
		.a(new_net_871),
		.b(new_net_1518),
		.c(_1368_)
	);

	and_bb _2333_ (
		.a(new_net_1408),
		.b(new_net_210),
		.c(_1369_)
	);

	and_bi _2334_ (
		.a(new_net_3064),
		.b(new_net_766),
		.c(_1370_)
	);

	and_bb _2335_ (
		.a(new_net_1476),
		.b(new_net_1798),
		.c(_1371_)
	);

	and_bi _2336_ (
		.a(new_net_1849),
		.b(new_net_501),
		.c(_1372_)
	);

	and_bb _2337_ (
		.a(new_net_3080),
		.b(new_net_1451),
		.c(_1373_)
	);

	and_bi _2338_ (
		.a(new_net_794),
		.b(new_net_1299),
		.c(_1374_)
	);

	and_bb _2339_ (
		.a(new_net_2346),
		.b(new_net_1247),
		.c(_1375_)
	);

	and_bi _2340_ (
		.a(new_net_1540),
		.b(new_net_69),
		.c(_1376_)
	);

	and_bb _2341_ (
		.a(new_net_3179),
		.b(new_net_2402),
		.c(_1377_)
	);

	and_bi _2342_ (
		.a(new_net_1274),
		.b(new_net_3134),
		.c(_1378_)
	);

	and_bb _2343_ (
		.a(new_net_398),
		.b(new_net_377),
		.c(_1379_)
	);

	and_bi _2344_ (
		.a(new_net_1351),
		.b(new_net_1899),
		.c(_1380_)
	);

	and_bb _2345_ (
		.a(new_net_2492),
		.b(new_net_47),
		.c(_1381_)
	);

	or_ii _2346_ (
		.a(new_net_1552),
		.b(new_net_3107),
		.c(_1382_)
	);

	and_bi _2347_ (
		.a(new_net_963),
		.b(new_net_582),
		.c(_1383_)
	);

	and_bb _2348_ (
		.a(new_net_1557),
		.b(new_net_2915),
		.c(_1384_)
	);

	and_bi _2349_ (
		.a(new_net_443),
		.b(new_net_958),
		.c(_1385_)
	);

	and_ii _2350_ (
		.a(new_net_3577),
		.b(new_net_807),
		.c(_1386_)
	);

	or_bb _2351_ (
		.a(new_net_2679),
		.b(new_net_632),
		.c(_1387_)
	);

	or_ii _2352_ (
		.a(new_net_2680),
		.b(new_net_631),
		.c(_1388_)
	);

	or_ii _2353_ (
		.a(new_net_3578),
		.b(new_net_1523),
		.c(_1389_)
	);

	and_ii _2354_ (
		.a(new_net_2775),
		.b(new_net_352),
		.c(_1390_)
	);

	and_bb _2355_ (
		.a(new_net_2776),
		.b(new_net_353),
		.c(_1391_)
	);

	or_bb _2356_ (
		.a(new_net_3579),
		.b(new_net_2038),
		.c(_1392_)
	);

	or_bb _2357_ (
		.a(new_net_2901),
		.b(new_net_188),
		.c(_1393_)
	);

	or_ii _2358_ (
		.a(new_net_2902),
		.b(new_net_189),
		.c(_1394_)
	);

	or_ii _2359_ (
		.a(new_net_3580),
		.b(new_net_2963),
		.c(_1395_)
	);

	and_ii _2360_ (
		.a(new_net_3075),
		.b(new_net_14),
		.c(_1396_)
	);

	and_bb _2361_ (
		.a(new_net_3076),
		.b(new_net_15),
		.c(_1397_)
	);

	or_bb _2362_ (
		.a(new_net_3581),
		.b(new_net_3109),
		.c(_1398_)
	);

	or_bb _2363_ (
		.a(new_net_360),
		.b(new_net_3067),
		.c(_1399_)
	);

	or_ii _2364_ (
		.a(new_net_361),
		.b(new_net_3068),
		.c(_1400_)
	);

	or_ii _2365_ (
		.a(new_net_3582),
		.b(new_net_3254),
		.c(_1401_)
	);

	and_ii _2366_ (
		.a(new_net_1644),
		.b(new_net_2825),
		.c(_1402_)
	);

	and_bb _2367_ (
		.a(new_net_1645),
		.b(new_net_2826),
		.c(_1403_)
	);

	or_bb _2368_ (
		.a(new_net_3583),
		.b(new_net_1692),
		.c(_1404_)
	);

	or_bb _2369_ (
		.a(new_net_1726),
		.b(new_net_2653),
		.c(_1405_)
	);

	or_ii _2370_ (
		.a(new_net_1727),
		.b(new_net_2654),
		.c(_1406_)
	);

	or_ii _2371_ (
		.a(new_net_3584),
		.b(new_net_832),
		.c(_1407_)
	);

	and_ii _2372_ (
		.a(new_net_1134),
		.b(new_net_2228),
		.c(_1408_)
	);

	and_bb _2373_ (
		.a(new_net_1135),
		.b(new_net_2229),
		.c(_1409_)
	);

	or_bb _2374_ (
		.a(new_net_3585),
		.b(new_net_1328),
		.c(_1410_)
	);

	or_bb _2375_ (
		.a(new_net_1944),
		.b(new_net_2248),
		.c(_1411_)
	);

	or_ii _2376_ (
		.a(new_net_1945),
		.b(new_net_2249),
		.c(_1412_)
	);

	or_ii _2377_ (
		.a(new_net_3586),
		.b(new_net_1982),
		.c(_1413_)
	);

	and_ii _2378_ (
		.a(new_net_2272),
		.b(new_net_2028),
		.c(_1414_)
	);

	and_bb _2379_ (
		.a(new_net_2273),
		.b(new_net_2029),
		.c(_1415_)
	);

	or_bb _2380_ (
		.a(new_net_3587),
		.b(new_net_2110),
		.c(_1416_)
	);

	or_bb _2381_ (
		.a(new_net_2878),
		.b(new_net_2118),
		.c(_1417_)
	);

	or_ii _2382_ (
		.a(new_net_2879),
		.b(new_net_2119),
		.c(_1418_)
	);

	or_ii _2383_ (
		.a(new_net_3588),
		.b(new_net_2236),
		.c(_1419_)
	);

	and_ii _2384_ (
		.a(new_net_222),
		.b(new_net_2076),
		.c(_1420_)
	);

	and_bb _2385_ (
		.a(new_net_223),
		.b(new_net_2077),
		.c(_1421_)
	);

	or_bb _2386_ (
		.a(new_net_3589),
		.b(new_net_2355),
		.c(_1422_)
	);

	or_bb _2387_ (
		.a(new_net_838),
		.b(new_net_1515),
		.c(_1423_)
	);

	or_ii _2388_ (
		.a(new_net_839),
		.b(new_net_1516),
		.c(_1424_)
	);

	or_ii _2389_ (
		.a(new_net_3590),
		.b(new_net_2464),
		.c(_1425_)
	);

	and_ii _2390_ (
		.a(new_net_2543),
		.b(new_net_1304),
		.c(_1426_)
	);

	and_bb _2391_ (
		.a(new_net_2544),
		.b(new_net_1305),
		.c(_1427_)
	);

	or_bb _2392_ (
		.a(new_net_3591),
		.b(new_net_2597),
		.c(_1428_)
	);

	or_bb _2393_ (
		.a(new_net_2677),
		.b(new_net_1946),
		.c(_1429_)
	);

	or_ii _2394_ (
		.a(new_net_2678),
		.b(new_net_1947),
		.c(_1430_)
	);

	or_ii _2395_ (
		.a(new_net_3592),
		.b(new_net_2084),
		.c(_1431_)
	);

	and_ii _2396_ (
		.a(new_net_2783),
		.b(new_net_1912),
		.c(_1432_)
	);

	and_bb _2397_ (
		.a(new_net_2784),
		.b(new_net_1913),
		.c(_1433_)
	);

	or_bb _2398_ (
		.a(new_net_3593),
		.b(new_net_2809),
		.c(_1434_)
	);

	or_bb _2399_ (
		.a(new_net_3125),
		.b(new_net_799),
		.c(_1435_)
	);

	or_ii _2400_ (
		.a(new_net_3126),
		.b(new_net_800),
		.c(_1436_)
	);

	or_ii _2401_ (
		.a(new_net_3594),
		.b(new_net_56),
		.c(_1437_)
	);

	and_ii _2402_ (
		.a(new_net_3049),
		.b(new_net_1836),
		.c(_1438_)
	);

	and_bb _2403_ (
		.a(new_net_3050),
		.b(new_net_1837),
		.c(_1439_)
	);

	or_bb _2404_ (
		.a(new_net_3595),
		.b(new_net_612),
		.c(_1440_)
	);

	or_bb _2405_ (
		.a(new_net_986),
		.b(new_net_1784),
		.c(_1441_)
	);

	or_ii _2406_ (
		.a(new_net_987),
		.b(new_net_1785),
		.c(_1442_)
	);

	or_ii _2407_ (
		.a(new_net_3596),
		.b(new_net_3258),
		.c(_1443_)
	);

	and_ii _2408_ (
		.a(new_net_3027),
		.b(new_net_1754),
		.c(_1444_)
	);

	and_bb _2409_ (
		.a(new_net_3028),
		.b(new_net_1755),
		.c(_1445_)
	);

	or_bb _2410_ (
		.a(new_net_3597),
		.b(new_net_104),
		.c(_1446_)
	);

	or_bb _2411_ (
		.a(new_net_178),
		.b(new_net_1730),
		.c(_1447_)
	);

	and_bb _2412_ (
		.a(new_net_179),
		.b(new_net_1731),
		.c(_1448_)
	);

	or_bi _2413_ (
		.a(new_net_3598),
		.b(new_net_542),
		.c(_1449_)
	);

	and_ii _2414_ (
		.a(new_net_277),
		.b(new_net_3059),
		.c(_1450_)
	);

	and_bb _2415_ (
		.a(new_net_278),
		.b(new_net_3060),
		.c(_1451_)
	);

	or_bb _2416_ (
		.a(new_net_3599),
		.b(new_net_1068),
		.c(new_net_3952)
	);

	and_bb _2417_ (
		.a(new_net_146),
		.b(new_net_2839),
		.c(_1452_)
	);

	and_bi _2418_ (
		.a(new_net_543),
		.b(new_net_1069),
		.c(_1453_)
	);

	and_bb _2419_ (
		.a(new_net_2556),
		.b(new_net_429),
		.c(_1454_)
	);

	and_bi _2420_ (
		.a(new_net_3259),
		.b(new_net_105),
		.c(_1455_)
	);

	and_bb _2421_ (
		.a(new_net_3012),
		.b(new_net_3239),
		.c(_1456_)
	);

	and_bi _2422_ (
		.a(new_net_57),
		.b(new_net_613),
		.c(_1457_)
	);

	and_bb _2423_ (
		.a(new_net_745),
		.b(new_net_2606),
		.c(_1459_)
	);

	and_bi _2424_ (
		.a(new_net_2085),
		.b(new_net_2810),
		.c(_1460_)
	);

	and_bb _2425_ (
		.a(new_net_1409),
		.b(new_net_266),
		.c(_1461_)
	);

	and_bi _2426_ (
		.a(new_net_2465),
		.b(new_net_2598),
		.c(_1462_)
	);

	and_bb _2427_ (
		.a(new_net_1477),
		.b(new_net_202),
		.c(_1463_)
	);

	and_bi _2428_ (
		.a(new_net_2237),
		.b(new_net_2356),
		.c(_1464_)
	);

	and_bb _2429_ (
		.a(new_net_3081),
		.b(new_net_1805),
		.c(_1465_)
	);

	and_bi _2430_ (
		.a(new_net_1983),
		.b(new_net_2111),
		.c(_1466_)
	);

	and_bb _2431_ (
		.a(new_net_2347),
		.b(new_net_1442),
		.c(_1467_)
	);

	and_bi _2432_ (
		.a(new_net_833),
		.b(new_net_1329),
		.c(_1468_)
	);

	and_bb _2433_ (
		.a(new_net_1248),
		.b(new_net_2404),
		.c(_1470_)
	);

	and_bi _2434_ (
		.a(new_net_3255),
		.b(new_net_1693),
		.c(_1471_)
	);

	and_bb _2435_ (
		.a(new_net_385),
		.b(new_net_3180),
		.c(_1472_)
	);

	and_bi _2436_ (
		.a(new_net_2964),
		.b(new_net_3110),
		.c(_1473_)
	);

	and_bb _2437_ (
		.a(new_net_2490),
		.b(new_net_399),
		.c(_1474_)
	);

	and_bi _2438_ (
		.a(new_net_1524),
		.b(new_net_2039),
		.c(_1475_)
	);

	and_bb _2439_ (
		.a(new_net_1122),
		.b(new_net_38),
		.c(_1476_)
	);

	or_ii _2440_ (
		.a(new_net_2712),
		.b(new_net_3099),
		.c(_1477_)
	);

	and_bi _2441_ (
		.a(new_net_959),
		.b(new_net_3037),
		.c(_1478_)
	);

	or_ii _2442_ (
		.a(new_net_2701),
		.b(new_net_2922),
		.c(_1479_)
	);

	and_bb _2443_ (
		.a(new_net_1372),
		.b(new_net_583),
		.c(_1481_)
	);

	and_ii _2444_ (
		.a(new_net_3600),
		.b(new_net_3),
		.c(_1482_)
	);

	or_bb _2445_ (
		.a(new_net_781),
		.b(new_net_808),
		.c(_1483_)
	);

	or_ii _2446_ (
		.a(new_net_782),
		.b(new_net_809),
		.c(_1484_)
	);

	or_ii _2447_ (
		.a(new_net_3601),
		.b(new_net_952),
		.c(_1485_)
	);

	and_ii _2448_ (
		.a(new_net_484),
		.b(new_net_1279),
		.c(_1486_)
	);

	and_bb _2449_ (
		.a(new_net_485),
		.b(new_net_1280),
		.c(_1487_)
	);

	or_bb _2450_ (
		.a(new_net_3602),
		.b(new_net_675),
		.c(_1488_)
	);

	or_bb _2451_ (
		.a(new_net_176),
		.b(new_net_2631),
		.c(_1489_)
	);

	or_ii _2452_ (
		.a(new_net_177),
		.b(new_net_2632),
		.c(_1490_)
	);

	or_ii _2453_ (
		.a(new_net_3603),
		.b(new_net_1198),
		.c(_1492_)
	);

	and_ii _2454_ (
		.a(new_net_305),
		.b(new_net_1182),
		.c(_1493_)
	);

	and_bb _2455_ (
		.a(new_net_306),
		.b(new_net_1183),
		.c(_1494_)
	);

	or_bb _2456_ (
		.a(new_net_3604),
		.b(new_net_1938),
		.c(_1495_)
	);

	or_bb _2457_ (
		.a(new_net_2372),
		.b(new_net_2218),
		.c(_1496_)
	);

	or_ii _2458_ (
		.a(new_net_2373),
		.b(new_net_2219),
		.c(_1497_)
	);

	or_ii _2459_ (
		.a(new_net_3605),
		.b(new_net_2567),
		.c(_1498_)
	);

	and_ii _2460_ (
		.a(new_net_560),
		.b(new_net_2000),
		.c(_1499_)
	);

	and_bb _2461_ (
		.a(new_net_561),
		.b(new_net_2001),
		.c(_1500_)
	);

	or_bb _2462_ (
		.a(new_net_3606),
		.b(new_net_3199),
		.c(_1501_)
	);

	or_bb _2463_ (
		.a(new_net_295),
		.b(new_net_1818),
		.c(_1503_)
	);

	or_ii _2464_ (
		.a(new_net_296),
		.b(new_net_1819),
		.c(_1504_)
	);

	or_ii _2465_ (
		.a(new_net_3607),
		.b(new_net_683),
		.c(_1505_)
	);

	and_ii _2466_ (
		.a(new_net_844),
		.b(new_net_1046),
		.c(_1506_)
	);

	and_bb _2467_ (
		.a(new_net_845),
		.b(new_net_1047),
		.c(_1507_)
	);

	or_bb _2468_ (
		.a(new_net_3608),
		.b(new_net_878),
		.c(_1508_)
	);

	or_bb _2469_ (
		.a(new_net_1624),
		.b(new_net_1285),
		.c(_1509_)
	);

	or_ii _2470_ (
		.a(new_net_1625),
		.b(new_net_1286),
		.c(_1510_)
	);

	or_ii _2471_ (
		.a(new_net_3609),
		.b(new_net_976),
		.c(_1511_)
	);

	and_ii _2472_ (
		.a(new_net_2170),
		.b(new_net_980),
		.c(_1512_)
	);

	and_bb _2473_ (
		.a(new_net_2171),
		.b(new_net_981),
		.c(_1514_)
	);

	or_bb _2474_ (
		.a(new_net_3610),
		.b(new_net_1058),
		.c(_1515_)
	);

	or_bb _2475_ (
		.a(new_net_2979),
		.b(new_net_940),
		.c(_1516_)
	);

	or_ii _2476_ (
		.a(new_net_2980),
		.b(new_net_941),
		.c(_1517_)
	);

	or_ii _2477_ (
		.a(new_net_3611),
		.b(new_net_3207),
		.c(_1518_)
	);

	and_ii _2478_ (
		.a(new_net_1277),
		.b(new_net_773),
		.c(_1519_)
	);

	and_bb _2479_ (
		.a(new_net_1278),
		.b(new_net_774),
		.c(_1520_)
	);

	or_bb _2480_ (
		.a(new_net_3612),
		.b(new_net_494),
		.c(_1521_)
	);

	or_bb _2481_ (
		.a(new_net_892),
		.b(new_net_566),
		.c(_1522_)
	);

	or_ii _2482_ (
		.a(new_net_893),
		.b(new_net_567),
		.c(_1523_)
	);

	or_ii _2483_ (
		.a(new_net_3613),
		.b(new_net_1040),
		.c(_1525_)
	);

	and_ii _2484_ (
		.a(new_net_1630),
		.b(new_net_339),
		.c(_1526_)
	);

	and_bb _2485_ (
		.a(new_net_1631),
		.b(new_net_340),
		.c(_1527_)
	);

	or_bb _2486_ (
		.a(new_net_3614),
		.b(new_net_1032),
		.c(_1528_)
	);

	or_bb _2487_ (
		.a(new_net_1388),
		.b(new_net_826),
		.c(_1529_)
	);

	or_ii _2488_ (
		.a(new_net_1389),
		.b(new_net_827),
		.c(_1530_)
	);

	or_ii _2489_ (
		.a(new_net_3615),
		.b(new_net_1700),
		.c(_1531_)
	);

	and_ii _2490_ (
		.a(new_net_1760),
		.b(new_net_769),
		.c(_1532_)
	);

	and_bb _2491_ (
		.a(new_net_1761),
		.b(new_net_770),
		.c(_1533_)
	);

	or_bb _2492_ (
		.a(new_net_3616),
		.b(new_net_2144),
		.c(_1534_)
	);

	or_bb _2493_ (
		.a(new_net_2531),
		.b(new_net_703),
		.c(_1536_)
	);

	or_ii _2494_ (
		.a(new_net_2532),
		.b(new_net_704),
		.c(_1537_)
	);

	or_ii _2495_ (
		.a(new_net_3617),
		.b(new_net_136),
		.c(_1538_)
	);

	and_ii _2496_ (
		.a(new_net_2008),
		.b(new_net_2795),
		.c(_1539_)
	);

	and_bb _2497_ (
		.a(new_net_2009),
		.b(new_net_2796),
		.c(_1540_)
	);

	or_bb _2498_ (
		.a(new_net_3618),
		.b(new_net_2068),
		.c(_1541_)
	);

	or_bb _2499_ (
		.a(new_net_677),
		.b(new_net_606),
		.c(_1542_)
	);

	or_ii _2500_ (
		.a(new_net_678),
		.b(new_net_607),
		.c(_1543_)
	);

	or_ii _2501_ (
		.a(new_net_3619),
		.b(new_net_2184),
		.c(_1544_)
	);

	and_ii _2502_ (
		.a(new_net_2264),
		.b(new_net_2210),
		.c(_1545_)
	);

	and_bb _2503_ (
		.a(new_net_2265),
		.b(new_net_2211),
		.c(_1546_)
	);

	or_bb _2504_ (
		.a(new_net_3620),
		.b(new_net_2307),
		.c(_1547_)
	);

	or_bb _2505_ (
		.a(new_net_2394),
		.b(new_net_1994),
		.c(_1548_)
	);

	or_ii _2506_ (
		.a(new_net_2395),
		.b(new_net_1995),
		.c(_1549_)
	);

	or_ii _2507_ (
		.a(new_net_3621),
		.b(new_net_1954),
		.c(_1550_)
	);

	and_ii _2508_ (
		.a(new_net_2509),
		.b(new_net_1812),
		.c(_1551_)
	);

	and_bb _2509_ (
		.a(new_net_2510),
		.b(new_net_1813),
		.c(_1552_)
	);

	or_bb _2510_ (
		.a(new_net_3622),
		.b(new_net_2569),
		.c(_1553_)
	);

	or_bb _2511_ (
		.a(new_net_2641),
		.b(new_net_1658),
		.c(_1554_)
	);

	and_bb _2512_ (
		.a(new_net_2642),
		.b(new_net_1659),
		.c(_1555_)
	);

	or_bi _2513_ (
		.a(new_net_3623),
		.b(new_net_3201),
		.c(_1557_)
	);

	and_ii _2514_ (
		.a(new_net_490),
		.b(new_net_1493),
		.c(_1558_)
	);

	and_bb _2515_ (
		.a(new_net_491),
		.b(new_net_1494),
		.c(_1559_)
	);

	or_bb _2516_ (
		.a(new_net_3624),
		.b(new_net_685),
		.c(new_net_3962)
	);

	and_bb _2517_ (
		.a(new_net_2831),
		.b(new_net_535),
		.c(_1560_)
	);

	and_bi _2518_ (
		.a(new_net_3202),
		.b(new_net_686),
		.c(_1561_)
	);

	and_bb _2519_ (
		.a(new_net_2557),
		.b(new_net_149),
		.c(_1562_)
	);

	and_bi _2520_ (
		.a(new_net_1955),
		.b(new_net_2570),
		.c(_1563_)
	);

	and_bb _2521_ (
		.a(new_net_427),
		.b(new_net_3240),
		.c(_1564_)
	);

	and_bi _2522_ (
		.a(new_net_2185),
		.b(new_net_2308),
		.c(_1565_)
	);

	and_bb _2523_ (
		.a(new_net_746),
		.b(new_net_3013),
		.c(_1567_)
	);

	and_bi _2524_ (
		.a(new_net_137),
		.b(new_net_2069),
		.c(_1568_)
	);

	and_bb _2525_ (
		.a(new_net_1410),
		.b(new_net_2615),
		.c(_1569_)
	);

	and_bi _2526_ (
		.a(new_net_1701),
		.b(new_net_2145),
		.c(_1570_)
	);

	and_bb _2527_ (
		.a(new_net_1478),
		.b(new_net_260),
		.c(_1571_)
	);

	and_bi _2528_ (
		.a(new_net_1041),
		.b(new_net_1033),
		.c(_1572_)
	);

	and_bb _2529_ (
		.a(new_net_3082),
		.b(new_net_211),
		.c(_1573_)
	);

	and_bi _2530_ (
		.a(new_net_3208),
		.b(new_net_495),
		.c(_1574_)
	);

	and_bb _2531_ (
		.a(new_net_2348),
		.b(new_net_1799),
		.c(_1575_)
	);

	and_bi _2532_ (
		.a(new_net_977),
		.b(new_net_1059),
		.c(_1576_)
	);

	and_bb _2533_ (
		.a(new_net_1443),
		.b(new_net_2405),
		.c(_1578_)
	);

	and_bi _2534_ (
		.a(new_net_684),
		.b(new_net_879),
		.c(_1579_)
	);

	and_bb _2535_ (
		.a(new_net_386),
		.b(new_net_1249),
		.c(_1580_)
	);

	and_bi _2536_ (
		.a(new_net_2568),
		.b(new_net_3200),
		.c(_1581_)
	);

	and_bb _2537_ (
		.a(new_net_2491),
		.b(new_net_3190),
		.c(_1582_)
	);

	and_bi _2538_ (
		.a(new_net_1199),
		.b(new_net_1939),
		.c(_1583_)
	);

	and_bb _2539_ (
		.a(new_net_1123),
		.b(new_net_394),
		.c(_1584_)
	);

	and_bi _2540_ (
		.a(new_net_953),
		.b(new_net_676),
		.c(_1585_)
	);

	and_bb _2541_ (
		.a(new_net_1547),
		.b(new_net_48),
		.c(_1586_)
	);

	or_ii _2542_ (
		.a(new_net_2046),
		.b(new_net_3108),
		.c(_1587_)
	);

	or_bb _2543_ (
		.a(new_net_2304),
		.b(new_net_1373),
		.c(_1589_)
	);

	and_bb _2544_ (
		.a(new_net_2054),
		.b(new_net_2916),
		.c(_1590_)
	);

	and_bi _2545_ (
		.a(new_net_3038),
		.b(new_net_1744),
		.c(_1591_)
	);

	and_bi _2546_ (
		.a(new_net_2386),
		.b(new_net_3625),
		.c(_1592_)
	);

	or_bb _2547_ (
		.a(new_net_2140),
		.b(new_net_4),
		.c(_1593_)
	);

	or_ii _2548_ (
		.a(new_net_2141),
		.b(new_net_5),
		.c(_1594_)
	);

	or_ii _2549_ (
		.a(new_net_3626),
		.b(new_net_2335),
		.c(_1595_)
	);

	and_ii _2550_ (
		.a(new_net_2744),
		.b(new_net_2262),
		.c(_1596_)
	);

	and_bb _2551_ (
		.a(new_net_2745),
		.b(new_net_2263),
		.c(_1597_)
	);

	or_bb _2552_ (
		.a(new_net_3627),
		.b(new_net_2953),
		.c(_1598_)
	);

	or_bb _2553_ (
		.a(new_net_114),
		.b(new_net_886),
		.c(_1600_)
	);

	or_ii _2554_ (
		.a(new_net_115),
		.b(new_net_887),
		.c(_1601_)
	);

	or_ii _2555_ (
		.a(new_net_3628),
		.b(new_net_482),
		.c(_1602_)
	);

	and_ii _2556_ (
		.a(new_net_2923),
		.b(new_net_671),
		.c(_1603_)
	);

	and_bb _2557_ (
		.a(new_net_2924),
		.b(new_net_672),
		.c(_1604_)
	);

	or_bb _2558_ (
		.a(new_net_3629),
		.b(new_net_2959),
		.c(_1605_)
	);

	or_bb _2559_ (
		.a(new_net_1392),
		.b(new_net_2162),
		.c(_1606_)
	);

	or_ii _2560_ (
		.a(new_net_1393),
		.b(new_net_2163),
		.c(_1607_)
	);

	or_ii _2561_ (
		.a(new_net_3630),
		.b(new_net_1608),
		.c(_1608_)
	);

	and_ii _2562_ (
		.a(new_net_1936),
		.b(new_net_2114),
		.c(_1609_)
	);

	and_bb _2563_ (
		.a(new_net_1937),
		.b(new_net_2115),
		.c(_1611_)
	);

	or_bb _2564_ (
		.a(new_net_3631),
		.b(new_net_2148),
		.c(_1612_)
	);

	or_bb _2565_ (
		.a(new_net_220),
		.b(new_net_2070),
		.c(_1613_)
	);

	or_ii _2566_ (
		.a(new_net_221),
		.b(new_net_2071),
		.c(_1614_)
	);

	or_ii _2567_ (
		.a(new_net_3632),
		.b(new_net_410),
		.c(_1615_)
	);

	and_ii _2568_ (
		.a(new_net_1750),
		.b(new_net_2018),
		.c(_1616_)
	);

	and_bb _2569_ (
		.a(new_net_1751),
		.b(new_net_2019),
		.c(_1617_)
	);

	or_bb _2570_ (
		.a(new_net_3633),
		.b(new_net_1788),
		.c(_1618_)
	);

	or_bb _2571_ (
		.a(new_net_1884),
		.b(new_net_2945),
		.c(_1619_)
	);

	or_ii _2572_ (
		.a(new_net_1885),
		.b(new_net_2946),
		.c(_1620_)
	);

	or_ii _2573_ (
		.a(new_net_3634),
		.b(new_net_1920),
		.c(_1622_)
	);

	and_ii _2574_ (
		.a(new_net_2078),
		.b(new_net_1948),
		.c(_1623_)
	);

	and_bb _2575_ (
		.a(new_net_2079),
		.b(new_net_1949),
		.c(_1624_)
	);

	or_bb _2576_ (
		.a(new_net_3635),
		.b(new_net_2072),
		.c(_1625_)
	);

	or_bb _2577_ (
		.a(new_net_2156),
		.b(new_net_2325),
		.c(_1626_)
	);

	or_ii _2578_ (
		.a(new_net_2157),
		.b(new_net_2326),
		.c(_1627_)
	);

	or_ii _2579_ (
		.a(new_net_3636),
		.b(new_net_2190),
		.c(_1628_)
	);

	and_ii _2580_ (
		.a(new_net_2258),
		.b(new_net_2132),
		.c(_1629_)
	);

	and_bb _2581_ (
		.a(new_net_2259),
		.b(new_net_2133),
		.c(_1630_)
	);

	or_bb _2582_ (
		.a(new_net_3637),
		.b(new_net_2298),
		.c(_1631_)
	);

	or_bb _2583_ (
		.a(new_net_610),
		.b(new_net_1928),
		.c(_1633_)
	);

	or_ii _2584_ (
		.a(new_net_611),
		.b(new_net_1929),
		.c(_1634_)
	);

	or_ii _2585_ (
		.a(new_net_3638),
		.b(new_net_2466),
		.c(_1635_)
	);

	and_ii _2586_ (
		.a(new_net_2533),
		.b(new_net_1740),
		.c(_1636_)
	);

	and_bb _2587_ (
		.a(new_net_2534),
		.b(new_net_1741),
		.c(_1637_)
	);

	or_bb _2588_ (
		.a(new_net_3639),
		.b(new_net_2595),
		.c(_1638_)
	);

	or_bb _2589_ (
		.a(new_net_2675),
		.b(new_net_1722),
		.c(_1639_)
	);

	or_ii _2590_ (
		.a(new_net_2676),
		.b(new_net_1723),
		.c(_1640_)
	);

	or_ii _2591_ (
		.a(new_net_3640),
		.b(new_net_2728),
		.c(_1641_)
	);

	and_ii _2592_ (
		.a(new_net_2474),
		.b(new_net_1708),
		.c(_1642_)
	);

	and_bb _2593_ (
		.a(new_net_2475),
		.b(new_net_1709),
		.c(_1644_)
	);

	or_bb _2594_ (
		.a(new_net_3641),
		.b(new_net_2811),
		.c(_1645_)
	);

	or_bb _2595_ (
		.a(new_net_54),
		.b(new_net_1188),
		.c(_1646_)
	);

	or_ii _2596_ (
		.a(new_net_55),
		.b(new_net_1189),
		.c(_1647_)
	);

	or_ii _2597_ (
		.a(new_net_3642),
		.b(new_net_2999),
		.c(_1648_)
	);

	and_ii _2598_ (
		.a(new_net_3121),
		.b(new_net_1648),
		.c(_1649_)
	);

	and_bb _2599_ (
		.a(new_net_3122),
		.b(new_net_1649),
		.c(_1650_)
	);

	or_bb _2600_ (
		.a(new_net_3643),
		.b(new_net_3139),
		.c(_1651_)
	);

	or_bb _2601_ (
		.a(new_net_1140),
		.b(new_net_1618),
		.c(_1652_)
	);

	or_ii _2602_ (
		.a(new_net_1141),
		.b(new_net_1619),
		.c(_1653_)
	);

	or_ii _2603_ (
		.a(new_net_3644),
		.b(new_net_24),
		.c(_1655_)
	);

	and_ii _2604_ (
		.a(new_net_578),
		.b(new_net_3250),
		.c(_1656_)
	);

	and_bb _2605_ (
		.a(new_net_579),
		.b(new_net_3251),
		.c(_1657_)
	);

	or_bb _2606_ (
		.a(new_net_3645),
		.b(new_net_791),
		.c(_1658_)
	);

	or_bb _2607_ (
		.a(new_net_1094),
		.b(new_net_3149),
		.c(_1659_)
	);

	or_ii _2608_ (
		.a(new_net_1095),
		.b(new_net_3150),
		.c(_1660_)
	);

	or_ii _2609_ (
		.a(new_net_3646),
		.b(new_net_1300),
		.c(_1661_)
	);

	and_ii _2610_ (
		.a(new_net_331),
		.b(new_net_3119),
		.c(_1662_)
	);

	and_bb _2611_ (
		.a(new_net_332),
		.b(new_net_3120),
		.c(_1663_)
	);

	or_bb _2612_ (
		.a(new_net_3647),
		.b(new_net_372),
		.c(_1664_)
	);

	or_bb _2613_ (
		.a(new_net_2242),
		.b(new_net_1626),
		.c(_1666_)
	);

	or_ii _2614_ (
		.a(new_net_2243),
		.b(new_net_1627),
		.c(_1667_)
	);

	or_ii _2615_ (
		.a(new_net_3648),
		.b(new_net_556),
		.c(_1668_)
	);

	and_ii _2616_ (
		.a(new_net_624),
		.b(new_net_3001),
		.c(_1669_)
	);

	and_bb _2617_ (
		.a(new_net_625),
		.b(new_net_3002),
		.c(_1670_)
	);

	or_bb _2618_ (
		.a(new_net_3649),
		.b(new_net_667),
		.c(_1671_)
	);

	or_bb _2619_ (
		.a(new_net_761),
		.b(new_net_2967),
		.c(_1672_)
	);

	and_bb _2620_ (
		.a(new_net_762),
		.b(new_net_2968),
		.c(_1673_)
	);

	or_bi _2621_ (
		.a(new_net_3650),
		.b(new_net_822),
		.c(_1674_)
	);

	and_ii _2622_ (
		.a(new_net_882),
		.b(new_net_2903),
		.c(_1675_)
	);

	and_bb _2623_ (
		.a(new_net_883),
		.b(new_net_2904),
		.c(_1677_)
	);

	or_bb _2624_ (
		.a(new_net_3651),
		.b(new_net_906),
		.c(new_net_3942)
	);

	and_bb _2625_ (
		.a(new_net_916),
		.b(new_net_2840),
		.c(_1678_)
	);

	and_bi _2626_ (
		.a(new_net_823),
		.b(new_net_907),
		.c(_1679_)
	);

	and_bb _2627_ (
		.a(new_net_2558),
		.b(new_net_528),
		.c(_1680_)
	);

	and_bi _2628_ (
		.a(new_net_557),
		.b(new_net_668),
		.c(_1681_)
	);

	and_bb _2629_ (
		.a(new_net_147),
		.b(new_net_3241),
		.c(_1682_)
	);

	and_bi _2630_ (
		.a(new_net_1301),
		.b(new_net_373),
		.c(_1683_)
	);

	and_bb _2631_ (
		.a(new_net_747),
		.b(new_net_428),
		.c(_1684_)
	);

	and_bi _2632_ (
		.a(new_net_25),
		.b(new_net_792),
		.c(_1685_)
	);

	and_bb _2633_ (
		.a(new_net_1411),
		.b(new_net_3018),
		.c(_1687_)
	);

	and_bi _2634_ (
		.a(new_net_3000),
		.b(new_net_3140),
		.c(_1688_)
	);

	and_bb _2635_ (
		.a(new_net_1479),
		.b(new_net_2609),
		.c(_1689_)
	);

	and_bi _2636_ (
		.a(new_net_2729),
		.b(new_net_2812),
		.c(_1690_)
	);

	and_bb _2637_ (
		.a(new_net_3083),
		.b(new_net_267),
		.c(_1691_)
	);

	and_bi _2638_ (
		.a(new_net_2467),
		.b(new_net_2596),
		.c(_1692_)
	);

	and_bb _2639_ (
		.a(new_net_2349),
		.b(new_net_203),
		.c(_1693_)
	);

	and_bi _2640_ (
		.a(new_net_2191),
		.b(new_net_2299),
		.c(_1694_)
	);

	and_bb _2641_ (
		.a(new_net_1800),
		.b(new_net_2406),
		.c(_1695_)
	);

	and_bi _2642_ (
		.a(new_net_1921),
		.b(new_net_2073),
		.c(_1696_)
	);

	and_bb _2643_ (
		.a(new_net_387),
		.b(new_net_1444),
		.c(_1698_)
	);

	and_bi _2644_ (
		.a(new_net_411),
		.b(new_net_1789),
		.c(_1699_)
	);

	and_bb _2645_ (
		.a(new_net_2493),
		.b(new_net_1255),
		.c(_1700_)
	);

	and_bi _2646_ (
		.a(new_net_1609),
		.b(new_net_2149),
		.c(_1701_)
	);

	and_bb _2647_ (
		.a(new_net_1124),
		.b(new_net_3181),
		.c(_1702_)
	);

	and_bi _2648_ (
		.a(new_net_483),
		.b(new_net_2960),
		.c(_1703_)
	);

	and_bb _2649_ (
		.a(new_net_1545),
		.b(new_net_400),
		.c(_1704_)
	);

	and_bi _2650_ (
		.a(new_net_2336),
		.b(new_net_2954),
		.c(_1705_)
	);

	and_bb _2651_ (
		.a(new_net_2706),
		.b(new_net_39),
		.c(_1706_)
	);

	and_ii _2652_ (
		.a(new_net_2387),
		.b(new_net_2870),
		.c(_1707_)
	);

	and_bb _2653_ (
		.a(new_net_2861),
		.b(new_net_2920),
		.c(_1709_)
	);

	and_bi _2654_ (
		.a(new_net_2306),
		.b(new_net_2374),
		.c(_1710_)
	);

	or_bb _2655_ (
		.a(new_net_2305),
		.b(new_net_2697),
		.c(_1711_)
	);

	and_bi _2656_ (
		.a(new_net_2375),
		.b(_1711_),
		.c(_1712_)
	);

	or_bb _2657_ (
		.a(_1712_),
		.b(new_net_3652),
		.c(_1713_)
	);

	or_bb _2658_ (
		.a(new_net_3203),
		.b(_1707_),
		.c(_1714_)
	);

	and_ii _2659_ (
		.a(new_net_2361),
		.b(new_net_2022),
		.c(_1715_)
	);

	and_bb _2660_ (
		.a(new_net_2362),
		.b(new_net_2023),
		.c(_1716_)
	);

	or_bb _2661_ (
		.a(new_net_3653),
		.b(new_net_297),
		.c(_1717_)
	);

	or_bb _2662_ (
		.a(new_net_687),
		.b(new_net_1984),
		.c(_1718_)
	);

	or_ii _2663_ (
		.a(new_net_688),
		.b(new_net_1985),
		.c(_1720_)
	);

	or_ii _2664_ (
		.a(new_net_3654),
		.b(new_net_2482),
		.c(_1721_)
	);

	and_ii _2665_ (
		.a(new_net_1396),
		.b(new_net_1394),
		.c(_1722_)
	);

	and_bb _2666_ (
		.a(new_net_1397),
		.b(new_net_1395),
		.c(_1723_)
	);

	or_bb _2667_ (
		.a(new_net_3655),
		.b(new_net_1628),
		.c(_1724_)
	);

	or_bb _2668_ (
		.a(new_net_1958),
		.b(new_net_1200),
		.c(_1725_)
	);

	or_ii _2669_ (
		.a(new_net_1959),
		.b(new_net_1201),
		.c(_1726_)
	);

	or_ii _2670_ (
		.a(new_net_3656),
		.b(new_net_2172),
		.c(_1727_)
	);

	and_ii _2671_ (
		.a(new_net_2853),
		.b(new_net_1880),
		.c(_1728_)
	);

	and_bb _2672_ (
		.a(new_net_2854),
		.b(new_net_1881),
		.c(_1729_)
	);

	or_bb _2673_ (
		.a(new_net_3657),
		.b(new_net_2763),
		.c(_1731_)
	);

	or_bb _2674_ (
		.a(new_net_3043),
		.b(new_net_1832),
		.c(_1732_)
	);

	or_ii _2675_ (
		.a(new_net_3044),
		.b(new_net_1833),
		.c(_1733_)
	);

	or_ii _2676_ (
		.a(new_net_3658),
		.b(new_net_3113),
		.c(_1734_)
	);

	and_ii _2677_ (
		.a(new_net_3195),
		.b(new_net_679),
		.c(_1735_)
	);

	and_bb _2678_ (
		.a(new_net_3196),
		.b(new_net_680),
		.c(_1736_)
	);

	or_bb _2679_ (
		.a(new_net_3659),
		.b(new_net_3252),
		.c(_1737_)
	);

	or_bb _2680_ (
		.a(new_net_1890),
		.b(new_net_1764),
		.c(_1738_)
	);

	or_ii _2681_ (
		.a(new_net_1891),
		.b(new_net_1765),
		.c(_1739_)
	);

	or_ii _2682_ (
		.a(new_net_3660),
		.b(new_net_2088),
		.c(_1740_)
	);

	and_ii _2683_ (
		.a(new_net_1724),
		.b(new_net_291),
		.c(_1742_)
	);

	and_bb _2684_ (
		.a(new_net_1725),
		.b(new_net_292),
		.c(_1743_)
	);

	or_bb _2685_ (
		.a(new_net_3661),
		.b(new_net_2884),
		.c(_1744_)
	);

	or_bb _2686_ (
		.a(new_net_1866),
		.b(new_net_3197),
		.c(_1745_)
	);

	or_ii _2687_ (
		.a(new_net_1867),
		.b(new_net_3198),
		.c(_1746_)
	);

	or_ii _2688_ (
		.a(new_net_3662),
		.b(new_net_1914),
		.c(_1747_)
	);

	and_ii _2689_ (
		.a(new_net_628),
		.b(new_net_2975),
		.c(_1748_)
	);

	and_bb _2690_ (
		.a(new_net_629),
		.b(new_net_2976),
		.c(_1749_)
	);

	or_bb _2691_ (
		.a(new_net_3663),
		.b(new_net_860),
		.c(_1750_)
	);

	or_bb _2692_ (
		.a(new_net_2120),
		.b(new_net_1620),
		.c(_1751_)
	);

	or_ii _2693_ (
		.a(new_net_2121),
		.b(new_net_1621),
		.c(_1753_)
	);

	or_ii _2694_ (
		.a(new_net_3664),
		.b(new_net_2164),
		.c(_1754_)
	);

	and_ii _2695_ (
		.a(new_net_1896),
		.b(new_net_1573),
		.c(_1755_)
	);

	and_bb _2696_ (
		.a(new_net_1897),
		.b(new_net_1574),
		.c(_1756_)
	);

	or_bb _2697_ (
		.a(new_net_3665),
		.b(new_net_2098),
		.c(_1757_)
	);

	or_bb _2698_ (
		.a(new_net_2388),
		.b(new_net_1533),
		.c(_1758_)
	);

	or_ii _2699_ (
		.a(new_net_2389),
		.b(new_net_1534),
		.c(_1759_)
	);

	or_ii _2700_ (
		.a(new_net_3666),
		.b(new_net_2691),
		.c(_1760_)
	);

	and_ii _2701_ (
		.a(new_net_3131),
		.b(new_net_1465),
		.c(_1761_)
	);

	and_bb _2702_ (
		.a(new_net_3132),
		.b(new_net_1466),
		.c(_1762_)
	);

	or_bb _2703_ (
		.a(new_net_3667),
		.b(new_net_2545),
		.c(_1764_)
	);

	or_bb _2704_ (
		.a(new_net_635),
		.b(new_net_812),
		.c(_1765_)
	);

	or_ii _2705_ (
		.a(new_net_636),
		.b(new_net_813),
		.c(_1766_)
	);

	or_ii _2706_ (
		.a(new_net_3668),
		.b(new_net_2695),
		.c(_1767_)
	);

	and_ii _2707_ (
		.a(new_net_1166),
		.b(new_net_584),
		.c(_1768_)
	);

	and_bb _2708_ (
		.a(new_net_1167),
		.b(new_net_585),
		.c(_1769_)
	);

	or_bb _2709_ (
		.a(new_net_3669),
		.b(new_net_1354),
		.c(_1770_)
	);

	or_bb _2710_ (
		.a(new_net_1720),
		.b(new_net_1344),
		.c(_1771_)
	);

	or_ii _2711_ (
		.a(new_net_1721),
		.b(new_net_1345),
		.c(_1772_)
	);

	or_ii _2712_ (
		.a(new_net_3670),
		.b(new_net_1904),
		.c(_1773_)
	);

	and_ii _2713_ (
		.a(new_net_2286),
		.b(new_net_190),
		.c(_1775_)
	);

	and_bb _2714_ (
		.a(new_net_2287),
		.b(new_net_191),
		.c(_1776_)
	);

	or_bb _2715_ (
		.a(new_net_3671),
		.b(new_net_3145),
		.c(_1777_)
	);

	or_bb _2716_ (
		.a(new_net_3137),
		.b(new_net_1218),
		.c(_1778_)
	);

	or_ii _2717_ (
		.a(new_net_3138),
		.b(new_net_1219),
		.c(_1779_)
	);

	or_ii _2718_ (
		.a(new_net_3672),
		.b(new_net_28),
		.c(_1780_)
	);

	and_ii _2719_ (
		.a(new_net_828),
		.b(new_net_2827),
		.c(_1781_)
	);

	and_bb _2720_ (
		.a(new_net_829),
		.b(new_net_2828),
		.c(_1782_)
	);

	or_bb _2721_ (
		.a(new_net_3673),
		.b(new_net_124),
		.c(_1783_)
	);

	or_bb _2722_ (
		.a(new_net_1322),
		.b(new_net_1148),
		.c(_1784_)
	);

	or_ii _2723_ (
		.a(new_net_1323),
		.b(new_net_1149),
		.c(_1786_)
	);

	or_ii _2724_ (
		.a(new_net_3674),
		.b(new_net_1543),
		.c(_1787_)
	);

	and_ii _2725_ (
		.a(new_net_2040),
		.b(new_net_1106),
		.c(_1788_)
	);

	and_bb _2726_ (
		.a(new_net_2041),
		.b(new_net_1107),
		.c(_1789_)
	);

	or_bb _2727_ (
		.a(new_net_3675),
		.b(new_net_368),
		.c(_1790_)
	);

	or_bb _2728_ (
		.a(new_net_2661),
		.b(new_net_2250),
		.c(_1791_)
	);

	or_ii _2729_ (
		.a(new_net_2662),
		.b(new_net_2251),
		.c(_1792_)
	);

	or_ii _2730_ (
		.a(new_net_3676),
		.b(new_net_2845),
		.c(_1793_)
	);

	and_ii _2731_ (
		.a(new_net_592),
		.b(new_net_1056),
		.c(_1794_)
	);

	and_bb _2732_ (
		.a(new_net_593),
		.b(new_net_1057),
		.c(_1795_)
	);

	or_bb _2733_ (
		.a(new_net_3677),
		.b(new_net_618),
		.c(_1797_)
	);

	and_ii _2734_ (
		.a(new_net_830),
		.b(new_net_1852),
		.c(_1798_)
	);

	and_bb _2735_ (
		.a(new_net_831),
		.b(new_net_1853),
		.c(_1799_)
	);

	or_bb _2736_ (
		.a(new_net_3678),
		.b(new_net_820),
		.c(_1800_)
	);

	and_ii _2737_ (
		.a(new_net_1324),
		.b(new_net_992),
		.c(_1801_)
	);

	and_bb _2738_ (
		.a(new_net_1325),
		.b(new_net_993),
		.c(_1802_)
	);

	or_bb _2739_ (
		.a(new_net_3679),
		.b(new_net_1561),
		.c(new_net_3920)
	);

	and_bi _2740_ (
		.a(new_net_2846),
		.b(new_net_619),
		.c(_1803_)
	);

	and_bb _2741_ (
		.a(new_net_527),
		.b(new_net_3242),
		.c(_1804_)
	);

	and_bi _2742_ (
		.a(new_net_1544),
		.b(new_net_369),
		.c(_1805_)
	);

	and_bb _2743_ (
		.a(new_net_748),
		.b(new_net_148),
		.c(_1807_)
	);

	and_bi _2744_ (
		.a(new_net_29),
		.b(new_net_125),
		.c(_1808_)
	);

	and_bb _2745_ (
		.a(new_net_1412),
		.b(new_net_436),
		.c(_1809_)
	);

	and_bi _2746_ (
		.a(new_net_1905),
		.b(new_net_3146),
		.c(_1810_)
	);

	and_bb _2747_ (
		.a(new_net_1480),
		.b(new_net_3015),
		.c(_1811_)
	);

	and_bi _2748_ (
		.a(new_net_2696),
		.b(new_net_1355),
		.c(_1812_)
	);

	and_bb _2749_ (
		.a(new_net_3084),
		.b(new_net_2616),
		.c(_1813_)
	);

	and_bi _2750_ (
		.a(new_net_2692),
		.b(new_net_2546),
		.c(_1814_)
	);

	and_bb _2751_ (
		.a(new_net_2350),
		.b(new_net_261),
		.c(_1815_)
	);

	and_bi _2752_ (
		.a(new_net_2165),
		.b(new_net_2099),
		.c(_1816_)
	);

	and_bb _2753_ (
		.a(new_net_204),
		.b(new_net_2407),
		.c(_1817_)
	);

	and_bi _2754_ (
		.a(new_net_1915),
		.b(new_net_861),
		.c(_1818_)
	);

	and_bb _2755_ (
		.a(new_net_1806),
		.b(new_net_379),
		.c(_1819_)
	);

	and_bi _2756_ (
		.a(new_net_2089),
		.b(new_net_2885),
		.c(_1820_)
	);

	and_bb _2757_ (
		.a(new_net_2494),
		.b(new_net_1452),
		.c(_1821_)
	);

	and_bi _2758_ (
		.a(new_net_3114),
		.b(new_net_3253),
		.c(_1822_)
	);

	and_bb _2759_ (
		.a(new_net_1125),
		.b(new_net_1250),
		.c(_1823_)
	);

	and_bi _2760_ (
		.a(new_net_2173),
		.b(new_net_2764),
		.c(_1824_)
	);

	and_bb _2761_ (
		.a(new_net_1546),
		.b(new_net_3191),
		.c(_1825_)
	);

	and_bi _2762_ (
		.a(new_net_2483),
		.b(new_net_1629),
		.c(_1826_)
	);

	and_bb _2763_ (
		.a(new_net_2707),
		.b(new_net_395),
		.c(_1828_)
	);

	and_ii _2764_ (
		.a(new_net_298),
		.b(new_net_3204),
		.c(_1829_)
	);

	or_ii _2765_ (
		.a(new_net_2863),
		.b(new_net_3104),
		.c(_1830_)
	);

	or_bb _2766_ (
		.a(new_net_1320),
		.b(new_net_1745),
		.c(_1831_)
	);

	and_bb _2767_ (
		.a(new_net_2051),
		.b(new_net_40),
		.c(_1832_)
	);

	and_ii _2768_ (
		.a(new_net_2020),
		.b(new_net_1541),
		.c(_1833_)
	);

	and_bb _2769_ (
		.a(new_net_2021),
		.b(new_net_1542),
		.c(_1834_)
	);

	or_bb _2770_ (
		.a(new_net_3680),
		.b(new_net_1860),
		.c(_1835_)
	);

	or_bb _2771_ (
		.a(new_net_2252),
		.b(new_net_1918),
		.c(_1836_)
	);

	or_ii _2772_ (
		.a(new_net_2253),
		.b(new_net_1919),
		.c(_1837_)
	);

	or_ii _2773_ (
		.a(new_net_3681),
		.b(new_net_2450),
		.c(_0001_)
	);

	and_ii _2774_ (
		.a(new_net_956),
		.b(new_net_1868),
		.c(_0002_)
	);

	and_bb _2775_ (
		.a(new_net_957),
		.b(new_net_1869),
		.c(_0003_)
	);

	or_bb _2776_ (
		.a(new_net_3682),
		.b(new_net_1006),
		.c(_0004_)
	);

	or_bb _2777_ (
		.a(new_net_1132),
		.b(new_net_588),
		.c(_0005_)
	);

	or_ii _2778_ (
		.a(new_net_1133),
		.b(new_net_589),
		.c(_0006_)
	);

	or_ii _2779_ (
		.a(new_net_3683),
		.b(new_net_1196),
		.c(_0007_)
	);

	and_ii _2780_ (
		.a(new_net_1314),
		.b(new_net_1762),
		.c(_0008_)
	);

	and_bb _2781_ (
		.a(new_net_1315),
		.b(new_net_1763),
		.c(_0009_)
	);

	or_bb _2782_ (
		.a(new_net_3684),
		.b(new_net_1336),
		.c(_0010_)
	);

	or_bb _2783_ (
		.a(new_net_1427),
		.b(new_net_192),
		.c(_0012_)
	);

	or_ii _2784_ (
		.a(new_net_1428),
		.b(new_net_193),
		.c(_0013_)
	);

	or_ii _2785_ (
		.a(new_net_3685),
		.b(new_net_1531),
		.c(_0014_)
	);

	and_ii _2786_ (
		.a(new_net_22),
		.b(new_net_18),
		.c(_0015_)
	);

	and_bb _2787_ (
		.a(new_net_23),
		.b(new_net_19),
		.c(_0016_)
	);

	or_bb _2788_ (
		.a(new_net_3686),
		.b(new_net_58),
		.c(_0017_)
	);

	or_bb _2789_ (
		.a(new_net_130),
		.b(new_net_3071),
		.c(_0018_)
	);

	or_ii _2790_ (
		.a(new_net_131),
		.b(new_net_3072),
		.c(_0019_)
	);

	or_ii _2791_ (
		.a(new_net_3687),
		.b(new_net_2319),
		.c(_0020_)
	);

	and_ii _2792_ (
		.a(new_net_234),
		.b(new_net_1646),
		.c(_0021_)
	);

	and_bb _2793_ (
		.a(new_net_235),
		.b(new_net_1647),
		.c(_0023_)
	);

	or_bb _2794_ (
		.a(new_net_3688),
		.b(new_net_2939),
		.c(_0024_)
	);

	or_bb _2795_ (
		.a(new_net_285),
		.b(new_net_1622),
		.c(_0025_)
	);

	or_ii _2796_ (
		.a(new_net_286),
		.b(new_net_1623),
		.c(_0026_)
	);

	or_ii _2797_ (
		.a(new_net_3689),
		.b(new_net_474),
		.c(_0027_)
	);

	and_ii _2798_ (
		.a(new_net_884),
		.b(new_net_1698),
		.c(_0028_)
	);

	and_bb _2799_ (
		.a(new_net_885),
		.b(new_net_1699),
		.c(_0029_)
	);

	or_bb _2800_ (
		.a(new_net_3690),
		.b(new_net_550),
		.c(_0030_)
	);

	or_bb _2801_ (
		.a(new_net_622),
		.b(new_net_1563),
		.c(_0031_)
	);

	or_ii _2802_ (
		.a(new_net_623),
		.b(new_net_1564),
		.c(_0032_)
	);

	or_ii _2803_ (
		.a(new_net_3691),
		.b(new_net_1604),
		.c(_0034_)
	);

	and_ii _2804_ (
		.a(new_net_818),
		.b(new_net_1326),
		.c(_0035_)
	);

	and_bb _2805_ (
		.a(new_net_819),
		.b(new_net_1327),
		.c(_0036_)
	);

	or_bb _2806_ (
		.a(new_net_3692),
		.b(new_net_2329),
		.c(_0037_)
	);

	or_bb _2807_ (
		.a(new_net_2738),
		.b(new_net_1429),
		.c(_0038_)
	);

	or_ii _2808_ (
		.a(new_net_2739),
		.b(new_net_1430),
		.c(_0039_)
	);

	or_ii _2809_ (
		.a(new_net_3693),
		.b(new_net_2947),
		.c(_0040_)
	);

	and_ii _2810_ (
		.a(new_net_108),
		.b(new_net_982),
		.c(_0041_)
	);

	and_bb _2811_ (
		.a(new_net_109),
		.b(new_net_983),
		.c(_0042_)
	);

	or_bb _2812_ (
		.a(new_net_3694),
		.b(new_net_1022),
		.c(_0043_)
	);

	or_bb _2813_ (
		.a(new_net_673),
		.b(new_net_1332),
		.c(_0045_)
	);

	or_ii _2814_ (
		.a(new_net_674),
		.b(new_net_1333),
		.c(_0046_)
	);

	or_ii _2815_ (
		.a(new_net_3695),
		.b(new_net_1030),
		.c(_0047_)
	);

	and_ii _2816_ (
		.a(new_net_1386),
		.b(new_net_608),
		.c(_0048_)
	);

	and_bb _2817_ (
		.a(new_net_1387),
		.b(new_net_609),
		.c(_0049_)
	);

	or_bb _2818_ (
		.a(new_net_3696),
		.b(new_net_1606),
		.c(_0050_)
	);

	or_bb _2819_ (
		.a(new_net_1932),
		.b(new_net_408),
		.c(_0051_)
	);

	or_ii _2820_ (
		.a(new_net_1933),
		.b(new_net_409),
		.c(_0052_)
	);

	or_ii _2821_ (
		.a(new_net_3697),
		.b(new_net_1378),
		.c(_0053_)
	);

	and_ii _2822_ (
		.a(new_net_2527),
		.b(new_net_218),
		.c(_0054_)
	);

	and_bb _2823_ (
		.a(new_net_2528),
		.b(new_net_219),
		.c(_0056_)
	);

	or_bb _2824_ (
		.a(new_net_3698),
		.b(new_net_2748),
		.c(_0057_)
	);

	or_bb _2825_ (
		.a(new_net_3209),
		.b(new_net_1172),
		.c(_0058_)
	);

	or_ii _2826_ (
		.a(new_net_3210),
		.b(new_net_1173),
		.c(_0059_)
	);

	or_ii _2827_ (
		.a(new_net_3699),
		.b(new_net_1688),
		.c(_0060_)
	);

	and_ii _2828_ (
		.a(new_net_1732),
		.b(new_net_1154),
		.c(_0061_)
	);

	and_bb _2829_ (
		.a(new_net_1733),
		.b(new_net_1155),
		.c(_0062_)
	);

	or_bb _2830_ (
		.a(new_net_3700),
		.b(new_net_691),
		.c(_0063_)
	);

	or_bb _2831_ (
		.a(new_net_1042),
		.b(new_net_2847),
		.c(_0064_)
	);

	or_ii _2832_ (
		.a(new_net_1043),
		.b(new_net_2848),
		.c(_0065_)
	);

	or_ii _2833_ (
		.a(new_net_3701),
		.b(new_net_1204),
		.c(_0067_)
	);

	and_ii _2834_ (
		.a(new_net_1978),
		.b(new_net_2663),
		.c(_0068_)
	);

	and_bb _2835_ (
		.a(new_net_1979),
		.b(new_net_2664),
		.c(_0069_)
	);

	or_bb _2836_ (
		.a(new_net_3702),
		.b(new_net_1960),
		.c(_0070_)
	);

	or_bb _2837_ (
		.a(new_net_2108),
		.b(new_net_2256),
		.c(_0071_)
	);

	or_ii _2838_ (
		.a(new_net_2109),
		.b(new_net_2257),
		.c(_0072_)
	);

	or_ii _2839_ (
		.a(new_net_3703),
		.b(new_net_2575),
		.c(_0073_)
	);

	and_ii _2840_ (
		.a(new_net_2983),
		.b(new_net_2058),
		.c(_0074_)
	);

	and_bb _2841_ (
		.a(new_net_2984),
		.b(new_net_2059),
		.c(_0075_)
	);

	or_bb _2842_ (
		.a(new_net_3704),
		.b(new_net_2268),
		.c(_0076_)
	);

	or_bb _2843_ (
		.a(new_net_2290),
		.b(new_net_1864),
		.c(_0078_)
	);

	and_bb _2844_ (
		.a(new_net_2562),
		.b(new_net_922),
		.c(_0079_)
	);

	or_ii _2845_ (
		.a(new_net_2291),
		.b(new_net_1865),
		.c(_0080_)
	);

	or_ii _2846_ (
		.a(new_net_3705),
		.b(new_net_2438),
		.c(_0081_)
	);

	and_ii _2847_ (
		.a(new_net_1228),
		.b(new_net_2460),
		.c(_0082_)
	);

	and_bi _2848_ (
		.a(new_net_2439),
		.b(new_net_1435),
		.c(_0083_)
	);

	and_bb _2849_ (
		.a(new_net_918),
		.b(new_net_3243),
		.c(_0084_)
	);

	and_bi _2850_ (
		.a(new_net_2576),
		.b(new_net_2269),
		.c(_0085_)
	);

	and_bb _2851_ (
		.a(new_net_749),
		.b(new_net_526),
		.c(_0086_)
	);

	and_bi _2852_ (
		.a(new_net_1205),
		.b(new_net_1961),
		.c(_0087_)
	);

	and_bb _2853_ (
		.a(new_net_1413),
		.b(new_net_157),
		.c(_0089_)
	);

	and_bi _2854_ (
		.a(new_net_1689),
		.b(new_net_692),
		.c(_0090_)
	);

	and_bb _2855_ (
		.a(new_net_1481),
		.b(new_net_430),
		.c(_0091_)
	);

	and_bi _2856_ (
		.a(new_net_1379),
		.b(new_net_2749),
		.c(_0092_)
	);

	and_bb _2857_ (
		.a(new_net_3085),
		.b(new_net_3019),
		.c(_0093_)
	);

	and_bi _2858_ (
		.a(new_net_1031),
		.b(new_net_1607),
		.c(_0094_)
	);

	and_bb _2859_ (
		.a(new_net_2351),
		.b(new_net_2610),
		.c(_0095_)
	);

	and_bi _2860_ (
		.a(new_net_2948),
		.b(new_net_1023),
		.c(_0096_)
	);

	and_bb _2861_ (
		.a(new_net_262),
		.b(new_net_2408),
		.c(_0097_)
	);

	and_bi _2862_ (
		.a(new_net_1605),
		.b(new_net_2330),
		.c(_0098_)
	);

	and_bb _2863_ (
		.a(new_net_212),
		.b(new_net_380),
		.c(_0100_)
	);

	and_bi _2864_ (
		.a(new_net_475),
		.b(new_net_551),
		.c(_0101_)
	);

	and_bb _2865_ (
		.a(new_net_2495),
		.b(new_net_1807),
		.c(_0102_)
	);

	and_bi _2866_ (
		.a(new_net_2320),
		.b(new_net_2940),
		.c(_0103_)
	);

	and_bb _2867_ (
		.a(new_net_1126),
		.b(new_net_1445),
		.c(_0104_)
	);

	and_bi _2868_ (
		.a(new_net_1532),
		.b(new_net_59),
		.c(_0105_)
	);

	and_bb _2869_ (
		.a(new_net_1548),
		.b(new_net_1256),
		.c(_0106_)
	);

	and_bi _2870_ (
		.a(new_net_1197),
		.b(new_net_1337),
		.c(_0107_)
	);

	and_bb _2871_ (
		.a(new_net_2708),
		.b(new_net_3182),
		.c(_0108_)
	);

	and_bi _2872_ (
		.a(new_net_2451),
		.b(new_net_1007),
		.c(_0109_)
	);

	and_bb _2873_ (
		.a(new_net_2042),
		.b(new_net_401),
		.c(_0111_)
	);

	and_bb _2874_ (
		.a(new_net_2871),
		.b(new_net_51),
		.c(_0112_)
	);

	and_ii _2875_ (
		.a(new_net_1861),
		.b(new_net_1321),
		.c(_0113_)
	);

	and_ii _2876_ (
		.a(new_net_2150),
		.b(new_net_3029),
		.c(_0114_)
	);

	and_bb _2877_ (
		.a(new_net_2151),
		.b(new_net_3030),
		.c(_0115_)
	);

	or_bb _2878_ (
		.a(new_net_3706),
		.b(new_net_2186),
		.c(_0116_)
	);

	and_ii _2879_ (
		.a(new_net_544),
		.b(new_net_2791),
		.c(_0117_)
	);

	and_bb _2880_ (
		.a(new_net_545),
		.b(new_net_2792),
		.c(_0118_)
	);

	or_bb _2881_ (
		.a(new_net_3707),
		.b(new_net_753),
		.c(_0119_)
	);

	or_bb _2882_ (
		.a(new_net_2390),
		.b(new_net_1974),
		.c(_0120_)
	);

	or_ii _2883_ (
		.a(new_net_2391),
		.b(new_net_1975),
		.c(_0122_)
	);

	or_ii _2884_ (
		.a(new_net_3708),
		.b(new_net_2432),
		.c(_0123_)
	);

	and_ii _2885_ (
		.a(new_net_1814),
		.b(new_net_2208),
		.c(_0124_)
	);

	and_bb _2886_ (
		.a(new_net_1815),
		.b(new_net_2209),
		.c(_0125_)
	);

	or_bb _2887_ (
		.a(new_net_3709),
		.b(new_net_2589),
		.c(_0126_)
	);

	or_bb _2888_ (
		.a(new_net_2665),
		.b(new_net_1992),
		.c(_0127_)
	);

	or_ii _2889_ (
		.a(new_net_2666),
		.b(new_net_1993),
		.c(_0128_)
	);

	or_ii _2890_ (
		.a(new_net_3710),
		.b(new_net_2627),
		.c(_0129_)
	);

	and_ii _2891_ (
		.a(new_net_3033),
		.b(new_net_1870),
		.c(_0130_)
	);

	and_bb _2892_ (
		.a(new_net_3034),
		.b(new_net_1871),
		.c(_0131_)
	);

	or_bb _2893_ (
		.a(new_net_3711),
		.b(new_net_2821),
		.c(_0133_)
	);

	or_bb _2894_ (
		.a(new_net_570),
		.b(new_net_1838),
		.c(_0134_)
	);

	or_ii _2895_ (
		.a(new_net_571),
		.b(new_net_1839),
		.c(_0135_)
	);

	or_ii _2896_ (
		.a(new_net_3712),
		.b(new_net_3003),
		.c(_0136_)
	);

	and_ii _2897_ (
		.a(new_net_1086),
		.b(new_net_1459),
		.c(_0137_)
	);

	and_bb _2898_ (
		.a(new_net_1087),
		.b(new_net_1460),
		.c(_0138_)
	);

	or_bb _2899_ (
		.a(new_net_3713),
		.b(new_net_3151),
		.c(_0139_)
	);

	or_bb _2900_ (
		.a(new_net_1660),
		.b(new_net_1758),
		.c(_0140_)
	);

	or_ii _2901_ (
		.a(new_net_1661),
		.b(new_net_1759),
		.c(_0141_)
	);

	or_ii _2902_ (
		.a(new_net_3714),
		.b(new_net_2122),
		.c(_0142_)
	);

	and_ii _2903_ (
		.a(new_net_2511),
		.b(new_net_1736),
		.c(_0144_)
	);

	and_bb _2904_ (
		.a(new_net_2512),
		.b(new_net_1737),
		.c(_0145_)
	);

	or_bb _2905_ (
		.a(new_net_3715),
		.b(new_net_2929),
		.c(_0146_)
	);

	or_bb _2906_ (
		.a(new_net_1782),
		.b(new_net_1704),
		.c(_0147_)
	);

	or_ii _2907_ (
		.a(new_net_1783),
		.b(new_net_1705),
		.c(_0148_)
	);

	or_ii _2908_ (
		.a(new_net_3716),
		.b(new_net_1834),
		.c(_0149_)
	);

	and_ii _2909_ (
		.a(new_net_1916),
		.b(new_net_735),
		.c(_0150_)
	);

	and_bb _2910_ (
		.a(new_net_1917),
		.b(new_net_736),
		.c(_0151_)
	);

	or_bb _2911_ (
		.a(new_net_3717),
		.b(new_net_1940),
		.c(_0152_)
	);

	or_bb _2912_ (
		.a(new_net_2012),
		.b(new_net_325),
		.c(_0153_)
	);

	or_ii _2913_ (
		.a(new_net_2013),
		.b(new_net_326),
		.c(_0155_)
	);

	or_ii _2914_ (
		.a(new_net_3718),
		.b(new_net_1364),
		.c(_0156_)
	);

	and_ii _2915_ (
		.a(new_net_2188),
		.b(new_net_3256),
		.c(_0157_)
	);

	and_bb _2916_ (
		.a(new_net_2189),
		.b(new_net_3257),
		.c(_0158_)
	);

	or_bb _2917_ (
		.a(new_net_3719),
		.b(new_net_2234),
		.c(_0159_)
	);

	or_bb _2918_ (
		.a(new_net_2515),
		.b(new_net_912),
		.c(_0160_)
	);

	or_ii _2919_ (
		.a(new_net_2516),
		.b(new_net_913),
		.c(_0161_)
	);

	or_ii _2920_ (
		.a(new_net_3720),
		.b(new_net_2366),
		.c(_0162_)
	);

	and_ii _2921_ (
		.a(new_net_3159),
		.b(new_net_721),
		.c(_0163_)
	);

	and_bb _2922_ (
		.a(new_net_3160),
		.b(new_net_722),
		.c(_0164_)
	);

	or_bb _2923_ (
		.a(new_net_3721),
		.b(new_net_2458),
		.c(_0166_)
	);

	or_bb _2924_ (
		.a(new_net_649),
		.b(new_net_516),
		.c(_0167_)
	);

	or_ii _2925_ (
		.a(new_net_650),
		.b(new_net_517),
		.c(_0168_)
	);

	or_ii _2926_ (
		.a(new_net_3722),
		.b(new_net_2639),
		.c(_0169_)
	);

	and_ii _2927_ (
		.a(new_net_2718),
		.b(new_net_3045),
		.c(_0170_)
	);

	and_bb _2928_ (
		.a(new_net_2719),
		.b(new_net_3046),
		.c(_0171_)
	);

	or_bb _2929_ (
		.a(new_net_3723),
		.b(new_net_1366),
		.c(_0172_)
	);

	or_bb _2930_ (
		.a(new_net_2805),
		.b(new_net_134),
		.c(_0173_)
	);

	or_ii _2931_ (
		.a(new_net_2806),
		.b(new_net_135),
		.c(_0174_)
	);

	or_ii _2932_ (
		.a(new_net_3724),
		.b(new_net_2859),
		.c(_0175_)
	);

	and_ii _2933_ (
		.a(new_net_2971),
		.b(new_net_3222),
		.c(_0177_)
	);

	and_bb _2934_ (
		.a(new_net_2972),
		.b(new_net_3223),
		.c(_0178_)
	);

	or_bb _2935_ (
		.a(new_net_3725),
		.b(new_net_3047),
		.c(_0179_)
	);

	or_bb _2936_ (
		.a(new_net_3163),
		.b(new_net_2927),
		.c(_0180_)
	);

	or_ii _2937_ (
		.a(new_net_3164),
		.b(new_net_2928),
		.c(_0181_)
	);

	or_ii _2938_ (
		.a(new_net_3726),
		.b(new_net_90),
		.c(_0182_)
	);

	and_ii _2939_ (
		.a(new_net_1612),
		.b(new_net_2857),
		.c(_0183_)
	);

	and_bb _2940_ (
		.a(new_net_1613),
		.b(new_net_2858),
		.c(_0184_)
	);

	or_bb _2941_ (
		.a(new_net_3727),
		.b(new_net_2519),
		.c(_0185_)
	);

	or_bb _2942_ (
		.a(new_net_2935),
		.b(new_net_2781),
		.c(_0186_)
	);

	or_ii _2943_ (
		.a(new_net_2936),
		.b(new_net_2782),
		.c(_0188_)
	);

	or_ii _2944_ (
		.a(new_net_3728),
		.b(new_net_1728),
		.c(_0189_)
	);

	and_ii _2945_ (
		.a(new_net_1844),
		.b(new_net_2180),
		.c(_0190_)
	);

	and_bb _2946_ (
		.a(new_net_1845),
		.b(new_net_2181),
		.c(_0191_)
	);

	or_bb _2947_ (
		.a(new_net_3729),
		.b(new_net_1876),
		.c(_0192_)
	);

	or_bb _2948_ (
		.a(new_net_1026),
		.b(new_net_1966),
		.c(_0193_)
	);

	or_ii _2949_ (
		.a(new_net_1027),
		.b(new_net_1967),
		.c(_0194_)
	);

	or_ii _2950_ (
		.a(new_net_3730),
		.b(new_net_1190),
		.c(_0195_)
	);

	and_ii _2951_ (
		.a(new_net_2064),
		.b(new_net_2667),
		.c(_0196_)
	);

	and_bb _2952_ (
		.a(new_net_2065),
		.b(new_net_2668),
		.c(_0197_)
	);

	or_bb _2953_ (
		.a(new_net_3731),
		.b(new_net_1738),
		.c(_0199_)
	);

	and_ii _2954_ (
		.a(new_net_2323),
		.b(new_net_1634),
		.c(_0200_)
	);

	and_bb _2955_ (
		.a(new_net_2324),
		.b(new_net_1635),
		.c(_0201_)
	);

	or_bb _2956_ (
		.a(new_net_3732),
		.b(new_net_2266),
		.c(_0202_)
	);

	or_bb _2957_ (
		.a(new_net_1562),
		.b(new_net_821),
		.c(_0203_)
	);

	and_bb _2958_ (
		.a(new_net_1229),
		.b(new_net_2461),
		.c(_0204_)
	);

	and_ii _2959_ (
		.a(new_net_3733),
		.b(new_net_1436),
		.c(_0205_)
	);

	or_bb _2960_ (
		.a(new_net_2468),
		.b(new_net_3167),
		.c(_0206_)
	);

	and_bi _2961_ (
		.a(new_net_2506),
		.b(new_net_2943),
		.c(_0207_)
	);

	and_bi _2962_ (
		.a(new_net_2944),
		.b(new_net_2508),
		.c(_0208_)
	);

	or_bb _2963_ (
		.a(new_net_3734),
		.b(new_net_669),
		.c(new_net_3936)
	);

	or_bb _2964_ (
		.a(new_net_670),
		.b(new_net_2267),
		.c(_0210_)
	);

	and_bi _2965_ (
		.a(new_net_1191),
		.b(new_net_1739),
		.c(_0211_)
	);

	and_bb _2966_ (
		.a(new_net_740),
		.b(new_net_929),
		.c(_0212_)
	);

	and_bi _2967_ (
		.a(new_net_1729),
		.b(new_net_1877),
		.c(_0213_)
	);

	and_bb _2968_ (
		.a(new_net_1420),
		.b(new_net_531),
		.c(_0214_)
	);

	and_bi _2969_ (
		.a(new_net_91),
		.b(new_net_2520),
		.c(_0215_)
	);

	and_bb _2970_ (
		.a(new_net_1472),
		.b(new_net_159),
		.c(_0216_)
	);

	and_bi _2971_ (
		.a(new_net_2860),
		.b(new_net_3048),
		.c(_0217_)
	);

	and_bb _2972_ (
		.a(new_net_3092),
		.b(new_net_432),
		.c(_0218_)
	);

	and_bi _2973_ (
		.a(new_net_2640),
		.b(new_net_1367),
		.c(_0220_)
	);

	and_bb _2974_ (
		.a(new_net_2341),
		.b(new_net_3023),
		.c(_0221_)
	);

	and_bi _2975_ (
		.a(new_net_2367),
		.b(new_net_2459),
		.c(_0222_)
	);

	and_bb _2976_ (
		.a(new_net_2618),
		.b(new_net_2398),
		.c(_0223_)
	);

	and_bi _2977_ (
		.a(new_net_1365),
		.b(new_net_2235),
		.c(_0224_)
	);

	and_bb _2978_ (
		.a(new_net_381),
		.b(new_net_270),
		.c(_0225_)
	);

	and_bi _2979_ (
		.a(new_net_1835),
		.b(new_net_1941),
		.c(_0226_)
	);

	and_bb _2980_ (
		.a(new_net_2503),
		.b(new_net_207),
		.c(_0227_)
	);

	and_bi _2981_ (
		.a(new_net_2123),
		.b(new_net_2930),
		.c(_0228_)
	);

	and_bb _2982_ (
		.a(new_net_1118),
		.b(new_net_1811),
		.c(_0229_)
	);

	and_bi _2983_ (
		.a(new_net_3004),
		.b(new_net_3152),
		.c(_0231_)
	);

	and_bb _2984_ (
		.a(new_net_1558),
		.b(new_net_1448),
		.c(_0232_)
	);

	and_bi _2985_ (
		.a(new_net_2628),
		.b(new_net_2822),
		.c(_0233_)
	);

	and_bb _2986_ (
		.a(new_net_2702),
		.b(new_net_1260),
		.c(_0234_)
	);

	and_bi _2987_ (
		.a(new_net_2433),
		.b(new_net_2590),
		.c(_0235_)
	);

	and_bb _2988_ (
		.a(new_net_2055),
		.b(new_net_3187),
		.c(_0236_)
	);

	and_bb _2989_ (
		.a(new_net_2862),
		.b(new_net_402),
		.c(_0237_)
	);

	and_ii _2990_ (
		.a(new_net_754),
		.b(new_net_2187),
		.c(_0238_)
	);

	and_ii _2991_ (
		.a(new_net_777),
		.b(new_net_568),
		.c(_0239_)
	);

	and_bb _2992_ (
		.a(new_net_778),
		.b(new_net_569),
		.c(_0240_)
	);

	or_bb _2993_ (
		.a(new_net_3735),
		.b(new_net_950),
		.c(_0242_)
	);

	and_ii _2994_ (
		.a(new_net_709),
		.b(new_net_466),
		.c(_0243_)
	);

	and_bb _2995_ (
		.a(new_net_710),
		.b(new_net_467),
		.c(_0244_)
	);

	or_bb _2996_ (
		.a(new_net_3736),
		.b(new_net_759),
		.c(_0245_)
	);

	and_ii _2997_ (
		.a(new_net_2004),
		.b(new_net_180),
		.c(_0246_)
	);

	and_bb _2998_ (
		.a(new_net_2005),
		.b(new_net_181),
		.c(_0247_)
	);

	or_bb _2999_ (
		.a(new_net_3737),
		.b(new_net_2220),
		.c(_0248_)
	);

	and_ii _3000_ (
		.a(new_net_942),
		.b(new_net_364),
		.c(_0249_)
	);

	and_bb _3001_ (
		.a(new_net_943),
		.b(new_net_365),
		.c(_0250_)
	);

	or_bb _3002_ (
		.a(new_net_3738),
		.b(new_net_2799),
		.c(_0251_)
	);

	and_ii _3003_ (
		.a(new_net_1012),
		.b(new_net_3031),
		.c(_0253_)
	);

	and_bb _3004_ (
		.a(new_net_1013),
		.b(new_net_3032),
		.c(_0254_)
	);

	or_bb _3005_ (
		.a(new_net_3739),
		.b(new_net_1080),
		.c(_0255_)
	);

	and_ii _3006_ (
		.a(new_net_785),
		.b(new_net_311),
		.c(_0256_)
	);

	and_bb _3007_ (
		.a(new_net_786),
		.b(new_net_312),
		.c(_0257_)
	);

	or_bb _3008_ (
		.a(new_net_3740),
		.b(new_net_954),
		.c(_0258_)
	);

	and_ii _3009_ (
		.a(new_net_1289),
		.b(new_net_279),
		.c(_0259_)
	);

	and_bb _3010_ (
		.a(new_net_1290),
		.b(new_net_280),
		.c(_0260_)
	);

	or_bb _3011_ (
		.a(new_net_3741),
		.b(new_net_1505),
		.c(_0261_)
	);

	and_ii _3012_ (
		.a(new_net_1824),
		.b(new_net_2214),
		.c(_0262_)
	);

	and_bb _3013_ (
		.a(new_net_1825),
		.b(new_net_2215),
		.c(_0264_)
	);

	or_bb _3014_ (
		.a(new_net_3742),
		.b(new_net_1421),
		.c(_0265_)
	);

	and_ii _3015_ (
		.a(new_net_2637),
		.b(new_net_174),
		.c(_0266_)
	);

	and_bb _3016_ (
		.a(new_net_2638),
		.b(new_net_175),
		.c(_0267_)
	);

	or_bb _3017_ (
		.a(new_net_3743),
		.b(new_net_1431),
		.c(_0268_)
	);

	and_ii _3018_ (
		.a(new_net_1690),
		.b(new_net_118),
		.c(_0269_)
	);

	and_bb _3019_ (
		.a(new_net_1691),
		.b(new_net_119),
		.c(_0270_)
	);

	or_bb _3020_ (
		.a(new_net_3744),
		.b(new_net_1962),
		.c(_0271_)
	);

	and_ii _3021_ (
		.a(new_net_2378),
		.b(new_net_94),
		.c(_0272_)
	);

	and_bb _3022_ (
		.a(new_net_2379),
		.b(new_net_95),
		.c(_0273_)
	);

	or_bb _3023_ (
		.a(new_net_3745),
		.b(new_net_2577),
		.c(_0275_)
	);

	and_ii _3024_ (
		.a(new_net_3215),
		.b(new_net_1491),
		.c(_0276_)
	);

	and_bb _3025_ (
		.a(new_net_3216),
		.b(new_net_1492),
		.c(_0277_)
	);

	or_bb _3026_ (
		.a(new_net_3746),
		.b(new_net_132),
		.c(_0278_)
	);

	and_ii _3027_ (
		.a(new_net_512),
		.b(new_net_1283),
		.c(_0279_)
	);

	and_bb _3028_ (
		.a(new_net_513),
		.b(new_net_1284),
		.c(_0280_)
	);

	or_bb _3029_ (
		.a(new_net_3747),
		.b(new_net_717),
		.c(_0281_)
	);

	and_ii _3030_ (
		.a(new_net_2158),
		.b(new_net_480),
		.c(_0282_)
	);

	and_bb _3031_ (
		.a(new_net_2159),
		.b(new_net_481),
		.c(_0283_)
	);

	or_bb _3032_ (
		.a(new_net_3748),
		.b(new_net_2192),
		.c(_0284_)
	);

	and_ii _3033_ (
		.a(new_net_1636),
		.b(new_net_3173),
		.c(_0286_)
	);

	and_bb _3034_ (
		.a(new_net_1637),
		.b(new_net_3174),
		.c(_0287_)
	);

	or_bb _3035_ (
		.a(new_net_3749),
		.b(new_net_2370),
		.c(_0288_)
	);

	and_ii _3036_ (
		.a(new_net_2426),
		.b(new_net_110),
		.c(_0289_)
	);

	and_bb _3037_ (
		.a(new_net_2427),
		.b(new_net_111),
		.c(_0290_)
	);

	or_bb _3038_ (
		.a(new_net_3750),
		.b(new_net_2462),
		.c(_0291_)
	);

	and_ii _3039_ (
		.a(new_net_2539),
		.b(new_net_3171),
		.c(_0292_)
	);

	and_bb _3040_ (
		.a(new_net_2540),
		.b(new_net_3172),
		.c(_0293_)
	);

	or_bb _3041_ (
		.a(new_net_3751),
		.b(new_net_3224),
		.c(_0294_)
	);

	and_ii _3042_ (
		.a(new_net_317),
		.b(new_net_2740),
		.c(_0295_)
	);

	and_bb _3043_ (
		.a(new_net_318),
		.b(new_net_2741),
		.c(_0297_)
	);

	or_bb _3044_ (
		.a(new_net_3752),
		.b(new_net_2726),
		.c(_0298_)
	);

	and_ii _3045_ (
		.a(new_net_1064),
		.b(new_net_2955),
		.c(_0299_)
	);

	and_bb _3046_ (
		.a(new_net_1065),
		.b(new_net_2956),
		.c(_0300_)
	);

	or_bb _3047_ (
		.a(new_net_3753),
		.b(new_net_1235),
		.c(_0301_)
	);

	and_ii _3048_ (
		.a(new_net_1638),
		.b(new_net_2331),
		.c(_0302_)
	);

	and_bb _3049_ (
		.a(new_net_1639),
		.b(new_net_2332),
		.c(_0303_)
	);

	or_bb _3050_ (
		.a(new_net_3754),
		.b(new_net_1774),
		.c(_0304_)
	);

	and_ii _3051_ (
		.a(new_net_3117),
		.b(new_net_2136),
		.c(_0305_)
	);

	and_bb _3052_ (
		.a(new_net_3118),
		.b(new_net_2137),
		.c(_0306_)
	);

	or_bb _3053_ (
		.a(new_net_3755),
		.b(new_net_2384),
		.c(_0308_)
	);

	and_ii _3054_ (
		.a(new_net_1602),
		.b(new_net_2815),
		.c(_0309_)
	);

	and_bb _3055_ (
		.a(new_net_1603),
		.b(new_net_2816),
		.c(_0310_)
	);

	or_bb _3056_ (
		.a(new_net_3756),
		.b(new_net_60),
		.c(_0311_)
	);

	and_ii _3057_ (
		.a(new_net_2130),
		.b(new_net_1742),
		.c(_0312_)
	);

	and_bb _3058_ (
		.a(new_net_2131),
		.b(new_net_1743),
		.c(_0313_)
	);

	or_bb _3059_ (
		.a(new_net_3757),
		.b(new_net_2321),
		.c(_0314_)
	);

	and_ii _3060_ (
		.a(new_net_232),
		.b(new_net_2752),
		.c(_0315_)
	);

	and_bb _3061_ (
		.a(new_net_233),
		.b(new_net_2753),
		.c(_0316_)
	);

	or_bb _3062_ (
		.a(new_net_3758),
		.b(new_net_2941),
		.c(_0317_)
	);

	and_ii _3063_ (
		.a(new_net_92),
		.b(new_net_1384),
		.c(_0319_)
	);

	and_bb _3064_ (
		.a(new_net_93),
		.b(new_net_1385),
		.c(_0320_)
	);

	or_bb _3065_ (
		.a(new_net_3759),
		.b(new_net_476),
		.c(_0321_)
	);

	and_bi _3066_ (
		.a(new_net_2673),
		.b(new_net_502),
		.c(_0322_)
	);

	and_bi _3067_ (
		.a(new_net_503),
		.b(new_net_2674),
		.c(_0323_)
	);

	or_bb _3068_ (
		.a(new_net_3760),
		.b(new_net_552),
		.c(new_net_3960)
	);

	or_bb _3069_ (
		.a(new_net_553),
		.b(new_net_477),
		.c(_0324_)
	);

	and_ii _3070_ (
		.a(new_net_2942),
		.b(new_net_2322),
		.c(_0325_)
	);

	and_bb _3071_ (
		.a(new_net_1417),
		.b(new_net_917),
		.c(_0326_)
	);

	and_ii _3072_ (
		.a(new_net_61),
		.b(new_net_2385),
		.c(_0327_)
	);

	and_bb _3073_ (
		.a(new_net_1470),
		.b(new_net_536),
		.c(_0329_)
	);

	and_ii _3074_ (
		.a(new_net_1775),
		.b(new_net_1236),
		.c(_0330_)
	);

	and_bb _3075_ (
		.a(new_net_3090),
		.b(new_net_150),
		.c(_0331_)
	);

	and_ii _3076_ (
		.a(new_net_2727),
		.b(new_net_3225),
		.c(_0332_)
	);

	and_bb _3077_ (
		.a(new_net_2340),
		.b(new_net_437),
		.c(_0333_)
	);

	and_ii _3078_ (
		.a(new_net_2463),
		.b(new_net_2371),
		.c(_0334_)
	);

	and_bb _3079_ (
		.a(new_net_3020),
		.b(new_net_2397),
		.c(_0335_)
	);

	and_ii _3080_ (
		.a(new_net_2193),
		.b(new_net_718),
		.c(_0336_)
	);

	and_bb _3081_ (
		.a(new_net_2611),
		.b(new_net_388),
		.c(_0337_)
	);

	and_ii _3082_ (
		.a(new_net_133),
		.b(new_net_2578),
		.c(_0338_)
	);

	and_bb _3083_ (
		.a(new_net_2501),
		.b(new_net_263),
		.c(_0340_)
	);

	and_ii _3084_ (
		.a(new_net_1963),
		.b(new_net_1432),
		.c(_0341_)
	);

	and_bb _3085_ (
		.a(new_net_1116),
		.b(new_net_213),
		.c(_0342_)
	);

	and_ii _3086_ (
		.a(new_net_1422),
		.b(new_net_1506),
		.c(_0343_)
	);

	and_bb _3087_ (
		.a(new_net_1555),
		.b(new_net_1801),
		.c(_0344_)
	);

	and_ii _3088_ (
		.a(new_net_955),
		.b(new_net_1081),
		.c(_0345_)
	);

	and_bb _3089_ (
		.a(new_net_2698),
		.b(new_net_1453),
		.c(_0346_)
	);

	and_ii _3090_ (
		.a(new_net_2800),
		.b(new_net_2221),
		.c(_0347_)
	);

	and_bb _3091_ (
		.a(new_net_2052),
		.b(new_net_1251),
		.c(_0348_)
	);

	and_bb _3092_ (
		.a(new_net_2875),
		.b(new_net_3188),
		.c(_0349_)
	);

	and_ii _3093_ (
		.a(new_net_760),
		.b(new_net_951),
		.c(_0351_)
	);

	and_ii _3094_ (
		.a(new_net_70),
		.b(new_net_1569),
		.c(_0352_)
	);

	and_bb _3095_ (
		.a(new_net_71),
		.b(new_net_1570),
		.c(_0353_)
	);

	or_bb _3096_ (
		.a(new_net_3761),
		.b(new_net_2767),
		.c(_0354_)
	);

	and_ii _3097_ (
		.a(new_net_170),
		.b(new_net_2746),
		.c(_0355_)
	);

	and_bb _3098_ (
		.a(new_net_171),
		.b(new_net_2747),
		.c(_0356_)
	);

	or_bb _3099_ (
		.a(new_net_3762),
		.b(new_net_196),
		.c(_0357_)
	);

	and_ii _3100_ (
		.a(new_net_281),
		.b(new_net_2529),
		.c(_0358_)
	);

	and_bb _3101_ (
		.a(new_net_282),
		.b(new_net_2530),
		.c(_0359_)
	);

	or_bb _3102_ (
		.a(new_net_3763),
		.b(new_net_723),
		.c(_0360_)
	);

	and_ii _3103_ (
		.a(new_net_374),
		.b(new_net_2337),
		.c(_0362_)
	);

	and_bb _3104_ (
		.a(new_net_375),
		.b(new_net_2338),
		.c(_0363_)
	);

	or_bb _3105_ (
		.a(new_net_3764),
		.b(new_net_472),
		.c(_0364_)
	);

	and_ii _3106_ (
		.a(new_net_558),
		.b(new_net_2142),
		.c(_0365_)
	);

	and_bb _3107_ (
		.a(new_net_559),
		.b(new_net_2143),
		.c(_0366_)
	);

	or_bb _3108_ (
		.a(new_net_3765),
		.b(new_net_1970),
		.c(_0367_)
	);

	and_ii _3109_ (
		.a(new_net_653),
		.b(new_net_1342),
		.c(_0368_)
	);

	and_bb _3110_ (
		.a(new_net_654),
		.b(new_net_1343),
		.c(_0369_)
	);

	or_bb _3111_ (
		.a(new_net_3766),
		.b(new_net_2583),
		.c(_0370_)
	);

	and_ii _3112_ (
		.a(new_net_2801),
		.b(new_net_1746),
		.c(_0371_)
	);

	and_bb _3113_ (
		.a(new_net_2802),
		.b(new_net_1747),
		.c(_0373_)
	);

	or_bb _3114_ (
		.a(new_net_3767),
		.b(new_net_3264),
		.c(_0374_)
	);

	and_ii _3115_ (
		.a(new_net_520),
		.b(new_net_1267),
		.c(_0375_)
	);

	and_bb _3116_ (
		.a(new_net_521),
		.b(new_net_1268),
		.c(_0376_)
	);

	or_bb _3117_ (
		.a(new_net_3768),
		.b(new_net_729),
		.c(_0377_)
	);

	and_ii _3118_ (
		.a(new_net_1018),
		.b(new_net_1220),
		.c(_0378_)
	);

	and_bb _3119_ (
		.a(new_net_1019),
		.b(new_net_1221),
		.c(_0379_)
	);

	or_bb _3120_ (
		.a(new_net_3769),
		.b(new_net_1239),
		.c(_0380_)
	);

	and_ii _3121_ (
		.a(new_net_1104),
		.b(new_net_1186),
		.c(_0381_)
	);

	and_bb _3122_ (
		.a(new_net_1105),
		.b(new_net_1187),
		.c(_0382_)
	);

	or_bb _3123_ (
		.a(new_net_3770),
		.b(new_net_1144),
		.c(_0384_)
	);

	and_ii _3124_ (
		.a(new_net_1265),
		.b(new_net_1108),
		.c(_0385_)
	);

	and_bb _3125_ (
		.a(new_net_1266),
		.b(new_net_1109),
		.c(_0386_)
	);

	or_bb _3126_ (
		.a(new_net_3771),
		.b(new_net_1316),
		.c(_0387_)
	);

	and_ii _3127_ (
		.a(new_net_3009),
		.b(new_net_1078),
		.c(_0388_)
	);

	and_bb _3128_ (
		.a(new_net_3010),
		.b(new_net_1079),
		.c(_0389_)
	);

	or_bb _3129_ (
		.a(new_net_3772),
		.b(new_net_3268),
		.c(_0390_)
	);

	and_ii _3130_ (
		.a(new_net_323),
		.b(new_net_478),
		.c(_0391_)
	);

	and_bb _3131_ (
		.a(new_net_324),
		.b(new_net_479),
		.c(_0392_)
	);

	or_bb _3132_ (
		.a(new_net_3773),
		.b(new_net_1571),
		.c(_0393_)
	);

	and_ii _3133_ (
		.a(new_net_908),
		.b(new_net_1024),
		.c(_0395_)
	);

	and_bb _3134_ (
		.a(new_net_909),
		.b(new_net_1025),
		.c(_0396_)
	);

	or_bb _3135_ (
		.a(new_net_3774),
		.b(new_net_1226),
		.c(_0397_)
	);

	and_ii _3136_ (
		.a(new_net_216),
		.b(new_net_996),
		.c(_0398_)
	);

	and_bb _3137_ (
		.a(new_net_217),
		.b(new_net_997),
		.c(_0399_)
	);

	or_bb _3138_ (
		.a(new_net_3775),
		.b(new_net_228),
		.c(_0400_)
	);

	and_ii _3139_ (
		.a(new_net_2178),
		.b(new_net_3169),
		.c(_0401_)
	);

	and_bb _3140_ (
		.a(new_net_2179),
		.b(new_net_3170),
		.c(_0402_)
	);

	or_bb _3141_ (
		.a(new_net_3776),
		.b(new_net_2380),
		.c(_0403_)
	);

	and_ii _3142_ (
		.a(new_net_2765),
		.b(new_net_944),
		.c(_0404_)
	);

	and_bb _3143_ (
		.a(new_net_2766),
		.b(new_net_945),
		.c(_0406_)
	);

	or_bb _3144_ (
		.a(new_net_3777),
		.b(new_net_2989),
		.c(_0407_)
	);

	and_ii _3145_ (
		.a(new_net_596),
		.b(new_net_900),
		.c(_0408_)
	);

	and_bb _3146_ (
		.a(new_net_597),
		.b(new_net_901),
		.c(_0409_)
	);

	or_bb _3147_ (
		.a(new_net_3778),
		.b(new_net_514),
		.c(_0410_)
	);

	and_ii _3148_ (
		.a(new_net_713),
		.b(new_net_2525),
		.c(_0411_)
	);

	and_bb _3149_ (
		.a(new_net_714),
		.b(new_net_2526),
		.c(_0412_)
	);

	or_bb _3150_ (
		.a(new_net_3779),
		.b(new_net_1062),
		.c(_0413_)
	);

	and_ii _3151_ (
		.a(new_net_848),
		.b(new_net_2327),
		.c(_0414_)
	);

	and_bb _3152_ (
		.a(new_net_849),
		.b(new_net_2328),
		.c(_0415_)
	);

	or_bb _3153_ (
		.a(new_net_3780),
		.b(new_net_880),
		.c(_0417_)
	);

	and_ii _3154_ (
		.a(new_net_2182),
		.b(new_net_1930),
		.c(_0418_)
	);

	and_bb _3155_ (
		.a(new_net_2183),
		.b(new_net_1931),
		.c(_0419_)
	);

	or_bb _3156_ (
		.a(new_net_3781),
		.b(new_net_990),
		.c(_0420_)
	);

	and_ii _3157_ (
		.a(new_net_1054),
		.b(new_net_711),
		.c(_0421_)
	);

	and_bb _3158_ (
		.a(new_net_1055),
		.b(new_net_712),
		.c(_0422_)
	);

	or_bb _3159_ (
		.a(new_net_3782),
		.b(new_net_2993),
		.c(_0423_)
	);

	and_ii _3160_ (
		.a(new_net_140),
		.b(new_net_651),
		.c(_0424_)
	);

	and_bb _3161_ (
		.a(new_net_141),
		.b(new_net_652),
		.c(_0425_)
	);

	or_bb _3162_ (
		.a(new_net_3783),
		.b(new_net_319),
		.c(_0426_)
	);

	and_bi _3163_ (
		.a(new_net_1382),
		.b(new_net_727),
		.c(_0428_)
	);

	and_bi _3164_ (
		.a(new_net_728),
		.b(new_net_1383),
		.c(_0429_)
	);

	or_bb _3165_ (
		.a(new_net_3784),
		.b(new_net_1338),
		.c(new_net_3934)
	);

	or_bb _3166_ (
		.a(new_net_1339),
		.b(new_net_320),
		.c(_0430_)
	);

	and_ii _3167_ (
		.a(new_net_2994),
		.b(new_net_991),
		.c(_0431_)
	);

	and_bb _3168_ (
		.a(new_net_1484),
		.b(new_net_923),
		.c(_0432_)
	);

	and_ii _3169_ (
		.a(new_net_881),
		.b(new_net_1063),
		.c(_0433_)
	);

	and_bb _3170_ (
		.a(new_net_3088),
		.b(new_net_539),
		.c(_0434_)
	);

	and_ii _3171_ (
		.a(new_net_515),
		.b(new_net_2990),
		.c(_0435_)
	);

	and_bb _3172_ (
		.a(new_net_2354),
		.b(new_net_153),
		.c(_0436_)
	);

	and_ii _3173_ (
		.a(new_net_2381),
		.b(new_net_229),
		.c(_0438_)
	);

	and_bb _3174_ (
		.a(new_net_433),
		.b(new_net_2410),
		.c(_0439_)
	);

	and_ii _3175_ (
		.a(new_net_1227),
		.b(new_net_1572),
		.c(_0440_)
	);

	and_bb _3176_ (
		.a(new_net_3024),
		.b(new_net_382),
		.c(_0441_)
	);

	and_ii _3177_ (
		.a(new_net_3269),
		.b(new_net_1317),
		.c(_0442_)
	);

	and_bb _3178_ (
		.a(new_net_2499),
		.b(new_net_2619),
		.c(_0443_)
	);

	and_ii _3179_ (
		.a(new_net_1145),
		.b(new_net_1240),
		.c(_0444_)
	);

	and_bb _3180_ (
		.a(new_net_1130),
		.b(new_net_265),
		.c(_0445_)
	);

	and_ii _3181_ (
		.a(new_net_730),
		.b(new_net_3265),
		.c(_0446_)
	);

	and_bb _3182_ (
		.a(new_net_1553),
		.b(new_net_214),
		.c(_0447_)
	);

	and_ii _3183_ (
		.a(new_net_2584),
		.b(new_net_1971),
		.c(_0449_)
	);

	and_bb _3184_ (
		.a(new_net_2713),
		.b(new_net_1803),
		.c(_0450_)
	);

	and_ii _3185_ (
		.a(new_net_473),
		.b(new_net_724),
		.c(_0451_)
	);

	and_bb _3186_ (
		.a(new_net_2047),
		.b(new_net_1455),
		.c(_0452_)
	);

	and_bb _3187_ (
		.a(new_net_2873),
		.b(new_net_1252),
		.c(_0453_)
	);

	and_ii _3188_ (
		.a(new_net_197),
		.b(new_net_2768),
		.c(_0454_)
	);

	and_ii _3189_ (
		.a(new_net_580),
		.b(new_net_350),
		.c(_0455_)
	);

	and_bb _3190_ (
		.a(new_net_581),
		.b(new_net_351),
		.c(_0456_)
	);

	or_bb _3191_ (
		.a(new_net_3785),
		.b(new_net_852),
		.c(_0457_)
	);

	and_ii _3192_ (
		.a(new_net_902),
		.b(new_net_184),
		.c(_0458_)
	);

	and_bb _3193_ (
		.a(new_net_903),
		.b(new_net_185),
		.c(_0460_)
	);

	or_bb _3194_ (
		.a(new_net_3786),
		.b(new_net_946),
		.c(_0461_)
	);

	and_ii _3195_ (
		.a(new_net_1854),
		.b(new_net_665),
		.c(_0462_)
	);

	and_bb _3196_ (
		.a(new_net_1855),
		.b(new_net_666),
		.c(_0463_)
	);

	or_bb _3197_ (
		.a(new_net_3787),
		.b(new_net_2032),
		.c(_0464_)
	);

	and_ii _3198_ (
		.a(new_net_2448),
		.b(new_net_3061),
		.c(_0465_)
	);

	and_bb _3199_ (
		.a(new_net_2449),
		.b(new_net_3062),
		.c(_0466_)
	);

	or_bb _3200_ (
		.a(new_net_3788),
		.b(new_net_1146),
		.c(_0467_)
	);

	and_ii _3201_ (
		.a(new_net_3069),
		.b(new_net_598),
		.c(_0468_)
	);

	and_bb _3202_ (
		.a(new_net_3070),
		.b(new_net_599),
		.c(_0469_)
	);

	or_bb _3203_ (
		.a(new_net_3789),
		.b(new_net_16),
		.c(_0471_)
	);

	and_ii _3204_ (
		.a(new_net_586),
		.b(new_net_498),
		.c(_0472_)
	);

	and_bb _3205_ (
		.a(new_net_587),
		.b(new_net_499),
		.c(_0473_)
	);

	or_bb _3206_ (
		.a(new_net_3790),
		.b(new_net_810),
		.c(_0474_)
	);

	and_ii _3207_ (
		.a(new_net_1100),
		.b(new_net_2244),
		.c(_0475_)
	);

	and_bb _3208_ (
		.a(new_net_1101),
		.b(new_net_2245),
		.c(_0476_)
	);

	or_bb _3209_ (
		.a(new_net_3791),
		.b(new_net_1308),
		.c(_0477_)
	);

	and_ii _3210_ (
		.a(new_net_74),
		.b(new_net_2026),
		.c(_0478_)
	);

	and_bb _3211_ (
		.a(new_net_75),
		.b(new_net_2027),
		.c(_0479_)
	);

	or_bb _3212_ (
		.a(new_net_3792),
		.b(new_net_2024),
		.c(_0480_)
	);

	and_ii _3213_ (
		.a(new_net_164),
		.b(new_net_1846),
		.c(_0482_)
	);

	and_bb _3214_ (
		.a(new_net_165),
		.b(new_net_1847),
		.c(_0483_)
	);

	or_bb _3215_ (
		.a(new_net_3793),
		.b(new_net_240),
		.c(_0484_)
	);

	and_ii _3216_ (
		.a(new_net_309),
		.b(new_net_1674),
		.c(_0485_)
	);

	and_bb _3217_ (
		.a(new_net_310),
		.b(new_net_1675),
		.c(_0486_)
	);

	or_bb _3218_ (
		.a(new_net_3794),
		.b(new_net_186),
		.c(_0487_)
	);

	and_ii _3219_ (
		.a(new_net_418),
		.b(new_net_1511),
		.c(_0488_)
	);

	and_bb _3220_ (
		.a(new_net_419),
		.b(new_net_1512),
		.c(_0489_)
	);

	or_bb _3221_ (
		.a(new_net_3795),
		.b(new_net_803),
		.c(_0490_)
	);

	and_ii _3222_ (
		.a(new_net_1098),
		.b(new_net_1302),
		.c(_0491_)
	);

	and_bb _3223_ (
		.a(new_net_1099),
		.b(new_net_1303),
		.c(_0493_)
	);

	or_bb _3224_ (
		.a(new_net_3796),
		.b(new_net_604),
		.c(_0494_)
	);

	and_ii _3225_ (
		.a(new_net_1858),
		.b(new_net_230),
		.c(_0495_)
	);

	and_bb _3226_ (
		.a(new_net_1859),
		.b(new_net_231),
		.c(_0496_)
	);

	or_bb _3227_ (
		.a(new_net_3797),
		.b(new_net_2034),
		.c(_0497_)
	);

	and_ii _3228_ (
		.a(new_net_846),
		.b(new_net_194),
		.c(_0498_)
	);

	and_bb _3229_ (
		.a(new_net_847),
		.b(new_net_195),
		.c(_0499_)
	);

	or_bb _3230_ (
		.a(new_net_3798),
		.b(new_net_2657),
		.c(_0500_)
	);

	and_ii _3231_ (
		.a(new_net_3073),
		.b(new_net_789),
		.c(_0501_)
	);

	and_bb _3232_ (
		.a(new_net_3074),
		.b(new_net_790),
		.c(_0502_)
	);

	or_bb _3233_ (
		.a(new_net_3799),
		.b(new_net_972),
		.c(_0504_)
	);

	and_ii _3234_ (
		.a(new_net_590),
		.b(new_net_106),
		.c(_0505_)
	);

	and_bb _3235_ (
		.a(new_net_591),
		.b(new_net_107),
		.c(_0506_)
	);

	or_bb _3236_ (
		.a(new_net_3800),
		.b(new_net_816),
		.c(_0507_)
	);

	and_ii _3237_ (
		.a(new_net_1150),
		.b(new_net_66),
		.c(_0508_)
	);

	and_bb _3238_ (
		.a(new_net_1151),
		.b(new_net_67),
		.c(_0509_)
	);

	or_bb _3239_ (
		.a(new_net_3801),
		.b(new_net_1180),
		.c(_0510_)
	);

	and_ii _3240_ (
		.a(new_net_1271),
		.b(new_net_26),
		.c(_0511_)
	);

	and_bb _3241_ (
		.a(new_net_1272),
		.b(new_net_27),
		.c(_0512_)
	);

	or_bb _3242_ (
		.a(new_net_3802),
		.b(new_net_1862),
		.c(_0513_)
	);

	and_ii _3243_ (
		.a(new_net_2254),
		.b(new_net_1972),
		.c(_0515_)
	);

	and_bb _3244_ (
		.a(new_net_2255),
		.b(new_net_1973),
		.c(_0516_)
	);

	or_bb _3245_ (
		.a(new_net_3803),
		.b(new_net_2659),
		.c(_0517_)
	);

	and_ii _3246_ (
		.a(new_net_1575),
		.b(new_net_1778),
		.c(_0518_)
	);

	and_bb _3247_ (
		.a(new_net_1576),
		.b(new_net_1779),
		.c(_0519_)
	);

	or_bb _3248_ (
		.a(new_net_3804),
		.b(new_net_1616),
		.c(_0520_)
	);

	and_ii _3249_ (
		.a(new_net_1684),
		.b(new_net_1463),
		.c(_0521_)
	);

	and_bb _3250_ (
		.a(new_net_1685),
		.b(new_net_1464),
		.c(_0522_)
	);

	and_ii _3251_ (
		.a(new_net_3805),
		.b(new_net_1293),
		.c(_0523_)
	);

	and_bb _3252_ (
		.a(new_net_1668),
		.b(new_net_1437),
		.c(_0524_)
	);

	and_ii _3253_ (
		.a(new_net_1669),
		.b(new_net_1438),
		.c(_0526_)
	);

	or_bb _3254_ (
		.a(new_net_3806),
		.b(new_net_1828),
		.c(new_net_3970)
	);

	or_bb _3255_ (
		.a(new_net_1829),
		.b(new_net_1294),
		.c(_0527_)
	);

	and_ii _3256_ (
		.a(new_net_1617),
		.b(new_net_2660),
		.c(_0528_)
	);

	and_bb _3257_ (
		.a(new_net_3086),
		.b(new_net_925),
		.c(_0529_)
	);

	and_ii _3258_ (
		.a(new_net_1863),
		.b(new_net_1181),
		.c(_0530_)
	);

	and_bb _3259_ (
		.a(new_net_2352),
		.b(new_net_529),
		.c(_0531_)
	);

	and_ii _3260_ (
		.a(new_net_817),
		.b(new_net_973),
		.c(_0532_)
	);

	and_bb _3261_ (
		.a(new_net_151),
		.b(new_net_2409),
		.c(_0533_)
	);

	and_ii _3262_ (
		.a(new_net_2658),
		.b(new_net_2035),
		.c(_0534_)
	);

	and_bb _3263_ (
		.a(new_net_390),
		.b(new_net_431),
		.c(_0536_)
	);

	and_ii _3264_ (
		.a(new_net_605),
		.b(new_net_804),
		.c(_0537_)
	);

	and_bb _3265_ (
		.a(new_net_2496),
		.b(new_net_3021),
		.c(_0538_)
	);

	and_ii _3266_ (
		.a(new_net_187),
		.b(new_net_241),
		.c(_0539_)
	);

	and_bb _3267_ (
		.a(new_net_1127),
		.b(new_net_2612),
		.c(_0540_)
	);

	and_ii _3268_ (
		.a(new_net_2025),
		.b(new_net_1309),
		.c(_0541_)
	);

	and_bb _3269_ (
		.a(new_net_1549),
		.b(new_net_268),
		.c(_0542_)
	);

	and_ii _3270_ (
		.a(new_net_811),
		.b(new_net_17),
		.c(_0543_)
	);

	and_bb _3271_ (
		.a(new_net_2709),
		.b(new_net_205),
		.c(_0544_)
	);

	and_ii _3272_ (
		.a(new_net_1147),
		.b(new_net_2033),
		.c(_0545_)
	);

	and_bb _3273_ (
		.a(new_net_2043),
		.b(new_net_1809),
		.c(_0547_)
	);

	and_bb _3274_ (
		.a(new_net_2872),
		.b(new_net_1456),
		.c(_0548_)
	);

	and_ii _3275_ (
		.a(new_net_947),
		.b(new_net_853),
		.c(_0549_)
	);

	and_ii _3276_ (
		.a(new_net_2771),
		.b(new_net_12),
		.c(_0550_)
	);

	and_bb _3277_ (
		.a(new_net_2772),
		.b(new_net_13),
		.c(_0551_)
	);

	or_bb _3278_ (
		.a(new_net_3807),
		.b(new_net_2817),
		.c(_0552_)
	);

	and_ii _3279_ (
		.a(new_net_805),
		.b(new_net_3065),
		.c(_0553_)
	);

	and_bb _3280_ (
		.a(new_net_806),
		.b(new_net_3066),
		.c(_0554_)
	);

	or_bb _3281_ (
		.a(new_net_3808),
		.b(new_net_2957),
		.c(_0555_)
	);

	and_ii _3282_ (
		.a(new_net_3051),
		.b(new_net_2645),
		.c(_0556_)
	);

	and_bb _3283_ (
		.a(new_net_3052),
		.b(new_net_2646),
		.c(_0558_)
	);

	or_bb _3284_ (
		.a(new_net_3809),
		.b(new_net_1521),
		.c(_0559_)
	);

	and_ii _3285_ (
		.a(new_net_2036),
		.b(new_net_2444),
		.c(_0560_)
	);

	and_bb _3286_ (
		.a(new_net_2037),
		.b(new_net_2445),
		.c(_0561_)
	);

	or_bb _3287_ (
		.a(new_net_3810),
		.b(new_net_1614),
		.c(_0562_)
	);

	and_ii _3288_ (
		.a(new_net_1682),
		.b(new_net_2565),
		.c(_0563_)
	);

	and_bb _3289_ (
		.a(new_net_1683),
		.b(new_net_2566),
		.c(_0564_)
	);

	or_bb _3290_ (
		.a(new_net_3811),
		.b(new_net_2732),
		.c(_0565_)
	);

	and_ii _3291_ (
		.a(new_net_3157),
		.b(new_net_2486),
		.c(_0566_)
	);

	and_bb _3292_ (
		.a(new_net_3158),
		.b(new_net_2487),
		.c(_0567_)
	);

	or_bb _3293_ (
		.a(new_net_3812),
		.b(new_net_82),
		.c(_0569_)
	);

	and_ii _3294_ (
		.a(new_net_645),
		.b(new_net_1850),
		.c(_0570_)
	);

	and_bb _3295_ (
		.a(new_net_646),
		.b(new_net_1851),
		.c(_0571_)
	);

	or_bb _3296_ (
		.a(new_net_3813),
		.b(new_net_1942),
		.c(_0572_)
	);

	and_ii _3297_ (
		.a(new_net_1170),
		.b(new_net_1696),
		.c(_0573_)
	);

	and_bb _3298_ (
		.a(new_net_1171),
		.b(new_net_1697),
		.c(_0574_)
	);

	or_bb _3299_ (
		.a(new_net_3814),
		.b(new_net_2074),
		.c(_0575_)
	);

	and_ii _3300_ (
		.a(new_net_2154),
		.b(new_net_1513),
		.c(_0576_)
	);

	and_bb _3301_ (
		.a(new_net_2155),
		.b(new_net_1514),
		.c(_0577_)
	);

	or_bb _3302_ (
		.a(new_net_3815),
		.b(new_net_1924),
		.c(_0578_)
	);

	and_ii _3303_ (
		.a(new_net_2270),
		.b(new_net_2359),
		.c(_0580_)
	);

	and_bb _3304_ (
		.a(new_net_2271),
		.b(new_net_2360),
		.c(_0581_)
	);

	or_bb _3305_ (
		.a(new_net_3816),
		.b(new_net_2368),
		.c(_0582_)
	);

	and_ii _3306_ (
		.a(new_net_2436),
		.b(new_net_2302),
		.c(_0583_)
	);

	and_bb _3307_ (
		.a(new_net_2437),
		.b(new_net_2303),
		.c(_0584_)
	);

	or_bb _3308_ (
		.a(new_net_3817),
		.b(new_net_2456),
		.c(_0585_)
	);

	and_ii _3309_ (
		.a(new_net_462),
		.b(new_net_2260),
		.c(_0586_)
	);

	and_bb _3310_ (
		.a(new_net_463),
		.b(new_net_2261),
		.c(_0587_)
	);

	or_bb _3311_ (
		.a(new_net_3818),
		.b(new_net_2587),
		.c(_0588_)
	);

	and_ii _3312_ (
		.a(new_net_1010),
		.b(new_net_2196),
		.c(_0589_)
	);

	and_bb _3313_ (
		.a(new_net_1011),
		.b(new_net_2197),
		.c(_0591_)
	);

	or_bb _3314_ (
		.a(new_net_3819),
		.b(new_net_2720),
		.c(_0592_)
	);

	and_ii _3315_ (
		.a(new_net_2807),
		.b(new_net_2160),
		.c(_0593_)
	);

	and_bb _3316_ (
		.a(new_net_2808),
		.b(new_net_2161),
		.c(_0594_)
	);

	or_bb _3317_ (
		.a(new_net_3820),
		.b(new_net_1926),
		.c(_0595_)
	);

	and_ii _3318_ (
		.a(new_net_2317),
		.b(new_net_2112),
		.c(_0596_)
	);

	and_bb _3319_ (
		.a(new_net_2318),
		.b(new_net_2113),
		.c(_0597_)
	);

	or_bb _3320_ (
		.a(new_net_3821),
		.b(new_net_2521),
		.c(_0598_)
	);

	and_ii _3321_ (
		.a(new_net_2937),
		.b(new_net_2060),
		.c(_0599_)
	);

	and_bb _3322_ (
		.a(new_net_2938),
		.b(new_net_2061),
		.c(_0600_)
	);

	or_bb _3323_ (
		.a(new_net_3822),
		.b(new_net_3161),
		.c(_0602_)
	);

	and_ii _3324_ (
		.a(new_net_2689),
		.b(new_net_3057),
		.c(_0603_)
	);

	and_bb _3325_ (
		.a(new_net_2690),
		.b(new_net_3058),
		.c(_0604_)
	);

	or_bb _3326_ (
		.a(new_net_3823),
		.b(new_net_2893),
		.c(_0605_)
	);

	and_ii _3327_ (
		.a(new_net_76),
		.b(new_net_1980),
		.c(_0606_)
	);

	and_bb _3328_ (
		.a(new_net_77),
		.b(new_net_1981),
		.c(_0607_)
	);

	or_bb _3329_ (
		.a(new_net_3824),
		.b(new_net_242),
		.c(_0608_)
	);

	and_ii _3330_ (
		.a(new_net_633),
		.b(new_net_1950),
		.c(_0609_)
	);

	and_bb _3331_ (
		.a(new_net_634),
		.b(new_net_1951),
		.c(_0610_)
	);

	and_ii _3332_ (
		.a(new_net_3825),
		.b(new_net_273),
		.c(_0611_)
	);

	and_bb _3333_ (
		.a(new_net_341),
		.b(new_net_2424),
		.c(_0613_)
	);

	and_ii _3334_ (
		.a(new_net_342),
		.b(new_net_2425),
		.c(_0614_)
	);

	or_bb _3335_ (
		.a(new_net_3826),
		.b(new_net_1592),
		.c(new_net_3966)
	);

	or_bb _3336_ (
		.a(new_net_1593),
		.b(new_net_274),
		.c(_0615_)
	);

	and_ii _3337_ (
		.a(new_net_243),
		.b(new_net_2894),
		.c(_0616_)
	);

	and_bb _3338_ (
		.a(new_net_2342),
		.b(new_net_930),
		.c(_0617_)
	);

	and_ii _3339_ (
		.a(new_net_3162),
		.b(new_net_2522),
		.c(_0618_)
	);

	and_bb _3340_ (
		.a(new_net_2411),
		.b(new_net_532),
		.c(_0619_)
	);

	and_ii _3341_ (
		.a(new_net_1927),
		.b(new_net_2721),
		.c(_0620_)
	);

	and_bb _3342_ (
		.a(new_net_154),
		.b(new_net_391),
		.c(_0621_)
	);

	and_ii _3343_ (
		.a(new_net_2588),
		.b(new_net_2457),
		.c(_0622_)
	);

	and_bb _3344_ (
		.a(new_net_2504),
		.b(new_net_434),
		.c(_0623_)
	);

	and_ii _3345_ (
		.a(new_net_2369),
		.b(new_net_1925),
		.c(_0624_)
	);

	and_bb _3346_ (
		.a(new_net_1119),
		.b(new_net_3025),
		.c(_0625_)
	);

	and_ii _3347_ (
		.a(new_net_2075),
		.b(new_net_1943),
		.c(_0626_)
	);

	and_bb _3348_ (
		.a(new_net_1559),
		.b(new_net_2614),
		.c(_0627_)
	);

	and_ii _3349_ (
		.a(new_net_83),
		.b(new_net_2733),
		.c(_0628_)
	);

	and_bb _3350_ (
		.a(new_net_2703),
		.b(new_net_271),
		.c(_0629_)
	);

	and_ii _3351_ (
		.a(new_net_1615),
		.b(new_net_1522),
		.c(_0630_)
	);

	and_bb _3352_ (
		.a(new_net_2056),
		.b(new_net_208),
		.c(_0631_)
	);

	and_bb _3353_ (
		.a(new_net_2864),
		.b(new_net_1808),
		.c(_0634_)
	);

	and_ii _3354_ (
		.a(new_net_2958),
		.b(new_net_2818),
		.c(_0635_)
	);

	and_ii _3355_ (
		.a(new_net_1222),
		.b(new_net_2311),
		.c(_0636_)
	);

	and_bb _3356_ (
		.a(new_net_1223),
		.b(new_net_2312),
		.c(_0637_)
	);

	or_bb _3357_ (
		.a(new_net_3827),
		.b(new_net_2730),
		.c(_0638_)
	);

	and_ii _3358_ (
		.a(new_net_3155),
		.b(new_net_1074),
		.c(_0639_)
	);

	and_bb _3359_ (
		.a(new_net_3156),
		.b(new_net_1075),
		.c(_0640_)
	);

	or_bb _3360_ (
		.a(new_net_3828),
		.b(new_net_80),
		.c(_0641_)
	);

	and_ii _3361_ (
		.a(new_net_456),
		.b(new_net_1044),
		.c(_0642_)
	);

	and_bb _3362_ (
		.a(new_net_457),
		.b(new_net_1045),
		.c(_0643_)
	);

	or_bb _3363_ (
		.a(new_net_3829),
		.b(new_net_643),
		.c(_0645_)
	);

	and_ii _3364_ (
		.a(new_net_2787),
		.b(new_net_1360),
		.c(_0646_)
	);

	and_bb _3365_ (
		.a(new_net_2788),
		.b(new_net_1361),
		.c(_0647_)
	);

	or_bb _3366_ (
		.a(new_net_3830),
		.b(new_net_3005),
		.c(_0648_)
	);

	and_ii _3367_ (
		.a(new_net_166),
		.b(new_net_1168),
		.c(_0649_)
	);

	and_bb _3368_ (
		.a(new_net_167),
		.b(new_net_1169),
		.c(_0650_)
	);

	or_bb _3369_ (
		.a(new_net_3831),
		.b(new_net_321),
		.c(_0651_)
	);

	and_ii _3370_ (
		.a(new_net_731),
		.b(new_net_978),
		.c(_0652_)
	);

	and_bb _3371_ (
		.a(new_net_732),
		.b(new_net_979),
		.c(_0653_)
	);

	or_bb _3372_ (
		.a(new_net_3832),
		.b(new_net_914),
		.c(_0654_)
	);

	and_ii _3373_ (
		.a(new_net_1241),
		.b(new_net_934),
		.c(_0656_)
	);

	and_bb _3374_ (
		.a(new_net_1242),
		.b(new_net_935),
		.c(_0657_)
	);

	or_bb _3375_ (
		.a(new_net_3833),
		.b(new_net_1654),
		.c(_0658_)
	);

	and_ii _3376_ (
		.a(new_net_1988),
		.b(new_net_637),
		.c(_0659_)
	);

	and_bb _3377_ (
		.a(new_net_1989),
		.b(new_net_638),
		.c(_0660_)
	);

	or_bb _3378_ (
		.a(new_net_3834),
		.b(new_net_2202),
		.c(_0661_)
	);

	and_ii _3379_ (
		.a(new_net_2603),
		.b(new_net_452),
		.c(_0662_)
	);

	and_bb _3380_ (
		.a(new_net_2604),
		.b(new_net_453),
		.c(_0663_)
	);

	or_bb _3381_ (
		.a(new_net_3835),
		.b(new_net_701),
		.c(_0664_)
	);

	and_ii _3382_ (
		.a(new_net_3272),
		.b(new_net_246),
		.c(_0665_)
	);

	and_bb _3383_ (
		.a(new_net_3273),
		.b(new_net_247),
		.c(_0667_)
	);

	or_bb _3384_ (
		.a(new_net_3836),
		.b(new_net_144),
		.c(_0668_)
	);

	and_ii _3385_ (
		.a(new_net_936),
		.b(new_net_78),
		.c(_0669_)
	);

	and_bb _3386_ (
		.a(new_net_937),
		.b(new_net_79),
		.c(_0670_)
	);

	or_bb _3387_ (
		.a(new_net_3837),
		.b(new_net_964),
		.c(_0671_)
	);

	and_ii _3388_ (
		.a(new_net_1263),
		.b(new_net_767),
		.c(_0672_)
	);

	and_bb _3389_ (
		.a(new_net_1264),
		.b(new_net_768),
		.c(_0673_)
	);

	or_bb _3390_ (
		.a(new_net_3838),
		.b(new_net_1461),
		.c(_0674_)
	);

	and_ii _3391_ (
		.a(new_net_1112),
		.b(new_net_2899),
		.c(_0675_)
	);

	and_bb _3392_ (
		.a(new_net_1113),
		.b(new_net_2900),
		.c(_0676_)
	);

	or_bb _3393_ (
		.a(new_net_3839),
		.b(new_net_1152),
		.c(_0678_)
	);

	and_ii _3394_ (
		.a(new_net_2623),
		.b(new_net_657),
		.c(_0679_)
	);

	and_bb _3395_ (
		.a(new_net_2624),
		.b(new_net_658),
		.c(_0680_)
	);

	or_bb _3396_ (
		.a(new_net_3840),
		.b(new_net_2793),
		.c(_0681_)
	);

	and_ii _3397_ (
		.a(new_net_1370),
		.b(new_net_616),
		.c(_0682_)
	);

	and_bb _3398_ (
		.a(new_net_1371),
		.b(new_net_617),
		.c(_0683_)
	);

	or_bb _3399_ (
		.a(new_net_3841),
		.b(new_net_162),
		.c(_0684_)
	);

	and_ii _3400_ (
		.a(new_net_546),
		.b(new_net_2284),
		.c(_0685_)
	);

	and_bb _3401_ (
		.a(new_net_547),
		.b(new_net_2285),
		.c(_0686_)
	);

	or_bb _3402_ (
		.a(new_net_3842),
		.b(new_net_755),
		.c(_0687_)
	);

	and_ii _3403_ (
		.a(new_net_64),
		.b(new_net_562),
		.c(_0689_)
	);

	and_bb _3404_ (
		.a(new_net_65),
		.b(new_net_563),
		.c(_0690_)
	);

	and_ii _3405_ (
		.a(new_net_3843),
		.b(new_net_122),
		.c(_0691_)
	);

	and_bb _3406_ (
		.a(new_net_639),
		.b(new_net_508),
		.c(_0692_)
	);

	and_ii _3407_ (
		.a(new_net_640),
		.b(new_net_509),
		.c(_0693_)
	);

	or_bb _3408_ (
		.a(new_net_3844),
		.b(new_net_866),
		.c(new_net_3944)
	);

	or_bb _3409_ (
		.a(new_net_867),
		.b(new_net_123),
		.c(_0694_)
	);

	and_ii _3410_ (
		.a(new_net_756),
		.b(new_net_163),
		.c(_0695_)
	);

	and_bb _3411_ (
		.a(new_net_931),
		.b(new_net_2399),
		.c(_0696_)
	);

	and_ii _3412_ (
		.a(new_net_2794),
		.b(new_net_1153),
		.c(_0697_)
	);

	and_bb _3413_ (
		.a(new_net_383),
		.b(new_net_533),
		.c(_0699_)
	);

	and_ii _3414_ (
		.a(new_net_1462),
		.b(new_net_965),
		.c(_0700_)
	);

	and_bb _3415_ (
		.a(new_net_2500),
		.b(new_net_152),
		.c(_0701_)
	);

	and_ii _3416_ (
		.a(new_net_145),
		.b(new_net_702),
		.c(_0702_)
	);

	and_bb _3417_ (
		.a(new_net_1120),
		.b(new_net_438),
		.c(_0703_)
	);

	and_ii _3418_ (
		.a(new_net_2203),
		.b(new_net_1655),
		.c(_0704_)
	);

	and_bb _3419_ (
		.a(new_net_1550),
		.b(new_net_3016),
		.c(_0705_)
	);

	and_ii _3420_ (
		.a(new_net_915),
		.b(new_net_322),
		.c(_0706_)
	);

	and_bb _3421_ (
		.a(new_net_2710),
		.b(new_net_2617),
		.c(_0707_)
	);

	and_ii _3422_ (
		.a(new_net_3006),
		.b(new_net_644),
		.c(_0708_)
	);

	and_bb _3423_ (
		.a(new_net_2053),
		.b(new_net_269),
		.c(_0710_)
	);

	and_bb _3424_ (
		.a(new_net_2865),
		.b(new_net_215),
		.c(_0711_)
	);

	and_ii _3425_ (
		.a(new_net_81),
		.b(new_net_2731),
		.c(_0712_)
	);

	and_ii _3426_ (
		.a(new_net_994),
		.b(new_net_974),
		.c(_0713_)
	);

	and_bb _3427_ (
		.a(new_net_995),
		.b(new_net_975),
		.c(_0714_)
	);

	or_bb _3428_ (
		.a(new_net_3845),
		.b(new_net_1014),
		.c(_0715_)
	);

	and_ii _3429_ (
		.a(new_net_1084),
		.b(new_net_1008),
		.c(_0716_)
	);

	and_bb _3430_ (
		.a(new_net_1085),
		.b(new_net_1009),
		.c(_0717_)
	);

	or_bb _3431_ (
		.a(new_net_3846),
		.b(new_net_2128),
		.c(_0718_)
	);

	and_ii _3432_ (
		.a(new_net_2517),
		.b(new_net_647),
		.c(_0719_)
	);

	and_bb _3433_ (
		.a(new_net_2518),
		.b(new_net_648),
		.c(_0721_)
	);

	or_bb _3434_ (
		.a(new_net_3847),
		.b(new_net_1208),
		.c(_0722_)
	);

	and_ii _3435_ (
		.a(new_net_1334),
		.b(new_net_458),
		.c(_0723_)
	);

	and_bb _3436_ (
		.a(new_net_1335),
		.b(new_net_459),
		.c(_0724_)
	);

	or_bb _3437_ (
		.a(new_net_3848),
		.b(new_net_252),
		.c(_0725_)
	);

	and_ii _3438_ (
		.a(new_net_1487),
		.b(new_net_250),
		.c(_0726_)
	);

	and_bb _3439_ (
		.a(new_net_1488),
		.b(new_net_251),
		.c(_0727_)
	);

	or_bb _3440_ (
		.a(new_net_3849),
		.b(new_net_1525),
		.c(_0728_)
	);

	and_ii _3441_ (
		.a(new_net_34),
		.b(new_net_84),
		.c(_0729_)
	);

	and_bb _3442_ (
		.a(new_net_35),
		.b(new_net_85),
		.c(_0730_)
	);

	or_bb _3443_ (
		.a(new_net_3850),
		.b(new_net_62),
		.c(_0732_)
	);

	and_ii _3444_ (
		.a(new_net_572),
		.b(new_net_705),
		.c(_0733_)
	);

	and_bb _3445_ (
		.a(new_net_573),
		.b(new_net_706),
		.c(_0734_)
	);

	or_bb _3446_ (
		.a(new_net_3851),
		.b(new_net_779),
		.c(_0735_)
	);

	and_ii _3447_ (
		.a(new_net_1088),
		.b(new_net_661),
		.c(_0736_)
	);

	and_bb _3448_ (
		.a(new_net_1089),
		.b(new_net_662),
		.c(_0737_)
	);

	or_bb _3449_ (
		.a(new_net_3852),
		.b(new_net_313),
		.c(_0738_)
	);

	and_ii _3450_ (
		.a(new_net_1662),
		.b(new_net_2734),
		.c(_0739_)
	);

	and_bb _3451_ (
		.a(new_net_1663),
		.b(new_net_2735),
		.c(_0740_)
	);

	or_bb _3452_ (
		.a(new_net_3853),
		.b(new_net_1820),
		.c(_0741_)
	);

	and_ii _3453_ (
		.a(new_net_2224),
		.b(new_net_2513),
		.c(_0743_)
	);

	and_bb _3454_ (
		.a(new_net_2225),
		.b(new_net_2514),
		.c(_0744_)
	);

	or_bb _3455_ (
		.a(new_net_3854),
		.b(new_net_594),
		.c(_0745_)
	);

	and_ii _3456_ (
		.a(new_net_3039),
		.b(new_net_2313),
		.c(_0746_)
	);

	and_bb _3457_ (
		.a(new_net_3040),
		.b(new_net_2314),
		.c(_0747_)
	);

	or_bb _3458_ (
		.a(new_net_3855),
		.b(new_net_8),
		.c(_0748_)
	);

	and_ii _3459_ (
		.a(new_net_824),
		.b(new_net_2124),
		.c(_0749_)
	);

	and_bb _3460_ (
		.a(new_net_825),
		.b(new_net_2125),
		.c(_0750_)
	);

	or_bb _3461_ (
		.a(new_net_3856),
		.b(new_net_576),
		.c(_0751_)
	);

	and_ii _3462_ (
		.a(new_net_898),
		.b(new_net_412),
		.c(_0752_)
	);

	and_bb _3463_ (
		.a(new_net_899),
		.b(new_net_413),
		.c(_0754_)
	);

	or_bb _3464_ (
		.a(new_net_3857),
		.b(new_net_1090),
		.c(_0755_)
	);

	and_ii _3465_ (
		.a(new_net_1670),
		.b(new_net_362),
		.c(_0756_)
	);

	and_bb _3466_ (
		.a(new_net_1671),
		.b(new_net_363),
		.c(_0757_)
	);

	or_bb _3467_ (
		.a(new_net_3858),
		.b(new_net_1050),
		.c(_0758_)
	);

	and_ii _3468_ (
		.a(new_net_2226),
		.b(new_net_1362),
		.c(_0759_)
	);

	and_bb _3469_ (
		.a(new_net_2227),
		.b(new_net_1363),
		.c(_0760_)
	);

	and_ii _3470_ (
		.a(new_net_3859),
		.b(new_net_2440),
		.c(_0761_)
	);

	and_bb _3471_ (
		.a(new_net_2823),
		.b(new_net_307),
		.c(_0762_)
	);

	and_ii _3472_ (
		.a(new_net_2824),
		.b(new_net_308),
		.c(_0763_)
	);

	or_bb _3473_ (
		.a(new_net_3860),
		.b(new_net_3055),
		.c(new_net_3918)
	);

	or_bb _3474_ (
		.a(new_net_3056),
		.b(new_net_2441),
		.c(_0765_)
	);

	and_ii _3475_ (
		.a(new_net_1051),
		.b(new_net_1091),
		.c(_0766_)
	);

	and_bb _3476_ (
		.a(new_net_924),
		.b(new_net_389),
		.c(_0767_)
	);

	and_ii _3477_ (
		.a(new_net_577),
		.b(new_net_9),
		.c(_0768_)
	);

	and_bb _3478_ (
		.a(new_net_2505),
		.b(new_net_537),
		.c(_0769_)
	);

	and_ii _3479_ (
		.a(new_net_595),
		.b(new_net_1821),
		.c(_0770_)
	);

	and_bb _3480_ (
		.a(new_net_1121),
		.b(new_net_160),
		.c(_0771_)
	);

	and_ii _3481_ (
		.a(new_net_314),
		.b(new_net_780),
		.c(_0772_)
	);

	and_bb _3482_ (
		.a(new_net_1554),
		.b(new_net_440),
		.c(_0773_)
	);

	and_ii _3483_ (
		.a(new_net_63),
		.b(new_net_1526),
		.c(_0775_)
	);

	and_bb _3484_ (
		.a(new_net_2711),
		.b(new_net_3022),
		.c(_0776_)
	);

	and_ii _3485_ (
		.a(new_net_253),
		.b(new_net_1209),
		.c(_0777_)
	);

	and_bb _3486_ (
		.a(new_net_2048),
		.b(new_net_2620),
		.c(_0778_)
	);

	and_bb _3487_ (
		.a(new_net_2866),
		.b(new_net_272),
		.c(_0779_)
	);

	and_ii _3488_ (
		.a(new_net_2129),
		.b(new_net_1015),
		.c(_0780_)
	);

	and_ii _3489_ (
		.a(new_net_370),
		.b(new_net_2472),
		.c(_0781_)
	);

	and_bb _3490_ (
		.a(new_net_371),
		.b(new_net_2473),
		.c(_0782_)
	);

	or_bb _3491_ (
		.a(new_net_3861),
		.b(new_net_416),
		.c(_0783_)
	);

	and_ii _3492_ (
		.a(new_net_52),
		.b(new_net_315),
		.c(_0784_)
	);

	and_bb _3493_ (
		.a(new_net_53),
		.b(new_net_316),
		.c(_0786_)
	);

	or_bb _3494_ (
		.a(new_net_3862),
		.b(new_net_554),
		.c(_0787_)
	);

	and_ii _3495_ (
		.a(new_net_840),
		.b(new_net_2082),
		.c(_0788_)
	);

	and_bb _3496_ (
		.a(new_net_841),
		.b(new_net_2083),
		.c(_0789_)
	);

	or_bb _3497_ (
		.a(new_net_3863),
		.b(new_net_695),
		.c(_0790_)
	);

	and_ii _3498_ (
		.a(new_net_2571),
		.b(new_net_1888),
		.c(_0791_)
	);

	and_bb _3499_ (
		.a(new_net_2572),
		.b(new_net_1889),
		.c(_0792_)
	);

	or_bb _3500_ (
		.a(new_net_3864),
		.b(new_net_850),
		.c(_0793_)
	);

	and_ii _3501_ (
		.a(new_net_904),
		.b(new_net_1712),
		.c(_0794_)
	);

	and_bb _3502_ (
		.a(new_net_905),
		.b(new_net_1713),
		.c(_0795_)
	);

	or_bb _3503_ (
		.a(new_net_3865),
		.b(new_net_2090),
		.c(_0797_)
	);

	and_ii _3504_ (
		.a(new_net_2685),
		.b(new_net_1330),
		.c(_0798_)
	);

	and_bb _3505_ (
		.a(new_net_2686),
		.b(new_net_1331),
		.c(_0799_)
	);

	or_bb _3506_ (
		.a(new_net_3866),
		.b(new_net_2886),
		.c(_0800_)
	);

	and_ii _3507_ (
		.a(new_net_1102),
		.b(new_net_1136),
		.c(_0801_)
	);

	and_bb _3508_ (
		.a(new_net_1103),
		.b(new_net_1137),
		.c(_0802_)
	);

	or_bb _3509_ (
		.a(new_net_3867),
		.b(new_net_1142),
		.c(_0803_)
	);

	and_ii _3510_ (
		.a(new_net_1216),
		.b(new_net_984),
		.c(_0804_)
	);

	and_bb _3511_ (
		.a(new_net_1217),
		.b(new_net_985),
		.c(_0805_)
	);

	or_bb _3512_ (
		.a(new_net_3868),
		.b(new_net_858),
		.c(_0806_)
	);

	and_ii _3513_ (
		.a(new_net_1160),
		.b(new_net_834),
		.c(_0808_)
	);

	and_bb _3514_ (
		.a(new_net_1161),
		.b(new_net_835),
		.c(_0809_)
	);

	or_bb _3515_ (
		.a(new_net_3869),
		.b(new_net_1588),
		.c(_0810_)
	);

	and_ii _3516_ (
		.a(new_net_1537),
		.b(new_net_1096),
		.c(_0811_)
	);

	and_bb _3517_ (
		.a(new_net_1538),
		.b(new_net_1097),
		.c(_0812_)
	);

	or_bb _3518_ (
		.a(new_net_3870),
		.b(new_net_2100),
		.c(_0813_)
	);

	and_ii _3519_ (
		.a(new_net_1642),
		.b(new_net_1529),
		.c(_0814_)
	);

	and_bb _3520_ (
		.a(new_net_1643),
		.b(new_net_1530),
		.c(_0815_)
	);

	or_bb _3521_ (
		.a(new_net_3871),
		.b(new_net_1676),
		.c(_0816_)
	);

	and_ii _3522_ (
		.a(new_net_1956),
		.b(new_net_797),
		.c(_0817_)
	);

	and_bb _3523_ (
		.a(new_net_1957),
		.b(new_net_798),
		.c(_0819_)
	);

	or_bb _3524_ (
		.a(new_net_3872),
		.b(new_net_2168),
		.c(_0820_)
	);

	and_ii _3525_ (
		.a(new_net_1882),
		.b(new_net_1423),
		.c(_0821_)
	);

	and_bb _3526_ (
		.a(new_net_1883),
		.b(new_net_1424),
		.c(_0822_)
	);

	and_ii _3527_ (
		.a(new_net_3873),
		.b(new_net_2977),
		.c(_0823_)
	);

	and_bb _3528_ (
		.a(new_net_1976),
		.b(new_net_1380),
		.c(_0824_)
	);

	and_ii _3529_ (
		.a(new_net_1977),
		.b(new_net_1381),
		.c(_0825_)
	);

	or_bb _3530_ (
		.a(new_net_3874),
		.b(new_net_2010),
		.c(new_net_3946)
	);

	or_bb _3531_ (
		.a(new_net_2011),
		.b(new_net_2978),
		.c(_0826_)
	);

	and_ii _3532_ (
		.a(new_net_2169),
		.b(new_net_1677),
		.c(_0827_)
	);

	and_bb _3533_ (
		.a(new_net_2497),
		.b(new_net_919),
		.c(_0829_)
	);

	and_ii _3534_ (
		.a(new_net_2101),
		.b(new_net_1589),
		.c(_0830_)
	);

	and_bb _3535_ (
		.a(new_net_1131),
		.b(new_net_534),
		.c(_0831_)
	);

	and_ii _3536_ (
		.a(new_net_859),
		.b(new_net_1143),
		.c(_0832_)
	);

	and_bb _3537_ (
		.a(new_net_1556),
		.b(new_net_155),
		.c(_0833_)
	);

	and_ii _3538_ (
		.a(new_net_2887),
		.b(new_net_2091),
		.c(_0834_)
	);

	and_bb _3539_ (
		.a(new_net_2699),
		.b(new_net_441),
		.c(_0835_)
	);

	and_ii _3540_ (
		.a(new_net_851),
		.b(new_net_696),
		.c(_0836_)
	);

	and_bb _3541_ (
		.a(new_net_2049),
		.b(new_net_3017),
		.c(_0837_)
	);

	and_bb _3542_ (
		.a(new_net_2874),
		.b(new_net_2613),
		.c(_0838_)
	);

	and_ii _3543_ (
		.a(new_net_555),
		.b(new_net_417),
		.c(_0840_)
	);

	and_ii _3544_ (
		.a(new_net_2671),
		.b(new_net_2593),
		.c(_0841_)
	);

	and_bb _3545_ (
		.a(new_net_2672),
		.b(new_net_2594),
		.c(_0842_)
	);

	or_bb _3546_ (
		.a(new_net_3875),
		.b(new_net_2724),
		.c(_0843_)
	);

	and_ii _3547_ (
		.a(new_net_715),
		.b(new_net_2535),
		.c(_0844_)
	);

	and_bb _3548_ (
		.a(new_net_716),
		.b(new_net_2536),
		.c(_0845_)
	);

	or_bb _3549_ (
		.a(new_net_3876),
		.b(new_net_910),
		.c(_0846_)
	);

	and_ii _3550_ (
		.a(new_net_1224),
		.b(new_net_2488),
		.c(_0847_)
	);

	and_bb _3551_ (
		.a(new_net_1225),
		.b(new_net_2489),
		.c(_0848_)
	);

	or_bb _3552_ (
		.a(new_net_3877),
		.b(new_net_1433),
		.c(_0849_)
	);

	and_ii _3553_ (
		.a(new_net_3053),
		.b(new_net_2376),
		.c(_0851_)
	);

	and_bb _3554_ (
		.a(new_net_3054),
		.b(new_net_2377),
		.c(_0852_)
	);

	or_bb _3555_ (
		.a(new_net_3878),
		.b(new_net_2176),
		.c(_0853_)
	);

	and_ii _3556_ (
		.a(new_net_2579),
		.b(new_net_2434),
		.c(_0854_)
	);

	and_bb _3557_ (
		.a(new_net_2580),
		.b(new_net_2435),
		.c(_0855_)
	);

	or_bb _3558_ (
		.a(new_net_3879),
		.b(new_net_1565),
		.c(_0856_)
	);

	and_ii _3559_ (
		.a(new_net_1694),
		.b(new_net_2392),
		.c(_0857_)
	);

	and_bb _3560_ (
		.a(new_net_1695),
		.b(new_net_2393),
		.c(_0858_)
	);

	or_bb _3561_ (
		.a(new_net_3880),
		.b(new_net_2080),
		.c(_0859_)
	);

	and_ii _3562_ (
		.a(new_net_1756),
		.b(new_net_1766),
		.c(_0860_)
	);

	and_bb _3563_ (
		.a(new_net_1757),
		.b(new_net_1767),
		.c(_0862_)
	);

	or_bb _3564_ (
		.a(new_net_3881),
		.b(new_net_1794),
		.c(_0863_)
	);

	and_ii _3565_ (
		.a(new_net_1910),
		.b(new_net_2294),
		.c(_0864_)
	);

	and_bb _3566_ (
		.a(new_net_1911),
		.b(new_net_2295),
		.c(_0865_)
	);

	or_bb _3567_ (
		.a(new_net_3882),
		.b(new_net_224),
		.c(_0866_)
	);

	and_ii _3568_ (
		.a(new_net_2016),
		.b(new_net_1398),
		.c(_0867_)
	);

	and_bb _3569_ (
		.a(new_net_2017),
		.b(new_net_1399),
		.c(_0868_)
	);

	or_bb _3570_ (
		.a(new_net_3883),
		.b(new_net_2062),
		.c(_0869_)
	);

	and_ii _3571_ (
		.a(new_net_1138),
		.b(new_net_2232),
		.c(_0870_)
	);

	and_bb _3572_ (
		.a(new_net_1139),
		.b(new_net_2233),
		.c(_0871_)
	);

	or_bb _3573_ (
		.a(new_net_3884),
		.b(new_net_2198),
		.c(_0873_)
	);

	and_ii _3574_ (
		.a(new_net_2300),
		.b(new_net_2152),
		.c(_0874_)
	);

	and_bb _3575_ (
		.a(new_net_2301),
		.b(new_net_2153),
		.c(_0875_)
	);

	and_ii _3576_ (
		.a(new_net_3885),
		.b(new_net_2086),
		.c(_0876_)
	);

	and_bb _3577_ (
		.a(new_net_2428),
		.b(new_net_689),
		.c(_0877_)
	);

	and_ii _3578_ (
		.a(new_net_2429),
		.b(new_net_690),
		.c(_0878_)
	);

	or_bb _3579_ (
		.a(new_net_3886),
		.b(new_net_2683),
		.c(new_net_3964)
	);

	or_bb _3580_ (
		.a(new_net_2684),
		.b(new_net_2087),
		.c(_0879_)
	);

	and_ii _3581_ (
		.a(new_net_2199),
		.b(new_net_2063),
		.c(_0880_)
	);

	and_bb _3582_ (
		.a(new_net_1128),
		.b(new_net_920),
		.c(_0881_)
	);

	and_ii _3583_ (
		.a(new_net_225),
		.b(new_net_1795),
		.c(_0883_)
	);

	and_bb _3584_ (
		.a(new_net_1560),
		.b(new_net_530),
		.c(_0884_)
	);

	and_ii _3585_ (
		.a(new_net_2081),
		.b(new_net_1566),
		.c(_0885_)
	);

	and_bb _3586_ (
		.a(new_net_2704),
		.b(new_net_161),
		.c(_0886_)
	);

	and_ii _3587_ (
		.a(new_net_2177),
		.b(new_net_1434),
		.c(_0887_)
	);

	and_bb _3588_ (
		.a(new_net_2044),
		.b(new_net_439),
		.c(_0888_)
	);

	and_bb _3589_ (
		.a(new_net_2876),
		.b(new_net_3026),
		.c(_0889_)
	);

	and_ii _3590_ (
		.a(new_net_911),
		.b(new_net_2725),
		.c(_0890_)
	);

	and_ii _3591_ (
		.a(new_net_2997),
		.b(new_net_1714),
		.c(_0891_)
	);

	and_bb _3592_ (
		.a(new_net_2998),
		.b(new_net_1715),
		.c(_0892_)
	);

	or_bb _3593_ (
		.a(new_net_3887),
		.b(new_net_2094),
		.c(_0894_)
	);

	and_ii _3594_ (
		.a(new_net_2687),
		.b(new_net_1582),
		.c(_0895_)
	);

	and_bb _3595_ (
		.a(new_net_2688),
		.b(new_net_1583),
		.c(_0896_)
	);

	or_bb _3596_ (
		.a(new_net_3888),
		.b(new_net_3260),
		.c(_0897_)
	);

	and_ii _3597_ (
		.a(new_net_1497),
		.b(new_net_1348),
		.c(_0898_)
	);

	and_bb _3598_ (
		.a(new_net_1498),
		.b(new_net_1349),
		.c(_0899_)
	);

	or_bb _3599_ (
		.a(new_net_3889),
		.b(new_net_100),
		.c(_0900_)
	);

	and_ii _3600_ (
		.a(new_net_1996),
		.b(new_net_2813),
		.c(_0901_)
	);

	and_bb _3601_ (
		.a(new_net_1997),
		.b(new_net_2814),
		.c(_0902_)
	);

	or_bb _3602_ (
		.a(new_net_3890),
		.b(new_net_198),
		.c(_0903_)
	);

	and_ii _3603_ (
		.a(new_net_283),
		.b(new_net_2779),
		.c(_0905_)
	);

	and_bb _3604_ (
		.a(new_net_284),
		.b(new_net_2780),
		.c(_0906_)
	);

	or_bb _3605_ (
		.a(new_net_3891),
		.b(new_net_333),
		.c(_0907_)
	);

	and_ii _3606_ (
		.a(new_net_414),
		.b(new_net_2750),
		.c(_0908_)
	);

	and_bb _3607_ (
		.a(new_net_415),
		.b(new_net_2751),
		.c(_0909_)
	);

	or_bb _3608_ (
		.a(new_net_3892),
		.b(new_net_468),
		.c(_0910_)
	);

	and_ii _3609_ (
		.a(new_net_775),
		.b(new_net_2722),
		.c(_0911_)
	);

	and_bb _3610_ (
		.a(new_net_776),
		.b(new_net_2723),
		.c(_0912_)
	);

	or_bb _3611_ (
		.a(new_net_3893),
		.b(new_net_948),
		.c(_0913_)
	);

	and_ii _3612_ (
		.a(new_net_659),
		.b(new_net_2643),
		.c(_0914_)
	);

	and_bb _3613_ (
		.a(new_net_660),
		.b(new_net_2644),
		.c(_0916_)
	);

	or_bb _3614_ (
		.a(new_net_3894),
		.b(new_net_1503),
		.c(_0917_)
	);

	and_ii _3615_ (
		.a(new_net_2002),
		.b(new_net_2591),
		.c(_0918_)
	);

	and_bb _3616_ (
		.a(new_net_2003),
		.b(new_net_2592),
		.c(_0919_)
	);

	and_ii _3617_ (
		.a(new_net_3895),
		.b(new_net_2222),
		.c(_0920_)
	);

	and_bb _3618_ (
		.a(new_net_2633),
		.b(new_net_3127),
		.c(_0921_)
	);

	and_ii _3619_ (
		.a(new_net_2634),
		.b(new_net_3128),
		.c(_0922_)
	);

	or_bb _3620_ (
		.a(new_net_3896),
		.b(new_net_2797),
		.c(new_net_3924)
	);

	or_bb _3621_ (
		.a(new_net_2798),
		.b(new_net_2223),
		.c(_0923_)
	);

	and_ii _3622_ (
		.a(new_net_1504),
		.b(new_net_949),
		.c(_0924_)
	);

	and_bb _3623_ (
		.a(new_net_1551),
		.b(new_net_926),
		.c(_0926_)
	);

	and_ii _3624_ (
		.a(new_net_469),
		.b(new_net_334),
		.c(_0927_)
	);

	and_bb _3625_ (
		.a(new_net_2705),
		.b(new_net_540),
		.c(_0928_)
	);

	and_ii _3626_ (
		.a(new_net_199),
		.b(new_net_101),
		.c(_0929_)
	);

	and_bb _3627_ (
		.a(new_net_2057),
		.b(new_net_156),
		.c(_0930_)
	);

	and_bb _3628_ (
		.a(new_net_2867),
		.b(new_net_435),
		.c(_0931_)
	);

	and_ii _3629_ (
		.a(new_net_3261),
		.b(new_net_2095),
		.c(_0932_)
	);

	and_ii _3630_ (
		.a(new_net_1666),
		.b(new_net_1507),
		.c(_0933_)
	);

	and_bb _3631_ (
		.a(new_net_1667),
		.b(new_net_1508),
		.c(_0934_)
	);

	or_bb _3632_ (
		.a(new_net_3897),
		.b(new_net_1826),
		.c(_0935_)
	);

	and_ii _3633_ (
		.a(new_net_1489),
		.b(new_net_1291),
		.c(_0937_)
	);

	and_bb _3634_ (
		.a(new_net_1490),
		.b(new_net_1292),
		.c(_0938_)
	);

	or_bb _3635_ (
		.a(new_net_3898),
		.b(new_net_2470),
		.c(_0939_)
	);

	and_ii _3636_ (
		.a(new_net_1772),
		.b(new_net_1210),
		.c(_0940_)
	);

	and_bb _3637_ (
		.a(new_net_1773),
		.b(new_net_1211),
		.c(_0941_)
	);

	or_bb _3638_ (
		.a(new_net_3899),
		.b(new_net_1968),
		.c(_0942_)
	);

	and_ii _3639_ (
		.a(new_net_2382),
		.b(new_net_1176),
		.c(_0943_)
	);

	and_bb _3640_ (
		.a(new_net_2383),
		.b(new_net_1177),
		.c(_0944_)
	);

	or_bb _3641_ (
		.a(new_net_3900),
		.b(new_net_2581),
		.c(_0945_)
	);

	and_ii _3642_ (
		.a(new_net_2991),
		.b(new_net_783),
		.c(_0946_)
	);

	and_bb _3643_ (
		.a(new_net_2992),
		.b(new_net_784),
		.c(_0948_)
	);

	or_bb _3644_ (
		.a(new_net_3901),
		.b(new_net_3228),
		.c(_0949_)
	);

	and_ii _3645_ (
		.a(new_net_518),
		.b(new_net_1114),
		.c(_0950_)
	);

	and_bb _3646_ (
		.a(new_net_519),
		.b(new_net_1115),
		.c(_0951_)
	);

	or_bb _3647_ (
		.a(new_net_3902),
		.b(new_net_725),
		.c(_0952_)
	);

	and_ii _3648_ (
		.a(new_net_2116),
		.b(new_net_1048),
		.c(_0953_)
	);

	and_bb _3649_ (
		.a(new_net_2117),
		.b(new_net_1049),
		.c(_0954_)
	);

	and_ii _3650_ (
		.a(new_net_3903),
		.b(new_net_1237),
		.c(_0955_)
	);

	and_bb _3651_ (
		.a(new_net_1640),
		.b(new_net_6),
		.c(_0956_)
	);

	and_ii _3652_ (
		.a(new_net_1641),
		.b(new_net_7),
		.c(_0957_)
	);

	or_bb _3653_ (
		.a(new_net_3904),
		.b(new_net_1776),
		.c(new_net_3948)
	);

	and_ii _3654_ (
		.a(new_net_1777),
		.b(new_net_1238),
		.c(_0959_)
	);

	and_ii _3655_ (
		.a(new_net_726),
		.b(new_net_3229),
		.c(_0960_)
	);

	and_bb _3656_ (
		.a(new_net_2700),
		.b(new_net_927),
		.c(_0961_)
	);

	and_ii _3657_ (
		.a(new_net_2582),
		.b(new_net_1969),
		.c(_0962_)
	);

	and_bb _3658_ (
		.a(new_net_2050),
		.b(new_net_538),
		.c(_0963_)
	);

	and_bb _3659_ (
		.a(new_net_2868),
		.b(new_net_158),
		.c(_0964_)
	);

	and_ii _3660_ (
		.a(new_net_2471),
		.b(new_net_1827),
		.c(_0965_)
	);

	and_ii _3661_ (
		.a(new_net_2647),
		.b(new_net_2585),
		.c(_0966_)
	);

	and_bb _3662_ (
		.a(new_net_2648),
		.b(new_net_2586),
		.c(_0967_)
	);

	or_bb _3663_ (
		.a(new_net_3905),
		.b(new_net_2681),
		.c(_0969_)
	);

	and_ii _3664_ (
		.a(new_net_1066),
		.b(new_net_3266),
		.c(_0970_)
	);

	and_bb _3665_ (
		.a(new_net_1067),
		.b(new_net_3267),
		.c(_0971_)
	);

	or_bb _3666_ (
		.a(new_net_3906),
		.b(new_net_1243),
		.c(_0972_)
	);

	and_ii _3667_ (
		.a(new_net_2925),
		.b(new_net_3007),
		.c(_0973_)
	);

	and_bb _3668_ (
		.a(new_net_2926),
		.b(new_net_3008),
		.c(_0974_)
	);

	or_bb _3669_ (
		.a(new_net_3907),
		.b(new_net_2961),
		.c(_0975_)
	);

	and_ii _3670_ (
		.a(new_net_2204),
		.b(new_net_2785),
		.c(_0976_)
	);

	and_bb _3671_ (
		.a(new_net_2205),
		.b(new_net_2786),
		.c(_0977_)
	);

	or_bb _3672_ (
		.a(new_net_3908),
		.b(new_net_2416),
		.c(_0978_)
	);

	and_ii _3673_ (
		.a(new_net_2789),
		.b(new_net_2601),
		.c(_0980_)
	);

	and_bb _3674_ (
		.a(new_net_2790),
		.b(new_net_2602),
		.c(_0981_)
	);

	and_ii _3675_ (
		.a(new_net_3909),
		.b(new_net_564),
		.c(_0982_)
	);

	and_bi _3676_ (
		.a(new_net_1680),
		.b(new_net_2414),
		.c(_0983_)
	);

	and_bi _3677_ (
		.a(new_net_2415),
		.b(new_net_1681),
		.c(_0984_)
	);

	or_bb _3678_ (
		.a(new_net_3910),
		.b(new_net_1710),
		.c(new_net_3972)
	);

	and_ii _3679_ (
		.a(new_net_1711),
		.b(new_net_565),
		.c(_0985_)
	);

	and_ii _3680_ (
		.a(new_net_2417),
		.b(new_net_2962),
		.c(_0986_)
	);

	and_bb _3681_ (
		.a(new_net_2045),
		.b(new_net_928),
		.c(_0987_)
	);

	and_bb _3682_ (
		.a(new_net_2869),
		.b(new_net_541),
		.c(_0988_)
	);

	and_ii _3683_ (
		.a(new_net_1244),
		.b(new_net_2682),
		.c(_0990_)
	);

	and_ii _3684_ (
		.a(new_net_2422),
		.b(new_net_1998),
		.c(_0991_)
	);

	and_bb _3685_ (
		.a(new_net_2423),
		.b(new_net_1999),
		.c(_0992_)
	);

	or_bb _3686_ (
		.a(new_net_3911),
		.b(new_net_2629),
		.c(_0993_)
	);

	and_ii _3687_ (
		.a(new_net_3035),
		.b(new_net_1816),
		.c(_0994_)
	);

	and_bb _3688_ (
		.a(new_net_3036),
		.b(new_net_1817),
		.c(_0995_)
	);

	or_bb _3689_ (
		.a(new_net_3912),
		.b(new_net_1),
		.c(_0996_)
	);

	and_ii _3690_ (
		.a(new_net_343),
		.b(new_net_1792),
		.c(_0997_)
	);

	and_bb _3691_ (
		.a(new_net_344),
		.b(new_net_1793),
		.c(_0998_)
	);

	and_ii _3692_ (
		.a(new_net_3913),
		.b(new_net_574),
		.c(_0999_)
	);

	and_bi _3693_ (
		.a(new_net_2296),
		.b(new_net_1501),
		.c(_1001_)
	);

	and_bi _3694_ (
		.a(new_net_1502),
		.b(new_net_2297),
		.c(_1002_)
	);

	or_bb _3695_ (
		.a(new_net_3914),
		.b(new_net_1287),
		.c(new_net_3938)
	);

	and_bb _3696_ (
		.a(new_net_2877),
		.b(new_net_921),
		.c(_1003_)
	);

	and_ii _3697_ (
		.a(new_net_2),
		.b(new_net_2630),
		.c(_1004_)
	);

	or_bb _3698_ (
		.a(new_net_1822),
		.b(new_net_1664),
		.c(_1005_)
	);

	and_ii _3699_ (
		.a(new_net_1288),
		.b(new_net_575),
		.c(_1006_)
	);

	and_bb _3700_ (
		.a(new_net_1823),
		.b(new_net_1665),
		.c(_1007_)
	);

	and_bi _3701_ (
		.a(new_net_2563),
		.b(new_net_3915),
		.c(_1008_)
	);

	and_bi _3702_ (
		.a(new_net_2635),
		.b(new_net_2599),
		.c(_1009_)
	);

	and_bi _3703_ (
		.a(new_net_2564),
		.b(new_net_2803),
		.c(N6287)
	);

	and_bi _3704_ (
		.a(new_net_2600),
		.b(new_net_2636),
		.c(_1011_)
	);

	or_bb _3705_ (
		.a(new_net_3916),
		.b(new_net_2804),
		.c(N6288)
	);

	and_bb _3706_ (
		.a(new_net_2469),
		.b(new_net_3168),
		.c(_1012_)
	);

	and_bi _3707_ (
		.a(new_net_2507),
		.b(new_net_3917),
		.c(new_net_3940)
	);

	spl2 _1009__v_fanout (
		.a(_1009_),
		.b(new_net_2803),
		.c(new_net_2804)
	);

	spl2 _1006__v_fanout (
		.a(_1006_),
		.b(new_net_2599),
		.c(new_net_2600)
	);

	spl2 _1001__v_fanout (
		.a(_1001_),
		.b(new_net_1287),
		.c(new_net_1288)
	);

	spl2 _0985__v_fanout (
		.a(_0985_),
		.b(new_net_1501),
		.c(new_net_1502)
	);

	spl2 _0983__v_fanout (
		.a(_0983_),
		.b(new_net_1710),
		.c(new_net_1711)
	);

	spl2 _0959__v_fanout (
		.a(_0959_),
		.b(new_net_2414),
		.c(new_net_2415)
	);

	spl2 _0956__v_fanout (
		.a(_0956_),
		.b(new_net_1776),
		.c(new_net_1777)
	);

	spl2 _0923__v_fanout (
		.a(_0923_),
		.b(new_net_6),
		.c(new_net_7)
	);

	spl2 _0921__v_fanout (
		.a(_0921_),
		.b(new_net_2797),
		.c(new_net_2798)
	);

	spl2 _0879__v_fanout (
		.a(_0879_),
		.b(new_net_3127),
		.c(new_net_3128)
	);

	spl2 _0877__v_fanout (
		.a(_0877_),
		.b(new_net_2683),
		.c(new_net_2684)
	);

	spl2 _0826__v_fanout (
		.a(_0826_),
		.b(new_net_689),
		.c(new_net_690)
	);

	spl2 _0824__v_fanout (
		.a(_0824_),
		.b(new_net_2010),
		.c(new_net_2011)
	);

	spl2 _0765__v_fanout (
		.a(_0765_),
		.b(new_net_1380),
		.c(new_net_1381)
	);

	spl2 _0762__v_fanout (
		.a(_0762_),
		.b(new_net_3055),
		.c(new_net_3056)
	);

	spl2 _0694__v_fanout (
		.a(_0694_),
		.b(new_net_307),
		.c(new_net_308)
	);

	spl2 _0692__v_fanout (
		.a(_0692_),
		.b(new_net_866),
		.c(new_net_867)
	);

	spl2 _0615__v_fanout (
		.a(_0615_),
		.b(new_net_508),
		.c(new_net_509)
	);

	spl2 _0613__v_fanout (
		.a(_0613_),
		.b(new_net_1592),
		.c(new_net_1593)
	);

	spl2 _0527__v_fanout (
		.a(_0527_),
		.b(new_net_2424),
		.c(new_net_2425)
	);

	spl2 _0524__v_fanout (
		.a(_0524_),
		.b(new_net_1828),
		.c(new_net_1829)
	);

	spl2 _0430__v_fanout (
		.a(_0430_),
		.b(new_net_1437),
		.c(new_net_1438)
	);

	spl2 _0428__v_fanout (
		.a(_0428_),
		.b(new_net_1338),
		.c(new_net_1339)
	);

	spl2 _0324__v_fanout (
		.a(_0324_),
		.b(new_net_1382),
		.c(new_net_1383)
	);

	spl2 _0322__v_fanout (
		.a(_0322_),
		.b(new_net_552),
		.c(new_net_553)
	);

	spl2 _0210__v_fanout (
		.a(_0210_),
		.b(new_net_2673),
		.c(new_net_2674)
	);

	spl2 _0207__v_fanout (
		.a(_0207_),
		.b(new_net_669),
		.c(new_net_670)
	);

	spl2 new_net_3454_v_fanout (
		.a(new_net_3454),
		.b(new_net_2506),
		.c(new_net_2508)
	);

	bfr new_net_3976_bfr_after (
		.din(_0955_),
		.dout(new_net_3976)
	);

	bfr new_net_3977_bfr_after (
		.din(new_net_3976),
		.dout(new_net_3977)
	);

	bfr new_net_3978_bfr_after (
		.din(new_net_3977),
		.dout(new_net_3978)
	);

	bfr new_net_3979_bfr_after (
		.din(new_net_3978),
		.dout(new_net_3979)
	);

	bfr new_net_3980_bfr_after (
		.din(new_net_3979),
		.dout(new_net_3980)
	);

	bfr new_net_3981_bfr_after (
		.din(new_net_3980),
		.dout(new_net_3981)
	);

	bfr new_net_3982_bfr_after (
		.din(new_net_3981),
		.dout(new_net_3982)
	);

	bfr new_net_3983_bfr_after (
		.din(new_net_3982),
		.dout(new_net_3983)
	);

	bfr new_net_3984_bfr_after (
		.din(new_net_3983),
		.dout(new_net_3984)
	);

	bfr new_net_3985_bfr_after (
		.din(new_net_3984),
		.dout(new_net_3985)
	);

	bfr new_net_3986_bfr_after (
		.din(new_net_3985),
		.dout(new_net_3986)
	);

	bfr new_net_3987_bfr_after (
		.din(new_net_3986),
		.dout(new_net_3987)
	);

	bfr new_net_3988_bfr_after (
		.din(new_net_3987),
		.dout(new_net_3988)
	);

	bfr new_net_3989_bfr_after (
		.din(new_net_3988),
		.dout(new_net_3989)
	);

	bfr new_net_3990_bfr_after (
		.din(new_net_3989),
		.dout(new_net_3990)
	);

	bfr new_net_3991_bfr_after (
		.din(new_net_3990),
		.dout(new_net_3991)
	);

	bfr new_net_3992_bfr_after (
		.din(new_net_3991),
		.dout(new_net_3992)
	);

	bfr new_net_3993_bfr_after (
		.din(new_net_3992),
		.dout(new_net_3993)
	);

	bfr new_net_3994_bfr_after (
		.din(new_net_3993),
		.dout(new_net_3994)
	);

	bfr new_net_3995_bfr_after (
		.din(new_net_3994),
		.dout(new_net_3995)
	);

	bfr new_net_3996_bfr_after (
		.din(new_net_3995),
		.dout(new_net_3996)
	);

	bfr new_net_3997_bfr_after (
		.din(new_net_3996),
		.dout(new_net_3997)
	);

	bfr new_net_3998_bfr_after (
		.din(new_net_3997),
		.dout(new_net_3998)
	);

	bfr new_net_3999_bfr_after (
		.din(new_net_3998),
		.dout(new_net_3999)
	);

	bfr new_net_4000_bfr_after (
		.din(new_net_3999),
		.dout(new_net_4000)
	);

	bfr new_net_4001_bfr_after (
		.din(new_net_4000),
		.dout(new_net_4001)
	);

	bfr new_net_4002_bfr_after (
		.din(new_net_4001),
		.dout(new_net_4002)
	);

	bfr new_net_4003_bfr_after (
		.din(new_net_4002),
		.dout(new_net_4003)
	);

	bfr new_net_4004_bfr_after (
		.din(new_net_4003),
		.dout(new_net_4004)
	);

	bfr new_net_4005_bfr_after (
		.din(new_net_4004),
		.dout(new_net_4005)
	);

	bfr new_net_4006_bfr_after (
		.din(new_net_4005),
		.dout(new_net_4006)
	);

	bfr new_net_4007_bfr_after (
		.din(new_net_4006),
		.dout(new_net_4007)
	);

	bfr new_net_4008_bfr_after (
		.din(new_net_4007),
		.dout(new_net_4008)
	);

	bfr new_net_4009_bfr_after (
		.din(new_net_4008),
		.dout(new_net_4009)
	);

	bfr new_net_4010_bfr_after (
		.din(new_net_4009),
		.dout(new_net_4010)
	);

	bfr new_net_4011_bfr_after (
		.din(new_net_4010),
		.dout(new_net_4011)
	);

	bfr new_net_4012_bfr_after (
		.din(new_net_4011),
		.dout(new_net_4012)
	);

	bfr new_net_4013_bfr_after (
		.din(new_net_4012),
		.dout(new_net_4013)
	);

	bfr new_net_4014_bfr_after (
		.din(new_net_4013),
		.dout(new_net_4014)
	);

	bfr new_net_4015_bfr_after (
		.din(new_net_4014),
		.dout(new_net_4015)
	);

	spl2 _0955__v_fanout (
		.a(new_net_4015),
		.b(new_net_1640),
		.c(new_net_1641)
	);

	bfr new_net_4016_bfr_after (
		.din(_0982_),
		.dout(new_net_4016)
	);

	bfr new_net_4017_bfr_after (
		.din(new_net_4016),
		.dout(new_net_4017)
	);

	bfr new_net_4018_bfr_after (
		.din(new_net_4017),
		.dout(new_net_4018)
	);

	bfr new_net_4019_bfr_after (
		.din(new_net_4018),
		.dout(new_net_4019)
	);

	bfr new_net_4020_bfr_after (
		.din(new_net_4019),
		.dout(new_net_4020)
	);

	bfr new_net_4021_bfr_after (
		.din(new_net_4020),
		.dout(new_net_4021)
	);

	bfr new_net_4022_bfr_after (
		.din(new_net_4021),
		.dout(new_net_4022)
	);

	bfr new_net_4023_bfr_after (
		.din(new_net_4022),
		.dout(new_net_4023)
	);

	bfr new_net_4024_bfr_after (
		.din(new_net_4023),
		.dout(new_net_4024)
	);

	bfr new_net_4025_bfr_after (
		.din(new_net_4024),
		.dout(new_net_4025)
	);

	bfr new_net_4026_bfr_after (
		.din(new_net_4025),
		.dout(new_net_4026)
	);

	bfr new_net_4027_bfr_after (
		.din(new_net_4026),
		.dout(new_net_4027)
	);

	bfr new_net_4028_bfr_after (
		.din(new_net_4027),
		.dout(new_net_4028)
	);

	bfr new_net_4029_bfr_after (
		.din(new_net_4028),
		.dout(new_net_4029)
	);

	bfr new_net_4030_bfr_after (
		.din(new_net_4029),
		.dout(new_net_4030)
	);

	bfr new_net_4031_bfr_after (
		.din(new_net_4030),
		.dout(new_net_4031)
	);

	bfr new_net_4032_bfr_after (
		.din(new_net_4031),
		.dout(new_net_4032)
	);

	bfr new_net_4033_bfr_after (
		.din(new_net_4032),
		.dout(new_net_4033)
	);

	bfr new_net_4034_bfr_after (
		.din(new_net_4033),
		.dout(new_net_4034)
	);

	bfr new_net_4035_bfr_after (
		.din(new_net_4034),
		.dout(new_net_4035)
	);

	bfr new_net_4036_bfr_after (
		.din(new_net_4035),
		.dout(new_net_4036)
	);

	bfr new_net_4037_bfr_after (
		.din(new_net_4036),
		.dout(new_net_4037)
	);

	bfr new_net_4038_bfr_after (
		.din(new_net_4037),
		.dout(new_net_4038)
	);

	bfr new_net_4039_bfr_after (
		.din(new_net_4038),
		.dout(new_net_4039)
	);

	bfr new_net_4040_bfr_after (
		.din(new_net_4039),
		.dout(new_net_4040)
	);

	bfr new_net_4041_bfr_after (
		.din(new_net_4040),
		.dout(new_net_4041)
	);

	bfr new_net_4042_bfr_after (
		.din(new_net_4041),
		.dout(new_net_4042)
	);

	bfr new_net_4043_bfr_after (
		.din(new_net_4042),
		.dout(new_net_4043)
	);

	bfr new_net_4044_bfr_after (
		.din(new_net_4043),
		.dout(new_net_4044)
	);

	bfr new_net_4045_bfr_after (
		.din(new_net_4044),
		.dout(new_net_4045)
	);

	bfr new_net_4046_bfr_after (
		.din(new_net_4045),
		.dout(new_net_4046)
	);

	bfr new_net_4047_bfr_after (
		.din(new_net_4046),
		.dout(new_net_4047)
	);

	bfr new_net_4048_bfr_after (
		.din(new_net_4047),
		.dout(new_net_4048)
	);

	bfr new_net_4049_bfr_after (
		.din(new_net_4048),
		.dout(new_net_4049)
	);

	bfr new_net_4050_bfr_after (
		.din(new_net_4049),
		.dout(new_net_4050)
	);

	bfr new_net_4051_bfr_after (
		.din(new_net_4050),
		.dout(new_net_4051)
	);

	bfr new_net_4052_bfr_after (
		.din(new_net_4051),
		.dout(new_net_4052)
	);

	bfr new_net_4053_bfr_after (
		.din(new_net_4052),
		.dout(new_net_4053)
	);

	bfr new_net_4054_bfr_after (
		.din(new_net_4053),
		.dout(new_net_4054)
	);

	bfr new_net_4055_bfr_after (
		.din(new_net_4054),
		.dout(new_net_4055)
	);

	bfr new_net_4056_bfr_after (
		.din(new_net_4055),
		.dout(new_net_4056)
	);

	bfr new_net_4057_bfr_after (
		.din(new_net_4056),
		.dout(new_net_4057)
	);

	bfr new_net_4058_bfr_after (
		.din(new_net_4057),
		.dout(new_net_4058)
	);

	bfr new_net_4059_bfr_after (
		.din(new_net_4058),
		.dout(new_net_4059)
	);

	spl2 _0982__v_fanout (
		.a(new_net_4059),
		.b(new_net_1680),
		.c(new_net_1681)
	);

	bfr new_net_4060_bfr_after (
		.din(_0761_),
		.dout(new_net_4060)
	);

	bfr new_net_4061_bfr_after (
		.din(new_net_4060),
		.dout(new_net_4061)
	);

	bfr new_net_4062_bfr_after (
		.din(new_net_4061),
		.dout(new_net_4062)
	);

	bfr new_net_4063_bfr_after (
		.din(new_net_4062),
		.dout(new_net_4063)
	);

	bfr new_net_4064_bfr_after (
		.din(new_net_4063),
		.dout(new_net_4064)
	);

	bfr new_net_4065_bfr_after (
		.din(new_net_4064),
		.dout(new_net_4065)
	);

	bfr new_net_4066_bfr_after (
		.din(new_net_4065),
		.dout(new_net_4066)
	);

	bfr new_net_4067_bfr_after (
		.din(new_net_4066),
		.dout(new_net_4067)
	);

	bfr new_net_4068_bfr_after (
		.din(new_net_4067),
		.dout(new_net_4068)
	);

	bfr new_net_4069_bfr_after (
		.din(new_net_4068),
		.dout(new_net_4069)
	);

	bfr new_net_4070_bfr_after (
		.din(new_net_4069),
		.dout(new_net_4070)
	);

	bfr new_net_4071_bfr_after (
		.din(new_net_4070),
		.dout(new_net_4071)
	);

	bfr new_net_4072_bfr_after (
		.din(new_net_4071),
		.dout(new_net_4072)
	);

	bfr new_net_4073_bfr_after (
		.din(new_net_4072),
		.dout(new_net_4073)
	);

	bfr new_net_4074_bfr_after (
		.din(new_net_4073),
		.dout(new_net_4074)
	);

	bfr new_net_4075_bfr_after (
		.din(new_net_4074),
		.dout(new_net_4075)
	);

	bfr new_net_4076_bfr_after (
		.din(new_net_4075),
		.dout(new_net_4076)
	);

	bfr new_net_4077_bfr_after (
		.din(new_net_4076),
		.dout(new_net_4077)
	);

	bfr new_net_4078_bfr_after (
		.din(new_net_4077),
		.dout(new_net_4078)
	);

	bfr new_net_4079_bfr_after (
		.din(new_net_4078),
		.dout(new_net_4079)
	);

	bfr new_net_4080_bfr_after (
		.din(new_net_4079),
		.dout(new_net_4080)
	);

	bfr new_net_4081_bfr_after (
		.din(new_net_4080),
		.dout(new_net_4081)
	);

	bfr new_net_4082_bfr_after (
		.din(new_net_4081),
		.dout(new_net_4082)
	);

	bfr new_net_4083_bfr_after (
		.din(new_net_4082),
		.dout(new_net_4083)
	);

	spl2 _0761__v_fanout (
		.a(new_net_4083),
		.b(new_net_2823),
		.c(new_net_2824)
	);

	bfr new_net_4084_bfr_after (
		.din(_0876_),
		.dout(new_net_4084)
	);

	bfr new_net_4085_bfr_after (
		.din(new_net_4084),
		.dout(new_net_4085)
	);

	bfr new_net_4086_bfr_after (
		.din(new_net_4085),
		.dout(new_net_4086)
	);

	bfr new_net_4087_bfr_after (
		.din(new_net_4086),
		.dout(new_net_4087)
	);

	bfr new_net_4088_bfr_after (
		.din(new_net_4087),
		.dout(new_net_4088)
	);

	bfr new_net_4089_bfr_after (
		.din(new_net_4088),
		.dout(new_net_4089)
	);

	bfr new_net_4090_bfr_after (
		.din(new_net_4089),
		.dout(new_net_4090)
	);

	bfr new_net_4091_bfr_after (
		.din(new_net_4090),
		.dout(new_net_4091)
	);

	bfr new_net_4092_bfr_after (
		.din(new_net_4091),
		.dout(new_net_4092)
	);

	bfr new_net_4093_bfr_after (
		.din(new_net_4092),
		.dout(new_net_4093)
	);

	bfr new_net_4094_bfr_after (
		.din(new_net_4093),
		.dout(new_net_4094)
	);

	bfr new_net_4095_bfr_after (
		.din(new_net_4094),
		.dout(new_net_4095)
	);

	bfr new_net_4096_bfr_after (
		.din(new_net_4095),
		.dout(new_net_4096)
	);

	bfr new_net_4097_bfr_after (
		.din(new_net_4096),
		.dout(new_net_4097)
	);

	bfr new_net_4098_bfr_after (
		.din(new_net_4097),
		.dout(new_net_4098)
	);

	bfr new_net_4099_bfr_after (
		.din(new_net_4098),
		.dout(new_net_4099)
	);

	bfr new_net_4100_bfr_after (
		.din(new_net_4099),
		.dout(new_net_4100)
	);

	bfr new_net_4101_bfr_after (
		.din(new_net_4100),
		.dout(new_net_4101)
	);

	bfr new_net_4102_bfr_after (
		.din(new_net_4101),
		.dout(new_net_4102)
	);

	bfr new_net_4103_bfr_after (
		.din(new_net_4102),
		.dout(new_net_4103)
	);

	bfr new_net_4104_bfr_after (
		.din(new_net_4103),
		.dout(new_net_4104)
	);

	bfr new_net_4105_bfr_after (
		.din(new_net_4104),
		.dout(new_net_4105)
	);

	bfr new_net_4106_bfr_after (
		.din(new_net_4105),
		.dout(new_net_4106)
	);

	bfr new_net_4107_bfr_after (
		.din(new_net_4106),
		.dout(new_net_4107)
	);

	bfr new_net_4108_bfr_after (
		.din(new_net_4107),
		.dout(new_net_4108)
	);

	bfr new_net_4109_bfr_after (
		.din(new_net_4108),
		.dout(new_net_4109)
	);

	bfr new_net_4110_bfr_after (
		.din(new_net_4109),
		.dout(new_net_4110)
	);

	bfr new_net_4111_bfr_after (
		.din(new_net_4110),
		.dout(new_net_4111)
	);

	bfr new_net_4112_bfr_after (
		.din(new_net_4111),
		.dout(new_net_4112)
	);

	bfr new_net_4113_bfr_after (
		.din(new_net_4112),
		.dout(new_net_4113)
	);

	bfr new_net_4114_bfr_after (
		.din(new_net_4113),
		.dout(new_net_4114)
	);

	bfr new_net_4115_bfr_after (
		.din(new_net_4114),
		.dout(new_net_4115)
	);

	spl2 _0876__v_fanout (
		.a(new_net_4115),
		.b(new_net_2428),
		.c(new_net_2429)
	);

	bfr new_net_4116_bfr_after (
		.din(_0321_),
		.dout(new_net_4116)
	);

	bfr new_net_4117_bfr_after (
		.din(new_net_4116),
		.dout(new_net_4117)
	);

	bfr new_net_4118_bfr_after (
		.din(new_net_4117),
		.dout(new_net_4118)
	);

	bfr new_net_4119_bfr_after (
		.din(new_net_4118),
		.dout(new_net_4119)
	);

	spl2 _0321__v_fanout (
		.a(new_net_4119),
		.b(new_net_502),
		.c(new_net_503)
	);

	bfr new_net_4120_bfr_after (
		.din(_0691_),
		.dout(new_net_4120)
	);

	bfr new_net_4121_bfr_after (
		.din(new_net_4120),
		.dout(new_net_4121)
	);

	bfr new_net_4122_bfr_after (
		.din(new_net_4121),
		.dout(new_net_4122)
	);

	bfr new_net_4123_bfr_after (
		.din(new_net_4122),
		.dout(new_net_4123)
	);

	bfr new_net_4124_bfr_after (
		.din(new_net_4123),
		.dout(new_net_4124)
	);

	bfr new_net_4125_bfr_after (
		.din(new_net_4124),
		.dout(new_net_4125)
	);

	bfr new_net_4126_bfr_after (
		.din(new_net_4125),
		.dout(new_net_4126)
	);

	bfr new_net_4127_bfr_after (
		.din(new_net_4126),
		.dout(new_net_4127)
	);

	bfr new_net_4128_bfr_after (
		.din(new_net_4127),
		.dout(new_net_4128)
	);

	bfr new_net_4129_bfr_after (
		.din(new_net_4128),
		.dout(new_net_4129)
	);

	bfr new_net_4130_bfr_after (
		.din(new_net_4129),
		.dout(new_net_4130)
	);

	bfr new_net_4131_bfr_after (
		.din(new_net_4130),
		.dout(new_net_4131)
	);

	bfr new_net_4132_bfr_after (
		.din(new_net_4131),
		.dout(new_net_4132)
	);

	bfr new_net_4133_bfr_after (
		.din(new_net_4132),
		.dout(new_net_4133)
	);

	bfr new_net_4134_bfr_after (
		.din(new_net_4133),
		.dout(new_net_4134)
	);

	bfr new_net_4135_bfr_after (
		.din(new_net_4134),
		.dout(new_net_4135)
	);

	bfr new_net_4136_bfr_after (
		.din(new_net_4135),
		.dout(new_net_4136)
	);

	bfr new_net_4137_bfr_after (
		.din(new_net_4136),
		.dout(new_net_4137)
	);

	bfr new_net_4138_bfr_after (
		.din(new_net_4137),
		.dout(new_net_4138)
	);

	bfr new_net_4139_bfr_after (
		.din(new_net_4138),
		.dout(new_net_4139)
	);

	spl2 _0691__v_fanout (
		.a(new_net_4139),
		.b(new_net_639),
		.c(new_net_640)
	);

	bfr new_net_4140_bfr_after (
		.din(_0611_),
		.dout(new_net_4140)
	);

	bfr new_net_4141_bfr_after (
		.din(new_net_4140),
		.dout(new_net_4141)
	);

	bfr new_net_4142_bfr_after (
		.din(new_net_4141),
		.dout(new_net_4142)
	);

	bfr new_net_4143_bfr_after (
		.din(new_net_4142),
		.dout(new_net_4143)
	);

	bfr new_net_4144_bfr_after (
		.din(new_net_4143),
		.dout(new_net_4144)
	);

	bfr new_net_4145_bfr_after (
		.din(new_net_4144),
		.dout(new_net_4145)
	);

	bfr new_net_4146_bfr_after (
		.din(new_net_4145),
		.dout(new_net_4146)
	);

	bfr new_net_4147_bfr_after (
		.din(new_net_4146),
		.dout(new_net_4147)
	);

	bfr new_net_4148_bfr_after (
		.din(new_net_4147),
		.dout(new_net_4148)
	);

	bfr new_net_4149_bfr_after (
		.din(new_net_4148),
		.dout(new_net_4149)
	);

	bfr new_net_4150_bfr_after (
		.din(new_net_4149),
		.dout(new_net_4150)
	);

	bfr new_net_4151_bfr_after (
		.din(new_net_4150),
		.dout(new_net_4151)
	);

	bfr new_net_4152_bfr_after (
		.din(new_net_4151),
		.dout(new_net_4152)
	);

	bfr new_net_4153_bfr_after (
		.din(new_net_4152),
		.dout(new_net_4153)
	);

	bfr new_net_4154_bfr_after (
		.din(new_net_4153),
		.dout(new_net_4154)
	);

	bfr new_net_4155_bfr_after (
		.din(new_net_4154),
		.dout(new_net_4155)
	);

	spl2 _0611__v_fanout (
		.a(new_net_4155),
		.b(new_net_341),
		.c(new_net_342)
	);

	bfr new_net_4156_bfr_after (
		.din(_0823_),
		.dout(new_net_4156)
	);

	bfr new_net_4157_bfr_after (
		.din(new_net_4156),
		.dout(new_net_4157)
	);

	bfr new_net_4158_bfr_after (
		.din(new_net_4157),
		.dout(new_net_4158)
	);

	bfr new_net_4159_bfr_after (
		.din(new_net_4158),
		.dout(new_net_4159)
	);

	bfr new_net_4160_bfr_after (
		.din(new_net_4159),
		.dout(new_net_4160)
	);

	bfr new_net_4161_bfr_after (
		.din(new_net_4160),
		.dout(new_net_4161)
	);

	bfr new_net_4162_bfr_after (
		.din(new_net_4161),
		.dout(new_net_4162)
	);

	bfr new_net_4163_bfr_after (
		.din(new_net_4162),
		.dout(new_net_4163)
	);

	bfr new_net_4164_bfr_after (
		.din(new_net_4163),
		.dout(new_net_4164)
	);

	bfr new_net_4165_bfr_after (
		.din(new_net_4164),
		.dout(new_net_4165)
	);

	bfr new_net_4166_bfr_after (
		.din(new_net_4165),
		.dout(new_net_4166)
	);

	bfr new_net_4167_bfr_after (
		.din(new_net_4166),
		.dout(new_net_4167)
	);

	bfr new_net_4168_bfr_after (
		.din(new_net_4167),
		.dout(new_net_4168)
	);

	bfr new_net_4169_bfr_after (
		.din(new_net_4168),
		.dout(new_net_4169)
	);

	bfr new_net_4170_bfr_after (
		.din(new_net_4169),
		.dout(new_net_4170)
	);

	bfr new_net_4171_bfr_after (
		.din(new_net_4170),
		.dout(new_net_4171)
	);

	bfr new_net_4172_bfr_after (
		.din(new_net_4171),
		.dout(new_net_4172)
	);

	bfr new_net_4173_bfr_after (
		.din(new_net_4172),
		.dout(new_net_4173)
	);

	bfr new_net_4174_bfr_after (
		.din(new_net_4173),
		.dout(new_net_4174)
	);

	bfr new_net_4175_bfr_after (
		.din(new_net_4174),
		.dout(new_net_4175)
	);

	bfr new_net_4176_bfr_after (
		.din(new_net_4175),
		.dout(new_net_4176)
	);

	bfr new_net_4177_bfr_after (
		.din(new_net_4176),
		.dout(new_net_4177)
	);

	bfr new_net_4178_bfr_after (
		.din(new_net_4177),
		.dout(new_net_4178)
	);

	bfr new_net_4179_bfr_after (
		.din(new_net_4178),
		.dout(new_net_4179)
	);

	bfr new_net_4180_bfr_after (
		.din(new_net_4179),
		.dout(new_net_4180)
	);

	bfr new_net_4181_bfr_after (
		.din(new_net_4180),
		.dout(new_net_4181)
	);

	bfr new_net_4182_bfr_after (
		.din(new_net_4181),
		.dout(new_net_4182)
	);

	bfr new_net_4183_bfr_after (
		.din(new_net_4182),
		.dout(new_net_4183)
	);

	spl2 _0823__v_fanout (
		.a(new_net_4183),
		.b(new_net_1976),
		.c(new_net_1977)
	);

	bfr new_net_4184_bfr_after (
		.din(_0920_),
		.dout(new_net_4184)
	);

	bfr new_net_4185_bfr_after (
		.din(new_net_4184),
		.dout(new_net_4185)
	);

	bfr new_net_4186_bfr_after (
		.din(new_net_4185),
		.dout(new_net_4186)
	);

	bfr new_net_4187_bfr_after (
		.din(new_net_4186),
		.dout(new_net_4187)
	);

	bfr new_net_4188_bfr_after (
		.din(new_net_4187),
		.dout(new_net_4188)
	);

	bfr new_net_4189_bfr_after (
		.din(new_net_4188),
		.dout(new_net_4189)
	);

	bfr new_net_4190_bfr_after (
		.din(new_net_4189),
		.dout(new_net_4190)
	);

	bfr new_net_4191_bfr_after (
		.din(new_net_4190),
		.dout(new_net_4191)
	);

	bfr new_net_4192_bfr_after (
		.din(new_net_4191),
		.dout(new_net_4192)
	);

	bfr new_net_4193_bfr_after (
		.din(new_net_4192),
		.dout(new_net_4193)
	);

	bfr new_net_4194_bfr_after (
		.din(new_net_4193),
		.dout(new_net_4194)
	);

	bfr new_net_4195_bfr_after (
		.din(new_net_4194),
		.dout(new_net_4195)
	);

	bfr new_net_4196_bfr_after (
		.din(new_net_4195),
		.dout(new_net_4196)
	);

	bfr new_net_4197_bfr_after (
		.din(new_net_4196),
		.dout(new_net_4197)
	);

	bfr new_net_4198_bfr_after (
		.din(new_net_4197),
		.dout(new_net_4198)
	);

	bfr new_net_4199_bfr_after (
		.din(new_net_4198),
		.dout(new_net_4199)
	);

	bfr new_net_4200_bfr_after (
		.din(new_net_4199),
		.dout(new_net_4200)
	);

	bfr new_net_4201_bfr_after (
		.din(new_net_4200),
		.dout(new_net_4201)
	);

	bfr new_net_4202_bfr_after (
		.din(new_net_4201),
		.dout(new_net_4202)
	);

	bfr new_net_4203_bfr_after (
		.din(new_net_4202),
		.dout(new_net_4203)
	);

	bfr new_net_4204_bfr_after (
		.din(new_net_4203),
		.dout(new_net_4204)
	);

	bfr new_net_4205_bfr_after (
		.din(new_net_4204),
		.dout(new_net_4205)
	);

	bfr new_net_4206_bfr_after (
		.din(new_net_4205),
		.dout(new_net_4206)
	);

	bfr new_net_4207_bfr_after (
		.din(new_net_4206),
		.dout(new_net_4207)
	);

	bfr new_net_4208_bfr_after (
		.din(new_net_4207),
		.dout(new_net_4208)
	);

	bfr new_net_4209_bfr_after (
		.din(new_net_4208),
		.dout(new_net_4209)
	);

	bfr new_net_4210_bfr_after (
		.din(new_net_4209),
		.dout(new_net_4210)
	);

	bfr new_net_4211_bfr_after (
		.din(new_net_4210),
		.dout(new_net_4211)
	);

	bfr new_net_4212_bfr_after (
		.din(new_net_4211),
		.dout(new_net_4212)
	);

	bfr new_net_4213_bfr_after (
		.din(new_net_4212),
		.dout(new_net_4213)
	);

	bfr new_net_4214_bfr_after (
		.din(new_net_4213),
		.dout(new_net_4214)
	);

	bfr new_net_4215_bfr_after (
		.din(new_net_4214),
		.dout(new_net_4215)
	);

	bfr new_net_4216_bfr_after (
		.din(new_net_4215),
		.dout(new_net_4216)
	);

	bfr new_net_4217_bfr_after (
		.din(new_net_4216),
		.dout(new_net_4217)
	);

	bfr new_net_4218_bfr_after (
		.din(new_net_4217),
		.dout(new_net_4218)
	);

	bfr new_net_4219_bfr_after (
		.din(new_net_4218),
		.dout(new_net_4219)
	);

	spl2 _0920__v_fanout (
		.a(new_net_4219),
		.b(new_net_2633),
		.c(new_net_2634)
	);

	bfr new_net_4220_bfr_after (
		.din(_0523_),
		.dout(new_net_4220)
	);

	bfr new_net_4221_bfr_after (
		.din(new_net_4220),
		.dout(new_net_4221)
	);

	bfr new_net_4222_bfr_after (
		.din(new_net_4221),
		.dout(new_net_4222)
	);

	bfr new_net_4223_bfr_after (
		.din(new_net_4222),
		.dout(new_net_4223)
	);

	bfr new_net_4224_bfr_after (
		.din(new_net_4223),
		.dout(new_net_4224)
	);

	bfr new_net_4225_bfr_after (
		.din(new_net_4224),
		.dout(new_net_4225)
	);

	bfr new_net_4226_bfr_after (
		.din(new_net_4225),
		.dout(new_net_4226)
	);

	bfr new_net_4227_bfr_after (
		.din(new_net_4226),
		.dout(new_net_4227)
	);

	bfr new_net_4228_bfr_after (
		.din(new_net_4227),
		.dout(new_net_4228)
	);

	bfr new_net_4229_bfr_after (
		.din(new_net_4228),
		.dout(new_net_4229)
	);

	bfr new_net_4230_bfr_after (
		.din(new_net_4229),
		.dout(new_net_4230)
	);

	bfr new_net_4231_bfr_after (
		.din(new_net_4230),
		.dout(new_net_4231)
	);

	spl2 _0523__v_fanout (
		.a(new_net_4231),
		.b(new_net_1668),
		.c(new_net_1669)
	);

	spl2 _0202__v_fanout (
		.a(_0202_),
		.b(new_net_2943),
		.c(new_net_2944)
	);

	bfr new_net_4232_bfr_after (
		.din(_0426_),
		.dout(new_net_4232)
	);

	bfr new_net_4233_bfr_after (
		.din(new_net_4232),
		.dout(new_net_4233)
	);

	bfr new_net_4234_bfr_after (
		.din(new_net_4233),
		.dout(new_net_4234)
	);

	bfr new_net_4235_bfr_after (
		.din(new_net_4234),
		.dout(new_net_4235)
	);

	bfr new_net_4236_bfr_after (
		.din(new_net_4235),
		.dout(new_net_4236)
	);

	bfr new_net_4237_bfr_after (
		.din(new_net_4236),
		.dout(new_net_4237)
	);

	bfr new_net_4238_bfr_after (
		.din(new_net_4237),
		.dout(new_net_4238)
	);

	bfr new_net_4239_bfr_after (
		.din(new_net_4238),
		.dout(new_net_4239)
	);

	spl2 _0426__v_fanout (
		.a(new_net_4239),
		.b(new_net_727),
		.c(new_net_728)
	);

	bfr new_net_4240_bfr_before (
		.din(new_net_4240),
		.dout(new_net_274)
	);

	bfr new_net_4241_bfr_before (
		.din(new_net_4241),
		.dout(new_net_4240)
	);

	bfr new_net_4242_bfr_before (
		.din(new_net_4242),
		.dout(new_net_4241)
	);

	bfr new_net_4243_bfr_before (
		.din(new_net_4243),
		.dout(new_net_4242)
	);

	bfr new_net_4244_bfr_before (
		.din(new_net_4244),
		.dout(new_net_4243)
	);

	bfr new_net_4245_bfr_before (
		.din(new_net_4245),
		.dout(new_net_4244)
	);

	bfr new_net_4246_bfr_before (
		.din(new_net_4246),
		.dout(new_net_4245)
	);

	bfr new_net_4247_bfr_before (
		.din(new_net_4247),
		.dout(new_net_4246)
	);

	bfr new_net_4248_bfr_before (
		.din(new_net_4248),
		.dout(new_net_4247)
	);

	bfr new_net_4249_bfr_before (
		.din(new_net_4249),
		.dout(new_net_4248)
	);

	bfr new_net_4250_bfr_before (
		.din(new_net_4250),
		.dout(new_net_4249)
	);

	bfr new_net_4251_bfr_before (
		.din(new_net_4251),
		.dout(new_net_4250)
	);

	bfr new_net_4252_bfr_before (
		.din(new_net_4252),
		.dout(new_net_4251)
	);

	bfr new_net_4253_bfr_before (
		.din(new_net_4253),
		.dout(new_net_4252)
	);

	bfr new_net_4254_bfr_before (
		.din(new_net_4254),
		.dout(new_net_4253)
	);

	bfr new_net_4255_bfr_before (
		.din(new_net_4255),
		.dout(new_net_4254)
	);

	bfr new_net_4256_bfr_before (
		.din(new_net_4256),
		.dout(new_net_4255)
	);

	bfr new_net_4257_bfr_before (
		.din(new_net_4257),
		.dout(new_net_4256)
	);

	bfr new_net_4258_bfr_before (
		.din(new_net_4258),
		.dout(new_net_4257)
	);

	bfr new_net_4259_bfr_before (
		.din(new_net_4259),
		.dout(new_net_4258)
	);

	spl2 _0609__v_fanout (
		.a(_0609_),
		.b(new_net_273),
		.c(new_net_4259)
	);

	bfr new_net_4260_bfr_before (
		.din(new_net_4260),
		.dout(new_net_3454)
	);

	spl2 _0206__v_fanout (
		.a(_0206_),
		.b(new_net_4260),
		.c(new_net_2507)
	);

	bfr new_net_4261_bfr_before (
		.din(new_net_4261),
		.dout(new_net_565)
	);

	bfr new_net_4262_bfr_before (
		.din(new_net_4262),
		.dout(new_net_4261)
	);

	bfr new_net_4263_bfr_before (
		.din(new_net_4263),
		.dout(new_net_4262)
	);

	bfr new_net_4264_bfr_before (
		.din(new_net_4264),
		.dout(new_net_4263)
	);

	bfr new_net_4265_bfr_before (
		.din(new_net_4265),
		.dout(new_net_4264)
	);

	bfr new_net_4266_bfr_before (
		.din(new_net_4266),
		.dout(new_net_4265)
	);

	bfr new_net_4267_bfr_before (
		.din(new_net_4267),
		.dout(new_net_4266)
	);

	bfr new_net_4268_bfr_before (
		.din(new_net_4268),
		.dout(new_net_4267)
	);

	bfr new_net_4269_bfr_before (
		.din(new_net_4269),
		.dout(new_net_4268)
	);

	bfr new_net_4270_bfr_before (
		.din(new_net_4270),
		.dout(new_net_4269)
	);

	bfr new_net_4271_bfr_before (
		.din(new_net_4271),
		.dout(new_net_4270)
	);

	bfr new_net_4272_bfr_before (
		.din(new_net_4272),
		.dout(new_net_4271)
	);

	bfr new_net_4273_bfr_before (
		.din(new_net_4273),
		.dout(new_net_4272)
	);

	bfr new_net_4274_bfr_before (
		.din(new_net_4274),
		.dout(new_net_4273)
	);

	bfr new_net_4275_bfr_before (
		.din(new_net_4275),
		.dout(new_net_4274)
	);

	bfr new_net_4276_bfr_before (
		.din(new_net_4276),
		.dout(new_net_4275)
	);

	bfr new_net_4277_bfr_before (
		.din(new_net_4277),
		.dout(new_net_4276)
	);

	bfr new_net_4278_bfr_before (
		.din(new_net_4278),
		.dout(new_net_4277)
	);

	bfr new_net_4279_bfr_before (
		.din(new_net_4279),
		.dout(new_net_4278)
	);

	bfr new_net_4280_bfr_before (
		.din(new_net_4280),
		.dout(new_net_4279)
	);

	bfr new_net_4281_bfr_before (
		.din(new_net_4281),
		.dout(new_net_4280)
	);

	bfr new_net_4282_bfr_before (
		.din(new_net_4282),
		.dout(new_net_4281)
	);

	bfr new_net_4283_bfr_before (
		.din(new_net_4283),
		.dout(new_net_4282)
	);

	bfr new_net_4284_bfr_before (
		.din(new_net_4284),
		.dout(new_net_4283)
	);

	bfr new_net_4285_bfr_before (
		.din(new_net_4285),
		.dout(new_net_4284)
	);

	bfr new_net_4286_bfr_before (
		.din(new_net_4286),
		.dout(new_net_4285)
	);

	bfr new_net_4287_bfr_before (
		.din(new_net_4287),
		.dout(new_net_4286)
	);

	bfr new_net_4288_bfr_before (
		.din(new_net_4288),
		.dout(new_net_4287)
	);

	bfr new_net_4289_bfr_before (
		.din(new_net_4289),
		.dout(new_net_4288)
	);

	bfr new_net_4290_bfr_before (
		.din(new_net_4290),
		.dout(new_net_4289)
	);

	bfr new_net_4291_bfr_before (
		.din(new_net_4291),
		.dout(new_net_4290)
	);

	bfr new_net_4292_bfr_before (
		.din(new_net_4292),
		.dout(new_net_4291)
	);

	bfr new_net_4293_bfr_before (
		.din(new_net_4293),
		.dout(new_net_4292)
	);

	bfr new_net_4294_bfr_before (
		.din(new_net_4294),
		.dout(new_net_4293)
	);

	bfr new_net_4295_bfr_before (
		.din(new_net_4295),
		.dout(new_net_4294)
	);

	bfr new_net_4296_bfr_before (
		.din(new_net_4296),
		.dout(new_net_4295)
	);

	bfr new_net_4297_bfr_before (
		.din(new_net_4297),
		.dout(new_net_4296)
	);

	bfr new_net_4298_bfr_before (
		.din(new_net_4298),
		.dout(new_net_4297)
	);

	bfr new_net_4299_bfr_before (
		.din(new_net_4299),
		.dout(new_net_4298)
	);

	bfr new_net_4300_bfr_before (
		.din(new_net_4300),
		.dout(new_net_4299)
	);

	bfr new_net_4301_bfr_before (
		.din(new_net_4301),
		.dout(new_net_4300)
	);

	bfr new_net_4302_bfr_before (
		.din(new_net_4302),
		.dout(new_net_4301)
	);

	bfr new_net_4303_bfr_before (
		.din(new_net_4303),
		.dout(new_net_4302)
	);

	bfr new_net_4304_bfr_before (
		.din(new_net_4304),
		.dout(new_net_4303)
	);

	bfr new_net_4305_bfr_before (
		.din(new_net_4305),
		.dout(new_net_4304)
	);

	bfr new_net_4306_bfr_before (
		.din(new_net_4306),
		.dout(new_net_4305)
	);

	bfr new_net_4307_bfr_before (
		.din(new_net_4307),
		.dout(new_net_4306)
	);

	bfr new_net_4308_bfr_before (
		.din(new_net_4308),
		.dout(new_net_4307)
	);

	spl2 _0980__v_fanout (
		.a(_0980_),
		.b(new_net_564),
		.c(new_net_4308)
	);

	bfr new_net_4309_bfr_before (
		.din(new_net_4309),
		.dout(new_net_2978)
	);

	bfr new_net_4310_bfr_before (
		.din(new_net_4310),
		.dout(new_net_4309)
	);

	bfr new_net_4311_bfr_before (
		.din(new_net_4311),
		.dout(new_net_4310)
	);

	bfr new_net_4312_bfr_before (
		.din(new_net_4312),
		.dout(new_net_4311)
	);

	bfr new_net_4313_bfr_before (
		.din(new_net_4313),
		.dout(new_net_4312)
	);

	bfr new_net_4314_bfr_before (
		.din(new_net_4314),
		.dout(new_net_4313)
	);

	bfr new_net_4315_bfr_before (
		.din(new_net_4315),
		.dout(new_net_4314)
	);

	bfr new_net_4316_bfr_before (
		.din(new_net_4316),
		.dout(new_net_4315)
	);

	bfr new_net_4317_bfr_before (
		.din(new_net_4317),
		.dout(new_net_4316)
	);

	bfr new_net_4318_bfr_before (
		.din(new_net_4318),
		.dout(new_net_4317)
	);

	bfr new_net_4319_bfr_before (
		.din(new_net_4319),
		.dout(new_net_4318)
	);

	bfr new_net_4320_bfr_before (
		.din(new_net_4320),
		.dout(new_net_4319)
	);

	bfr new_net_4321_bfr_before (
		.din(new_net_4321),
		.dout(new_net_4320)
	);

	bfr new_net_4322_bfr_before (
		.din(new_net_4322),
		.dout(new_net_4321)
	);

	bfr new_net_4323_bfr_before (
		.din(new_net_4323),
		.dout(new_net_4322)
	);

	bfr new_net_4324_bfr_before (
		.din(new_net_4324),
		.dout(new_net_4323)
	);

	bfr new_net_4325_bfr_before (
		.din(new_net_4325),
		.dout(new_net_4324)
	);

	bfr new_net_4326_bfr_before (
		.din(new_net_4326),
		.dout(new_net_4325)
	);

	bfr new_net_4327_bfr_before (
		.din(new_net_4327),
		.dout(new_net_4326)
	);

	bfr new_net_4328_bfr_before (
		.din(new_net_4328),
		.dout(new_net_4327)
	);

	bfr new_net_4329_bfr_before (
		.din(new_net_4329),
		.dout(new_net_4328)
	);

	bfr new_net_4330_bfr_before (
		.din(new_net_4330),
		.dout(new_net_4329)
	);

	bfr new_net_4331_bfr_before (
		.din(new_net_4331),
		.dout(new_net_4330)
	);

	bfr new_net_4332_bfr_before (
		.din(new_net_4332),
		.dout(new_net_4331)
	);

	bfr new_net_4333_bfr_before (
		.din(new_net_4333),
		.dout(new_net_4332)
	);

	bfr new_net_4334_bfr_before (
		.din(new_net_4334),
		.dout(new_net_4333)
	);

	bfr new_net_4335_bfr_before (
		.din(new_net_4335),
		.dout(new_net_4334)
	);

	bfr new_net_4336_bfr_before (
		.din(new_net_4336),
		.dout(new_net_4335)
	);

	bfr new_net_4337_bfr_before (
		.din(new_net_4337),
		.dout(new_net_4336)
	);

	bfr new_net_4338_bfr_before (
		.din(new_net_4338),
		.dout(new_net_4337)
	);

	bfr new_net_4339_bfr_before (
		.din(new_net_4339),
		.dout(new_net_4338)
	);

	bfr new_net_4340_bfr_before (
		.din(new_net_4340),
		.dout(new_net_4339)
	);

	spl2 _0821__v_fanout (
		.a(_0821_),
		.b(new_net_2977),
		.c(new_net_4340)
	);

	bfr new_net_4341_bfr_before (
		.din(new_net_4341),
		.dout(new_net_1238)
	);

	bfr new_net_4342_bfr_before (
		.din(new_net_4342),
		.dout(new_net_4341)
	);

	bfr new_net_4343_bfr_before (
		.din(new_net_4343),
		.dout(new_net_4342)
	);

	bfr new_net_4344_bfr_before (
		.din(new_net_4344),
		.dout(new_net_4343)
	);

	bfr new_net_4345_bfr_before (
		.din(new_net_4345),
		.dout(new_net_4344)
	);

	bfr new_net_4346_bfr_before (
		.din(new_net_4346),
		.dout(new_net_4345)
	);

	bfr new_net_4347_bfr_before (
		.din(new_net_4347),
		.dout(new_net_4346)
	);

	bfr new_net_4348_bfr_before (
		.din(new_net_4348),
		.dout(new_net_4347)
	);

	bfr new_net_4349_bfr_before (
		.din(new_net_4349),
		.dout(new_net_4348)
	);

	bfr new_net_4350_bfr_before (
		.din(new_net_4350),
		.dout(new_net_4349)
	);

	bfr new_net_4351_bfr_before (
		.din(new_net_4351),
		.dout(new_net_4350)
	);

	bfr new_net_4352_bfr_before (
		.din(new_net_4352),
		.dout(new_net_4351)
	);

	bfr new_net_4353_bfr_before (
		.din(new_net_4353),
		.dout(new_net_4352)
	);

	bfr new_net_4354_bfr_before (
		.din(new_net_4354),
		.dout(new_net_4353)
	);

	bfr new_net_4355_bfr_before (
		.din(new_net_4355),
		.dout(new_net_4354)
	);

	bfr new_net_4356_bfr_before (
		.din(new_net_4356),
		.dout(new_net_4355)
	);

	bfr new_net_4357_bfr_before (
		.din(new_net_4357),
		.dout(new_net_4356)
	);

	bfr new_net_4358_bfr_before (
		.din(new_net_4358),
		.dout(new_net_4357)
	);

	bfr new_net_4359_bfr_before (
		.din(new_net_4359),
		.dout(new_net_4358)
	);

	bfr new_net_4360_bfr_before (
		.din(new_net_4360),
		.dout(new_net_4359)
	);

	bfr new_net_4361_bfr_before (
		.din(new_net_4361),
		.dout(new_net_4360)
	);

	bfr new_net_4362_bfr_before (
		.din(new_net_4362),
		.dout(new_net_4361)
	);

	bfr new_net_4363_bfr_before (
		.din(new_net_4363),
		.dout(new_net_4362)
	);

	bfr new_net_4364_bfr_before (
		.din(new_net_4364),
		.dout(new_net_4363)
	);

	bfr new_net_4365_bfr_before (
		.din(new_net_4365),
		.dout(new_net_4364)
	);

	bfr new_net_4366_bfr_before (
		.din(new_net_4366),
		.dout(new_net_4365)
	);

	bfr new_net_4367_bfr_before (
		.din(new_net_4367),
		.dout(new_net_4366)
	);

	bfr new_net_4368_bfr_before (
		.din(new_net_4368),
		.dout(new_net_4367)
	);

	bfr new_net_4369_bfr_before (
		.din(new_net_4369),
		.dout(new_net_4368)
	);

	bfr new_net_4370_bfr_before (
		.din(new_net_4370),
		.dout(new_net_4369)
	);

	bfr new_net_4371_bfr_before (
		.din(new_net_4371),
		.dout(new_net_4370)
	);

	bfr new_net_4372_bfr_before (
		.din(new_net_4372),
		.dout(new_net_4371)
	);

	bfr new_net_4373_bfr_before (
		.din(new_net_4373),
		.dout(new_net_4372)
	);

	bfr new_net_4374_bfr_before (
		.din(new_net_4374),
		.dout(new_net_4373)
	);

	bfr new_net_4375_bfr_before (
		.din(new_net_4375),
		.dout(new_net_4374)
	);

	bfr new_net_4376_bfr_before (
		.din(new_net_4376),
		.dout(new_net_4375)
	);

	bfr new_net_4377_bfr_before (
		.din(new_net_4377),
		.dout(new_net_4376)
	);

	bfr new_net_4378_bfr_before (
		.din(new_net_4378),
		.dout(new_net_4377)
	);

	bfr new_net_4379_bfr_before (
		.din(new_net_4379),
		.dout(new_net_4378)
	);

	bfr new_net_4380_bfr_before (
		.din(new_net_4380),
		.dout(new_net_4379)
	);

	bfr new_net_4381_bfr_before (
		.din(new_net_4381),
		.dout(new_net_4380)
	);

	bfr new_net_4382_bfr_before (
		.din(new_net_4382),
		.dout(new_net_4381)
	);

	bfr new_net_4383_bfr_before (
		.din(new_net_4383),
		.dout(new_net_4382)
	);

	bfr new_net_4384_bfr_before (
		.din(new_net_4384),
		.dout(new_net_4383)
	);

	spl2 _0953__v_fanout (
		.a(_0953_),
		.b(new_net_1237),
		.c(new_net_4384)
	);

	bfr new_net_4385_bfr_before (
		.din(new_net_4385),
		.dout(new_net_2267)
	);

	bfr new_net_4386_bfr_before (
		.din(new_net_4386),
		.dout(new_net_4385)
	);

	bfr new_net_4387_bfr_before (
		.din(new_net_4387),
		.dout(new_net_4386)
	);

	bfr new_net_4388_bfr_before (
		.din(new_net_4388),
		.dout(new_net_4387)
	);

	spl2 _0200__v_fanout (
		.a(_0200_),
		.b(new_net_2266),
		.c(new_net_4388)
	);

	bfr new_net_4389_bfr_before (
		.din(new_net_4389),
		.dout(new_net_2087)
	);

	bfr new_net_4390_bfr_before (
		.din(new_net_4390),
		.dout(new_net_4389)
	);

	bfr new_net_4391_bfr_before (
		.din(new_net_4391),
		.dout(new_net_4390)
	);

	bfr new_net_4392_bfr_before (
		.din(new_net_4392),
		.dout(new_net_4391)
	);

	bfr new_net_4393_bfr_before (
		.din(new_net_4393),
		.dout(new_net_4392)
	);

	bfr new_net_4394_bfr_before (
		.din(new_net_4394),
		.dout(new_net_4393)
	);

	bfr new_net_4395_bfr_before (
		.din(new_net_4395),
		.dout(new_net_4394)
	);

	bfr new_net_4396_bfr_before (
		.din(new_net_4396),
		.dout(new_net_4395)
	);

	bfr new_net_4397_bfr_before (
		.din(new_net_4397),
		.dout(new_net_4396)
	);

	bfr new_net_4398_bfr_before (
		.din(new_net_4398),
		.dout(new_net_4397)
	);

	bfr new_net_4399_bfr_before (
		.din(new_net_4399),
		.dout(new_net_4398)
	);

	bfr new_net_4400_bfr_before (
		.din(new_net_4400),
		.dout(new_net_4399)
	);

	bfr new_net_4401_bfr_before (
		.din(new_net_4401),
		.dout(new_net_4400)
	);

	bfr new_net_4402_bfr_before (
		.din(new_net_4402),
		.dout(new_net_4401)
	);

	bfr new_net_4403_bfr_before (
		.din(new_net_4403),
		.dout(new_net_4402)
	);

	bfr new_net_4404_bfr_before (
		.din(new_net_4404),
		.dout(new_net_4403)
	);

	bfr new_net_4405_bfr_before (
		.din(new_net_4405),
		.dout(new_net_4404)
	);

	bfr new_net_4406_bfr_before (
		.din(new_net_4406),
		.dout(new_net_4405)
	);

	bfr new_net_4407_bfr_before (
		.din(new_net_4407),
		.dout(new_net_4406)
	);

	bfr new_net_4408_bfr_before (
		.din(new_net_4408),
		.dout(new_net_4407)
	);

	bfr new_net_4409_bfr_before (
		.din(new_net_4409),
		.dout(new_net_4408)
	);

	bfr new_net_4410_bfr_before (
		.din(new_net_4410),
		.dout(new_net_4409)
	);

	bfr new_net_4411_bfr_before (
		.din(new_net_4411),
		.dout(new_net_4410)
	);

	bfr new_net_4412_bfr_before (
		.din(new_net_4412),
		.dout(new_net_4411)
	);

	bfr new_net_4413_bfr_before (
		.din(new_net_4413),
		.dout(new_net_4412)
	);

	bfr new_net_4414_bfr_before (
		.din(new_net_4414),
		.dout(new_net_4413)
	);

	bfr new_net_4415_bfr_before (
		.din(new_net_4415),
		.dout(new_net_4414)
	);

	bfr new_net_4416_bfr_before (
		.din(new_net_4416),
		.dout(new_net_4415)
	);

	bfr new_net_4417_bfr_before (
		.din(new_net_4417),
		.dout(new_net_4416)
	);

	bfr new_net_4418_bfr_before (
		.din(new_net_4418),
		.dout(new_net_4417)
	);

	bfr new_net_4419_bfr_before (
		.din(new_net_4419),
		.dout(new_net_4418)
	);

	bfr new_net_4420_bfr_before (
		.din(new_net_4420),
		.dout(new_net_4419)
	);

	bfr new_net_4421_bfr_before (
		.din(new_net_4421),
		.dout(new_net_4420)
	);

	bfr new_net_4422_bfr_before (
		.din(new_net_4422),
		.dout(new_net_4421)
	);

	bfr new_net_4423_bfr_before (
		.din(new_net_4423),
		.dout(new_net_4422)
	);

	bfr new_net_4424_bfr_before (
		.din(new_net_4424),
		.dout(new_net_4423)
	);

	spl2 _0874__v_fanout (
		.a(_0874_),
		.b(new_net_2086),
		.c(new_net_4424)
	);

	bfr new_net_4425_bfr_before (
		.din(new_net_4425),
		.dout(new_net_2223)
	);

	bfr new_net_4426_bfr_before (
		.din(new_net_4426),
		.dout(new_net_4425)
	);

	bfr new_net_4427_bfr_before (
		.din(new_net_4427),
		.dout(new_net_4426)
	);

	bfr new_net_4428_bfr_before (
		.din(new_net_4428),
		.dout(new_net_4427)
	);

	bfr new_net_4429_bfr_before (
		.din(new_net_4429),
		.dout(new_net_4428)
	);

	bfr new_net_4430_bfr_before (
		.din(new_net_4430),
		.dout(new_net_4429)
	);

	bfr new_net_4431_bfr_before (
		.din(new_net_4431),
		.dout(new_net_4430)
	);

	bfr new_net_4432_bfr_before (
		.din(new_net_4432),
		.dout(new_net_4431)
	);

	bfr new_net_4433_bfr_before (
		.din(new_net_4433),
		.dout(new_net_4432)
	);

	bfr new_net_4434_bfr_before (
		.din(new_net_4434),
		.dout(new_net_4433)
	);

	bfr new_net_4435_bfr_before (
		.din(new_net_4435),
		.dout(new_net_4434)
	);

	bfr new_net_4436_bfr_before (
		.din(new_net_4436),
		.dout(new_net_4435)
	);

	bfr new_net_4437_bfr_before (
		.din(new_net_4437),
		.dout(new_net_4436)
	);

	bfr new_net_4438_bfr_before (
		.din(new_net_4438),
		.dout(new_net_4437)
	);

	bfr new_net_4439_bfr_before (
		.din(new_net_4439),
		.dout(new_net_4438)
	);

	bfr new_net_4440_bfr_before (
		.din(new_net_4440),
		.dout(new_net_4439)
	);

	bfr new_net_4441_bfr_before (
		.din(new_net_4441),
		.dout(new_net_4440)
	);

	bfr new_net_4442_bfr_before (
		.din(new_net_4442),
		.dout(new_net_4441)
	);

	bfr new_net_4443_bfr_before (
		.din(new_net_4443),
		.dout(new_net_4442)
	);

	bfr new_net_4444_bfr_before (
		.din(new_net_4444),
		.dout(new_net_4443)
	);

	bfr new_net_4445_bfr_before (
		.din(new_net_4445),
		.dout(new_net_4444)
	);

	bfr new_net_4446_bfr_before (
		.din(new_net_4446),
		.dout(new_net_4445)
	);

	bfr new_net_4447_bfr_before (
		.din(new_net_4447),
		.dout(new_net_4446)
	);

	bfr new_net_4448_bfr_before (
		.din(new_net_4448),
		.dout(new_net_4447)
	);

	bfr new_net_4449_bfr_before (
		.din(new_net_4449),
		.dout(new_net_4448)
	);

	bfr new_net_4450_bfr_before (
		.din(new_net_4450),
		.dout(new_net_4449)
	);

	bfr new_net_4451_bfr_before (
		.din(new_net_4451),
		.dout(new_net_4450)
	);

	bfr new_net_4452_bfr_before (
		.din(new_net_4452),
		.dout(new_net_4451)
	);

	bfr new_net_4453_bfr_before (
		.din(new_net_4453),
		.dout(new_net_4452)
	);

	bfr new_net_4454_bfr_before (
		.din(new_net_4454),
		.dout(new_net_4453)
	);

	bfr new_net_4455_bfr_before (
		.din(new_net_4455),
		.dout(new_net_4454)
	);

	bfr new_net_4456_bfr_before (
		.din(new_net_4456),
		.dout(new_net_4455)
	);

	bfr new_net_4457_bfr_before (
		.din(new_net_4457),
		.dout(new_net_4456)
	);

	bfr new_net_4458_bfr_before (
		.din(new_net_4458),
		.dout(new_net_4457)
	);

	bfr new_net_4459_bfr_before (
		.din(new_net_4459),
		.dout(new_net_4458)
	);

	bfr new_net_4460_bfr_before (
		.din(new_net_4460),
		.dout(new_net_4459)
	);

	bfr new_net_4461_bfr_before (
		.din(new_net_4461),
		.dout(new_net_4460)
	);

	bfr new_net_4462_bfr_before (
		.din(new_net_4462),
		.dout(new_net_4461)
	);

	bfr new_net_4463_bfr_before (
		.din(new_net_4463),
		.dout(new_net_4462)
	);

	bfr new_net_4464_bfr_before (
		.din(new_net_4464),
		.dout(new_net_4463)
	);

	spl2 _0918__v_fanout (
		.a(_0918_),
		.b(new_net_2222),
		.c(new_net_4464)
	);

	bfr new_net_4465_bfr_before (
		.din(new_net_4465),
		.dout(new_net_123)
	);

	bfr new_net_4466_bfr_before (
		.din(new_net_4466),
		.dout(new_net_4465)
	);

	bfr new_net_4467_bfr_before (
		.din(new_net_4467),
		.dout(new_net_4466)
	);

	bfr new_net_4468_bfr_before (
		.din(new_net_4468),
		.dout(new_net_4467)
	);

	bfr new_net_4469_bfr_before (
		.din(new_net_4469),
		.dout(new_net_4468)
	);

	bfr new_net_4470_bfr_before (
		.din(new_net_4470),
		.dout(new_net_4469)
	);

	bfr new_net_4471_bfr_before (
		.din(new_net_4471),
		.dout(new_net_4470)
	);

	bfr new_net_4472_bfr_before (
		.din(new_net_4472),
		.dout(new_net_4471)
	);

	bfr new_net_4473_bfr_before (
		.din(new_net_4473),
		.dout(new_net_4472)
	);

	bfr new_net_4474_bfr_before (
		.din(new_net_4474),
		.dout(new_net_4473)
	);

	bfr new_net_4475_bfr_before (
		.din(new_net_4475),
		.dout(new_net_4474)
	);

	bfr new_net_4476_bfr_before (
		.din(new_net_4476),
		.dout(new_net_4475)
	);

	bfr new_net_4477_bfr_before (
		.din(new_net_4477),
		.dout(new_net_4476)
	);

	bfr new_net_4478_bfr_before (
		.din(new_net_4478),
		.dout(new_net_4477)
	);

	bfr new_net_4479_bfr_before (
		.din(new_net_4479),
		.dout(new_net_4478)
	);

	bfr new_net_4480_bfr_before (
		.din(new_net_4480),
		.dout(new_net_4479)
	);

	bfr new_net_4481_bfr_before (
		.din(new_net_4481),
		.dout(new_net_4480)
	);

	bfr new_net_4482_bfr_before (
		.din(new_net_4482),
		.dout(new_net_4481)
	);

	bfr new_net_4483_bfr_before (
		.din(new_net_4483),
		.dout(new_net_4482)
	);

	bfr new_net_4484_bfr_before (
		.din(new_net_4484),
		.dout(new_net_4483)
	);

	bfr new_net_4485_bfr_before (
		.din(new_net_4485),
		.dout(new_net_4484)
	);

	bfr new_net_4486_bfr_before (
		.din(new_net_4486),
		.dout(new_net_4485)
	);

	bfr new_net_4487_bfr_before (
		.din(new_net_4487),
		.dout(new_net_4486)
	);

	bfr new_net_4488_bfr_before (
		.din(new_net_4488),
		.dout(new_net_4487)
	);

	spl2 _0689__v_fanout (
		.a(_0689_),
		.b(new_net_122),
		.c(new_net_4488)
	);

	bfr new_net_4489_bfr_before (
		.din(new_net_4489),
		.dout(new_net_320)
	);

	bfr new_net_4490_bfr_before (
		.din(new_net_4490),
		.dout(new_net_4489)
	);

	bfr new_net_4491_bfr_before (
		.din(new_net_4491),
		.dout(new_net_4490)
	);

	bfr new_net_4492_bfr_before (
		.din(new_net_4492),
		.dout(new_net_4491)
	);

	bfr new_net_4493_bfr_before (
		.din(new_net_4493),
		.dout(new_net_4492)
	);

	bfr new_net_4494_bfr_before (
		.din(new_net_4494),
		.dout(new_net_4493)
	);

	bfr new_net_4495_bfr_before (
		.din(new_net_4495),
		.dout(new_net_4494)
	);

	bfr new_net_4496_bfr_before (
		.din(new_net_4496),
		.dout(new_net_4495)
	);

	bfr new_net_4497_bfr_before (
		.din(new_net_4497),
		.dout(new_net_4496)
	);

	bfr new_net_4498_bfr_before (
		.din(new_net_4498),
		.dout(new_net_4497)
	);

	bfr new_net_4499_bfr_before (
		.din(new_net_4499),
		.dout(new_net_4498)
	);

	bfr new_net_4500_bfr_before (
		.din(new_net_4500),
		.dout(new_net_4499)
	);

	spl2 _0424__v_fanout (
		.a(_0424_),
		.b(new_net_319),
		.c(new_net_4500)
	);

	bfr new_net_4501_bfr_before (
		.din(new_net_4501),
		.dout(new_net_2441)
	);

	bfr new_net_4502_bfr_before (
		.din(new_net_4502),
		.dout(new_net_4501)
	);

	bfr new_net_4503_bfr_before (
		.din(new_net_4503),
		.dout(new_net_4502)
	);

	bfr new_net_4504_bfr_before (
		.din(new_net_4504),
		.dout(new_net_4503)
	);

	bfr new_net_4505_bfr_before (
		.din(new_net_4505),
		.dout(new_net_4504)
	);

	bfr new_net_4506_bfr_before (
		.din(new_net_4506),
		.dout(new_net_4505)
	);

	bfr new_net_4507_bfr_before (
		.din(new_net_4507),
		.dout(new_net_4506)
	);

	bfr new_net_4508_bfr_before (
		.din(new_net_4508),
		.dout(new_net_4507)
	);

	bfr new_net_4509_bfr_before (
		.din(new_net_4509),
		.dout(new_net_4508)
	);

	bfr new_net_4510_bfr_before (
		.din(new_net_4510),
		.dout(new_net_4509)
	);

	bfr new_net_4511_bfr_before (
		.din(new_net_4511),
		.dout(new_net_4510)
	);

	bfr new_net_4512_bfr_before (
		.din(new_net_4512),
		.dout(new_net_4511)
	);

	bfr new_net_4513_bfr_before (
		.din(new_net_4513),
		.dout(new_net_4512)
	);

	bfr new_net_4514_bfr_before (
		.din(new_net_4514),
		.dout(new_net_4513)
	);

	bfr new_net_4515_bfr_before (
		.din(new_net_4515),
		.dout(new_net_4514)
	);

	bfr new_net_4516_bfr_before (
		.din(new_net_4516),
		.dout(new_net_4515)
	);

	bfr new_net_4517_bfr_before (
		.din(new_net_4517),
		.dout(new_net_4516)
	);

	bfr new_net_4518_bfr_before (
		.din(new_net_4518),
		.dout(new_net_4517)
	);

	bfr new_net_4519_bfr_before (
		.din(new_net_4519),
		.dout(new_net_4518)
	);

	bfr new_net_4520_bfr_before (
		.din(new_net_4520),
		.dout(new_net_4519)
	);

	bfr new_net_4521_bfr_before (
		.din(new_net_4521),
		.dout(new_net_4520)
	);

	bfr new_net_4522_bfr_before (
		.din(new_net_4522),
		.dout(new_net_4521)
	);

	bfr new_net_4523_bfr_before (
		.din(new_net_4523),
		.dout(new_net_4522)
	);

	bfr new_net_4524_bfr_before (
		.din(new_net_4524),
		.dout(new_net_4523)
	);

	bfr new_net_4525_bfr_before (
		.din(new_net_4525),
		.dout(new_net_4524)
	);

	bfr new_net_4526_bfr_before (
		.din(new_net_4526),
		.dout(new_net_4525)
	);

	bfr new_net_4527_bfr_before (
		.din(new_net_4527),
		.dout(new_net_4526)
	);

	bfr new_net_4528_bfr_before (
		.din(new_net_4528),
		.dout(new_net_4527)
	);

	spl2 _0759__v_fanout (
		.a(_0759_),
		.b(new_net_2440),
		.c(new_net_4528)
	);

	bfr new_net_4529_bfr_before (
		.din(new_net_4529),
		.dout(new_net_477)
	);

	bfr new_net_4530_bfr_before (
		.din(new_net_4530),
		.dout(new_net_4529)
	);

	bfr new_net_4531_bfr_before (
		.din(new_net_4531),
		.dout(new_net_4530)
	);

	bfr new_net_4532_bfr_before (
		.din(new_net_4532),
		.dout(new_net_4531)
	);

	bfr new_net_4533_bfr_before (
		.din(new_net_4533),
		.dout(new_net_4532)
	);

	bfr new_net_4534_bfr_before (
		.din(new_net_4534),
		.dout(new_net_4533)
	);

	bfr new_net_4535_bfr_before (
		.din(new_net_4535),
		.dout(new_net_4534)
	);

	bfr new_net_4536_bfr_before (
		.din(new_net_4536),
		.dout(new_net_4535)
	);

	spl2 _0319__v_fanout (
		.a(_0319_),
		.b(new_net_476),
		.c(new_net_4536)
	);

	bfr new_net_4537_bfr_before (
		.din(new_net_4537),
		.dout(new_net_1294)
	);

	bfr new_net_4538_bfr_before (
		.din(new_net_4538),
		.dout(new_net_4537)
	);

	bfr new_net_4539_bfr_before (
		.din(new_net_4539),
		.dout(new_net_4538)
	);

	bfr new_net_4540_bfr_before (
		.din(new_net_4540),
		.dout(new_net_4539)
	);

	bfr new_net_4541_bfr_before (
		.din(new_net_4541),
		.dout(new_net_4540)
	);

	bfr new_net_4542_bfr_before (
		.din(new_net_4542),
		.dout(new_net_4541)
	);

	bfr new_net_4543_bfr_before (
		.din(new_net_4543),
		.dout(new_net_4542)
	);

	bfr new_net_4544_bfr_before (
		.din(new_net_4544),
		.dout(new_net_4543)
	);

	bfr new_net_4545_bfr_before (
		.din(new_net_4545),
		.dout(new_net_4544)
	);

	bfr new_net_4546_bfr_before (
		.din(new_net_4546),
		.dout(new_net_4545)
	);

	bfr new_net_4547_bfr_before (
		.din(new_net_4547),
		.dout(new_net_4546)
	);

	bfr new_net_4548_bfr_before (
		.din(new_net_4548),
		.dout(new_net_4547)
	);

	bfr new_net_4549_bfr_before (
		.din(new_net_4549),
		.dout(new_net_4548)
	);

	bfr new_net_4550_bfr_before (
		.din(new_net_4550),
		.dout(new_net_4549)
	);

	bfr new_net_4551_bfr_before (
		.din(new_net_4551),
		.dout(new_net_4550)
	);

	bfr new_net_4552_bfr_before (
		.din(new_net_4552),
		.dout(new_net_4551)
	);

	spl2 _0521__v_fanout (
		.a(_0521_),
		.b(new_net_1293),
		.c(new_net_4552)
	);

	bfr new_net_4553_bfr_after (
		.din(_0999_),
		.dout(new_net_4553)
	);

	bfr new_net_4554_bfr_after (
		.din(new_net_4553),
		.dout(new_net_4554)
	);

	bfr new_net_4555_bfr_after (
		.din(new_net_4554),
		.dout(new_net_4555)
	);

	bfr new_net_4556_bfr_after (
		.din(new_net_4555),
		.dout(new_net_4556)
	);

	bfr new_net_4557_bfr_after (
		.din(new_net_4556),
		.dout(new_net_4557)
	);

	bfr new_net_4558_bfr_after (
		.din(new_net_4557),
		.dout(new_net_4558)
	);

	bfr new_net_4559_bfr_after (
		.din(new_net_4558),
		.dout(new_net_4559)
	);

	bfr new_net_4560_bfr_after (
		.din(new_net_4559),
		.dout(new_net_4560)
	);

	bfr new_net_4561_bfr_after (
		.din(new_net_4560),
		.dout(new_net_4561)
	);

	bfr new_net_4562_bfr_after (
		.din(new_net_4561),
		.dout(new_net_4562)
	);

	bfr new_net_4563_bfr_after (
		.din(new_net_4562),
		.dout(new_net_4563)
	);

	bfr new_net_4564_bfr_after (
		.din(new_net_4563),
		.dout(new_net_4564)
	);

	bfr new_net_4565_bfr_after (
		.din(new_net_4564),
		.dout(new_net_4565)
	);

	bfr new_net_4566_bfr_after (
		.din(new_net_4565),
		.dout(new_net_4566)
	);

	bfr new_net_4567_bfr_after (
		.din(new_net_4566),
		.dout(new_net_4567)
	);

	bfr new_net_4568_bfr_after (
		.din(new_net_4567),
		.dout(new_net_4568)
	);

	bfr new_net_4569_bfr_after (
		.din(new_net_4568),
		.dout(new_net_4569)
	);

	bfr new_net_4570_bfr_after (
		.din(new_net_4569),
		.dout(new_net_4570)
	);

	bfr new_net_4571_bfr_after (
		.din(new_net_4570),
		.dout(new_net_4571)
	);

	bfr new_net_4572_bfr_after (
		.din(new_net_4571),
		.dout(new_net_4572)
	);

	bfr new_net_4573_bfr_after (
		.din(new_net_4572),
		.dout(new_net_4573)
	);

	bfr new_net_4574_bfr_after (
		.din(new_net_4573),
		.dout(new_net_4574)
	);

	bfr new_net_4575_bfr_after (
		.din(new_net_4574),
		.dout(new_net_4575)
	);

	bfr new_net_4576_bfr_after (
		.din(new_net_4575),
		.dout(new_net_4576)
	);

	bfr new_net_4577_bfr_after (
		.din(new_net_4576),
		.dout(new_net_4577)
	);

	bfr new_net_4578_bfr_after (
		.din(new_net_4577),
		.dout(new_net_4578)
	);

	bfr new_net_4579_bfr_after (
		.din(new_net_4578),
		.dout(new_net_4579)
	);

	bfr new_net_4580_bfr_after (
		.din(new_net_4579),
		.dout(new_net_4580)
	);

	bfr new_net_4581_bfr_after (
		.din(new_net_4580),
		.dout(new_net_4581)
	);

	bfr new_net_4582_bfr_after (
		.din(new_net_4581),
		.dout(new_net_4582)
	);

	bfr new_net_4583_bfr_after (
		.din(new_net_4582),
		.dout(new_net_4583)
	);

	bfr new_net_4584_bfr_after (
		.din(new_net_4583),
		.dout(new_net_4584)
	);

	bfr new_net_4585_bfr_after (
		.din(new_net_4584),
		.dout(new_net_4585)
	);

	bfr new_net_4586_bfr_after (
		.din(new_net_4585),
		.dout(new_net_4586)
	);

	bfr new_net_4587_bfr_after (
		.din(new_net_4586),
		.dout(new_net_4587)
	);

	bfr new_net_4588_bfr_after (
		.din(new_net_4587),
		.dout(new_net_4588)
	);

	bfr new_net_4589_bfr_after (
		.din(new_net_4588),
		.dout(new_net_4589)
	);

	bfr new_net_4590_bfr_after (
		.din(new_net_4589),
		.dout(new_net_4590)
	);

	bfr new_net_4591_bfr_after (
		.din(new_net_4590),
		.dout(new_net_4591)
	);

	bfr new_net_4592_bfr_after (
		.din(new_net_4591),
		.dout(new_net_4592)
	);

	bfr new_net_4593_bfr_after (
		.din(new_net_4592),
		.dout(new_net_4593)
	);

	bfr new_net_4594_bfr_after (
		.din(new_net_4593),
		.dout(new_net_4594)
	);

	bfr new_net_4595_bfr_after (
		.din(new_net_4594),
		.dout(new_net_4595)
	);

	bfr new_net_4596_bfr_after (
		.din(new_net_4595),
		.dout(new_net_4596)
	);

	bfr new_net_4597_bfr_after (
		.din(new_net_4596),
		.dout(new_net_4597)
	);

	bfr new_net_4598_bfr_after (
		.din(new_net_4597),
		.dout(new_net_4598)
	);

	bfr new_net_4599_bfr_after (
		.din(new_net_4598),
		.dout(new_net_4599)
	);

	bfr new_net_4600_bfr_after (
		.din(new_net_4599),
		.dout(new_net_4600)
	);

	bfr new_net_4601_bfr_after (
		.din(new_net_4600),
		.dout(new_net_4601)
	);

	bfr new_net_4602_bfr_after (
		.din(new_net_4601),
		.dout(new_net_4602)
	);

	spl2 _0999__v_fanout (
		.a(new_net_4602),
		.b(new_net_2296),
		.c(new_net_2297)
	);

	spl2 _0924__v_fanout (
		.a(_0924_),
		.b(new_net_1048),
		.c(new_net_1049)
	);

	spl2 _0687__v_fanout (
		.a(_0687_),
		.b(new_net_64),
		.c(new_net_65)
	);

	spl2 _0431__v_fanout (
		.a(_0431_),
		.b(new_net_1463),
		.c(new_net_1464)
	);

	spl2 _0317__v_fanout (
		.a(_0317_),
		.b(new_net_92),
		.c(new_net_93)
	);

	spl2 _0880__v_fanout (
		.a(_0880_),
		.b(new_net_2591),
		.c(new_net_2592)
	);

	spl2 _0758__v_fanout (
		.a(_0758_),
		.b(new_net_2226),
		.c(new_net_2227)
	);

	spl2 _0203__v_fanout (
		.a(_0203_),
		.b(new_net_3167),
		.c(new_net_3168)
	);

	spl2 _0873__v_fanout (
		.a(_0873_),
		.b(new_net_2300),
		.c(new_net_2301)
	);

	spl2 _0827__v_fanout (
		.a(_0827_),
		.b(new_net_2152),
		.c(new_net_2153)
	);

	spl2 _0520__v_fanout (
		.a(_0520_),
		.b(new_net_1684),
		.c(new_net_1685)
	);

	spl2 _0616__v_fanout (
		.a(_0616_),
		.b(new_net_562),
		.c(new_net_563)
	);

	spl2 _0960__v_fanout (
		.a(_0960_),
		.b(new_net_2601),
		.c(new_net_2602)
	);

	bfr new_net_4603_bfr_before (
		.din(new_net_4603),
		.dout(new_net_575)
	);

	bfr new_net_4604_bfr_before (
		.din(new_net_4604),
		.dout(new_net_4603)
	);

	bfr new_net_4605_bfr_before (
		.din(new_net_4605),
		.dout(new_net_4604)
	);

	bfr new_net_4606_bfr_before (
		.din(new_net_4606),
		.dout(new_net_4605)
	);

	bfr new_net_4607_bfr_before (
		.din(new_net_4607),
		.dout(new_net_4606)
	);

	bfr new_net_4608_bfr_before (
		.din(new_net_4608),
		.dout(new_net_4607)
	);

	bfr new_net_4609_bfr_before (
		.din(new_net_4609),
		.dout(new_net_4608)
	);

	bfr new_net_4610_bfr_before (
		.din(new_net_4610),
		.dout(new_net_4609)
	);

	bfr new_net_4611_bfr_before (
		.din(new_net_4611),
		.dout(new_net_4610)
	);

	bfr new_net_4612_bfr_before (
		.din(new_net_4612),
		.dout(new_net_4611)
	);

	bfr new_net_4613_bfr_before (
		.din(new_net_4613),
		.dout(new_net_4612)
	);

	bfr new_net_4614_bfr_before (
		.din(new_net_4614),
		.dout(new_net_4613)
	);

	bfr new_net_4615_bfr_before (
		.din(new_net_4615),
		.dout(new_net_4614)
	);

	bfr new_net_4616_bfr_before (
		.din(new_net_4616),
		.dout(new_net_4615)
	);

	bfr new_net_4617_bfr_before (
		.din(new_net_4617),
		.dout(new_net_4616)
	);

	bfr new_net_4618_bfr_before (
		.din(new_net_4618),
		.dout(new_net_4617)
	);

	bfr new_net_4619_bfr_before (
		.din(new_net_4619),
		.dout(new_net_4618)
	);

	bfr new_net_4620_bfr_before (
		.din(new_net_4620),
		.dout(new_net_4619)
	);

	bfr new_net_4621_bfr_before (
		.din(new_net_4621),
		.dout(new_net_4620)
	);

	bfr new_net_4622_bfr_before (
		.din(new_net_4622),
		.dout(new_net_4621)
	);

	bfr new_net_4623_bfr_before (
		.din(new_net_4623),
		.dout(new_net_4622)
	);

	bfr new_net_4624_bfr_before (
		.din(new_net_4624),
		.dout(new_net_4623)
	);

	bfr new_net_4625_bfr_before (
		.din(new_net_4625),
		.dout(new_net_4624)
	);

	bfr new_net_4626_bfr_before (
		.din(new_net_4626),
		.dout(new_net_4625)
	);

	bfr new_net_4627_bfr_before (
		.din(new_net_4627),
		.dout(new_net_4626)
	);

	bfr new_net_4628_bfr_before (
		.din(new_net_4628),
		.dout(new_net_4627)
	);

	bfr new_net_4629_bfr_before (
		.din(new_net_4629),
		.dout(new_net_4628)
	);

	bfr new_net_4630_bfr_before (
		.din(new_net_4630),
		.dout(new_net_4629)
	);

	bfr new_net_4631_bfr_before (
		.din(new_net_4631),
		.dout(new_net_4630)
	);

	bfr new_net_4632_bfr_before (
		.din(new_net_4632),
		.dout(new_net_4631)
	);

	bfr new_net_4633_bfr_before (
		.din(new_net_4633),
		.dout(new_net_4632)
	);

	bfr new_net_4634_bfr_before (
		.din(new_net_4634),
		.dout(new_net_4633)
	);

	bfr new_net_4635_bfr_before (
		.din(new_net_4635),
		.dout(new_net_4634)
	);

	bfr new_net_4636_bfr_before (
		.din(new_net_4636),
		.dout(new_net_4635)
	);

	bfr new_net_4637_bfr_before (
		.din(new_net_4637),
		.dout(new_net_4636)
	);

	bfr new_net_4638_bfr_before (
		.din(new_net_4638),
		.dout(new_net_4637)
	);

	bfr new_net_4639_bfr_before (
		.din(new_net_4639),
		.dout(new_net_4638)
	);

	bfr new_net_4640_bfr_before (
		.din(new_net_4640),
		.dout(new_net_4639)
	);

	bfr new_net_4641_bfr_before (
		.din(new_net_4641),
		.dout(new_net_4640)
	);

	bfr new_net_4642_bfr_before (
		.din(new_net_4642),
		.dout(new_net_4641)
	);

	bfr new_net_4643_bfr_before (
		.din(new_net_4643),
		.dout(new_net_4642)
	);

	bfr new_net_4644_bfr_before (
		.din(new_net_4644),
		.dout(new_net_4643)
	);

	bfr new_net_4645_bfr_before (
		.din(new_net_4645),
		.dout(new_net_4644)
	);

	bfr new_net_4646_bfr_before (
		.din(new_net_4646),
		.dout(new_net_4645)
	);

	bfr new_net_4647_bfr_before (
		.din(new_net_4647),
		.dout(new_net_4646)
	);

	bfr new_net_4648_bfr_before (
		.din(new_net_4648),
		.dout(new_net_4647)
	);

	bfr new_net_4649_bfr_before (
		.din(new_net_4649),
		.dout(new_net_4648)
	);

	bfr new_net_4650_bfr_before (
		.din(new_net_4650),
		.dout(new_net_4649)
	);

	bfr new_net_4651_bfr_before (
		.din(new_net_4651),
		.dout(new_net_4650)
	);

	bfr new_net_4652_bfr_before (
		.din(new_net_4652),
		.dout(new_net_4651)
	);

	bfr new_net_4653_bfr_before (
		.din(new_net_4653),
		.dout(new_net_4652)
	);

	bfr new_net_4654_bfr_before (
		.din(new_net_4654),
		.dout(new_net_4653)
	);

	bfr new_net_4655_bfr_before (
		.din(new_net_4655),
		.dout(new_net_4654)
	);

	bfr new_net_4656_bfr_before (
		.din(new_net_4656),
		.dout(new_net_4655)
	);

	spl2 _0997__v_fanout (
		.a(_0997_),
		.b(new_net_574),
		.c(new_net_4656)
	);

	spl2 _0083__v_fanout (
		.a(_0083_),
		.b(new_net_1634),
		.c(new_net_1635)
	);

	spl2 _0211__v_fanout (
		.a(_0211_),
		.b(new_net_1384),
		.c(new_net_1385)
	);

	spl2 _0917__v_fanout (
		.a(_0917_),
		.b(new_net_2002),
		.c(new_net_2003)
	);

	spl2 _0199__v_fanout (
		.a(_0199_),
		.b(new_net_2323),
		.c(new_net_2324)
	);

	spl2 _0325__v_fanout (
		.a(_0325_),
		.b(new_net_651),
		.c(new_net_652)
	);

	spl2 _0695__v_fanout (
		.a(_0695_),
		.b(new_net_1362),
		.c(new_net_1363)
	);

	spl2 _0205__v_fanout (
		.a(_0205_),
		.b(new_net_2468),
		.c(new_net_2469)
	);

	spl2 _0766__v_fanout (
		.a(_0766_),
		.b(new_net_1423),
		.c(new_net_1424)
	);

	spl2 _0820__v_fanout (
		.a(_0820_),
		.b(new_net_1882),
		.c(new_net_1883)
	);

	spl2 _0952__v_fanout (
		.a(_0952_),
		.b(new_net_2116),
		.c(new_net_2117)
	);

	spl2 _0608__v_fanout (
		.a(_0608_),
		.b(new_net_633),
		.c(new_net_634)
	);

	spl2 _0423__v_fanout (
		.a(_0423_),
		.b(new_net_140),
		.c(new_net_141)
	);

	spl2 _0528__v_fanout (
		.a(_0528_),
		.b(new_net_1950),
		.c(new_net_1951)
	);

	spl2 _0421__v_fanout (
		.a(_0421_),
		.b(new_net_2993),
		.c(new_net_2994)
	);

	spl2 _0315__v_fanout (
		.a(_0315_),
		.b(new_net_2941),
		.c(new_net_2942)
	);

	spl2 _0914__v_fanout (
		.a(_0914_),
		.b(new_net_1503),
		.c(new_net_1504)
	);

	bfr new_net_4657_bfr_after (
		.din(_1008_),
		.dout(new_net_4657)
	);

	bfr new_net_4658_bfr_after (
		.din(new_net_4657),
		.dout(new_net_4658)
	);

	bfr new_net_4659_bfr_after (
		.din(new_net_4658),
		.dout(new_net_4659)
	);

	bfr new_net_4660_bfr_after (
		.din(new_net_4659),
		.dout(new_net_4660)
	);

	bfr new_net_4661_bfr_after (
		.din(new_net_4660),
		.dout(new_net_4661)
	);

	bfr new_net_4662_bfr_after (
		.din(new_net_4661),
		.dout(new_net_4662)
	);

	bfr new_net_4663_bfr_after (
		.din(new_net_4662),
		.dout(new_net_4663)
	);

	bfr new_net_4664_bfr_after (
		.din(new_net_4663),
		.dout(new_net_4664)
	);

	bfr new_net_4665_bfr_after (
		.din(new_net_4664),
		.dout(new_net_4665)
	);

	bfr new_net_4666_bfr_after (
		.din(new_net_4665),
		.dout(new_net_4666)
	);

	bfr new_net_4667_bfr_after (
		.din(new_net_4666),
		.dout(new_net_4667)
	);

	bfr new_net_4668_bfr_after (
		.din(new_net_4667),
		.dout(new_net_4668)
	);

	bfr new_net_4669_bfr_after (
		.din(new_net_4668),
		.dout(new_net_4669)
	);

	bfr new_net_4670_bfr_after (
		.din(new_net_4669),
		.dout(new_net_4670)
	);

	bfr new_net_4671_bfr_after (
		.din(new_net_4670),
		.dout(new_net_4671)
	);

	bfr new_net_4672_bfr_after (
		.din(new_net_4671),
		.dout(new_net_4672)
	);

	bfr new_net_4673_bfr_after (
		.din(new_net_4672),
		.dout(new_net_4673)
	);

	bfr new_net_4674_bfr_after (
		.din(new_net_4673),
		.dout(new_net_4674)
	);

	bfr new_net_4675_bfr_after (
		.din(new_net_4674),
		.dout(new_net_4675)
	);

	bfr new_net_4676_bfr_after (
		.din(new_net_4675),
		.dout(new_net_4676)
	);

	bfr new_net_4677_bfr_after (
		.din(new_net_4676),
		.dout(new_net_4677)
	);

	bfr new_net_4678_bfr_after (
		.din(new_net_4677),
		.dout(new_net_4678)
	);

	bfr new_net_4679_bfr_after (
		.din(new_net_4678),
		.dout(new_net_4679)
	);

	bfr new_net_4680_bfr_after (
		.din(new_net_4679),
		.dout(new_net_4680)
	);

	bfr new_net_4681_bfr_after (
		.din(new_net_4680),
		.dout(new_net_4681)
	);

	bfr new_net_4682_bfr_after (
		.din(new_net_4681),
		.dout(new_net_4682)
	);

	bfr new_net_4683_bfr_after (
		.din(new_net_4682),
		.dout(new_net_4683)
	);

	bfr new_net_4684_bfr_after (
		.din(new_net_4683),
		.dout(new_net_4684)
	);

	bfr new_net_4685_bfr_after (
		.din(new_net_4684),
		.dout(new_net_4685)
	);

	bfr new_net_4686_bfr_after (
		.din(new_net_4685),
		.dout(new_net_4686)
	);

	bfr new_net_4687_bfr_after (
		.din(new_net_4686),
		.dout(new_net_4687)
	);

	bfr new_net_4688_bfr_after (
		.din(new_net_4687),
		.dout(new_net_4688)
	);

	bfr new_net_4689_bfr_after (
		.din(new_net_4688),
		.dout(new_net_4689)
	);

	bfr new_net_4690_bfr_after (
		.din(new_net_4689),
		.dout(new_net_4690)
	);

	bfr new_net_4691_bfr_after (
		.din(new_net_4690),
		.dout(new_net_4691)
	);

	bfr new_net_4692_bfr_after (
		.din(new_net_4691),
		.dout(new_net_4692)
	);

	bfr new_net_4693_bfr_after (
		.din(new_net_4692),
		.dout(new_net_4693)
	);

	bfr new_net_4694_bfr_after (
		.din(new_net_4693),
		.dout(new_net_4694)
	);

	bfr new_net_4695_bfr_after (
		.din(new_net_4694),
		.dout(new_net_4695)
	);

	bfr new_net_4696_bfr_after (
		.din(new_net_4695),
		.dout(new_net_4696)
	);

	bfr new_net_4697_bfr_after (
		.din(new_net_4696),
		.dout(new_net_4697)
	);

	bfr new_net_4698_bfr_after (
		.din(new_net_4697),
		.dout(new_net_4698)
	);

	bfr new_net_4699_bfr_after (
		.din(new_net_4698),
		.dout(new_net_4699)
	);

	bfr new_net_4700_bfr_after (
		.din(new_net_4699),
		.dout(new_net_4700)
	);

	bfr new_net_4701_bfr_after (
		.din(new_net_4700),
		.dout(new_net_4701)
	);

	bfr new_net_4702_bfr_after (
		.din(new_net_4701),
		.dout(new_net_4702)
	);

	bfr new_net_4703_bfr_after (
		.din(new_net_4702),
		.dout(new_net_4703)
	);

	bfr new_net_4704_bfr_after (
		.din(new_net_4703),
		.dout(new_net_4704)
	);

	bfr new_net_4705_bfr_after (
		.din(new_net_4704),
		.dout(new_net_4705)
	);

	bfr new_net_4706_bfr_after (
		.din(new_net_4705),
		.dout(new_net_4706)
	);

	bfr new_net_4707_bfr_after (
		.din(new_net_4706),
		.dout(new_net_4707)
	);

	bfr new_net_4708_bfr_after (
		.din(new_net_4707),
		.dout(new_net_4708)
	);

	bfr new_net_4709_bfr_after (
		.din(new_net_4708),
		.dout(new_net_4709)
	);

	bfr new_net_4710_bfr_after (
		.din(new_net_4709),
		.dout(new_net_4710)
	);

	bfr new_net_4711_bfr_after (
		.din(new_net_4710),
		.dout(new_net_4711)
	);

	bfr new_net_4712_bfr_after (
		.din(new_net_4711),
		.dout(new_net_4712)
	);

	bfr new_net_4713_bfr_after (
		.din(new_net_4712),
		.dout(new_net_4713)
	);

	bfr new_net_4714_bfr_after (
		.din(new_net_4713),
		.dout(new_net_4714)
	);

	spl2 _1008__v_fanout (
		.a(new_net_4714),
		.b(new_net_2635),
		.c(new_net_2636)
	);

	spl2 _1801__v_fanout (
		.a(_1801_),
		.b(new_net_1561),
		.c(new_net_1562)
	);

	bfr new_net_4715_bfr_after (
		.din(_0978_),
		.dout(new_net_4715)
	);

	bfr new_net_4716_bfr_after (
		.din(new_net_4715),
		.dout(new_net_4716)
	);

	spl2 _0978__v_fanout (
		.a(new_net_4716),
		.b(new_net_2789),
		.c(new_net_2790)
	);

	spl2 _0870__v_fanout (
		.a(_0870_),
		.b(new_net_2198),
		.c(new_net_2199)
	);

	spl2 _0606__v_fanout (
		.a(_0606_),
		.b(new_net_242),
		.c(new_net_243)
	);

	spl2 _0817__v_fanout (
		.a(_0817_),
		.b(new_net_2168),
		.c(new_net_2169)
	);

	spl2 _0518__v_fanout (
		.a(_0518_),
		.b(new_net_1616),
		.c(new_net_1617)
	);

	spl2 _0756__v_fanout (
		.a(_0756_),
		.b(new_net_1050),
		.c(new_net_1051)
	);

	spl2 _0685__v_fanout (
		.a(_0685_),
		.b(new_net_755),
		.c(new_net_756)
	);

	spl2 _0950__v_fanout (
		.a(_0950_),
		.b(new_net_725),
		.c(new_net_726)
	);

	spl2 _0082__v_fanout (
		.a(_0082_),
		.b(new_net_1435),
		.c(new_net_1436)
	);

	spl2 _0196__v_fanout (
		.a(_0196_),
		.b(new_net_1738),
		.c(new_net_1739)
	);

	spl2 _0986__v_fanout (
		.a(_0986_),
		.b(new_net_1792),
		.c(new_net_1793)
	);

	spl2 _1800__v_fanout (
		.a(_1800_),
		.b(new_net_1324),
		.c(new_net_1325)
	);

	spl2 _0976__v_fanout (
		.a(_0976_),
		.b(new_net_2416),
		.c(new_net_2417)
	);

	spl2 _0605__v_fanout (
		.a(_0605_),
		.b(new_net_76),
		.c(new_net_77)
	);

	spl2 _0684__v_fanout (
		.a(_0684_),
		.b(new_net_546),
		.c(new_net_547)
	);

	spl2 _0420__v_fanout (
		.a(_0420_),
		.b(new_net_1054),
		.c(new_net_1055)
	);

	spl2 _0081__v_fanout (
		.a(_0081_),
		.b(new_net_1228),
		.c(new_net_1229)
	);

	spl2 _0949__v_fanout (
		.a(_0949_),
		.b(new_net_518),
		.c(new_net_519)
	);

	spl2 _0314__v_fanout (
		.a(_0314_),
		.b(new_net_232),
		.c(new_net_233)
	);

	spl2 _0755__v_fanout (
		.a(_0755_),
		.b(new_net_1670),
		.c(new_net_1671)
	);

	spl2 _0517__v_fanout (
		.a(_0517_),
		.b(new_net_1575),
		.c(new_net_1576)
	);

	spl2 _0195__v_fanout (
		.a(_0195_),
		.b(new_net_2064),
		.c(new_net_2065)
	);

	spl2 _0869__v_fanout (
		.a(_0869_),
		.b(new_net_1138),
		.c(new_net_1139)
	);

	spl2 _0816__v_fanout (
		.a(_0816_),
		.b(new_net_1956),
		.c(new_net_1957)
	);

	spl2 _0913__v_fanout (
		.a(_0913_),
		.b(new_net_659),
		.c(new_net_660)
	);

	bfr new_net_4717_bfr_before (
		.din(new_net_4717),
		.dout(new_net_2564)
	);

	bfr new_net_4718_bfr_before (
		.din(new_net_4718),
		.dout(new_net_4717)
	);

	bfr new_net_4719_bfr_before (
		.din(new_net_4719),
		.dout(new_net_4718)
	);

	bfr new_net_4720_bfr_before (
		.din(new_net_4720),
		.dout(new_net_4719)
	);

	bfr new_net_4721_bfr_before (
		.din(new_net_4721),
		.dout(new_net_4720)
	);

	bfr new_net_4722_bfr_before (
		.din(new_net_4722),
		.dout(new_net_4721)
	);

	bfr new_net_4723_bfr_before (
		.din(new_net_4723),
		.dout(new_net_4722)
	);

	bfr new_net_4724_bfr_before (
		.din(new_net_4724),
		.dout(new_net_4723)
	);

	bfr new_net_4725_bfr_before (
		.din(new_net_4725),
		.dout(new_net_4724)
	);

	bfr new_net_4726_bfr_before (
		.din(new_net_4726),
		.dout(new_net_4725)
	);

	bfr new_net_4727_bfr_before (
		.din(new_net_4727),
		.dout(new_net_4726)
	);

	bfr new_net_4728_bfr_before (
		.din(new_net_4728),
		.dout(new_net_4727)
	);

	bfr new_net_4729_bfr_before (
		.din(new_net_4729),
		.dout(new_net_4728)
	);

	bfr new_net_4730_bfr_before (
		.din(new_net_4730),
		.dout(new_net_4729)
	);

	bfr new_net_4731_bfr_before (
		.din(new_net_4731),
		.dout(new_net_4730)
	);

	bfr new_net_4732_bfr_before (
		.din(new_net_4732),
		.dout(new_net_4731)
	);

	bfr new_net_4733_bfr_before (
		.din(new_net_4733),
		.dout(new_net_4732)
	);

	bfr new_net_4734_bfr_before (
		.din(new_net_4734),
		.dout(new_net_4733)
	);

	bfr new_net_4735_bfr_before (
		.din(new_net_4735),
		.dout(new_net_4734)
	);

	bfr new_net_4736_bfr_before (
		.din(new_net_4736),
		.dout(new_net_4735)
	);

	bfr new_net_4737_bfr_before (
		.din(new_net_4737),
		.dout(new_net_4736)
	);

	bfr new_net_4738_bfr_before (
		.din(new_net_4738),
		.dout(new_net_4737)
	);

	bfr new_net_4739_bfr_before (
		.din(new_net_4739),
		.dout(new_net_4738)
	);

	bfr new_net_4740_bfr_before (
		.din(new_net_4740),
		.dout(new_net_4739)
	);

	bfr new_net_4741_bfr_before (
		.din(new_net_4741),
		.dout(new_net_4740)
	);

	bfr new_net_4742_bfr_before (
		.din(new_net_4742),
		.dout(new_net_4741)
	);

	bfr new_net_4743_bfr_before (
		.din(new_net_4743),
		.dout(new_net_4742)
	);

	bfr new_net_4744_bfr_before (
		.din(new_net_4744),
		.dout(new_net_4743)
	);

	bfr new_net_4745_bfr_before (
		.din(new_net_4745),
		.dout(new_net_4744)
	);

	bfr new_net_4746_bfr_before (
		.din(new_net_4746),
		.dout(new_net_4745)
	);

	bfr new_net_4747_bfr_before (
		.din(new_net_4747),
		.dout(new_net_4746)
	);

	bfr new_net_4748_bfr_before (
		.din(new_net_4748),
		.dout(new_net_4747)
	);

	bfr new_net_4749_bfr_before (
		.din(new_net_4749),
		.dout(new_net_4748)
	);

	bfr new_net_4750_bfr_before (
		.din(new_net_4750),
		.dout(new_net_4749)
	);

	bfr new_net_4751_bfr_before (
		.din(new_net_4751),
		.dout(new_net_4750)
	);

	bfr new_net_4752_bfr_before (
		.din(new_net_4752),
		.dout(new_net_4751)
	);

	bfr new_net_4753_bfr_before (
		.din(new_net_4753),
		.dout(new_net_4752)
	);

	bfr new_net_4754_bfr_before (
		.din(new_net_4754),
		.dout(new_net_4753)
	);

	bfr new_net_4755_bfr_before (
		.din(new_net_4755),
		.dout(new_net_4754)
	);

	bfr new_net_4756_bfr_before (
		.din(new_net_4756),
		.dout(new_net_4755)
	);

	bfr new_net_4757_bfr_before (
		.din(new_net_4757),
		.dout(new_net_4756)
	);

	bfr new_net_4758_bfr_before (
		.din(new_net_4758),
		.dout(new_net_4757)
	);

	bfr new_net_4759_bfr_before (
		.din(new_net_4759),
		.dout(new_net_4758)
	);

	bfr new_net_4760_bfr_before (
		.din(new_net_4760),
		.dout(new_net_4759)
	);

	bfr new_net_4761_bfr_before (
		.din(new_net_4761),
		.dout(new_net_4760)
	);

	bfr new_net_4762_bfr_before (
		.din(new_net_4762),
		.dout(new_net_4761)
	);

	bfr new_net_4763_bfr_before (
		.din(new_net_4763),
		.dout(new_net_4762)
	);

	bfr new_net_4764_bfr_before (
		.din(new_net_4764),
		.dout(new_net_4763)
	);

	bfr new_net_4765_bfr_before (
		.din(new_net_4765),
		.dout(new_net_4764)
	);

	bfr new_net_4766_bfr_before (
		.din(new_net_4766),
		.dout(new_net_4765)
	);

	bfr new_net_4767_bfr_before (
		.din(new_net_4767),
		.dout(new_net_4766)
	);

	bfr new_net_4768_bfr_before (
		.din(new_net_4768),
		.dout(new_net_4767)
	);

	bfr new_net_4769_bfr_before (
		.din(new_net_4769),
		.dout(new_net_4768)
	);

	bfr new_net_4770_bfr_before (
		.din(new_net_4770),
		.dout(new_net_4769)
	);

	bfr new_net_4771_bfr_before (
		.din(new_net_4771),
		.dout(new_net_4770)
	);

	bfr new_net_4772_bfr_before (
		.din(new_net_4772),
		.dout(new_net_4771)
	);

	bfr new_net_4773_bfr_before (
		.din(new_net_4773),
		.dout(new_net_4772)
	);

	bfr new_net_4774_bfr_before (
		.din(new_net_4774),
		.dout(new_net_4773)
	);

	bfr new_net_4775_bfr_before (
		.din(new_net_4775),
		.dout(new_net_4774)
	);

	bfr new_net_4776_bfr_before (
		.din(new_net_4776),
		.dout(new_net_4775)
	);

	bfr new_net_4777_bfr_before (
		.din(new_net_4777),
		.dout(new_net_4776)
	);

	bfr new_net_4778_bfr_before (
		.din(new_net_4778),
		.dout(new_net_4777)
	);

	spl2 _1005__v_fanout (
		.a(_1005_),
		.b(new_net_2563),
		.c(new_net_4778)
	);

	bfr new_net_4779_bfr_before (
		.din(new_net_4779),
		.dout(new_net_3229)
	);

	bfr new_net_4780_bfr_before (
		.din(new_net_4780),
		.dout(new_net_4779)
	);

	bfr new_net_4781_bfr_before (
		.din(new_net_4781),
		.dout(new_net_4780)
	);

	bfr new_net_4782_bfr_before (
		.din(new_net_4782),
		.dout(new_net_4781)
	);

	spl2 _0946__v_fanout (
		.a(_0946_),
		.b(new_net_3228),
		.c(new_net_4782)
	);

	bfr new_net_4783_bfr_before (
		.din(new_net_4783),
		.dout(new_net_2894)
	);

	bfr new_net_4784_bfr_before (
		.din(new_net_4784),
		.dout(new_net_4783)
	);

	bfr new_net_4785_bfr_before (
		.din(new_net_4785),
		.dout(new_net_4784)
	);

	bfr new_net_4786_bfr_before (
		.din(new_net_4786),
		.dout(new_net_4785)
	);

	spl2 _0603__v_fanout (
		.a(_0603_),
		.b(new_net_2893),
		.c(new_net_4786)
	);

	bfr new_net_4787_bfr_before (
		.din(new_net_4787),
		.dout(new_net_1677)
	);

	bfr new_net_4788_bfr_before (
		.din(new_net_4788),
		.dout(new_net_4787)
	);

	bfr new_net_4789_bfr_before (
		.din(new_net_4789),
		.dout(new_net_4788)
	);

	bfr new_net_4790_bfr_before (
		.din(new_net_4790),
		.dout(new_net_4789)
	);

	spl2 _0814__v_fanout (
		.a(_0814_),
		.b(new_net_1676),
		.c(new_net_4790)
	);

	bfr new_net_4791_bfr_before (
		.din(new_net_4791),
		.dout(new_net_2439)
	);

	bfr new_net_4792_bfr_before (
		.din(new_net_4792),
		.dout(new_net_4791)
	);

	bfr new_net_4793_bfr_before (
		.din(new_net_4793),
		.dout(new_net_4792)
	);

	bfr new_net_4794_bfr_before (
		.din(new_net_4794),
		.dout(new_net_4793)
	);

	spl2 _0078__v_fanout (
		.a(_0078_),
		.b(new_net_2438),
		.c(new_net_4794)
	);

	bfr new_net_4795_bfr_before (
		.din(new_net_4795),
		.dout(new_net_2322)
	);

	bfr new_net_4796_bfr_before (
		.din(new_net_4796),
		.dout(new_net_4795)
	);

	bfr new_net_4797_bfr_before (
		.din(new_net_4797),
		.dout(new_net_4796)
	);

	bfr new_net_4798_bfr_before (
		.din(new_net_4798),
		.dout(new_net_4797)
	);

	spl2 _0312__v_fanout (
		.a(_0312_),
		.b(new_net_2321),
		.c(new_net_4798)
	);

	bfr new_net_4799_bfr_before (
		.din(new_net_4799),
		.dout(new_net_2063)
	);

	bfr new_net_4800_bfr_before (
		.din(new_net_4800),
		.dout(new_net_4799)
	);

	bfr new_net_4801_bfr_before (
		.din(new_net_4801),
		.dout(new_net_4800)
	);

	bfr new_net_4802_bfr_before (
		.din(new_net_4802),
		.dout(new_net_4801)
	);

	spl2 _0867__v_fanout (
		.a(_0867_),
		.b(new_net_2062),
		.c(new_net_4802)
	);

	bfr new_net_4803_bfr_after (
		.din(_0996_),
		.dout(new_net_4803)
	);

	bfr new_net_4804_bfr_after (
		.din(new_net_4803),
		.dout(new_net_4804)
	);

	bfr new_net_4805_bfr_after (
		.din(new_net_4804),
		.dout(new_net_4805)
	);

	bfr new_net_4806_bfr_after (
		.din(new_net_4805),
		.dout(new_net_4806)
	);

	spl2 _0996__v_fanout (
		.a(new_net_4806),
		.b(new_net_343),
		.c(new_net_344)
	);

	spl2 _0975__v_fanout (
		.a(_0975_),
		.b(new_net_2204),
		.c(new_net_2205)
	);

	bfr new_net_4807_bfr_before (
		.din(new_net_4807),
		.dout(new_net_2660)
	);

	bfr new_net_4808_bfr_before (
		.din(new_net_4808),
		.dout(new_net_4807)
	);

	bfr new_net_4809_bfr_before (
		.din(new_net_4809),
		.dout(new_net_4808)
	);

	bfr new_net_4810_bfr_before (
		.din(new_net_4810),
		.dout(new_net_4809)
	);

	spl2 _0515__v_fanout (
		.a(_0515_),
		.b(new_net_2659),
		.c(new_net_4810)
	);

	bfr new_net_4811_bfr_before (
		.din(new_net_4811),
		.dout(new_net_163)
	);

	bfr new_net_4812_bfr_before (
		.din(new_net_4812),
		.dout(new_net_4811)
	);

	bfr new_net_4813_bfr_before (
		.din(new_net_4813),
		.dout(new_net_4812)
	);

	bfr new_net_4814_bfr_before (
		.din(new_net_4814),
		.dout(new_net_4813)
	);

	spl2 _0682__v_fanout (
		.a(_0682_),
		.b(new_net_162),
		.c(new_net_4814)
	);

	bfr new_net_4815_bfr_before (
		.din(new_net_4815),
		.dout(new_net_1191)
	);

	bfr new_net_4816_bfr_before (
		.din(new_net_4816),
		.dout(new_net_4815)
	);

	bfr new_net_4817_bfr_before (
		.din(new_net_4817),
		.dout(new_net_4816)
	);

	bfr new_net_4818_bfr_before (
		.din(new_net_4818),
		.dout(new_net_4817)
	);

	spl2 _0193__v_fanout (
		.a(_0193_),
		.b(new_net_1190),
		.c(new_net_4818)
	);

	bfr new_net_4819_bfr_before (
		.din(new_net_4819),
		.dout(new_net_821)
	);

	bfr new_net_4820_bfr_before (
		.din(new_net_4820),
		.dout(new_net_4819)
	);

	bfr new_net_4821_bfr_before (
		.din(new_net_4821),
		.dout(new_net_4820)
	);

	bfr new_net_4822_bfr_before (
		.din(new_net_4822),
		.dout(new_net_4821)
	);

	spl2 _1798__v_fanout (
		.a(_1798_),
		.b(new_net_820),
		.c(new_net_4822)
	);

	bfr new_net_4823_bfr_before (
		.din(new_net_4823),
		.dout(new_net_1091)
	);

	bfr new_net_4824_bfr_before (
		.din(new_net_4824),
		.dout(new_net_4823)
	);

	bfr new_net_4825_bfr_before (
		.din(new_net_4825),
		.dout(new_net_4824)
	);

	bfr new_net_4826_bfr_before (
		.din(new_net_4826),
		.dout(new_net_4825)
	);

	spl2 _0752__v_fanout (
		.a(_0752_),
		.b(new_net_1090),
		.c(new_net_4826)
	);

	bfr new_net_4827_bfr_before (
		.din(new_net_4827),
		.dout(new_net_991)
	);

	bfr new_net_4828_bfr_before (
		.din(new_net_4828),
		.dout(new_net_4827)
	);

	bfr new_net_4829_bfr_before (
		.din(new_net_4829),
		.dout(new_net_4828)
	);

	bfr new_net_4830_bfr_before (
		.din(new_net_4830),
		.dout(new_net_4829)
	);

	spl2 _0418__v_fanout (
		.a(_0418_),
		.b(new_net_990),
		.c(new_net_4830)
	);

	spl2 _1004__v_fanout (
		.a(_1004_),
		.b(new_net_1822),
		.c(new_net_1823)
	);

	bfr new_net_4831_bfr_before (
		.din(new_net_4831),
		.dout(new_net_949)
	);

	bfr new_net_4832_bfr_before (
		.din(new_net_4832),
		.dout(new_net_4831)
	);

	bfr new_net_4833_bfr_before (
		.din(new_net_4833),
		.dout(new_net_4832)
	);

	bfr new_net_4834_bfr_before (
		.din(new_net_4834),
		.dout(new_net_4833)
	);

	spl2 _0911__v_fanout (
		.a(_0911_),
		.b(new_net_948),
		.c(new_net_4834)
	);

	spl2 _0697__v_fanout (
		.a(_0697_),
		.b(new_net_412),
		.c(new_net_413)
	);

	spl2 _0327__v_fanout (
		.a(_0327_),
		.b(new_net_1930),
		.c(new_net_1931)
	);

	spl2 _0813__v_fanout (
		.a(_0813_),
		.b(new_net_1642),
		.c(new_net_1643)
	);

	spl2 _0311__v_fanout (
		.a(_0311_),
		.b(new_net_2130),
		.c(new_net_2131)
	);

	spl2 _1679__v_fanout (
		.a(_1679_),
		.b(new_net_1852),
		.c(new_net_1853)
	);

	spl2 _0076__v_fanout (
		.a(_0076_),
		.b(new_net_2290),
		.c(new_net_2291)
	);

	spl2 _0530__v_fanout (
		.a(_0530_),
		.b(new_net_3057),
		.c(new_net_3058)
	);

	spl2 _0927__v_fanout (
		.a(_0927_),
		.b(new_net_783),
		.c(new_net_784)
	);

	spl2 _0681__v_fanout (
		.a(_0681_),
		.b(new_net_1370),
		.c(new_net_1371)
	);

	spl2 _0213__v_fanout (
		.a(_0213_),
		.b(new_net_1742),
		.c(new_net_1743)
	);

	spl2 _0618__v_fanout (
		.a(_0618_),
		.b(new_net_616),
		.c(new_net_617)
	);

	spl2 _1803__v_fanout (
		.a(_1803_),
		.b(new_net_1864),
		.c(new_net_1865)
	);

	spl2 _0192__v_fanout (
		.a(_0192_),
		.b(new_net_1026),
		.c(new_net_1027)
	);

	spl2 _0085__v_fanout (
		.a(_0085_),
		.b(new_net_1966),
		.c(new_net_1967)
	);

	spl2 _0751__v_fanout (
		.a(_0751_),
		.b(new_net_898),
		.c(new_net_899)
	);

	spl2 _1797__v_fanout (
		.a(_1797_),
		.b(new_net_830),
		.c(new_net_831)
	);

	spl2 _0417__v_fanout (
		.a(_0417_),
		.b(new_net_2182),
		.c(new_net_2183)
	);

	spl2 _0768__v_fanout (
		.a(_0768_),
		.b(new_net_1529),
		.c(new_net_1530)
	);

	spl2 _0866__v_fanout (
		.a(_0866_),
		.b(new_net_2016),
		.c(new_net_2017)
	);

	spl2 _0433__v_fanout (
		.a(_0433_),
		.b(new_net_1972),
		.c(new_net_1973)
	);

	spl2 _0883__v_fanout (
		.a(_0883_),
		.b(new_net_2722),
		.c(new_net_2723)
	);

	spl2 _0830__v_fanout (
		.a(_0830_),
		.b(new_net_1398),
		.c(new_net_1399)
	);

	spl2 _0602__v_fanout (
		.a(_0602_),
		.b(new_net_2689),
		.c(new_net_2690)
	);

	spl2 _0513__v_fanout (
		.a(_0513_),
		.b(new_net_2254),
		.c(new_net_2255)
	);

	spl2 _0994__v_fanout (
		.a(_0994_),
		.b(new_net_1),
		.c(new_net_2)
	);

	spl2 _0910__v_fanout (
		.a(_0910_),
		.b(new_net_775),
		.c(new_net_776)
	);

	bfr new_net_4835_bfr_before (
		.din(new_net_4835),
		.dout(new_net_2962)
	);

	bfr new_net_4836_bfr_before (
		.din(new_net_4836),
		.dout(new_net_4835)
	);

	bfr new_net_4837_bfr_before (
		.din(new_net_4837),
		.dout(new_net_4836)
	);

	bfr new_net_4838_bfr_before (
		.din(new_net_4838),
		.dout(new_net_4837)
	);

	spl2 _0973__v_fanout (
		.a(_0973_),
		.b(new_net_2961),
		.c(new_net_4838)
	);

	spl2 _1675__v_fanout (
		.a(_1675_),
		.b(new_net_906),
		.c(new_net_907)
	);

	spl2 _0414__v_fanout (
		.a(_0414_),
		.b(new_net_880),
		.c(new_net_881)
	);

	spl2 _0749__v_fanout (
		.a(_0749_),
		.b(new_net_576),
		.c(new_net_577)
	);

	spl2 _0190__v_fanout (
		.a(_0190_),
		.b(new_net_1876),
		.c(new_net_1877)
	);

	spl2 _0599__v_fanout (
		.a(_0599_),
		.b(new_net_3161),
		.c(new_net_3162)
	);

	spl2 _0679__v_fanout (
		.a(_0679_),
		.b(new_net_2793),
		.c(new_net_2794)
	);

	spl2 _0309__v_fanout (
		.a(_0309_),
		.b(new_net_60),
		.c(new_net_61)
	);

	spl2 _0074__v_fanout (
		.a(_0074_),
		.b(new_net_2268),
		.c(new_net_2269)
	);

	bfr new_net_4839_bfr_after (
		.din(_0945_),
		.dout(new_net_4839)
	);

	bfr new_net_4840_bfr_after (
		.din(new_net_4839),
		.dout(new_net_4840)
	);

	spl2 _0945__v_fanout (
		.a(new_net_4840),
		.b(new_net_2991),
		.c(new_net_2992)
	);

	spl2 _0962__v_fanout (
		.a(_0962_),
		.b(new_net_3007),
		.c(new_net_3008)
	);

	spl2 _0511__v_fanout (
		.a(_0511_),
		.b(new_net_1862),
		.c(new_net_1863)
	);

	spl2 _0993__v_fanout (
		.a(_0993_),
		.b(new_net_3035),
		.c(new_net_3036)
	);

	spl2 _0908__v_fanout (
		.a(_0908_),
		.b(new_net_468),
		.c(new_net_469)
	);

	spl2 _0864__v_fanout (
		.a(_0864_),
		.b(new_net_224),
		.c(new_net_225)
	);

	spl2 _1794__v_fanout (
		.a(_1794_),
		.b(new_net_618),
		.c(new_net_619)
	);

	spl2 _0811__v_fanout (
		.a(_0811_),
		.b(new_net_2100),
		.c(new_net_2101)
	);

	bfr new_net_4841_bfr_before (
		.din(new_net_4841),
		.dout(new_net_2630)
	);

	bfr new_net_4842_bfr_before (
		.din(new_net_4842),
		.dout(new_net_4841)
	);

	bfr new_net_4843_bfr_before (
		.din(new_net_4843),
		.dout(new_net_4842)
	);

	bfr new_net_4844_bfr_before (
		.din(new_net_4844),
		.dout(new_net_4843)
	);

	spl2 _0991__v_fanout (
		.a(_0991_),
		.b(new_net_2629),
		.c(new_net_4844)
	);

	spl2 _0598__v_fanout (
		.a(_0598_),
		.b(new_net_2937),
		.c(new_net_2938)
	);

	spl2 _0907__v_fanout (
		.a(_0907_),
		.b(new_net_414),
		.c(new_net_415)
	);

	spl2 _0308__v_fanout (
		.a(_0308_),
		.b(new_net_1602),
		.c(new_net_1603)
	);

	spl2 _0413__v_fanout (
		.a(_0413_),
		.b(new_net_848),
		.c(new_net_849)
	);

	spl2 _0678__v_fanout (
		.a(_0678_),
		.b(new_net_2623),
		.c(new_net_2624)
	);

	spl2 _0748__v_fanout (
		.a(_0748_),
		.b(new_net_824),
		.c(new_net_825)
	);

	spl2 _0863__v_fanout (
		.a(_0863_),
		.b(new_net_1910),
		.c(new_net_1911)
	);

	spl2 _1793__v_fanout (
		.a(_1793_),
		.b(new_net_592),
		.c(new_net_593)
	);

	spl2 _0510__v_fanout (
		.a(_0510_),
		.b(new_net_1271),
		.c(new_net_1272)
	);

	spl2 _0073__v_fanout (
		.a(_0073_),
		.b(new_net_2983),
		.c(new_net_2984)
	);

	spl2 _1674__v_fanout (
		.a(_1674_),
		.b(new_net_882),
		.c(new_net_883)
	);

	spl2 _0810__v_fanout (
		.a(_0810_),
		.b(new_net_1537),
		.c(new_net_1538)
	);

	spl2 _0943__v_fanout (
		.a(_0943_),
		.b(new_net_2581),
		.c(new_net_2582)
	);

	spl2 _0189__v_fanout (
		.a(_0189_),
		.b(new_net_1844),
		.c(new_net_1845)
	);

	bfr new_net_4845_bfr_after (
		.din(_0972_),
		.dout(new_net_4845)
	);

	bfr new_net_4846_bfr_after (
		.din(new_net_4845),
		.dout(new_net_4846)
	);

	bfr new_net_4847_bfr_after (
		.din(new_net_4846),
		.dout(new_net_4847)
	);

	bfr new_net_4848_bfr_after (
		.din(new_net_4847),
		.dout(new_net_4848)
	);

	spl2 _0972__v_fanout (
		.a(new_net_4848),
		.b(new_net_2925),
		.c(new_net_2926)
	);

	bfr new_net_4849_bfr_before (
		.din(new_net_4849),
		.dout(new_net_2522)
	);

	bfr new_net_4850_bfr_before (
		.din(new_net_4850),
		.dout(new_net_4849)
	);

	bfr new_net_4851_bfr_before (
		.din(new_net_4851),
		.dout(new_net_4850)
	);

	bfr new_net_4852_bfr_before (
		.din(new_net_4852),
		.dout(new_net_4851)
	);

	spl2 _0596__v_fanout (
		.a(_0596_),
		.b(new_net_2521),
		.c(new_net_4852)
	);

	bfr new_net_4853_bfr_before (
		.din(new_net_4853),
		.dout(new_net_1181)
	);

	bfr new_net_4854_bfr_before (
		.din(new_net_4854),
		.dout(new_net_4853)
	);

	bfr new_net_4855_bfr_before (
		.din(new_net_4855),
		.dout(new_net_4854)
	);

	bfr new_net_4856_bfr_before (
		.din(new_net_4856),
		.dout(new_net_4855)
	);

	spl2 _0508__v_fanout (
		.a(_0508_),
		.b(new_net_1180),
		.c(new_net_4856)
	);

	bfr new_net_4857_bfr_before (
		.din(new_net_4857),
		.dout(new_net_2846)
	);

	bfr new_net_4858_bfr_before (
		.din(new_net_4858),
		.dout(new_net_4857)
	);

	bfr new_net_4859_bfr_before (
		.din(new_net_4859),
		.dout(new_net_4858)
	);

	bfr new_net_4860_bfr_before (
		.din(new_net_4860),
		.dout(new_net_4859)
	);

	spl2 _1791__v_fanout (
		.a(_1791_),
		.b(new_net_2845),
		.c(new_net_4860)
	);

	bfr new_net_4861_bfr_before (
		.din(new_net_4861),
		.dout(new_net_2576)
	);

	bfr new_net_4862_bfr_before (
		.din(new_net_4862),
		.dout(new_net_4861)
	);

	bfr new_net_4863_bfr_before (
		.din(new_net_4863),
		.dout(new_net_4862)
	);

	bfr new_net_4864_bfr_before (
		.din(new_net_4864),
		.dout(new_net_4863)
	);

	spl2 _0071__v_fanout (
		.a(_0071_),
		.b(new_net_2575),
		.c(new_net_4864)
	);

	bfr new_net_4865_bfr_before (
		.din(new_net_4865),
		.dout(new_net_1153)
	);

	bfr new_net_4866_bfr_before (
		.din(new_net_4866),
		.dout(new_net_4865)
	);

	bfr new_net_4867_bfr_before (
		.din(new_net_4867),
		.dout(new_net_4866)
	);

	bfr new_net_4868_bfr_before (
		.din(new_net_4868),
		.dout(new_net_4867)
	);

	spl2 _0675__v_fanout (
		.a(_0675_),
		.b(new_net_1152),
		.c(new_net_4868)
	);

	bfr new_net_4869_bfr_before (
		.din(new_net_4869),
		.dout(new_net_1589)
	);

	bfr new_net_4870_bfr_before (
		.din(new_net_4870),
		.dout(new_net_4869)
	);

	bfr new_net_4871_bfr_before (
		.din(new_net_4871),
		.dout(new_net_4870)
	);

	bfr new_net_4872_bfr_before (
		.din(new_net_4872),
		.dout(new_net_4871)
	);

	spl2 _0808__v_fanout (
		.a(_0808_),
		.b(new_net_1588),
		.c(new_net_4872)
	);

	bfr new_net_4873_bfr_before (
		.din(new_net_4873),
		.dout(new_net_823)
	);

	bfr new_net_4874_bfr_before (
		.din(new_net_4874),
		.dout(new_net_4873)
	);

	bfr new_net_4875_bfr_before (
		.din(new_net_4875),
		.dout(new_net_4874)
	);

	bfr new_net_4876_bfr_before (
		.din(new_net_4876),
		.dout(new_net_4875)
	);

	spl2 _1672__v_fanout (
		.a(_1672_),
		.b(new_net_822),
		.c(new_net_4876)
	);

	bfr new_net_4877_bfr_before (
		.din(new_net_4877),
		.dout(new_net_9)
	);

	bfr new_net_4878_bfr_before (
		.din(new_net_4878),
		.dout(new_net_4877)
	);

	bfr new_net_4879_bfr_before (
		.din(new_net_4879),
		.dout(new_net_4878)
	);

	bfr new_net_4880_bfr_before (
		.din(new_net_4880),
		.dout(new_net_4879)
	);

	spl2 _0746__v_fanout (
		.a(_0746_),
		.b(new_net_8),
		.c(new_net_4880)
	);

	bfr new_net_4881_bfr_before (
		.din(new_net_4881),
		.dout(new_net_2385)
	);

	bfr new_net_4882_bfr_before (
		.din(new_net_4882),
		.dout(new_net_4881)
	);

	bfr new_net_4883_bfr_before (
		.din(new_net_4883),
		.dout(new_net_4882)
	);

	bfr new_net_4884_bfr_before (
		.din(new_net_4884),
		.dout(new_net_4883)
	);

	spl2 _0305__v_fanout (
		.a(_0305_),
		.b(new_net_2384),
		.c(new_net_4884)
	);

	bfr new_net_4885_bfr_before (
		.din(new_net_4885),
		.dout(new_net_334)
	);

	bfr new_net_4886_bfr_before (
		.din(new_net_4886),
		.dout(new_net_4885)
	);

	bfr new_net_4887_bfr_before (
		.din(new_net_4887),
		.dout(new_net_4886)
	);

	bfr new_net_4888_bfr_before (
		.din(new_net_4888),
		.dout(new_net_4887)
	);

	spl2 _0905__v_fanout (
		.a(_0905_),
		.b(new_net_333),
		.c(new_net_4888)
	);

	spl2 _0942__v_fanout (
		.a(_0942_),
		.b(new_net_2382),
		.c(new_net_2383)
	);

	bfr new_net_4889_bfr_before (
		.din(new_net_4889),
		.dout(new_net_1795)
	);

	bfr new_net_4890_bfr_before (
		.din(new_net_4890),
		.dout(new_net_4889)
	);

	bfr new_net_4891_bfr_before (
		.din(new_net_4891),
		.dout(new_net_4890)
	);

	bfr new_net_4892_bfr_before (
		.din(new_net_4892),
		.dout(new_net_4891)
	);

	spl2 _0860__v_fanout (
		.a(_0860_),
		.b(new_net_1794),
		.c(new_net_4892)
	);

	bfr new_net_4893_bfr_before (
		.din(new_net_4893),
		.dout(new_net_1729)
	);

	bfr new_net_4894_bfr_before (
		.din(new_net_4894),
		.dout(new_net_4893)
	);

	bfr new_net_4895_bfr_before (
		.din(new_net_4895),
		.dout(new_net_4894)
	);

	bfr new_net_4896_bfr_before (
		.din(new_net_4896),
		.dout(new_net_4895)
	);

	spl2 _0186__v_fanout (
		.a(_0186_),
		.b(new_net_1728),
		.c(new_net_4896)
	);

	spl2 _0990__v_fanout (
		.a(_0990_),
		.b(new_net_2422),
		.c(new_net_2423)
	);

	bfr new_net_4897_bfr_before (
		.din(new_net_4897),
		.dout(new_net_1063)
	);

	bfr new_net_4898_bfr_before (
		.din(new_net_4898),
		.dout(new_net_4897)
	);

	bfr new_net_4899_bfr_before (
		.din(new_net_4899),
		.dout(new_net_4898)
	);

	bfr new_net_4900_bfr_before (
		.din(new_net_4900),
		.dout(new_net_4899)
	);

	spl2 _0411__v_fanout (
		.a(_0411_),
		.b(new_net_1062),
		.c(new_net_4900)
	);

	spl2 _0806__v_fanout (
		.a(_0806_),
		.b(new_net_1160),
		.c(new_net_1161)
	);

	spl2 _0304__v_fanout (
		.a(_0304_),
		.b(new_net_3117),
		.c(new_net_3118)
	);

	spl2 _0215__v_fanout (
		.a(_0215_),
		.b(new_net_2136),
		.c(new_net_2137)
	);

	spl2 _1671__v_fanout (
		.a(_1671_),
		.b(new_net_761),
		.c(new_net_762)
	);

	spl2 _0970__v_fanout (
		.a(_0970_),
		.b(new_net_1243),
		.c(new_net_1244)
	);

	spl2 _0070__v_fanout (
		.a(_0070_),
		.b(new_net_2108),
		.c(new_net_2109)
	);

	spl2 _0185__v_fanout (
		.a(_0185_),
		.b(new_net_2935),
		.c(new_net_2936)
	);

	spl2 _0674__v_fanout (
		.a(_0674_),
		.b(new_net_1112),
		.c(new_net_1113)
	);

	spl2 _0435__v_fanout (
		.a(_0435_),
		.b(new_net_66),
		.c(new_net_67)
	);

	spl2 _0620__v_fanout (
		.a(_0620_),
		.b(new_net_2899),
		.c(new_net_2900)
	);

	spl2 _0745__v_fanout (
		.a(_0745_),
		.b(new_net_3039),
		.c(new_net_3040)
	);

	spl2 _1805__v_fanout (
		.a(_1805_),
		.b(new_net_2256),
		.c(new_net_2257)
	);

	spl2 _0595__v_fanout (
		.a(_0595_),
		.b(new_net_2317),
		.c(new_net_2318)
	);

	bfr new_net_4901_bfr_before (
		.din(new_net_4901),
		.dout(new_net_1969)
	);

	bfr new_net_4902_bfr_before (
		.din(new_net_4902),
		.dout(new_net_4901)
	);

	bfr new_net_4903_bfr_before (
		.din(new_net_4903),
		.dout(new_net_4902)
	);

	bfr new_net_4904_bfr_before (
		.din(new_net_4904),
		.dout(new_net_4903)
	);

	spl2 _0940__v_fanout (
		.a(_0940_),
		.b(new_net_1968),
		.c(new_net_4904)
	);

	spl2 _0700__v_fanout (
		.a(_0700_),
		.b(new_net_2313),
		.c(new_net_2314)
	);

	spl2 _0770__v_fanout (
		.a(_0770_),
		.b(new_net_834),
		.c(new_net_835)
	);

	spl2 _1561__v_fanout (
		.a(_1561_),
		.b(new_net_2967),
		.c(new_net_2968)
	);

	spl2 _0410__v_fanout (
		.a(_0410_),
		.b(new_net_713),
		.c(new_net_714)
	);

	spl2 _0087__v_fanout (
		.a(_0087_),
		.b(new_net_2781),
		.c(new_net_2782)
	);

	spl2 _0507__v_fanout (
		.a(_0507_),
		.b(new_net_1150),
		.c(new_net_1151)
	);

	spl2 _0532__v_fanout (
		.a(_0532_),
		.b(new_net_2112),
		.c(new_net_2113)
	);

	spl2 _1790__v_fanout (
		.a(_1790_),
		.b(new_net_2661),
		.c(new_net_2662)
	);

	spl2 _0885__v_fanout (
		.a(_0885_),
		.b(new_net_2779),
		.c(new_net_2780)
	);

	spl2 _0330__v_fanout (
		.a(_0330_),
		.b(new_net_2525),
		.c(new_net_2526)
	);

	spl2 _0859__v_fanout (
		.a(_0859_),
		.b(new_net_1756),
		.c(new_net_1757)
	);

	spl2 _1681__v_fanout (
		.a(_1681_),
		.b(new_net_2250),
		.c(new_net_2251)
	);

	spl2 _0832__v_fanout (
		.a(_0832_),
		.b(new_net_1766),
		.c(new_net_1767)
	);

	spl2 _0068__v_fanout (
		.a(_0068_),
		.b(new_net_1960),
		.c(new_net_1961)
	);

	spl2 _1788__v_fanout (
		.a(_1788_),
		.b(new_net_368),
		.c(new_net_369)
	);

	spl2 _1669__v_fanout (
		.a(_1669_),
		.b(new_net_667),
		.c(new_net_668)
	);

	spl2 _0408__v_fanout (
		.a(_0408_),
		.b(new_net_514),
		.c(new_net_515)
	);

	spl2 _0302__v_fanout (
		.a(_0302_),
		.b(new_net_1774),
		.c(new_net_1775)
	);

	spl2 _0969__v_fanout (
		.a(_0969_),
		.b(new_net_1066),
		.c(new_net_1067)
	);

	spl2 _0505__v_fanout (
		.a(_0505_),
		.b(new_net_816),
		.c(new_net_817)
	);

	bfr new_net_4905_bfr_after (
		.din(_0903_),
		.dout(new_net_4905)
	);

	bfr new_net_4906_bfr_after (
		.din(new_net_4905),
		.dout(new_net_4906)
	);

	spl2 _0903__v_fanout (
		.a(new_net_4906),
		.b(new_net_283),
		.c(new_net_284)
	);

	spl2 _0672__v_fanout (
		.a(_0672_),
		.b(new_net_1461),
		.c(new_net_1462)
	);

	spl2 _0183__v_fanout (
		.a(_0183_),
		.b(new_net_2519),
		.c(new_net_2520)
	);

	spl2 _0743__v_fanout (
		.a(_0743_),
		.b(new_net_594),
		.c(new_net_595)
	);

	spl2 _0804__v_fanout (
		.a(_0804_),
		.b(new_net_858),
		.c(new_net_859)
	);

	spl2 _1558__v_fanout (
		.a(_1558_),
		.b(new_net_685),
		.c(new_net_686)
	);

	spl2 _0929__v_fanout (
		.a(_0929_),
		.b(new_net_1210),
		.c(new_net_1211)
	);

	spl2 _0857__v_fanout (
		.a(_0857_),
		.b(new_net_2080),
		.c(new_net_2081)
	);

	spl2 _0593__v_fanout (
		.a(_0593_),
		.b(new_net_1926),
		.c(new_net_1927)
	);

	bfr new_net_4907_bfr_before (
		.din(new_net_4907),
		.dout(new_net_2682)
	);

	bfr new_net_4908_bfr_before (
		.din(new_net_4908),
		.dout(new_net_4907)
	);

	bfr new_net_4909_bfr_before (
		.din(new_net_4909),
		.dout(new_net_4908)
	);

	bfr new_net_4910_bfr_before (
		.din(new_net_4910),
		.dout(new_net_4909)
	);

	spl2 _0966__v_fanout (
		.a(_0966_),
		.b(new_net_2681),
		.c(new_net_4910)
	);

	spl2 _0671__v_fanout (
		.a(_0671_),
		.b(new_net_1263),
		.c(new_net_1264)
	);

	spl2 _1557__v_fanout (
		.a(_1557_),
		.b(new_net_490),
		.c(new_net_491)
	);

	spl2 _1787__v_fanout (
		.a(_1787_),
		.b(new_net_2040),
		.c(new_net_2041)
	);

	spl2 _0301__v_fanout (
		.a(_0301_),
		.b(new_net_1638),
		.c(new_net_1639)
	);

	spl2 _0592__v_fanout (
		.a(_0592_),
		.b(new_net_2807),
		.c(new_net_2808)
	);

	spl2 _0803__v_fanout (
		.a(_0803_),
		.b(new_net_1216),
		.c(new_net_1217)
	);

	spl2 _0901__v_fanout (
		.a(_0901_),
		.b(new_net_198),
		.c(new_net_199)
	);

	spl2 _1668__v_fanout (
		.a(_1668_),
		.b(new_net_624),
		.c(new_net_625)
	);

	spl2 _0504__v_fanout (
		.a(_0504_),
		.b(new_net_590),
		.c(new_net_591)
	);

	spl2 _0067__v_fanout (
		.a(_0067_),
		.b(new_net_1978),
		.c(new_net_1979)
	);

	spl2 _0741__v_fanout (
		.a(_0741_),
		.b(new_net_2224),
		.c(new_net_2225)
	);

	spl2 _0407__v_fanout (
		.a(_0407_),
		.b(new_net_596),
		.c(new_net_597)
	);

	spl2 _0182__v_fanout (
		.a(_0182_),
		.b(new_net_1612),
		.c(new_net_1613)
	);

	spl2 _0856__v_fanout (
		.a(_0856_),
		.b(new_net_1694),
		.c(new_net_1695)
	);

	bfr new_net_4911_bfr_before (
		.din(new_net_4911),
		.dout(new_net_965)
	);

	bfr new_net_4912_bfr_before (
		.din(new_net_4912),
		.dout(new_net_4911)
	);

	bfr new_net_4913_bfr_before (
		.din(new_net_4913),
		.dout(new_net_4912)
	);

	bfr new_net_4914_bfr_before (
		.din(new_net_4914),
		.dout(new_net_4913)
	);

	spl2 _0669__v_fanout (
		.a(_0669_),
		.b(new_net_964),
		.c(new_net_4914)
	);

	bfr new_net_4915_bfr_before (
		.din(new_net_4915),
		.dout(new_net_1236)
	);

	bfr new_net_4916_bfr_before (
		.din(new_net_4916),
		.dout(new_net_4915)
	);

	bfr new_net_4917_bfr_before (
		.din(new_net_4917),
		.dout(new_net_4916)
	);

	bfr new_net_4918_bfr_before (
		.din(new_net_4918),
		.dout(new_net_4917)
	);

	spl2 _0299__v_fanout (
		.a(_0299_),
		.b(new_net_1235),
		.c(new_net_4918)
	);

	bfr new_net_4919_bfr_before (
		.din(new_net_4919),
		.dout(new_net_557)
	);

	bfr new_net_4920_bfr_before (
		.din(new_net_4920),
		.dout(new_net_4919)
	);

	bfr new_net_4921_bfr_before (
		.din(new_net_4921),
		.dout(new_net_4920)
	);

	bfr new_net_4922_bfr_before (
		.din(new_net_4922),
		.dout(new_net_4921)
	);

	spl2 _1666__v_fanout (
		.a(_1666_),
		.b(new_net_556),
		.c(new_net_4922)
	);

	bfr new_net_4923_bfr_before (
		.din(new_net_4923),
		.dout(new_net_1544)
	);

	bfr new_net_4924_bfr_before (
		.din(new_net_4924),
		.dout(new_net_4923)
	);

	bfr new_net_4925_bfr_before (
		.din(new_net_4925),
		.dout(new_net_4924)
	);

	bfr new_net_4926_bfr_before (
		.din(new_net_4926),
		.dout(new_net_4925)
	);

	spl2 _1784__v_fanout (
		.a(_1784_),
		.b(new_net_1543),
		.c(new_net_4926)
	);

	spl2 _0900__v_fanout (
		.a(_0900_),
		.b(new_net_1996),
		.c(new_net_1997)
	);

	bfr new_net_4927_bfr_before (
		.din(new_net_4927),
		.dout(new_net_973)
	);

	bfr new_net_4928_bfr_before (
		.din(new_net_4928),
		.dout(new_net_4927)
	);

	bfr new_net_4929_bfr_before (
		.din(new_net_4929),
		.dout(new_net_4928)
	);

	bfr new_net_4930_bfr_before (
		.din(new_net_4930),
		.dout(new_net_4929)
	);

	spl2 _0501__v_fanout (
		.a(_0501_),
		.b(new_net_972),
		.c(new_net_4930)
	);

	bfr new_net_4931_bfr_after (
		.din(_0939_),
		.dout(new_net_4931)
	);

	bfr new_net_4932_bfr_after (
		.din(new_net_4931),
		.dout(new_net_4932)
	);

	bfr new_net_4933_bfr_after (
		.din(new_net_4932),
		.dout(new_net_4933)
	);

	bfr new_net_4934_bfr_after (
		.din(new_net_4933),
		.dout(new_net_4934)
	);

	spl2 _0939__v_fanout (
		.a(new_net_4934),
		.b(new_net_1772),
		.c(new_net_1773)
	);

	bfr new_net_4935_bfr_before (
		.din(new_net_4935),
		.dout(new_net_1143)
	);

	bfr new_net_4936_bfr_before (
		.din(new_net_4936),
		.dout(new_net_4935)
	);

	bfr new_net_4937_bfr_before (
		.din(new_net_4937),
		.dout(new_net_4936)
	);

	bfr new_net_4938_bfr_before (
		.din(new_net_4938),
		.dout(new_net_4937)
	);

	spl2 _0801__v_fanout (
		.a(_0801_),
		.b(new_net_1142),
		.c(new_net_4938)
	);

	bfr new_net_4939_bfr_before (
		.din(new_net_4939),
		.dout(new_net_91)
	);

	bfr new_net_4940_bfr_before (
		.din(new_net_4940),
		.dout(new_net_4939)
	);

	bfr new_net_4941_bfr_before (
		.din(new_net_4941),
		.dout(new_net_4940)
	);

	bfr new_net_4942_bfr_before (
		.din(new_net_4942),
		.dout(new_net_4941)
	);

	spl2 _0180__v_fanout (
		.a(_0180_),
		.b(new_net_90),
		.c(new_net_4942)
	);

	bfr new_net_4943_bfr_before (
		.din(new_net_4943),
		.dout(new_net_1205)
	);

	bfr new_net_4944_bfr_before (
		.din(new_net_4944),
		.dout(new_net_4943)
	);

	bfr new_net_4945_bfr_before (
		.din(new_net_4945),
		.dout(new_net_4944)
	);

	bfr new_net_4946_bfr_before (
		.din(new_net_4946),
		.dout(new_net_4945)
	);

	spl2 _0064__v_fanout (
		.a(_0064_),
		.b(new_net_1204),
		.c(new_net_4946)
	);

	spl2 _0965__v_fanout (
		.a(_0965_),
		.b(new_net_2647),
		.c(new_net_2648)
	);

	bfr new_net_4947_bfr_before (
		.din(new_net_4947),
		.dout(new_net_1566)
	);

	bfr new_net_4948_bfr_before (
		.din(new_net_4948),
		.dout(new_net_4947)
	);

	bfr new_net_4949_bfr_before (
		.din(new_net_4949),
		.dout(new_net_4948)
	);

	bfr new_net_4950_bfr_before (
		.din(new_net_4950),
		.dout(new_net_4949)
	);

	spl2 _0854__v_fanout (
		.a(_0854_),
		.b(new_net_1565),
		.c(new_net_4950)
	);

	bfr new_net_4951_bfr_before (
		.din(new_net_4951),
		.dout(new_net_1821)
	);

	bfr new_net_4952_bfr_before (
		.din(new_net_4952),
		.dout(new_net_4951)
	);

	bfr new_net_4953_bfr_before (
		.din(new_net_4953),
		.dout(new_net_4952)
	);

	bfr new_net_4954_bfr_before (
		.din(new_net_4954),
		.dout(new_net_4953)
	);

	spl2 _0739__v_fanout (
		.a(_0739_),
		.b(new_net_1820),
		.c(new_net_4954)
	);

	bfr new_net_4955_bfr_before (
		.din(new_net_4955),
		.dout(new_net_3202)
	);

	bfr new_net_4956_bfr_before (
		.din(new_net_4956),
		.dout(new_net_4955)
	);

	bfr new_net_4957_bfr_before (
		.din(new_net_4957),
		.dout(new_net_4956)
	);

	bfr new_net_4958_bfr_before (
		.din(new_net_4958),
		.dout(new_net_4957)
	);

	spl2 _1554__v_fanout (
		.a(_1554_),
		.b(new_net_3201),
		.c(new_net_4958)
	);

	bfr new_net_4959_bfr_before (
		.din(new_net_4959),
		.dout(new_net_2990)
	);

	bfr new_net_4960_bfr_before (
		.din(new_net_4960),
		.dout(new_net_4959)
	);

	bfr new_net_4961_bfr_before (
		.din(new_net_4961),
		.dout(new_net_4960)
	);

	bfr new_net_4962_bfr_before (
		.din(new_net_4962),
		.dout(new_net_4961)
	);

	spl2 _0404__v_fanout (
		.a(_0404_),
		.b(new_net_2989),
		.c(new_net_4962)
	);

	bfr new_net_4963_bfr_before (
		.din(new_net_4963),
		.dout(new_net_2721)
	);

	bfr new_net_4964_bfr_before (
		.din(new_net_4964),
		.dout(new_net_4963)
	);

	bfr new_net_4965_bfr_before (
		.din(new_net_4965),
		.dout(new_net_4964)
	);

	bfr new_net_4966_bfr_before (
		.din(new_net_4966),
		.dout(new_net_4965)
	);

	spl2 _0589__v_fanout (
		.a(_0589_),
		.b(new_net_2720),
		.c(new_net_4966)
	);

	spl2 _0668__v_fanout (
		.a(_0668_),
		.b(new_net_936),
		.c(new_net_937)
	);

	spl2 _0298__v_fanout (
		.a(_0298_),
		.b(new_net_1064),
		.c(new_net_1065)
	);

	spl2 _0179__v_fanout (
		.a(_0179_),
		.b(new_net_3163),
		.c(new_net_3164)
	);

	spl2 _0332__v_fanout (
		.a(_0332_),
		.b(new_net_944),
		.c(new_net_945)
	);

	spl2 _0534__v_fanout (
		.a(_0534_),
		.b(new_net_2196),
		.c(new_net_2197)
	);

	spl2 _1683__v_fanout (
		.a(_1683_),
		.b(new_net_1148),
		.c(new_net_1149)
	);

	bfr new_net_4967_bfr_before (
		.din(new_net_4967),
		.dout(new_net_101)
	);

	bfr new_net_4968_bfr_before (
		.din(new_net_4968),
		.dout(new_net_4967)
	);

	bfr new_net_4969_bfr_before (
		.din(new_net_4969),
		.dout(new_net_4968)
	);

	bfr new_net_4970_bfr_before (
		.din(new_net_4970),
		.dout(new_net_4969)
	);

	spl2 _0898__v_fanout (
		.a(_0898_),
		.b(new_net_100),
		.c(new_net_4970)
	);

	spl2 _0834__v_fanout (
		.a(_0834_),
		.b(new_net_2434),
		.c(new_net_2435)
	);

	spl2 _1808__v_fanout (
		.a(_1808_),
		.b(new_net_2847),
		.c(new_net_2848)
	);

	spl2 _1553__v_fanout (
		.a(_1553_),
		.b(new_net_2641),
		.c(new_net_2642)
	);

	spl2 _0772__v_fanout (
		.a(_0772_),
		.b(new_net_1136),
		.c(new_net_1137)
	);

	spl2 _1783__v_fanout (
		.a(_1783_),
		.b(new_net_1322),
		.c(new_net_1323)
	);

	spl2 _0800__v_fanout (
		.a(_0800_),
		.b(new_net_1102),
		.c(new_net_1103)
	);

	spl2 _1664__v_fanout (
		.a(_1664_),
		.b(new_net_2242),
		.c(new_net_2243)
	);

	spl2 _0588__v_fanout (
		.a(_0588_),
		.b(new_net_1010),
		.c(new_net_1011)
	);

	spl2 _0063__v_fanout (
		.a(_0063_),
		.b(new_net_1042),
		.c(new_net_1043)
	);

	spl2 _1563__v_fanout (
		.a(_1563_),
		.b(new_net_1626),
		.c(new_net_1627)
	);

	spl2 _0403__v_fanout (
		.a(_0403_),
		.b(new_net_2765),
		.c(new_net_2766)
	);

	spl2 _0622__v_fanout (
		.a(_0622_),
		.b(new_net_78),
		.c(new_net_79)
	);

	spl2 _0738__v_fanout (
		.a(_0738_),
		.b(new_net_1662),
		.c(new_net_1663)
	);

	spl2 _0090__v_fanout (
		.a(_0090_),
		.b(new_net_2927),
		.c(new_net_2928)
	);

	spl2 _0702__v_fanout (
		.a(_0702_),
		.b(new_net_2734),
		.c(new_net_2735)
	);

	spl2 _0438__v_fanout (
		.a(_0438_),
		.b(new_net_789),
		.c(new_net_790)
	);

	spl2 _1453__v_fanout (
		.a(_1453_),
		.b(new_net_1658),
		.c(new_net_1659)
	);

	spl2 _0500__v_fanout (
		.a(_0500_),
		.b(new_net_3073),
		.c(new_net_3074)
	);

	spl2 _0937__v_fanout (
		.a(_0937_),
		.b(new_net_2470),
		.c(new_net_2471)
	);

	spl2 _0217__v_fanout (
		.a(_0217_),
		.b(new_net_2955),
		.c(new_net_2956)
	);

	spl2 _0935__v_fanout (
		.a(_0935_),
		.b(new_net_1489),
		.c(new_net_1490)
	);

	spl2 _0586__v_fanout (
		.a(_0586_),
		.b(new_net_2587),
		.c(new_net_2588)
	);

	spl2 _0177__v_fanout (
		.a(_0177_),
		.b(new_net_3047),
		.c(new_net_3048)
	);

	spl2 _0665__v_fanout (
		.a(_0665_),
		.b(new_net_144),
		.c(new_net_145)
	);

	spl2 _0061__v_fanout (
		.a(_0061_),
		.b(new_net_691),
		.c(new_net_692)
	);

	spl2 _0887__v_fanout (
		.a(_0887_),
		.b(new_net_1348),
		.c(new_net_1349)
	);

	spl2 _1450__v_fanout (
		.a(_1450_),
		.b(new_net_1068),
		.c(new_net_1069)
	);

	spl2 _1662__v_fanout (
		.a(_1662_),
		.b(new_net_372),
		.c(new_net_373)
	);

	spl2 _0798__v_fanout (
		.a(_0798_),
		.b(new_net_2886),
		.c(new_net_2887)
	);

	spl2 _0736__v_fanout (
		.a(_0736_),
		.b(new_net_313),
		.c(new_net_314)
	);

	spl2 _0498__v_fanout (
		.a(_0498_),
		.b(new_net_2657),
		.c(new_net_2658)
	);

	spl2 _0401__v_fanout (
		.a(_0401_),
		.b(new_net_2380),
		.c(new_net_2381)
	);

	bfr new_net_4971_bfr_after (
		.din(_0853_),
		.dout(new_net_4971)
	);

	bfr new_net_4972_bfr_after (
		.din(new_net_4971),
		.dout(new_net_4972)
	);

	spl2 _0853__v_fanout (
		.a(new_net_4972),
		.b(new_net_2579),
		.c(new_net_2580)
	);

	spl2 _1781__v_fanout (
		.a(_1781_),
		.b(new_net_124),
		.c(new_net_125)
	);

	spl2 _0295__v_fanout (
		.a(_0295_),
		.b(new_net_2726),
		.c(new_net_2727)
	);

	spl2 _1551__v_fanout (
		.a(_1551_),
		.b(new_net_2569),
		.c(new_net_2570)
	);

	bfr new_net_4973_bfr_before (
		.din(new_net_4973),
		.dout(new_net_1827)
	);

	bfr new_net_4974_bfr_before (
		.din(new_net_4974),
		.dout(new_net_4973)
	);

	bfr new_net_4975_bfr_before (
		.din(new_net_4975),
		.dout(new_net_4974)
	);

	bfr new_net_4976_bfr_before (
		.din(new_net_4976),
		.dout(new_net_4975)
	);

	spl2 _0933__v_fanout (
		.a(_0933_),
		.b(new_net_1826),
		.c(new_net_4976)
	);

	spl2 _0175__v_fanout (
		.a(_0175_),
		.b(new_net_2971),
		.c(new_net_2972)
	);

	spl2 _0735__v_fanout (
		.a(_0735_),
		.b(new_net_1088),
		.c(new_net_1089)
	);

	spl2 _0400__v_fanout (
		.a(_0400_),
		.b(new_net_2178),
		.c(new_net_2179)
	);

	spl2 _0585__v_fanout (
		.a(_0585_),
		.b(new_net_462),
		.c(new_net_463)
	);

	spl2 _1661__v_fanout (
		.a(_1661_),
		.b(new_net_331),
		.c(new_net_332)
	);

	spl2 _0664__v_fanout (
		.a(_0664_),
		.b(new_net_3272),
		.c(new_net_3273)
	);

	spl2 _0497__v_fanout (
		.a(_0497_),
		.b(new_net_846),
		.c(new_net_847)
	);

	spl2 _0060__v_fanout (
		.a(_0060_),
		.b(new_net_1732),
		.c(new_net_1733)
	);

	spl2 _0797__v_fanout (
		.a(_0797_),
		.b(new_net_2685),
		.c(new_net_2686)
	);

	spl2 _1780__v_fanout (
		.a(_1780_),
		.b(new_net_828),
		.c(new_net_829)
	);

	spl2 _0851__v_fanout (
		.a(_0851_),
		.b(new_net_2176),
		.c(new_net_2177)
	);

	spl2 _1449__v_fanout (
		.a(_1449_),
		.b(new_net_277),
		.c(new_net_278)
	);

	spl2 _0294__v_fanout (
		.a(_0294_),
		.b(new_net_317),
		.c(new_net_318)
	);

	spl2 _1550__v_fanout (
		.a(_1550_),
		.b(new_net_2509),
		.c(new_net_2510)
	);

	bfr new_net_4977_bfr_before (
		.din(new_net_4977),
		.dout(new_net_1301)
	);

	bfr new_net_4978_bfr_before (
		.din(new_net_4978),
		.dout(new_net_4977)
	);

	bfr new_net_4979_bfr_before (
		.din(new_net_4979),
		.dout(new_net_4978)
	);

	bfr new_net_4980_bfr_before (
		.din(new_net_4980),
		.dout(new_net_4979)
	);

	spl2 _1659__v_fanout (
		.a(_1659_),
		.b(new_net_1300),
		.c(new_net_4980)
	);

	bfr new_net_4981_bfr_after (
		.din(_0897_),
		.dout(new_net_4981)
	);

	bfr new_net_4982_bfr_after (
		.din(new_net_4981),
		.dout(new_net_4982)
	);

	bfr new_net_4983_bfr_after (
		.din(new_net_4982),
		.dout(new_net_4983)
	);

	bfr new_net_4984_bfr_after (
		.din(new_net_4983),
		.dout(new_net_4984)
	);

	spl2 _0897__v_fanout (
		.a(new_net_4984),
		.b(new_net_1497),
		.c(new_net_1498)
	);

	bfr new_net_4985_bfr_before (
		.din(new_net_4985),
		.dout(new_net_2457)
	);

	bfr new_net_4986_bfr_before (
		.din(new_net_4986),
		.dout(new_net_4985)
	);

	bfr new_net_4987_bfr_before (
		.din(new_net_4987),
		.dout(new_net_4986)
	);

	bfr new_net_4988_bfr_before (
		.din(new_net_4988),
		.dout(new_net_4987)
	);

	spl2 _0583__v_fanout (
		.a(_0583_),
		.b(new_net_2456),
		.c(new_net_4988)
	);

	bfr new_net_4989_bfr_before (
		.din(new_net_4989),
		.dout(new_net_1955)
	);

	bfr new_net_4990_bfr_before (
		.din(new_net_4990),
		.dout(new_net_4989)
	);

	bfr new_net_4991_bfr_before (
		.din(new_net_4991),
		.dout(new_net_4990)
	);

	bfr new_net_4992_bfr_before (
		.din(new_net_4992),
		.dout(new_net_4991)
	);

	spl2 _1548__v_fanout (
		.a(_1548_),
		.b(new_net_1954),
		.c(new_net_4992)
	);

	bfr new_net_4993_bfr_before (
		.din(new_net_4993),
		.dout(new_net_780)
	);

	bfr new_net_4994_bfr_before (
		.din(new_net_4994),
		.dout(new_net_4993)
	);

	bfr new_net_4995_bfr_before (
		.din(new_net_4995),
		.dout(new_net_4994)
	);

	bfr new_net_4996_bfr_before (
		.din(new_net_4996),
		.dout(new_net_4995)
	);

	spl2 _0733__v_fanout (
		.a(_0733_),
		.b(new_net_779),
		.c(new_net_4996)
	);

	bfr new_net_4997_bfr_before (
		.din(new_net_4997),
		.dout(new_net_29)
	);

	bfr new_net_4998_bfr_before (
		.din(new_net_4998),
		.dout(new_net_4997)
	);

	bfr new_net_4999_bfr_before (
		.din(new_net_4999),
		.dout(new_net_4998)
	);

	bfr new_net_5000_bfr_before (
		.din(new_net_5000),
		.dout(new_net_4999)
	);

	spl2 _1778__v_fanout (
		.a(_1778_),
		.b(new_net_28),
		.c(new_net_5000)
	);

	bfr new_net_5001_bfr_before (
		.din(new_net_5001),
		.dout(new_net_3225)
	);

	bfr new_net_5002_bfr_before (
		.din(new_net_5002),
		.dout(new_net_5001)
	);

	bfr new_net_5003_bfr_before (
		.din(new_net_5003),
		.dout(new_net_5002)
	);

	bfr new_net_5004_bfr_before (
		.din(new_net_5004),
		.dout(new_net_5003)
	);

	spl2 _0292__v_fanout (
		.a(_0292_),
		.b(new_net_3224),
		.c(new_net_5004)
	);

	spl2 _0932__v_fanout (
		.a(_0932_),
		.b(new_net_1666),
		.c(new_net_1667)
	);

	spl2 _0849__v_fanout (
		.a(_0849_),
		.b(new_net_3053),
		.c(new_net_3054)
	);

	bfr new_net_5005_bfr_before (
		.din(new_net_5005),
		.dout(new_net_2035)
	);

	bfr new_net_5006_bfr_before (
		.din(new_net_5006),
		.dout(new_net_5005)
	);

	bfr new_net_5007_bfr_before (
		.din(new_net_5007),
		.dout(new_net_5006)
	);

	bfr new_net_5008_bfr_before (
		.din(new_net_5008),
		.dout(new_net_5007)
	);

	spl2 _0495__v_fanout (
		.a(_0495_),
		.b(new_net_2034),
		.c(new_net_5008)
	);

	bfr new_net_5009_bfr_before (
		.din(new_net_5009),
		.dout(new_net_702)
	);

	bfr new_net_5010_bfr_before (
		.din(new_net_5010),
		.dout(new_net_5009)
	);

	bfr new_net_5011_bfr_before (
		.din(new_net_5011),
		.dout(new_net_5010)
	);

	bfr new_net_5012_bfr_before (
		.din(new_net_5012),
		.dout(new_net_5011)
	);

	spl2 _0662__v_fanout (
		.a(_0662_),
		.b(new_net_701),
		.c(new_net_5012)
	);

	bfr new_net_5013_bfr_before (
		.din(new_net_5013),
		.dout(new_net_2091)
	);

	bfr new_net_5014_bfr_before (
		.din(new_net_5014),
		.dout(new_net_5013)
	);

	bfr new_net_5015_bfr_before (
		.din(new_net_5015),
		.dout(new_net_5014)
	);

	bfr new_net_5016_bfr_before (
		.din(new_net_5016),
		.dout(new_net_5015)
	);

	spl2 _0794__v_fanout (
		.a(_0794_),
		.b(new_net_2090),
		.c(new_net_5016)
	);

	bfr new_net_5017_bfr_before (
		.din(new_net_5017),
		.dout(new_net_229)
	);

	bfr new_net_5018_bfr_before (
		.din(new_net_5018),
		.dout(new_net_5017)
	);

	bfr new_net_5019_bfr_before (
		.din(new_net_5019),
		.dout(new_net_5018)
	);

	bfr new_net_5020_bfr_before (
		.din(new_net_5020),
		.dout(new_net_5019)
	);

	spl2 _0398__v_fanout (
		.a(_0398_),
		.b(new_net_228),
		.c(new_net_5020)
	);

	bfr new_net_5021_bfr_before (
		.din(new_net_5021),
		.dout(new_net_2860)
	);

	bfr new_net_5022_bfr_before (
		.din(new_net_5022),
		.dout(new_net_5021)
	);

	bfr new_net_5023_bfr_before (
		.din(new_net_5023),
		.dout(new_net_5022)
	);

	bfr new_net_5024_bfr_before (
		.din(new_net_5024),
		.dout(new_net_5023)
	);

	spl2 _0173__v_fanout (
		.a(_0173_),
		.b(new_net_2859),
		.c(new_net_5024)
	);

	bfr new_net_5025_bfr_before (
		.din(new_net_5025),
		.dout(new_net_543)
	);

	bfr new_net_5026_bfr_before (
		.din(new_net_5026),
		.dout(new_net_5025)
	);

	bfr new_net_5027_bfr_before (
		.din(new_net_5027),
		.dout(new_net_5026)
	);

	bfr new_net_5028_bfr_before (
		.din(new_net_5028),
		.dout(new_net_5027)
	);

	spl2 _1447__v_fanout (
		.a(_1447_),
		.b(new_net_542),
		.c(new_net_5028)
	);

	bfr new_net_5029_bfr_before (
		.din(new_net_5029),
		.dout(new_net_1689)
	);

	bfr new_net_5030_bfr_before (
		.din(new_net_5030),
		.dout(new_net_5029)
	);

	bfr new_net_5031_bfr_before (
		.din(new_net_5031),
		.dout(new_net_5030)
	);

	bfr new_net_5032_bfr_before (
		.din(new_net_5032),
		.dout(new_net_5031)
	);

	spl2 _0058__v_fanout (
		.a(_0058_),
		.b(new_net_1688),
		.c(new_net_5032)
	);

	spl2 _1810__v_fanout (
		.a(_1810_),
		.b(new_net_1172),
		.c(new_net_1173)
	);

	spl2 _1455__v_fanout (
		.a(_1455_),
		.b(new_net_1994),
		.c(new_net_1995)
	);

	spl2 _1446__v_fanout (
		.a(_1446_),
		.b(new_net_178),
		.c(new_net_179)
	);

	spl2 _0172__v_fanout (
		.a(_0172_),
		.b(new_net_2805),
		.c(new_net_2806)
	);

	spl2 _0440__v_fanout (
		.a(_0440_),
		.b(new_net_230),
		.c(new_net_231)
	);

	spl2 _0291__v_fanout (
		.a(_0291_),
		.b(new_net_2539),
		.c(new_net_2540)
	);

	spl2 _1565__v_fanout (
		.a(_1565_),
		.b(new_net_3149),
		.c(new_net_3150)
	);

	spl2 _0057__v_fanout (
		.a(_0057_),
		.b(new_net_3209),
		.c(new_net_3210)
	);

	spl2 _0397__v_fanout (
		.a(_0397_),
		.b(new_net_216),
		.c(new_net_217)
	);

	spl2 _1685__v_fanout (
		.a(_1685_),
		.b(new_net_1218),
		.c(new_net_1219)
	);

	spl2 _0494__v_fanout (
		.a(_0494_),
		.b(new_net_1858),
		.c(new_net_1859)
	);

	spl2 _0895__v_fanout (
		.a(_0895_),
		.b(new_net_3260),
		.c(new_net_3261)
	);

	spl2 _0661__v_fanout (
		.a(_0661_),
		.b(new_net_2603),
		.c(new_net_2604)
	);

	spl2 _0220__v_fanout (
		.a(_0220_),
		.b(new_net_3171),
		.c(new_net_3172)
	);

	spl2 _1547__v_fanout (
		.a(_1547_),
		.b(new_net_2394),
		.c(new_net_2395)
	);

	spl2 _0624__v_fanout (
		.a(_0624_),
		.b(new_net_452),
		.c(new_net_453)
	);

	spl2 _1362__v_fanout (
		.a(_1362_),
		.b(new_net_1730),
		.c(new_net_1731)
	);

	spl2 _0775__v_fanout (
		.a(_0775_),
		.b(new_net_1712),
		.c(new_net_1713)
	);

	spl2 _0092__v_fanout (
		.a(_0092_),
		.b(new_net_134),
		.c(new_net_135)
	);

	spl2 _0732__v_fanout (
		.a(_0732_),
		.b(new_net_572),
		.c(new_net_573)
	);

	spl2 _0537__v_fanout (
		.a(_0537_),
		.b(new_net_2302),
		.c(new_net_2303)
	);

	spl2 _1777__v_fanout (
		.a(_1777_),
		.b(new_net_3137),
		.c(new_net_3138)
	);

	spl2 _0582__v_fanout (
		.a(_0582_),
		.b(new_net_2436),
		.c(new_net_2437)
	);

	spl2 _1658__v_fanout (
		.a(_1658_),
		.b(new_net_1094),
		.c(new_net_1095)
	);

	spl2 _0704__v_fanout (
		.a(_0704_),
		.b(new_net_705),
		.c(new_net_706)
	);

	spl2 _0334__v_fanout (
		.a(_0334_),
		.b(new_net_996),
		.c(new_net_997)
	);

	bfr new_net_5033_bfr_before (
		.din(new_net_5033),
		.dout(new_net_1434)
	);

	bfr new_net_5034_bfr_before (
		.din(new_net_5034),
		.dout(new_net_5033)
	);

	bfr new_net_5035_bfr_before (
		.din(new_net_5035),
		.dout(new_net_5034)
	);

	bfr new_net_5036_bfr_before (
		.din(new_net_5036),
		.dout(new_net_5035)
	);

	spl2 _0847__v_fanout (
		.a(_0847_),
		.b(new_net_1433),
		.c(new_net_5036)
	);

	spl2 _0894__v_fanout (
		.a(_0894_),
		.b(new_net_2687),
		.c(new_net_2688)
	);

	spl2 _1656__v_fanout (
		.a(_1656_),
		.b(new_net_791),
		.c(new_net_792)
	);

	spl2 _0836__v_fanout (
		.a(_0836_),
		.b(new_net_2488),
		.c(new_net_2489)
	);

	spl2 _0491__v_fanout (
		.a(_0491_),
		.b(new_net_604),
		.c(new_net_605)
	);

	spl2 _1545__v_fanout (
		.a(_1545_),
		.b(new_net_2307),
		.c(new_net_2308)
	);

	spl2 _0170__v_fanout (
		.a(_0170_),
		.b(new_net_1366),
		.c(new_net_1367)
	);

	spl2 _0054__v_fanout (
		.a(_0054_),
		.b(new_net_2748),
		.c(new_net_2749)
	);

	bfr new_net_5037_bfr_after (
		.din(_0793_),
		.dout(new_net_5037)
	);

	bfr new_net_5038_bfr_after (
		.din(new_net_5037),
		.dout(new_net_5038)
	);

	spl2 _0793__v_fanout (
		.a(new_net_5038),
		.b(new_net_904),
		.c(new_net_905)
	);

	spl2 _1359__v_fanout (
		.a(_1359_),
		.b(new_net_2651),
		.c(new_net_2652)
	);

	spl2 _0395__v_fanout (
		.a(_0395_),
		.b(new_net_1226),
		.c(new_net_1227)
	);

	spl2 _0659__v_fanout (
		.a(_0659_),
		.b(new_net_2202),
		.c(new_net_2203)
	);

	spl2 _0289__v_fanout (
		.a(_0289_),
		.b(new_net_2462),
		.c(new_net_2463)
	);

	spl2 _1444__v_fanout (
		.a(_1444_),
		.b(new_net_104),
		.c(new_net_105)
	);

	spl2 _1775__v_fanout (
		.a(_1775_),
		.b(new_net_3145),
		.c(new_net_3146)
	);

	spl2 _0729__v_fanout (
		.a(_0729_),
		.b(new_net_62),
		.c(new_net_63)
	);

	spl2 _0580__v_fanout (
		.a(_0580_),
		.b(new_net_2368),
		.c(new_net_2369)
	);

	spl2 _0658__v_fanout (
		.a(_0658_),
		.b(new_net_1988),
		.c(new_net_1989)
	);

	spl2 _0791__v_fanout (
		.a(_0791_),
		.b(new_net_850),
		.c(new_net_851)
	);

	spl2 _0578__v_fanout (
		.a(_0578_),
		.b(new_net_2270),
		.c(new_net_2271)
	);

	spl2 _1655__v_fanout (
		.a(_1655_),
		.b(new_net_578),
		.c(new_net_579)
	);

	spl2 _0053__v_fanout (
		.a(_0053_),
		.b(new_net_2527),
		.c(new_net_2528)
	);

	spl2 _1443__v_fanout (
		.a(_1443_),
		.b(new_net_3027),
		.c(new_net_3028)
	);

	spl2 _0490__v_fanout (
		.a(_0490_),
		.b(new_net_1098),
		.c(new_net_1099)
	);

	spl2 _0288__v_fanout (
		.a(_0288_),
		.b(new_net_2426),
		.c(new_net_2427)
	);

	spl2 _1773__v_fanout (
		.a(_1773_),
		.b(new_net_2286),
		.c(new_net_2287)
	);

	spl2 _1544__v_fanout (
		.a(_1544_),
		.b(new_net_2264),
		.c(new_net_2265)
	);

	spl2 _0393__v_fanout (
		.a(_0393_),
		.b(new_net_908),
		.c(new_net_909)
	);

	spl2 _0728__v_fanout (
		.a(_0728_),
		.b(new_net_34),
		.c(new_net_35)
	);

	spl2 _0169__v_fanout (
		.a(_0169_),
		.b(new_net_2718),
		.c(new_net_2719)
	);

	bfr new_net_5039_bfr_before (
		.din(new_net_5039),
		.dout(new_net_2095)
	);

	bfr new_net_5040_bfr_before (
		.din(new_net_5040),
		.dout(new_net_5039)
	);

	bfr new_net_5041_bfr_before (
		.din(new_net_5041),
		.dout(new_net_5040)
	);

	bfr new_net_5042_bfr_before (
		.din(new_net_5042),
		.dout(new_net_5041)
	);

	spl2 _0891__v_fanout (
		.a(_0891_),
		.b(new_net_2094),
		.c(new_net_5042)
	);

	spl2 _1358__v_fanout (
		.a(_1358_),
		.b(new_net_1610),
		.c(new_net_1611)
	);

	bfr new_net_5043_bfr_before (
		.din(new_net_5043),
		.dout(new_net_1905)
	);

	bfr new_net_5044_bfr_before (
		.din(new_net_5044),
		.dout(new_net_5043)
	);

	bfr new_net_5045_bfr_before (
		.din(new_net_5045),
		.dout(new_net_5044)
	);

	bfr new_net_5046_bfr_before (
		.din(new_net_5046),
		.dout(new_net_5045)
	);

	spl2 _1771__v_fanout (
		.a(_1771_),
		.b(new_net_1904),
		.c(new_net_5046)
	);

	bfr new_net_5047_bfr_before (
		.din(new_net_5047),
		.dout(new_net_2640)
	);

	bfr new_net_5048_bfr_before (
		.din(new_net_5048),
		.dout(new_net_5047)
	);

	bfr new_net_5049_bfr_before (
		.din(new_net_5049),
		.dout(new_net_5048)
	);

	bfr new_net_5050_bfr_before (
		.din(new_net_5050),
		.dout(new_net_5049)
	);

	spl2 _0167__v_fanout (
		.a(_0167_),
		.b(new_net_2639),
		.c(new_net_5050)
	);

	bfr new_net_5051_bfr_before (
		.din(new_net_5051),
		.dout(new_net_2371)
	);

	bfr new_net_5052_bfr_before (
		.din(new_net_5052),
		.dout(new_net_5051)
	);

	bfr new_net_5053_bfr_before (
		.din(new_net_5053),
		.dout(new_net_5052)
	);

	bfr new_net_5054_bfr_before (
		.din(new_net_5054),
		.dout(new_net_5053)
	);

	spl2 _0286__v_fanout (
		.a(_0286_),
		.b(new_net_2370),
		.c(new_net_5054)
	);

	bfr new_net_5055_bfr_before (
		.din(new_net_5055),
		.dout(new_net_3259)
	);

	bfr new_net_5056_bfr_before (
		.din(new_net_5056),
		.dout(new_net_5055)
	);

	bfr new_net_5057_bfr_before (
		.din(new_net_5057),
		.dout(new_net_5056)
	);

	bfr new_net_5058_bfr_before (
		.din(new_net_5058),
		.dout(new_net_5057)
	);

	spl2 _1441__v_fanout (
		.a(_1441_),
		.b(new_net_3258),
		.c(new_net_5058)
	);

	bfr new_net_5059_bfr_before (
		.din(new_net_5059),
		.dout(new_net_1572)
	);

	bfr new_net_5060_bfr_before (
		.din(new_net_5060),
		.dout(new_net_5059)
	);

	bfr new_net_5061_bfr_before (
		.din(new_net_5061),
		.dout(new_net_5060)
	);

	bfr new_net_5062_bfr_before (
		.din(new_net_5062),
		.dout(new_net_5061)
	);

	spl2 _0391__v_fanout (
		.a(_0391_),
		.b(new_net_1571),
		.c(new_net_5062)
	);

	bfr new_net_5063_bfr_before (
		.din(new_net_5063),
		.dout(new_net_1536)
	);

	bfr new_net_5064_bfr_before (
		.din(new_net_5064),
		.dout(new_net_5063)
	);

	bfr new_net_5065_bfr_before (
		.din(new_net_5065),
		.dout(new_net_5064)
	);

	bfr new_net_5066_bfr_before (
		.din(new_net_5066),
		.dout(new_net_5065)
	);

	spl2 _1356__v_fanout (
		.a(_1356_),
		.b(new_net_1535),
		.c(new_net_5066)
	);

	bfr new_net_5067_bfr_before (
		.din(new_net_5067),
		.dout(new_net_1655)
	);

	bfr new_net_5068_bfr_before (
		.din(new_net_5068),
		.dout(new_net_5067)
	);

	bfr new_net_5069_bfr_before (
		.din(new_net_5069),
		.dout(new_net_5068)
	);

	bfr new_net_5070_bfr_before (
		.din(new_net_5070),
		.dout(new_net_5069)
	);

	spl2 _0656__v_fanout (
		.a(_0656_),
		.b(new_net_1654),
		.c(new_net_5070)
	);

	bfr new_net_5071_bfr_after (
		.din(_0846_),
		.dout(new_net_5071)
	);

	bfr new_net_5072_bfr_after (
		.din(new_net_5071),
		.dout(new_net_5072)
	);

	bfr new_net_5073_bfr_after (
		.din(new_net_5072),
		.dout(new_net_5073)
	);

	bfr new_net_5074_bfr_after (
		.din(new_net_5073),
		.dout(new_net_5074)
	);

	spl2 _0846__v_fanout (
		.a(new_net_5074),
		.b(new_net_1224),
		.c(new_net_1225)
	);

	bfr new_net_5075_bfr_before (
		.din(new_net_5075),
		.dout(new_net_25)
	);

	bfr new_net_5076_bfr_before (
		.din(new_net_5076),
		.dout(new_net_5075)
	);

	bfr new_net_5077_bfr_before (
		.din(new_net_5077),
		.dout(new_net_5076)
	);

	bfr new_net_5078_bfr_before (
		.din(new_net_5078),
		.dout(new_net_5077)
	);

	spl2 _1652__v_fanout (
		.a(_1652_),
		.b(new_net_24),
		.c(new_net_5078)
	);

	spl2 _0790__v_fanout (
		.a(_0790_),
		.b(new_net_2571),
		.c(new_net_2572)
	);

	spl2 _0890__v_fanout (
		.a(_0890_),
		.b(new_net_2997),
		.c(new_net_2998)
	);

	bfr new_net_5079_bfr_before (
		.din(new_net_5079),
		.dout(new_net_804)
	);

	bfr new_net_5080_bfr_before (
		.din(new_net_5080),
		.dout(new_net_5079)
	);

	bfr new_net_5081_bfr_before (
		.din(new_net_5081),
		.dout(new_net_5080)
	);

	bfr new_net_5082_bfr_before (
		.din(new_net_5082),
		.dout(new_net_5081)
	);

	spl2 _0488__v_fanout (
		.a(_0488_),
		.b(new_net_803),
		.c(new_net_5082)
	);

	bfr new_net_5083_bfr_before (
		.din(new_net_5083),
		.dout(new_net_1379)
	);

	bfr new_net_5084_bfr_before (
		.din(new_net_5084),
		.dout(new_net_5083)
	);

	bfr new_net_5085_bfr_before (
		.din(new_net_5085),
		.dout(new_net_5084)
	);

	bfr new_net_5086_bfr_before (
		.din(new_net_5086),
		.dout(new_net_5085)
	);

	spl2 _0051__v_fanout (
		.a(_0051_),
		.b(new_net_1378),
		.c(new_net_5086)
	);

	bfr new_net_5087_bfr_before (
		.din(new_net_5087),
		.dout(new_net_1925)
	);

	bfr new_net_5088_bfr_before (
		.din(new_net_5088),
		.dout(new_net_5087)
	);

	bfr new_net_5089_bfr_before (
		.din(new_net_5089),
		.dout(new_net_5088)
	);

	bfr new_net_5090_bfr_before (
		.din(new_net_5090),
		.dout(new_net_5089)
	);

	spl2 _0576__v_fanout (
		.a(_0576_),
		.b(new_net_1924),
		.c(new_net_5090)
	);

	bfr new_net_5091_bfr_before (
		.din(new_net_5091),
		.dout(new_net_1526)
	);

	bfr new_net_5092_bfr_before (
		.din(new_net_5092),
		.dout(new_net_5091)
	);

	bfr new_net_5093_bfr_before (
		.din(new_net_5093),
		.dout(new_net_5092)
	);

	bfr new_net_5094_bfr_before (
		.din(new_net_5094),
		.dout(new_net_5093)
	);

	spl2 _0726__v_fanout (
		.a(_0726_),
		.b(new_net_1525),
		.c(new_net_5094)
	);

	bfr new_net_5095_bfr_before (
		.din(new_net_5095),
		.dout(new_net_2185)
	);

	bfr new_net_5096_bfr_before (
		.din(new_net_5096),
		.dout(new_net_5095)
	);

	bfr new_net_5097_bfr_before (
		.din(new_net_5097),
		.dout(new_net_5096)
	);

	bfr new_net_5098_bfr_before (
		.din(new_net_5098),
		.dout(new_net_5097)
	);

	spl2 _1542__v_fanout (
		.a(_1542_),
		.b(new_net_2184),
		.c(new_net_5098)
	);

	spl2 _0442__v_fanout (
		.a(_0442_),
		.b(new_net_1511),
		.c(new_net_1512)
	);

	spl2 _1279__v_fanout (
		.a(_1279_),
		.b(new_net_226),
		.c(new_net_227)
	);

	spl2 _1355__v_fanout (
		.a(_1355_),
		.b(new_net_960),
		.c(new_net_961)
	);

	spl2 _1812__v_fanout (
		.a(_1812_),
		.b(new_net_408),
		.c(new_net_409)
	);

	spl2 _1568__v_fanout (
		.a(_1568_),
		.b(new_net_1618),
		.c(new_net_1619)
	);

	spl2 _0336__v_fanout (
		.a(_0336_),
		.b(new_net_478),
		.c(new_net_479)
	);

	spl2 _1364__v_fanout (
		.a(_1364_),
		.b(new_net_1784),
		.c(new_net_1785)
	);

	spl2 _1440__v_fanout (
		.a(_1440_),
		.b(new_net_986),
		.c(new_net_987)
	);

	spl2 _1770__v_fanout (
		.a(_1770_),
		.b(new_net_1720),
		.c(new_net_1721)
	);

	spl2 _0166__v_fanout (
		.a(_0166_),
		.b(new_net_649),
		.c(new_net_650)
	);

	spl2 _0050__v_fanout (
		.a(_0050_),
		.b(new_net_1932),
		.c(new_net_1933)
	);

	spl2 _0487__v_fanout (
		.a(_0487_),
		.b(new_net_418),
		.c(new_net_419)
	);

	spl2 _0539__v_fanout (
		.a(_0539_),
		.b(new_net_1513),
		.c(new_net_1514)
	);

	spl2 _0284__v_fanout (
		.a(_0284_),
		.b(new_net_1636),
		.c(new_net_1637)
	);

	spl2 _0390__v_fanout (
		.a(_0390_),
		.b(new_net_323),
		.c(new_net_324)
	);

	spl2 _0575__v_fanout (
		.a(_0575_),
		.b(new_net_2154),
		.c(new_net_2155)
	);

	spl2 _0654__v_fanout (
		.a(_0654_),
		.b(new_net_1241),
		.c(new_net_1242)
	);

	spl2 _0844__v_fanout (
		.a(_0844_),
		.b(new_net_910),
		.c(new_net_911)
	);

	spl2 _1541__v_fanout (
		.a(_1541_),
		.b(new_net_677),
		.c(new_net_678)
	);

	spl2 _0706__v_fanout (
		.a(_0706_),
		.b(new_net_250),
		.c(new_net_251)
	);

	spl2 _0626__v_fanout (
		.a(_0626_),
		.b(new_net_934),
		.c(new_net_935)
	);

	spl2 _1688__v_fanout (
		.a(_1688_),
		.b(new_net_1344),
		.c(new_net_1345)
	);

	spl2 _1651__v_fanout (
		.a(_1651_),
		.b(new_net_1140),
		.c(new_net_1141)
	);

	spl2 _1457__v_fanout (
		.a(_1457_),
		.b(new_net_606),
		.c(new_net_607)
	);

	spl2 _0094__v_fanout (
		.a(_0094_),
		.b(new_net_516),
		.c(new_net_517)
	);

	bfr new_net_5099_bfr_before (
		.din(new_net_5099),
		.dout(new_net_696)
	);

	bfr new_net_5100_bfr_before (
		.din(new_net_5100),
		.dout(new_net_5099)
	);

	bfr new_net_5101_bfr_before (
		.din(new_net_5101),
		.dout(new_net_5100)
	);

	bfr new_net_5102_bfr_before (
		.din(new_net_5102),
		.dout(new_net_5101)
	);

	spl2 _0788__v_fanout (
		.a(_0788_),
		.b(new_net_695),
		.c(new_net_5102)
	);

	spl2 _0222__v_fanout (
		.a(_0222_),
		.b(new_net_3173),
		.c(new_net_3174)
	);

	spl2 _0388__v_fanout (
		.a(_0388_),
		.b(new_net_3268),
		.c(new_net_3269)
	);

	spl2 _0652__v_fanout (
		.a(_0652_),
		.b(new_net_914),
		.c(new_net_915)
	);

	spl2 _1276__v_fanout (
		.a(_1276_),
		.b(new_net_2882),
		.c(new_net_2883)
	);

	spl2 _0282__v_fanout (
		.a(_0282_),
		.b(new_net_2192),
		.c(new_net_2193)
	);

	spl2 _0777__v_fanout (
		.a(_0777_),
		.b(new_net_2082),
		.c(new_net_2083)
	);

	spl2 _1438__v_fanout (
		.a(_1438_),
		.b(new_net_612),
		.c(new_net_613)
	);

	spl2 _1539__v_fanout (
		.a(_1539_),
		.b(new_net_2068),
		.c(new_net_2069)
	);

	spl2 _1649__v_fanout (
		.a(_1649_),
		.b(new_net_3139),
		.c(new_net_3140)
	);

	spl2 _1768__v_fanout (
		.a(_1768_),
		.b(new_net_1354),
		.c(new_net_1355)
	);

	spl2 _0163__v_fanout (
		.a(_0163_),
		.b(new_net_2458),
		.c(new_net_2459)
	);

	spl2 _0048__v_fanout (
		.a(_0048_),
		.b(new_net_1606),
		.c(new_net_1607)
	);

	spl2 _0573__v_fanout (
		.a(_0573_),
		.b(new_net_2074),
		.c(new_net_2075)
	);

	bfr new_net_5103_bfr_after (
		.din(_0725_),
		.dout(new_net_5103)
	);

	bfr new_net_5104_bfr_after (
		.din(new_net_5103),
		.dout(new_net_5104)
	);

	spl2 _0725__v_fanout (
		.a(new_net_5104),
		.b(new_net_1487),
		.c(new_net_1488)
	);

	spl2 _0843__v_fanout (
		.a(_0843_),
		.b(new_net_715),
		.c(new_net_716)
	);

	spl2 _0485__v_fanout (
		.a(_0485_),
		.b(new_net_186),
		.c(new_net_187)
	);

	spl2 _1353__v_fanout (
		.a(_1353_),
		.b(new_net_1376),
		.c(new_net_1377)
	);

	spl2 _0651__v_fanout (
		.a(_0651_),
		.b(new_net_731),
		.c(new_net_732)
	);

	spl2 _0572__v_fanout (
		.a(_0572_),
		.b(new_net_1170),
		.c(new_net_1171)
	);

	spl2 _0162__v_fanout (
		.a(_0162_),
		.b(new_net_3159),
		.c(new_net_3160)
	);

	spl2 _0281__v_fanout (
		.a(_0281_),
		.b(new_net_2158),
		.c(new_net_2159)
	);

	spl2 _1767__v_fanout (
		.a(_1767_),
		.b(new_net_1166),
		.c(new_net_1167)
	);

	spl2 _1437__v_fanout (
		.a(_1437_),
		.b(new_net_3049),
		.c(new_net_3050)
	);

	spl2 _0484__v_fanout (
		.a(_0484_),
		.b(new_net_309),
		.c(new_net_310)
	);

	spl2 _0723__v_fanout (
		.a(_0723_),
		.b(new_net_252),
		.c(new_net_253)
	);

	spl2 _1538__v_fanout (
		.a(_1538_),
		.b(new_net_2008),
		.c(new_net_2009)
	);

	spl2 _1352__v_fanout (
		.a(_1352_),
		.b(new_net_354),
		.c(new_net_355)
	);

	spl2 _0047__v_fanout (
		.a(_0047_),
		.b(new_net_1386),
		.c(new_net_1387)
	);

	bfr new_net_5105_bfr_before (
		.din(new_net_5105),
		.dout(new_net_2725)
	);

	bfr new_net_5106_bfr_before (
		.din(new_net_5106),
		.dout(new_net_5105)
	);

	bfr new_net_5107_bfr_before (
		.din(new_net_5107),
		.dout(new_net_5106)
	);

	bfr new_net_5108_bfr_before (
		.din(new_net_5108),
		.dout(new_net_5107)
	);

	spl2 _0841__v_fanout (
		.a(_0841_),
		.b(new_net_2724),
		.c(new_net_5108)
	);

	spl2 _1275__v_fanout (
		.a(_1275_),
		.b(new_net_72),
		.c(new_net_73)
	);

	spl2 _0387__v_fanout (
		.a(_0387_),
		.b(new_net_3009),
		.c(new_net_3010)
	);

	spl2 _1648__v_fanout (
		.a(_1648_),
		.b(new_net_3121),
		.c(new_net_3122)
	);

	bfr new_net_5109_bfr_before (
		.din(new_net_5109),
		.dout(new_net_322)
	);

	bfr new_net_5110_bfr_before (
		.din(new_net_5110),
		.dout(new_net_5109)
	);

	bfr new_net_5111_bfr_before (
		.din(new_net_5111),
		.dout(new_net_5110)
	);

	bfr new_net_5112_bfr_before (
		.din(new_net_5112),
		.dout(new_net_5111)
	);

	spl2 _0649__v_fanout (
		.a(_0649_),
		.b(new_net_321),
		.c(new_net_5112)
	);

	spl2 _0722__v_fanout (
		.a(_0722_),
		.b(new_net_1334),
		.c(new_net_1335)
	);

	bfr new_net_5113_bfr_before (
		.din(new_net_5113),
		.dout(new_net_1317)
	);

	bfr new_net_5114_bfr_before (
		.din(new_net_5114),
		.dout(new_net_5113)
	);

	bfr new_net_5115_bfr_before (
		.din(new_net_5115),
		.dout(new_net_5114)
	);

	bfr new_net_5116_bfr_before (
		.din(new_net_5116),
		.dout(new_net_5115)
	);

	spl2 _0385__v_fanout (
		.a(_0385_),
		.b(new_net_1316),
		.c(new_net_5116)
	);

	bfr new_net_5117_bfr_before (
		.din(new_net_5117),
		.dout(new_net_718)
	);

	bfr new_net_5118_bfr_before (
		.din(new_net_5118),
		.dout(new_net_5117)
	);

	bfr new_net_5119_bfr_before (
		.din(new_net_5119),
		.dout(new_net_5118)
	);

	bfr new_net_5120_bfr_before (
		.din(new_net_5120),
		.dout(new_net_5119)
	);

	spl2 _0279__v_fanout (
		.a(_0279_),
		.b(new_net_717),
		.c(new_net_5120)
	);

	bfr new_net_5121_bfr_before (
		.din(new_net_5121),
		.dout(new_net_241)
	);

	bfr new_net_5122_bfr_before (
		.din(new_net_5122),
		.dout(new_net_5121)
	);

	bfr new_net_5123_bfr_before (
		.din(new_net_5123),
		.dout(new_net_5122)
	);

	bfr new_net_5124_bfr_before (
		.din(new_net_5124),
		.dout(new_net_5123)
	);

	spl2 _0482__v_fanout (
		.a(_0482_),
		.b(new_net_240),
		.c(new_net_5124)
	);

	bfr new_net_5125_bfr_before (
		.din(new_net_5125),
		.dout(new_net_2367)
	);

	bfr new_net_5126_bfr_before (
		.din(new_net_5126),
		.dout(new_net_5125)
	);

	bfr new_net_5127_bfr_before (
		.din(new_net_5127),
		.dout(new_net_5126)
	);

	bfr new_net_5128_bfr_before (
		.din(new_net_5128),
		.dout(new_net_5127)
	);

	spl2 _0160__v_fanout (
		.a(_0160_),
		.b(new_net_2366),
		.c(new_net_5128)
	);

	bfr new_net_5129_bfr_before (
		.din(new_net_5129),
		.dout(new_net_137)
	);

	bfr new_net_5130_bfr_before (
		.din(new_net_5130),
		.dout(new_net_5129)
	);

	bfr new_net_5131_bfr_before (
		.din(new_net_5131),
		.dout(new_net_5130)
	);

	bfr new_net_5132_bfr_before (
		.din(new_net_5132),
		.dout(new_net_5131)
	);

	spl2 _1536__v_fanout (
		.a(_1536_),
		.b(new_net_136),
		.c(new_net_5132)
	);

	bfr new_net_5133_bfr_before (
		.din(new_net_5133),
		.dout(new_net_3231)
	);

	bfr new_net_5134_bfr_before (
		.din(new_net_5134),
		.dout(new_net_5133)
	);

	bfr new_net_5135_bfr_before (
		.din(new_net_5135),
		.dout(new_net_5134)
	);

	bfr new_net_5136_bfr_before (
		.din(new_net_5136),
		.dout(new_net_5135)
	);

	spl2 _1273__v_fanout (
		.a(_1273_),
		.b(new_net_3230),
		.c(new_net_5136)
	);

	bfr new_net_5137_bfr_after (
		.din(_0787_),
		.dout(new_net_5137)
	);

	bfr new_net_5138_bfr_after (
		.din(new_net_5137),
		.dout(new_net_5138)
	);

	bfr new_net_5139_bfr_after (
		.din(new_net_5138),
		.dout(new_net_5139)
	);

	bfr new_net_5140_bfr_after (
		.din(new_net_5139),
		.dout(new_net_5140)
	);

	spl2 _0787__v_fanout (
		.a(new_net_5140),
		.b(new_net_840),
		.c(new_net_841)
	);

	spl2 _0840__v_fanout (
		.a(_0840_),
		.b(new_net_2671),
		.c(new_net_2672)
	);

	bfr new_net_5141_bfr_before (
		.din(new_net_5141),
		.dout(new_net_1031)
	);

	bfr new_net_5142_bfr_before (
		.din(new_net_5142),
		.dout(new_net_5141)
	);

	bfr new_net_5143_bfr_before (
		.din(new_net_5143),
		.dout(new_net_5142)
	);

	bfr new_net_5144_bfr_before (
		.din(new_net_5144),
		.dout(new_net_5143)
	);

	spl2 _0045__v_fanout (
		.a(_0045_),
		.b(new_net_1030),
		.c(new_net_5144)
	);

	bfr new_net_5145_bfr_before (
		.din(new_net_5145),
		.dout(new_net_2696)
	);

	bfr new_net_5146_bfr_before (
		.din(new_net_5146),
		.dout(new_net_5145)
	);

	bfr new_net_5147_bfr_before (
		.din(new_net_5147),
		.dout(new_net_5146)
	);

	bfr new_net_5148_bfr_before (
		.din(new_net_5148),
		.dout(new_net_5147)
	);

	spl2 _1765__v_fanout (
		.a(_1765_),
		.b(new_net_2695),
		.c(new_net_5148)
	);

	bfr new_net_5149_bfr_before (
		.din(new_net_5149),
		.dout(new_net_57)
	);

	bfr new_net_5150_bfr_before (
		.din(new_net_5150),
		.dout(new_net_5149)
	);

	bfr new_net_5151_bfr_before (
		.din(new_net_5151),
		.dout(new_net_5150)
	);

	bfr new_net_5152_bfr_before (
		.din(new_net_5152),
		.dout(new_net_5151)
	);

	spl2 _1435__v_fanout (
		.a(_1435_),
		.b(new_net_56),
		.c(new_net_5152)
	);

	bfr new_net_5153_bfr_before (
		.din(new_net_5153),
		.dout(new_net_1282)
	);

	bfr new_net_5154_bfr_before (
		.din(new_net_5154),
		.dout(new_net_5153)
	);

	bfr new_net_5155_bfr_before (
		.din(new_net_5155),
		.dout(new_net_5154)
	);

	bfr new_net_5156_bfr_before (
		.din(new_net_5156),
		.dout(new_net_5155)
	);

	spl2 _1350__v_fanout (
		.a(_1350_),
		.b(new_net_1281),
		.c(new_net_5156)
	);

	bfr new_net_5157_bfr_before (
		.din(new_net_5157),
		.dout(new_net_3000)
	);

	bfr new_net_5158_bfr_before (
		.din(new_net_5158),
		.dout(new_net_5157)
	);

	bfr new_net_5159_bfr_before (
		.din(new_net_5159),
		.dout(new_net_5158)
	);

	bfr new_net_5160_bfr_before (
		.din(new_net_5160),
		.dout(new_net_5159)
	);

	spl2 _1646__v_fanout (
		.a(_1646_),
		.b(new_net_2999),
		.c(new_net_5160)
	);

	bfr new_net_5161_bfr_before (
		.din(new_net_5161),
		.dout(new_net_1943)
	);

	bfr new_net_5162_bfr_before (
		.din(new_net_5162),
		.dout(new_net_5161)
	);

	bfr new_net_5163_bfr_before (
		.din(new_net_5163),
		.dout(new_net_5162)
	);

	bfr new_net_5164_bfr_before (
		.din(new_net_5164),
		.dout(new_net_5163)
	);

	spl2 _0570__v_fanout (
		.a(_0570_),
		.b(new_net_1942),
		.c(new_net_5164)
	);

	spl2 _1281__v_fanout (
		.a(_1281_),
		.b(new_net_614),
		.c(new_net_615)
	);

	spl2 _0384__v_fanout (
		.a(_0384_),
		.b(new_net_1265),
		.c(new_net_1266)
	);

	spl2 _1814__v_fanout (
		.a(_1814_),
		.b(new_net_1332),
		.c(new_net_1333)
	);

	spl2 _0784__v_fanout (
		.a(_0784_),
		.b(new_net_554),
		.c(new_net_555)
	);

	spl2 _0043__v_fanout (
		.a(_0043_),
		.b(new_net_673),
		.c(new_net_674)
	);

	spl2 _0628__v_fanout (
		.a(_0628_),
		.b(new_net_1168),
		.c(new_net_1169)
	);

	bfr new_net_5165_bfr_before (
		.din(new_net_5165),
		.dout(new_net_1209)
	);

	bfr new_net_5166_bfr_before (
		.din(new_net_5166),
		.dout(new_net_5165)
	);

	bfr new_net_5167_bfr_before (
		.din(new_net_5167),
		.dout(new_net_5166)
	);

	bfr new_net_5168_bfr_before (
		.din(new_net_5168),
		.dout(new_net_5167)
	);

	spl2 _0719__v_fanout (
		.a(_0719_),
		.b(new_net_1208),
		.c(new_net_5168)
	);

	spl2 _0096__v_fanout (
		.a(_0096_),
		.b(new_net_912),
		.c(new_net_913)
	);

	spl2 _0224__v_fanout (
		.a(_0224_),
		.b(new_net_1283),
		.c(new_net_1284)
	);

	spl2 _1764__v_fanout (
		.a(_1764_),
		.b(new_net_635),
		.c(new_net_636)
	);

	spl2 _0159__v_fanout (
		.a(_0159_),
		.b(new_net_2515),
		.c(new_net_2516)
	);

	spl2 _1349__v_fanout (
		.a(_1349_),
		.b(new_net_1214),
		.c(new_net_1215)
	);

	spl2 _1570__v_fanout (
		.a(_1570_),
		.b(new_net_1188),
		.c(new_net_1189)
	);

	spl2 _1272__v_fanout (
		.a(_1272_),
		.b(new_net_3175),
		.c(new_net_3176)
	);

	spl2 _1534__v_fanout (
		.a(_1534_),
		.b(new_net_2531),
		.c(new_net_2532)
	);

	spl2 _0569__v_fanout (
		.a(_0569_),
		.b(new_net_645),
		.c(new_net_646)
	);

	spl2 _1366__v_fanout (
		.a(_1366_),
		.b(new_net_799),
		.c(new_net_800)
	);

	spl2 _1690__v_fanout (
		.a(_1690_),
		.b(new_net_812),
		.c(new_net_813)
	);

	spl2 _0278__v_fanout (
		.a(_0278_),
		.b(new_net_512),
		.c(new_net_513)
	);

	spl2 _1204__v_fanout (
		.a(_1204_),
		.b(new_net_3211),
		.c(new_net_3212)
	);

	spl2 _1460__v_fanout (
		.a(_1460_),
		.b(new_net_703),
		.c(new_net_704)
	);

	spl2 _0444__v_fanout (
		.a(_0444_),
		.b(new_net_1846),
		.c(new_net_1847)
	);

	spl2 _0480__v_fanout (
		.a(_0480_),
		.b(new_net_164),
		.c(new_net_165)
	);

	spl2 _1434__v_fanout (
		.a(_1434_),
		.b(new_net_3125),
		.c(new_net_3126)
	);

	spl2 _0338__v_fanout (
		.a(_0338_),
		.b(new_net_1108),
		.c(new_net_1109)
	);

	spl2 _0541__v_fanout (
		.a(_0541_),
		.b(new_net_1850),
		.c(new_net_1851)
	);

	spl2 _1645__v_fanout (
		.a(_1645_),
		.b(new_net_54),
		.c(new_net_55)
	);

	spl2 _1642__v_fanout (
		.a(_1642_),
		.b(new_net_2811),
		.c(new_net_2812)
	);

	spl2 _0783__v_fanout (
		.a(_0783_),
		.b(new_net_52),
		.c(new_net_53)
	);

	spl2 _0041__v_fanout (
		.a(_0041_),
		.b(new_net_1022),
		.c(new_net_1023)
	);

	spl2 _1532__v_fanout (
		.a(_1532_),
		.b(new_net_2144),
		.c(new_net_2145)
	);

	spl2 _1270__v_fanout (
		.a(_1270_),
		.b(new_net_3111),
		.c(new_net_3112)
	);

	spl2 _1761__v_fanout (
		.a(_1761_),
		.b(new_net_2545),
		.c(new_net_2546)
	);

	spl2 _0381__v_fanout (
		.a(_0381_),
		.b(new_net_1144),
		.c(new_net_1145)
	);

	spl2 _0478__v_fanout (
		.a(_0478_),
		.b(new_net_2024),
		.c(new_net_2025)
	);

	spl2 _0566__v_fanout (
		.a(_0566_),
		.b(new_net_82),
		.c(new_net_83)
	);

	spl2 _0708__v_fanout (
		.a(_0708_),
		.b(new_net_647),
		.c(new_net_648)
	);

	spl2 _0157__v_fanout (
		.a(_0157_),
		.b(new_net_2234),
		.c(new_net_2235)
	);

	spl2 _1193__v_fanout (
		.a(_1193_),
		.b(new_net_1036),
		.c(new_net_1037)
	);

	spl2 _1432__v_fanout (
		.a(_1432_),
		.b(new_net_2809),
		.c(new_net_2810)
	);

	bfr new_net_5169_bfr_after (
		.din(_0648_),
		.dout(new_net_5169)
	);

	bfr new_net_5170_bfr_after (
		.din(new_net_5169),
		.dout(new_net_5170)
	);

	spl2 _0648__v_fanout (
		.a(new_net_5170),
		.b(new_net_166),
		.c(new_net_167)
	);

	spl2 _1347__v_fanout (
		.a(_1347_),
		.b(new_net_2655),
		.c(new_net_2656)
	);

	spl2 _0276__v_fanout (
		.a(_0276_),
		.b(new_net_132),
		.c(new_net_133)
	);

	spl2 _0040__v_fanout (
		.a(_0040_),
		.b(new_net_108),
		.c(new_net_109)
	);

	spl2 _0380__v_fanout (
		.a(_0380_),
		.b(new_net_1104),
		.c(new_net_1105)
	);

	bfr new_net_5171_bfr_before (
		.din(new_net_5171),
		.dout(new_net_417)
	);

	bfr new_net_5172_bfr_before (
		.din(new_net_5172),
		.dout(new_net_5171)
	);

	bfr new_net_5173_bfr_before (
		.din(new_net_5173),
		.dout(new_net_5172)
	);

	bfr new_net_5174_bfr_before (
		.din(new_net_5174),
		.dout(new_net_5173)
	);

	spl2 _0781__v_fanout (
		.a(_0781_),
		.b(new_net_416),
		.c(new_net_5174)
	);

	spl2 _0477__v_fanout (
		.a(_0477_),
		.b(new_net_74),
		.c(new_net_75)
	);

	spl2 _1269__v_fanout (
		.a(_1269_),
		.b(new_net_864),
		.c(new_net_865)
	);

	spl2 _0156__v_fanout (
		.a(_0156_),
		.b(new_net_2188),
		.c(new_net_2189)
	);

	spl2 _0646__v_fanout (
		.a(_0646_),
		.b(new_net_3005),
		.c(new_net_3006)
	);

	spl2 _0565__v_fanout (
		.a(_0565_),
		.b(new_net_3157),
		.c(new_net_3158)
	);

	spl2 _1346__v_fanout (
		.a(_1346_),
		.b(new_net_2446),
		.c(new_net_2447)
	);

	spl2 _1431__v_fanout (
		.a(_1431_),
		.b(new_net_2783),
		.c(new_net_2784)
	);

	spl2 _1760__v_fanout (
		.a(_1760_),
		.b(new_net_3131),
		.c(new_net_3132)
	);

	spl2 _1531__v_fanout (
		.a(_1531_),
		.b(new_net_1760),
		.c(new_net_1761)
	);

	spl2 _1192__v_fanout (
		.a(_1192_),
		.b(new_net_98),
		.c(new_net_99)
	);

	spl2 _1641__v_fanout (
		.a(_1641_),
		.b(new_net_2474),
		.c(new_net_2475)
	);

	spl2 _0275__v_fanout (
		.a(_0275_),
		.b(new_net_3215),
		.c(new_net_3216)
	);

	bfr new_net_5175_bfr_before (
		.din(new_net_5175),
		.dout(new_net_1365)
	);

	bfr new_net_5176_bfr_before (
		.din(new_net_5176),
		.dout(new_net_5175)
	);

	bfr new_net_5177_bfr_before (
		.din(new_net_5177),
		.dout(new_net_5176)
	);

	bfr new_net_5178_bfr_before (
		.din(new_net_5178),
		.dout(new_net_5177)
	);

	spl2 _0153__v_fanout (
		.a(_0153_),
		.b(new_net_1364),
		.c(new_net_5178)
	);

	bfr new_net_5179_bfr_before (
		.din(new_net_5179),
		.dout(new_net_493)
	);

	bfr new_net_5180_bfr_before (
		.din(new_net_5180),
		.dout(new_net_5179)
	);

	bfr new_net_5181_bfr_before (
		.din(new_net_5181),
		.dout(new_net_5180)
	);

	bfr new_net_5182_bfr_before (
		.din(new_net_5182),
		.dout(new_net_5181)
	);

	spl2 _1190__v_fanout (
		.a(_1190_),
		.b(new_net_492),
		.c(new_net_5182)
	);

	bfr new_net_5183_bfr_before (
		.din(new_net_5183),
		.dout(new_net_2729)
	);

	bfr new_net_5184_bfr_before (
		.din(new_net_5184),
		.dout(new_net_5183)
	);

	bfr new_net_5185_bfr_before (
		.din(new_net_5185),
		.dout(new_net_5184)
	);

	bfr new_net_5186_bfr_before (
		.din(new_net_5186),
		.dout(new_net_5185)
	);

	spl2 _1639__v_fanout (
		.a(_1639_),
		.b(new_net_2728),
		.c(new_net_5186)
	);

	bfr new_net_5187_bfr_before (
		.din(new_net_5187),
		.dout(new_net_2031)
	);

	bfr new_net_5188_bfr_before (
		.din(new_net_5188),
		.dout(new_net_5187)
	);

	bfr new_net_5189_bfr_before (
		.din(new_net_5189),
		.dout(new_net_5188)
	);

	bfr new_net_5190_bfr_before (
		.din(new_net_5190),
		.dout(new_net_5189)
	);

	spl2 _1344__v_fanout (
		.a(_1344_),
		.b(new_net_2030),
		.c(new_net_5190)
	);

	spl2 _0645__v_fanout (
		.a(_0645_),
		.b(new_net_2787),
		.c(new_net_2788)
	);

	bfr new_net_5191_bfr_before (
		.din(new_net_5191),
		.dout(new_net_2948)
	);

	bfr new_net_5192_bfr_before (
		.din(new_net_5192),
		.dout(new_net_5191)
	);

	bfr new_net_5193_bfr_before (
		.din(new_net_5193),
		.dout(new_net_5192)
	);

	bfr new_net_5194_bfr_before (
		.din(new_net_5194),
		.dout(new_net_5193)
	);

	spl2 _0038__v_fanout (
		.a(_0038_),
		.b(new_net_2947),
		.c(new_net_5194)
	);

	bfr new_net_5195_bfr_before (
		.din(new_net_5195),
		.dout(new_net_1309)
	);

	bfr new_net_5196_bfr_before (
		.din(new_net_5196),
		.dout(new_net_5195)
	);

	bfr new_net_5197_bfr_before (
		.din(new_net_5197),
		.dout(new_net_5196)
	);

	bfr new_net_5198_bfr_before (
		.din(new_net_5198),
		.dout(new_net_5197)
	);

	spl2 _0475__v_fanout (
		.a(_0475_),
		.b(new_net_1308),
		.c(new_net_5198)
	);

	bfr new_net_5199_bfr_after (
		.din(_0718_),
		.dout(new_net_5199)
	);

	bfr new_net_5200_bfr_after (
		.din(new_net_5199),
		.dout(new_net_5200)
	);

	bfr new_net_5201_bfr_after (
		.din(new_net_5200),
		.dout(new_net_5201)
	);

	bfr new_net_5202_bfr_after (
		.din(new_net_5201),
		.dout(new_net_5202)
	);

	spl2 _0718__v_fanout (
		.a(new_net_5202),
		.b(new_net_2517),
		.c(new_net_2518)
	);

	bfr new_net_5203_bfr_before (
		.din(new_net_5203),
		.dout(new_net_1701)
	);

	bfr new_net_5204_bfr_before (
		.din(new_net_5204),
		.dout(new_net_5203)
	);

	bfr new_net_5205_bfr_before (
		.din(new_net_5205),
		.dout(new_net_5204)
	);

	bfr new_net_5206_bfr_before (
		.din(new_net_5206),
		.dout(new_net_5205)
	);

	spl2 _1529__v_fanout (
		.a(_1529_),
		.b(new_net_1700),
		.c(new_net_5206)
	);

	spl2 _0780__v_fanout (
		.a(_0780_),
		.b(new_net_370),
		.c(new_net_371)
	);

	bfr new_net_5207_bfr_before (
		.din(new_net_5207),
		.dout(new_net_2733)
	);

	bfr new_net_5208_bfr_before (
		.din(new_net_5208),
		.dout(new_net_5207)
	);

	bfr new_net_5209_bfr_before (
		.din(new_net_5209),
		.dout(new_net_5208)
	);

	bfr new_net_5210_bfr_before (
		.din(new_net_5210),
		.dout(new_net_5209)
	);

	spl2 _0563__v_fanout (
		.a(_0563_),
		.b(new_net_2732),
		.c(new_net_5210)
	);

	bfr new_net_5211_bfr_before (
		.din(new_net_5211),
		.dout(new_net_2578)
	);

	bfr new_net_5212_bfr_before (
		.din(new_net_5212),
		.dout(new_net_5211)
	);

	bfr new_net_5213_bfr_before (
		.din(new_net_5213),
		.dout(new_net_5212)
	);

	bfr new_net_5214_bfr_before (
		.din(new_net_5214),
		.dout(new_net_5213)
	);

	spl2 _0272__v_fanout (
		.a(_0272_),
		.b(new_net_2577),
		.c(new_net_5214)
	);

	bfr new_net_5215_bfr_before (
		.din(new_net_5215),
		.dout(new_net_2692)
	);

	bfr new_net_5216_bfr_before (
		.din(new_net_5216),
		.dout(new_net_5215)
	);

	bfr new_net_5217_bfr_before (
		.din(new_net_5217),
		.dout(new_net_5216)
	);

	bfr new_net_5218_bfr_before (
		.din(new_net_5218),
		.dout(new_net_5217)
	);

	spl2 _1758__v_fanout (
		.a(_1758_),
		.b(new_net_2691),
		.c(new_net_5218)
	);

	bfr new_net_5219_bfr_before (
		.din(new_net_5219),
		.dout(new_net_2966)
	);

	bfr new_net_5220_bfr_before (
		.din(new_net_5220),
		.dout(new_net_5219)
	);

	bfr new_net_5221_bfr_before (
		.din(new_net_5221),
		.dout(new_net_5220)
	);

	bfr new_net_5222_bfr_before (
		.din(new_net_5222),
		.dout(new_net_5221)
	);

	spl2 _1267__v_fanout (
		.a(_1267_),
		.b(new_net_2965),
		.c(new_net_5222)
	);

	bfr new_net_5223_bfr_before (
		.din(new_net_5223),
		.dout(new_net_1240)
	);

	bfr new_net_5224_bfr_before (
		.din(new_net_5224),
		.dout(new_net_5223)
	);

	bfr new_net_5225_bfr_before (
		.din(new_net_5225),
		.dout(new_net_5224)
	);

	bfr new_net_5226_bfr_before (
		.din(new_net_5226),
		.dout(new_net_5225)
	);

	spl2 _0378__v_fanout (
		.a(_0378_),
		.b(new_net_1239),
		.c(new_net_5226)
	);

	bfr new_net_5227_bfr_before (
		.din(new_net_5227),
		.dout(new_net_2085)
	);

	bfr new_net_5228_bfr_before (
		.din(new_net_5228),
		.dout(new_net_5227)
	);

	bfr new_net_5229_bfr_before (
		.din(new_net_5229),
		.dout(new_net_5228)
	);

	bfr new_net_5230_bfr_before (
		.din(new_net_5230),
		.dout(new_net_5229)
	);

	spl2 _1429__v_fanout (
		.a(_1429_),
		.b(new_net_2084),
		.c(new_net_5230)
	);

	spl2 _0716__v_fanout (
		.a(_0716_),
		.b(new_net_2128),
		.c(new_net_2129)
	);

	spl2 _0271__v_fanout (
		.a(_0271_),
		.b(new_net_2378),
		.c(new_net_2379)
	);

	spl2 _1266__v_fanout (
		.a(_1266_),
		.b(new_net_248),
		.c(new_net_249)
	);

	bfr new_net_5231_bfr_before (
		.din(new_net_5231),
		.dout(new_net_644)
	);

	bfr new_net_5232_bfr_before (
		.din(new_net_5232),
		.dout(new_net_5231)
	);

	bfr new_net_5233_bfr_before (
		.din(new_net_5233),
		.dout(new_net_5232)
	);

	bfr new_net_5234_bfr_before (
		.din(new_net_5234),
		.dout(new_net_5233)
	);

	spl2 _0642__v_fanout (
		.a(_0642_),
		.b(new_net_643),
		.c(new_net_5234)
	);

	spl2 _1189__v_fanout (
		.a(_1189_),
		.b(new_net_86),
		.c(new_net_87)
	);

	spl2 _1757__v_fanout (
		.a(_1757_),
		.b(new_net_2388),
		.c(new_net_2389)
	);

	spl2 _1528__v_fanout (
		.a(_1528_),
		.b(new_net_1388),
		.c(new_net_1389)
	);

	spl2 _1368__v_fanout (
		.a(_1368_),
		.b(new_net_1946),
		.c(new_net_1947)
	);

	spl2 _1462__v_fanout (
		.a(_1462_),
		.b(new_net_826),
		.c(new_net_827)
	);

	spl2 _1428__v_fanout (
		.a(_1428_),
		.b(new_net_2677),
		.c(new_net_2678)
	);

	spl2 _0341__v_fanout (
		.a(_0341_),
		.b(new_net_1220),
		.c(new_net_1221)
	);

	spl2 _0474__v_fanout (
		.a(_0474_),
		.b(new_net_1100),
		.c(new_net_1101)
	);

	spl2 _0098__v_fanout (
		.a(_0098_),
		.b(new_net_325),
		.c(new_net_326)
	);

	spl2 _0377__v_fanout (
		.a(_0377_),
		.b(new_net_1018),
		.c(new_net_1019)
	);

	spl2 _1816__v_fanout (
		.a(_1816_),
		.b(new_net_1429),
		.c(new_net_1430)
	);

	spl2 _1343__v_fanout (
		.a(_1343_),
		.b(new_net_1856),
		.c(new_net_1857)
	);

	spl2 _0152__v_fanout (
		.a(_0152_),
		.b(new_net_2012),
		.c(new_net_2013)
	);

	spl2 _1692__v_fanout (
		.a(_1692_),
		.b(new_net_1533),
		.c(new_net_1534)
	);

	spl2 _1572__v_fanout (
		.a(_1572_),
		.b(new_net_1722),
		.c(new_net_1723)
	);

	spl2 _1129__v_fanout (
		.a(_1129_),
		.b(new_net_2973),
		.c(new_net_2974)
	);

	spl2 _0543__v_fanout (
		.a(_0543_),
		.b(new_net_2565),
		.c(new_net_2566)
	);

	spl2 _0037__v_fanout (
		.a(_0037_),
		.b(new_net_2738),
		.c(new_net_2739)
	);

	spl2 _0446__v_fanout (
		.a(_0446_),
		.b(new_net_2244),
		.c(new_net_2245)
	);

	spl2 _1638__v_fanout (
		.a(_1638_),
		.b(new_net_2675),
		.c(new_net_2676)
	);

	spl2 _1206__v_fanout (
		.a(_1206_),
		.b(new_net_299),
		.c(new_net_300)
	);

	spl2 _1283__v_fanout (
		.a(_1283_),
		.b(new_net_988),
		.c(new_net_989)
	);

	spl2 _0226__v_fanout (
		.a(_0226_),
		.b(new_net_94),
		.c(new_net_95)
	);

	spl2 _1341__v_fanout (
		.a(_1341_),
		.b(new_net_1517),
		.c(new_net_1518)
	);

	spl2 _0269__v_fanout (
		.a(_0269_),
		.b(new_net_1962),
		.c(new_net_1963)
	);

	spl2 _1187__v_fanout (
		.a(_1187_),
		.b(new_net_2931),
		.c(new_net_2932)
	);

	spl2 _0035__v_fanout (
		.a(_0035_),
		.b(new_net_2329),
		.c(new_net_2330)
	);

	spl2 _0630__v_fanout (
		.a(_0630_),
		.b(new_net_1044),
		.c(new_net_1045)
	);

	spl2 _1426__v_fanout (
		.a(_1426_),
		.b(new_net_2597),
		.c(new_net_2598)
	);

	spl2 _1526__v_fanout (
		.a(_1526_),
		.b(new_net_1032),
		.c(new_net_1033)
	);

	spl2 _0472__v_fanout (
		.a(_0472_),
		.b(new_net_810),
		.c(new_net_811)
	);

	spl2 _0375__v_fanout (
		.a(_0375_),
		.b(new_net_729),
		.c(new_net_730)
	);

	spl2 _1755__v_fanout (
		.a(_1755_),
		.b(new_net_2098),
		.c(new_net_2099)
	);

	bfr new_net_5235_bfr_after (
		.din(_0562_),
		.dout(new_net_5235)
	);

	bfr new_net_5236_bfr_after (
		.din(new_net_5235),
		.dout(new_net_5236)
	);

	spl2 _0562__v_fanout (
		.a(new_net_5236),
		.b(new_net_1682),
		.c(new_net_1683)
	);

	spl2 _1128__v_fanout (
		.a(_1128_),
		.b(new_net_876),
		.c(new_net_877)
	);

	spl2 _1636__v_fanout (
		.a(_1636_),
		.b(new_net_2595),
		.c(new_net_2596)
	);

	spl2 _1264__v_fanout (
		.a(_1264_),
		.b(new_net_3153),
		.c(new_net_3154)
	);

	spl2 _0150__v_fanout (
		.a(_0150_),
		.b(new_net_1940),
		.c(new_net_1941)
	);

	spl2 _0715__v_fanout (
		.a(_0715_),
		.b(new_net_1084),
		.c(new_net_1085)
	);

	spl2 _1635__v_fanout (
		.a(_1635_),
		.b(new_net_2533),
		.c(new_net_2534)
	);

	spl2 _0268__v_fanout (
		.a(_0268_),
		.b(new_net_1690),
		.c(new_net_1691)
	);

	spl2 _1186__v_fanout (
		.a(_1186_),
		.b(new_net_2736),
		.c(new_net_2737)
	);

	spl2 _0560__v_fanout (
		.a(_0560_),
		.b(new_net_1614),
		.c(new_net_1615)
	);

	spl2 _1525__v_fanout (
		.a(_1525_),
		.b(new_net_1630),
		.c(new_net_1631)
	);

	spl2 _1340__v_fanout (
		.a(_1340_),
		.b(new_net_1306),
		.c(new_net_1307)
	);

	spl2 _0149__v_fanout (
		.a(_0149_),
		.b(new_net_1916),
		.c(new_net_1917)
	);

	spl2 _1425__v_fanout (
		.a(_1425_),
		.b(new_net_2543),
		.c(new_net_2544)
	);

	spl2 _0374__v_fanout (
		.a(_0374_),
		.b(new_net_520),
		.c(new_net_521)
	);

	spl2 _1754__v_fanout (
		.a(_1754_),
		.b(new_net_1896),
		.c(new_net_1897)
	);

	spl2 _1127__v_fanout (
		.a(_1127_),
		.b(new_net_856),
		.c(new_net_857)
	);

	spl2 _0034__v_fanout (
		.a(_0034_),
		.b(new_net_818),
		.c(new_net_819)
	);

	spl2 _1263__v_fanout (
		.a(_1263_),
		.b(new_net_2777),
		.c(new_net_2778)
	);

	bfr new_net_5237_bfr_before (
		.din(new_net_5237),
		.dout(new_net_1015)
	);

	bfr new_net_5238_bfr_before (
		.din(new_net_5238),
		.dout(new_net_5237)
	);

	bfr new_net_5239_bfr_before (
		.din(new_net_5239),
		.dout(new_net_5238)
	);

	bfr new_net_5240_bfr_before (
		.din(new_net_5240),
		.dout(new_net_5239)
	);

	spl2 _0713__v_fanout (
		.a(_0713_),
		.b(new_net_1014),
		.c(new_net_5240)
	);

	spl2 _0471__v_fanout (
		.a(_0471_),
		.b(new_net_586),
		.c(new_net_587)
	);

	bfr new_net_5241_bfr_before (
		.din(new_net_5241),
		.dout(new_net_17)
	);

	bfr new_net_5242_bfr_before (
		.din(new_net_5242),
		.dout(new_net_5241)
	);

	bfr new_net_5243_bfr_before (
		.din(new_net_5243),
		.dout(new_net_5242)
	);

	bfr new_net_5244_bfr_before (
		.din(new_net_5244),
		.dout(new_net_5243)
	);

	spl2 _0468__v_fanout (
		.a(_0468_),
		.b(new_net_16),
		.c(new_net_5244)
	);

	bfr new_net_5245_bfr_before (
		.din(new_net_5245),
		.dout(new_net_871)
	);

	bfr new_net_5246_bfr_before (
		.din(new_net_5246),
		.dout(new_net_5245)
	);

	bfr new_net_5247_bfr_before (
		.din(new_net_5247),
		.dout(new_net_5246)
	);

	bfr new_net_5248_bfr_before (
		.din(new_net_5248),
		.dout(new_net_5247)
	);

	spl2 _1338__v_fanout (
		.a(_1338_),
		.b(new_net_870),
		.c(new_net_5248)
	);

	spl2 _0559__v_fanout (
		.a(_0559_),
		.b(new_net_2036),
		.c(new_net_2037)
	);

	bfr new_net_5249_bfr_before (
		.din(new_net_5249),
		.dout(new_net_1605)
	);

	bfr new_net_5250_bfr_before (
		.din(new_net_5250),
		.dout(new_net_5249)
	);

	bfr new_net_5251_bfr_before (
		.din(new_net_5251),
		.dout(new_net_5250)
	);

	bfr new_net_5252_bfr_before (
		.din(new_net_5252),
		.dout(new_net_5251)
	);

	spl2 _0031__v_fanout (
		.a(_0031_),
		.b(new_net_1604),
		.c(new_net_5252)
	);

	bfr new_net_5253_bfr_before (
		.din(new_net_5253),
		.dout(new_net_2316)
	);

	bfr new_net_5254_bfr_before (
		.din(new_net_5254),
		.dout(new_net_5253)
	);

	bfr new_net_5255_bfr_before (
		.din(new_net_5255),
		.dout(new_net_5254)
	);

	bfr new_net_5256_bfr_before (
		.din(new_net_5256),
		.dout(new_net_5255)
	);

	spl2 _1184__v_fanout (
		.a(_1184_),
		.b(new_net_2315),
		.c(new_net_5256)
	);

	bfr new_net_5257_bfr_before (
		.din(new_net_5257),
		.dout(new_net_2465)
	);

	bfr new_net_5258_bfr_before (
		.din(new_net_5258),
		.dout(new_net_5257)
	);

	bfr new_net_5259_bfr_before (
		.din(new_net_5259),
		.dout(new_net_5258)
	);

	bfr new_net_5260_bfr_before (
		.din(new_net_5260),
		.dout(new_net_5259)
	);

	spl2 _1423__v_fanout (
		.a(_1423_),
		.b(new_net_2464),
		.c(new_net_5260)
	);

	bfr new_net_5261_bfr_before (
		.din(new_net_5261),
		.dout(new_net_1041)
	);

	bfr new_net_5262_bfr_before (
		.din(new_net_5262),
		.dout(new_net_5261)
	);

	bfr new_net_5263_bfr_before (
		.din(new_net_5263),
		.dout(new_net_5262)
	);

	bfr new_net_5264_bfr_before (
		.din(new_net_5264),
		.dout(new_net_5263)
	);

	spl2 _1522__v_fanout (
		.a(_1522_),
		.b(new_net_1040),
		.c(new_net_5264)
	);

	bfr new_net_5265_bfr_before (
		.din(new_net_5265),
		.dout(new_net_1432)
	);

	bfr new_net_5266_bfr_before (
		.din(new_net_5266),
		.dout(new_net_5265)
	);

	bfr new_net_5267_bfr_before (
		.din(new_net_5267),
		.dout(new_net_5266)
	);

	bfr new_net_5268_bfr_before (
		.din(new_net_5268),
		.dout(new_net_5267)
	);

	spl2 _0266__v_fanout (
		.a(_0266_),
		.b(new_net_1431),
		.c(new_net_5268)
	);

	spl2 _0712__v_fanout (
		.a(_0712_),
		.b(new_net_994),
		.c(new_net_995)
	);

	bfr new_net_5269_bfr_before (
		.din(new_net_5269),
		.dout(new_net_1935)
	);

	bfr new_net_5270_bfr_before (
		.din(new_net_5270),
		.dout(new_net_5269)
	);

	bfr new_net_5271_bfr_before (
		.din(new_net_5271),
		.dout(new_net_5270)
	);

	bfr new_net_5272_bfr_before (
		.din(new_net_5272),
		.dout(new_net_5271)
	);

	spl2 _1124__v_fanout (
		.a(_1124_),
		.b(new_net_1934),
		.c(new_net_5272)
	);

	bfr new_net_5273_bfr_before (
		.din(new_net_5273),
		.dout(new_net_2467)
	);

	bfr new_net_5274_bfr_before (
		.din(new_net_5274),
		.dout(new_net_5273)
	);

	bfr new_net_5275_bfr_before (
		.din(new_net_5275),
		.dout(new_net_5274)
	);

	bfr new_net_5276_bfr_before (
		.din(new_net_5276),
		.dout(new_net_5275)
	);

	spl2 _1633__v_fanout (
		.a(_1633_),
		.b(new_net_2466),
		.c(new_net_5276)
	);

	bfr new_net_5277_bfr_before (
		.din(new_net_5277),
		.dout(new_net_2715)
	);

	bfr new_net_5278_bfr_before (
		.din(new_net_5278),
		.dout(new_net_5277)
	);

	bfr new_net_5279_bfr_before (
		.din(new_net_5279),
		.dout(new_net_5278)
	);

	bfr new_net_5280_bfr_before (
		.din(new_net_5280),
		.dout(new_net_5279)
	);

	spl2 _1261__v_fanout (
		.a(_1261_),
		.b(new_net_2714),
		.c(new_net_5280)
	);

	bfr new_net_5281_bfr_before (
		.din(new_net_5281),
		.dout(new_net_3265)
	);

	bfr new_net_5282_bfr_before (
		.din(new_net_5282),
		.dout(new_net_5281)
	);

	bfr new_net_5283_bfr_before (
		.din(new_net_5283),
		.dout(new_net_5282)
	);

	bfr new_net_5284_bfr_before (
		.din(new_net_5284),
		.dout(new_net_5283)
	);

	spl2 _0371__v_fanout (
		.a(_0371_),
		.b(new_net_3264),
		.c(new_net_5284)
	);

	bfr new_net_5285_bfr_after (
		.din(_0641_),
		.dout(new_net_5285)
	);

	bfr new_net_5286_bfr_after (
		.din(new_net_5285),
		.dout(new_net_5286)
	);

	bfr new_net_5287_bfr_after (
		.din(new_net_5286),
		.dout(new_net_5287)
	);

	bfr new_net_5288_bfr_after (
		.din(new_net_5287),
		.dout(new_net_5288)
	);

	spl2 _0641__v_fanout (
		.a(new_net_5288),
		.b(new_net_456),
		.c(new_net_457)
	);

	bfr new_net_5289_bfr_before (
		.din(new_net_5289),
		.dout(new_net_2165)
	);

	bfr new_net_5290_bfr_before (
		.din(new_net_5290),
		.dout(new_net_5289)
	);

	bfr new_net_5291_bfr_before (
		.din(new_net_5291),
		.dout(new_net_5290)
	);

	bfr new_net_5292_bfr_before (
		.din(new_net_5292),
		.dout(new_net_5291)
	);

	spl2 _1751__v_fanout (
		.a(_1751_),
		.b(new_net_2164),
		.c(new_net_5292)
	);

	bfr new_net_5293_bfr_before (
		.din(new_net_5293),
		.dout(new_net_1835)
	);

	bfr new_net_5294_bfr_before (
		.din(new_net_5294),
		.dout(new_net_5293)
	);

	bfr new_net_5295_bfr_before (
		.din(new_net_5295),
		.dout(new_net_5294)
	);

	bfr new_net_5296_bfr_before (
		.din(new_net_5296),
		.dout(new_net_5295)
	);

	spl2 _0147__v_fanout (
		.a(_0147_),
		.b(new_net_1834),
		.c(new_net_5296)
	);

	spl2 _0101__v_fanout (
		.a(_0101_),
		.b(new_net_1704),
		.c(new_net_1705)
	);

	spl2 _1574__v_fanout (
		.a(_1574_),
		.b(new_net_1928),
		.c(new_net_1929)
	);

	spl2 _1337__v_fanout (
		.a(_1337_),
		.b(new_net_801),
		.c(new_net_802)
	);

	spl2 _1422__v_fanout (
		.a(_1422_),
		.b(new_net_838),
		.c(new_net_839)
	);

	spl2 _0265__v_fanout (
		.a(_0265_),
		.b(new_net_2637),
		.c(new_net_2638)
	);

	bfr new_net_5297_bfr_before (
		.din(new_net_5297),
		.dout(new_net_1522)
	);

	bfr new_net_5298_bfr_before (
		.din(new_net_5298),
		.dout(new_net_5297)
	);

	bfr new_net_5299_bfr_before (
		.din(new_net_5299),
		.dout(new_net_5298)
	);

	bfr new_net_5300_bfr_before (
		.din(new_net_5300),
		.dout(new_net_5299)
	);

	spl2 _0556__v_fanout (
		.a(_0556_),
		.b(new_net_1521),
		.c(new_net_5300)
	);

	spl2 _0639__v_fanout (
		.a(_0639_),
		.b(new_net_80),
		.c(new_net_81)
	);

	spl2 _1208__v_fanout (
		.a(_1208_),
		.b(new_net_693),
		.c(new_net_694)
	);

	spl2 _1123__v_fanout (
		.a(_1123_),
		.b(new_net_1748),
		.c(new_net_1749)
	);

	spl2 _1521__v_fanout (
		.a(_1521_),
		.b(new_net_892),
		.c(new_net_893)
	);

	spl2 _1131__v_fanout (
		.a(_1131_),
		.b(new_net_966),
		.c(new_net_967)
	);

	spl2 _1071__v_fanout (
		.a(_1071_),
		.b(new_net_3270),
		.c(new_net_3271)
	);

	spl2 _0449__v_fanout (
		.a(_0449_),
		.b(new_net_598),
		.c(new_net_599)
	);

	spl2 _0228__v_fanout (
		.a(_0228_),
		.b(new_net_174),
		.c(new_net_175)
	);

	spl2 _0370__v_fanout (
		.a(_0370_),
		.b(new_net_2801),
		.c(new_net_2802)
	);

	spl2 _1370__v_fanout (
		.a(_1370_),
		.b(new_net_1515),
		.c(new_net_1516)
	);

	spl2 _1694__v_fanout (
		.a(_1694_),
		.b(new_net_1620),
		.c(new_net_1621)
	);

	spl2 _0030__v_fanout (
		.a(_0030_),
		.b(new_net_622),
		.c(new_net_623)
	);

	spl2 _1464__v_fanout (
		.a(_1464_),
		.b(new_net_566),
		.c(new_net_567)
	);

	spl2 _1183__v_fanout (
		.a(_1183_),
		.b(new_net_2126),
		.c(new_net_2127)
	);

	spl2 _1631__v_fanout (
		.a(_1631_),
		.b(new_net_610),
		.c(new_net_611)
	);

	spl2 _1750__v_fanout (
		.a(_1750_),
		.b(new_net_2120),
		.c(new_net_2121)
	);

	spl2 _0146__v_fanout (
		.a(_0146_),
		.b(new_net_1782),
		.c(new_net_1783)
	);

	spl2 _0343__v_fanout (
		.a(_0343_),
		.b(new_net_1746),
		.c(new_net_1747)
	);

	spl2 _1285__v_fanout (
		.a(_1285_),
		.b(new_net_420),
		.c(new_net_421)
	);

	spl2 _1260__v_fanout (
		.a(_1260_),
		.b(new_net_2288),
		.c(new_net_2289)
	);

	spl2 _1818__v_fanout (
		.a(_1818_),
		.b(new_net_1563),
		.c(new_net_1564)
	);

	spl2 _0144__v_fanout (
		.a(_0144_),
		.b(new_net_2929),
		.c(new_net_2930)
	);

	spl2 _0262__v_fanout (
		.a(_0262_),
		.b(new_net_1421),
		.c(new_net_1422)
	);

	spl2 _0638__v_fanout (
		.a(_0638_),
		.b(new_net_3155),
		.c(new_net_3156)
	);

	spl2 _1070__v_fanout (
		.a(_1070_),
		.b(new_net_1790),
		.c(new_net_1791)
	);

	spl2 _0368__v_fanout (
		.a(_0368_),
		.b(new_net_2583),
		.c(new_net_2584)
	);

	spl2 _0545__v_fanout (
		.a(_0545_),
		.b(new_net_2645),
		.c(new_net_2646)
	);

	spl2 _1748__v_fanout (
		.a(_1748_),
		.b(new_net_860),
		.c(new_net_861)
	);

	spl2 _1258__v_fanout (
		.a(_1258_),
		.b(new_net_1906),
		.c(new_net_1907)
	);

	spl2 _0028__v_fanout (
		.a(_0028_),
		.b(new_net_550),
		.c(new_net_551)
	);

	spl2 _1629__v_fanout (
		.a(_1629_),
		.b(new_net_2298),
		.c(new_net_2299)
	);

	spl2 _1181__v_fanout (
		.a(_1181_),
		.b(new_net_2851),
		.c(new_net_2852)
	);

	spl2 _1420__v_fanout (
		.a(_1420_),
		.b(new_net_2355),
		.c(new_net_2356)
	);

	spl2 _1519__v_fanout (
		.a(_1519_),
		.b(new_net_494),
		.c(new_net_495)
	);

	spl2 _1335__v_fanout (
		.a(_1335_),
		.b(new_net_765),
		.c(new_net_766)
	);

	spl2 _1121__v_fanout (
		.a(_1121_),
		.b(new_net_1390),
		.c(new_net_1391)
	);

	bfr new_net_5301_bfr_after (
		.din(_0467_),
		.dout(new_net_5301)
	);

	bfr new_net_5302_bfr_after (
		.din(new_net_5301),
		.dout(new_net_5302)
	);

	spl2 _0467__v_fanout (
		.a(new_net_5302),
		.b(new_net_3069),
		.c(new_net_3070)
	);

	spl2 _1257__v_fanout (
		.a(_1257_),
		.b(new_net_2541),
		.c(new_net_2542)
	);

	spl2 _1628__v_fanout (
		.a(_1628_),
		.b(new_net_2258),
		.c(new_net_2259)
	);

	spl2 _0465__v_fanout (
		.a(_0465_),
		.b(new_net_1146),
		.c(new_net_1147)
	);

	bfr new_net_5303_bfr_before (
		.din(new_net_5303),
		.dout(new_net_2731)
	);

	bfr new_net_5304_bfr_before (
		.din(new_net_5304),
		.dout(new_net_5303)
	);

	bfr new_net_5305_bfr_before (
		.din(new_net_5305),
		.dout(new_net_5304)
	);

	bfr new_net_5306_bfr_before (
		.din(new_net_5306),
		.dout(new_net_5305)
	);

	spl2 _0636__v_fanout (
		.a(_0636_),
		.b(new_net_2730),
		.c(new_net_5306)
	);

	spl2 _0142__v_fanout (
		.a(_0142_),
		.b(new_net_2511),
		.c(new_net_2512)
	);

	spl2 _1334__v_fanout (
		.a(_1334_),
		.b(new_net_697),
		.c(new_net_698)
	);

	spl2 _1120__v_fanout (
		.a(_1120_),
		.b(new_net_1192),
		.c(new_net_1193)
	);

	spl2 _1069__v_fanout (
		.a(_1069_),
		.b(new_net_1752),
		.c(new_net_1753)
	);

	spl2 _1180__v_fanout (
		.a(_1180_),
		.b(new_net_1598),
		.c(new_net_1599)
	);

	spl2 _0367__v_fanout (
		.a(_0367_),
		.b(new_net_653),
		.c(new_net_654)
	);

	spl2 _1419__v_fanout (
		.a(_1419_),
		.b(new_net_222),
		.c(new_net_223)
	);

	spl2 _0027__v_fanout (
		.a(_0027_),
		.b(new_net_884),
		.c(new_net_885)
	);

	spl2 _0261__v_fanout (
		.a(_0261_),
		.b(new_net_1824),
		.c(new_net_1825)
	);

	spl2 _1518__v_fanout (
		.a(_1518_),
		.b(new_net_1277),
		.c(new_net_1278)
	);

	spl2 _1747__v_fanout (
		.a(_1747_),
		.b(new_net_628),
		.c(new_net_629)
	);

	bfr new_net_5307_bfr_before (
		.din(new_net_5307),
		.dout(new_net_3208)
	);

	bfr new_net_5308_bfr_before (
		.din(new_net_5308),
		.dout(new_net_5307)
	);

	bfr new_net_5309_bfr_before (
		.din(new_net_5309),
		.dout(new_net_5308)
	);

	bfr new_net_5310_bfr_before (
		.din(new_net_5310),
		.dout(new_net_5309)
	);

	spl2 _1516__v_fanout (
		.a(_1516_),
		.b(new_net_3207),
		.c(new_net_5310)
	);

	bfr new_net_5311_bfr_before (
		.din(new_net_5311),
		.dout(new_net_2758)
	);

	bfr new_net_5312_bfr_before (
		.din(new_net_5312),
		.dout(new_net_5311)
	);

	bfr new_net_5313_bfr_before (
		.din(new_net_5313),
		.dout(new_net_5312)
	);

	bfr new_net_5314_bfr_before (
		.din(new_net_5314),
		.dout(new_net_5313)
	);

	spl2 _1178__v_fanout (
		.a(_1178_),
		.b(new_net_2757),
		.c(new_net_5314)
	);

	bfr new_net_5315_bfr_before (
		.din(new_net_5315),
		.dout(new_net_1971)
	);

	bfr new_net_5316_bfr_before (
		.din(new_net_5316),
		.dout(new_net_5315)
	);

	bfr new_net_5317_bfr_before (
		.din(new_net_5317),
		.dout(new_net_5316)
	);

	bfr new_net_5318_bfr_before (
		.din(new_net_5318),
		.dout(new_net_5317)
	);

	spl2 _0365__v_fanout (
		.a(_0365_),
		.b(new_net_1970),
		.c(new_net_5318)
	);

	bfr new_net_5319_bfr_before (
		.din(new_net_5319),
		.dout(new_net_3064)
	);

	bfr new_net_5320_bfr_before (
		.din(new_net_5320),
		.dout(new_net_5319)
	);

	bfr new_net_5321_bfr_before (
		.din(new_net_5321),
		.dout(new_net_5320)
	);

	bfr new_net_5322_bfr_before (
		.din(new_net_5322),
		.dout(new_net_5321)
	);

	spl2 _1332__v_fanout (
		.a(_1332_),
		.b(new_net_3063),
		.c(new_net_5322)
	);

	bfr new_net_5323_bfr_before (
		.din(new_net_5323),
		.dout(new_net_1915)
	);

	bfr new_net_5324_bfr_before (
		.din(new_net_5324),
		.dout(new_net_5323)
	);

	bfr new_net_5325_bfr_before (
		.din(new_net_5325),
		.dout(new_net_5324)
	);

	bfr new_net_5326_bfr_before (
		.din(new_net_5326),
		.dout(new_net_5325)
	);

	spl2 _1745__v_fanout (
		.a(_1745_),
		.b(new_net_1914),
		.c(new_net_5326)
	);

	bfr new_net_5327_bfr_before (
		.din(new_net_5327),
		.dout(new_net_465)
	);

	bfr new_net_5328_bfr_before (
		.din(new_net_5328),
		.dout(new_net_5327)
	);

	bfr new_net_5329_bfr_before (
		.din(new_net_5329),
		.dout(new_net_5328)
	);

	bfr new_net_5330_bfr_before (
		.din(new_net_5330),
		.dout(new_net_5329)
	);

	spl2 _1118__v_fanout (
		.a(_1118_),
		.b(new_net_464),
		.c(new_net_5330)
	);

	bfr new_net_5331_bfr_after (
		.din(_0555_),
		.dout(new_net_5331)
	);

	bfr new_net_5332_bfr_after (
		.din(new_net_5331),
		.dout(new_net_5332)
	);

	bfr new_net_5333_bfr_after (
		.din(new_net_5332),
		.dout(new_net_5333)
	);

	bfr new_net_5334_bfr_after (
		.din(new_net_5333),
		.dout(new_net_5334)
	);

	spl2 _0555__v_fanout (
		.a(new_net_5334),
		.b(new_net_3051),
		.c(new_net_3052)
	);

	spl2 _0464__v_fanout (
		.a(_0464_),
		.b(new_net_2448),
		.c(new_net_2449)
	);

	bfr new_net_5335_bfr_before (
		.din(new_net_5335),
		.dout(new_net_1687)
	);

	bfr new_net_5336_bfr_before (
		.din(new_net_5336),
		.dout(new_net_5335)
	);

	bfr new_net_5337_bfr_before (
		.din(new_net_5337),
		.dout(new_net_5336)
	);

	bfr new_net_5338_bfr_before (
		.din(new_net_5338),
		.dout(new_net_5337)
	);

	spl2 _1066__v_fanout (
		.a(_1066_),
		.b(new_net_1686),
		.c(new_net_5338)
	);

	spl2 _0635__v_fanout (
		.a(_0635_),
		.b(new_net_1222),
		.c(new_net_1223)
	);

	bfr new_net_5339_bfr_before (
		.din(new_net_5339),
		.dout(new_net_1357)
	);

	bfr new_net_5340_bfr_before (
		.din(new_net_5340),
		.dout(new_net_5339)
	);

	bfr new_net_5341_bfr_before (
		.din(new_net_5341),
		.dout(new_net_5340)
	);

	bfr new_net_5342_bfr_before (
		.din(new_net_5342),
		.dout(new_net_5341)
	);

	spl2 _1255__v_fanout (
		.a(_1255_),
		.b(new_net_1356),
		.c(new_net_5342)
	);

	bfr new_net_5343_bfr_before (
		.din(new_net_5343),
		.dout(new_net_475)
	);

	bfr new_net_5344_bfr_before (
		.din(new_net_5344),
		.dout(new_net_5343)
	);

	bfr new_net_5345_bfr_before (
		.din(new_net_5345),
		.dout(new_net_5344)
	);

	bfr new_net_5346_bfr_before (
		.din(new_net_5346),
		.dout(new_net_5345)
	);

	spl2 _0025__v_fanout (
		.a(_0025_),
		.b(new_net_474),
		.c(new_net_5346)
	);

	bfr new_net_5347_bfr_before (
		.din(new_net_5347),
		.dout(new_net_2123)
	);

	bfr new_net_5348_bfr_before (
		.din(new_net_5348),
		.dout(new_net_5347)
	);

	bfr new_net_5349_bfr_before (
		.din(new_net_5349),
		.dout(new_net_5348)
	);

	bfr new_net_5350_bfr_before (
		.din(new_net_5350),
		.dout(new_net_5349)
	);

	spl2 _0140__v_fanout (
		.a(_0140_),
		.b(new_net_2122),
		.c(new_net_5350)
	);

	bfr new_net_5351_bfr_before (
		.din(new_net_5351),
		.dout(new_net_2237)
	);

	bfr new_net_5352_bfr_before (
		.din(new_net_5352),
		.dout(new_net_5351)
	);

	bfr new_net_5353_bfr_before (
		.din(new_net_5353),
		.dout(new_net_5352)
	);

	bfr new_net_5354_bfr_before (
		.din(new_net_5354),
		.dout(new_net_5353)
	);

	spl2 _1417__v_fanout (
		.a(_1417_),
		.b(new_net_2236),
		.c(new_net_5354)
	);

	bfr new_net_5355_bfr_before (
		.din(new_net_5355),
		.dout(new_net_2191)
	);

	bfr new_net_5356_bfr_before (
		.din(new_net_5356),
		.dout(new_net_5355)
	);

	bfr new_net_5357_bfr_before (
		.din(new_net_5357),
		.dout(new_net_5356)
	);

	bfr new_net_5358_bfr_before (
		.din(new_net_5358),
		.dout(new_net_5357)
	);

	spl2 _1626__v_fanout (
		.a(_1626_),
		.b(new_net_2190),
		.c(new_net_5358)
	);

	bfr new_net_5359_bfr_before (
		.din(new_net_5359),
		.dout(new_net_1506)
	);

	bfr new_net_5360_bfr_before (
		.din(new_net_5360),
		.dout(new_net_5359)
	);

	bfr new_net_5361_bfr_before (
		.din(new_net_5361),
		.dout(new_net_5360)
	);

	bfr new_net_5362_bfr_before (
		.din(new_net_5362),
		.dout(new_net_5361)
	);

	spl2 _0259__v_fanout (
		.a(_0259_),
		.b(new_net_1505),
		.c(new_net_5362)
	);

	spl2 _1515__v_fanout (
		.a(_1515_),
		.b(new_net_2979),
		.c(new_net_2980)
	);

	spl2 _0345__v_fanout (
		.a(_0345_),
		.b(new_net_2142),
		.c(new_net_2143)
	);

	spl2 _1820__v_fanout (
		.a(_1820_),
		.b(new_net_1622),
		.c(new_net_1623)
	);

	spl2 _0231__v_fanout (
		.a(_0231_),
		.b(new_net_279),
		.c(new_net_280)
	);

	spl2 _1625__v_fanout (
		.a(_1625_),
		.b(new_net_2156),
		.c(new_net_2157)
	);

	spl2 _0139__v_fanout (
		.a(_0139_),
		.b(new_net_1660),
		.c(new_net_1661)
	);

	spl2 _0024__v_fanout (
		.a(_0024_),
		.b(new_net_285),
		.c(new_net_286)
	);

	spl2 _1021__v_fanout (
		.a(_1021_),
		.b(new_net_1830),
		.c(new_net_1831)
	);

	spl2 _1117__v_fanout (
		.a(_1117_),
		.b(new_net_424),
		.c(new_net_425)
	);

	spl2 _1466__v_fanout (
		.a(_1466_),
		.b(new_net_940),
		.c(new_net_941)
	);

	spl2 _1254__v_fanout (
		.a(_1254_),
		.b(new_net_2430),
		.c(new_net_2431)
	);

	spl2 _0103__v_fanout (
		.a(_0103_),
		.b(new_net_1758),
		.c(new_net_1759)
	);

	spl2 _1287__v_fanout (
		.a(_1287_),
		.b(new_net_504),
		.c(new_net_505)
	);

	spl2 _0258__v_fanout (
		.a(_0258_),
		.b(new_net_1289),
		.c(new_net_1290)
	);

	bfr new_net_5363_bfr_before (
		.din(new_net_5363),
		.dout(new_net_2033)
	);

	bfr new_net_5364_bfr_before (
		.din(new_net_5364),
		.dout(new_net_5363)
	);

	bfr new_net_5365_bfr_before (
		.din(new_net_5365),
		.dout(new_net_5364)
	);

	bfr new_net_5366_bfr_before (
		.din(new_net_5366),
		.dout(new_net_5365)
	);

	spl2 _0462__v_fanout (
		.a(_0462_),
		.b(new_net_2032),
		.c(new_net_5366)
	);

	spl2 _1416__v_fanout (
		.a(_1416_),
		.b(new_net_2878),
		.c(new_net_2879)
	);

	spl2 _1331__v_fanout (
		.a(_1331_),
		.b(new_net_600),
		.c(new_net_601)
	);

	spl2 _1576__v_fanout (
		.a(_1576_),
		.b(new_net_2325),
		.c(new_net_2326)
	);

	spl2 _1210__v_fanout (
		.a(_1210_),
		.b(new_net_1034),
		.c(new_net_1035)
	);

	spl2 _1372__v_fanout (
		.a(_1372_),
		.b(new_net_2118),
		.c(new_net_2119)
	);

	spl2 _1177__v_fanout (
		.a(_1177_),
		.b(new_net_2716),
		.c(new_net_2717)
	);

	spl2 _1744__v_fanout (
		.a(_1744_),
		.b(new_net_1866),
		.c(new_net_1867)
	);

	spl2 _1073__v_fanout (
		.a(_1073_),
		.b(new_net_1922),
		.c(new_net_1923)
	);

	spl2 _0553__v_fanout (
		.a(_0553_),
		.b(new_net_2957),
		.c(new_net_2958)
	);

	spl2 _1065__v_fanout (
		.a(_1065_),
		.b(new_net_1650),
		.c(new_net_1651)
	);

	spl2 _1696__v_fanout (
		.a(_1696_),
		.b(new_net_3197),
		.c(new_net_3198)
	);

	spl2 _1133__v_fanout (
		.a(_1133_),
		.b(new_net_486),
		.c(new_net_487)
	);

	spl2 _1414__v_fanout (
		.a(_1414_),
		.b(new_net_2110),
		.c(new_net_2111)
	);

	spl2 _1063__v_fanout (
		.a(_1063_),
		.b(new_net_2292),
		.c(new_net_2293)
	);

	spl2 _1623__v_fanout (
		.a(_1623_),
		.b(new_net_2072),
		.c(new_net_2073)
	);

	spl2 _0137__v_fanout (
		.a(_0137_),
		.b(new_net_3151),
		.c(new_net_3152)
	);

	spl2 _0021__v_fanout (
		.a(_0021_),
		.b(new_net_2939),
		.c(new_net_2940)
	);

	spl2 _1252__v_fanout (
		.a(_1252_),
		.b(new_net_862),
		.c(new_net_863)
	);

	bfr new_net_5367_bfr_after (
		.din(_0364_),
		.dout(new_net_5367)
	);

	bfr new_net_5368_bfr_after (
		.din(new_net_5367),
		.dout(new_net_5368)
	);

	spl2 _0364__v_fanout (
		.a(new_net_5368),
		.b(new_net_558),
		.c(new_net_559)
	);

	spl2 _1329__v_fanout (
		.a(_1329_),
		.b(new_net_500),
		.c(new_net_501)
	);

	spl2 _0552__v_fanout (
		.a(_0552_),
		.b(new_net_805),
		.c(new_net_806)
	);

	spl2 _0451__v_fanout (
		.a(_0451_),
		.b(new_net_665),
		.c(new_net_666)
	);

	spl2 _1020__v_fanout (
		.a(_1020_),
		.b(new_net_1672),
		.c(new_net_1673)
	);

	spl2 _0256__v_fanout (
		.a(_0256_),
		.b(new_net_954),
		.c(new_net_955)
	);

	spl2 _1742__v_fanout (
		.a(_1742_),
		.b(new_net_2884),
		.c(new_net_2885)
	);

	spl2 _1115__v_fanout (
		.a(_1115_),
		.b(new_net_289),
		.c(new_net_290)
	);

	spl2 _1512__v_fanout (
		.a(_1512_),
		.b(new_net_1058),
		.c(new_net_1059)
	);

	spl2 _1175__v_fanout (
		.a(_1175_),
		.b(new_net_641),
		.c(new_net_642)
	);

	spl2 _1740__v_fanout (
		.a(_1740_),
		.b(new_net_1724),
		.c(new_net_1725)
	);

	spl2 _1114__v_fanout (
		.a(_1114_),
		.b(new_net_112),
		.c(new_net_113)
	);

	spl2 _0362__v_fanout (
		.a(_0362_),
		.b(new_net_472),
		.c(new_net_473)
	);

	spl2 _0136__v_fanout (
		.a(_0136_),
		.b(new_net_1086),
		.c(new_net_1087)
	);

	bfr new_net_5369_bfr_before (
		.din(new_net_5369),
		.dout(new_net_2818)
	);

	bfr new_net_5370_bfr_before (
		.din(new_net_5370),
		.dout(new_net_5369)
	);

	bfr new_net_5371_bfr_before (
		.din(new_net_5371),
		.dout(new_net_5370)
	);

	bfr new_net_5372_bfr_before (
		.din(new_net_5372),
		.dout(new_net_5371)
	);

	spl2 _0550__v_fanout (
		.a(_0550_),
		.b(new_net_2817),
		.c(new_net_5372)
	);

	spl2 _0255__v_fanout (
		.a(_0255_),
		.b(new_net_785),
		.c(new_net_786)
	);

	spl2 _0020__v_fanout (
		.a(_0020_),
		.b(new_net_234),
		.c(new_net_235)
	);

	spl2 _1413__v_fanout (
		.a(_1413_),
		.b(new_net_2272),
		.c(new_net_2273)
	);

	spl2 _1062__v_fanout (
		.a(_1062_),
		.b(new_net_2106),
		.c(new_net_2107)
	);

	spl2 _1622__v_fanout (
		.a(_1622_),
		.b(new_net_2078),
		.c(new_net_2079)
	);

	spl2 _1174__v_fanout (
		.a(_1174_),
		.b(new_net_454),
		.c(new_net_455)
	);

	spl2 _1251__v_fanout (
		.a(_1251_),
		.b(new_net_2309),
		.c(new_net_2310)
	);

	spl2 _1511__v_fanout (
		.a(_1511_),
		.b(new_net_2170),
		.c(new_net_2171)
	);

	spl2 _1328__v_fanout (
		.a(_1328_),
		.b(new_net_2246),
		.c(new_net_2247)
	);

	spl2 _1019__v_fanout (
		.a(_1019_),
		.b(new_net_1509),
		.c(new_net_1510)
	);

	bfr new_net_5373_bfr_before (
		.din(new_net_5373),
		.dout(new_net_2996)
	);

	bfr new_net_5374_bfr_before (
		.din(new_net_5374),
		.dout(new_net_5373)
	);

	bfr new_net_5375_bfr_before (
		.din(new_net_5375),
		.dout(new_net_5374)
	);

	bfr new_net_5376_bfr_before (
		.din(new_net_5376),
		.dout(new_net_5375)
	);

	spl2 _1016__v_fanout (
		.a(_1016_),
		.b(new_net_2995),
		.c(new_net_5376)
	);

	bfr new_net_5377_bfr_before (
		.din(new_net_5377),
		.dout(new_net_1983)
	);

	bfr new_net_5378_bfr_before (
		.din(new_net_5378),
		.dout(new_net_5377)
	);

	bfr new_net_5379_bfr_before (
		.din(new_net_5379),
		.dout(new_net_5378)
	);

	bfr new_net_5380_bfr_before (
		.din(new_net_5380),
		.dout(new_net_5379)
	);

	spl2 _1411__v_fanout (
		.a(_1411_),
		.b(new_net_1982),
		.c(new_net_5380)
	);

	bfr new_net_5381_bfr_before (
		.din(new_net_5381),
		.dout(new_net_977)
	);

	bfr new_net_5382_bfr_before (
		.din(new_net_5382),
		.dout(new_net_5381)
	);

	bfr new_net_5383_bfr_before (
		.din(new_net_5383),
		.dout(new_net_5382)
	);

	bfr new_net_5384_bfr_before (
		.din(new_net_5384),
		.dout(new_net_5383)
	);

	spl2 _1509__v_fanout (
		.a(_1509_),
		.b(new_net_976),
		.c(new_net_5384)
	);

	bfr new_net_5385_bfr_before (
		.din(new_net_5385),
		.dout(new_net_1849)
	);

	bfr new_net_5386_bfr_before (
		.din(new_net_5386),
		.dout(new_net_5385)
	);

	bfr new_net_5387_bfr_before (
		.din(new_net_5387),
		.dout(new_net_5386)
	);

	bfr new_net_5388_bfr_before (
		.din(new_net_5388),
		.dout(new_net_5387)
	);

	spl2 _1326__v_fanout (
		.a(_1326_),
		.b(new_net_1848),
		.c(new_net_5388)
	);

	bfr new_net_5389_bfr_before (
		.din(new_net_5389),
		.dout(new_net_3004)
	);

	bfr new_net_5390_bfr_before (
		.din(new_net_5390),
		.dout(new_net_5389)
	);

	bfr new_net_5391_bfr_before (
		.din(new_net_5391),
		.dout(new_net_5390)
	);

	bfr new_net_5392_bfr_before (
		.din(new_net_5392),
		.dout(new_net_5391)
	);

	spl2 _0134__v_fanout (
		.a(_0134_),
		.b(new_net_3003),
		.c(new_net_5392)
	);

	bfr new_net_5393_bfr_before (
		.din(new_net_5393),
		.dout(new_net_2952)
	);

	bfr new_net_5394_bfr_before (
		.din(new_net_5394),
		.dout(new_net_5393)
	);

	bfr new_net_5395_bfr_before (
		.din(new_net_5395),
		.dout(new_net_5394)
	);

	bfr new_net_5396_bfr_before (
		.din(new_net_5396),
		.dout(new_net_5395)
	);

	spl2 _1112__v_fanout (
		.a(_1112_),
		.b(new_net_2951),
		.c(new_net_5396)
	);

	bfr new_net_5397_bfr_before (
		.din(new_net_5397),
		.dout(new_net_1921)
	);

	bfr new_net_5398_bfr_before (
		.din(new_net_5398),
		.dout(new_net_5397)
	);

	bfr new_net_5399_bfr_before (
		.din(new_net_5399),
		.dout(new_net_5398)
	);

	bfr new_net_5400_bfr_before (
		.din(new_net_5400),
		.dout(new_net_5399)
	);

	spl2 _1619__v_fanout (
		.a(_1619_),
		.b(new_net_1920),
		.c(new_net_5400)
	);

	bfr new_net_5401_bfr_before (
		.din(new_net_5401),
		.dout(new_net_2485)
	);

	bfr new_net_5402_bfr_before (
		.din(new_net_5402),
		.dout(new_net_5401)
	);

	bfr new_net_5403_bfr_before (
		.din(new_net_5403),
		.dout(new_net_5402)
	);

	bfr new_net_5404_bfr_before (
		.din(new_net_5404),
		.dout(new_net_5403)
	);

	spl2 _1172__v_fanout (
		.a(_1172_),
		.b(new_net_2484),
		.c(new_net_5404)
	);

	bfr new_net_5405_bfr_before (
		.din(new_net_5405),
		.dout(new_net_2239)
	);

	bfr new_net_5406_bfr_before (
		.din(new_net_5406),
		.dout(new_net_5405)
	);

	bfr new_net_5407_bfr_before (
		.din(new_net_5407),
		.dout(new_net_5406)
	);

	bfr new_net_5408_bfr_before (
		.din(new_net_5408),
		.dout(new_net_5407)
	);

	spl2 _1249__v_fanout (
		.a(_1249_),
		.b(new_net_2238),
		.c(new_net_5408)
	);

	bfr new_net_5409_bfr_before (
		.din(new_net_5409),
		.dout(new_net_1081)
	);

	bfr new_net_5410_bfr_before (
		.din(new_net_5410),
		.dout(new_net_5409)
	);

	bfr new_net_5411_bfr_before (
		.din(new_net_5411),
		.dout(new_net_5410)
	);

	bfr new_net_5412_bfr_before (
		.din(new_net_5412),
		.dout(new_net_5411)
	);

	spl2 _0253__v_fanout (
		.a(_0253_),
		.b(new_net_1080),
		.c(new_net_5412)
	);

	bfr new_net_5413_bfr_before (
		.din(new_net_5413),
		.dout(new_net_1404)
	);

	bfr new_net_5414_bfr_before (
		.din(new_net_5414),
		.dout(new_net_5413)
	);

	bfr new_net_5415_bfr_before (
		.din(new_net_5415),
		.dout(new_net_5414)
	);

	bfr new_net_5416_bfr_before (
		.din(new_net_5416),
		.dout(new_net_5415)
	);

	spl2 _1060__v_fanout (
		.a(_1060_),
		.b(new_net_1403),
		.c(new_net_5416)
	);

	spl2 _0549__v_fanout (
		.a(_0549_),
		.b(new_net_2771),
		.c(new_net_2772)
	);

	bfr new_net_5417_bfr_after (
		.din(_0461_),
		.dout(new_net_5417)
	);

	bfr new_net_5418_bfr_after (
		.din(new_net_5417),
		.dout(new_net_5418)
	);

	bfr new_net_5419_bfr_after (
		.din(new_net_5418),
		.dout(new_net_5419)
	);

	bfr new_net_5420_bfr_after (
		.din(new_net_5419),
		.dout(new_net_5420)
	);

	spl2 _0461__v_fanout (
		.a(new_net_5420),
		.b(new_net_1854),
		.c(new_net_1855)
	);

	spl2 _0360__v_fanout (
		.a(_0360_),
		.b(new_net_374),
		.c(new_net_375)
	);

	bfr new_net_5421_bfr_before (
		.din(new_net_5421),
		.dout(new_net_2320)
	);

	bfr new_net_5422_bfr_before (
		.din(new_net_5422),
		.dout(new_net_5421)
	);

	bfr new_net_5423_bfr_before (
		.din(new_net_5423),
		.dout(new_net_5422)
	);

	bfr new_net_5424_bfr_before (
		.din(new_net_5424),
		.dout(new_net_5423)
	);

	spl2 _0018__v_fanout (
		.a(_0018_),
		.b(new_net_2319),
		.c(new_net_5424)
	);

	bfr new_net_5425_bfr_before (
		.din(new_net_5425),
		.dout(new_net_2089)
	);

	bfr new_net_5426_bfr_before (
		.din(new_net_5426),
		.dout(new_net_5425)
	);

	bfr new_net_5427_bfr_before (
		.din(new_net_5427),
		.dout(new_net_5426)
	);

	bfr new_net_5428_bfr_before (
		.din(new_net_5428),
		.dout(new_net_5427)
	);

	spl2 _1738__v_fanout (
		.a(_1738_),
		.b(new_net_2088),
		.c(new_net_5428)
	);

	spl2 _0233__v_fanout (
		.a(_0233_),
		.b(new_net_3031),
		.c(new_net_3032)
	);

	spl2 _1075__v_fanout (
		.a(_1075_),
		.b(new_net_733),
		.c(new_net_734)
	);

	spl2 _0105__v_fanout (
		.a(_0105_),
		.b(new_net_1838),
		.c(new_net_1839)
	);

	spl2 _1468__v_fanout (
		.a(_1468_),
		.b(new_net_1285),
		.c(new_net_1286)
	);

	spl2 _1737__v_fanout (
		.a(_1737_),
		.b(new_net_1890),
		.c(new_net_1891)
	);

	spl2 _0655__v_fanout (
		.a(_0655_),
		.b(new_net_1439),
		.c(new_net_1440)
	);

	spl2 _1135__v_fanout (
		.a(_1135_),
		.b(new_net_1072),
		.c(new_net_1073)
	);

	spl2 _1374__v_fanout (
		.a(_1374_),
		.b(new_net_2248),
		.c(new_net_2249)
	);

	spl2 _1212__v_fanout (
		.a(_1212_),
		.b(new_net_872),
		.c(new_net_873)
	);

	spl2 _1508__v_fanout (
		.a(_1508_),
		.b(new_net_1624),
		.c(new_net_1625)
	);

	spl2 _0133__v_fanout (
		.a(_0133_),
		.b(new_net_570),
		.c(new_net_571)
	);

	spl2 _1618__v_fanout (
		.a(_1618_),
		.b(new_net_1884),
		.c(new_net_1885)
	);

	spl2 _1699__v_fanout (
		.a(_1699_),
		.b(new_net_1764),
		.c(new_net_1765)
	);

	spl2 _1289__v_fanout (
		.a(_1289_),
		.b(new_net_2092),
		.c(new_net_2093)
	);

	spl2 _1023__v_fanout (
		.a(_1023_),
		.b(new_net_1158),
		.c(new_net_1159)
	);

	spl2 _1579__v_fanout (
		.a(_1579_),
		.b(new_net_2945),
		.c(new_net_2946)
	);

	spl2 _1015__v_fanout (
		.a(_1015_),
		.b(new_net_787),
		.c(new_net_788)
	);

	spl2 _0017__v_fanout (
		.a(_0017_),
		.b(new_net_130),
		.c(new_net_131)
	);

	spl2 _1248__v_fanout (
		.a(_1248_),
		.b(new_net_2200),
		.c(new_net_2201)
	);

	spl2 _0458__v_fanout (
		.a(_0458_),
		.b(new_net_946),
		.c(new_net_947)
	);

	spl2 _1325__v_fanout (
		.a(_1325_),
		.b(new_net_337),
		.c(new_net_338)
	);

	spl2 _1059__v_fanout (
		.a(_1059_),
		.b(new_net_1596),
		.c(new_net_1597)
	);

	spl2 _1822__v_fanout (
		.a(_1822_),
		.b(new_net_3071),
		.c(new_net_3072)
	);

	spl2 _1171__v_fanout (
		.a(_1171_),
		.b(new_net_2454),
		.c(new_net_2455)
	);

	spl2 _1410__v_fanout (
		.a(_1410_),
		.b(new_net_1944),
		.c(new_net_1945)
	);

	spl2 _1111__v_fanout (
		.a(_1111_),
		.b(new_net_2742),
		.c(new_net_2743)
	);

	bfr new_net_5429_bfr_before (
		.din(new_net_5429),
		.dout(new_net_724)
	);

	bfr new_net_5430_bfr_before (
		.din(new_net_5430),
		.dout(new_net_5429)
	);

	bfr new_net_5431_bfr_before (
		.din(new_net_5431),
		.dout(new_net_5430)
	);

	bfr new_net_5432_bfr_before (
		.din(new_net_5432),
		.dout(new_net_5431)
	);

	spl2 _0358__v_fanout (
		.a(_0358_),
		.b(new_net_723),
		.c(new_net_5432)
	);

	spl2 _1057__v_fanout (
		.a(_1057_),
		.b(new_net_1312),
		.c(new_net_1313)
	);

	spl2 _1408__v_fanout (
		.a(_1408_),
		.b(new_net_1328),
		.c(new_net_1329)
	);

	spl2 _1013__v_fanout (
		.a(_1013_),
		.b(new_net_2855),
		.c(new_net_2856)
	);

	spl2 _1246__v_fanout (
		.a(_1246_),
		.b(new_net_2895),
		.c(new_net_2896)
	);

	spl2 _0457__v_fanout (
		.a(_0457_),
		.b(new_net_902),
		.c(new_net_903)
	);

	bfr new_net_5433_bfr_after (
		.din(_0251_),
		.dout(new_net_5433)
	);

	bfr new_net_5434_bfr_after (
		.din(new_net_5433),
		.dout(new_net_5434)
	);

	spl2 _0251__v_fanout (
		.a(new_net_5434),
		.b(new_net_1012),
		.c(new_net_1013)
	);

	spl2 _0130__v_fanout (
		.a(_0130_),
		.b(new_net_2821),
		.c(new_net_2822)
	);

	spl2 _1109__v_fanout (
		.a(_1109_),
		.b(new_net_2333),
		.c(new_net_2334)
	);

	spl2 _1506__v_fanout (
		.a(_1506_),
		.b(new_net_878),
		.c(new_net_879)
	);

	spl2 _1616__v_fanout (
		.a(_1616_),
		.b(new_net_1788),
		.c(new_net_1789)
	);

	spl2 _1169__v_fanout (
		.a(_1169_),
		.b(new_net_2412),
		.c(new_net_2413)
	);

	spl2 _1323__v_fanout (
		.a(_1323_),
		.b(new_net_1298),
		.c(new_net_1299)
	);

	spl2 _0347__v_fanout (
		.a(_0347_),
		.b(new_net_2529),
		.c(new_net_2530)
	);

	spl2 _0644__v_fanout (
		.a(_0644_),
		.b(new_net_30),
		.c(new_net_31)
	);

	spl2 _1735__v_fanout (
		.a(_1735_),
		.b(new_net_3252),
		.c(new_net_3253)
	);

	spl2 _0015__v_fanout (
		.a(_0015_),
		.b(new_net_58),
		.c(new_net_59)
	);

	spl2 _1505__v_fanout (
		.a(_1505_),
		.b(new_net_844),
		.c(new_net_845)
	);

	spl2 _1108__v_fanout (
		.a(_1108_),
		.b(new_net_2138),
		.c(new_net_2139)
	);

	spl2 _1615__v_fanout (
		.a(_1615_),
		.b(new_net_1750),
		.c(new_net_1751)
	);

	spl2 _0633__v_fanout (
		.a(_0633_),
		.b(new_net_1156),
		.c(new_net_1157)
	);

	bfr new_net_5435_bfr_before (
		.din(new_net_5435),
		.dout(new_net_853)
	);

	bfr new_net_5436_bfr_before (
		.din(new_net_5436),
		.dout(new_net_5435)
	);

	bfr new_net_5437_bfr_before (
		.din(new_net_5437),
		.dout(new_net_5436)
	);

	bfr new_net_5438_bfr_before (
		.din(new_net_5438),
		.dout(new_net_5437)
	);

	spl2 _0455__v_fanout (
		.a(_0455_),
		.b(new_net_852),
		.c(new_net_5438)
	);

	spl2 _1322__v_fanout (
		.a(_1322_),
		.b(new_net_236),
		.c(new_net_237)
	);

	spl2 _1407__v_fanout (
		.a(_1407_),
		.b(new_net_1134),
		.c(new_net_1135)
	);

	spl2 _0014__v_fanout (
		.a(_0014_),
		.b(new_net_22),
		.c(new_net_23)
	);

	spl2 _1168__v_fanout (
		.a(_1168_),
		.b(new_net_2357),
		.c(new_net_2358)
	);

	spl2 _1010__v_fanout (
		.a(_1010_),
		.b(new_net_3041),
		.c(new_net_3042)
	);

	spl2 _1734__v_fanout (
		.a(_1734_),
		.b(new_net_3195),
		.c(new_net_3196)
	);

	spl2 _0129__v_fanout (
		.a(_0129_),
		.b(new_net_3033),
		.c(new_net_3034)
	);

	spl2 _0249__v_fanout (
		.a(_0249_),
		.b(new_net_2799),
		.c(new_net_2800)
	);

	spl2 _1245__v_fanout (
		.a(_1245_),
		.b(new_net_2693),
		.c(new_net_2694)
	);

	spl2 _1056__v_fanout (
		.a(_1056_),
		.b(new_net_1004),
		.c(new_net_1005)
	);

	spl2 _0454__v_fanout (
		.a(_0454_),
		.b(new_net_580),
		.c(new_net_581)
	);

	bfr new_net_5439_bfr_before (
		.din(new_net_5439),
		.dout(new_net_833)
	);

	bfr new_net_5440_bfr_before (
		.din(new_net_5440),
		.dout(new_net_5439)
	);

	bfr new_net_5441_bfr_before (
		.din(new_net_5441),
		.dout(new_net_5440)
	);

	bfr new_net_5442_bfr_before (
		.din(new_net_5442),
		.dout(new_net_5441)
	);

	spl2 _1405__v_fanout (
		.a(_1405_),
		.b(new_net_832),
		.c(new_net_5442)
	);

	spl2 _0248__v_fanout (
		.a(_0248_),
		.b(new_net_942),
		.c(new_net_943)
	);

	bfr new_net_5443_bfr_before (
		.din(new_net_5443),
		.dout(new_net_1532)
	);

	bfr new_net_5444_bfr_before (
		.din(new_net_5444),
		.dout(new_net_5443)
	);

	bfr new_net_5445_bfr_before (
		.din(new_net_5445),
		.dout(new_net_5444)
	);

	bfr new_net_5446_bfr_before (
		.din(new_net_5446),
		.dout(new_net_5445)
	);

	spl2 _0012__v_fanout (
		.a(_0012_),
		.b(new_net_1531),
		.c(new_net_5446)
	);

	bfr new_net_5447_bfr_before (
		.din(new_net_5447),
		.dout(new_net_794)
	);

	bfr new_net_5448_bfr_before (
		.din(new_net_5448),
		.dout(new_net_5447)
	);

	bfr new_net_5449_bfr_before (
		.din(new_net_5449),
		.dout(new_net_5448)
	);

	bfr new_net_5450_bfr_before (
		.din(new_net_5450),
		.dout(new_net_5449)
	);

	spl2 _1320__v_fanout (
		.a(_1320_),
		.b(new_net_793),
		.c(new_net_5450)
	);

	bfr new_net_5451_bfr_before (
		.din(new_net_5451),
		.dout(new_net_2105)
	);

	bfr new_net_5452_bfr_before (
		.din(new_net_5452),
		.dout(new_net_5451)
	);

	bfr new_net_5453_bfr_before (
		.din(new_net_5453),
		.dout(new_net_5452)
	);

	bfr new_net_5454_bfr_before (
		.din(new_net_5454),
		.dout(new_net_5453)
	);

	spl2 _1166__v_fanout (
		.a(_1166_),
		.b(new_net_2104),
		.c(new_net_5454)
	);

	bfr new_net_5455_bfr_before (
		.din(new_net_5455),
		.dout(new_net_2279)
	);

	bfr new_net_5456_bfr_before (
		.din(new_net_5456),
		.dout(new_net_5455)
	);

	bfr new_net_5457_bfr_before (
		.din(new_net_5457),
		.dout(new_net_5456)
	);

	bfr new_net_5458_bfr_before (
		.din(new_net_5458),
		.dout(new_net_5457)
	);

	spl2 _1243__v_fanout (
		.a(_1243_),
		.b(new_net_2278),
		.c(new_net_5458)
	);

	bfr new_net_5459_bfr_before (
		.din(new_net_5459),
		.dout(new_net_3114)
	);

	bfr new_net_5460_bfr_before (
		.din(new_net_5460),
		.dout(new_net_5459)
	);

	bfr new_net_5461_bfr_before (
		.din(new_net_5461),
		.dout(new_net_5460)
	);

	bfr new_net_5462_bfr_before (
		.din(new_net_5462),
		.dout(new_net_5461)
	);

	spl2 _1732__v_fanout (
		.a(_1732_),
		.b(new_net_3113),
		.c(new_net_5462)
	);

	bfr new_net_5463_bfr_before (
		.din(new_net_5463),
		.dout(new_net_302)
	);

	bfr new_net_5464_bfr_before (
		.din(new_net_5464),
		.dout(new_net_5463)
	);

	bfr new_net_5465_bfr_before (
		.din(new_net_5465),
		.dout(new_net_5464)
	);

	bfr new_net_5466_bfr_before (
		.din(new_net_5466),
		.dout(new_net_5465)
	);

	spl2 _0601__v_fanout (
		.a(_0601_),
		.b(new_net_301),
		.c(new_net_5466)
	);

	bfr new_net_5467_bfr_before (
		.din(new_net_5467),
		.dout(new_net_1185)
	);

	bfr new_net_5468_bfr_before (
		.din(new_net_5468),
		.dout(new_net_5467)
	);

	bfr new_net_5469_bfr_before (
		.din(new_net_5469),
		.dout(new_net_5468)
	);

	bfr new_net_5470_bfr_before (
		.din(new_net_5470),
		.dout(new_net_5469)
	);

	spl2 _1054__v_fanout (
		.a(_1054_),
		.b(new_net_1184),
		.c(new_net_5470)
	);

	bfr new_net_5471_bfr_before (
		.din(new_net_5471),
		.dout(new_net_411)
	);

	bfr new_net_5472_bfr_before (
		.din(new_net_5472),
		.dout(new_net_5471)
	);

	bfr new_net_5473_bfr_before (
		.din(new_net_5473),
		.dout(new_net_5472)
	);

	bfr new_net_5474_bfr_before (
		.din(new_net_5474),
		.dout(new_net_5473)
	);

	spl2 _1613__v_fanout (
		.a(_1613_),
		.b(new_net_410),
		.c(new_net_5474)
	);

	bfr new_net_5475_bfr_before (
		.din(new_net_5475),
		.dout(new_net_2217)
	);

	bfr new_net_5476_bfr_before (
		.din(new_net_5476),
		.dout(new_net_5475)
	);

	bfr new_net_5477_bfr_before (
		.din(new_net_5477),
		.dout(new_net_5476)
	);

	bfr new_net_5478_bfr_before (
		.din(new_net_5478),
		.dout(new_net_5477)
	);

	spl2 _0989__v_fanout (
		.a(_0989_),
		.b(new_net_2216),
		.c(new_net_5478)
	);

	bfr new_net_5479_bfr_before (
		.din(new_net_5479),
		.dout(new_net_684)
	);

	bfr new_net_5480_bfr_before (
		.din(new_net_5480),
		.dout(new_net_5479)
	);

	bfr new_net_5481_bfr_before (
		.din(new_net_5481),
		.dout(new_net_5480)
	);

	bfr new_net_5482_bfr_before (
		.din(new_net_5482),
		.dout(new_net_5481)
	);

	spl2 _1503__v_fanout (
		.a(_1503_),
		.b(new_net_683),
		.c(new_net_5482)
	);

	bfr new_net_5483_bfr_before (
		.din(new_net_5483),
		.dout(new_net_2628)
	);

	bfr new_net_5484_bfr_before (
		.din(new_net_5484),
		.dout(new_net_5483)
	);

	bfr new_net_5485_bfr_before (
		.din(new_net_5485),
		.dout(new_net_5484)
	);

	bfr new_net_5486_bfr_before (
		.din(new_net_5486),
		.dout(new_net_5485)
	);

	spl2 _0127__v_fanout (
		.a(_0127_),
		.b(new_net_2627),
		.c(new_net_5486)
	);

	bfr new_net_5487_bfr_before (
		.din(new_net_5487),
		.dout(new_net_33)
	);

	bfr new_net_5488_bfr_before (
		.din(new_net_5488),
		.dout(new_net_5487)
	);

	bfr new_net_5489_bfr_before (
		.din(new_net_5489),
		.dout(new_net_5488)
	);

	bfr new_net_5490_bfr_before (
		.din(new_net_5490),
		.dout(new_net_5489)
	);

	spl2 _1106__v_fanout (
		.a(_1106_),
		.b(new_net_32),
		.c(new_net_5490)
	);

	bfr new_net_5491_bfr_after (
		.din(_0357_),
		.dout(new_net_5491)
	);

	bfr new_net_5492_bfr_after (
		.din(new_net_5491),
		.dout(new_net_5492)
	);

	bfr new_net_5493_bfr_after (
		.din(new_net_5492),
		.dout(new_net_5493)
	);

	bfr new_net_5494_bfr_after (
		.din(new_net_5493),
		.dout(new_net_5494)
	);

	spl2 _0357__v_fanout (
		.a(new_net_5494),
		.b(new_net_281),
		.c(new_net_282)
	);

	spl2 _0677__v_fanout (
		.a(_0677_),
		.b(new_net_2418),
		.c(new_net_2419)
	);

	spl2 _0285__v_fanout (
		.a(_0285_),
		.b(new_net_1770),
		.c(new_net_1771)
	);

	spl2 _1319__v_fanout (
		.a(_1319_),
		.b(new_net_128),
		.c(new_net_129)
	);

	spl2 _1025__v_fanout (
		.a(_1025_),
		.b(new_net_1584),
		.c(new_net_1585)
	);

	spl2 _0107__v_fanout (
		.a(_0107_),
		.b(new_net_1992),
		.c(new_net_1993)
	);

	spl2 _0010__v_fanout (
		.a(_0010_),
		.b(new_net_1427),
		.c(new_net_1428)
	);

	spl2 _0979__v_fanout (
		.a(_0979_),
		.b(new_net_3262),
		.c(new_net_3263)
	);

	spl2 _1581__v_fanout (
		.a(_1581_),
		.b(new_net_2070),
		.c(new_net_2071)
	);

	spl2 _1291__v_fanout (
		.a(_1291_),
		.b(new_net_2478),
		.c(new_net_2479)
	);

	spl2 _1404__v_fanout (
		.a(_1404_),
		.b(new_net_1726),
		.c(new_net_1727)
	);

	spl2 _1376__v_fanout (
		.a(_1376_),
		.b(new_net_2653),
		.c(new_net_2654)
	);

	spl2 _0355__v_fanout (
		.a(_0355_),
		.b(new_net_196),
		.c(new_net_197)
	);

	spl2 _1612__v_fanout (
		.a(_1612_),
		.b(new_net_220),
		.c(new_net_221)
	);

	spl2 _1077__v_fanout (
		.a(_1077_),
		.b(new_net_2066),
		.c(new_net_2067)
	);

	spl2 _1105__v_fanout (
		.a(_1105_),
		.b(new_net_3248),
		.c(new_net_3249)
	);

	spl2 _1053__v_fanout (
		.a(_1053_),
		.b(new_net_450),
		.c(new_net_451)
	);

	spl2 _1501__v_fanout (
		.a(_1501_),
		.b(new_net_295),
		.c(new_net_296)
	);

	spl2 _1701__v_fanout (
		.a(_1701_),
		.b(new_net_1832),
		.c(new_net_1833)
	);

	spl2 _1471__v_fanout (
		.a(_1471_),
		.b(new_net_1818),
		.c(new_net_1819)
	);

	bfr new_net_5495_bfr_before (
		.din(new_net_5495),
		.dout(new_net_2221)
	);

	bfr new_net_5496_bfr_before (
		.din(new_net_5496),
		.dout(new_net_5495)
	);

	bfr new_net_5497_bfr_before (
		.din(new_net_5497),
		.dout(new_net_5496)
	);

	bfr new_net_5498_bfr_before (
		.din(new_net_5498),
		.dout(new_net_5497)
	);

	spl2 _0246__v_fanout (
		.a(_0246_),
		.b(new_net_2220),
		.c(new_net_5498)
	);

	spl2 _1242__v_fanout (
		.a(_1242_),
		.b(new_net_1952),
		.c(new_net_1953)
	);

	spl2 _0590__v_fanout (
		.a(_0590_),
		.b(new_net_2761),
		.c(new_net_2762)
	);

	spl2 _1137__v_fanout (
		.a(_1137_),
		.b(new_net_1202),
		.c(new_net_1203)
	);

	spl2 _1165__v_fanout (
		.a(_1165_),
		.b(new_net_2240),
		.c(new_net_2241)
	);

	spl2 _1824__v_fanout (
		.a(_1824_),
		.b(new_net_192),
		.c(new_net_193)
	);

	spl2 _1731__v_fanout (
		.a(_1731_),
		.b(new_net_3043),
		.c(new_net_3044)
	);

	spl2 _1214__v_fanout (
		.a(_1214_),
		.b(new_net_1768),
		.c(new_net_1769)
	);

	spl2 _0958__v_fanout (
		.a(_0958_),
		.b(new_net_358),
		.c(new_net_359)
	);

	spl2 _1240__v_fanout (
		.a(_1240_),
		.b(new_net_1716),
		.c(new_net_1717)
	);

	spl2 _1103__v_fanout (
		.a(_1103_),
		.b(new_net_3147),
		.c(new_net_3148)
	);

	spl2 _1499__v_fanout (
		.a(_1499_),
		.b(new_net_3199),
		.c(new_net_3200)
	);

	spl2 _0274__v_fanout (
		.a(_0274_),
		.b(new_net_2985),
		.c(new_net_2986)
	);

	spl2 _0354__v_fanout (
		.a(_0354_),
		.b(new_net_170),
		.c(new_net_171)
	);

	spl2 _0235__v_fanout (
		.a(_0235_),
		.b(new_net_180),
		.c(new_net_181)
	);

	spl2 _1609__v_fanout (
		.a(_1609_),
		.b(new_net_2148),
		.c(new_net_2149)
	);

	spl2 _1051__v_fanout (
		.a(_1051_),
		.b(new_net_1076),
		.c(new_net_1077)
	);

	spl2 _1317__v_fanout (
		.a(_1317_),
		.b(new_net_68),
		.c(new_net_69)
	);

	spl2 _0008__v_fanout (
		.a(_0008_),
		.b(new_net_1336),
		.c(new_net_1337)
	);

	spl2 _1163__v_fanout (
		.a(_1163_),
		.b(new_net_1594),
		.c(new_net_1595)
	);

	bfr new_net_5499_bfr_after (
		.din(_0126_),
		.dout(new_net_5499)
	);

	bfr new_net_5500_bfr_after (
		.din(new_net_5499),
		.dout(new_net_5500)
	);

	spl2 _0126__v_fanout (
		.a(new_net_5500),
		.b(new_net_2665),
		.c(new_net_2666)
	);

	spl2 _0568__v_fanout (
		.a(_0568_),
		.b(new_net_1878),
		.c(new_net_1879)
	);

	spl2 _1402__v_fanout (
		.a(_1402_),
		.b(new_net_1692),
		.c(new_net_1693)
	);

	spl2 _1728__v_fanout (
		.a(_1728_),
		.b(new_net_2763),
		.c(new_net_2764)
	);

	spl2 _1162__v_fanout (
		.a(_1162_),
		.b(new_net_1358),
		.c(new_net_1359)
	);

	spl2 _1239__v_fanout (
		.a(_1239_),
		.b(new_net_1842),
		.c(new_net_1843)
	);

	spl2 _0007__v_fanout (
		.a(_0007_),
		.b(new_net_1314),
		.c(new_net_1315)
	);

	spl2 _1608__v_fanout (
		.a(_1608_),
		.b(new_net_1936),
		.c(new_net_1937)
	);

	spl2 _1050__v_fanout (
		.a(_1050_),
		.b(new_net_3135),
		.c(new_net_3136)
	);

	spl2 _1316__v_fanout (
		.a(_1316_),
		.b(new_net_10),
		.c(new_net_11)
	);

	spl2 _1727__v_fanout (
		.a(_1727_),
		.b(new_net_2853),
		.c(new_net_2854)
	);

	spl2 _0557__v_fanout (
		.a(_0557_),
		.b(new_net_3141),
		.c(new_net_3142)
	);

	bfr new_net_5501_bfr_before (
		.din(new_net_5501),
		.dout(new_net_2768)
	);

	bfr new_net_5502_bfr_before (
		.din(new_net_5502),
		.dout(new_net_5501)
	);

	bfr new_net_5503_bfr_before (
		.din(new_net_5503),
		.dout(new_net_5502)
	);

	bfr new_net_5504_bfr_before (
		.din(new_net_5504),
		.dout(new_net_5503)
	);

	spl2 _0352__v_fanout (
		.a(_0352_),
		.b(new_net_2767),
		.c(new_net_5504)
	);

	spl2 _1102__v_fanout (
		.a(_1102_),
		.b(new_net_2625),
		.c(new_net_2626)
	);

	spl2 _0124__v_fanout (
		.a(_0124_),
		.b(new_net_2589),
		.c(new_net_2590)
	);

	spl2 _0263__v_fanout (
		.a(_0263_),
		.b(new_net_1485),
		.c(new_net_1486)
	);

	spl2 _1401__v_fanout (
		.a(_1401_),
		.b(new_net_1644),
		.c(new_net_1645)
	);

	spl2 _0947__v_fanout (
		.a(_0947_),
		.b(new_net_138),
		.c(new_net_139)
	);

	spl2 _1498__v_fanout (
		.a(_1498_),
		.b(new_net_560),
		.c(new_net_561)
	);

	spl2 _0351__v_fanout (
		.a(_0351_),
		.b(new_net_70),
		.c(new_net_71)
	);

	bfr new_net_5505_bfr_before (
		.din(new_net_5505),
		.dout(new_net_2568)
	);

	bfr new_net_5506_bfr_before (
		.din(new_net_5506),
		.dout(new_net_5505)
	);

	bfr new_net_5507_bfr_before (
		.din(new_net_5507),
		.dout(new_net_5506)
	);

	bfr new_net_5508_bfr_before (
		.din(new_net_5508),
		.dout(new_net_5507)
	);

	spl2 _1496__v_fanout (
		.a(_1496_),
		.b(new_net_2567),
		.c(new_net_5508)
	);

	bfr new_net_5509_bfr_before (
		.din(new_net_5509),
		.dout(new_net_2421)
	);

	bfr new_net_5510_bfr_before (
		.din(new_net_5510),
		.dout(new_net_5509)
	);

	bfr new_net_5511_bfr_before (
		.din(new_net_5511),
		.dout(new_net_5510)
	);

	bfr new_net_5512_bfr_before (
		.din(new_net_5512),
		.dout(new_net_5511)
	);

	spl2 _0230__v_fanout (
		.a(_0230_),
		.b(new_net_2420),
		.c(new_net_5512)
	);

	bfr new_net_5513_bfr_before (
		.din(new_net_5513),
		.dout(new_net_346)
	);

	bfr new_net_5514_bfr_before (
		.din(new_net_5514),
		.dout(new_net_5513)
	);

	bfr new_net_5515_bfr_before (
		.din(new_net_5515),
		.dout(new_net_5514)
	);

	bfr new_net_5516_bfr_before (
		.din(new_net_5516),
		.dout(new_net_5515)
	);

	spl2 _0925__v_fanout (
		.a(_0925_),
		.b(new_net_345),
		.c(new_net_5516)
	);

	bfr new_net_5517_bfr_before (
		.din(new_net_5517),
		.dout(new_net_1540)
	);

	bfr new_net_5518_bfr_before (
		.din(new_net_5518),
		.dout(new_net_5517)
	);

	bfr new_net_5519_bfr_before (
		.din(new_net_5519),
		.dout(new_net_5518)
	);

	bfr new_net_5520_bfr_before (
		.din(new_net_5520),
		.dout(new_net_5519)
	);

	spl2 _1314__v_fanout (
		.a(_1314_),
		.b(new_net_1539),
		.c(new_net_5520)
	);

	spl2 _0123__v_fanout (
		.a(_0123_),
		.b(new_net_1814),
		.c(new_net_1815)
	);

	bfr new_net_5521_bfr_before (
		.din(new_net_5521),
		.dout(new_net_1163)
	);

	bfr new_net_5522_bfr_before (
		.din(new_net_5522),
		.dout(new_net_5521)
	);

	bfr new_net_5523_bfr_before (
		.din(new_net_5523),
		.dout(new_net_5522)
	);

	bfr new_net_5524_bfr_before (
		.din(new_net_5524),
		.dout(new_net_5523)
	);

	spl2 _1237__v_fanout (
		.a(_1237_),
		.b(new_net_1162),
		.c(new_net_5524)
	);

	bfr new_net_5525_bfr_before (
		.din(new_net_5525),
		.dout(new_net_2213)
	);

	bfr new_net_5526_bfr_before (
		.din(new_net_5526),
		.dout(new_net_5525)
	);

	bfr new_net_5527_bfr_before (
		.din(new_net_5527),
		.dout(new_net_5526)
	);

	bfr new_net_5528_bfr_before (
		.din(new_net_5528),
		.dout(new_net_5527)
	);

	spl2 _1100__v_fanout (
		.a(_1100_),
		.b(new_net_2212),
		.c(new_net_5528)
	);

	bfr new_net_5529_bfr_before (
		.din(new_net_5529),
		.dout(new_net_1001)
	);

	bfr new_net_5530_bfr_before (
		.din(new_net_5530),
		.dout(new_net_5529)
	);

	bfr new_net_5531_bfr_before (
		.din(new_net_5531),
		.dout(new_net_5530)
	);

	bfr new_net_5532_bfr_before (
		.din(new_net_5532),
		.dout(new_net_5531)
	);

	spl2 _1048__v_fanout (
		.a(_1048_),
		.b(new_net_1000),
		.c(new_net_5532)
	);

	bfr new_net_5533_bfr_before (
		.din(new_net_5533),
		.dout(new_net_1197)
	);

	bfr new_net_5534_bfr_before (
		.din(new_net_5534),
		.dout(new_net_5533)
	);

	bfr new_net_5535_bfr_before (
		.din(new_net_5535),
		.dout(new_net_5534)
	);

	bfr new_net_5536_bfr_before (
		.din(new_net_5536),
		.dout(new_net_5535)
	);

	spl2 _0005__v_fanout (
		.a(_0005_),
		.b(new_net_1196),
		.c(new_net_5536)
	);

	bfr new_net_5537_bfr_before (
		.din(new_net_5537),
		.dout(new_net_3255)
	);

	bfr new_net_5538_bfr_before (
		.din(new_net_5538),
		.dout(new_net_5537)
	);

	bfr new_net_5539_bfr_before (
		.din(new_net_5539),
		.dout(new_net_5538)
	);

	bfr new_net_5540_bfr_before (
		.din(new_net_5540),
		.dout(new_net_5539)
	);

	spl2 _1399__v_fanout (
		.a(_1399_),
		.b(new_net_3254),
		.c(new_net_5540)
	);

	bfr new_net_5541_bfr_before (
		.din(new_net_5541),
		.dout(new_net_2173)
	);

	bfr new_net_5542_bfr_before (
		.din(new_net_5542),
		.dout(new_net_5541)
	);

	bfr new_net_5543_bfr_before (
		.din(new_net_5543),
		.dout(new_net_5542)
	);

	bfr new_net_5544_bfr_before (
		.din(new_net_5544),
		.dout(new_net_5543)
	);

	spl2 _1725__v_fanout (
		.a(_1725_),
		.b(new_net_2172),
		.c(new_net_5544)
	);

	bfr new_net_5545_bfr_before (
		.din(new_net_5545),
		.dout(new_net_1003)
	);

	bfr new_net_5546_bfr_before (
		.din(new_net_5546),
		.dout(new_net_5545)
	);

	bfr new_net_5547_bfr_before (
		.din(new_net_5547),
		.dout(new_net_5546)
	);

	bfr new_net_5548_bfr_before (
		.din(new_net_5548),
		.dout(new_net_5547)
	);

	spl2 _1160__v_fanout (
		.a(_1160_),
		.b(new_net_1002),
		.c(new_net_5548)
	);

	bfr new_net_5549_bfr_before (
		.din(new_net_5549),
		.dout(new_net_1609)
	);

	bfr new_net_5550_bfr_before (
		.din(new_net_5550),
		.dout(new_net_5549)
	);

	bfr new_net_5551_bfr_before (
		.din(new_net_5551),
		.dout(new_net_5550)
	);

	bfr new_net_5552_bfr_before (
		.din(new_net_5552),
		.dout(new_net_5551)
	);

	spl2 _1606__v_fanout (
		.a(_1606_),
		.b(new_net_1608),
		.c(new_net_5552)
	);

	bfr new_net_5553_bfr_after (
		.din(_0245_),
		.dout(new_net_5553)
	);

	bfr new_net_5554_bfr_after (
		.din(new_net_5553),
		.dout(new_net_5554)
	);

	bfr new_net_5555_bfr_after (
		.din(new_net_5554),
		.dout(new_net_5555)
	);

	bfr new_net_5556_bfr_after (
		.din(new_net_5555),
		.dout(new_net_5556)
	);

	spl2 _0245__v_fanout (
		.a(new_net_5556),
		.b(new_net_2004),
		.c(new_net_2005)
	);

	bfr new_net_5557_bfr_before (
		.din(new_net_5557),
		.dout(new_net_796)
	);

	bfr new_net_5558_bfr_before (
		.din(new_net_5558),
		.dout(new_net_5557)
	);

	bfr new_net_5559_bfr_before (
		.din(new_net_5559),
		.dout(new_net_5558)
	);

	bfr new_net_5560_bfr_before (
		.din(new_net_5560),
		.dout(new_net_5559)
	);

	spl2 _0535__v_fanout (
		.a(_0535_),
		.b(new_net_795),
		.c(new_net_5560)
	);

	spl2 _0243__v_fanout (
		.a(_0243_),
		.b(new_net_759),
		.c(new_net_760)
	);

	spl2 _0307__v_fanout (
		.a(_0307_),
		.b(new_net_2769),
		.c(new_net_2770)
	);

	spl2 _0000__v_fanout (
		.a(_0000_),
		.b(new_net_890),
		.c(new_net_891)
	);

	spl2 _1293__v_fanout (
		.a(_1293_),
		.b(new_net_2888),
		.c(new_net_2889)
	);

	spl2 _1605__v_fanout (
		.a(_1605_),
		.b(new_net_1392),
		.c(new_net_1393)
	);

	spl2 _1495__v_fanout (
		.a(_1495_),
		.b(new_net_2372),
		.c(new_net_2373)
	);

	spl2 _1236__v_fanout (
		.a(_1236_),
		.b(new_net_1734),
		.c(new_net_1735)
	);

	spl2 _1216__v_fanout (
		.a(_1216_),
		.b(new_net_2174),
		.c(new_net_2175)
	);

	spl2 _1398__v_fanout (
		.a(_1398_),
		.b(new_net_360),
		.c(new_net_361)
	);

	spl2 _1378__v_fanout (
		.a(_1378_),
		.b(new_net_3067),
		.c(new_net_3068)
	);

	spl2 _1313__v_fanout (
		.a(_1313_),
		.b(new_net_244),
		.c(new_net_245)
	);

	spl2 _0698__v_fanout (
		.a(_0698_),
		.b(new_net_470),
		.c(new_net_471)
	);

	spl2 _1099__v_fanout (
		.a(_1099_),
		.b(new_net_2969),
		.c(new_net_2970)
	);

	spl2 _1703__v_fanout (
		.a(_1703_),
		.b(new_net_1200),
		.c(new_net_1201)
	);

	spl2 _1079__v_fanout (
		.a(_1079_),
		.b(new_net_1457),
		.c(new_net_1458)
	);

	spl2 _1027__v_fanout (
		.a(_1027_),
		.b(new_net_1894),
		.c(new_net_1895)
	);

	spl2 _0525__v_fanout (
		.a(_0525_),
		.b(new_net_2006),
		.c(new_net_2007)
	);

	spl2 _1139__v_fanout (
		.a(_1139_),
		.b(new_net_1206),
		.c(new_net_1207)
	);

	bfr new_net_5561_bfr_before (
		.din(new_net_5561),
		.dout(new_net_2433)
	);

	bfr new_net_5562_bfr_before (
		.din(new_net_5562),
		.dout(new_net_5561)
	);

	bfr new_net_5563_bfr_before (
		.din(new_net_5563),
		.dout(new_net_5562)
	);

	bfr new_net_5564_bfr_before (
		.din(new_net_5564),
		.dout(new_net_5563)
	);

	spl2 _0120__v_fanout (
		.a(_0120_),
		.b(new_net_2432),
		.c(new_net_5564)
	);

	spl2 _1826__v_fanout (
		.a(_1826_),
		.b(new_net_588),
		.c(new_net_589)
	);

	spl2 _1473__v_fanout (
		.a(_1473_),
		.b(new_net_2218),
		.c(new_net_2219)
	);

	spl2 _0915__v_fanout (
		.a(_0915_),
		.b(new_net_757),
		.c(new_net_758)
	);

	spl2 _0219__v_fanout (
		.a(_0219_),
		.b(new_net_2949),
		.c(new_net_2950)
	);

	spl2 _1047__v_fanout (
		.a(_1047_),
		.b(new_net_968),
		.c(new_net_969)
	);

	spl2 _1159__v_fanout (
		.a(_1159_),
		.b(new_net_1986),
		.c(new_net_1987)
	);

	spl2 _1724__v_fanout (
		.a(_1724_),
		.b(new_net_1958),
		.c(new_net_1959)
	);

	spl2 _1583__v_fanout (
		.a(_1583_),
		.b(new_net_2162),
		.c(new_net_2163)
	);

	spl2 _0893__v_fanout (
		.a(_0893_),
		.b(new_net_3143),
		.c(new_net_3144)
	);

	spl2 _1796__v_fanout (
		.a(_1796_),
		.b(new_net_707),
		.c(new_net_708)
	);

	spl2 _1234__v_fanout (
		.a(_1234_),
		.b(new_net_1678),
		.c(new_net_1679)
	);

	spl2 _1603__v_fanout (
		.a(_1603_),
		.b(new_net_2959),
		.c(new_net_2960)
	);

	spl2 _1722__v_fanout (
		.a(_1722_),
		.b(new_net_1628),
		.c(new_net_1629)
	);

	spl2 _0198__v_fanout (
		.a(_0198_),
		.b(new_net_2194),
		.c(new_net_2195)
	);

	spl2 _0503__v_fanout (
		.a(_0503_),
		.b(new_net_356),
		.c(new_net_357)
	);

	spl2 _1311__v_fanout (
		.a(_1311_),
		.b(new_net_3133),
		.c(new_net_3134)
	);

	spl2 _1157__v_fanout (
		.a(_1157_),
		.b(new_net_448),
		.c(new_net_449)
	);

	bfr new_net_5565_bfr_after (
		.din(_0004_),
		.dout(new_net_5565)
	);

	bfr new_net_5566_bfr_after (
		.din(new_net_5565),
		.dout(new_net_5566)
	);

	spl2 _0004__v_fanout (
		.a(new_net_5566),
		.b(new_net_1132),
		.c(new_net_1133)
	);

	spl2 _0242__v_fanout (
		.a(_0242_),
		.b(new_net_709),
		.c(new_net_710)
	);

	spl2 _1097__v_fanout (
		.a(_1097_),
		.b(new_net_2849),
		.c(new_net_2850)
	);

	spl2 _0109__v_fanout (
		.a(_0109_),
		.b(new_net_1974),
		.c(new_net_1975)
	);

	spl2 _1493__v_fanout (
		.a(_1493_),
		.b(new_net_1938),
		.c(new_net_1939)
	);

	spl2 _1045__v_fanout (
		.a(_1045_),
		.b(new_net_2102),
		.c(new_net_2103)
	);

	spl2 _1396__v_fanout (
		.a(_1396_),
		.b(new_net_3109),
		.c(new_net_3110)
	);

	spl2 _0002__v_fanout (
		.a(_0002_),
		.b(new_net_1006),
		.c(new_net_1007)
	);

	spl2 _1310__v_fanout (
		.a(_1310_),
		.b(new_net_1346),
		.c(new_net_1347)
	);

	spl2 _0187__v_fanout (
		.a(_0187_),
		.b(new_net_88),
		.c(new_net_89)
	);

	spl2 _0492__v_fanout (
		.a(_0492_),
		.b(new_net_1519),
		.c(new_net_1520)
	);

	spl2 _1785__v_fanout (
		.a(_1785_),
		.b(new_net_275),
		.c(new_net_276)
	);

	spl2 _1721__v_fanout (
		.a(_1721_),
		.b(new_net_1396),
		.c(new_net_1397)
	);

	spl2 _1233__v_fanout (
		.a(_1233_),
		.b(new_net_1652),
		.c(new_net_1653)
	);

	spl2 _1156__v_fanout (
		.a(_1156_),
		.b(new_net_1872),
		.c(new_net_1873)
	);

	spl2 _1096__v_fanout (
		.a(_1096_),
		.b(new_net_1495),
		.c(new_net_1496)
	);

	spl2 _1492__v_fanout (
		.a(_1492_),
		.b(new_net_305),
		.c(new_net_306)
	);

	spl2 _1395__v_fanout (
		.a(_1395_),
		.b(new_net_3075),
		.c(new_net_3076)
	);

	spl2 _1044__v_fanout (
		.a(_1044_),
		.b(new_net_1902),
		.c(new_net_1903)
	);

	spl2 _0882__v_fanout (
		.a(_0882_),
		.b(new_net_2669),
		.c(new_net_2670)
	);

	spl2 _1602__v_fanout (
		.a(_1602_),
		.b(new_net_2923),
		.c(new_net_2924)
	);

	bfr new_net_5567_bfr_before (
		.din(new_net_5567),
		.dout(new_net_951)
	);

	bfr new_net_5568_bfr_before (
		.din(new_net_5568),
		.dout(new_net_5567)
	);

	bfr new_net_5569_bfr_before (
		.din(new_net_5569),
		.dout(new_net_5568)
	);

	bfr new_net_5570_bfr_before (
		.din(new_net_5570),
		.dout(new_net_5569)
	);

	spl2 _0239__v_fanout (
		.a(_0239_),
		.b(new_net_950),
		.c(new_net_5570)
	);

	bfr new_net_5571_bfr_after (
		.din(_0119_),
		.dout(new_net_5571)
	);

	bfr new_net_5572_bfr_after (
		.din(new_net_5571),
		.dout(new_net_5572)
	);

	bfr new_net_5573_bfr_after (
		.din(new_net_5572),
		.dout(new_net_5573)
	);

	bfr new_net_5574_bfr_after (
		.din(new_net_5573),
		.dout(new_net_5574)
	);

	spl2 _0119__v_fanout (
		.a(new_net_5574),
		.b(new_net_2390),
		.c(new_net_2391)
	);

	bfr new_net_5575_bfr_before (
		.din(new_net_5575),
		.dout(new_net_1341)
	);

	bfr new_net_5576_bfr_before (
		.din(new_net_5576),
		.dout(new_net_5575)
	);

	bfr new_net_5577_bfr_before (
		.din(new_net_5577),
		.dout(new_net_5576)
	);

	bfr new_net_5578_bfr_before (
		.din(new_net_5578),
		.dout(new_net_5577)
	);

	spl2 _0470__v_fanout (
		.a(_0470_),
		.b(new_net_1340),
		.c(new_net_5578)
	);

	bfr new_net_5579_bfr_before (
		.din(new_net_5579),
		.dout(new_net_1787)
	);

	bfr new_net_5580_bfr_before (
		.din(new_net_5580),
		.dout(new_net_5579)
	);

	bfr new_net_5581_bfr_before (
		.din(new_net_5581),
		.dout(new_net_5580)
	);

	bfr new_net_5582_bfr_before (
		.din(new_net_5582),
		.dout(new_net_5581)
	);

	spl2 _1154__v_fanout (
		.a(_1154_),
		.b(new_net_1786),
		.c(new_net_5582)
	);

	bfr new_net_5583_bfr_before (
		.din(new_net_5583),
		.dout(new_net_2483)
	);

	bfr new_net_5584_bfr_before (
		.din(new_net_5584),
		.dout(new_net_5583)
	);

	bfr new_net_5585_bfr_before (
		.din(new_net_5585),
		.dout(new_net_5584)
	);

	bfr new_net_5586_bfr_before (
		.din(new_net_5586),
		.dout(new_net_5585)
	);

	spl2 _1718__v_fanout (
		.a(_1718_),
		.b(new_net_2482),
		.c(new_net_5586)
	);

	bfr new_net_5587_bfr_before (
		.din(new_net_5587),
		.dout(new_net_1568)
	);

	bfr new_net_5588_bfr_before (
		.din(new_net_5588),
		.dout(new_net_5587)
	);

	bfr new_net_5589_bfr_before (
		.din(new_net_5589),
		.dout(new_net_5588)
	);

	bfr new_net_5590_bfr_before (
		.din(new_net_5590),
		.dout(new_net_5589)
	);

	spl2 _1231__v_fanout (
		.a(_1231_),
		.b(new_net_1567),
		.c(new_net_5590)
	);

	bfr new_net_5591_bfr_before (
		.din(new_net_5591),
		.dout(new_net_483)
	);

	bfr new_net_5592_bfr_before (
		.din(new_net_5592),
		.dout(new_net_5591)
	);

	bfr new_net_5593_bfr_before (
		.din(new_net_5593),
		.dout(new_net_5592)
	);

	bfr new_net_5594_bfr_before (
		.din(new_net_5594),
		.dout(new_net_5593)
	);

	spl2 _1600__v_fanout (
		.a(_1600_),
		.b(new_net_482),
		.c(new_net_5594)
	);

	bfr new_net_5595_bfr_before (
		.din(new_net_5595),
		.dout(new_net_1071)
	);

	bfr new_net_5596_bfr_before (
		.din(new_net_5596),
		.dout(new_net_5595)
	);

	bfr new_net_5597_bfr_before (
		.din(new_net_5597),
		.dout(new_net_5596)
	);

	bfr new_net_5598_bfr_before (
		.din(new_net_5598),
		.dout(new_net_5597)
	);

	spl2 _1094__v_fanout (
		.a(_1094_),
		.b(new_net_1070),
		.c(new_net_5598)
	);

	bfr new_net_5599_bfr_before (
		.din(new_net_5599),
		.dout(new_net_1591)
	);

	bfr new_net_5600_bfr_before (
		.din(new_net_5600),
		.dout(new_net_5599)
	);

	bfr new_net_5601_bfr_before (
		.din(new_net_5601),
		.dout(new_net_5600)
	);

	bfr new_net_5602_bfr_before (
		.din(new_net_5602),
		.dout(new_net_5601)
	);

	spl2 _1042__v_fanout (
		.a(_1042_),
		.b(new_net_1590),
		.c(new_net_5602)
	);

	bfr new_net_5603_bfr_before (
		.din(new_net_5603),
		.dout(new_net_1841)
	);

	bfr new_net_5604_bfr_before (
		.din(new_net_5604),
		.dout(new_net_5603)
	);

	bfr new_net_5605_bfr_before (
		.din(new_net_5605),
		.dout(new_net_5604)
	);

	bfr new_net_5606_bfr_before (
		.din(new_net_5606),
		.dout(new_net_5605)
	);

	spl2 _0861__v_fanout (
		.a(_0861_),
		.b(new_net_1840),
		.c(new_net_5606)
	);

	spl2 _0001__v_fanout (
		.a(_0001_),
		.b(new_net_956),
		.c(new_net_957)
	);

	bfr new_net_5607_bfr_before (
		.din(new_net_5607),
		.dout(new_net_2964)
	);

	bfr new_net_5608_bfr_before (
		.din(new_net_5608),
		.dout(new_net_5607)
	);

	bfr new_net_5609_bfr_before (
		.din(new_net_5609),
		.dout(new_net_5608)
	);

	bfr new_net_5610_bfr_before (
		.din(new_net_5610),
		.dout(new_net_5609)
	);

	spl2 _1393__v_fanout (
		.a(_1393_),
		.b(new_net_2963),
		.c(new_net_5610)
	);

	spl2 _0238__v_fanout (
		.a(_0238_),
		.b(new_net_777),
		.c(new_net_778)
	);

	bfr new_net_5611_bfr_before (
		.din(new_net_5611),
		.dout(new_net_447)
	);

	bfr new_net_5612_bfr_before (
		.din(new_net_5612),
		.dout(new_net_5611)
	);

	bfr new_net_5613_bfr_before (
		.din(new_net_5613),
		.dout(new_net_5612)
	);

	bfr new_net_5614_bfr_before (
		.din(new_net_5614),
		.dout(new_net_5613)
	);

	spl2 _1763__v_fanout (
		.a(_1763_),
		.b(new_net_446),
		.c(new_net_5614)
	);

	bfr new_net_5615_bfr_before (
		.din(new_net_5615),
		.dout(new_net_1274)
	);

	bfr new_net_5616_bfr_before (
		.din(new_net_5616),
		.dout(new_net_5615)
	);

	bfr new_net_5617_bfr_before (
		.din(new_net_5617),
		.dout(new_net_5616)
	);

	bfr new_net_5618_bfr_before (
		.din(new_net_5618),
		.dout(new_net_5617)
	);

	spl2 _1308__v_fanout (
		.a(_1308_),
		.b(new_net_1273),
		.c(new_net_5618)
	);

	bfr new_net_5619_bfr_before (
		.din(new_net_5619),
		.dout(new_net_461)
	);

	bfr new_net_5620_bfr_before (
		.din(new_net_5620),
		.dout(new_net_5619)
	);

	bfr new_net_5621_bfr_before (
		.din(new_net_5621),
		.dout(new_net_5620)
	);

	bfr new_net_5622_bfr_before (
		.din(new_net_5622),
		.dout(new_net_5621)
	);

	spl2 _0165__v_fanout (
		.a(_0165_),
		.b(new_net_460),
		.c(new_net_5622)
	);

	bfr new_net_5623_bfr_before (
		.din(new_net_5623),
		.dout(new_net_1199)
	);

	bfr new_net_5624_bfr_before (
		.din(new_net_5624),
		.dout(new_net_5623)
	);

	bfr new_net_5625_bfr_before (
		.din(new_net_5625),
		.dout(new_net_5624)
	);

	bfr new_net_5626_bfr_before (
		.din(new_net_5626),
		.dout(new_net_5625)
	);

	spl2 _1489__v_fanout (
		.a(_1489_),
		.b(new_net_1198),
		.c(new_net_5626)
	);

	spl2 _1093__v_fanout (
		.a(_1093_),
		.b(new_net_932),
		.c(new_net_933)
	);

	spl2 _1218__v_fanout (
		.a(_1218_),
		.b(new_net_1052),
		.c(new_net_1053)
	);

	spl2 _1230__v_fanout (
		.a(_1230_),
		.b(new_net_1527),
		.c(new_net_1528)
	);

	spl2 _1488__v_fanout (
		.a(_1488_),
		.b(new_net_176),
		.c(new_net_177)
	);

	spl2 _1307__v_fanout (
		.a(_1307_),
		.b(new_net_2280),
		.c(new_net_2281)
	);

	spl2 _1621__v_fanout (
		.a(_1621_),
		.b(new_net_1886),
		.c(new_net_1887)
	);

	spl2 _1475__v_fanout (
		.a(_1475_),
		.b(new_net_2631),
		.c(new_net_2632)
	);

	spl2 _1041__v_fanout (
		.a(_1041_),
		.b(new_net_771),
		.c(new_net_772)
	);

	spl2 _0720__v_fanout (
		.a(_0720_),
		.b(new_net_2933),
		.c(new_net_2934)
	);

	spl2 _1752__v_fanout (
		.a(_1752_),
		.b(new_net_1586),
		.c(new_net_1587)
	);

	spl2 _1081__v_fanout (
		.a(_1081_),
		.b(new_net_2230),
		.c(new_net_2231)
	);

	bfr new_net_5627_bfr_before (
		.din(new_net_5627),
		.dout(new_net_2451)
	);

	bfr new_net_5628_bfr_before (
		.din(new_net_5628),
		.dout(new_net_5627)
	);

	bfr new_net_5629_bfr_before (
		.din(new_net_5629),
		.dout(new_net_5628)
	);

	bfr new_net_5630_bfr_before (
		.din(new_net_5630),
		.dout(new_net_5629)
	);

	spl2 _1836__v_fanout (
		.a(_1836_),
		.b(new_net_2450),
		.c(new_net_5630)
	);

	spl2 _0154__v_fanout (
		.a(_0154_),
		.b(new_net_1600),
		.c(new_net_1601)
	);

	spl2 _1380__v_fanout (
		.a(_1380_),
		.b(new_net_188),
		.c(new_net_189)
	);

	spl2 _0459__v_fanout (
		.a(_0459_),
		.b(new_net_970),
		.c(new_net_971)
	);

	spl2 _1141__v_fanout (
		.a(_1141_),
		.b(new_net_1318),
		.c(new_net_1319)
	);

	spl2 _0117__v_fanout (
		.a(_0117_),
		.b(new_net_753),
		.c(new_net_754)
	);

	spl2 _0022__v_fanout (
		.a(_0022_),
		.b(new_net_3165),
		.c(new_net_3166)
	);

	spl2 _1598__v_fanout (
		.a(_1598_),
		.b(new_net_114),
		.c(new_net_115)
	);

	spl2 _1585__v_fanout (
		.a(_1585_),
		.b(new_net_886),
		.c(new_net_887)
	);

	spl2 _0328__v_fanout (
		.a(_0328_),
		.b(new_net_2134),
		.c(new_net_2135)
	);

	spl2 _1153__v_fanout (
		.a(_1153_),
		.b(new_net_2897),
		.c(new_net_2898)
	);

	spl2 _1705__v_fanout (
		.a(_1705_),
		.b(new_net_1984),
		.c(new_net_1985)
	);

	spl2 _1029__v_fanout (
		.a(_1029_),
		.b(new_net_2276),
		.c(new_net_2277)
	);

	spl2 _1392__v_fanout (
		.a(_1392_),
		.b(new_net_2901),
		.c(new_net_2902)
	);

	spl2 _0850__v_fanout (
		.a(_0850_),
		.b(new_net_3115),
		.c(new_net_3116)
	);

	spl2 _1295__v_fanout (
		.a(_1295_),
		.b(new_net_854),
		.c(new_net_855)
	);

	spl2 _0828__v_fanout (
		.a(_0828_),
		.b(new_net_1038),
		.c(new_net_1039)
	);

	spl2 _1829__v_fanout (
		.a(_1829_),
		.b(new_net_1918),
		.c(new_net_1919)
	);

	spl2 _1486__v_fanout (
		.a(_1486_),
		.b(new_net_675),
		.c(new_net_676)
	);

	bfr new_net_5631_bfr_after (
		.din(_1717_),
		.dout(new_net_5631)
	);

	bfr new_net_5632_bfr_after (
		.din(new_net_5631),
		.dout(new_net_5632)
	);

	spl2 _1717__v_fanout (
		.a(new_net_5632),
		.b(new_net_687),
		.c(new_net_688)
	);

	spl2 _1091__v_fanout (
		.a(_1091_),
		.b(new_net_2649),
		.c(new_net_2650)
	);

	spl2 _0132__v_fanout (
		.a(_0132_),
		.b(new_net_2905),
		.c(new_net_2906)
	);

	spl2 _1228__v_fanout (
		.a(_1228_),
		.b(new_net_1230),
		.c(new_net_1231)
	);

	spl2 _1610__v_fanout (
		.a(_1610_),
		.b(new_net_3123),
		.c(new_net_3124)
	);

	spl2 _1039__v_fanout (
		.a(_1039_),
		.b(new_net_655),
		.c(new_net_656)
	);

	spl2 _1151__v_fanout (
		.a(_1151_),
		.b(new_net_2480),
		.c(new_net_2481)
	);

	spl2 _1730__v_fanout (
		.a(_1730_),
		.b(new_net_3213),
		.c(new_net_3214)
	);

	spl2 _0116__v_fanout (
		.a(_0116_),
		.b(new_net_544),
		.c(new_net_545)
	);

	spl2 _0437__v_fanout (
		.a(_0437_),
		.b(new_net_120),
		.c(new_net_121)
	);

	spl2 _1596__v_fanout (
		.a(_1596_),
		.b(new_net_2953),
		.c(new_net_2954)
	);

	spl2 _1305__v_fanout (
		.a(_1305_),
		.b(new_net_1898),
		.c(new_net_1899)
	);

	spl2 _1390__v_fanout (
		.a(_1390_),
		.b(new_net_2038),
		.c(new_net_2039)
	);

	spl2 _1227__v_fanout (
		.a(_1227_),
		.b(new_net_1374),
		.c(new_net_1375)
	);

	spl2 _1389__v_fanout (
		.a(_1389_),
		.b(new_net_2775),
		.c(new_net_2776)
	);

	spl2 _1719__v_fanout (
		.a(_1719_),
		.b(new_net_2537),
		.c(new_net_2538)
	);

	spl2 _1038__v_fanout (
		.a(_1038_),
		.b(new_net_626),
		.c(new_net_627)
	);

	spl2 _0818__v_fanout (
		.a(_0818_),
		.b(new_net_1780),
		.c(new_net_1781)
	);

	spl2 _1304__v_fanout (
		.a(_1304_),
		.b(new_net_1718),
		.c(new_net_1719)
	);

	spl2 _0121__v_fanout (
		.a(_0121_),
		.b(new_net_1499),
		.c(new_net_1500)
	);

	spl2 _1599__v_fanout (
		.a(_1599_),
		.b(new_net_2773),
		.c(new_net_2774)
	);

	spl2 _1150__v_fanout (
		.a(_1150_),
		.b(new_net_2282),
		.c(new_net_2283)
	);

	spl2 _1090__v_fanout (
		.a(_1090_),
		.b(new_net_329),
		.c(new_net_330)
	);

	spl2 _1595__v_fanout (
		.a(_1595_),
		.b(new_net_2744),
		.c(new_net_2745)
	);

	bfr new_net_5633_bfr_before (
		.din(new_net_5633),
		.dout(new_net_2187)
	);

	bfr new_net_5634_bfr_before (
		.din(new_net_5634),
		.dout(new_net_5633)
	);

	bfr new_net_5635_bfr_before (
		.din(new_net_5635),
		.dout(new_net_5634)
	);

	bfr new_net_5636_bfr_before (
		.din(new_net_5636),
		.dout(new_net_5635)
	);

	spl2 _0114__v_fanout (
		.a(_0114_),
		.b(new_net_2186),
		.c(new_net_5636)
	);

	spl2 _0427__v_fanout (
		.a(_0427_),
		.b(new_net_1310),
		.c(new_net_1311)
	);

	spl2 _1485__v_fanout (
		.a(_1485_),
		.b(new_net_484),
		.c(new_net_485)
	);

	spl2 _1715__v_fanout (
		.a(_1715_),
		.b(new_net_297),
		.c(new_net_298)
	);

	bfr new_net_5637_bfr_before (
		.din(new_net_5637),
		.dout(new_net_3221)
	);

	bfr new_net_5638_bfr_before (
		.din(new_net_5638),
		.dout(new_net_5637)
	);

	bfr new_net_5639_bfr_before (
		.din(new_net_5639),
		.dout(new_net_5638)
	);

	bfr new_net_5640_bfr_before (
		.din(new_net_5640),
		.dout(new_net_5639)
	);

	spl2 _0405__v_fanout (
		.a(_0405_),
		.b(new_net_3220),
		.c(new_net_5640)
	);

	bfr new_net_5641_bfr_before (
		.din(new_net_5641),
		.dout(new_net_3194)
	);

	bfr new_net_5642_bfr_before (
		.din(new_net_5642),
		.dout(new_net_5641)
	);

	bfr new_net_5643_bfr_before (
		.din(new_net_5643),
		.dout(new_net_5642)
	);

	bfr new_net_5644_bfr_before (
		.din(new_net_5644),
		.dout(new_net_5643)
	);

	spl2 _1566__v_fanout (
		.a(_1566_),
		.b(new_net_3193),
		.c(new_net_5644)
	);

	bfr new_net_5645_bfr_before (
		.din(new_net_5645),
		.dout(new_net_720)
	);

	bfr new_net_5646_bfr_before (
		.din(new_net_5646),
		.dout(new_net_5645)
	);

	bfr new_net_5647_bfr_before (
		.din(new_net_5647),
		.dout(new_net_5646)
	);

	bfr new_net_5648_bfr_before (
		.din(new_net_5648),
		.dout(new_net_5647)
	);

	spl2 _1225__v_fanout (
		.a(_1225_),
		.b(new_net_719),
		.c(new_net_5648)
	);

	bfr new_net_5649_bfr_before (
		.din(new_net_5649),
		.dout(new_net_1351)
	);

	bfr new_net_5650_bfr_before (
		.din(new_net_5650),
		.dout(new_net_5649)
	);

	bfr new_net_5651_bfr_before (
		.din(new_net_5651),
		.dout(new_net_5650)
	);

	bfr new_net_5652_bfr_before (
		.din(new_net_5652),
		.dout(new_net_5651)
	);

	spl2 _1302__v_fanout (
		.a(_1302_),
		.b(new_net_1350),
		.c(new_net_5652)
	);

	bfr new_net_5653_bfr_before (
		.din(new_net_5653),
		.dout(new_net_2477)
	);

	bfr new_net_5654_bfr_before (
		.din(new_net_5654),
		.dout(new_net_5653)
	);

	bfr new_net_5655_bfr_before (
		.din(new_net_5655),
		.dout(new_net_5654)
	);

	bfr new_net_5656_bfr_before (
		.din(new_net_5656),
		.dout(new_net_5655)
	);

	spl2 _0796__v_fanout (
		.a(_0796_),
		.b(new_net_2476),
		.c(new_net_5656)
	);

	bfr new_net_5657_bfr_after (
		.din(_1835_),
		.dout(new_net_5657)
	);

	bfr new_net_5658_bfr_after (
		.din(new_net_5657),
		.dout(new_net_5658)
	);

	bfr new_net_5659_bfr_after (
		.din(new_net_5658),
		.dout(new_net_5659)
	);

	bfr new_net_5660_bfr_after (
		.din(new_net_5659),
		.dout(new_net_5660)
	);

	spl2 _1835__v_fanout (
		.a(new_net_5660),
		.b(new_net_2252),
		.c(new_net_2253)
	);

	spl2 _1714__v_fanout (
		.a(_1714_),
		.b(new_net_2361),
		.c(new_net_2362)
	);

	bfr new_net_5661_bfr_before (
		.din(new_net_5661),
		.dout(new_net_445)
	);

	bfr new_net_5662_bfr_before (
		.din(new_net_5662),
		.dout(new_net_5661)
	);

	bfr new_net_5663_bfr_before (
		.din(new_net_5663),
		.dout(new_net_5662)
	);

	bfr new_net_5664_bfr_before (
		.din(new_net_5664),
		.dout(new_net_5663)
	);

	spl2 _1036__v_fanout (
		.a(_1036_),
		.b(new_net_444),
		.c(new_net_5664)
	);

	spl2 _0113__v_fanout (
		.a(_0113_),
		.b(new_net_2150),
		.c(new_net_2151)
	);

	bfr new_net_5665_bfr_before (
		.din(new_net_5665),
		.dout(new_net_2336)
	);

	bfr new_net_5666_bfr_before (
		.din(new_net_5666),
		.dout(new_net_5665)
	);

	bfr new_net_5667_bfr_before (
		.din(new_net_5667),
		.dout(new_net_5666)
	);

	bfr new_net_5668_bfr_before (
		.din(new_net_5668),
		.dout(new_net_5667)
	);

	spl2 _1593__v_fanout (
		.a(_1593_),
		.b(new_net_2335),
		.c(new_net_5668)
	);

	bfr new_net_5669_bfr_before (
		.din(new_net_5669),
		.dout(new_net_525)
	);

	bfr new_net_5670_bfr_before (
		.din(new_net_5670),
		.dout(new_net_5669)
	);

	bfr new_net_5671_bfr_before (
		.din(new_net_5671),
		.dout(new_net_5670)
	);

	bfr new_net_5672_bfr_before (
		.din(new_net_5672),
		.dout(new_net_5671)
	);

	spl2 _0099__v_fanout (
		.a(_0099_),
		.b(new_net_524),
		.c(new_net_5672)
	);

	bfr new_net_5673_bfr_before (
		.din(new_net_5673),
		.dout(new_net_953)
	);

	bfr new_net_5674_bfr_before (
		.din(new_net_5674),
		.dout(new_net_5673)
	);

	bfr new_net_5675_bfr_before (
		.din(new_net_5675),
		.dout(new_net_5674)
	);

	bfr new_net_5676_bfr_before (
		.din(new_net_5676),
		.dout(new_net_5675)
	);

	spl2 _1483__v_fanout (
		.a(_1483_),
		.b(new_net_952),
		.c(new_net_5676)
	);

	bfr new_net_5677_bfr_before (
		.din(new_net_5677),
		.dout(new_net_3275)
	);

	bfr new_net_5678_bfr_before (
		.din(new_net_5678),
		.dout(new_net_5677)
	);

	bfr new_net_5679_bfr_before (
		.din(new_net_5679),
		.dout(new_net_5678)
	);

	bfr new_net_5680_bfr_before (
		.din(new_net_5680),
		.dout(new_net_5679)
	);

	spl2 _1088__v_fanout (
		.a(_1088_),
		.b(new_net_3274),
		.c(new_net_5680)
	);

	bfr new_net_5681_bfr_before (
		.din(new_net_5681),
		.dout(new_net_1524)
	);

	bfr new_net_5682_bfr_before (
		.din(new_net_5682),
		.dout(new_net_5681)
	);

	bfr new_net_5683_bfr_before (
		.din(new_net_5683),
		.dout(new_net_5682)
	);

	bfr new_net_5684_bfr_before (
		.din(new_net_5684),
		.dout(new_net_5683)
	);

	spl2 _1387__v_fanout (
		.a(_1387_),
		.b(new_net_1523),
		.c(new_net_5684)
	);

	bfr new_net_5685_bfr_before (
		.din(new_net_5685),
		.dout(new_net_1901)
	);

	bfr new_net_5686_bfr_before (
		.din(new_net_5686),
		.dout(new_net_5685)
	);

	bfr new_net_5687_bfr_before (
		.din(new_net_5687),
		.dout(new_net_5686)
	);

	bfr new_net_5688_bfr_before (
		.din(new_net_5688),
		.dout(new_net_5687)
	);

	spl2 _1148__v_fanout (
		.a(_1148_),
		.b(new_net_1900),
		.c(new_net_5688)
	);

	bfr new_net_5689_bfr_before (
		.din(new_net_5689),
		.dout(new_net_1707)
	);

	bfr new_net_5690_bfr_before (
		.din(new_net_5690),
		.dout(new_net_5689)
	);

	bfr new_net_5691_bfr_before (
		.din(new_net_5691),
		.dout(new_net_5690)
	);

	bfr new_net_5692_bfr_before (
		.din(new_net_5692),
		.dout(new_net_5691)
	);

	spl2 _1697__v_fanout (
		.a(_1697_),
		.b(new_net_1706),
		.c(new_net_5692)
	);

	spl2 new_net_3442_v_fanout (
		.a(new_net_3442),
		.b(new_net_256),
		.c(new_net_255)
	);

	spl2 _0088__v_fanout (
		.a(_0088_),
		.b(new_net_2819),
		.c(new_net_2820)
	);

	spl2 new_net_3446_v_fanout (
		.a(new_net_3446),
		.b(new_net_1401),
		.c(new_net_1402)
	);

	spl2 _1087__v_fanout (
		.a(_1087_),
		.b(new_net_2452),
		.c(new_net_2453)
	);

	spl2 _1035__v_fanout (
		.a(_1035_),
		.b(new_net_506),
		.c(new_net_507)
	);

	spl2 _1386__v_fanout (
		.a(_1386_),
		.b(new_net_2679),
		.c(new_net_2680)
	);

	spl2 _1147__v_fanout (
		.a(_1147_),
		.b(new_net_3205),
		.c(new_net_3206)
	);

	spl2 _1224__v_fanout (
		.a(_1224_),
		.b(new_net_510),
		.c(new_net_511)
	);

	spl2 _1535__v_fanout (
		.a(_1535_),
		.b(new_net_1908),
		.c(new_net_1909)
	);

	spl2 _1686__v_fanout (
		.a(_1686_),
		.b(new_net_1269),
		.c(new_net_1270)
	);

	bfr new_net_5693_bfr_before (
		.din(new_net_5693),
		.dout(new_net_3204)
	);

	bfr new_net_5694_bfr_before (
		.din(new_net_5694),
		.dout(new_net_5693)
	);

	bfr new_net_5695_bfr_before (
		.din(new_net_5695),
		.dout(new_net_5694)
	);

	bfr new_net_5696_bfr_before (
		.din(new_net_5696),
		.dout(new_net_5695)
	);

	spl2 _1713__v_fanout (
		.a(_1713_),
		.b(new_net_3203),
		.c(new_net_5696)
	);

	spl2 new_net_3444_v_fanout (
		.a(new_net_3444),
		.b(new_net_1578),
		.c(new_net_1579)
	);

	spl2 _1301__v_fanout (
		.a(_1301_),
		.b(new_net_1164),
		.c(new_net_1165)
	);

	spl2 new_net_3448_v_fanout (
		.a(new_net_3448),
		.b(new_net_808),
		.c(new_net_809)
	);

	spl2 new_net_3445_v_fanout (
		.a(new_net_3445),
		.b(new_net_1234),
		.c(new_net_1233)
	);

	spl2 new_net_3452_v_fanout (
		.a(new_net_3452),
		.b(new_net_3219),
		.c(new_net_3218)
	);

	spl2 new_net_3453_v_fanout (
		.a(new_net_3453),
		.b(new_net_5),
		.c(new_net_4)
	);

	spl2 new_net_3441_v_fanout (
		.a(new_net_3441),
		.b(new_net_631),
		.c(new_net_632)
	);

	spl2 _0785__v_fanout (
		.a(_0785_),
		.b(new_net_602),
		.c(new_net_603)
	);

	spl2 _0394__v_fanout (
		.a(_0394_),
		.b(new_net_1060),
		.c(new_net_1061)
	);

	spl2 new_net_3443_v_fanout (
		.a(new_net_3443),
		.b(new_net_348),
		.c(new_net_349)
	);

	spl2 new_net_3449_v_fanout (
		.a(new_net_3449),
		.b(new_net_2892),
		.c(new_net_2891)
	);

	spl2 _1482__v_fanout (
		.a(_1482_),
		.b(new_net_781),
		.c(new_net_782)
	);

	spl2 new_net_3447_v_fanout (
		.a(new_net_3447),
		.b(new_net_1296),
		.c(new_net_1297)
	);

	spl2 _1833__v_fanout (
		.a(_1833_),
		.b(new_net_1860),
		.c(new_net_1861)
	);

	spl2 new_net_3451_v_fanout (
		.a(new_net_3451),
		.b(new_net_2754),
		.c(new_net_2756)
	);

	spl2 _1592__v_fanout (
		.a(_1592_),
		.b(new_net_2140),
		.c(new_net_2141)
	);

	spl2 new_net_3450_v_fanout (
		.a(new_net_3450),
		.b(new_net_2364),
		.c(new_net_2365)
	);

	bfr new_net_5697_bfr_before (
		.din(new_net_5697),
		.dout(new_net_3442)
	);

	spl2 _1491__v_fanout (
		.a(_1491_),
		.b(new_net_254),
		.c(new_net_5697)
	);

	bfr new_net_5698_bfr_before (
		.din(new_net_5698),
		.dout(new_net_3449)
	);

	spl2 _1032__v_fanout (
		.a(_1032_),
		.b(new_net_2890),
		.c(new_net_5698)
	);

	bfr new_net_5699_bfr_before (
		.din(new_net_5699),
		.dout(new_net_3451)
	);

	spl2 _1556__v_fanout (
		.a(_1556_),
		.b(new_net_5699),
		.c(new_net_2755)
	);

	bfr new_net_5700_bfr_before (
		.din(new_net_5700),
		.dout(new_net_3453)
	);

	spl2 _1478__v_fanout (
		.a(_1478_),
		.b(new_net_3),
		.c(new_net_5700)
	);

	bfr new_net_5701_bfr_before (
		.din(new_net_5701),
		.dout(new_net_3448)
	);

	spl2 _1383__v_fanout (
		.a(_1383_),
		.b(new_net_807),
		.c(new_net_5701)
	);

	bfr new_net_5702_bfr_before (
		.din(new_net_5702),
		.dout(new_net_3447)
	);

	spl2 _0753__v_fanout (
		.a(_0753_),
		.b(new_net_1295),
		.c(new_net_5702)
	);

	bfr new_net_5703_bfr_before (
		.din(new_net_5703),
		.dout(new_net_3446)
	);

	spl2 _1144__v_fanout (
		.a(_1144_),
		.b(new_net_1400),
		.c(new_net_5703)
	);

	bfr new_net_5704_bfr_before (
		.din(new_net_5704),
		.dout(new_net_3443)
	);

	spl2 _1654__v_fanout (
		.a(_1654_),
		.b(new_net_347),
		.c(new_net_5704)
	);

	bfr new_net_5705_bfr_before (
		.din(new_net_5705),
		.dout(new_net_3441)
	);

	spl2 _1298__v_fanout (
		.a(_1298_),
		.b(new_net_630),
		.c(new_net_5705)
	);

	bfr new_net_5706_bfr_before (
		.din(new_net_5706),
		.dout(new_net_3445)
	);

	spl2 _0361__v_fanout (
		.a(_0361_),
		.b(new_net_1232),
		.c(new_net_5706)
	);

	bfr new_net_5707_bfr_before (
		.din(new_net_5707),
		.dout(new_net_3450)
	);

	spl2 _1084__v_fanout (
		.a(_1084_),
		.b(new_net_2363),
		.c(new_net_5707)
	);

	bfr new_net_5708_bfr_before (
		.din(new_net_5708),
		.dout(new_net_3444)
	);

	spl2 _0055__v_fanout (
		.a(_0055_),
		.b(new_net_1577),
		.c(new_net_5708)
	);

	bfr new_net_5709_bfr_before (
		.din(new_net_5709),
		.dout(new_net_3452)
	);

	spl2 _1221__v_fanout (
		.a(_1221_),
		.b(new_net_3217),
		.c(new_net_5709)
	);

	bfr new_net_5710_bfr_before (
		.din(new_net_5710),
		.dout(new_net_2387)
	);

	spl2 _1589__v_fanout (
		.a(_1589_),
		.b(new_net_2386),
		.c(new_net_5710)
	);

	spl2 _1831__v_fanout (
		.a(_1831_),
		.b(new_net_1541),
		.c(new_net_1542)
	);

	bfr new_net_5711_bfr_after (
		.din(_1474_),
		.dout(new_net_5711)
	);

	bfr new_net_5712_bfr_after (
		.din(new_net_5711),
		.dout(new_net_5712)
	);

	bfr new_net_5713_bfr_after (
		.din(new_net_5712),
		.dout(new_net_5713)
	);

	bfr new_net_5714_bfr_after (
		.din(new_net_5713),
		.dout(new_net_5714)
	);

	bfr new_net_5715_bfr_after (
		.din(new_net_5714),
		.dout(new_net_5715)
	);

	bfr new_net_5716_bfr_after (
		.din(new_net_5715),
		.dout(new_net_5716)
	);

	bfr new_net_5717_bfr_after (
		.din(new_net_5716),
		.dout(new_net_5717)
	);

	bfr new_net_5718_bfr_after (
		.din(new_net_5717),
		.dout(new_net_5718)
	);

	bfr new_net_5719_bfr_after (
		.din(new_net_5718),
		.dout(new_net_5719)
	);

	bfr new_net_5720_bfr_after (
		.din(new_net_5719),
		.dout(new_net_5720)
	);

	bfr new_net_5721_bfr_after (
		.din(new_net_5720),
		.dout(new_net_5721)
	);

	bfr new_net_5722_bfr_after (
		.din(new_net_5721),
		.dout(new_net_5722)
	);

	bfr new_net_5723_bfr_after (
		.din(new_net_5722),
		.dout(new_net_5723)
	);

	bfr new_net_5724_bfr_after (
		.din(new_net_5723),
		.dout(new_net_5724)
	);

	bfr new_net_5725_bfr_after (
		.din(new_net_5724),
		.dout(new_net_5725)
	);

	bfr new_net_5726_bfr_after (
		.din(new_net_5725),
		.dout(new_net_5726)
	);

	spl2 _1474__v_fanout (
		.a(new_net_5726),
		.b(new_net_1182),
		.c(new_net_1183)
	);

	bfr new_net_5727_bfr_after (
		.din(_0703_),
		.dout(new_net_5727)
	);

	bfr new_net_5728_bfr_after (
		.din(new_net_5727),
		.dout(new_net_5728)
	);

	bfr new_net_5729_bfr_after (
		.din(new_net_5728),
		.dout(new_net_5729)
	);

	bfr new_net_5730_bfr_after (
		.din(new_net_5729),
		.dout(new_net_5730)
	);

	bfr new_net_5731_bfr_after (
		.din(new_net_5730),
		.dout(new_net_5731)
	);

	bfr new_net_5732_bfr_after (
		.din(new_net_5731),
		.dout(new_net_5732)
	);

	bfr new_net_5733_bfr_after (
		.din(new_net_5732),
		.dout(new_net_5733)
	);

	bfr new_net_5734_bfr_after (
		.din(new_net_5733),
		.dout(new_net_5734)
	);

	bfr new_net_5735_bfr_after (
		.din(new_net_5734),
		.dout(new_net_5735)
	);

	bfr new_net_5736_bfr_after (
		.din(new_net_5735),
		.dout(new_net_5736)
	);

	bfr new_net_5737_bfr_after (
		.din(new_net_5736),
		.dout(new_net_5737)
	);

	bfr new_net_5738_bfr_after (
		.din(new_net_5737),
		.dout(new_net_5738)
	);

	bfr new_net_5739_bfr_after (
		.din(new_net_5738),
		.dout(new_net_5739)
	);

	bfr new_net_5740_bfr_after (
		.din(new_net_5739),
		.dout(new_net_5740)
	);

	bfr new_net_5741_bfr_after (
		.din(new_net_5740),
		.dout(new_net_5741)
	);

	bfr new_net_5742_bfr_after (
		.din(new_net_5741),
		.dout(new_net_5742)
	);

	bfr new_net_5743_bfr_after (
		.din(new_net_5742),
		.dout(new_net_5743)
	);

	bfr new_net_5744_bfr_after (
		.din(new_net_5743),
		.dout(new_net_5744)
	);

	bfr new_net_5745_bfr_after (
		.din(new_net_5744),
		.dout(new_net_5745)
	);

	bfr new_net_5746_bfr_after (
		.din(new_net_5745),
		.dout(new_net_5746)
	);

	bfr new_net_5747_bfr_after (
		.din(new_net_5746),
		.dout(new_net_5747)
	);

	bfr new_net_5748_bfr_after (
		.din(new_net_5747),
		.dout(new_net_5748)
	);

	bfr new_net_5749_bfr_after (
		.din(new_net_5748),
		.dout(new_net_5749)
	);

	bfr new_net_5750_bfr_after (
		.din(new_net_5749),
		.dout(new_net_5750)
	);

	bfr new_net_5751_bfr_after (
		.din(new_net_5750),
		.dout(new_net_5751)
	);

	bfr new_net_5752_bfr_after (
		.din(new_net_5751),
		.dout(new_net_5752)
	);

	bfr new_net_5753_bfr_after (
		.din(new_net_5752),
		.dout(new_net_5753)
	);

	bfr new_net_5754_bfr_after (
		.din(new_net_5753),
		.dout(new_net_5754)
	);

	bfr new_net_5755_bfr_after (
		.din(new_net_5754),
		.dout(new_net_5755)
	);

	bfr new_net_5756_bfr_after (
		.din(new_net_5755),
		.dout(new_net_5756)
	);

	bfr new_net_5757_bfr_after (
		.din(new_net_5756),
		.dout(new_net_5757)
	);

	bfr new_net_5758_bfr_after (
		.din(new_net_5757),
		.dout(new_net_5758)
	);

	bfr new_net_5759_bfr_after (
		.din(new_net_5758),
		.dout(new_net_5759)
	);

	bfr new_net_5760_bfr_after (
		.din(new_net_5759),
		.dout(new_net_5760)
	);

	bfr new_net_5761_bfr_after (
		.din(new_net_5760),
		.dout(new_net_5761)
	);

	bfr new_net_5762_bfr_after (
		.din(new_net_5761),
		.dout(new_net_5762)
	);

	bfr new_net_5763_bfr_after (
		.din(new_net_5762),
		.dout(new_net_5763)
	);

	bfr new_net_5764_bfr_after (
		.din(new_net_5763),
		.dout(new_net_5764)
	);

	bfr new_net_5765_bfr_after (
		.din(new_net_5764),
		.dout(new_net_5765)
	);

	bfr new_net_5766_bfr_after (
		.din(new_net_5765),
		.dout(new_net_5766)
	);

	bfr new_net_5767_bfr_after (
		.din(new_net_5766),
		.dout(new_net_5767)
	);

	bfr new_net_5768_bfr_after (
		.din(new_net_5767),
		.dout(new_net_5768)
	);

	bfr new_net_5769_bfr_after (
		.din(new_net_5768),
		.dout(new_net_5769)
	);

	bfr new_net_5770_bfr_after (
		.din(new_net_5769),
		.dout(new_net_5770)
	);

	bfr new_net_5771_bfr_after (
		.din(new_net_5770),
		.dout(new_net_5771)
	);

	bfr new_net_5772_bfr_after (
		.din(new_net_5771),
		.dout(new_net_5772)
	);

	bfr new_net_5773_bfr_after (
		.din(new_net_5772),
		.dout(new_net_5773)
	);

	bfr new_net_5774_bfr_after (
		.din(new_net_5773),
		.dout(new_net_5774)
	);

	bfr new_net_5775_bfr_after (
		.din(new_net_5774),
		.dout(new_net_5775)
	);

	bfr new_net_5776_bfr_after (
		.din(new_net_5775),
		.dout(new_net_5776)
	);

	bfr new_net_5777_bfr_after (
		.din(new_net_5776),
		.dout(new_net_5777)
	);

	bfr new_net_5778_bfr_after (
		.din(new_net_5777),
		.dout(new_net_5778)
	);

	bfr new_net_5779_bfr_after (
		.din(new_net_5778),
		.dout(new_net_5779)
	);

	bfr new_net_5780_bfr_after (
		.din(new_net_5779),
		.dout(new_net_5780)
	);

	bfr new_net_5781_bfr_after (
		.din(new_net_5780),
		.dout(new_net_5781)
	);

	bfr new_net_5782_bfr_after (
		.din(new_net_5781),
		.dout(new_net_5782)
	);

	bfr new_net_5783_bfr_after (
		.din(new_net_5782),
		.dout(new_net_5783)
	);

	bfr new_net_5784_bfr_after (
		.din(new_net_5783),
		.dout(new_net_5784)
	);

	bfr new_net_5785_bfr_after (
		.din(new_net_5784),
		.dout(new_net_5785)
	);

	bfr new_net_5786_bfr_after (
		.din(new_net_5785),
		.dout(new_net_5786)
	);

	bfr new_net_5787_bfr_after (
		.din(new_net_5786),
		.dout(new_net_5787)
	);

	bfr new_net_5788_bfr_after (
		.din(new_net_5787),
		.dout(new_net_5788)
	);

	bfr new_net_5789_bfr_after (
		.din(new_net_5788),
		.dout(new_net_5789)
	);

	bfr new_net_5790_bfr_after (
		.din(new_net_5789),
		.dout(new_net_5790)
	);

	bfr new_net_5791_bfr_after (
		.din(new_net_5790),
		.dout(new_net_5791)
	);

	bfr new_net_5792_bfr_after (
		.din(new_net_5791),
		.dout(new_net_5792)
	);

	bfr new_net_5793_bfr_after (
		.din(new_net_5792),
		.dout(new_net_5793)
	);

	bfr new_net_5794_bfr_after (
		.din(new_net_5793),
		.dout(new_net_5794)
	);

	bfr new_net_5795_bfr_after (
		.din(new_net_5794),
		.dout(new_net_5795)
	);

	bfr new_net_5796_bfr_after (
		.din(new_net_5795),
		.dout(new_net_5796)
	);

	bfr new_net_5797_bfr_after (
		.din(new_net_5796),
		.dout(new_net_5797)
	);

	bfr new_net_5798_bfr_after (
		.din(new_net_5797),
		.dout(new_net_5798)
	);

	bfr new_net_5799_bfr_after (
		.din(new_net_5798),
		.dout(new_net_5799)
	);

	bfr new_net_5800_bfr_after (
		.din(new_net_5799),
		.dout(new_net_5800)
	);

	bfr new_net_5801_bfr_after (
		.din(new_net_5800),
		.dout(new_net_5801)
	);

	bfr new_net_5802_bfr_after (
		.din(new_net_5801),
		.dout(new_net_5802)
	);

	bfr new_net_5803_bfr_after (
		.din(new_net_5802),
		.dout(new_net_5803)
	);

	bfr new_net_5804_bfr_after (
		.din(new_net_5803),
		.dout(new_net_5804)
	);

	bfr new_net_5805_bfr_after (
		.din(new_net_5804),
		.dout(new_net_5805)
	);

	bfr new_net_5806_bfr_after (
		.din(new_net_5805),
		.dout(new_net_5806)
	);

	bfr new_net_5807_bfr_after (
		.din(new_net_5806),
		.dout(new_net_5807)
	);

	bfr new_net_5808_bfr_after (
		.din(new_net_5807),
		.dout(new_net_5808)
	);

	bfr new_net_5809_bfr_after (
		.din(new_net_5808),
		.dout(new_net_5809)
	);

	bfr new_net_5810_bfr_after (
		.din(new_net_5809),
		.dout(new_net_5810)
	);

	bfr new_net_5811_bfr_after (
		.din(new_net_5810),
		.dout(new_net_5811)
	);

	bfr new_net_5812_bfr_after (
		.din(new_net_5811),
		.dout(new_net_5812)
	);

	bfr new_net_5813_bfr_after (
		.din(new_net_5812),
		.dout(new_net_5813)
	);

	bfr new_net_5814_bfr_after (
		.din(new_net_5813),
		.dout(new_net_5814)
	);

	spl2 _0703__v_fanout (
		.a(new_net_5814),
		.b(new_net_661),
		.c(new_net_662)
	);

	bfr new_net_5815_bfr_after (
		.din(_0707_),
		.dout(new_net_5815)
	);

	bfr new_net_5816_bfr_after (
		.din(new_net_5815),
		.dout(new_net_5816)
	);

	bfr new_net_5817_bfr_after (
		.din(new_net_5816),
		.dout(new_net_5817)
	);

	bfr new_net_5818_bfr_after (
		.din(new_net_5817),
		.dout(new_net_5818)
	);

	bfr new_net_5819_bfr_after (
		.din(new_net_5818),
		.dout(new_net_5819)
	);

	bfr new_net_5820_bfr_after (
		.din(new_net_5819),
		.dout(new_net_5820)
	);

	bfr new_net_5821_bfr_after (
		.din(new_net_5820),
		.dout(new_net_5821)
	);

	bfr new_net_5822_bfr_after (
		.din(new_net_5821),
		.dout(new_net_5822)
	);

	bfr new_net_5823_bfr_after (
		.din(new_net_5822),
		.dout(new_net_5823)
	);

	bfr new_net_5824_bfr_after (
		.din(new_net_5823),
		.dout(new_net_5824)
	);

	bfr new_net_5825_bfr_after (
		.din(new_net_5824),
		.dout(new_net_5825)
	);

	bfr new_net_5826_bfr_after (
		.din(new_net_5825),
		.dout(new_net_5826)
	);

	bfr new_net_5827_bfr_after (
		.din(new_net_5826),
		.dout(new_net_5827)
	);

	bfr new_net_5828_bfr_after (
		.din(new_net_5827),
		.dout(new_net_5828)
	);

	bfr new_net_5829_bfr_after (
		.din(new_net_5828),
		.dout(new_net_5829)
	);

	bfr new_net_5830_bfr_after (
		.din(new_net_5829),
		.dout(new_net_5830)
	);

	bfr new_net_5831_bfr_after (
		.din(new_net_5830),
		.dout(new_net_5831)
	);

	bfr new_net_5832_bfr_after (
		.din(new_net_5831),
		.dout(new_net_5832)
	);

	bfr new_net_5833_bfr_after (
		.din(new_net_5832),
		.dout(new_net_5833)
	);

	bfr new_net_5834_bfr_after (
		.din(new_net_5833),
		.dout(new_net_5834)
	);

	bfr new_net_5835_bfr_after (
		.din(new_net_5834),
		.dout(new_net_5835)
	);

	bfr new_net_5836_bfr_after (
		.din(new_net_5835),
		.dout(new_net_5836)
	);

	bfr new_net_5837_bfr_after (
		.din(new_net_5836),
		.dout(new_net_5837)
	);

	bfr new_net_5838_bfr_after (
		.din(new_net_5837),
		.dout(new_net_5838)
	);

	bfr new_net_5839_bfr_after (
		.din(new_net_5838),
		.dout(new_net_5839)
	);

	bfr new_net_5840_bfr_after (
		.din(new_net_5839),
		.dout(new_net_5840)
	);

	bfr new_net_5841_bfr_after (
		.din(new_net_5840),
		.dout(new_net_5841)
	);

	bfr new_net_5842_bfr_after (
		.din(new_net_5841),
		.dout(new_net_5842)
	);

	bfr new_net_5843_bfr_after (
		.din(new_net_5842),
		.dout(new_net_5843)
	);

	bfr new_net_5844_bfr_after (
		.din(new_net_5843),
		.dout(new_net_5844)
	);

	bfr new_net_5845_bfr_after (
		.din(new_net_5844),
		.dout(new_net_5845)
	);

	bfr new_net_5846_bfr_after (
		.din(new_net_5845),
		.dout(new_net_5846)
	);

	bfr new_net_5847_bfr_after (
		.din(new_net_5846),
		.dout(new_net_5847)
	);

	bfr new_net_5848_bfr_after (
		.din(new_net_5847),
		.dout(new_net_5848)
	);

	bfr new_net_5849_bfr_after (
		.din(new_net_5848),
		.dout(new_net_5849)
	);

	bfr new_net_5850_bfr_after (
		.din(new_net_5849),
		.dout(new_net_5850)
	);

	bfr new_net_5851_bfr_after (
		.din(new_net_5850),
		.dout(new_net_5851)
	);

	bfr new_net_5852_bfr_after (
		.din(new_net_5851),
		.dout(new_net_5852)
	);

	bfr new_net_5853_bfr_after (
		.din(new_net_5852),
		.dout(new_net_5853)
	);

	bfr new_net_5854_bfr_after (
		.din(new_net_5853),
		.dout(new_net_5854)
	);

	bfr new_net_5855_bfr_after (
		.din(new_net_5854),
		.dout(new_net_5855)
	);

	bfr new_net_5856_bfr_after (
		.din(new_net_5855),
		.dout(new_net_5856)
	);

	bfr new_net_5857_bfr_after (
		.din(new_net_5856),
		.dout(new_net_5857)
	);

	bfr new_net_5858_bfr_after (
		.din(new_net_5857),
		.dout(new_net_5858)
	);

	bfr new_net_5859_bfr_after (
		.din(new_net_5858),
		.dout(new_net_5859)
	);

	bfr new_net_5860_bfr_after (
		.din(new_net_5859),
		.dout(new_net_5860)
	);

	bfr new_net_5861_bfr_after (
		.din(new_net_5860),
		.dout(new_net_5861)
	);

	bfr new_net_5862_bfr_after (
		.din(new_net_5861),
		.dout(new_net_5862)
	);

	bfr new_net_5863_bfr_after (
		.din(new_net_5862),
		.dout(new_net_5863)
	);

	bfr new_net_5864_bfr_after (
		.din(new_net_5863),
		.dout(new_net_5864)
	);

	bfr new_net_5865_bfr_after (
		.din(new_net_5864),
		.dout(new_net_5865)
	);

	bfr new_net_5866_bfr_after (
		.din(new_net_5865),
		.dout(new_net_5866)
	);

	bfr new_net_5867_bfr_after (
		.din(new_net_5866),
		.dout(new_net_5867)
	);

	bfr new_net_5868_bfr_after (
		.din(new_net_5867),
		.dout(new_net_5868)
	);

	bfr new_net_5869_bfr_after (
		.din(new_net_5868),
		.dout(new_net_5869)
	);

	bfr new_net_5870_bfr_after (
		.din(new_net_5869),
		.dout(new_net_5870)
	);

	bfr new_net_5871_bfr_after (
		.din(new_net_5870),
		.dout(new_net_5871)
	);

	bfr new_net_5872_bfr_after (
		.din(new_net_5871),
		.dout(new_net_5872)
	);

	bfr new_net_5873_bfr_after (
		.din(new_net_5872),
		.dout(new_net_5873)
	);

	bfr new_net_5874_bfr_after (
		.din(new_net_5873),
		.dout(new_net_5874)
	);

	bfr new_net_5875_bfr_after (
		.din(new_net_5874),
		.dout(new_net_5875)
	);

	bfr new_net_5876_bfr_after (
		.din(new_net_5875),
		.dout(new_net_5876)
	);

	bfr new_net_5877_bfr_after (
		.din(new_net_5876),
		.dout(new_net_5877)
	);

	bfr new_net_5878_bfr_after (
		.din(new_net_5877),
		.dout(new_net_5878)
	);

	bfr new_net_5879_bfr_after (
		.din(new_net_5878),
		.dout(new_net_5879)
	);

	bfr new_net_5880_bfr_after (
		.din(new_net_5879),
		.dout(new_net_5880)
	);

	bfr new_net_5881_bfr_after (
		.din(new_net_5880),
		.dout(new_net_5881)
	);

	bfr new_net_5882_bfr_after (
		.din(new_net_5881),
		.dout(new_net_5882)
	);

	bfr new_net_5883_bfr_after (
		.din(new_net_5882),
		.dout(new_net_5883)
	);

	bfr new_net_5884_bfr_after (
		.din(new_net_5883),
		.dout(new_net_5884)
	);

	spl2 _0707__v_fanout (
		.a(new_net_5884),
		.b(new_net_458),
		.c(new_net_459)
	);

	bfr new_net_5885_bfr_after (
		.din(_1704_),
		.dout(new_net_5885)
	);

	bfr new_net_5886_bfr_after (
		.din(new_net_5885),
		.dout(new_net_5886)
	);

	bfr new_net_5887_bfr_after (
		.din(new_net_5886),
		.dout(new_net_5887)
	);

	bfr new_net_5888_bfr_after (
		.din(new_net_5887),
		.dout(new_net_5888)
	);

	bfr new_net_5889_bfr_after (
		.din(new_net_5888),
		.dout(new_net_5889)
	);

	bfr new_net_5890_bfr_after (
		.din(new_net_5889),
		.dout(new_net_5890)
	);

	bfr new_net_5891_bfr_after (
		.din(new_net_5890),
		.dout(new_net_5891)
	);

	bfr new_net_5892_bfr_after (
		.din(new_net_5891),
		.dout(new_net_5892)
	);

	bfr new_net_5893_bfr_after (
		.din(new_net_5892),
		.dout(new_net_5893)
	);

	bfr new_net_5894_bfr_after (
		.din(new_net_5893),
		.dout(new_net_5894)
	);

	bfr new_net_5895_bfr_after (
		.din(new_net_5894),
		.dout(new_net_5895)
	);

	bfr new_net_5896_bfr_after (
		.din(new_net_5895),
		.dout(new_net_5896)
	);

	bfr new_net_5897_bfr_after (
		.din(new_net_5896),
		.dout(new_net_5897)
	);

	bfr new_net_5898_bfr_after (
		.din(new_net_5897),
		.dout(new_net_5898)
	);

	bfr new_net_5899_bfr_after (
		.din(new_net_5898),
		.dout(new_net_5899)
	);

	bfr new_net_5900_bfr_after (
		.din(new_net_5899),
		.dout(new_net_5900)
	);

	spl2 _1704__v_fanout (
		.a(new_net_5900),
		.b(new_net_1394),
		.c(new_net_1395)
	);

	bfr new_net_5901_bfr_after (
		.din(_0831_),
		.dout(new_net_5901)
	);

	bfr new_net_5902_bfr_after (
		.din(new_net_5901),
		.dout(new_net_5902)
	);

	bfr new_net_5903_bfr_after (
		.din(new_net_5902),
		.dout(new_net_5903)
	);

	bfr new_net_5904_bfr_after (
		.din(new_net_5903),
		.dout(new_net_5904)
	);

	bfr new_net_5905_bfr_after (
		.din(new_net_5904),
		.dout(new_net_5905)
	);

	bfr new_net_5906_bfr_after (
		.din(new_net_5905),
		.dout(new_net_5906)
	);

	bfr new_net_5907_bfr_after (
		.din(new_net_5906),
		.dout(new_net_5907)
	);

	bfr new_net_5908_bfr_after (
		.din(new_net_5907),
		.dout(new_net_5908)
	);

	bfr new_net_5909_bfr_after (
		.din(new_net_5908),
		.dout(new_net_5909)
	);

	bfr new_net_5910_bfr_after (
		.din(new_net_5909),
		.dout(new_net_5910)
	);

	bfr new_net_5911_bfr_after (
		.din(new_net_5910),
		.dout(new_net_5911)
	);

	bfr new_net_5912_bfr_after (
		.din(new_net_5911),
		.dout(new_net_5912)
	);

	bfr new_net_5913_bfr_after (
		.din(new_net_5912),
		.dout(new_net_5913)
	);

	bfr new_net_5914_bfr_after (
		.din(new_net_5913),
		.dout(new_net_5914)
	);

	bfr new_net_5915_bfr_after (
		.din(new_net_5914),
		.dout(new_net_5915)
	);

	bfr new_net_5916_bfr_after (
		.din(new_net_5915),
		.dout(new_net_5916)
	);

	bfr new_net_5917_bfr_after (
		.din(new_net_5916),
		.dout(new_net_5917)
	);

	bfr new_net_5918_bfr_after (
		.din(new_net_5917),
		.dout(new_net_5918)
	);

	bfr new_net_5919_bfr_after (
		.din(new_net_5918),
		.dout(new_net_5919)
	);

	bfr new_net_5920_bfr_after (
		.din(new_net_5919),
		.dout(new_net_5920)
	);

	bfr new_net_5921_bfr_after (
		.din(new_net_5920),
		.dout(new_net_5921)
	);

	bfr new_net_5922_bfr_after (
		.din(new_net_5921),
		.dout(new_net_5922)
	);

	bfr new_net_5923_bfr_after (
		.din(new_net_5922),
		.dout(new_net_5923)
	);

	bfr new_net_5924_bfr_after (
		.din(new_net_5923),
		.dout(new_net_5924)
	);

	bfr new_net_5925_bfr_after (
		.din(new_net_5924),
		.dout(new_net_5925)
	);

	bfr new_net_5926_bfr_after (
		.din(new_net_5925),
		.dout(new_net_5926)
	);

	bfr new_net_5927_bfr_after (
		.din(new_net_5926),
		.dout(new_net_5927)
	);

	bfr new_net_5928_bfr_after (
		.din(new_net_5927),
		.dout(new_net_5928)
	);

	bfr new_net_5929_bfr_after (
		.din(new_net_5928),
		.dout(new_net_5929)
	);

	bfr new_net_5930_bfr_after (
		.din(new_net_5929),
		.dout(new_net_5930)
	);

	bfr new_net_5931_bfr_after (
		.din(new_net_5930),
		.dout(new_net_5931)
	);

	bfr new_net_5932_bfr_after (
		.din(new_net_5931),
		.dout(new_net_5932)
	);

	bfr new_net_5933_bfr_after (
		.din(new_net_5932),
		.dout(new_net_5933)
	);

	bfr new_net_5934_bfr_after (
		.din(new_net_5933),
		.dout(new_net_5934)
	);

	bfr new_net_5935_bfr_after (
		.din(new_net_5934),
		.dout(new_net_5935)
	);

	bfr new_net_5936_bfr_after (
		.din(new_net_5935),
		.dout(new_net_5936)
	);

	bfr new_net_5937_bfr_after (
		.din(new_net_5936),
		.dout(new_net_5937)
	);

	bfr new_net_5938_bfr_after (
		.din(new_net_5937),
		.dout(new_net_5938)
	);

	bfr new_net_5939_bfr_after (
		.din(new_net_5938),
		.dout(new_net_5939)
	);

	bfr new_net_5940_bfr_after (
		.din(new_net_5939),
		.dout(new_net_5940)
	);

	bfr new_net_5941_bfr_after (
		.din(new_net_5940),
		.dout(new_net_5941)
	);

	bfr new_net_5942_bfr_after (
		.din(new_net_5941),
		.dout(new_net_5942)
	);

	bfr new_net_5943_bfr_after (
		.din(new_net_5942),
		.dout(new_net_5943)
	);

	bfr new_net_5944_bfr_after (
		.din(new_net_5943),
		.dout(new_net_5944)
	);

	bfr new_net_5945_bfr_after (
		.din(new_net_5944),
		.dout(new_net_5945)
	);

	bfr new_net_5946_bfr_after (
		.din(new_net_5945),
		.dout(new_net_5946)
	);

	bfr new_net_5947_bfr_after (
		.din(new_net_5946),
		.dout(new_net_5947)
	);

	bfr new_net_5948_bfr_after (
		.din(new_net_5947),
		.dout(new_net_5948)
	);

	bfr new_net_5949_bfr_after (
		.din(new_net_5948),
		.dout(new_net_5949)
	);

	bfr new_net_5950_bfr_after (
		.din(new_net_5949),
		.dout(new_net_5950)
	);

	bfr new_net_5951_bfr_after (
		.din(new_net_5950),
		.dout(new_net_5951)
	);

	bfr new_net_5952_bfr_after (
		.din(new_net_5951),
		.dout(new_net_5952)
	);

	bfr new_net_5953_bfr_after (
		.din(new_net_5952),
		.dout(new_net_5953)
	);

	bfr new_net_5954_bfr_after (
		.din(new_net_5953),
		.dout(new_net_5954)
	);

	bfr new_net_5955_bfr_after (
		.din(new_net_5954),
		.dout(new_net_5955)
	);

	bfr new_net_5956_bfr_after (
		.din(new_net_5955),
		.dout(new_net_5956)
	);

	bfr new_net_5957_bfr_after (
		.din(new_net_5956),
		.dout(new_net_5957)
	);

	bfr new_net_5958_bfr_after (
		.din(new_net_5957),
		.dout(new_net_5958)
	);

	bfr new_net_5959_bfr_after (
		.din(new_net_5958),
		.dout(new_net_5959)
	);

	bfr new_net_5960_bfr_after (
		.din(new_net_5959),
		.dout(new_net_5960)
	);

	bfr new_net_5961_bfr_after (
		.din(new_net_5960),
		.dout(new_net_5961)
	);

	bfr new_net_5962_bfr_after (
		.din(new_net_5961),
		.dout(new_net_5962)
	);

	bfr new_net_5963_bfr_after (
		.din(new_net_5962),
		.dout(new_net_5963)
	);

	bfr new_net_5964_bfr_after (
		.din(new_net_5963),
		.dout(new_net_5964)
	);

	bfr new_net_5965_bfr_after (
		.din(new_net_5964),
		.dout(new_net_5965)
	);

	bfr new_net_5966_bfr_after (
		.din(new_net_5965),
		.dout(new_net_5966)
	);

	bfr new_net_5967_bfr_after (
		.din(new_net_5966),
		.dout(new_net_5967)
	);

	bfr new_net_5968_bfr_after (
		.din(new_net_5967),
		.dout(new_net_5968)
	);

	bfr new_net_5969_bfr_after (
		.din(new_net_5968),
		.dout(new_net_5969)
	);

	bfr new_net_5970_bfr_after (
		.din(new_net_5969),
		.dout(new_net_5970)
	);

	bfr new_net_5971_bfr_after (
		.din(new_net_5970),
		.dout(new_net_5971)
	);

	bfr new_net_5972_bfr_after (
		.din(new_net_5971),
		.dout(new_net_5972)
	);

	bfr new_net_5973_bfr_after (
		.din(new_net_5972),
		.dout(new_net_5973)
	);

	bfr new_net_5974_bfr_after (
		.din(new_net_5973),
		.dout(new_net_5974)
	);

	bfr new_net_5975_bfr_after (
		.din(new_net_5974),
		.dout(new_net_5975)
	);

	bfr new_net_5976_bfr_after (
		.din(new_net_5975),
		.dout(new_net_5976)
	);

	bfr new_net_5977_bfr_after (
		.din(new_net_5976),
		.dout(new_net_5977)
	);

	bfr new_net_5978_bfr_after (
		.din(new_net_5977),
		.dout(new_net_5978)
	);

	bfr new_net_5979_bfr_after (
		.din(new_net_5978),
		.dout(new_net_5979)
	);

	bfr new_net_5980_bfr_after (
		.din(new_net_5979),
		.dout(new_net_5980)
	);

	bfr new_net_5981_bfr_after (
		.din(new_net_5980),
		.dout(new_net_5981)
	);

	bfr new_net_5982_bfr_after (
		.din(new_net_5981),
		.dout(new_net_5982)
	);

	bfr new_net_5983_bfr_after (
		.din(new_net_5982),
		.dout(new_net_5983)
	);

	bfr new_net_5984_bfr_after (
		.din(new_net_5983),
		.dout(new_net_5984)
	);

	bfr new_net_5985_bfr_after (
		.din(new_net_5984),
		.dout(new_net_5985)
	);

	bfr new_net_5986_bfr_after (
		.din(new_net_5985),
		.dout(new_net_5986)
	);

	bfr new_net_5987_bfr_after (
		.din(new_net_5986),
		.dout(new_net_5987)
	);

	bfr new_net_5988_bfr_after (
		.din(new_net_5987),
		.dout(new_net_5988)
	);

	bfr new_net_5989_bfr_after (
		.din(new_net_5988),
		.dout(new_net_5989)
	);

	bfr new_net_5990_bfr_after (
		.din(new_net_5989),
		.dout(new_net_5990)
	);

	bfr new_net_5991_bfr_after (
		.din(new_net_5990),
		.dout(new_net_5991)
	);

	bfr new_net_5992_bfr_after (
		.din(new_net_5991),
		.dout(new_net_5992)
	);

	bfr new_net_5993_bfr_after (
		.din(new_net_5992),
		.dout(new_net_5993)
	);

	bfr new_net_5994_bfr_after (
		.din(new_net_5993),
		.dout(new_net_5994)
	);

	bfr new_net_5995_bfr_after (
		.din(new_net_5994),
		.dout(new_net_5995)
	);

	bfr new_net_5996_bfr_after (
		.din(new_net_5995),
		.dout(new_net_5996)
	);

	bfr new_net_5997_bfr_after (
		.din(new_net_5996),
		.dout(new_net_5997)
	);

	bfr new_net_5998_bfr_after (
		.din(new_net_5997),
		.dout(new_net_5998)
	);

	bfr new_net_5999_bfr_after (
		.din(new_net_5998),
		.dout(new_net_5999)
	);

	bfr new_net_6000_bfr_after (
		.din(new_net_5999),
		.dout(new_net_6000)
	);

	bfr new_net_6001_bfr_after (
		.din(new_net_6000),
		.dout(new_net_6001)
	);

	bfr new_net_6002_bfr_after (
		.din(new_net_6001),
		.dout(new_net_6002)
	);

	bfr new_net_6003_bfr_after (
		.din(new_net_6002),
		.dout(new_net_6003)
	);

	bfr new_net_6004_bfr_after (
		.din(new_net_6003),
		.dout(new_net_6004)
	);

	spl2 _0831__v_fanout (
		.a(new_net_6004),
		.b(new_net_2294),
		.c(new_net_2295)
	);

	bfr new_net_6005_bfr_after (
		.din(_0778_),
		.dout(new_net_6005)
	);

	bfr new_net_6006_bfr_after (
		.din(new_net_6005),
		.dout(new_net_6006)
	);

	bfr new_net_6007_bfr_after (
		.din(new_net_6006),
		.dout(new_net_6007)
	);

	bfr new_net_6008_bfr_after (
		.din(new_net_6007),
		.dout(new_net_6008)
	);

	bfr new_net_6009_bfr_after (
		.din(new_net_6008),
		.dout(new_net_6009)
	);

	bfr new_net_6010_bfr_after (
		.din(new_net_6009),
		.dout(new_net_6010)
	);

	bfr new_net_6011_bfr_after (
		.din(new_net_6010),
		.dout(new_net_6011)
	);

	bfr new_net_6012_bfr_after (
		.din(new_net_6011),
		.dout(new_net_6012)
	);

	bfr new_net_6013_bfr_after (
		.din(new_net_6012),
		.dout(new_net_6013)
	);

	bfr new_net_6014_bfr_after (
		.din(new_net_6013),
		.dout(new_net_6014)
	);

	bfr new_net_6015_bfr_after (
		.din(new_net_6014),
		.dout(new_net_6015)
	);

	bfr new_net_6016_bfr_after (
		.din(new_net_6015),
		.dout(new_net_6016)
	);

	bfr new_net_6017_bfr_after (
		.din(new_net_6016),
		.dout(new_net_6017)
	);

	bfr new_net_6018_bfr_after (
		.din(new_net_6017),
		.dout(new_net_6018)
	);

	bfr new_net_6019_bfr_after (
		.din(new_net_6018),
		.dout(new_net_6019)
	);

	bfr new_net_6020_bfr_after (
		.din(new_net_6019),
		.dout(new_net_6020)
	);

	bfr new_net_6021_bfr_after (
		.din(new_net_6020),
		.dout(new_net_6021)
	);

	bfr new_net_6022_bfr_after (
		.din(new_net_6021),
		.dout(new_net_6022)
	);

	bfr new_net_6023_bfr_after (
		.din(new_net_6022),
		.dout(new_net_6023)
	);

	bfr new_net_6024_bfr_after (
		.din(new_net_6023),
		.dout(new_net_6024)
	);

	bfr new_net_6025_bfr_after (
		.din(new_net_6024),
		.dout(new_net_6025)
	);

	bfr new_net_6026_bfr_after (
		.din(new_net_6025),
		.dout(new_net_6026)
	);

	bfr new_net_6027_bfr_after (
		.din(new_net_6026),
		.dout(new_net_6027)
	);

	bfr new_net_6028_bfr_after (
		.din(new_net_6027),
		.dout(new_net_6028)
	);

	bfr new_net_6029_bfr_after (
		.din(new_net_6028),
		.dout(new_net_6029)
	);

	bfr new_net_6030_bfr_after (
		.din(new_net_6029),
		.dout(new_net_6030)
	);

	bfr new_net_6031_bfr_after (
		.din(new_net_6030),
		.dout(new_net_6031)
	);

	bfr new_net_6032_bfr_after (
		.din(new_net_6031),
		.dout(new_net_6032)
	);

	bfr new_net_6033_bfr_after (
		.din(new_net_6032),
		.dout(new_net_6033)
	);

	bfr new_net_6034_bfr_after (
		.din(new_net_6033),
		.dout(new_net_6034)
	);

	bfr new_net_6035_bfr_after (
		.din(new_net_6034),
		.dout(new_net_6035)
	);

	bfr new_net_6036_bfr_after (
		.din(new_net_6035),
		.dout(new_net_6036)
	);

	bfr new_net_6037_bfr_after (
		.din(new_net_6036),
		.dout(new_net_6037)
	);

	bfr new_net_6038_bfr_after (
		.din(new_net_6037),
		.dout(new_net_6038)
	);

	bfr new_net_6039_bfr_after (
		.din(new_net_6038),
		.dout(new_net_6039)
	);

	bfr new_net_6040_bfr_after (
		.din(new_net_6039),
		.dout(new_net_6040)
	);

	bfr new_net_6041_bfr_after (
		.din(new_net_6040),
		.dout(new_net_6041)
	);

	bfr new_net_6042_bfr_after (
		.din(new_net_6041),
		.dout(new_net_6042)
	);

	bfr new_net_6043_bfr_after (
		.din(new_net_6042),
		.dout(new_net_6043)
	);

	bfr new_net_6044_bfr_after (
		.din(new_net_6043),
		.dout(new_net_6044)
	);

	bfr new_net_6045_bfr_after (
		.din(new_net_6044),
		.dout(new_net_6045)
	);

	bfr new_net_6046_bfr_after (
		.din(new_net_6045),
		.dout(new_net_6046)
	);

	bfr new_net_6047_bfr_after (
		.din(new_net_6046),
		.dout(new_net_6047)
	);

	bfr new_net_6048_bfr_after (
		.din(new_net_6047),
		.dout(new_net_6048)
	);

	bfr new_net_6049_bfr_after (
		.din(new_net_6048),
		.dout(new_net_6049)
	);

	bfr new_net_6050_bfr_after (
		.din(new_net_6049),
		.dout(new_net_6050)
	);

	bfr new_net_6051_bfr_after (
		.din(new_net_6050),
		.dout(new_net_6051)
	);

	bfr new_net_6052_bfr_after (
		.din(new_net_6051),
		.dout(new_net_6052)
	);

	bfr new_net_6053_bfr_after (
		.din(new_net_6052),
		.dout(new_net_6053)
	);

	bfr new_net_6054_bfr_after (
		.din(new_net_6053),
		.dout(new_net_6054)
	);

	bfr new_net_6055_bfr_after (
		.din(new_net_6054),
		.dout(new_net_6055)
	);

	bfr new_net_6056_bfr_after (
		.din(new_net_6055),
		.dout(new_net_6056)
	);

	bfr new_net_6057_bfr_after (
		.din(new_net_6056),
		.dout(new_net_6057)
	);

	bfr new_net_6058_bfr_after (
		.din(new_net_6057),
		.dout(new_net_6058)
	);

	bfr new_net_6059_bfr_after (
		.din(new_net_6058),
		.dout(new_net_6059)
	);

	bfr new_net_6060_bfr_after (
		.din(new_net_6059),
		.dout(new_net_6060)
	);

	bfr new_net_6061_bfr_after (
		.din(new_net_6060),
		.dout(new_net_6061)
	);

	bfr new_net_6062_bfr_after (
		.din(new_net_6061),
		.dout(new_net_6062)
	);

	bfr new_net_6063_bfr_after (
		.din(new_net_6062),
		.dout(new_net_6063)
	);

	bfr new_net_6064_bfr_after (
		.din(new_net_6063),
		.dout(new_net_6064)
	);

	bfr new_net_6065_bfr_after (
		.din(new_net_6064),
		.dout(new_net_6065)
	);

	bfr new_net_6066_bfr_after (
		.din(new_net_6065),
		.dout(new_net_6066)
	);

	bfr new_net_6067_bfr_after (
		.din(new_net_6066),
		.dout(new_net_6067)
	);

	bfr new_net_6068_bfr_after (
		.din(new_net_6067),
		.dout(new_net_6068)
	);

	bfr new_net_6069_bfr_after (
		.din(new_net_6068),
		.dout(new_net_6069)
	);

	bfr new_net_6070_bfr_after (
		.din(new_net_6069),
		.dout(new_net_6070)
	);

	spl2 _0778__v_fanout (
		.a(new_net_6070),
		.b(new_net_315),
		.c(new_net_316)
	);

	bfr new_net_6071_bfr_after (
		.din(_0095_),
		.dout(new_net_6071)
	);

	bfr new_net_6072_bfr_after (
		.din(new_net_6071),
		.dout(new_net_6072)
	);

	bfr new_net_6073_bfr_after (
		.din(new_net_6072),
		.dout(new_net_6073)
	);

	bfr new_net_6074_bfr_after (
		.din(new_net_6073),
		.dout(new_net_6074)
	);

	bfr new_net_6075_bfr_after (
		.din(new_net_6074),
		.dout(new_net_6075)
	);

	bfr new_net_6076_bfr_after (
		.din(new_net_6075),
		.dout(new_net_6076)
	);

	bfr new_net_6077_bfr_after (
		.din(new_net_6076),
		.dout(new_net_6077)
	);

	bfr new_net_6078_bfr_after (
		.din(new_net_6077),
		.dout(new_net_6078)
	);

	bfr new_net_6079_bfr_after (
		.din(new_net_6078),
		.dout(new_net_6079)
	);

	bfr new_net_6080_bfr_after (
		.din(new_net_6079),
		.dout(new_net_6080)
	);

	bfr new_net_6081_bfr_after (
		.din(new_net_6080),
		.dout(new_net_6081)
	);

	bfr new_net_6082_bfr_after (
		.din(new_net_6081),
		.dout(new_net_6082)
	);

	bfr new_net_6083_bfr_after (
		.din(new_net_6082),
		.dout(new_net_6083)
	);

	bfr new_net_6084_bfr_after (
		.din(new_net_6083),
		.dout(new_net_6084)
	);

	bfr new_net_6085_bfr_after (
		.din(new_net_6084),
		.dout(new_net_6085)
	);

	bfr new_net_6086_bfr_after (
		.din(new_net_6085),
		.dout(new_net_6086)
	);

	bfr new_net_6087_bfr_after (
		.din(new_net_6086),
		.dout(new_net_6087)
	);

	bfr new_net_6088_bfr_after (
		.din(new_net_6087),
		.dout(new_net_6088)
	);

	bfr new_net_6089_bfr_after (
		.din(new_net_6088),
		.dout(new_net_6089)
	);

	bfr new_net_6090_bfr_after (
		.din(new_net_6089),
		.dout(new_net_6090)
	);

	bfr new_net_6091_bfr_after (
		.din(new_net_6090),
		.dout(new_net_6091)
	);

	bfr new_net_6092_bfr_after (
		.din(new_net_6091),
		.dout(new_net_6092)
	);

	bfr new_net_6093_bfr_after (
		.din(new_net_6092),
		.dout(new_net_6093)
	);

	bfr new_net_6094_bfr_after (
		.din(new_net_6093),
		.dout(new_net_6094)
	);

	bfr new_net_6095_bfr_after (
		.din(new_net_6094),
		.dout(new_net_6095)
	);

	bfr new_net_6096_bfr_after (
		.din(new_net_6095),
		.dout(new_net_6096)
	);

	bfr new_net_6097_bfr_after (
		.din(new_net_6096),
		.dout(new_net_6097)
	);

	bfr new_net_6098_bfr_after (
		.din(new_net_6097),
		.dout(new_net_6098)
	);

	bfr new_net_6099_bfr_after (
		.din(new_net_6098),
		.dout(new_net_6099)
	);

	bfr new_net_6100_bfr_after (
		.din(new_net_6099),
		.dout(new_net_6100)
	);

	bfr new_net_6101_bfr_after (
		.din(new_net_6100),
		.dout(new_net_6101)
	);

	bfr new_net_6102_bfr_after (
		.din(new_net_6101),
		.dout(new_net_6102)
	);

	bfr new_net_6103_bfr_after (
		.din(new_net_6102),
		.dout(new_net_6103)
	);

	bfr new_net_6104_bfr_after (
		.din(new_net_6103),
		.dout(new_net_6104)
	);

	bfr new_net_6105_bfr_after (
		.din(new_net_6104),
		.dout(new_net_6105)
	);

	bfr new_net_6106_bfr_after (
		.din(new_net_6105),
		.dout(new_net_6106)
	);

	bfr new_net_6107_bfr_after (
		.din(new_net_6106),
		.dout(new_net_6107)
	);

	bfr new_net_6108_bfr_after (
		.din(new_net_6107),
		.dout(new_net_6108)
	);

	bfr new_net_6109_bfr_after (
		.din(new_net_6108),
		.dout(new_net_6109)
	);

	bfr new_net_6110_bfr_after (
		.din(new_net_6109),
		.dout(new_net_6110)
	);

	bfr new_net_6111_bfr_after (
		.din(new_net_6110),
		.dout(new_net_6111)
	);

	bfr new_net_6112_bfr_after (
		.din(new_net_6111),
		.dout(new_net_6112)
	);

	bfr new_net_6113_bfr_after (
		.din(new_net_6112),
		.dout(new_net_6113)
	);

	bfr new_net_6114_bfr_after (
		.din(new_net_6113),
		.dout(new_net_6114)
	);

	bfr new_net_6115_bfr_after (
		.din(new_net_6114),
		.dout(new_net_6115)
	);

	bfr new_net_6116_bfr_after (
		.din(new_net_6115),
		.dout(new_net_6116)
	);

	bfr new_net_6117_bfr_after (
		.din(new_net_6116),
		.dout(new_net_6117)
	);

	bfr new_net_6118_bfr_after (
		.din(new_net_6117),
		.dout(new_net_6118)
	);

	bfr new_net_6119_bfr_after (
		.din(new_net_6118),
		.dout(new_net_6119)
	);

	bfr new_net_6120_bfr_after (
		.din(new_net_6119),
		.dout(new_net_6120)
	);

	bfr new_net_6121_bfr_after (
		.din(new_net_6120),
		.dout(new_net_6121)
	);

	bfr new_net_6122_bfr_after (
		.din(new_net_6121),
		.dout(new_net_6122)
	);

	bfr new_net_6123_bfr_after (
		.din(new_net_6122),
		.dout(new_net_6123)
	);

	bfr new_net_6124_bfr_after (
		.din(new_net_6123),
		.dout(new_net_6124)
	);

	bfr new_net_6125_bfr_after (
		.din(new_net_6124),
		.dout(new_net_6125)
	);

	bfr new_net_6126_bfr_after (
		.din(new_net_6125),
		.dout(new_net_6126)
	);

	bfr new_net_6127_bfr_after (
		.din(new_net_6126),
		.dout(new_net_6127)
	);

	bfr new_net_6128_bfr_after (
		.din(new_net_6127),
		.dout(new_net_6128)
	);

	bfr new_net_6129_bfr_after (
		.din(new_net_6128),
		.dout(new_net_6129)
	);

	bfr new_net_6130_bfr_after (
		.din(new_net_6129),
		.dout(new_net_6130)
	);

	bfr new_net_6131_bfr_after (
		.din(new_net_6130),
		.dout(new_net_6131)
	);

	bfr new_net_6132_bfr_after (
		.din(new_net_6131),
		.dout(new_net_6132)
	);

	bfr new_net_6133_bfr_after (
		.din(new_net_6132),
		.dout(new_net_6133)
	);

	bfr new_net_6134_bfr_after (
		.din(new_net_6133),
		.dout(new_net_6134)
	);

	bfr new_net_6135_bfr_after (
		.din(new_net_6134),
		.dout(new_net_6135)
	);

	bfr new_net_6136_bfr_after (
		.din(new_net_6135),
		.dout(new_net_6136)
	);

	bfr new_net_6137_bfr_after (
		.din(new_net_6136),
		.dout(new_net_6137)
	);

	bfr new_net_6138_bfr_after (
		.din(new_net_6137),
		.dout(new_net_6138)
	);

	bfr new_net_6139_bfr_after (
		.din(new_net_6138),
		.dout(new_net_6139)
	);

	bfr new_net_6140_bfr_after (
		.din(new_net_6139),
		.dout(new_net_6140)
	);

	bfr new_net_6141_bfr_after (
		.din(new_net_6140),
		.dout(new_net_6141)
	);

	bfr new_net_6142_bfr_after (
		.din(new_net_6141),
		.dout(new_net_6142)
	);

	spl2 _0095__v_fanout (
		.a(new_net_6142),
		.b(new_net_721),
		.c(new_net_722)
	);

	bfr new_net_6143_bfr_after (
		.din(_0333_),
		.dout(new_net_6143)
	);

	bfr new_net_6144_bfr_after (
		.din(new_net_6143),
		.dout(new_net_6144)
	);

	bfr new_net_6145_bfr_after (
		.din(new_net_6144),
		.dout(new_net_6145)
	);

	bfr new_net_6146_bfr_after (
		.din(new_net_6145),
		.dout(new_net_6146)
	);

	bfr new_net_6147_bfr_after (
		.din(new_net_6146),
		.dout(new_net_6147)
	);

	bfr new_net_6148_bfr_after (
		.din(new_net_6147),
		.dout(new_net_6148)
	);

	bfr new_net_6149_bfr_after (
		.din(new_net_6148),
		.dout(new_net_6149)
	);

	bfr new_net_6150_bfr_after (
		.din(new_net_6149),
		.dout(new_net_6150)
	);

	bfr new_net_6151_bfr_after (
		.din(new_net_6150),
		.dout(new_net_6151)
	);

	bfr new_net_6152_bfr_after (
		.din(new_net_6151),
		.dout(new_net_6152)
	);

	bfr new_net_6153_bfr_after (
		.din(new_net_6152),
		.dout(new_net_6153)
	);

	bfr new_net_6154_bfr_after (
		.din(new_net_6153),
		.dout(new_net_6154)
	);

	bfr new_net_6155_bfr_after (
		.din(new_net_6154),
		.dout(new_net_6155)
	);

	bfr new_net_6156_bfr_after (
		.din(new_net_6155),
		.dout(new_net_6156)
	);

	bfr new_net_6157_bfr_after (
		.din(new_net_6156),
		.dout(new_net_6157)
	);

	bfr new_net_6158_bfr_after (
		.din(new_net_6157),
		.dout(new_net_6158)
	);

	bfr new_net_6159_bfr_after (
		.din(new_net_6158),
		.dout(new_net_6159)
	);

	bfr new_net_6160_bfr_after (
		.din(new_net_6159),
		.dout(new_net_6160)
	);

	bfr new_net_6161_bfr_after (
		.din(new_net_6160),
		.dout(new_net_6161)
	);

	bfr new_net_6162_bfr_after (
		.din(new_net_6161),
		.dout(new_net_6162)
	);

	bfr new_net_6163_bfr_after (
		.din(new_net_6162),
		.dout(new_net_6163)
	);

	bfr new_net_6164_bfr_after (
		.din(new_net_6163),
		.dout(new_net_6164)
	);

	bfr new_net_6165_bfr_after (
		.din(new_net_6164),
		.dout(new_net_6165)
	);

	bfr new_net_6166_bfr_after (
		.din(new_net_6165),
		.dout(new_net_6166)
	);

	bfr new_net_6167_bfr_after (
		.din(new_net_6166),
		.dout(new_net_6167)
	);

	bfr new_net_6168_bfr_after (
		.din(new_net_6167),
		.dout(new_net_6168)
	);

	bfr new_net_6169_bfr_after (
		.din(new_net_6168),
		.dout(new_net_6169)
	);

	bfr new_net_6170_bfr_after (
		.din(new_net_6169),
		.dout(new_net_6170)
	);

	bfr new_net_6171_bfr_after (
		.din(new_net_6170),
		.dout(new_net_6171)
	);

	bfr new_net_6172_bfr_after (
		.din(new_net_6171),
		.dout(new_net_6172)
	);

	bfr new_net_6173_bfr_after (
		.din(new_net_6172),
		.dout(new_net_6173)
	);

	bfr new_net_6174_bfr_after (
		.din(new_net_6173),
		.dout(new_net_6174)
	);

	bfr new_net_6175_bfr_after (
		.din(new_net_6174),
		.dout(new_net_6175)
	);

	bfr new_net_6176_bfr_after (
		.din(new_net_6175),
		.dout(new_net_6176)
	);

	bfr new_net_6177_bfr_after (
		.din(new_net_6176),
		.dout(new_net_6177)
	);

	bfr new_net_6178_bfr_after (
		.din(new_net_6177),
		.dout(new_net_6178)
	);

	bfr new_net_6179_bfr_after (
		.din(new_net_6178),
		.dout(new_net_6179)
	);

	bfr new_net_6180_bfr_after (
		.din(new_net_6179),
		.dout(new_net_6180)
	);

	bfr new_net_6181_bfr_after (
		.din(new_net_6180),
		.dout(new_net_6181)
	);

	bfr new_net_6182_bfr_after (
		.din(new_net_6181),
		.dout(new_net_6182)
	);

	bfr new_net_6183_bfr_after (
		.din(new_net_6182),
		.dout(new_net_6183)
	);

	bfr new_net_6184_bfr_after (
		.din(new_net_6183),
		.dout(new_net_6184)
	);

	bfr new_net_6185_bfr_after (
		.din(new_net_6184),
		.dout(new_net_6185)
	);

	bfr new_net_6186_bfr_after (
		.din(new_net_6185),
		.dout(new_net_6186)
	);

	bfr new_net_6187_bfr_after (
		.din(new_net_6186),
		.dout(new_net_6187)
	);

	bfr new_net_6188_bfr_after (
		.din(new_net_6187),
		.dout(new_net_6188)
	);

	bfr new_net_6189_bfr_after (
		.din(new_net_6188),
		.dout(new_net_6189)
	);

	bfr new_net_6190_bfr_after (
		.din(new_net_6189),
		.dout(new_net_6190)
	);

	bfr new_net_6191_bfr_after (
		.din(new_net_6190),
		.dout(new_net_6191)
	);

	bfr new_net_6192_bfr_after (
		.din(new_net_6191),
		.dout(new_net_6192)
	);

	bfr new_net_6193_bfr_after (
		.din(new_net_6192),
		.dout(new_net_6193)
	);

	bfr new_net_6194_bfr_after (
		.din(new_net_6193),
		.dout(new_net_6194)
	);

	bfr new_net_6195_bfr_after (
		.din(new_net_6194),
		.dout(new_net_6195)
	);

	bfr new_net_6196_bfr_after (
		.din(new_net_6195),
		.dout(new_net_6196)
	);

	bfr new_net_6197_bfr_after (
		.din(new_net_6196),
		.dout(new_net_6197)
	);

	bfr new_net_6198_bfr_after (
		.din(new_net_6197),
		.dout(new_net_6198)
	);

	bfr new_net_6199_bfr_after (
		.din(new_net_6198),
		.dout(new_net_6199)
	);

	bfr new_net_6200_bfr_after (
		.din(new_net_6199),
		.dout(new_net_6200)
	);

	bfr new_net_6201_bfr_after (
		.din(new_net_6200),
		.dout(new_net_6201)
	);

	bfr new_net_6202_bfr_after (
		.din(new_net_6201),
		.dout(new_net_6202)
	);

	bfr new_net_6203_bfr_after (
		.din(new_net_6202),
		.dout(new_net_6203)
	);

	bfr new_net_6204_bfr_after (
		.din(new_net_6203),
		.dout(new_net_6204)
	);

	bfr new_net_6205_bfr_after (
		.din(new_net_6204),
		.dout(new_net_6205)
	);

	bfr new_net_6206_bfr_after (
		.din(new_net_6205),
		.dout(new_net_6206)
	);

	bfr new_net_6207_bfr_after (
		.din(new_net_6206),
		.dout(new_net_6207)
	);

	bfr new_net_6208_bfr_after (
		.din(new_net_6207),
		.dout(new_net_6208)
	);

	bfr new_net_6209_bfr_after (
		.din(new_net_6208),
		.dout(new_net_6209)
	);

	bfr new_net_6210_bfr_after (
		.din(new_net_6209),
		.dout(new_net_6210)
	);

	bfr new_net_6211_bfr_after (
		.din(new_net_6210),
		.dout(new_net_6211)
	);

	bfr new_net_6212_bfr_after (
		.din(new_net_6211),
		.dout(new_net_6212)
	);

	bfr new_net_6213_bfr_after (
		.din(new_net_6212),
		.dout(new_net_6213)
	);

	bfr new_net_6214_bfr_after (
		.din(new_net_6213),
		.dout(new_net_6214)
	);

	bfr new_net_6215_bfr_after (
		.din(new_net_6214),
		.dout(new_net_6215)
	);

	bfr new_net_6216_bfr_after (
		.din(new_net_6215),
		.dout(new_net_6216)
	);

	bfr new_net_6217_bfr_after (
		.din(new_net_6216),
		.dout(new_net_6217)
	);

	bfr new_net_6218_bfr_after (
		.din(new_net_6217),
		.dout(new_net_6218)
	);

	bfr new_net_6219_bfr_after (
		.din(new_net_6218),
		.dout(new_net_6219)
	);

	bfr new_net_6220_bfr_after (
		.din(new_net_6219),
		.dout(new_net_6220)
	);

	bfr new_net_6221_bfr_after (
		.din(new_net_6220),
		.dout(new_net_6221)
	);

	bfr new_net_6222_bfr_after (
		.din(new_net_6221),
		.dout(new_net_6222)
	);

	bfr new_net_6223_bfr_after (
		.din(new_net_6222),
		.dout(new_net_6223)
	);

	bfr new_net_6224_bfr_after (
		.din(new_net_6223),
		.dout(new_net_6224)
	);

	bfr new_net_6225_bfr_after (
		.din(new_net_6224),
		.dout(new_net_6225)
	);

	bfr new_net_6226_bfr_after (
		.din(new_net_6225),
		.dout(new_net_6226)
	);

	bfr new_net_6227_bfr_after (
		.din(new_net_6226),
		.dout(new_net_6227)
	);

	bfr new_net_6228_bfr_after (
		.din(new_net_6227),
		.dout(new_net_6228)
	);

	bfr new_net_6229_bfr_after (
		.din(new_net_6228),
		.dout(new_net_6229)
	);

	bfr new_net_6230_bfr_after (
		.din(new_net_6229),
		.dout(new_net_6230)
	);

	spl2 _0333__v_fanout (
		.a(new_net_6230),
		.b(new_net_3169),
		.c(new_net_3170)
	);

	bfr new_net_6231_bfr_after (
		.din(_1472_),
		.dout(new_net_6231)
	);

	bfr new_net_6232_bfr_after (
		.din(new_net_6231),
		.dout(new_net_6232)
	);

	bfr new_net_6233_bfr_after (
		.din(new_net_6232),
		.dout(new_net_6233)
	);

	bfr new_net_6234_bfr_after (
		.din(new_net_6233),
		.dout(new_net_6234)
	);

	bfr new_net_6235_bfr_after (
		.din(new_net_6234),
		.dout(new_net_6235)
	);

	bfr new_net_6236_bfr_after (
		.din(new_net_6235),
		.dout(new_net_6236)
	);

	bfr new_net_6237_bfr_after (
		.din(new_net_6236),
		.dout(new_net_6237)
	);

	bfr new_net_6238_bfr_after (
		.din(new_net_6237),
		.dout(new_net_6238)
	);

	bfr new_net_6239_bfr_after (
		.din(new_net_6238),
		.dout(new_net_6239)
	);

	bfr new_net_6240_bfr_after (
		.din(new_net_6239),
		.dout(new_net_6240)
	);

	bfr new_net_6241_bfr_after (
		.din(new_net_6240),
		.dout(new_net_6241)
	);

	bfr new_net_6242_bfr_after (
		.din(new_net_6241),
		.dout(new_net_6242)
	);

	bfr new_net_6243_bfr_after (
		.din(new_net_6242),
		.dout(new_net_6243)
	);

	bfr new_net_6244_bfr_after (
		.din(new_net_6243),
		.dout(new_net_6244)
	);

	bfr new_net_6245_bfr_after (
		.din(new_net_6244),
		.dout(new_net_6245)
	);

	bfr new_net_6246_bfr_after (
		.din(new_net_6245),
		.dout(new_net_6246)
	);

	bfr new_net_6247_bfr_after (
		.din(new_net_6246),
		.dout(new_net_6247)
	);

	bfr new_net_6248_bfr_after (
		.din(new_net_6247),
		.dout(new_net_6248)
	);

	bfr new_net_6249_bfr_after (
		.din(new_net_6248),
		.dout(new_net_6249)
	);

	bfr new_net_6250_bfr_after (
		.din(new_net_6249),
		.dout(new_net_6250)
	);

	bfr new_net_6251_bfr_after (
		.din(new_net_6250),
		.dout(new_net_6251)
	);

	bfr new_net_6252_bfr_after (
		.din(new_net_6251),
		.dout(new_net_6252)
	);

	bfr new_net_6253_bfr_after (
		.din(new_net_6252),
		.dout(new_net_6253)
	);

	bfr new_net_6254_bfr_after (
		.din(new_net_6253),
		.dout(new_net_6254)
	);

	spl2 _1472__v_fanout (
		.a(new_net_6254),
		.b(new_net_2000),
		.c(new_net_2001)
	);

	spl2 _0742__v_fanout (
		.a(_0742_),
		.b(new_net_548),
		.c(new_net_549)
	);

	bfr new_net_6255_bfr_after (
		.din(_1207_),
		.dout(new_net_6255)
	);

	bfr new_net_6256_bfr_after (
		.din(new_net_6255),
		.dout(new_net_6256)
	);

	bfr new_net_6257_bfr_after (
		.din(new_net_6256),
		.dout(new_net_6257)
	);

	bfr new_net_6258_bfr_after (
		.din(new_net_6257),
		.dout(new_net_6258)
	);

	bfr new_net_6259_bfr_after (
		.din(new_net_6258),
		.dout(new_net_6259)
	);

	bfr new_net_6260_bfr_after (
		.din(new_net_6259),
		.dout(new_net_6260)
	);

	bfr new_net_6261_bfr_after (
		.din(new_net_6260),
		.dout(new_net_6261)
	);

	bfr new_net_6262_bfr_after (
		.din(new_net_6261),
		.dout(new_net_6262)
	);

	bfr new_net_6263_bfr_after (
		.din(new_net_6262),
		.dout(new_net_6263)
	);

	bfr new_net_6264_bfr_after (
		.din(new_net_6263),
		.dout(new_net_6264)
	);

	bfr new_net_6265_bfr_after (
		.din(new_net_6264),
		.dout(new_net_6265)
	);

	bfr new_net_6266_bfr_after (
		.din(new_net_6265),
		.dout(new_net_6266)
	);

	bfr new_net_6267_bfr_after (
		.din(new_net_6266),
		.dout(new_net_6267)
	);

	bfr new_net_6268_bfr_after (
		.din(new_net_6267),
		.dout(new_net_6268)
	);

	bfr new_net_6269_bfr_after (
		.din(new_net_6268),
		.dout(new_net_6269)
	);

	bfr new_net_6270_bfr_after (
		.din(new_net_6269),
		.dout(new_net_6270)
	);

	bfr new_net_6271_bfr_after (
		.din(new_net_6270),
		.dout(new_net_6271)
	);

	bfr new_net_6272_bfr_after (
		.din(new_net_6271),
		.dout(new_net_6272)
	);

	bfr new_net_6273_bfr_after (
		.din(new_net_6272),
		.dout(new_net_6273)
	);

	bfr new_net_6274_bfr_after (
		.din(new_net_6273),
		.dout(new_net_6274)
	);

	bfr new_net_6275_bfr_after (
		.din(new_net_6274),
		.dout(new_net_6275)
	);

	bfr new_net_6276_bfr_after (
		.din(new_net_6275),
		.dout(new_net_6276)
	);

	bfr new_net_6277_bfr_after (
		.din(new_net_6276),
		.dout(new_net_6277)
	);

	bfr new_net_6278_bfr_after (
		.din(new_net_6277),
		.dout(new_net_6278)
	);

	bfr new_net_6279_bfr_after (
		.din(new_net_6278),
		.dout(new_net_6279)
	);

	bfr new_net_6280_bfr_after (
		.din(new_net_6279),
		.dout(new_net_6280)
	);

	bfr new_net_6281_bfr_after (
		.din(new_net_6280),
		.dout(new_net_6281)
	);

	bfr new_net_6282_bfr_after (
		.din(new_net_6281),
		.dout(new_net_6282)
	);

	bfr new_net_6283_bfr_after (
		.din(new_net_6282),
		.dout(new_net_6283)
	);

	bfr new_net_6284_bfr_after (
		.din(new_net_6283),
		.dout(new_net_6284)
	);

	bfr new_net_6285_bfr_after (
		.din(new_net_6284),
		.dout(new_net_6285)
	);

	bfr new_net_6286_bfr_after (
		.din(new_net_6285),
		.dout(new_net_6286)
	);

	bfr new_net_6287_bfr_after (
		.din(new_net_6286),
		.dout(new_net_6287)
	);

	bfr new_net_6288_bfr_after (
		.din(new_net_6287),
		.dout(new_net_6288)
	);

	bfr new_net_6289_bfr_after (
		.din(new_net_6288),
		.dout(new_net_6289)
	);

	bfr new_net_6290_bfr_after (
		.din(new_net_6289),
		.dout(new_net_6290)
	);

	bfr new_net_6291_bfr_after (
		.din(new_net_6290),
		.dout(new_net_6291)
	);

	bfr new_net_6292_bfr_after (
		.din(new_net_6291),
		.dout(new_net_6292)
	);

	bfr new_net_6293_bfr_after (
		.din(new_net_6292),
		.dout(new_net_6293)
	);

	bfr new_net_6294_bfr_after (
		.din(new_net_6293),
		.dout(new_net_6294)
	);

	bfr new_net_6295_bfr_after (
		.din(new_net_6294),
		.dout(new_net_6295)
	);

	bfr new_net_6296_bfr_after (
		.din(new_net_6295),
		.dout(new_net_6296)
	);

	bfr new_net_6297_bfr_after (
		.din(new_net_6296),
		.dout(new_net_6297)
	);

	bfr new_net_6298_bfr_after (
		.din(new_net_6297),
		.dout(new_net_6298)
	);

	bfr new_net_6299_bfr_after (
		.din(new_net_6298),
		.dout(new_net_6299)
	);

	bfr new_net_6300_bfr_after (
		.din(new_net_6299),
		.dout(new_net_6300)
	);

	bfr new_net_6301_bfr_after (
		.din(new_net_6300),
		.dout(new_net_6301)
	);

	bfr new_net_6302_bfr_after (
		.din(new_net_6301),
		.dout(new_net_6302)
	);

	bfr new_net_6303_bfr_after (
		.din(new_net_6302),
		.dout(new_net_6303)
	);

	bfr new_net_6304_bfr_after (
		.din(new_net_6303),
		.dout(new_net_6304)
	);

	bfr new_net_6305_bfr_after (
		.din(new_net_6304),
		.dout(new_net_6305)
	);

	bfr new_net_6306_bfr_after (
		.din(new_net_6305),
		.dout(new_net_6306)
	);

	bfr new_net_6307_bfr_after (
		.din(new_net_6306),
		.dout(new_net_6307)
	);

	bfr new_net_6308_bfr_after (
		.din(new_net_6307),
		.dout(new_net_6308)
	);

	bfr new_net_6309_bfr_after (
		.din(new_net_6308),
		.dout(new_net_6309)
	);

	bfr new_net_6310_bfr_after (
		.din(new_net_6309),
		.dout(new_net_6310)
	);

	spl2 _1207__v_fanout (
		.a(new_net_6310),
		.b(new_net_496),
		.c(new_net_497)
	);

	bfr new_net_6311_bfr_after (
		.din(_1571_),
		.dout(new_net_6311)
	);

	bfr new_net_6312_bfr_after (
		.din(new_net_6311),
		.dout(new_net_6312)
	);

	bfr new_net_6313_bfr_after (
		.din(new_net_6312),
		.dout(new_net_6313)
	);

	bfr new_net_6314_bfr_after (
		.din(new_net_6313),
		.dout(new_net_6314)
	);

	bfr new_net_6315_bfr_after (
		.din(new_net_6314),
		.dout(new_net_6315)
	);

	bfr new_net_6316_bfr_after (
		.din(new_net_6315),
		.dout(new_net_6316)
	);

	bfr new_net_6317_bfr_after (
		.din(new_net_6316),
		.dout(new_net_6317)
	);

	bfr new_net_6318_bfr_after (
		.din(new_net_6317),
		.dout(new_net_6318)
	);

	bfr new_net_6319_bfr_after (
		.din(new_net_6318),
		.dout(new_net_6319)
	);

	bfr new_net_6320_bfr_after (
		.din(new_net_6319),
		.dout(new_net_6320)
	);

	bfr new_net_6321_bfr_after (
		.din(new_net_6320),
		.dout(new_net_6321)
	);

	bfr new_net_6322_bfr_after (
		.din(new_net_6321),
		.dout(new_net_6322)
	);

	bfr new_net_6323_bfr_after (
		.din(new_net_6322),
		.dout(new_net_6323)
	);

	bfr new_net_6324_bfr_after (
		.din(new_net_6323),
		.dout(new_net_6324)
	);

	bfr new_net_6325_bfr_after (
		.din(new_net_6324),
		.dout(new_net_6325)
	);

	bfr new_net_6326_bfr_after (
		.din(new_net_6325),
		.dout(new_net_6326)
	);

	bfr new_net_6327_bfr_after (
		.din(new_net_6326),
		.dout(new_net_6327)
	);

	bfr new_net_6328_bfr_after (
		.din(new_net_6327),
		.dout(new_net_6328)
	);

	bfr new_net_6329_bfr_after (
		.din(new_net_6328),
		.dout(new_net_6329)
	);

	bfr new_net_6330_bfr_after (
		.din(new_net_6329),
		.dout(new_net_6330)
	);

	bfr new_net_6331_bfr_after (
		.din(new_net_6330),
		.dout(new_net_6331)
	);

	bfr new_net_6332_bfr_after (
		.din(new_net_6331),
		.dout(new_net_6332)
	);

	bfr new_net_6333_bfr_after (
		.din(new_net_6332),
		.dout(new_net_6333)
	);

	bfr new_net_6334_bfr_after (
		.din(new_net_6333),
		.dout(new_net_6334)
	);

	bfr new_net_6335_bfr_after (
		.din(new_net_6334),
		.dout(new_net_6335)
	);

	bfr new_net_6336_bfr_after (
		.din(new_net_6335),
		.dout(new_net_6336)
	);

	bfr new_net_6337_bfr_after (
		.din(new_net_6336),
		.dout(new_net_6337)
	);

	bfr new_net_6338_bfr_after (
		.din(new_net_6337),
		.dout(new_net_6338)
	);

	bfr new_net_6339_bfr_after (
		.din(new_net_6338),
		.dout(new_net_6339)
	);

	bfr new_net_6340_bfr_after (
		.din(new_net_6339),
		.dout(new_net_6340)
	);

	bfr new_net_6341_bfr_after (
		.din(new_net_6340),
		.dout(new_net_6341)
	);

	bfr new_net_6342_bfr_after (
		.din(new_net_6341),
		.dout(new_net_6342)
	);

	bfr new_net_6343_bfr_after (
		.din(new_net_6342),
		.dout(new_net_6343)
	);

	bfr new_net_6344_bfr_after (
		.din(new_net_6343),
		.dout(new_net_6344)
	);

	bfr new_net_6345_bfr_after (
		.din(new_net_6344),
		.dout(new_net_6345)
	);

	bfr new_net_6346_bfr_after (
		.din(new_net_6345),
		.dout(new_net_6346)
	);

	bfr new_net_6347_bfr_after (
		.din(new_net_6346),
		.dout(new_net_6347)
	);

	bfr new_net_6348_bfr_after (
		.din(new_net_6347),
		.dout(new_net_6348)
	);

	bfr new_net_6349_bfr_after (
		.din(new_net_6348),
		.dout(new_net_6349)
	);

	bfr new_net_6350_bfr_after (
		.din(new_net_6349),
		.dout(new_net_6350)
	);

	bfr new_net_6351_bfr_after (
		.din(new_net_6350),
		.dout(new_net_6351)
	);

	bfr new_net_6352_bfr_after (
		.din(new_net_6351),
		.dout(new_net_6352)
	);

	bfr new_net_6353_bfr_after (
		.din(new_net_6352),
		.dout(new_net_6353)
	);

	bfr new_net_6354_bfr_after (
		.din(new_net_6353),
		.dout(new_net_6354)
	);

	bfr new_net_6355_bfr_after (
		.din(new_net_6354),
		.dout(new_net_6355)
	);

	bfr new_net_6356_bfr_after (
		.din(new_net_6355),
		.dout(new_net_6356)
	);

	bfr new_net_6357_bfr_after (
		.din(new_net_6356),
		.dout(new_net_6357)
	);

	bfr new_net_6358_bfr_after (
		.din(new_net_6357),
		.dout(new_net_6358)
	);

	bfr new_net_6359_bfr_after (
		.din(new_net_6358),
		.dout(new_net_6359)
	);

	bfr new_net_6360_bfr_after (
		.din(new_net_6359),
		.dout(new_net_6360)
	);

	bfr new_net_6361_bfr_after (
		.din(new_net_6360),
		.dout(new_net_6361)
	);

	bfr new_net_6362_bfr_after (
		.din(new_net_6361),
		.dout(new_net_6362)
	);

	bfr new_net_6363_bfr_after (
		.din(new_net_6362),
		.dout(new_net_6363)
	);

	bfr new_net_6364_bfr_after (
		.din(new_net_6363),
		.dout(new_net_6364)
	);

	bfr new_net_6365_bfr_after (
		.din(new_net_6364),
		.dout(new_net_6365)
	);

	bfr new_net_6366_bfr_after (
		.din(new_net_6365),
		.dout(new_net_6366)
	);

	bfr new_net_6367_bfr_after (
		.din(new_net_6366),
		.dout(new_net_6367)
	);

	bfr new_net_6368_bfr_after (
		.din(new_net_6367),
		.dout(new_net_6368)
	);

	bfr new_net_6369_bfr_after (
		.din(new_net_6368),
		.dout(new_net_6369)
	);

	bfr new_net_6370_bfr_after (
		.din(new_net_6369),
		.dout(new_net_6370)
	);

	bfr new_net_6371_bfr_after (
		.din(new_net_6370),
		.dout(new_net_6371)
	);

	bfr new_net_6372_bfr_after (
		.din(new_net_6371),
		.dout(new_net_6372)
	);

	bfr new_net_6373_bfr_after (
		.din(new_net_6372),
		.dout(new_net_6373)
	);

	bfr new_net_6374_bfr_after (
		.din(new_net_6373),
		.dout(new_net_6374)
	);

	spl2 _1571__v_fanout (
		.a(new_net_6374),
		.b(new_net_1708),
		.c(new_net_1709)
	);

	bfr new_net_6375_bfr_after (
		.din(_0884_),
		.dout(new_net_6375)
	);

	bfr new_net_6376_bfr_after (
		.din(new_net_6375),
		.dout(new_net_6376)
	);

	bfr new_net_6377_bfr_after (
		.din(new_net_6376),
		.dout(new_net_6377)
	);

	bfr new_net_6378_bfr_after (
		.din(new_net_6377),
		.dout(new_net_6378)
	);

	bfr new_net_6379_bfr_after (
		.din(new_net_6378),
		.dout(new_net_6379)
	);

	bfr new_net_6380_bfr_after (
		.din(new_net_6379),
		.dout(new_net_6380)
	);

	bfr new_net_6381_bfr_after (
		.din(new_net_6380),
		.dout(new_net_6381)
	);

	bfr new_net_6382_bfr_after (
		.din(new_net_6381),
		.dout(new_net_6382)
	);

	bfr new_net_6383_bfr_after (
		.din(new_net_6382),
		.dout(new_net_6383)
	);

	bfr new_net_6384_bfr_after (
		.din(new_net_6383),
		.dout(new_net_6384)
	);

	bfr new_net_6385_bfr_after (
		.din(new_net_6384),
		.dout(new_net_6385)
	);

	bfr new_net_6386_bfr_after (
		.din(new_net_6385),
		.dout(new_net_6386)
	);

	bfr new_net_6387_bfr_after (
		.din(new_net_6386),
		.dout(new_net_6387)
	);

	bfr new_net_6388_bfr_after (
		.din(new_net_6387),
		.dout(new_net_6388)
	);

	bfr new_net_6389_bfr_after (
		.din(new_net_6388),
		.dout(new_net_6389)
	);

	bfr new_net_6390_bfr_after (
		.din(new_net_6389),
		.dout(new_net_6390)
	);

	bfr new_net_6391_bfr_after (
		.din(new_net_6390),
		.dout(new_net_6391)
	);

	bfr new_net_6392_bfr_after (
		.din(new_net_6391),
		.dout(new_net_6392)
	);

	bfr new_net_6393_bfr_after (
		.din(new_net_6392),
		.dout(new_net_6393)
	);

	bfr new_net_6394_bfr_after (
		.din(new_net_6393),
		.dout(new_net_6394)
	);

	bfr new_net_6395_bfr_after (
		.din(new_net_6394),
		.dout(new_net_6395)
	);

	bfr new_net_6396_bfr_after (
		.din(new_net_6395),
		.dout(new_net_6396)
	);

	bfr new_net_6397_bfr_after (
		.din(new_net_6396),
		.dout(new_net_6397)
	);

	bfr new_net_6398_bfr_after (
		.din(new_net_6397),
		.dout(new_net_6398)
	);

	bfr new_net_6399_bfr_after (
		.din(new_net_6398),
		.dout(new_net_6399)
	);

	bfr new_net_6400_bfr_after (
		.din(new_net_6399),
		.dout(new_net_6400)
	);

	bfr new_net_6401_bfr_after (
		.din(new_net_6400),
		.dout(new_net_6401)
	);

	bfr new_net_6402_bfr_after (
		.din(new_net_6401),
		.dout(new_net_6402)
	);

	bfr new_net_6403_bfr_after (
		.din(new_net_6402),
		.dout(new_net_6403)
	);

	bfr new_net_6404_bfr_after (
		.din(new_net_6403),
		.dout(new_net_6404)
	);

	bfr new_net_6405_bfr_after (
		.din(new_net_6404),
		.dout(new_net_6405)
	);

	bfr new_net_6406_bfr_after (
		.din(new_net_6405),
		.dout(new_net_6406)
	);

	bfr new_net_6407_bfr_after (
		.din(new_net_6406),
		.dout(new_net_6407)
	);

	bfr new_net_6408_bfr_after (
		.din(new_net_6407),
		.dout(new_net_6408)
	);

	bfr new_net_6409_bfr_after (
		.din(new_net_6408),
		.dout(new_net_6409)
	);

	bfr new_net_6410_bfr_after (
		.din(new_net_6409),
		.dout(new_net_6410)
	);

	bfr new_net_6411_bfr_after (
		.din(new_net_6410),
		.dout(new_net_6411)
	);

	bfr new_net_6412_bfr_after (
		.din(new_net_6411),
		.dout(new_net_6412)
	);

	bfr new_net_6413_bfr_after (
		.din(new_net_6412),
		.dout(new_net_6413)
	);

	bfr new_net_6414_bfr_after (
		.din(new_net_6413),
		.dout(new_net_6414)
	);

	bfr new_net_6415_bfr_after (
		.din(new_net_6414),
		.dout(new_net_6415)
	);

	bfr new_net_6416_bfr_after (
		.din(new_net_6415),
		.dout(new_net_6416)
	);

	bfr new_net_6417_bfr_after (
		.din(new_net_6416),
		.dout(new_net_6417)
	);

	bfr new_net_6418_bfr_after (
		.din(new_net_6417),
		.dout(new_net_6418)
	);

	bfr new_net_6419_bfr_after (
		.din(new_net_6418),
		.dout(new_net_6419)
	);

	bfr new_net_6420_bfr_after (
		.din(new_net_6419),
		.dout(new_net_6420)
	);

	bfr new_net_6421_bfr_after (
		.din(new_net_6420),
		.dout(new_net_6421)
	);

	bfr new_net_6422_bfr_after (
		.din(new_net_6421),
		.dout(new_net_6422)
	);

	bfr new_net_6423_bfr_after (
		.din(new_net_6422),
		.dout(new_net_6423)
	);

	bfr new_net_6424_bfr_after (
		.din(new_net_6423),
		.dout(new_net_6424)
	);

	bfr new_net_6425_bfr_after (
		.din(new_net_6424),
		.dout(new_net_6425)
	);

	bfr new_net_6426_bfr_after (
		.din(new_net_6425),
		.dout(new_net_6426)
	);

	bfr new_net_6427_bfr_after (
		.din(new_net_6426),
		.dout(new_net_6427)
	);

	bfr new_net_6428_bfr_after (
		.din(new_net_6427),
		.dout(new_net_6428)
	);

	bfr new_net_6429_bfr_after (
		.din(new_net_6428),
		.dout(new_net_6429)
	);

	bfr new_net_6430_bfr_after (
		.din(new_net_6429),
		.dout(new_net_6430)
	);

	bfr new_net_6431_bfr_after (
		.din(new_net_6430),
		.dout(new_net_6431)
	);

	bfr new_net_6432_bfr_after (
		.din(new_net_6431),
		.dout(new_net_6432)
	);

	bfr new_net_6433_bfr_after (
		.din(new_net_6432),
		.dout(new_net_6433)
	);

	bfr new_net_6434_bfr_after (
		.din(new_net_6433),
		.dout(new_net_6434)
	);

	bfr new_net_6435_bfr_after (
		.din(new_net_6434),
		.dout(new_net_6435)
	);

	bfr new_net_6436_bfr_after (
		.din(new_net_6435),
		.dout(new_net_6436)
	);

	bfr new_net_6437_bfr_after (
		.din(new_net_6436),
		.dout(new_net_6437)
	);

	bfr new_net_6438_bfr_after (
		.din(new_net_6437),
		.dout(new_net_6438)
	);

	bfr new_net_6439_bfr_after (
		.din(new_net_6438),
		.dout(new_net_6439)
	);

	bfr new_net_6440_bfr_after (
		.din(new_net_6439),
		.dout(new_net_6440)
	);

	bfr new_net_6441_bfr_after (
		.din(new_net_6440),
		.dout(new_net_6441)
	);

	bfr new_net_6442_bfr_after (
		.din(new_net_6441),
		.dout(new_net_6442)
	);

	bfr new_net_6443_bfr_after (
		.din(new_net_6442),
		.dout(new_net_6443)
	);

	bfr new_net_6444_bfr_after (
		.din(new_net_6443),
		.dout(new_net_6444)
	);

	bfr new_net_6445_bfr_after (
		.din(new_net_6444),
		.dout(new_net_6445)
	);

	bfr new_net_6446_bfr_after (
		.din(new_net_6445),
		.dout(new_net_6446)
	);

	bfr new_net_6447_bfr_after (
		.din(new_net_6446),
		.dout(new_net_6447)
	);

	bfr new_net_6448_bfr_after (
		.din(new_net_6447),
		.dout(new_net_6448)
	);

	bfr new_net_6449_bfr_after (
		.din(new_net_6448),
		.dout(new_net_6449)
	);

	bfr new_net_6450_bfr_after (
		.din(new_net_6449),
		.dout(new_net_6450)
	);

	bfr new_net_6451_bfr_after (
		.din(new_net_6450),
		.dout(new_net_6451)
	);

	bfr new_net_6452_bfr_after (
		.din(new_net_6451),
		.dout(new_net_6452)
	);

	bfr new_net_6453_bfr_after (
		.din(new_net_6452),
		.dout(new_net_6453)
	);

	bfr new_net_6454_bfr_after (
		.din(new_net_6453),
		.dout(new_net_6454)
	);

	bfr new_net_6455_bfr_after (
		.din(new_net_6454),
		.dout(new_net_6455)
	);

	bfr new_net_6456_bfr_after (
		.din(new_net_6455),
		.dout(new_net_6456)
	);

	bfr new_net_6457_bfr_after (
		.din(new_net_6456),
		.dout(new_net_6457)
	);

	bfr new_net_6458_bfr_after (
		.din(new_net_6457),
		.dout(new_net_6458)
	);

	bfr new_net_6459_bfr_after (
		.din(new_net_6458),
		.dout(new_net_6459)
	);

	bfr new_net_6460_bfr_after (
		.din(new_net_6459),
		.dout(new_net_6460)
	);

	bfr new_net_6461_bfr_after (
		.din(new_net_6460),
		.dout(new_net_6461)
	);

	bfr new_net_6462_bfr_after (
		.din(new_net_6461),
		.dout(new_net_6462)
	);

	bfr new_net_6463_bfr_after (
		.din(new_net_6462),
		.dout(new_net_6463)
	);

	bfr new_net_6464_bfr_after (
		.din(new_net_6463),
		.dout(new_net_6464)
	);

	bfr new_net_6465_bfr_after (
		.din(new_net_6464),
		.dout(new_net_6465)
	);

	bfr new_net_6466_bfr_after (
		.din(new_net_6465),
		.dout(new_net_6466)
	);

	bfr new_net_6467_bfr_after (
		.din(new_net_6466),
		.dout(new_net_6467)
	);

	bfr new_net_6468_bfr_after (
		.din(new_net_6467),
		.dout(new_net_6468)
	);

	bfr new_net_6469_bfr_after (
		.din(new_net_6468),
		.dout(new_net_6469)
	);

	bfr new_net_6470_bfr_after (
		.din(new_net_6469),
		.dout(new_net_6470)
	);

	bfr new_net_6471_bfr_after (
		.din(new_net_6470),
		.dout(new_net_6471)
	);

	bfr new_net_6472_bfr_after (
		.din(new_net_6471),
		.dout(new_net_6472)
	);

	bfr new_net_6473_bfr_after (
		.din(new_net_6472),
		.dout(new_net_6473)
	);

	bfr new_net_6474_bfr_after (
		.din(new_net_6473),
		.dout(new_net_6474)
	);

	bfr new_net_6475_bfr_after (
		.din(new_net_6474),
		.dout(new_net_6475)
	);

	bfr new_net_6476_bfr_after (
		.din(new_net_6475),
		.dout(new_net_6476)
	);

	bfr new_net_6477_bfr_after (
		.din(new_net_6476),
		.dout(new_net_6477)
	);

	bfr new_net_6478_bfr_after (
		.din(new_net_6477),
		.dout(new_net_6478)
	);

	spl2 _0884__v_fanout (
		.a(new_net_6478),
		.b(new_net_2750),
		.c(new_net_2751)
	);

	bfr new_net_6479_bfr_after (
		.din(_1134_),
		.dout(new_net_6479)
	);

	bfr new_net_6480_bfr_after (
		.din(new_net_6479),
		.dout(new_net_6480)
	);

	bfr new_net_6481_bfr_after (
		.din(new_net_6480),
		.dout(new_net_6481)
	);

	bfr new_net_6482_bfr_after (
		.din(new_net_6481),
		.dout(new_net_6482)
	);

	bfr new_net_6483_bfr_after (
		.din(new_net_6482),
		.dout(new_net_6483)
	);

	bfr new_net_6484_bfr_after (
		.din(new_net_6483),
		.dout(new_net_6484)
	);

	bfr new_net_6485_bfr_after (
		.din(new_net_6484),
		.dout(new_net_6485)
	);

	bfr new_net_6486_bfr_after (
		.din(new_net_6485),
		.dout(new_net_6486)
	);

	bfr new_net_6487_bfr_after (
		.din(new_net_6486),
		.dout(new_net_6487)
	);

	bfr new_net_6488_bfr_after (
		.din(new_net_6487),
		.dout(new_net_6488)
	);

	bfr new_net_6489_bfr_after (
		.din(new_net_6488),
		.dout(new_net_6489)
	);

	bfr new_net_6490_bfr_after (
		.din(new_net_6489),
		.dout(new_net_6490)
	);

	bfr new_net_6491_bfr_after (
		.din(new_net_6490),
		.dout(new_net_6491)
	);

	bfr new_net_6492_bfr_after (
		.din(new_net_6491),
		.dout(new_net_6492)
	);

	bfr new_net_6493_bfr_after (
		.din(new_net_6492),
		.dout(new_net_6493)
	);

	bfr new_net_6494_bfr_after (
		.din(new_net_6493),
		.dout(new_net_6494)
	);

	bfr new_net_6495_bfr_after (
		.din(new_net_6494),
		.dout(new_net_6495)
	);

	bfr new_net_6496_bfr_after (
		.din(new_net_6495),
		.dout(new_net_6496)
	);

	bfr new_net_6497_bfr_after (
		.din(new_net_6496),
		.dout(new_net_6497)
	);

	bfr new_net_6498_bfr_after (
		.din(new_net_6497),
		.dout(new_net_6498)
	);

	bfr new_net_6499_bfr_after (
		.din(new_net_6498),
		.dout(new_net_6499)
	);

	bfr new_net_6500_bfr_after (
		.din(new_net_6499),
		.dout(new_net_6500)
	);

	bfr new_net_6501_bfr_after (
		.din(new_net_6500),
		.dout(new_net_6501)
	);

	bfr new_net_6502_bfr_after (
		.din(new_net_6501),
		.dout(new_net_6502)
	);

	bfr new_net_6503_bfr_after (
		.din(new_net_6502),
		.dout(new_net_6503)
	);

	bfr new_net_6504_bfr_after (
		.din(new_net_6503),
		.dout(new_net_6504)
	);

	bfr new_net_6505_bfr_after (
		.din(new_net_6504),
		.dout(new_net_6505)
	);

	bfr new_net_6506_bfr_after (
		.din(new_net_6505),
		.dout(new_net_6506)
	);

	bfr new_net_6507_bfr_after (
		.din(new_net_6506),
		.dout(new_net_6507)
	);

	bfr new_net_6508_bfr_after (
		.din(new_net_6507),
		.dout(new_net_6508)
	);

	bfr new_net_6509_bfr_after (
		.din(new_net_6508),
		.dout(new_net_6509)
	);

	bfr new_net_6510_bfr_after (
		.din(new_net_6509),
		.dout(new_net_6510)
	);

	bfr new_net_6511_bfr_after (
		.din(new_net_6510),
		.dout(new_net_6511)
	);

	bfr new_net_6512_bfr_after (
		.din(new_net_6511),
		.dout(new_net_6512)
	);

	bfr new_net_6513_bfr_after (
		.din(new_net_6512),
		.dout(new_net_6513)
	);

	bfr new_net_6514_bfr_after (
		.din(new_net_6513),
		.dout(new_net_6514)
	);

	bfr new_net_6515_bfr_after (
		.din(new_net_6514),
		.dout(new_net_6515)
	);

	bfr new_net_6516_bfr_after (
		.din(new_net_6515),
		.dout(new_net_6516)
	);

	bfr new_net_6517_bfr_after (
		.din(new_net_6516),
		.dout(new_net_6517)
	);

	bfr new_net_6518_bfr_after (
		.din(new_net_6517),
		.dout(new_net_6518)
	);

	spl2 _1134__v_fanout (
		.a(new_net_6518),
		.b(new_net_681),
		.c(new_net_682)
	);

	bfr new_net_6519_bfr_after (
		.din(_1217_),
		.dout(new_net_6519)
	);

	bfr new_net_6520_bfr_after (
		.din(new_net_6519),
		.dout(new_net_6520)
	);

	bfr new_net_6521_bfr_after (
		.din(new_net_6520),
		.dout(new_net_6521)
	);

	bfr new_net_6522_bfr_after (
		.din(new_net_6521),
		.dout(new_net_6522)
	);

	bfr new_net_6523_bfr_after (
		.din(new_net_6522),
		.dout(new_net_6523)
	);

	bfr new_net_6524_bfr_after (
		.din(new_net_6523),
		.dout(new_net_6524)
	);

	bfr new_net_6525_bfr_after (
		.din(new_net_6524),
		.dout(new_net_6525)
	);

	bfr new_net_6526_bfr_after (
		.din(new_net_6525),
		.dout(new_net_6526)
	);

	bfr new_net_6527_bfr_after (
		.din(new_net_6526),
		.dout(new_net_6527)
	);

	bfr new_net_6528_bfr_after (
		.din(new_net_6527),
		.dout(new_net_6528)
	);

	bfr new_net_6529_bfr_after (
		.din(new_net_6528),
		.dout(new_net_6529)
	);

	bfr new_net_6530_bfr_after (
		.din(new_net_6529),
		.dout(new_net_6530)
	);

	bfr new_net_6531_bfr_after (
		.din(new_net_6530),
		.dout(new_net_6531)
	);

	bfr new_net_6532_bfr_after (
		.din(new_net_6531),
		.dout(new_net_6532)
	);

	bfr new_net_6533_bfr_after (
		.din(new_net_6532),
		.dout(new_net_6533)
	);

	bfr new_net_6534_bfr_after (
		.din(new_net_6533),
		.dout(new_net_6534)
	);

	spl2 _1217__v_fanout (
		.a(new_net_6534),
		.b(new_net_1016),
		.c(new_net_1017)
	);

	bfr new_net_6535_bfr_after (
		.din(_1456_),
		.dout(new_net_6535)
	);

	bfr new_net_6536_bfr_after (
		.din(new_net_6535),
		.dout(new_net_6536)
	);

	bfr new_net_6537_bfr_after (
		.din(new_net_6536),
		.dout(new_net_6537)
	);

	bfr new_net_6538_bfr_after (
		.din(new_net_6537),
		.dout(new_net_6538)
	);

	bfr new_net_6539_bfr_after (
		.din(new_net_6538),
		.dout(new_net_6539)
	);

	bfr new_net_6540_bfr_after (
		.din(new_net_6539),
		.dout(new_net_6540)
	);

	bfr new_net_6541_bfr_after (
		.din(new_net_6540),
		.dout(new_net_6541)
	);

	bfr new_net_6542_bfr_after (
		.din(new_net_6541),
		.dout(new_net_6542)
	);

	bfr new_net_6543_bfr_after (
		.din(new_net_6542),
		.dout(new_net_6543)
	);

	bfr new_net_6544_bfr_after (
		.din(new_net_6543),
		.dout(new_net_6544)
	);

	bfr new_net_6545_bfr_after (
		.din(new_net_6544),
		.dout(new_net_6545)
	);

	bfr new_net_6546_bfr_after (
		.din(new_net_6545),
		.dout(new_net_6546)
	);

	bfr new_net_6547_bfr_after (
		.din(new_net_6546),
		.dout(new_net_6547)
	);

	bfr new_net_6548_bfr_after (
		.din(new_net_6547),
		.dout(new_net_6548)
	);

	bfr new_net_6549_bfr_after (
		.din(new_net_6548),
		.dout(new_net_6549)
	);

	bfr new_net_6550_bfr_after (
		.din(new_net_6549),
		.dout(new_net_6550)
	);

	bfr new_net_6551_bfr_after (
		.din(new_net_6550),
		.dout(new_net_6551)
	);

	bfr new_net_6552_bfr_after (
		.din(new_net_6551),
		.dout(new_net_6552)
	);

	bfr new_net_6553_bfr_after (
		.din(new_net_6552),
		.dout(new_net_6553)
	);

	bfr new_net_6554_bfr_after (
		.din(new_net_6553),
		.dout(new_net_6554)
	);

	bfr new_net_6555_bfr_after (
		.din(new_net_6554),
		.dout(new_net_6555)
	);

	bfr new_net_6556_bfr_after (
		.din(new_net_6555),
		.dout(new_net_6556)
	);

	bfr new_net_6557_bfr_after (
		.din(new_net_6556),
		.dout(new_net_6557)
	);

	bfr new_net_6558_bfr_after (
		.din(new_net_6557),
		.dout(new_net_6558)
	);

	bfr new_net_6559_bfr_after (
		.din(new_net_6558),
		.dout(new_net_6559)
	);

	bfr new_net_6560_bfr_after (
		.din(new_net_6559),
		.dout(new_net_6560)
	);

	bfr new_net_6561_bfr_after (
		.din(new_net_6560),
		.dout(new_net_6561)
	);

	bfr new_net_6562_bfr_after (
		.din(new_net_6561),
		.dout(new_net_6562)
	);

	bfr new_net_6563_bfr_after (
		.din(new_net_6562),
		.dout(new_net_6563)
	);

	bfr new_net_6564_bfr_after (
		.din(new_net_6563),
		.dout(new_net_6564)
	);

	bfr new_net_6565_bfr_after (
		.din(new_net_6564),
		.dout(new_net_6565)
	);

	bfr new_net_6566_bfr_after (
		.din(new_net_6565),
		.dout(new_net_6566)
	);

	bfr new_net_6567_bfr_after (
		.din(new_net_6566),
		.dout(new_net_6567)
	);

	bfr new_net_6568_bfr_after (
		.din(new_net_6567),
		.dout(new_net_6568)
	);

	bfr new_net_6569_bfr_after (
		.din(new_net_6568),
		.dout(new_net_6569)
	);

	bfr new_net_6570_bfr_after (
		.din(new_net_6569),
		.dout(new_net_6570)
	);

	bfr new_net_6571_bfr_after (
		.din(new_net_6570),
		.dout(new_net_6571)
	);

	bfr new_net_6572_bfr_after (
		.din(new_net_6571),
		.dout(new_net_6572)
	);

	bfr new_net_6573_bfr_after (
		.din(new_net_6572),
		.dout(new_net_6573)
	);

	bfr new_net_6574_bfr_after (
		.din(new_net_6573),
		.dout(new_net_6574)
	);

	bfr new_net_6575_bfr_after (
		.din(new_net_6574),
		.dout(new_net_6575)
	);

	bfr new_net_6576_bfr_after (
		.din(new_net_6575),
		.dout(new_net_6576)
	);

	bfr new_net_6577_bfr_after (
		.din(new_net_6576),
		.dout(new_net_6577)
	);

	bfr new_net_6578_bfr_after (
		.din(new_net_6577),
		.dout(new_net_6578)
	);

	bfr new_net_6579_bfr_after (
		.din(new_net_6578),
		.dout(new_net_6579)
	);

	bfr new_net_6580_bfr_after (
		.din(new_net_6579),
		.dout(new_net_6580)
	);

	bfr new_net_6581_bfr_after (
		.din(new_net_6580),
		.dout(new_net_6581)
	);

	bfr new_net_6582_bfr_after (
		.din(new_net_6581),
		.dout(new_net_6582)
	);

	bfr new_net_6583_bfr_after (
		.din(new_net_6582),
		.dout(new_net_6583)
	);

	bfr new_net_6584_bfr_after (
		.din(new_net_6583),
		.dout(new_net_6584)
	);

	bfr new_net_6585_bfr_after (
		.din(new_net_6584),
		.dout(new_net_6585)
	);

	bfr new_net_6586_bfr_after (
		.din(new_net_6585),
		.dout(new_net_6586)
	);

	bfr new_net_6587_bfr_after (
		.din(new_net_6586),
		.dout(new_net_6587)
	);

	bfr new_net_6588_bfr_after (
		.din(new_net_6587),
		.dout(new_net_6588)
	);

	bfr new_net_6589_bfr_after (
		.din(new_net_6588),
		.dout(new_net_6589)
	);

	bfr new_net_6590_bfr_after (
		.din(new_net_6589),
		.dout(new_net_6590)
	);

	bfr new_net_6591_bfr_after (
		.din(new_net_6590),
		.dout(new_net_6591)
	);

	bfr new_net_6592_bfr_after (
		.din(new_net_6591),
		.dout(new_net_6592)
	);

	bfr new_net_6593_bfr_after (
		.din(new_net_6592),
		.dout(new_net_6593)
	);

	bfr new_net_6594_bfr_after (
		.din(new_net_6593),
		.dout(new_net_6594)
	);

	bfr new_net_6595_bfr_after (
		.din(new_net_6594),
		.dout(new_net_6595)
	);

	bfr new_net_6596_bfr_after (
		.din(new_net_6595),
		.dout(new_net_6596)
	);

	bfr new_net_6597_bfr_after (
		.din(new_net_6596),
		.dout(new_net_6597)
	);

	bfr new_net_6598_bfr_after (
		.din(new_net_6597),
		.dout(new_net_6598)
	);

	bfr new_net_6599_bfr_after (
		.din(new_net_6598),
		.dout(new_net_6599)
	);

	bfr new_net_6600_bfr_after (
		.din(new_net_6599),
		.dout(new_net_6600)
	);

	bfr new_net_6601_bfr_after (
		.din(new_net_6600),
		.dout(new_net_6601)
	);

	bfr new_net_6602_bfr_after (
		.din(new_net_6601),
		.dout(new_net_6602)
	);

	bfr new_net_6603_bfr_after (
		.din(new_net_6602),
		.dout(new_net_6603)
	);

	bfr new_net_6604_bfr_after (
		.din(new_net_6603),
		.dout(new_net_6604)
	);

	bfr new_net_6605_bfr_after (
		.din(new_net_6604),
		.dout(new_net_6605)
	);

	bfr new_net_6606_bfr_after (
		.din(new_net_6605),
		.dout(new_net_6606)
	);

	bfr new_net_6607_bfr_after (
		.din(new_net_6606),
		.dout(new_net_6607)
	);

	bfr new_net_6608_bfr_after (
		.din(new_net_6607),
		.dout(new_net_6608)
	);

	bfr new_net_6609_bfr_after (
		.din(new_net_6608),
		.dout(new_net_6609)
	);

	bfr new_net_6610_bfr_after (
		.din(new_net_6609),
		.dout(new_net_6610)
	);

	bfr new_net_6611_bfr_after (
		.din(new_net_6610),
		.dout(new_net_6611)
	);

	bfr new_net_6612_bfr_after (
		.din(new_net_6611),
		.dout(new_net_6612)
	);

	bfr new_net_6613_bfr_after (
		.din(new_net_6612),
		.dout(new_net_6613)
	);

	bfr new_net_6614_bfr_after (
		.din(new_net_6613),
		.dout(new_net_6614)
	);

	spl2 _1456__v_fanout (
		.a(new_net_6614),
		.b(new_net_2210),
		.c(new_net_2211)
	);

	bfr new_net_6615_bfr_after (
		.din(_0111_),
		.dout(new_net_6615)
	);

	bfr new_net_6616_bfr_after (
		.din(new_net_6615),
		.dout(new_net_6616)
	);

	bfr new_net_6617_bfr_after (
		.din(new_net_6616),
		.dout(new_net_6617)
	);

	bfr new_net_6618_bfr_after (
		.din(new_net_6617),
		.dout(new_net_6618)
	);

	bfr new_net_6619_bfr_after (
		.din(new_net_6618),
		.dout(new_net_6619)
	);

	bfr new_net_6620_bfr_after (
		.din(new_net_6619),
		.dout(new_net_6620)
	);

	bfr new_net_6621_bfr_after (
		.din(new_net_6620),
		.dout(new_net_6621)
	);

	bfr new_net_6622_bfr_after (
		.din(new_net_6621),
		.dout(new_net_6622)
	);

	bfr new_net_6623_bfr_after (
		.din(new_net_6622),
		.dout(new_net_6623)
	);

	bfr new_net_6624_bfr_after (
		.din(new_net_6623),
		.dout(new_net_6624)
	);

	spl2 _0111__v_fanout (
		.a(new_net_6624),
		.b(new_net_2791),
		.c(new_net_2792)
	);

	bfr new_net_6625_bfr_after (
		.din(_0886_),
		.dout(new_net_6625)
	);

	bfr new_net_6626_bfr_after (
		.din(new_net_6625),
		.dout(new_net_6626)
	);

	bfr new_net_6627_bfr_after (
		.din(new_net_6626),
		.dout(new_net_6627)
	);

	bfr new_net_6628_bfr_after (
		.din(new_net_6627),
		.dout(new_net_6628)
	);

	bfr new_net_6629_bfr_after (
		.din(new_net_6628),
		.dout(new_net_6629)
	);

	bfr new_net_6630_bfr_after (
		.din(new_net_6629),
		.dout(new_net_6630)
	);

	bfr new_net_6631_bfr_after (
		.din(new_net_6630),
		.dout(new_net_6631)
	);

	bfr new_net_6632_bfr_after (
		.din(new_net_6631),
		.dout(new_net_6632)
	);

	bfr new_net_6633_bfr_after (
		.din(new_net_6632),
		.dout(new_net_6633)
	);

	bfr new_net_6634_bfr_after (
		.din(new_net_6633),
		.dout(new_net_6634)
	);

	bfr new_net_6635_bfr_after (
		.din(new_net_6634),
		.dout(new_net_6635)
	);

	bfr new_net_6636_bfr_after (
		.din(new_net_6635),
		.dout(new_net_6636)
	);

	bfr new_net_6637_bfr_after (
		.din(new_net_6636),
		.dout(new_net_6637)
	);

	bfr new_net_6638_bfr_after (
		.din(new_net_6637),
		.dout(new_net_6638)
	);

	bfr new_net_6639_bfr_after (
		.din(new_net_6638),
		.dout(new_net_6639)
	);

	bfr new_net_6640_bfr_after (
		.din(new_net_6639),
		.dout(new_net_6640)
	);

	bfr new_net_6641_bfr_after (
		.din(new_net_6640),
		.dout(new_net_6641)
	);

	bfr new_net_6642_bfr_after (
		.din(new_net_6641),
		.dout(new_net_6642)
	);

	bfr new_net_6643_bfr_after (
		.din(new_net_6642),
		.dout(new_net_6643)
	);

	bfr new_net_6644_bfr_after (
		.din(new_net_6643),
		.dout(new_net_6644)
	);

	bfr new_net_6645_bfr_after (
		.din(new_net_6644),
		.dout(new_net_6645)
	);

	bfr new_net_6646_bfr_after (
		.din(new_net_6645),
		.dout(new_net_6646)
	);

	bfr new_net_6647_bfr_after (
		.din(new_net_6646),
		.dout(new_net_6647)
	);

	bfr new_net_6648_bfr_after (
		.din(new_net_6647),
		.dout(new_net_6648)
	);

	bfr new_net_6649_bfr_after (
		.din(new_net_6648),
		.dout(new_net_6649)
	);

	bfr new_net_6650_bfr_after (
		.din(new_net_6649),
		.dout(new_net_6650)
	);

	bfr new_net_6651_bfr_after (
		.din(new_net_6650),
		.dout(new_net_6651)
	);

	bfr new_net_6652_bfr_after (
		.din(new_net_6651),
		.dout(new_net_6652)
	);

	bfr new_net_6653_bfr_after (
		.din(new_net_6652),
		.dout(new_net_6653)
	);

	bfr new_net_6654_bfr_after (
		.din(new_net_6653),
		.dout(new_net_6654)
	);

	bfr new_net_6655_bfr_after (
		.din(new_net_6654),
		.dout(new_net_6655)
	);

	bfr new_net_6656_bfr_after (
		.din(new_net_6655),
		.dout(new_net_6656)
	);

	bfr new_net_6657_bfr_after (
		.din(new_net_6656),
		.dout(new_net_6657)
	);

	bfr new_net_6658_bfr_after (
		.din(new_net_6657),
		.dout(new_net_6658)
	);

	bfr new_net_6659_bfr_after (
		.din(new_net_6658),
		.dout(new_net_6659)
	);

	bfr new_net_6660_bfr_after (
		.din(new_net_6659),
		.dout(new_net_6660)
	);

	bfr new_net_6661_bfr_after (
		.din(new_net_6660),
		.dout(new_net_6661)
	);

	bfr new_net_6662_bfr_after (
		.din(new_net_6661),
		.dout(new_net_6662)
	);

	bfr new_net_6663_bfr_after (
		.din(new_net_6662),
		.dout(new_net_6663)
	);

	bfr new_net_6664_bfr_after (
		.din(new_net_6663),
		.dout(new_net_6664)
	);

	bfr new_net_6665_bfr_after (
		.din(new_net_6664),
		.dout(new_net_6665)
	);

	bfr new_net_6666_bfr_after (
		.din(new_net_6665),
		.dout(new_net_6666)
	);

	bfr new_net_6667_bfr_after (
		.din(new_net_6666),
		.dout(new_net_6667)
	);

	bfr new_net_6668_bfr_after (
		.din(new_net_6667),
		.dout(new_net_6668)
	);

	bfr new_net_6669_bfr_after (
		.din(new_net_6668),
		.dout(new_net_6669)
	);

	bfr new_net_6670_bfr_after (
		.din(new_net_6669),
		.dout(new_net_6670)
	);

	bfr new_net_6671_bfr_after (
		.din(new_net_6670),
		.dout(new_net_6671)
	);

	bfr new_net_6672_bfr_after (
		.din(new_net_6671),
		.dout(new_net_6672)
	);

	bfr new_net_6673_bfr_after (
		.din(new_net_6672),
		.dout(new_net_6673)
	);

	bfr new_net_6674_bfr_after (
		.din(new_net_6673),
		.dout(new_net_6674)
	);

	bfr new_net_6675_bfr_after (
		.din(new_net_6674),
		.dout(new_net_6675)
	);

	bfr new_net_6676_bfr_after (
		.din(new_net_6675),
		.dout(new_net_6676)
	);

	bfr new_net_6677_bfr_after (
		.din(new_net_6676),
		.dout(new_net_6677)
	);

	bfr new_net_6678_bfr_after (
		.din(new_net_6677),
		.dout(new_net_6678)
	);

	bfr new_net_6679_bfr_after (
		.din(new_net_6678),
		.dout(new_net_6679)
	);

	bfr new_net_6680_bfr_after (
		.din(new_net_6679),
		.dout(new_net_6680)
	);

	bfr new_net_6681_bfr_after (
		.din(new_net_6680),
		.dout(new_net_6681)
	);

	bfr new_net_6682_bfr_after (
		.din(new_net_6681),
		.dout(new_net_6682)
	);

	bfr new_net_6683_bfr_after (
		.din(new_net_6682),
		.dout(new_net_6683)
	);

	bfr new_net_6684_bfr_after (
		.din(new_net_6683),
		.dout(new_net_6684)
	);

	bfr new_net_6685_bfr_after (
		.din(new_net_6684),
		.dout(new_net_6685)
	);

	bfr new_net_6686_bfr_after (
		.din(new_net_6685),
		.dout(new_net_6686)
	);

	bfr new_net_6687_bfr_after (
		.din(new_net_6686),
		.dout(new_net_6687)
	);

	bfr new_net_6688_bfr_after (
		.din(new_net_6687),
		.dout(new_net_6688)
	);

	bfr new_net_6689_bfr_after (
		.din(new_net_6688),
		.dout(new_net_6689)
	);

	bfr new_net_6690_bfr_after (
		.din(new_net_6689),
		.dout(new_net_6690)
	);

	bfr new_net_6691_bfr_after (
		.din(new_net_6690),
		.dout(new_net_6691)
	);

	bfr new_net_6692_bfr_after (
		.din(new_net_6691),
		.dout(new_net_6692)
	);

	bfr new_net_6693_bfr_after (
		.din(new_net_6692),
		.dout(new_net_6693)
	);

	bfr new_net_6694_bfr_after (
		.din(new_net_6693),
		.dout(new_net_6694)
	);

	bfr new_net_6695_bfr_after (
		.din(new_net_6694),
		.dout(new_net_6695)
	);

	bfr new_net_6696_bfr_after (
		.din(new_net_6695),
		.dout(new_net_6696)
	);

	bfr new_net_6697_bfr_after (
		.din(new_net_6696),
		.dout(new_net_6697)
	);

	bfr new_net_6698_bfr_after (
		.din(new_net_6697),
		.dout(new_net_6698)
	);

	bfr new_net_6699_bfr_after (
		.din(new_net_6698),
		.dout(new_net_6699)
	);

	bfr new_net_6700_bfr_after (
		.din(new_net_6699),
		.dout(new_net_6700)
	);

	bfr new_net_6701_bfr_after (
		.din(new_net_6700),
		.dout(new_net_6701)
	);

	bfr new_net_6702_bfr_after (
		.din(new_net_6701),
		.dout(new_net_6702)
	);

	bfr new_net_6703_bfr_after (
		.din(new_net_6702),
		.dout(new_net_6703)
	);

	bfr new_net_6704_bfr_after (
		.din(new_net_6703),
		.dout(new_net_6704)
	);

	bfr new_net_6705_bfr_after (
		.din(new_net_6704),
		.dout(new_net_6705)
	);

	bfr new_net_6706_bfr_after (
		.din(new_net_6705),
		.dout(new_net_6706)
	);

	bfr new_net_6707_bfr_after (
		.din(new_net_6706),
		.dout(new_net_6707)
	);

	bfr new_net_6708_bfr_after (
		.din(new_net_6707),
		.dout(new_net_6708)
	);

	bfr new_net_6709_bfr_after (
		.din(new_net_6708),
		.dout(new_net_6709)
	);

	bfr new_net_6710_bfr_after (
		.din(new_net_6709),
		.dout(new_net_6710)
	);

	bfr new_net_6711_bfr_after (
		.din(new_net_6710),
		.dout(new_net_6711)
	);

	bfr new_net_6712_bfr_after (
		.din(new_net_6711),
		.dout(new_net_6712)
	);

	bfr new_net_6713_bfr_after (
		.din(new_net_6712),
		.dout(new_net_6713)
	);

	bfr new_net_6714_bfr_after (
		.din(new_net_6713),
		.dout(new_net_6714)
	);

	bfr new_net_6715_bfr_after (
		.din(new_net_6714),
		.dout(new_net_6715)
	);

	bfr new_net_6716_bfr_after (
		.din(new_net_6715),
		.dout(new_net_6716)
	);

	bfr new_net_6717_bfr_after (
		.din(new_net_6716),
		.dout(new_net_6717)
	);

	bfr new_net_6718_bfr_after (
		.din(new_net_6717),
		.dout(new_net_6718)
	);

	spl2 _0886__v_fanout (
		.a(new_net_6718),
		.b(new_net_2813),
		.c(new_net_2814)
	);

	spl2 _1382__v_fanout (
		.a(_1382_),
		.b(new_net_582),
		.c(new_net_583)
	);

	bfr new_net_6719_bfr_after (
		.din(_1379_),
		.dout(new_net_6719)
	);

	bfr new_net_6720_bfr_after (
		.din(new_net_6719),
		.dout(new_net_6720)
	);

	bfr new_net_6721_bfr_after (
		.din(new_net_6720),
		.dout(new_net_6721)
	);

	bfr new_net_6722_bfr_after (
		.din(new_net_6721),
		.dout(new_net_6722)
	);

	bfr new_net_6723_bfr_after (
		.din(new_net_6722),
		.dout(new_net_6723)
	);

	bfr new_net_6724_bfr_after (
		.din(new_net_6723),
		.dout(new_net_6724)
	);

	bfr new_net_6725_bfr_after (
		.din(new_net_6724),
		.dout(new_net_6725)
	);

	bfr new_net_6726_bfr_after (
		.din(new_net_6725),
		.dout(new_net_6726)
	);

	bfr new_net_6727_bfr_after (
		.din(new_net_6726),
		.dout(new_net_6727)
	);

	bfr new_net_6728_bfr_after (
		.din(new_net_6727),
		.dout(new_net_6728)
	);

	bfr new_net_6729_bfr_after (
		.din(new_net_6728),
		.dout(new_net_6729)
	);

	bfr new_net_6730_bfr_after (
		.din(new_net_6729),
		.dout(new_net_6730)
	);

	bfr new_net_6731_bfr_after (
		.din(new_net_6730),
		.dout(new_net_6731)
	);

	bfr new_net_6732_bfr_after (
		.din(new_net_6731),
		.dout(new_net_6732)
	);

	bfr new_net_6733_bfr_after (
		.din(new_net_6732),
		.dout(new_net_6733)
	);

	bfr new_net_6734_bfr_after (
		.din(new_net_6733),
		.dout(new_net_6734)
	);

	spl2 _1379__v_fanout (
		.a(new_net_6734),
		.b(new_net_14),
		.c(new_net_15)
	);

	bfr new_net_6735_bfr_after (
		.din(_0447_),
		.dout(new_net_6735)
	);

	bfr new_net_6736_bfr_after (
		.din(new_net_6735),
		.dout(new_net_6736)
	);

	bfr new_net_6737_bfr_after (
		.din(new_net_6736),
		.dout(new_net_6737)
	);

	bfr new_net_6738_bfr_after (
		.din(new_net_6737),
		.dout(new_net_6738)
	);

	bfr new_net_6739_bfr_after (
		.din(new_net_6738),
		.dout(new_net_6739)
	);

	bfr new_net_6740_bfr_after (
		.din(new_net_6739),
		.dout(new_net_6740)
	);

	bfr new_net_6741_bfr_after (
		.din(new_net_6740),
		.dout(new_net_6741)
	);

	bfr new_net_6742_bfr_after (
		.din(new_net_6741),
		.dout(new_net_6742)
	);

	bfr new_net_6743_bfr_after (
		.din(new_net_6742),
		.dout(new_net_6743)
	);

	bfr new_net_6744_bfr_after (
		.din(new_net_6743),
		.dout(new_net_6744)
	);

	bfr new_net_6745_bfr_after (
		.din(new_net_6744),
		.dout(new_net_6745)
	);

	bfr new_net_6746_bfr_after (
		.din(new_net_6745),
		.dout(new_net_6746)
	);

	bfr new_net_6747_bfr_after (
		.din(new_net_6746),
		.dout(new_net_6747)
	);

	bfr new_net_6748_bfr_after (
		.din(new_net_6747),
		.dout(new_net_6748)
	);

	bfr new_net_6749_bfr_after (
		.din(new_net_6748),
		.dout(new_net_6749)
	);

	bfr new_net_6750_bfr_after (
		.din(new_net_6749),
		.dout(new_net_6750)
	);

	bfr new_net_6751_bfr_after (
		.din(new_net_6750),
		.dout(new_net_6751)
	);

	bfr new_net_6752_bfr_after (
		.din(new_net_6751),
		.dout(new_net_6752)
	);

	bfr new_net_6753_bfr_after (
		.din(new_net_6752),
		.dout(new_net_6753)
	);

	bfr new_net_6754_bfr_after (
		.din(new_net_6753),
		.dout(new_net_6754)
	);

	bfr new_net_6755_bfr_after (
		.din(new_net_6754),
		.dout(new_net_6755)
	);

	bfr new_net_6756_bfr_after (
		.din(new_net_6755),
		.dout(new_net_6756)
	);

	bfr new_net_6757_bfr_after (
		.din(new_net_6756),
		.dout(new_net_6757)
	);

	bfr new_net_6758_bfr_after (
		.din(new_net_6757),
		.dout(new_net_6758)
	);

	bfr new_net_6759_bfr_after (
		.din(new_net_6758),
		.dout(new_net_6759)
	);

	bfr new_net_6760_bfr_after (
		.din(new_net_6759),
		.dout(new_net_6760)
	);

	bfr new_net_6761_bfr_after (
		.din(new_net_6760),
		.dout(new_net_6761)
	);

	bfr new_net_6762_bfr_after (
		.din(new_net_6761),
		.dout(new_net_6762)
	);

	bfr new_net_6763_bfr_after (
		.din(new_net_6762),
		.dout(new_net_6763)
	);

	bfr new_net_6764_bfr_after (
		.din(new_net_6763),
		.dout(new_net_6764)
	);

	bfr new_net_6765_bfr_after (
		.din(new_net_6764),
		.dout(new_net_6765)
	);

	bfr new_net_6766_bfr_after (
		.din(new_net_6765),
		.dout(new_net_6766)
	);

	bfr new_net_6767_bfr_after (
		.din(new_net_6766),
		.dout(new_net_6767)
	);

	bfr new_net_6768_bfr_after (
		.din(new_net_6767),
		.dout(new_net_6768)
	);

	bfr new_net_6769_bfr_after (
		.din(new_net_6768),
		.dout(new_net_6769)
	);

	bfr new_net_6770_bfr_after (
		.din(new_net_6769),
		.dout(new_net_6770)
	);

	bfr new_net_6771_bfr_after (
		.din(new_net_6770),
		.dout(new_net_6771)
	);

	bfr new_net_6772_bfr_after (
		.din(new_net_6771),
		.dout(new_net_6772)
	);

	bfr new_net_6773_bfr_after (
		.din(new_net_6772),
		.dout(new_net_6773)
	);

	bfr new_net_6774_bfr_after (
		.din(new_net_6773),
		.dout(new_net_6774)
	);

	bfr new_net_6775_bfr_after (
		.din(new_net_6774),
		.dout(new_net_6775)
	);

	bfr new_net_6776_bfr_after (
		.din(new_net_6775),
		.dout(new_net_6776)
	);

	bfr new_net_6777_bfr_after (
		.din(new_net_6776),
		.dout(new_net_6777)
	);

	bfr new_net_6778_bfr_after (
		.din(new_net_6777),
		.dout(new_net_6778)
	);

	bfr new_net_6779_bfr_after (
		.din(new_net_6778),
		.dout(new_net_6779)
	);

	bfr new_net_6780_bfr_after (
		.din(new_net_6779),
		.dout(new_net_6780)
	);

	bfr new_net_6781_bfr_after (
		.din(new_net_6780),
		.dout(new_net_6781)
	);

	bfr new_net_6782_bfr_after (
		.din(new_net_6781),
		.dout(new_net_6782)
	);

	bfr new_net_6783_bfr_after (
		.din(new_net_6782),
		.dout(new_net_6783)
	);

	bfr new_net_6784_bfr_after (
		.din(new_net_6783),
		.dout(new_net_6784)
	);

	bfr new_net_6785_bfr_after (
		.din(new_net_6784),
		.dout(new_net_6785)
	);

	bfr new_net_6786_bfr_after (
		.din(new_net_6785),
		.dout(new_net_6786)
	);

	bfr new_net_6787_bfr_after (
		.din(new_net_6786),
		.dout(new_net_6787)
	);

	bfr new_net_6788_bfr_after (
		.din(new_net_6787),
		.dout(new_net_6788)
	);

	bfr new_net_6789_bfr_after (
		.din(new_net_6788),
		.dout(new_net_6789)
	);

	bfr new_net_6790_bfr_after (
		.din(new_net_6789),
		.dout(new_net_6790)
	);

	spl2 _0447__v_fanout (
		.a(new_net_6790),
		.b(new_net_498),
		.c(new_net_499)
	);

	spl2 _1297__v_fanout (
		.a(_1297_),
		.b(new_net_442),
		.c(new_net_443)
	);

	bfr new_net_6791_bfr_after (
		.din(_1465_),
		.dout(new_net_6791)
	);

	bfr new_net_6792_bfr_after (
		.din(new_net_6791),
		.dout(new_net_6792)
	);

	bfr new_net_6793_bfr_after (
		.din(new_net_6792),
		.dout(new_net_6793)
	);

	bfr new_net_6794_bfr_after (
		.din(new_net_6793),
		.dout(new_net_6794)
	);

	bfr new_net_6795_bfr_after (
		.din(new_net_6794),
		.dout(new_net_6795)
	);

	bfr new_net_6796_bfr_after (
		.din(new_net_6795),
		.dout(new_net_6796)
	);

	bfr new_net_6797_bfr_after (
		.din(new_net_6796),
		.dout(new_net_6797)
	);

	bfr new_net_6798_bfr_after (
		.din(new_net_6797),
		.dout(new_net_6798)
	);

	bfr new_net_6799_bfr_after (
		.din(new_net_6798),
		.dout(new_net_6799)
	);

	bfr new_net_6800_bfr_after (
		.din(new_net_6799),
		.dout(new_net_6800)
	);

	bfr new_net_6801_bfr_after (
		.din(new_net_6800),
		.dout(new_net_6801)
	);

	bfr new_net_6802_bfr_after (
		.din(new_net_6801),
		.dout(new_net_6802)
	);

	bfr new_net_6803_bfr_after (
		.din(new_net_6802),
		.dout(new_net_6803)
	);

	bfr new_net_6804_bfr_after (
		.din(new_net_6803),
		.dout(new_net_6804)
	);

	bfr new_net_6805_bfr_after (
		.din(new_net_6804),
		.dout(new_net_6805)
	);

	bfr new_net_6806_bfr_after (
		.din(new_net_6805),
		.dout(new_net_6806)
	);

	bfr new_net_6807_bfr_after (
		.din(new_net_6806),
		.dout(new_net_6807)
	);

	bfr new_net_6808_bfr_after (
		.din(new_net_6807),
		.dout(new_net_6808)
	);

	bfr new_net_6809_bfr_after (
		.din(new_net_6808),
		.dout(new_net_6809)
	);

	bfr new_net_6810_bfr_after (
		.din(new_net_6809),
		.dout(new_net_6810)
	);

	bfr new_net_6811_bfr_after (
		.din(new_net_6810),
		.dout(new_net_6811)
	);

	bfr new_net_6812_bfr_after (
		.din(new_net_6811),
		.dout(new_net_6812)
	);

	bfr new_net_6813_bfr_after (
		.din(new_net_6812),
		.dout(new_net_6813)
	);

	bfr new_net_6814_bfr_after (
		.din(new_net_6813),
		.dout(new_net_6814)
	);

	bfr new_net_6815_bfr_after (
		.din(new_net_6814),
		.dout(new_net_6815)
	);

	bfr new_net_6816_bfr_after (
		.din(new_net_6815),
		.dout(new_net_6816)
	);

	bfr new_net_6817_bfr_after (
		.din(new_net_6816),
		.dout(new_net_6817)
	);

	bfr new_net_6818_bfr_after (
		.din(new_net_6817),
		.dout(new_net_6818)
	);

	bfr new_net_6819_bfr_after (
		.din(new_net_6818),
		.dout(new_net_6819)
	);

	bfr new_net_6820_bfr_after (
		.din(new_net_6819),
		.dout(new_net_6820)
	);

	bfr new_net_6821_bfr_after (
		.din(new_net_6820),
		.dout(new_net_6821)
	);

	bfr new_net_6822_bfr_after (
		.din(new_net_6821),
		.dout(new_net_6822)
	);

	bfr new_net_6823_bfr_after (
		.din(new_net_6822),
		.dout(new_net_6823)
	);

	bfr new_net_6824_bfr_after (
		.din(new_net_6823),
		.dout(new_net_6824)
	);

	bfr new_net_6825_bfr_after (
		.din(new_net_6824),
		.dout(new_net_6825)
	);

	bfr new_net_6826_bfr_after (
		.din(new_net_6825),
		.dout(new_net_6826)
	);

	bfr new_net_6827_bfr_after (
		.din(new_net_6826),
		.dout(new_net_6827)
	);

	bfr new_net_6828_bfr_after (
		.din(new_net_6827),
		.dout(new_net_6828)
	);

	bfr new_net_6829_bfr_after (
		.din(new_net_6828),
		.dout(new_net_6829)
	);

	bfr new_net_6830_bfr_after (
		.din(new_net_6829),
		.dout(new_net_6830)
	);

	bfr new_net_6831_bfr_after (
		.din(new_net_6830),
		.dout(new_net_6831)
	);

	bfr new_net_6832_bfr_after (
		.din(new_net_6831),
		.dout(new_net_6832)
	);

	bfr new_net_6833_bfr_after (
		.din(new_net_6832),
		.dout(new_net_6833)
	);

	bfr new_net_6834_bfr_after (
		.din(new_net_6833),
		.dout(new_net_6834)
	);

	bfr new_net_6835_bfr_after (
		.din(new_net_6834),
		.dout(new_net_6835)
	);

	bfr new_net_6836_bfr_after (
		.din(new_net_6835),
		.dout(new_net_6836)
	);

	bfr new_net_6837_bfr_after (
		.din(new_net_6836),
		.dout(new_net_6837)
	);

	bfr new_net_6838_bfr_after (
		.din(new_net_6837),
		.dout(new_net_6838)
	);

	spl2 _1465__v_fanout (
		.a(new_net_6838),
		.b(new_net_773),
		.c(new_net_774)
	);

	bfr new_net_6839_bfr_after (
		.din(_0547_),
		.dout(new_net_6839)
	);

	bfr new_net_6840_bfr_after (
		.din(new_net_6839),
		.dout(new_net_6840)
	);

	bfr new_net_6841_bfr_after (
		.din(new_net_6840),
		.dout(new_net_6841)
	);

	bfr new_net_6842_bfr_after (
		.din(new_net_6841),
		.dout(new_net_6842)
	);

	bfr new_net_6843_bfr_after (
		.din(new_net_6842),
		.dout(new_net_6843)
	);

	bfr new_net_6844_bfr_after (
		.din(new_net_6843),
		.dout(new_net_6844)
	);

	bfr new_net_6845_bfr_after (
		.din(new_net_6844),
		.dout(new_net_6845)
	);

	bfr new_net_6846_bfr_after (
		.din(new_net_6845),
		.dout(new_net_6846)
	);

	bfr new_net_6847_bfr_after (
		.din(new_net_6846),
		.dout(new_net_6847)
	);

	bfr new_net_6848_bfr_after (
		.din(new_net_6847),
		.dout(new_net_6848)
	);

	bfr new_net_6849_bfr_after (
		.din(new_net_6848),
		.dout(new_net_6849)
	);

	bfr new_net_6850_bfr_after (
		.din(new_net_6849),
		.dout(new_net_6850)
	);

	bfr new_net_6851_bfr_after (
		.din(new_net_6850),
		.dout(new_net_6851)
	);

	bfr new_net_6852_bfr_after (
		.din(new_net_6851),
		.dout(new_net_6852)
	);

	bfr new_net_6853_bfr_after (
		.din(new_net_6852),
		.dout(new_net_6853)
	);

	bfr new_net_6854_bfr_after (
		.din(new_net_6853),
		.dout(new_net_6854)
	);

	bfr new_net_6855_bfr_after (
		.din(new_net_6854),
		.dout(new_net_6855)
	);

	bfr new_net_6856_bfr_after (
		.din(new_net_6855),
		.dout(new_net_6856)
	);

	bfr new_net_6857_bfr_after (
		.din(new_net_6856),
		.dout(new_net_6857)
	);

	bfr new_net_6858_bfr_after (
		.din(new_net_6857),
		.dout(new_net_6858)
	);

	bfr new_net_6859_bfr_after (
		.din(new_net_6858),
		.dout(new_net_6859)
	);

	bfr new_net_6860_bfr_after (
		.din(new_net_6859),
		.dout(new_net_6860)
	);

	bfr new_net_6861_bfr_after (
		.din(new_net_6860),
		.dout(new_net_6861)
	);

	bfr new_net_6862_bfr_after (
		.din(new_net_6861),
		.dout(new_net_6862)
	);

	bfr new_net_6863_bfr_after (
		.din(new_net_6862),
		.dout(new_net_6863)
	);

	bfr new_net_6864_bfr_after (
		.din(new_net_6863),
		.dout(new_net_6864)
	);

	bfr new_net_6865_bfr_after (
		.din(new_net_6864),
		.dout(new_net_6865)
	);

	bfr new_net_6866_bfr_after (
		.din(new_net_6865),
		.dout(new_net_6866)
	);

	bfr new_net_6867_bfr_after (
		.din(new_net_6866),
		.dout(new_net_6867)
	);

	bfr new_net_6868_bfr_after (
		.din(new_net_6867),
		.dout(new_net_6868)
	);

	bfr new_net_6869_bfr_after (
		.din(new_net_6868),
		.dout(new_net_6869)
	);

	bfr new_net_6870_bfr_after (
		.din(new_net_6869),
		.dout(new_net_6870)
	);

	bfr new_net_6871_bfr_after (
		.din(new_net_6870),
		.dout(new_net_6871)
	);

	bfr new_net_6872_bfr_after (
		.din(new_net_6871),
		.dout(new_net_6872)
	);

	bfr new_net_6873_bfr_after (
		.din(new_net_6872),
		.dout(new_net_6873)
	);

	bfr new_net_6874_bfr_after (
		.din(new_net_6873),
		.dout(new_net_6874)
	);

	bfr new_net_6875_bfr_after (
		.din(new_net_6874),
		.dout(new_net_6875)
	);

	bfr new_net_6876_bfr_after (
		.din(new_net_6875),
		.dout(new_net_6876)
	);

	bfr new_net_6877_bfr_after (
		.din(new_net_6876),
		.dout(new_net_6877)
	);

	bfr new_net_6878_bfr_after (
		.din(new_net_6877),
		.dout(new_net_6878)
	);

	bfr new_net_6879_bfr_after (
		.din(new_net_6878),
		.dout(new_net_6879)
	);

	bfr new_net_6880_bfr_after (
		.din(new_net_6879),
		.dout(new_net_6880)
	);

	spl2 _0547__v_fanout (
		.a(new_net_6880),
		.b(new_net_3065),
		.c(new_net_3066)
	);

	bfr new_net_6881_bfr_after (
		.din(_0346_),
		.dout(new_net_6881)
	);

	bfr new_net_6882_bfr_after (
		.din(new_net_6881),
		.dout(new_net_6882)
	);

	bfr new_net_6883_bfr_after (
		.din(new_net_6882),
		.dout(new_net_6883)
	);

	bfr new_net_6884_bfr_after (
		.din(new_net_6883),
		.dout(new_net_6884)
	);

	bfr new_net_6885_bfr_after (
		.din(new_net_6884),
		.dout(new_net_6885)
	);

	bfr new_net_6886_bfr_after (
		.din(new_net_6885),
		.dout(new_net_6886)
	);

	bfr new_net_6887_bfr_after (
		.din(new_net_6886),
		.dout(new_net_6887)
	);

	bfr new_net_6888_bfr_after (
		.din(new_net_6887),
		.dout(new_net_6888)
	);

	bfr new_net_6889_bfr_after (
		.din(new_net_6888),
		.dout(new_net_6889)
	);

	bfr new_net_6890_bfr_after (
		.din(new_net_6889),
		.dout(new_net_6890)
	);

	bfr new_net_6891_bfr_after (
		.din(new_net_6890),
		.dout(new_net_6891)
	);

	bfr new_net_6892_bfr_after (
		.din(new_net_6891),
		.dout(new_net_6892)
	);

	bfr new_net_6893_bfr_after (
		.din(new_net_6892),
		.dout(new_net_6893)
	);

	bfr new_net_6894_bfr_after (
		.din(new_net_6893),
		.dout(new_net_6894)
	);

	bfr new_net_6895_bfr_after (
		.din(new_net_6894),
		.dout(new_net_6895)
	);

	bfr new_net_6896_bfr_after (
		.din(new_net_6895),
		.dout(new_net_6896)
	);

	bfr new_net_6897_bfr_after (
		.din(new_net_6896),
		.dout(new_net_6897)
	);

	bfr new_net_6898_bfr_after (
		.din(new_net_6897),
		.dout(new_net_6898)
	);

	bfr new_net_6899_bfr_after (
		.din(new_net_6898),
		.dout(new_net_6899)
	);

	bfr new_net_6900_bfr_after (
		.din(new_net_6899),
		.dout(new_net_6900)
	);

	bfr new_net_6901_bfr_after (
		.din(new_net_6900),
		.dout(new_net_6901)
	);

	bfr new_net_6902_bfr_after (
		.din(new_net_6901),
		.dout(new_net_6902)
	);

	bfr new_net_6903_bfr_after (
		.din(new_net_6902),
		.dout(new_net_6903)
	);

	bfr new_net_6904_bfr_after (
		.din(new_net_6903),
		.dout(new_net_6904)
	);

	bfr new_net_6905_bfr_after (
		.din(new_net_6904),
		.dout(new_net_6905)
	);

	bfr new_net_6906_bfr_after (
		.din(new_net_6905),
		.dout(new_net_6906)
	);

	bfr new_net_6907_bfr_after (
		.din(new_net_6906),
		.dout(new_net_6907)
	);

	bfr new_net_6908_bfr_after (
		.din(new_net_6907),
		.dout(new_net_6908)
	);

	bfr new_net_6909_bfr_after (
		.din(new_net_6908),
		.dout(new_net_6909)
	);

	bfr new_net_6910_bfr_after (
		.din(new_net_6909),
		.dout(new_net_6910)
	);

	bfr new_net_6911_bfr_after (
		.din(new_net_6910),
		.dout(new_net_6911)
	);

	bfr new_net_6912_bfr_after (
		.din(new_net_6911),
		.dout(new_net_6912)
	);

	bfr new_net_6913_bfr_after (
		.din(new_net_6912),
		.dout(new_net_6913)
	);

	bfr new_net_6914_bfr_after (
		.din(new_net_6913),
		.dout(new_net_6914)
	);

	bfr new_net_6915_bfr_after (
		.din(new_net_6914),
		.dout(new_net_6915)
	);

	bfr new_net_6916_bfr_after (
		.din(new_net_6915),
		.dout(new_net_6916)
	);

	bfr new_net_6917_bfr_after (
		.din(new_net_6916),
		.dout(new_net_6917)
	);

	bfr new_net_6918_bfr_after (
		.din(new_net_6917),
		.dout(new_net_6918)
	);

	spl2 _0346__v_fanout (
		.a(new_net_6918),
		.b(new_net_2337),
		.c(new_net_2338)
	);

	bfr new_net_6919_bfr_after (
		.din(_0237_),
		.dout(new_net_6919)
	);

	bfr new_net_6920_bfr_after (
		.din(new_net_6919),
		.dout(new_net_6920)
	);

	bfr new_net_6921_bfr_after (
		.din(new_net_6920),
		.dout(new_net_6921)
	);

	bfr new_net_6922_bfr_after (
		.din(new_net_6921),
		.dout(new_net_6922)
	);

	bfr new_net_6923_bfr_after (
		.din(new_net_6922),
		.dout(new_net_6923)
	);

	bfr new_net_6924_bfr_after (
		.din(new_net_6923),
		.dout(new_net_6924)
	);

	bfr new_net_6925_bfr_after (
		.din(new_net_6924),
		.dout(new_net_6925)
	);

	bfr new_net_6926_bfr_after (
		.din(new_net_6925),
		.dout(new_net_6926)
	);

	bfr new_net_6927_bfr_after (
		.din(new_net_6926),
		.dout(new_net_6927)
	);

	bfr new_net_6928_bfr_after (
		.din(new_net_6927),
		.dout(new_net_6928)
	);

	bfr new_net_6929_bfr_after (
		.din(new_net_6928),
		.dout(new_net_6929)
	);

	bfr new_net_6930_bfr_after (
		.din(new_net_6929),
		.dout(new_net_6930)
	);

	bfr new_net_6931_bfr_after (
		.din(new_net_6930),
		.dout(new_net_6931)
	);

	bfr new_net_6932_bfr_after (
		.din(new_net_6931),
		.dout(new_net_6932)
	);

	spl2 _0237__v_fanout (
		.a(new_net_6932),
		.b(new_net_568),
		.c(new_net_569)
	);

	bfr new_net_6933_bfr_after (
		.din(_1205_),
		.dout(new_net_6933)
	);

	bfr new_net_6934_bfr_after (
		.din(new_net_6933),
		.dout(new_net_6934)
	);

	bfr new_net_6935_bfr_after (
		.din(new_net_6934),
		.dout(new_net_6935)
	);

	bfr new_net_6936_bfr_after (
		.din(new_net_6935),
		.dout(new_net_6936)
	);

	bfr new_net_6937_bfr_after (
		.din(new_net_6936),
		.dout(new_net_6937)
	);

	bfr new_net_6938_bfr_after (
		.din(new_net_6937),
		.dout(new_net_6938)
	);

	bfr new_net_6939_bfr_after (
		.din(new_net_6938),
		.dout(new_net_6939)
	);

	bfr new_net_6940_bfr_after (
		.din(new_net_6939),
		.dout(new_net_6940)
	);

	bfr new_net_6941_bfr_after (
		.din(new_net_6940),
		.dout(new_net_6941)
	);

	bfr new_net_6942_bfr_after (
		.din(new_net_6941),
		.dout(new_net_6942)
	);

	bfr new_net_6943_bfr_after (
		.din(new_net_6942),
		.dout(new_net_6943)
	);

	bfr new_net_6944_bfr_after (
		.din(new_net_6943),
		.dout(new_net_6944)
	);

	bfr new_net_6945_bfr_after (
		.din(new_net_6944),
		.dout(new_net_6945)
	);

	bfr new_net_6946_bfr_after (
		.din(new_net_6945),
		.dout(new_net_6946)
	);

	bfr new_net_6947_bfr_after (
		.din(new_net_6946),
		.dout(new_net_6947)
	);

	bfr new_net_6948_bfr_after (
		.din(new_net_6947),
		.dout(new_net_6948)
	);

	bfr new_net_6949_bfr_after (
		.din(new_net_6948),
		.dout(new_net_6949)
	);

	bfr new_net_6950_bfr_after (
		.din(new_net_6949),
		.dout(new_net_6950)
	);

	bfr new_net_6951_bfr_after (
		.din(new_net_6950),
		.dout(new_net_6951)
	);

	bfr new_net_6952_bfr_after (
		.din(new_net_6951),
		.dout(new_net_6952)
	);

	bfr new_net_6953_bfr_after (
		.din(new_net_6952),
		.dout(new_net_6953)
	);

	bfr new_net_6954_bfr_after (
		.din(new_net_6953),
		.dout(new_net_6954)
	);

	bfr new_net_6955_bfr_after (
		.din(new_net_6954),
		.dout(new_net_6955)
	);

	bfr new_net_6956_bfr_after (
		.din(new_net_6955),
		.dout(new_net_6956)
	);

	bfr new_net_6957_bfr_after (
		.din(new_net_6956),
		.dout(new_net_6957)
	);

	bfr new_net_6958_bfr_after (
		.din(new_net_6957),
		.dout(new_net_6958)
	);

	bfr new_net_6959_bfr_after (
		.din(new_net_6958),
		.dout(new_net_6959)
	);

	bfr new_net_6960_bfr_after (
		.din(new_net_6959),
		.dout(new_net_6960)
	);

	bfr new_net_6961_bfr_after (
		.din(new_net_6960),
		.dout(new_net_6961)
	);

	bfr new_net_6962_bfr_after (
		.din(new_net_6961),
		.dout(new_net_6962)
	);

	bfr new_net_6963_bfr_after (
		.din(new_net_6962),
		.dout(new_net_6963)
	);

	bfr new_net_6964_bfr_after (
		.din(new_net_6963),
		.dout(new_net_6964)
	);

	bfr new_net_6965_bfr_after (
		.din(new_net_6964),
		.dout(new_net_6965)
	);

	bfr new_net_6966_bfr_after (
		.din(new_net_6965),
		.dout(new_net_6966)
	);

	bfr new_net_6967_bfr_after (
		.din(new_net_6966),
		.dout(new_net_6967)
	);

	bfr new_net_6968_bfr_after (
		.din(new_net_6967),
		.dout(new_net_6968)
	);

	bfr new_net_6969_bfr_after (
		.din(new_net_6968),
		.dout(new_net_6969)
	);

	bfr new_net_6970_bfr_after (
		.din(new_net_6969),
		.dout(new_net_6970)
	);

	bfr new_net_6971_bfr_after (
		.din(new_net_6970),
		.dout(new_net_6971)
	);

	bfr new_net_6972_bfr_after (
		.din(new_net_6971),
		.dout(new_net_6972)
	);

	bfr new_net_6973_bfr_after (
		.din(new_net_6972),
		.dout(new_net_6973)
	);

	bfr new_net_6974_bfr_after (
		.din(new_net_6973),
		.dout(new_net_6974)
	);

	bfr new_net_6975_bfr_after (
		.din(new_net_6974),
		.dout(new_net_6975)
	);

	bfr new_net_6976_bfr_after (
		.din(new_net_6975),
		.dout(new_net_6976)
	);

	bfr new_net_6977_bfr_after (
		.din(new_net_6976),
		.dout(new_net_6977)
	);

	bfr new_net_6978_bfr_after (
		.din(new_net_6977),
		.dout(new_net_6978)
	);

	bfr new_net_6979_bfr_after (
		.din(new_net_6978),
		.dout(new_net_6979)
	);

	bfr new_net_6980_bfr_after (
		.din(new_net_6979),
		.dout(new_net_6980)
	);

	bfr new_net_6981_bfr_after (
		.din(new_net_6980),
		.dout(new_net_6981)
	);

	bfr new_net_6982_bfr_after (
		.din(new_net_6981),
		.dout(new_net_6982)
	);

	bfr new_net_6983_bfr_after (
		.din(new_net_6982),
		.dout(new_net_6983)
	);

	bfr new_net_6984_bfr_after (
		.din(new_net_6983),
		.dout(new_net_6984)
	);

	bfr new_net_6985_bfr_after (
		.din(new_net_6984),
		.dout(new_net_6985)
	);

	bfr new_net_6986_bfr_after (
		.din(new_net_6985),
		.dout(new_net_6986)
	);

	bfr new_net_6987_bfr_after (
		.din(new_net_6986),
		.dout(new_net_6987)
	);

	bfr new_net_6988_bfr_after (
		.din(new_net_6987),
		.dout(new_net_6988)
	);

	bfr new_net_6989_bfr_after (
		.din(new_net_6988),
		.dout(new_net_6989)
	);

	bfr new_net_6990_bfr_after (
		.din(new_net_6989),
		.dout(new_net_6990)
	);

	bfr new_net_6991_bfr_after (
		.din(new_net_6990),
		.dout(new_net_6991)
	);

	bfr new_net_6992_bfr_after (
		.din(new_net_6991),
		.dout(new_net_6992)
	);

	bfr new_net_6993_bfr_after (
		.din(new_net_6992),
		.dout(new_net_6993)
	);

	bfr new_net_6994_bfr_after (
		.din(new_net_6993),
		.dout(new_net_6994)
	);

	bfr new_net_6995_bfr_after (
		.din(new_net_6994),
		.dout(new_net_6995)
	);

	bfr new_net_6996_bfr_after (
		.din(new_net_6995),
		.dout(new_net_6996)
	);

	spl2 _1205__v_fanout (
		.a(new_net_6996),
		.b(new_net_116),
		.c(new_net_117)
	);

	bfr new_net_6997_bfr_after (
		.din(_0443_),
		.dout(new_net_6997)
	);

	bfr new_net_6998_bfr_after (
		.din(new_net_6997),
		.dout(new_net_6998)
	);

	bfr new_net_6999_bfr_after (
		.din(new_net_6998),
		.dout(new_net_6999)
	);

	bfr new_net_7000_bfr_after (
		.din(new_net_6999),
		.dout(new_net_7000)
	);

	bfr new_net_7001_bfr_after (
		.din(new_net_7000),
		.dout(new_net_7001)
	);

	bfr new_net_7002_bfr_after (
		.din(new_net_7001),
		.dout(new_net_7002)
	);

	bfr new_net_7003_bfr_after (
		.din(new_net_7002),
		.dout(new_net_7003)
	);

	bfr new_net_7004_bfr_after (
		.din(new_net_7003),
		.dout(new_net_7004)
	);

	bfr new_net_7005_bfr_after (
		.din(new_net_7004),
		.dout(new_net_7005)
	);

	bfr new_net_7006_bfr_after (
		.din(new_net_7005),
		.dout(new_net_7006)
	);

	bfr new_net_7007_bfr_after (
		.din(new_net_7006),
		.dout(new_net_7007)
	);

	bfr new_net_7008_bfr_after (
		.din(new_net_7007),
		.dout(new_net_7008)
	);

	bfr new_net_7009_bfr_after (
		.din(new_net_7008),
		.dout(new_net_7009)
	);

	bfr new_net_7010_bfr_after (
		.din(new_net_7009),
		.dout(new_net_7010)
	);

	bfr new_net_7011_bfr_after (
		.din(new_net_7010),
		.dout(new_net_7011)
	);

	bfr new_net_7012_bfr_after (
		.din(new_net_7011),
		.dout(new_net_7012)
	);

	bfr new_net_7013_bfr_after (
		.din(new_net_7012),
		.dout(new_net_7013)
	);

	bfr new_net_7014_bfr_after (
		.din(new_net_7013),
		.dout(new_net_7014)
	);

	bfr new_net_7015_bfr_after (
		.din(new_net_7014),
		.dout(new_net_7015)
	);

	bfr new_net_7016_bfr_after (
		.din(new_net_7015),
		.dout(new_net_7016)
	);

	bfr new_net_7017_bfr_after (
		.din(new_net_7016),
		.dout(new_net_7017)
	);

	bfr new_net_7018_bfr_after (
		.din(new_net_7017),
		.dout(new_net_7018)
	);

	bfr new_net_7019_bfr_after (
		.din(new_net_7018),
		.dout(new_net_7019)
	);

	bfr new_net_7020_bfr_after (
		.din(new_net_7019),
		.dout(new_net_7020)
	);

	bfr new_net_7021_bfr_after (
		.din(new_net_7020),
		.dout(new_net_7021)
	);

	bfr new_net_7022_bfr_after (
		.din(new_net_7021),
		.dout(new_net_7022)
	);

	bfr new_net_7023_bfr_after (
		.din(new_net_7022),
		.dout(new_net_7023)
	);

	bfr new_net_7024_bfr_after (
		.din(new_net_7023),
		.dout(new_net_7024)
	);

	bfr new_net_7025_bfr_after (
		.din(new_net_7024),
		.dout(new_net_7025)
	);

	bfr new_net_7026_bfr_after (
		.din(new_net_7025),
		.dout(new_net_7026)
	);

	bfr new_net_7027_bfr_after (
		.din(new_net_7026),
		.dout(new_net_7027)
	);

	bfr new_net_7028_bfr_after (
		.din(new_net_7027),
		.dout(new_net_7028)
	);

	bfr new_net_7029_bfr_after (
		.din(new_net_7028),
		.dout(new_net_7029)
	);

	bfr new_net_7030_bfr_after (
		.din(new_net_7029),
		.dout(new_net_7030)
	);

	bfr new_net_7031_bfr_after (
		.din(new_net_7030),
		.dout(new_net_7031)
	);

	bfr new_net_7032_bfr_after (
		.din(new_net_7031),
		.dout(new_net_7032)
	);

	bfr new_net_7033_bfr_after (
		.din(new_net_7032),
		.dout(new_net_7033)
	);

	bfr new_net_7034_bfr_after (
		.din(new_net_7033),
		.dout(new_net_7034)
	);

	bfr new_net_7035_bfr_after (
		.din(new_net_7034),
		.dout(new_net_7035)
	);

	bfr new_net_7036_bfr_after (
		.din(new_net_7035),
		.dout(new_net_7036)
	);

	bfr new_net_7037_bfr_after (
		.din(new_net_7036),
		.dout(new_net_7037)
	);

	bfr new_net_7038_bfr_after (
		.din(new_net_7037),
		.dout(new_net_7038)
	);

	bfr new_net_7039_bfr_after (
		.din(new_net_7038),
		.dout(new_net_7039)
	);

	bfr new_net_7040_bfr_after (
		.din(new_net_7039),
		.dout(new_net_7040)
	);

	bfr new_net_7041_bfr_after (
		.din(new_net_7040),
		.dout(new_net_7041)
	);

	bfr new_net_7042_bfr_after (
		.din(new_net_7041),
		.dout(new_net_7042)
	);

	bfr new_net_7043_bfr_after (
		.din(new_net_7042),
		.dout(new_net_7043)
	);

	bfr new_net_7044_bfr_after (
		.din(new_net_7043),
		.dout(new_net_7044)
	);

	bfr new_net_7045_bfr_after (
		.din(new_net_7044),
		.dout(new_net_7045)
	);

	bfr new_net_7046_bfr_after (
		.din(new_net_7045),
		.dout(new_net_7046)
	);

	bfr new_net_7047_bfr_after (
		.din(new_net_7046),
		.dout(new_net_7047)
	);

	bfr new_net_7048_bfr_after (
		.din(new_net_7047),
		.dout(new_net_7048)
	);

	bfr new_net_7049_bfr_after (
		.din(new_net_7048),
		.dout(new_net_7049)
	);

	bfr new_net_7050_bfr_after (
		.din(new_net_7049),
		.dout(new_net_7050)
	);

	bfr new_net_7051_bfr_after (
		.din(new_net_7050),
		.dout(new_net_7051)
	);

	bfr new_net_7052_bfr_after (
		.din(new_net_7051),
		.dout(new_net_7052)
	);

	bfr new_net_7053_bfr_after (
		.din(new_net_7052),
		.dout(new_net_7053)
	);

	bfr new_net_7054_bfr_after (
		.din(new_net_7053),
		.dout(new_net_7054)
	);

	bfr new_net_7055_bfr_after (
		.din(new_net_7054),
		.dout(new_net_7055)
	);

	bfr new_net_7056_bfr_after (
		.din(new_net_7055),
		.dout(new_net_7056)
	);

	bfr new_net_7057_bfr_after (
		.din(new_net_7056),
		.dout(new_net_7057)
	);

	bfr new_net_7058_bfr_after (
		.din(new_net_7057),
		.dout(new_net_7058)
	);

	bfr new_net_7059_bfr_after (
		.din(new_net_7058),
		.dout(new_net_7059)
	);

	bfr new_net_7060_bfr_after (
		.din(new_net_7059),
		.dout(new_net_7060)
	);

	bfr new_net_7061_bfr_after (
		.din(new_net_7060),
		.dout(new_net_7061)
	);

	bfr new_net_7062_bfr_after (
		.din(new_net_7061),
		.dout(new_net_7062)
	);

	bfr new_net_7063_bfr_after (
		.din(new_net_7062),
		.dout(new_net_7063)
	);

	bfr new_net_7064_bfr_after (
		.din(new_net_7063),
		.dout(new_net_7064)
	);

	bfr new_net_7065_bfr_after (
		.din(new_net_7064),
		.dout(new_net_7065)
	);

	bfr new_net_7066_bfr_after (
		.din(new_net_7065),
		.dout(new_net_7066)
	);

	bfr new_net_7067_bfr_after (
		.din(new_net_7066),
		.dout(new_net_7067)
	);

	bfr new_net_7068_bfr_after (
		.din(new_net_7067),
		.dout(new_net_7068)
	);

	spl2 _0443__v_fanout (
		.a(new_net_7068),
		.b(new_net_1674),
		.c(new_net_1675)
	);

	bfr new_net_7069_bfr_after (
		.din(_1680_),
		.dout(new_net_7069)
	);

	bfr new_net_7070_bfr_after (
		.din(new_net_7069),
		.dout(new_net_7070)
	);

	bfr new_net_7071_bfr_after (
		.din(new_net_7070),
		.dout(new_net_7071)
	);

	bfr new_net_7072_bfr_after (
		.din(new_net_7071),
		.dout(new_net_7072)
	);

	bfr new_net_7073_bfr_after (
		.din(new_net_7072),
		.dout(new_net_7073)
	);

	bfr new_net_7074_bfr_after (
		.din(new_net_7073),
		.dout(new_net_7074)
	);

	bfr new_net_7075_bfr_after (
		.din(new_net_7074),
		.dout(new_net_7075)
	);

	bfr new_net_7076_bfr_after (
		.din(new_net_7075),
		.dout(new_net_7076)
	);

	bfr new_net_7077_bfr_after (
		.din(new_net_7076),
		.dout(new_net_7077)
	);

	bfr new_net_7078_bfr_after (
		.din(new_net_7077),
		.dout(new_net_7078)
	);

	bfr new_net_7079_bfr_after (
		.din(new_net_7078),
		.dout(new_net_7079)
	);

	bfr new_net_7080_bfr_after (
		.din(new_net_7079),
		.dout(new_net_7080)
	);

	bfr new_net_7081_bfr_after (
		.din(new_net_7080),
		.dout(new_net_7081)
	);

	bfr new_net_7082_bfr_after (
		.din(new_net_7081),
		.dout(new_net_7082)
	);

	bfr new_net_7083_bfr_after (
		.din(new_net_7082),
		.dout(new_net_7083)
	);

	bfr new_net_7084_bfr_after (
		.din(new_net_7083),
		.dout(new_net_7084)
	);

	bfr new_net_7085_bfr_after (
		.din(new_net_7084),
		.dout(new_net_7085)
	);

	bfr new_net_7086_bfr_after (
		.din(new_net_7085),
		.dout(new_net_7086)
	);

	bfr new_net_7087_bfr_after (
		.din(new_net_7086),
		.dout(new_net_7087)
	);

	bfr new_net_7088_bfr_after (
		.din(new_net_7087),
		.dout(new_net_7088)
	);

	bfr new_net_7089_bfr_after (
		.din(new_net_7088),
		.dout(new_net_7089)
	);

	bfr new_net_7090_bfr_after (
		.din(new_net_7089),
		.dout(new_net_7090)
	);

	bfr new_net_7091_bfr_after (
		.din(new_net_7090),
		.dout(new_net_7091)
	);

	bfr new_net_7092_bfr_after (
		.din(new_net_7091),
		.dout(new_net_7092)
	);

	bfr new_net_7093_bfr_after (
		.din(new_net_7092),
		.dout(new_net_7093)
	);

	bfr new_net_7094_bfr_after (
		.din(new_net_7093),
		.dout(new_net_7094)
	);

	bfr new_net_7095_bfr_after (
		.din(new_net_7094),
		.dout(new_net_7095)
	);

	bfr new_net_7096_bfr_after (
		.din(new_net_7095),
		.dout(new_net_7096)
	);

	bfr new_net_7097_bfr_after (
		.din(new_net_7096),
		.dout(new_net_7097)
	);

	bfr new_net_7098_bfr_after (
		.din(new_net_7097),
		.dout(new_net_7098)
	);

	bfr new_net_7099_bfr_after (
		.din(new_net_7098),
		.dout(new_net_7099)
	);

	bfr new_net_7100_bfr_after (
		.din(new_net_7099),
		.dout(new_net_7100)
	);

	bfr new_net_7101_bfr_after (
		.din(new_net_7100),
		.dout(new_net_7101)
	);

	bfr new_net_7102_bfr_after (
		.din(new_net_7101),
		.dout(new_net_7102)
	);

	bfr new_net_7103_bfr_after (
		.din(new_net_7102),
		.dout(new_net_7103)
	);

	bfr new_net_7104_bfr_after (
		.din(new_net_7103),
		.dout(new_net_7104)
	);

	bfr new_net_7105_bfr_after (
		.din(new_net_7104),
		.dout(new_net_7105)
	);

	bfr new_net_7106_bfr_after (
		.din(new_net_7105),
		.dout(new_net_7106)
	);

	bfr new_net_7107_bfr_after (
		.din(new_net_7106),
		.dout(new_net_7107)
	);

	bfr new_net_7108_bfr_after (
		.din(new_net_7107),
		.dout(new_net_7108)
	);

	bfr new_net_7109_bfr_after (
		.din(new_net_7108),
		.dout(new_net_7109)
	);

	bfr new_net_7110_bfr_after (
		.din(new_net_7109),
		.dout(new_net_7110)
	);

	bfr new_net_7111_bfr_after (
		.din(new_net_7110),
		.dout(new_net_7111)
	);

	bfr new_net_7112_bfr_after (
		.din(new_net_7111),
		.dout(new_net_7112)
	);

	bfr new_net_7113_bfr_after (
		.din(new_net_7112),
		.dout(new_net_7113)
	);

	bfr new_net_7114_bfr_after (
		.din(new_net_7113),
		.dout(new_net_7114)
	);

	bfr new_net_7115_bfr_after (
		.din(new_net_7114),
		.dout(new_net_7115)
	);

	bfr new_net_7116_bfr_after (
		.din(new_net_7115),
		.dout(new_net_7116)
	);

	bfr new_net_7117_bfr_after (
		.din(new_net_7116),
		.dout(new_net_7117)
	);

	bfr new_net_7118_bfr_after (
		.din(new_net_7117),
		.dout(new_net_7118)
	);

	bfr new_net_7119_bfr_after (
		.din(new_net_7118),
		.dout(new_net_7119)
	);

	bfr new_net_7120_bfr_after (
		.din(new_net_7119),
		.dout(new_net_7120)
	);

	bfr new_net_7121_bfr_after (
		.din(new_net_7120),
		.dout(new_net_7121)
	);

	bfr new_net_7122_bfr_after (
		.din(new_net_7121),
		.dout(new_net_7122)
	);

	bfr new_net_7123_bfr_after (
		.din(new_net_7122),
		.dout(new_net_7123)
	);

	bfr new_net_7124_bfr_after (
		.din(new_net_7123),
		.dout(new_net_7124)
	);

	bfr new_net_7125_bfr_after (
		.din(new_net_7124),
		.dout(new_net_7125)
	);

	bfr new_net_7126_bfr_after (
		.din(new_net_7125),
		.dout(new_net_7126)
	);

	bfr new_net_7127_bfr_after (
		.din(new_net_7126),
		.dout(new_net_7127)
	);

	bfr new_net_7128_bfr_after (
		.din(new_net_7127),
		.dout(new_net_7128)
	);

	bfr new_net_7129_bfr_after (
		.din(new_net_7128),
		.dout(new_net_7129)
	);

	bfr new_net_7130_bfr_after (
		.din(new_net_7129),
		.dout(new_net_7130)
	);

	bfr new_net_7131_bfr_after (
		.din(new_net_7130),
		.dout(new_net_7131)
	);

	bfr new_net_7132_bfr_after (
		.din(new_net_7131),
		.dout(new_net_7132)
	);

	bfr new_net_7133_bfr_after (
		.din(new_net_7132),
		.dout(new_net_7133)
	);

	bfr new_net_7134_bfr_after (
		.din(new_net_7133),
		.dout(new_net_7134)
	);

	bfr new_net_7135_bfr_after (
		.din(new_net_7134),
		.dout(new_net_7135)
	);

	bfr new_net_7136_bfr_after (
		.din(new_net_7135),
		.dout(new_net_7136)
	);

	bfr new_net_7137_bfr_after (
		.din(new_net_7136),
		.dout(new_net_7137)
	);

	bfr new_net_7138_bfr_after (
		.din(new_net_7137),
		.dout(new_net_7138)
	);

	bfr new_net_7139_bfr_after (
		.din(new_net_7138),
		.dout(new_net_7139)
	);

	bfr new_net_7140_bfr_after (
		.din(new_net_7139),
		.dout(new_net_7140)
	);

	bfr new_net_7141_bfr_after (
		.din(new_net_7140),
		.dout(new_net_7141)
	);

	bfr new_net_7142_bfr_after (
		.din(new_net_7141),
		.dout(new_net_7142)
	);

	bfr new_net_7143_bfr_after (
		.din(new_net_7142),
		.dout(new_net_7143)
	);

	bfr new_net_7144_bfr_after (
		.din(new_net_7143),
		.dout(new_net_7144)
	);

	bfr new_net_7145_bfr_after (
		.din(new_net_7144),
		.dout(new_net_7145)
	);

	bfr new_net_7146_bfr_after (
		.din(new_net_7145),
		.dout(new_net_7146)
	);

	bfr new_net_7147_bfr_after (
		.din(new_net_7146),
		.dout(new_net_7147)
	);

	bfr new_net_7148_bfr_after (
		.din(new_net_7147),
		.dout(new_net_7148)
	);

	bfr new_net_7149_bfr_after (
		.din(new_net_7148),
		.dout(new_net_7149)
	);

	bfr new_net_7150_bfr_after (
		.din(new_net_7149),
		.dout(new_net_7150)
	);

	bfr new_net_7151_bfr_after (
		.din(new_net_7150),
		.dout(new_net_7151)
	);

	bfr new_net_7152_bfr_after (
		.din(new_net_7151),
		.dout(new_net_7152)
	);

	bfr new_net_7153_bfr_after (
		.din(new_net_7152),
		.dout(new_net_7153)
	);

	bfr new_net_7154_bfr_after (
		.din(new_net_7153),
		.dout(new_net_7154)
	);

	bfr new_net_7155_bfr_after (
		.din(new_net_7154),
		.dout(new_net_7155)
	);

	bfr new_net_7156_bfr_after (
		.din(new_net_7155),
		.dout(new_net_7156)
	);

	bfr new_net_7157_bfr_after (
		.din(new_net_7156),
		.dout(new_net_7157)
	);

	bfr new_net_7158_bfr_after (
		.din(new_net_7157),
		.dout(new_net_7158)
	);

	bfr new_net_7159_bfr_after (
		.din(new_net_7158),
		.dout(new_net_7159)
	);

	bfr new_net_7160_bfr_after (
		.din(new_net_7159),
		.dout(new_net_7160)
	);

	bfr new_net_7161_bfr_after (
		.din(new_net_7160),
		.dout(new_net_7161)
	);

	bfr new_net_7162_bfr_after (
		.din(new_net_7161),
		.dout(new_net_7162)
	);

	bfr new_net_7163_bfr_after (
		.din(new_net_7162),
		.dout(new_net_7163)
	);

	bfr new_net_7164_bfr_after (
		.din(new_net_7163),
		.dout(new_net_7164)
	);

	bfr new_net_7165_bfr_after (
		.din(new_net_7164),
		.dout(new_net_7165)
	);

	bfr new_net_7166_bfr_after (
		.din(new_net_7165),
		.dout(new_net_7166)
	);

	bfr new_net_7167_bfr_after (
		.din(new_net_7166),
		.dout(new_net_7167)
	);

	bfr new_net_7168_bfr_after (
		.din(new_net_7167),
		.dout(new_net_7168)
	);

	bfr new_net_7169_bfr_after (
		.din(new_net_7168),
		.dout(new_net_7169)
	);

	bfr new_net_7170_bfr_after (
		.din(new_net_7169),
		.dout(new_net_7170)
	);

	bfr new_net_7171_bfr_after (
		.din(new_net_7170),
		.dout(new_net_7171)
	);

	bfr new_net_7172_bfr_after (
		.din(new_net_7171),
		.dout(new_net_7172)
	);

	spl2 _1680__v_fanout (
		.a(new_net_7172),
		.b(new_net_1056),
		.c(new_net_1057)
	);

	bfr new_net_7173_bfr_after (
		.din(_0779_),
		.dout(new_net_7173)
	);

	bfr new_net_7174_bfr_after (
		.din(new_net_7173),
		.dout(new_net_7174)
	);

	bfr new_net_7175_bfr_after (
		.din(new_net_7174),
		.dout(new_net_7175)
	);

	bfr new_net_7176_bfr_after (
		.din(new_net_7175),
		.dout(new_net_7176)
	);

	bfr new_net_7177_bfr_after (
		.din(new_net_7176),
		.dout(new_net_7177)
	);

	bfr new_net_7178_bfr_after (
		.din(new_net_7177),
		.dout(new_net_7178)
	);

	bfr new_net_7179_bfr_after (
		.din(new_net_7178),
		.dout(new_net_7179)
	);

	bfr new_net_7180_bfr_after (
		.din(new_net_7179),
		.dout(new_net_7180)
	);

	bfr new_net_7181_bfr_after (
		.din(new_net_7180),
		.dout(new_net_7181)
	);

	bfr new_net_7182_bfr_after (
		.din(new_net_7181),
		.dout(new_net_7182)
	);

	bfr new_net_7183_bfr_after (
		.din(new_net_7182),
		.dout(new_net_7183)
	);

	bfr new_net_7184_bfr_after (
		.din(new_net_7183),
		.dout(new_net_7184)
	);

	bfr new_net_7185_bfr_after (
		.din(new_net_7184),
		.dout(new_net_7185)
	);

	bfr new_net_7186_bfr_after (
		.din(new_net_7185),
		.dout(new_net_7186)
	);

	bfr new_net_7187_bfr_after (
		.din(new_net_7186),
		.dout(new_net_7187)
	);

	bfr new_net_7188_bfr_after (
		.din(new_net_7187),
		.dout(new_net_7188)
	);

	bfr new_net_7189_bfr_after (
		.din(new_net_7188),
		.dout(new_net_7189)
	);

	bfr new_net_7190_bfr_after (
		.din(new_net_7189),
		.dout(new_net_7190)
	);

	bfr new_net_7191_bfr_after (
		.din(new_net_7190),
		.dout(new_net_7191)
	);

	bfr new_net_7192_bfr_after (
		.din(new_net_7191),
		.dout(new_net_7192)
	);

	bfr new_net_7193_bfr_after (
		.din(new_net_7192),
		.dout(new_net_7193)
	);

	bfr new_net_7194_bfr_after (
		.din(new_net_7193),
		.dout(new_net_7194)
	);

	bfr new_net_7195_bfr_after (
		.din(new_net_7194),
		.dout(new_net_7195)
	);

	bfr new_net_7196_bfr_after (
		.din(new_net_7195),
		.dout(new_net_7196)
	);

	bfr new_net_7197_bfr_after (
		.din(new_net_7196),
		.dout(new_net_7197)
	);

	bfr new_net_7198_bfr_after (
		.din(new_net_7197),
		.dout(new_net_7198)
	);

	bfr new_net_7199_bfr_after (
		.din(new_net_7198),
		.dout(new_net_7199)
	);

	bfr new_net_7200_bfr_after (
		.din(new_net_7199),
		.dout(new_net_7200)
	);

	bfr new_net_7201_bfr_after (
		.din(new_net_7200),
		.dout(new_net_7201)
	);

	bfr new_net_7202_bfr_after (
		.din(new_net_7201),
		.dout(new_net_7202)
	);

	bfr new_net_7203_bfr_after (
		.din(new_net_7202),
		.dout(new_net_7203)
	);

	bfr new_net_7204_bfr_after (
		.din(new_net_7203),
		.dout(new_net_7204)
	);

	bfr new_net_7205_bfr_after (
		.din(new_net_7204),
		.dout(new_net_7205)
	);

	bfr new_net_7206_bfr_after (
		.din(new_net_7205),
		.dout(new_net_7206)
	);

	bfr new_net_7207_bfr_after (
		.din(new_net_7206),
		.dout(new_net_7207)
	);

	bfr new_net_7208_bfr_after (
		.din(new_net_7207),
		.dout(new_net_7208)
	);

	bfr new_net_7209_bfr_after (
		.din(new_net_7208),
		.dout(new_net_7209)
	);

	bfr new_net_7210_bfr_after (
		.din(new_net_7209),
		.dout(new_net_7210)
	);

	bfr new_net_7211_bfr_after (
		.din(new_net_7210),
		.dout(new_net_7211)
	);

	bfr new_net_7212_bfr_after (
		.din(new_net_7211),
		.dout(new_net_7212)
	);

	bfr new_net_7213_bfr_after (
		.din(new_net_7212),
		.dout(new_net_7213)
	);

	bfr new_net_7214_bfr_after (
		.din(new_net_7213),
		.dout(new_net_7214)
	);

	bfr new_net_7215_bfr_after (
		.din(new_net_7214),
		.dout(new_net_7215)
	);

	bfr new_net_7216_bfr_after (
		.din(new_net_7215),
		.dout(new_net_7216)
	);

	bfr new_net_7217_bfr_after (
		.din(new_net_7216),
		.dout(new_net_7217)
	);

	bfr new_net_7218_bfr_after (
		.din(new_net_7217),
		.dout(new_net_7218)
	);

	bfr new_net_7219_bfr_after (
		.din(new_net_7218),
		.dout(new_net_7219)
	);

	bfr new_net_7220_bfr_after (
		.din(new_net_7219),
		.dout(new_net_7220)
	);

	bfr new_net_7221_bfr_after (
		.din(new_net_7220),
		.dout(new_net_7221)
	);

	bfr new_net_7222_bfr_after (
		.din(new_net_7221),
		.dout(new_net_7222)
	);

	bfr new_net_7223_bfr_after (
		.din(new_net_7222),
		.dout(new_net_7223)
	);

	bfr new_net_7224_bfr_after (
		.din(new_net_7223),
		.dout(new_net_7224)
	);

	bfr new_net_7225_bfr_after (
		.din(new_net_7224),
		.dout(new_net_7225)
	);

	bfr new_net_7226_bfr_after (
		.din(new_net_7225),
		.dout(new_net_7226)
	);

	bfr new_net_7227_bfr_after (
		.din(new_net_7226),
		.dout(new_net_7227)
	);

	bfr new_net_7228_bfr_after (
		.din(new_net_7227),
		.dout(new_net_7228)
	);

	bfr new_net_7229_bfr_after (
		.din(new_net_7228),
		.dout(new_net_7229)
	);

	bfr new_net_7230_bfr_after (
		.din(new_net_7229),
		.dout(new_net_7230)
	);

	bfr new_net_7231_bfr_after (
		.din(new_net_7230),
		.dout(new_net_7231)
	);

	bfr new_net_7232_bfr_after (
		.din(new_net_7231),
		.dout(new_net_7232)
	);

	bfr new_net_7233_bfr_after (
		.din(new_net_7232),
		.dout(new_net_7233)
	);

	bfr new_net_7234_bfr_after (
		.din(new_net_7233),
		.dout(new_net_7234)
	);

	spl2 _0779__v_fanout (
		.a(new_net_7234),
		.b(new_net_2472),
		.c(new_net_2473)
	);

	bfr new_net_7235_bfr_after (
		.din(_1577_),
		.dout(new_net_7235)
	);

	bfr new_net_7236_bfr_after (
		.din(new_net_7235),
		.dout(new_net_7236)
	);

	bfr new_net_7237_bfr_after (
		.din(new_net_7236),
		.dout(new_net_7237)
	);

	bfr new_net_7238_bfr_after (
		.din(new_net_7237),
		.dout(new_net_7238)
	);

	bfr new_net_7239_bfr_after (
		.din(new_net_7238),
		.dout(new_net_7239)
	);

	bfr new_net_7240_bfr_after (
		.din(new_net_7239),
		.dout(new_net_7240)
	);

	bfr new_net_7241_bfr_after (
		.din(new_net_7240),
		.dout(new_net_7241)
	);

	bfr new_net_7242_bfr_after (
		.din(new_net_7241),
		.dout(new_net_7242)
	);

	spl2 _1577__v_fanout (
		.a(new_net_7242),
		.b(new_net_2523),
		.c(new_net_2524)
	);

	bfr new_net_7243_bfr_after (
		.din(_0033_),
		.dout(new_net_7243)
	);

	bfr new_net_7244_bfr_after (
		.din(new_net_7243),
		.dout(new_net_7244)
	);

	bfr new_net_7245_bfr_after (
		.din(new_net_7244),
		.dout(new_net_7245)
	);

	bfr new_net_7246_bfr_after (
		.din(new_net_7245),
		.dout(new_net_7246)
	);

	bfr new_net_7247_bfr_after (
		.din(new_net_7246),
		.dout(new_net_7247)
	);

	bfr new_net_7248_bfr_after (
		.din(new_net_7247),
		.dout(new_net_7248)
	);

	bfr new_net_7249_bfr_after (
		.din(new_net_7248),
		.dout(new_net_7249)
	);

	bfr new_net_7250_bfr_after (
		.din(new_net_7249),
		.dout(new_net_7250)
	);

	spl2 _0033__v_fanout (
		.a(new_net_7250),
		.b(new_net_763),
		.c(new_net_764)
	);

	bfr new_net_7251_bfr_after (
		.din(_1573_),
		.dout(new_net_7251)
	);

	bfr new_net_7252_bfr_after (
		.din(new_net_7251),
		.dout(new_net_7252)
	);

	bfr new_net_7253_bfr_after (
		.din(new_net_7252),
		.dout(new_net_7253)
	);

	bfr new_net_7254_bfr_after (
		.din(new_net_7253),
		.dout(new_net_7254)
	);

	bfr new_net_7255_bfr_after (
		.din(new_net_7254),
		.dout(new_net_7255)
	);

	bfr new_net_7256_bfr_after (
		.din(new_net_7255),
		.dout(new_net_7256)
	);

	bfr new_net_7257_bfr_after (
		.din(new_net_7256),
		.dout(new_net_7257)
	);

	bfr new_net_7258_bfr_after (
		.din(new_net_7257),
		.dout(new_net_7258)
	);

	bfr new_net_7259_bfr_after (
		.din(new_net_7258),
		.dout(new_net_7259)
	);

	bfr new_net_7260_bfr_after (
		.din(new_net_7259),
		.dout(new_net_7260)
	);

	bfr new_net_7261_bfr_after (
		.din(new_net_7260),
		.dout(new_net_7261)
	);

	bfr new_net_7262_bfr_after (
		.din(new_net_7261),
		.dout(new_net_7262)
	);

	bfr new_net_7263_bfr_after (
		.din(new_net_7262),
		.dout(new_net_7263)
	);

	bfr new_net_7264_bfr_after (
		.din(new_net_7263),
		.dout(new_net_7264)
	);

	bfr new_net_7265_bfr_after (
		.din(new_net_7264),
		.dout(new_net_7265)
	);

	bfr new_net_7266_bfr_after (
		.din(new_net_7265),
		.dout(new_net_7266)
	);

	bfr new_net_7267_bfr_after (
		.din(new_net_7266),
		.dout(new_net_7267)
	);

	bfr new_net_7268_bfr_after (
		.din(new_net_7267),
		.dout(new_net_7268)
	);

	bfr new_net_7269_bfr_after (
		.din(new_net_7268),
		.dout(new_net_7269)
	);

	bfr new_net_7270_bfr_after (
		.din(new_net_7269),
		.dout(new_net_7270)
	);

	bfr new_net_7271_bfr_after (
		.din(new_net_7270),
		.dout(new_net_7271)
	);

	bfr new_net_7272_bfr_after (
		.din(new_net_7271),
		.dout(new_net_7272)
	);

	bfr new_net_7273_bfr_after (
		.din(new_net_7272),
		.dout(new_net_7273)
	);

	bfr new_net_7274_bfr_after (
		.din(new_net_7273),
		.dout(new_net_7274)
	);

	bfr new_net_7275_bfr_after (
		.din(new_net_7274),
		.dout(new_net_7275)
	);

	bfr new_net_7276_bfr_after (
		.din(new_net_7275),
		.dout(new_net_7276)
	);

	bfr new_net_7277_bfr_after (
		.din(new_net_7276),
		.dout(new_net_7277)
	);

	bfr new_net_7278_bfr_after (
		.din(new_net_7277),
		.dout(new_net_7278)
	);

	bfr new_net_7279_bfr_after (
		.din(new_net_7278),
		.dout(new_net_7279)
	);

	bfr new_net_7280_bfr_after (
		.din(new_net_7279),
		.dout(new_net_7280)
	);

	bfr new_net_7281_bfr_after (
		.din(new_net_7280),
		.dout(new_net_7281)
	);

	bfr new_net_7282_bfr_after (
		.din(new_net_7281),
		.dout(new_net_7282)
	);

	bfr new_net_7283_bfr_after (
		.din(new_net_7282),
		.dout(new_net_7283)
	);

	bfr new_net_7284_bfr_after (
		.din(new_net_7283),
		.dout(new_net_7284)
	);

	bfr new_net_7285_bfr_after (
		.din(new_net_7284),
		.dout(new_net_7285)
	);

	bfr new_net_7286_bfr_after (
		.din(new_net_7285),
		.dout(new_net_7286)
	);

	bfr new_net_7287_bfr_after (
		.din(new_net_7286),
		.dout(new_net_7287)
	);

	bfr new_net_7288_bfr_after (
		.din(new_net_7287),
		.dout(new_net_7288)
	);

	bfr new_net_7289_bfr_after (
		.din(new_net_7288),
		.dout(new_net_7289)
	);

	bfr new_net_7290_bfr_after (
		.din(new_net_7289),
		.dout(new_net_7290)
	);

	bfr new_net_7291_bfr_after (
		.din(new_net_7290),
		.dout(new_net_7291)
	);

	bfr new_net_7292_bfr_after (
		.din(new_net_7291),
		.dout(new_net_7292)
	);

	bfr new_net_7293_bfr_after (
		.din(new_net_7292),
		.dout(new_net_7293)
	);

	bfr new_net_7294_bfr_after (
		.din(new_net_7293),
		.dout(new_net_7294)
	);

	bfr new_net_7295_bfr_after (
		.din(new_net_7294),
		.dout(new_net_7295)
	);

	bfr new_net_7296_bfr_after (
		.din(new_net_7295),
		.dout(new_net_7296)
	);

	bfr new_net_7297_bfr_after (
		.din(new_net_7296),
		.dout(new_net_7297)
	);

	bfr new_net_7298_bfr_after (
		.din(new_net_7297),
		.dout(new_net_7298)
	);

	bfr new_net_7299_bfr_after (
		.din(new_net_7298),
		.dout(new_net_7299)
	);

	bfr new_net_7300_bfr_after (
		.din(new_net_7299),
		.dout(new_net_7300)
	);

	bfr new_net_7301_bfr_after (
		.din(new_net_7300),
		.dout(new_net_7301)
	);

	bfr new_net_7302_bfr_after (
		.din(new_net_7301),
		.dout(new_net_7302)
	);

	bfr new_net_7303_bfr_after (
		.din(new_net_7302),
		.dout(new_net_7303)
	);

	bfr new_net_7304_bfr_after (
		.din(new_net_7303),
		.dout(new_net_7304)
	);

	bfr new_net_7305_bfr_after (
		.din(new_net_7304),
		.dout(new_net_7305)
	);

	bfr new_net_7306_bfr_after (
		.din(new_net_7305),
		.dout(new_net_7306)
	);

	spl2 _1573__v_fanout (
		.a(new_net_7306),
		.b(new_net_1740),
		.c(new_net_1741)
	);

	bfr new_net_7307_bfr_after (
		.din(_1815_),
		.dout(new_net_7307)
	);

	bfr new_net_7308_bfr_after (
		.din(new_net_7307),
		.dout(new_net_7308)
	);

	bfr new_net_7309_bfr_after (
		.din(new_net_7308),
		.dout(new_net_7309)
	);

	bfr new_net_7310_bfr_after (
		.din(new_net_7309),
		.dout(new_net_7310)
	);

	bfr new_net_7311_bfr_after (
		.din(new_net_7310),
		.dout(new_net_7311)
	);

	bfr new_net_7312_bfr_after (
		.din(new_net_7311),
		.dout(new_net_7312)
	);

	bfr new_net_7313_bfr_after (
		.din(new_net_7312),
		.dout(new_net_7313)
	);

	bfr new_net_7314_bfr_after (
		.din(new_net_7313),
		.dout(new_net_7314)
	);

	bfr new_net_7315_bfr_after (
		.din(new_net_7314),
		.dout(new_net_7315)
	);

	bfr new_net_7316_bfr_after (
		.din(new_net_7315),
		.dout(new_net_7316)
	);

	bfr new_net_7317_bfr_after (
		.din(new_net_7316),
		.dout(new_net_7317)
	);

	bfr new_net_7318_bfr_after (
		.din(new_net_7317),
		.dout(new_net_7318)
	);

	bfr new_net_7319_bfr_after (
		.din(new_net_7318),
		.dout(new_net_7319)
	);

	bfr new_net_7320_bfr_after (
		.din(new_net_7319),
		.dout(new_net_7320)
	);

	bfr new_net_7321_bfr_after (
		.din(new_net_7320),
		.dout(new_net_7321)
	);

	bfr new_net_7322_bfr_after (
		.din(new_net_7321),
		.dout(new_net_7322)
	);

	bfr new_net_7323_bfr_after (
		.din(new_net_7322),
		.dout(new_net_7323)
	);

	bfr new_net_7324_bfr_after (
		.din(new_net_7323),
		.dout(new_net_7324)
	);

	bfr new_net_7325_bfr_after (
		.din(new_net_7324),
		.dout(new_net_7325)
	);

	bfr new_net_7326_bfr_after (
		.din(new_net_7325),
		.dout(new_net_7326)
	);

	bfr new_net_7327_bfr_after (
		.din(new_net_7326),
		.dout(new_net_7327)
	);

	bfr new_net_7328_bfr_after (
		.din(new_net_7327),
		.dout(new_net_7328)
	);

	bfr new_net_7329_bfr_after (
		.din(new_net_7328),
		.dout(new_net_7329)
	);

	bfr new_net_7330_bfr_after (
		.din(new_net_7329),
		.dout(new_net_7330)
	);

	bfr new_net_7331_bfr_after (
		.din(new_net_7330),
		.dout(new_net_7331)
	);

	bfr new_net_7332_bfr_after (
		.din(new_net_7331),
		.dout(new_net_7332)
	);

	bfr new_net_7333_bfr_after (
		.din(new_net_7332),
		.dout(new_net_7333)
	);

	bfr new_net_7334_bfr_after (
		.din(new_net_7333),
		.dout(new_net_7334)
	);

	bfr new_net_7335_bfr_after (
		.din(new_net_7334),
		.dout(new_net_7335)
	);

	bfr new_net_7336_bfr_after (
		.din(new_net_7335),
		.dout(new_net_7336)
	);

	bfr new_net_7337_bfr_after (
		.din(new_net_7336),
		.dout(new_net_7337)
	);

	bfr new_net_7338_bfr_after (
		.din(new_net_7337),
		.dout(new_net_7338)
	);

	bfr new_net_7339_bfr_after (
		.din(new_net_7338),
		.dout(new_net_7339)
	);

	bfr new_net_7340_bfr_after (
		.din(new_net_7339),
		.dout(new_net_7340)
	);

	bfr new_net_7341_bfr_after (
		.din(new_net_7340),
		.dout(new_net_7341)
	);

	bfr new_net_7342_bfr_after (
		.din(new_net_7341),
		.dout(new_net_7342)
	);

	bfr new_net_7343_bfr_after (
		.din(new_net_7342),
		.dout(new_net_7343)
	);

	bfr new_net_7344_bfr_after (
		.din(new_net_7343),
		.dout(new_net_7344)
	);

	bfr new_net_7345_bfr_after (
		.din(new_net_7344),
		.dout(new_net_7345)
	);

	bfr new_net_7346_bfr_after (
		.din(new_net_7345),
		.dout(new_net_7346)
	);

	bfr new_net_7347_bfr_after (
		.din(new_net_7346),
		.dout(new_net_7347)
	);

	bfr new_net_7348_bfr_after (
		.din(new_net_7347),
		.dout(new_net_7348)
	);

	bfr new_net_7349_bfr_after (
		.din(new_net_7348),
		.dout(new_net_7349)
	);

	bfr new_net_7350_bfr_after (
		.din(new_net_7349),
		.dout(new_net_7350)
	);

	bfr new_net_7351_bfr_after (
		.din(new_net_7350),
		.dout(new_net_7351)
	);

	bfr new_net_7352_bfr_after (
		.din(new_net_7351),
		.dout(new_net_7352)
	);

	bfr new_net_7353_bfr_after (
		.din(new_net_7352),
		.dout(new_net_7353)
	);

	bfr new_net_7354_bfr_after (
		.din(new_net_7353),
		.dout(new_net_7354)
	);

	bfr new_net_7355_bfr_after (
		.din(new_net_7354),
		.dout(new_net_7355)
	);

	bfr new_net_7356_bfr_after (
		.din(new_net_7355),
		.dout(new_net_7356)
	);

	bfr new_net_7357_bfr_after (
		.din(new_net_7356),
		.dout(new_net_7357)
	);

	bfr new_net_7358_bfr_after (
		.din(new_net_7357),
		.dout(new_net_7358)
	);

	bfr new_net_7359_bfr_after (
		.din(new_net_7358),
		.dout(new_net_7359)
	);

	bfr new_net_7360_bfr_after (
		.din(new_net_7359),
		.dout(new_net_7360)
	);

	bfr new_net_7361_bfr_after (
		.din(new_net_7360),
		.dout(new_net_7361)
	);

	bfr new_net_7362_bfr_after (
		.din(new_net_7361),
		.dout(new_net_7362)
	);

	bfr new_net_7363_bfr_after (
		.din(new_net_7362),
		.dout(new_net_7363)
	);

	bfr new_net_7364_bfr_after (
		.din(new_net_7363),
		.dout(new_net_7364)
	);

	bfr new_net_7365_bfr_after (
		.din(new_net_7364),
		.dout(new_net_7365)
	);

	bfr new_net_7366_bfr_after (
		.din(new_net_7365),
		.dout(new_net_7366)
	);

	bfr new_net_7367_bfr_after (
		.din(new_net_7366),
		.dout(new_net_7367)
	);

	bfr new_net_7368_bfr_after (
		.din(new_net_7367),
		.dout(new_net_7368)
	);

	bfr new_net_7369_bfr_after (
		.din(new_net_7368),
		.dout(new_net_7369)
	);

	bfr new_net_7370_bfr_after (
		.din(new_net_7369),
		.dout(new_net_7370)
	);

	spl2 _1815__v_fanout (
		.a(new_net_7370),
		.b(new_net_982),
		.c(new_net_983)
	);

	bfr new_net_7371_bfr_after (
		.din(_0963_),
		.dout(new_net_7371)
	);

	bfr new_net_7372_bfr_after (
		.din(new_net_7371),
		.dout(new_net_7372)
	);

	bfr new_net_7373_bfr_after (
		.din(new_net_7372),
		.dout(new_net_7373)
	);

	bfr new_net_7374_bfr_after (
		.din(new_net_7373),
		.dout(new_net_7374)
	);

	bfr new_net_7375_bfr_after (
		.din(new_net_7374),
		.dout(new_net_7375)
	);

	bfr new_net_7376_bfr_after (
		.din(new_net_7375),
		.dout(new_net_7376)
	);

	bfr new_net_7377_bfr_after (
		.din(new_net_7376),
		.dout(new_net_7377)
	);

	bfr new_net_7378_bfr_after (
		.din(new_net_7377),
		.dout(new_net_7378)
	);

	bfr new_net_7379_bfr_after (
		.din(new_net_7378),
		.dout(new_net_7379)
	);

	bfr new_net_7380_bfr_after (
		.din(new_net_7379),
		.dout(new_net_7380)
	);

	bfr new_net_7381_bfr_after (
		.din(new_net_7380),
		.dout(new_net_7381)
	);

	bfr new_net_7382_bfr_after (
		.din(new_net_7381),
		.dout(new_net_7382)
	);

	bfr new_net_7383_bfr_after (
		.din(new_net_7382),
		.dout(new_net_7383)
	);

	bfr new_net_7384_bfr_after (
		.din(new_net_7383),
		.dout(new_net_7384)
	);

	bfr new_net_7385_bfr_after (
		.din(new_net_7384),
		.dout(new_net_7385)
	);

	bfr new_net_7386_bfr_after (
		.din(new_net_7385),
		.dout(new_net_7386)
	);

	bfr new_net_7387_bfr_after (
		.din(new_net_7386),
		.dout(new_net_7387)
	);

	bfr new_net_7388_bfr_after (
		.din(new_net_7387),
		.dout(new_net_7388)
	);

	bfr new_net_7389_bfr_after (
		.din(new_net_7388),
		.dout(new_net_7389)
	);

	bfr new_net_7390_bfr_after (
		.din(new_net_7389),
		.dout(new_net_7390)
	);

	bfr new_net_7391_bfr_after (
		.din(new_net_7390),
		.dout(new_net_7391)
	);

	bfr new_net_7392_bfr_after (
		.din(new_net_7391),
		.dout(new_net_7392)
	);

	bfr new_net_7393_bfr_after (
		.din(new_net_7392),
		.dout(new_net_7393)
	);

	bfr new_net_7394_bfr_after (
		.din(new_net_7393),
		.dout(new_net_7394)
	);

	bfr new_net_7395_bfr_after (
		.din(new_net_7394),
		.dout(new_net_7395)
	);

	bfr new_net_7396_bfr_after (
		.din(new_net_7395),
		.dout(new_net_7396)
	);

	bfr new_net_7397_bfr_after (
		.din(new_net_7396),
		.dout(new_net_7397)
	);

	bfr new_net_7398_bfr_after (
		.din(new_net_7397),
		.dout(new_net_7398)
	);

	bfr new_net_7399_bfr_after (
		.din(new_net_7398),
		.dout(new_net_7399)
	);

	bfr new_net_7400_bfr_after (
		.din(new_net_7399),
		.dout(new_net_7400)
	);

	bfr new_net_7401_bfr_after (
		.din(new_net_7400),
		.dout(new_net_7401)
	);

	bfr new_net_7402_bfr_after (
		.din(new_net_7401),
		.dout(new_net_7402)
	);

	bfr new_net_7403_bfr_after (
		.din(new_net_7402),
		.dout(new_net_7403)
	);

	bfr new_net_7404_bfr_after (
		.din(new_net_7403),
		.dout(new_net_7404)
	);

	bfr new_net_7405_bfr_after (
		.din(new_net_7404),
		.dout(new_net_7405)
	);

	bfr new_net_7406_bfr_after (
		.din(new_net_7405),
		.dout(new_net_7406)
	);

	bfr new_net_7407_bfr_after (
		.din(new_net_7406),
		.dout(new_net_7407)
	);

	bfr new_net_7408_bfr_after (
		.din(new_net_7407),
		.dout(new_net_7408)
	);

	bfr new_net_7409_bfr_after (
		.din(new_net_7408),
		.dout(new_net_7409)
	);

	bfr new_net_7410_bfr_after (
		.din(new_net_7409),
		.dout(new_net_7410)
	);

	bfr new_net_7411_bfr_after (
		.din(new_net_7410),
		.dout(new_net_7411)
	);

	bfr new_net_7412_bfr_after (
		.din(new_net_7411),
		.dout(new_net_7412)
	);

	bfr new_net_7413_bfr_after (
		.din(new_net_7412),
		.dout(new_net_7413)
	);

	bfr new_net_7414_bfr_after (
		.din(new_net_7413),
		.dout(new_net_7414)
	);

	bfr new_net_7415_bfr_after (
		.din(new_net_7414),
		.dout(new_net_7415)
	);

	bfr new_net_7416_bfr_after (
		.din(new_net_7415),
		.dout(new_net_7416)
	);

	bfr new_net_7417_bfr_after (
		.din(new_net_7416),
		.dout(new_net_7417)
	);

	bfr new_net_7418_bfr_after (
		.din(new_net_7417),
		.dout(new_net_7418)
	);

	bfr new_net_7419_bfr_after (
		.din(new_net_7418),
		.dout(new_net_7419)
	);

	bfr new_net_7420_bfr_after (
		.din(new_net_7419),
		.dout(new_net_7420)
	);

	bfr new_net_7421_bfr_after (
		.din(new_net_7420),
		.dout(new_net_7421)
	);

	bfr new_net_7422_bfr_after (
		.din(new_net_7421),
		.dout(new_net_7422)
	);

	bfr new_net_7423_bfr_after (
		.din(new_net_7422),
		.dout(new_net_7423)
	);

	bfr new_net_7424_bfr_after (
		.din(new_net_7423),
		.dout(new_net_7424)
	);

	bfr new_net_7425_bfr_after (
		.din(new_net_7424),
		.dout(new_net_7425)
	);

	bfr new_net_7426_bfr_after (
		.din(new_net_7425),
		.dout(new_net_7426)
	);

	bfr new_net_7427_bfr_after (
		.din(new_net_7426),
		.dout(new_net_7427)
	);

	bfr new_net_7428_bfr_after (
		.din(new_net_7427),
		.dout(new_net_7428)
	);

	bfr new_net_7429_bfr_after (
		.din(new_net_7428),
		.dout(new_net_7429)
	);

	bfr new_net_7430_bfr_after (
		.din(new_net_7429),
		.dout(new_net_7430)
	);

	bfr new_net_7431_bfr_after (
		.din(new_net_7430),
		.dout(new_net_7431)
	);

	bfr new_net_7432_bfr_after (
		.din(new_net_7431),
		.dout(new_net_7432)
	);

	bfr new_net_7433_bfr_after (
		.din(new_net_7432),
		.dout(new_net_7433)
	);

	bfr new_net_7434_bfr_after (
		.din(new_net_7433),
		.dout(new_net_7434)
	);

	bfr new_net_7435_bfr_after (
		.din(new_net_7434),
		.dout(new_net_7435)
	);

	bfr new_net_7436_bfr_after (
		.din(new_net_7435),
		.dout(new_net_7436)
	);

	bfr new_net_7437_bfr_after (
		.din(new_net_7436),
		.dout(new_net_7437)
	);

	bfr new_net_7438_bfr_after (
		.din(new_net_7437),
		.dout(new_net_7438)
	);

	bfr new_net_7439_bfr_after (
		.din(new_net_7438),
		.dout(new_net_7439)
	);

	bfr new_net_7440_bfr_after (
		.din(new_net_7439),
		.dout(new_net_7440)
	);

	bfr new_net_7441_bfr_after (
		.din(new_net_7440),
		.dout(new_net_7441)
	);

	bfr new_net_7442_bfr_after (
		.din(new_net_7441),
		.dout(new_net_7442)
	);

	bfr new_net_7443_bfr_after (
		.din(new_net_7442),
		.dout(new_net_7443)
	);

	bfr new_net_7444_bfr_after (
		.din(new_net_7443),
		.dout(new_net_7444)
	);

	bfr new_net_7445_bfr_after (
		.din(new_net_7444),
		.dout(new_net_7445)
	);

	bfr new_net_7446_bfr_after (
		.din(new_net_7445),
		.dout(new_net_7446)
	);

	bfr new_net_7447_bfr_after (
		.din(new_net_7446),
		.dout(new_net_7447)
	);

	bfr new_net_7448_bfr_after (
		.din(new_net_7447),
		.dout(new_net_7448)
	);

	bfr new_net_7449_bfr_after (
		.din(new_net_7448),
		.dout(new_net_7449)
	);

	bfr new_net_7450_bfr_after (
		.din(new_net_7449),
		.dout(new_net_7450)
	);

	bfr new_net_7451_bfr_after (
		.din(new_net_7450),
		.dout(new_net_7451)
	);

	bfr new_net_7452_bfr_after (
		.din(new_net_7451),
		.dout(new_net_7452)
	);

	bfr new_net_7453_bfr_after (
		.din(new_net_7452),
		.dout(new_net_7453)
	);

	bfr new_net_7454_bfr_after (
		.din(new_net_7453),
		.dout(new_net_7454)
	);

	bfr new_net_7455_bfr_after (
		.din(new_net_7454),
		.dout(new_net_7455)
	);

	bfr new_net_7456_bfr_after (
		.din(new_net_7455),
		.dout(new_net_7456)
	);

	bfr new_net_7457_bfr_after (
		.din(new_net_7456),
		.dout(new_net_7457)
	);

	bfr new_net_7458_bfr_after (
		.din(new_net_7457),
		.dout(new_net_7458)
	);

	bfr new_net_7459_bfr_after (
		.din(new_net_7458),
		.dout(new_net_7459)
	);

	bfr new_net_7460_bfr_after (
		.din(new_net_7459),
		.dout(new_net_7460)
	);

	bfr new_net_7461_bfr_after (
		.din(new_net_7460),
		.dout(new_net_7461)
	);

	bfr new_net_7462_bfr_after (
		.din(new_net_7461),
		.dout(new_net_7462)
	);

	bfr new_net_7463_bfr_after (
		.din(new_net_7462),
		.dout(new_net_7463)
	);

	bfr new_net_7464_bfr_after (
		.din(new_net_7463),
		.dout(new_net_7464)
	);

	bfr new_net_7465_bfr_after (
		.din(new_net_7464),
		.dout(new_net_7465)
	);

	bfr new_net_7466_bfr_after (
		.din(new_net_7465),
		.dout(new_net_7466)
	);

	bfr new_net_7467_bfr_after (
		.din(new_net_7466),
		.dout(new_net_7467)
	);

	bfr new_net_7468_bfr_after (
		.din(new_net_7467),
		.dout(new_net_7468)
	);

	spl2 _0963__v_fanout (
		.a(new_net_7468),
		.b(new_net_3266),
		.c(new_net_3267)
	);

	bfr new_net_7469_bfr_after (
		.din(_0621_),
		.dout(new_net_7469)
	);

	bfr new_net_7470_bfr_after (
		.din(new_net_7469),
		.dout(new_net_7470)
	);

	bfr new_net_7471_bfr_after (
		.din(new_net_7470),
		.dout(new_net_7471)
	);

	bfr new_net_7472_bfr_after (
		.din(new_net_7471),
		.dout(new_net_7472)
	);

	bfr new_net_7473_bfr_after (
		.din(new_net_7472),
		.dout(new_net_7473)
	);

	bfr new_net_7474_bfr_after (
		.din(new_net_7473),
		.dout(new_net_7474)
	);

	bfr new_net_7475_bfr_after (
		.din(new_net_7474),
		.dout(new_net_7475)
	);

	bfr new_net_7476_bfr_after (
		.din(new_net_7475),
		.dout(new_net_7476)
	);

	bfr new_net_7477_bfr_after (
		.din(new_net_7476),
		.dout(new_net_7477)
	);

	bfr new_net_7478_bfr_after (
		.din(new_net_7477),
		.dout(new_net_7478)
	);

	bfr new_net_7479_bfr_after (
		.din(new_net_7478),
		.dout(new_net_7479)
	);

	bfr new_net_7480_bfr_after (
		.din(new_net_7479),
		.dout(new_net_7480)
	);

	bfr new_net_7481_bfr_after (
		.din(new_net_7480),
		.dout(new_net_7481)
	);

	bfr new_net_7482_bfr_after (
		.din(new_net_7481),
		.dout(new_net_7482)
	);

	bfr new_net_7483_bfr_after (
		.din(new_net_7482),
		.dout(new_net_7483)
	);

	bfr new_net_7484_bfr_after (
		.din(new_net_7483),
		.dout(new_net_7484)
	);

	bfr new_net_7485_bfr_after (
		.din(new_net_7484),
		.dout(new_net_7485)
	);

	bfr new_net_7486_bfr_after (
		.din(new_net_7485),
		.dout(new_net_7486)
	);

	bfr new_net_7487_bfr_after (
		.din(new_net_7486),
		.dout(new_net_7487)
	);

	bfr new_net_7488_bfr_after (
		.din(new_net_7487),
		.dout(new_net_7488)
	);

	bfr new_net_7489_bfr_after (
		.din(new_net_7488),
		.dout(new_net_7489)
	);

	bfr new_net_7490_bfr_after (
		.din(new_net_7489),
		.dout(new_net_7490)
	);

	bfr new_net_7491_bfr_after (
		.din(new_net_7490),
		.dout(new_net_7491)
	);

	bfr new_net_7492_bfr_after (
		.din(new_net_7491),
		.dout(new_net_7492)
	);

	bfr new_net_7493_bfr_after (
		.din(new_net_7492),
		.dout(new_net_7493)
	);

	bfr new_net_7494_bfr_after (
		.din(new_net_7493),
		.dout(new_net_7494)
	);

	bfr new_net_7495_bfr_after (
		.din(new_net_7494),
		.dout(new_net_7495)
	);

	bfr new_net_7496_bfr_after (
		.din(new_net_7495),
		.dout(new_net_7496)
	);

	bfr new_net_7497_bfr_after (
		.din(new_net_7496),
		.dout(new_net_7497)
	);

	bfr new_net_7498_bfr_after (
		.din(new_net_7497),
		.dout(new_net_7498)
	);

	bfr new_net_7499_bfr_after (
		.din(new_net_7498),
		.dout(new_net_7499)
	);

	bfr new_net_7500_bfr_after (
		.din(new_net_7499),
		.dout(new_net_7500)
	);

	bfr new_net_7501_bfr_after (
		.din(new_net_7500),
		.dout(new_net_7501)
	);

	bfr new_net_7502_bfr_after (
		.din(new_net_7501),
		.dout(new_net_7502)
	);

	bfr new_net_7503_bfr_after (
		.din(new_net_7502),
		.dout(new_net_7503)
	);

	bfr new_net_7504_bfr_after (
		.din(new_net_7503),
		.dout(new_net_7504)
	);

	bfr new_net_7505_bfr_after (
		.din(new_net_7504),
		.dout(new_net_7505)
	);

	bfr new_net_7506_bfr_after (
		.din(new_net_7505),
		.dout(new_net_7506)
	);

	bfr new_net_7507_bfr_after (
		.din(new_net_7506),
		.dout(new_net_7507)
	);

	bfr new_net_7508_bfr_after (
		.din(new_net_7507),
		.dout(new_net_7508)
	);

	bfr new_net_7509_bfr_after (
		.din(new_net_7508),
		.dout(new_net_7509)
	);

	bfr new_net_7510_bfr_after (
		.din(new_net_7509),
		.dout(new_net_7510)
	);

	bfr new_net_7511_bfr_after (
		.din(new_net_7510),
		.dout(new_net_7511)
	);

	bfr new_net_7512_bfr_after (
		.din(new_net_7511),
		.dout(new_net_7512)
	);

	bfr new_net_7513_bfr_after (
		.din(new_net_7512),
		.dout(new_net_7513)
	);

	bfr new_net_7514_bfr_after (
		.din(new_net_7513),
		.dout(new_net_7514)
	);

	bfr new_net_7515_bfr_after (
		.din(new_net_7514),
		.dout(new_net_7515)
	);

	bfr new_net_7516_bfr_after (
		.din(new_net_7515),
		.dout(new_net_7516)
	);

	bfr new_net_7517_bfr_after (
		.din(new_net_7516),
		.dout(new_net_7517)
	);

	bfr new_net_7518_bfr_after (
		.din(new_net_7517),
		.dout(new_net_7518)
	);

	bfr new_net_7519_bfr_after (
		.din(new_net_7518),
		.dout(new_net_7519)
	);

	bfr new_net_7520_bfr_after (
		.din(new_net_7519),
		.dout(new_net_7520)
	);

	bfr new_net_7521_bfr_after (
		.din(new_net_7520),
		.dout(new_net_7521)
	);

	bfr new_net_7522_bfr_after (
		.din(new_net_7521),
		.dout(new_net_7522)
	);

	bfr new_net_7523_bfr_after (
		.din(new_net_7522),
		.dout(new_net_7523)
	);

	bfr new_net_7524_bfr_after (
		.din(new_net_7523),
		.dout(new_net_7524)
	);

	bfr new_net_7525_bfr_after (
		.din(new_net_7524),
		.dout(new_net_7525)
	);

	bfr new_net_7526_bfr_after (
		.din(new_net_7525),
		.dout(new_net_7526)
	);

	bfr new_net_7527_bfr_after (
		.din(new_net_7526),
		.dout(new_net_7527)
	);

	bfr new_net_7528_bfr_after (
		.din(new_net_7527),
		.dout(new_net_7528)
	);

	bfr new_net_7529_bfr_after (
		.din(new_net_7528),
		.dout(new_net_7529)
	);

	bfr new_net_7530_bfr_after (
		.din(new_net_7529),
		.dout(new_net_7530)
	);

	bfr new_net_7531_bfr_after (
		.din(new_net_7530),
		.dout(new_net_7531)
	);

	bfr new_net_7532_bfr_after (
		.din(new_net_7531),
		.dout(new_net_7532)
	);

	bfr new_net_7533_bfr_after (
		.din(new_net_7532),
		.dout(new_net_7533)
	);

	bfr new_net_7534_bfr_after (
		.din(new_net_7533),
		.dout(new_net_7534)
	);

	bfr new_net_7535_bfr_after (
		.din(new_net_7534),
		.dout(new_net_7535)
	);

	bfr new_net_7536_bfr_after (
		.din(new_net_7535),
		.dout(new_net_7536)
	);

	bfr new_net_7537_bfr_after (
		.din(new_net_7536),
		.dout(new_net_7537)
	);

	bfr new_net_7538_bfr_after (
		.din(new_net_7537),
		.dout(new_net_7538)
	);

	bfr new_net_7539_bfr_after (
		.din(new_net_7538),
		.dout(new_net_7539)
	);

	bfr new_net_7540_bfr_after (
		.din(new_net_7539),
		.dout(new_net_7540)
	);

	bfr new_net_7541_bfr_after (
		.din(new_net_7540),
		.dout(new_net_7541)
	);

	bfr new_net_7542_bfr_after (
		.din(new_net_7541),
		.dout(new_net_7542)
	);

	bfr new_net_7543_bfr_after (
		.din(new_net_7542),
		.dout(new_net_7543)
	);

	bfr new_net_7544_bfr_after (
		.din(new_net_7543),
		.dout(new_net_7544)
	);

	bfr new_net_7545_bfr_after (
		.din(new_net_7544),
		.dout(new_net_7545)
	);

	bfr new_net_7546_bfr_after (
		.din(new_net_7545),
		.dout(new_net_7546)
	);

	bfr new_net_7547_bfr_after (
		.din(new_net_7546),
		.dout(new_net_7547)
	);

	bfr new_net_7548_bfr_after (
		.din(new_net_7547),
		.dout(new_net_7548)
	);

	bfr new_net_7549_bfr_after (
		.din(new_net_7548),
		.dout(new_net_7549)
	);

	bfr new_net_7550_bfr_after (
		.din(new_net_7549),
		.dout(new_net_7550)
	);

	bfr new_net_7551_bfr_after (
		.din(new_net_7550),
		.dout(new_net_7551)
	);

	bfr new_net_7552_bfr_after (
		.din(new_net_7551),
		.dout(new_net_7552)
	);

	bfr new_net_7553_bfr_after (
		.din(new_net_7552),
		.dout(new_net_7553)
	);

	bfr new_net_7554_bfr_after (
		.din(new_net_7553),
		.dout(new_net_7554)
	);

	bfr new_net_7555_bfr_after (
		.din(new_net_7554),
		.dout(new_net_7555)
	);

	bfr new_net_7556_bfr_after (
		.din(new_net_7555),
		.dout(new_net_7556)
	);

	bfr new_net_7557_bfr_after (
		.din(new_net_7556),
		.dout(new_net_7557)
	);

	bfr new_net_7558_bfr_after (
		.din(new_net_7557),
		.dout(new_net_7558)
	);

	bfr new_net_7559_bfr_after (
		.din(new_net_7558),
		.dout(new_net_7559)
	);

	bfr new_net_7560_bfr_after (
		.din(new_net_7559),
		.dout(new_net_7560)
	);

	bfr new_net_7561_bfr_after (
		.din(new_net_7560),
		.dout(new_net_7561)
	);

	bfr new_net_7562_bfr_after (
		.din(new_net_7561),
		.dout(new_net_7562)
	);

	bfr new_net_7563_bfr_after (
		.din(new_net_7562),
		.dout(new_net_7563)
	);

	bfr new_net_7564_bfr_after (
		.din(new_net_7563),
		.dout(new_net_7564)
	);

	spl2 _0621__v_fanout (
		.a(new_net_7564),
		.b(new_net_767),
		.c(new_net_768)
	);

	bfr new_net_7565_bfr_after (
		.din(_0091_),
		.dout(new_net_7565)
	);

	bfr new_net_7566_bfr_after (
		.din(new_net_7565),
		.dout(new_net_7566)
	);

	bfr new_net_7567_bfr_after (
		.din(new_net_7566),
		.dout(new_net_7567)
	);

	bfr new_net_7568_bfr_after (
		.din(new_net_7567),
		.dout(new_net_7568)
	);

	bfr new_net_7569_bfr_after (
		.din(new_net_7568),
		.dout(new_net_7569)
	);

	bfr new_net_7570_bfr_after (
		.din(new_net_7569),
		.dout(new_net_7570)
	);

	bfr new_net_7571_bfr_after (
		.din(new_net_7570),
		.dout(new_net_7571)
	);

	bfr new_net_7572_bfr_after (
		.din(new_net_7571),
		.dout(new_net_7572)
	);

	bfr new_net_7573_bfr_after (
		.din(new_net_7572),
		.dout(new_net_7573)
	);

	bfr new_net_7574_bfr_after (
		.din(new_net_7573),
		.dout(new_net_7574)
	);

	bfr new_net_7575_bfr_after (
		.din(new_net_7574),
		.dout(new_net_7575)
	);

	bfr new_net_7576_bfr_after (
		.din(new_net_7575),
		.dout(new_net_7576)
	);

	bfr new_net_7577_bfr_after (
		.din(new_net_7576),
		.dout(new_net_7577)
	);

	bfr new_net_7578_bfr_after (
		.din(new_net_7577),
		.dout(new_net_7578)
	);

	bfr new_net_7579_bfr_after (
		.din(new_net_7578),
		.dout(new_net_7579)
	);

	bfr new_net_7580_bfr_after (
		.din(new_net_7579),
		.dout(new_net_7580)
	);

	bfr new_net_7581_bfr_after (
		.din(new_net_7580),
		.dout(new_net_7581)
	);

	bfr new_net_7582_bfr_after (
		.din(new_net_7581),
		.dout(new_net_7582)
	);

	bfr new_net_7583_bfr_after (
		.din(new_net_7582),
		.dout(new_net_7583)
	);

	bfr new_net_7584_bfr_after (
		.din(new_net_7583),
		.dout(new_net_7584)
	);

	bfr new_net_7585_bfr_after (
		.din(new_net_7584),
		.dout(new_net_7585)
	);

	bfr new_net_7586_bfr_after (
		.din(new_net_7585),
		.dout(new_net_7586)
	);

	bfr new_net_7587_bfr_after (
		.din(new_net_7586),
		.dout(new_net_7587)
	);

	bfr new_net_7588_bfr_after (
		.din(new_net_7587),
		.dout(new_net_7588)
	);

	bfr new_net_7589_bfr_after (
		.din(new_net_7588),
		.dout(new_net_7589)
	);

	bfr new_net_7590_bfr_after (
		.din(new_net_7589),
		.dout(new_net_7590)
	);

	bfr new_net_7591_bfr_after (
		.din(new_net_7590),
		.dout(new_net_7591)
	);

	bfr new_net_7592_bfr_after (
		.din(new_net_7591),
		.dout(new_net_7592)
	);

	bfr new_net_7593_bfr_after (
		.din(new_net_7592),
		.dout(new_net_7593)
	);

	bfr new_net_7594_bfr_after (
		.din(new_net_7593),
		.dout(new_net_7594)
	);

	bfr new_net_7595_bfr_after (
		.din(new_net_7594),
		.dout(new_net_7595)
	);

	bfr new_net_7596_bfr_after (
		.din(new_net_7595),
		.dout(new_net_7596)
	);

	bfr new_net_7597_bfr_after (
		.din(new_net_7596),
		.dout(new_net_7597)
	);

	bfr new_net_7598_bfr_after (
		.din(new_net_7597),
		.dout(new_net_7598)
	);

	bfr new_net_7599_bfr_after (
		.din(new_net_7598),
		.dout(new_net_7599)
	);

	bfr new_net_7600_bfr_after (
		.din(new_net_7599),
		.dout(new_net_7600)
	);

	bfr new_net_7601_bfr_after (
		.din(new_net_7600),
		.dout(new_net_7601)
	);

	bfr new_net_7602_bfr_after (
		.din(new_net_7601),
		.dout(new_net_7602)
	);

	bfr new_net_7603_bfr_after (
		.din(new_net_7602),
		.dout(new_net_7603)
	);

	bfr new_net_7604_bfr_after (
		.din(new_net_7603),
		.dout(new_net_7604)
	);

	bfr new_net_7605_bfr_after (
		.din(new_net_7604),
		.dout(new_net_7605)
	);

	bfr new_net_7606_bfr_after (
		.din(new_net_7605),
		.dout(new_net_7606)
	);

	bfr new_net_7607_bfr_after (
		.din(new_net_7606),
		.dout(new_net_7607)
	);

	bfr new_net_7608_bfr_after (
		.din(new_net_7607),
		.dout(new_net_7608)
	);

	bfr new_net_7609_bfr_after (
		.din(new_net_7608),
		.dout(new_net_7609)
	);

	bfr new_net_7610_bfr_after (
		.din(new_net_7609),
		.dout(new_net_7610)
	);

	bfr new_net_7611_bfr_after (
		.din(new_net_7610),
		.dout(new_net_7611)
	);

	bfr new_net_7612_bfr_after (
		.din(new_net_7611),
		.dout(new_net_7612)
	);

	bfr new_net_7613_bfr_after (
		.din(new_net_7612),
		.dout(new_net_7613)
	);

	bfr new_net_7614_bfr_after (
		.din(new_net_7613),
		.dout(new_net_7614)
	);

	bfr new_net_7615_bfr_after (
		.din(new_net_7614),
		.dout(new_net_7615)
	);

	bfr new_net_7616_bfr_after (
		.din(new_net_7615),
		.dout(new_net_7616)
	);

	bfr new_net_7617_bfr_after (
		.din(new_net_7616),
		.dout(new_net_7617)
	);

	bfr new_net_7618_bfr_after (
		.din(new_net_7617),
		.dout(new_net_7618)
	);

	bfr new_net_7619_bfr_after (
		.din(new_net_7618),
		.dout(new_net_7619)
	);

	bfr new_net_7620_bfr_after (
		.din(new_net_7619),
		.dout(new_net_7620)
	);

	bfr new_net_7621_bfr_after (
		.din(new_net_7620),
		.dout(new_net_7621)
	);

	bfr new_net_7622_bfr_after (
		.din(new_net_7621),
		.dout(new_net_7622)
	);

	bfr new_net_7623_bfr_after (
		.din(new_net_7622),
		.dout(new_net_7623)
	);

	bfr new_net_7624_bfr_after (
		.din(new_net_7623),
		.dout(new_net_7624)
	);

	bfr new_net_7625_bfr_after (
		.din(new_net_7624),
		.dout(new_net_7625)
	);

	bfr new_net_7626_bfr_after (
		.din(new_net_7625),
		.dout(new_net_7626)
	);

	bfr new_net_7627_bfr_after (
		.din(new_net_7626),
		.dout(new_net_7627)
	);

	bfr new_net_7628_bfr_after (
		.din(new_net_7627),
		.dout(new_net_7628)
	);

	bfr new_net_7629_bfr_after (
		.din(new_net_7628),
		.dout(new_net_7629)
	);

	bfr new_net_7630_bfr_after (
		.din(new_net_7629),
		.dout(new_net_7630)
	);

	bfr new_net_7631_bfr_after (
		.din(new_net_7630),
		.dout(new_net_7631)
	);

	bfr new_net_7632_bfr_after (
		.din(new_net_7631),
		.dout(new_net_7632)
	);

	bfr new_net_7633_bfr_after (
		.din(new_net_7632),
		.dout(new_net_7633)
	);

	bfr new_net_7634_bfr_after (
		.din(new_net_7633),
		.dout(new_net_7634)
	);

	bfr new_net_7635_bfr_after (
		.din(new_net_7634),
		.dout(new_net_7635)
	);

	bfr new_net_7636_bfr_after (
		.din(new_net_7635),
		.dout(new_net_7636)
	);

	bfr new_net_7637_bfr_after (
		.din(new_net_7636),
		.dout(new_net_7637)
	);

	bfr new_net_7638_bfr_after (
		.din(new_net_7637),
		.dout(new_net_7638)
	);

	bfr new_net_7639_bfr_after (
		.din(new_net_7638),
		.dout(new_net_7639)
	);

	bfr new_net_7640_bfr_after (
		.din(new_net_7639),
		.dout(new_net_7640)
	);

	bfr new_net_7641_bfr_after (
		.din(new_net_7640),
		.dout(new_net_7641)
	);

	bfr new_net_7642_bfr_after (
		.din(new_net_7641),
		.dout(new_net_7642)
	);

	bfr new_net_7643_bfr_after (
		.din(new_net_7642),
		.dout(new_net_7643)
	);

	bfr new_net_7644_bfr_after (
		.din(new_net_7643),
		.dout(new_net_7644)
	);

	bfr new_net_7645_bfr_after (
		.din(new_net_7644),
		.dout(new_net_7645)
	);

	bfr new_net_7646_bfr_after (
		.din(new_net_7645),
		.dout(new_net_7646)
	);

	bfr new_net_7647_bfr_after (
		.din(new_net_7646),
		.dout(new_net_7647)
	);

	bfr new_net_7648_bfr_after (
		.din(new_net_7647),
		.dout(new_net_7648)
	);

	bfr new_net_7649_bfr_after (
		.din(new_net_7648),
		.dout(new_net_7649)
	);

	bfr new_net_7650_bfr_after (
		.din(new_net_7649),
		.dout(new_net_7650)
	);

	bfr new_net_7651_bfr_after (
		.din(new_net_7650),
		.dout(new_net_7651)
	);

	bfr new_net_7652_bfr_after (
		.din(new_net_7651),
		.dout(new_net_7652)
	);

	spl2 _0091__v_fanout (
		.a(new_net_7652),
		.b(new_net_3222),
		.c(new_net_3223)
	);

	bfr new_net_7653_bfr_after (
		.din(_1813_),
		.dout(new_net_7653)
	);

	bfr new_net_7654_bfr_after (
		.din(new_net_7653),
		.dout(new_net_7654)
	);

	bfr new_net_7655_bfr_after (
		.din(new_net_7654),
		.dout(new_net_7655)
	);

	bfr new_net_7656_bfr_after (
		.din(new_net_7655),
		.dout(new_net_7656)
	);

	bfr new_net_7657_bfr_after (
		.din(new_net_7656),
		.dout(new_net_7657)
	);

	bfr new_net_7658_bfr_after (
		.din(new_net_7657),
		.dout(new_net_7658)
	);

	bfr new_net_7659_bfr_after (
		.din(new_net_7658),
		.dout(new_net_7659)
	);

	bfr new_net_7660_bfr_after (
		.din(new_net_7659),
		.dout(new_net_7660)
	);

	bfr new_net_7661_bfr_after (
		.din(new_net_7660),
		.dout(new_net_7661)
	);

	bfr new_net_7662_bfr_after (
		.din(new_net_7661),
		.dout(new_net_7662)
	);

	bfr new_net_7663_bfr_after (
		.din(new_net_7662),
		.dout(new_net_7663)
	);

	bfr new_net_7664_bfr_after (
		.din(new_net_7663),
		.dout(new_net_7664)
	);

	bfr new_net_7665_bfr_after (
		.din(new_net_7664),
		.dout(new_net_7665)
	);

	bfr new_net_7666_bfr_after (
		.din(new_net_7665),
		.dout(new_net_7666)
	);

	bfr new_net_7667_bfr_after (
		.din(new_net_7666),
		.dout(new_net_7667)
	);

	bfr new_net_7668_bfr_after (
		.din(new_net_7667),
		.dout(new_net_7668)
	);

	bfr new_net_7669_bfr_after (
		.din(new_net_7668),
		.dout(new_net_7669)
	);

	bfr new_net_7670_bfr_after (
		.din(new_net_7669),
		.dout(new_net_7670)
	);

	bfr new_net_7671_bfr_after (
		.din(new_net_7670),
		.dout(new_net_7671)
	);

	bfr new_net_7672_bfr_after (
		.din(new_net_7671),
		.dout(new_net_7672)
	);

	bfr new_net_7673_bfr_after (
		.din(new_net_7672),
		.dout(new_net_7673)
	);

	bfr new_net_7674_bfr_after (
		.din(new_net_7673),
		.dout(new_net_7674)
	);

	bfr new_net_7675_bfr_after (
		.din(new_net_7674),
		.dout(new_net_7675)
	);

	bfr new_net_7676_bfr_after (
		.din(new_net_7675),
		.dout(new_net_7676)
	);

	bfr new_net_7677_bfr_after (
		.din(new_net_7676),
		.dout(new_net_7677)
	);

	bfr new_net_7678_bfr_after (
		.din(new_net_7677),
		.dout(new_net_7678)
	);

	bfr new_net_7679_bfr_after (
		.din(new_net_7678),
		.dout(new_net_7679)
	);

	bfr new_net_7680_bfr_after (
		.din(new_net_7679),
		.dout(new_net_7680)
	);

	bfr new_net_7681_bfr_after (
		.din(new_net_7680),
		.dout(new_net_7681)
	);

	bfr new_net_7682_bfr_after (
		.din(new_net_7681),
		.dout(new_net_7682)
	);

	bfr new_net_7683_bfr_after (
		.din(new_net_7682),
		.dout(new_net_7683)
	);

	bfr new_net_7684_bfr_after (
		.din(new_net_7683),
		.dout(new_net_7684)
	);

	bfr new_net_7685_bfr_after (
		.din(new_net_7684),
		.dout(new_net_7685)
	);

	bfr new_net_7686_bfr_after (
		.din(new_net_7685),
		.dout(new_net_7686)
	);

	bfr new_net_7687_bfr_after (
		.din(new_net_7686),
		.dout(new_net_7687)
	);

	bfr new_net_7688_bfr_after (
		.din(new_net_7687),
		.dout(new_net_7688)
	);

	bfr new_net_7689_bfr_after (
		.din(new_net_7688),
		.dout(new_net_7689)
	);

	bfr new_net_7690_bfr_after (
		.din(new_net_7689),
		.dout(new_net_7690)
	);

	bfr new_net_7691_bfr_after (
		.din(new_net_7690),
		.dout(new_net_7691)
	);

	bfr new_net_7692_bfr_after (
		.din(new_net_7691),
		.dout(new_net_7692)
	);

	bfr new_net_7693_bfr_after (
		.din(new_net_7692),
		.dout(new_net_7693)
	);

	bfr new_net_7694_bfr_after (
		.din(new_net_7693),
		.dout(new_net_7694)
	);

	bfr new_net_7695_bfr_after (
		.din(new_net_7694),
		.dout(new_net_7695)
	);

	bfr new_net_7696_bfr_after (
		.din(new_net_7695),
		.dout(new_net_7696)
	);

	bfr new_net_7697_bfr_after (
		.din(new_net_7696),
		.dout(new_net_7697)
	);

	bfr new_net_7698_bfr_after (
		.din(new_net_7697),
		.dout(new_net_7698)
	);

	bfr new_net_7699_bfr_after (
		.din(new_net_7698),
		.dout(new_net_7699)
	);

	bfr new_net_7700_bfr_after (
		.din(new_net_7699),
		.dout(new_net_7700)
	);

	bfr new_net_7701_bfr_after (
		.din(new_net_7700),
		.dout(new_net_7701)
	);

	bfr new_net_7702_bfr_after (
		.din(new_net_7701),
		.dout(new_net_7702)
	);

	bfr new_net_7703_bfr_after (
		.din(new_net_7702),
		.dout(new_net_7703)
	);

	bfr new_net_7704_bfr_after (
		.din(new_net_7703),
		.dout(new_net_7704)
	);

	bfr new_net_7705_bfr_after (
		.din(new_net_7704),
		.dout(new_net_7705)
	);

	bfr new_net_7706_bfr_after (
		.din(new_net_7705),
		.dout(new_net_7706)
	);

	bfr new_net_7707_bfr_after (
		.din(new_net_7706),
		.dout(new_net_7707)
	);

	bfr new_net_7708_bfr_after (
		.din(new_net_7707),
		.dout(new_net_7708)
	);

	bfr new_net_7709_bfr_after (
		.din(new_net_7708),
		.dout(new_net_7709)
	);

	bfr new_net_7710_bfr_after (
		.din(new_net_7709),
		.dout(new_net_7710)
	);

	bfr new_net_7711_bfr_after (
		.din(new_net_7710),
		.dout(new_net_7711)
	);

	bfr new_net_7712_bfr_after (
		.din(new_net_7711),
		.dout(new_net_7712)
	);

	bfr new_net_7713_bfr_after (
		.din(new_net_7712),
		.dout(new_net_7713)
	);

	bfr new_net_7714_bfr_after (
		.din(new_net_7713),
		.dout(new_net_7714)
	);

	bfr new_net_7715_bfr_after (
		.din(new_net_7714),
		.dout(new_net_7715)
	);

	bfr new_net_7716_bfr_after (
		.din(new_net_7715),
		.dout(new_net_7716)
	);

	bfr new_net_7717_bfr_after (
		.din(new_net_7716),
		.dout(new_net_7717)
	);

	bfr new_net_7718_bfr_after (
		.din(new_net_7717),
		.dout(new_net_7718)
	);

	bfr new_net_7719_bfr_after (
		.din(new_net_7718),
		.dout(new_net_7719)
	);

	bfr new_net_7720_bfr_after (
		.din(new_net_7719),
		.dout(new_net_7720)
	);

	bfr new_net_7721_bfr_after (
		.din(new_net_7720),
		.dout(new_net_7721)
	);

	bfr new_net_7722_bfr_after (
		.din(new_net_7721),
		.dout(new_net_7722)
	);

	bfr new_net_7723_bfr_after (
		.din(new_net_7722),
		.dout(new_net_7723)
	);

	bfr new_net_7724_bfr_after (
		.din(new_net_7723),
		.dout(new_net_7724)
	);

	spl2 _1813__v_fanout (
		.a(new_net_7724),
		.b(new_net_608),
		.c(new_net_609)
	);

	bfr new_net_7725_bfr_after (
		.din(_0106_),
		.dout(new_net_7725)
	);

	bfr new_net_7726_bfr_after (
		.din(new_net_7725),
		.dout(new_net_7726)
	);

	bfr new_net_7727_bfr_after (
		.din(new_net_7726),
		.dout(new_net_7727)
	);

	bfr new_net_7728_bfr_after (
		.din(new_net_7727),
		.dout(new_net_7728)
	);

	bfr new_net_7729_bfr_after (
		.din(new_net_7728),
		.dout(new_net_7729)
	);

	bfr new_net_7730_bfr_after (
		.din(new_net_7729),
		.dout(new_net_7730)
	);

	bfr new_net_7731_bfr_after (
		.din(new_net_7730),
		.dout(new_net_7731)
	);

	bfr new_net_7732_bfr_after (
		.din(new_net_7731),
		.dout(new_net_7732)
	);

	bfr new_net_7733_bfr_after (
		.din(new_net_7732),
		.dout(new_net_7733)
	);

	bfr new_net_7734_bfr_after (
		.din(new_net_7733),
		.dout(new_net_7734)
	);

	bfr new_net_7735_bfr_after (
		.din(new_net_7734),
		.dout(new_net_7735)
	);

	bfr new_net_7736_bfr_after (
		.din(new_net_7735),
		.dout(new_net_7736)
	);

	bfr new_net_7737_bfr_after (
		.din(new_net_7736),
		.dout(new_net_7737)
	);

	bfr new_net_7738_bfr_after (
		.din(new_net_7737),
		.dout(new_net_7738)
	);

	bfr new_net_7739_bfr_after (
		.din(new_net_7738),
		.dout(new_net_7739)
	);

	bfr new_net_7740_bfr_after (
		.din(new_net_7739),
		.dout(new_net_7740)
	);

	bfr new_net_7741_bfr_after (
		.din(new_net_7740),
		.dout(new_net_7741)
	);

	bfr new_net_7742_bfr_after (
		.din(new_net_7741),
		.dout(new_net_7742)
	);

	bfr new_net_7743_bfr_after (
		.din(new_net_7742),
		.dout(new_net_7743)
	);

	bfr new_net_7744_bfr_after (
		.din(new_net_7743),
		.dout(new_net_7744)
	);

	bfr new_net_7745_bfr_after (
		.din(new_net_7744),
		.dout(new_net_7745)
	);

	bfr new_net_7746_bfr_after (
		.din(new_net_7745),
		.dout(new_net_7746)
	);

	bfr new_net_7747_bfr_after (
		.din(new_net_7746),
		.dout(new_net_7747)
	);

	bfr new_net_7748_bfr_after (
		.din(new_net_7747),
		.dout(new_net_7748)
	);

	bfr new_net_7749_bfr_after (
		.din(new_net_7748),
		.dout(new_net_7749)
	);

	bfr new_net_7750_bfr_after (
		.din(new_net_7749),
		.dout(new_net_7750)
	);

	bfr new_net_7751_bfr_after (
		.din(new_net_7750),
		.dout(new_net_7751)
	);

	bfr new_net_7752_bfr_after (
		.din(new_net_7751),
		.dout(new_net_7752)
	);

	bfr new_net_7753_bfr_after (
		.din(new_net_7752),
		.dout(new_net_7753)
	);

	bfr new_net_7754_bfr_after (
		.din(new_net_7753),
		.dout(new_net_7754)
	);

	bfr new_net_7755_bfr_after (
		.din(new_net_7754),
		.dout(new_net_7755)
	);

	bfr new_net_7756_bfr_after (
		.din(new_net_7755),
		.dout(new_net_7756)
	);

	spl2 _0106__v_fanout (
		.a(new_net_7756),
		.b(new_net_1870),
		.c(new_net_1871)
	);

	bfr new_net_7757_bfr_after (
		.din(_1827_),
		.dout(new_net_7757)
	);

	bfr new_net_7758_bfr_after (
		.din(new_net_7757),
		.dout(new_net_7758)
	);

	bfr new_net_7759_bfr_after (
		.din(new_net_7758),
		.dout(new_net_7759)
	);

	bfr new_net_7760_bfr_after (
		.din(new_net_7759),
		.dout(new_net_7760)
	);

	bfr new_net_7761_bfr_after (
		.din(new_net_7760),
		.dout(new_net_7761)
	);

	bfr new_net_7762_bfr_after (
		.din(new_net_7761),
		.dout(new_net_7762)
	);

	bfr new_net_7763_bfr_after (
		.din(new_net_7762),
		.dout(new_net_7763)
	);

	bfr new_net_7764_bfr_after (
		.din(new_net_7763),
		.dout(new_net_7764)
	);

	bfr new_net_7765_bfr_after (
		.din(new_net_7764),
		.dout(new_net_7765)
	);

	bfr new_net_7766_bfr_after (
		.din(new_net_7765),
		.dout(new_net_7766)
	);

	bfr new_net_7767_bfr_after (
		.din(new_net_7766),
		.dout(new_net_7767)
	);

	bfr new_net_7768_bfr_after (
		.din(new_net_7767),
		.dout(new_net_7768)
	);

	bfr new_net_7769_bfr_after (
		.din(new_net_7768),
		.dout(new_net_7769)
	);

	bfr new_net_7770_bfr_after (
		.din(new_net_7769),
		.dout(new_net_7770)
	);

	bfr new_net_7771_bfr_after (
		.din(new_net_7770),
		.dout(new_net_7771)
	);

	bfr new_net_7772_bfr_after (
		.din(new_net_7771),
		.dout(new_net_7772)
	);

	bfr new_net_7773_bfr_after (
		.din(new_net_7772),
		.dout(new_net_7773)
	);

	bfr new_net_7774_bfr_after (
		.din(new_net_7773),
		.dout(new_net_7774)
	);

	bfr new_net_7775_bfr_after (
		.din(new_net_7774),
		.dout(new_net_7775)
	);

	bfr new_net_7776_bfr_after (
		.din(new_net_7775),
		.dout(new_net_7776)
	);

	bfr new_net_7777_bfr_after (
		.din(new_net_7776),
		.dout(new_net_7777)
	);

	bfr new_net_7778_bfr_after (
		.din(new_net_7777),
		.dout(new_net_7778)
	);

	bfr new_net_7779_bfr_after (
		.din(new_net_7778),
		.dout(new_net_7779)
	);

	bfr new_net_7780_bfr_after (
		.din(new_net_7779),
		.dout(new_net_7780)
	);

	bfr new_net_7781_bfr_after (
		.din(new_net_7780),
		.dout(new_net_7781)
	);

	bfr new_net_7782_bfr_after (
		.din(new_net_7781),
		.dout(new_net_7782)
	);

	bfr new_net_7783_bfr_after (
		.din(new_net_7782),
		.dout(new_net_7783)
	);

	bfr new_net_7784_bfr_after (
		.din(new_net_7783),
		.dout(new_net_7784)
	);

	bfr new_net_7785_bfr_after (
		.din(new_net_7784),
		.dout(new_net_7785)
	);

	bfr new_net_7786_bfr_after (
		.din(new_net_7785),
		.dout(new_net_7786)
	);

	bfr new_net_7787_bfr_after (
		.din(new_net_7786),
		.dout(new_net_7787)
	);

	bfr new_net_7788_bfr_after (
		.din(new_net_7787),
		.dout(new_net_7788)
	);

	bfr new_net_7789_bfr_after (
		.din(new_net_7788),
		.dout(new_net_7789)
	);

	bfr new_net_7790_bfr_after (
		.din(new_net_7789),
		.dout(new_net_7790)
	);

	bfr new_net_7791_bfr_after (
		.din(new_net_7790),
		.dout(new_net_7791)
	);

	bfr new_net_7792_bfr_after (
		.din(new_net_7791),
		.dout(new_net_7792)
	);

	bfr new_net_7793_bfr_after (
		.din(new_net_7792),
		.dout(new_net_7793)
	);

	bfr new_net_7794_bfr_after (
		.din(new_net_7793),
		.dout(new_net_7794)
	);

	bfr new_net_7795_bfr_after (
		.din(new_net_7794),
		.dout(new_net_7795)
	);

	bfr new_net_7796_bfr_after (
		.din(new_net_7795),
		.dout(new_net_7796)
	);

	bfr new_net_7797_bfr_after (
		.din(new_net_7796),
		.dout(new_net_7797)
	);

	bfr new_net_7798_bfr_after (
		.din(new_net_7797),
		.dout(new_net_7798)
	);

	bfr new_net_7799_bfr_after (
		.din(new_net_7798),
		.dout(new_net_7799)
	);

	bfr new_net_7800_bfr_after (
		.din(new_net_7799),
		.dout(new_net_7800)
	);

	bfr new_net_7801_bfr_after (
		.din(new_net_7800),
		.dout(new_net_7801)
	);

	bfr new_net_7802_bfr_after (
		.din(new_net_7801),
		.dout(new_net_7802)
	);

	bfr new_net_7803_bfr_after (
		.din(new_net_7802),
		.dout(new_net_7803)
	);

	bfr new_net_7804_bfr_after (
		.din(new_net_7803),
		.dout(new_net_7804)
	);

	bfr new_net_7805_bfr_after (
		.din(new_net_7804),
		.dout(new_net_7805)
	);

	bfr new_net_7806_bfr_after (
		.din(new_net_7805),
		.dout(new_net_7806)
	);

	bfr new_net_7807_bfr_after (
		.din(new_net_7806),
		.dout(new_net_7807)
	);

	bfr new_net_7808_bfr_after (
		.din(new_net_7807),
		.dout(new_net_7808)
	);

	bfr new_net_7809_bfr_after (
		.din(new_net_7808),
		.dout(new_net_7809)
	);

	bfr new_net_7810_bfr_after (
		.din(new_net_7809),
		.dout(new_net_7810)
	);

	bfr new_net_7811_bfr_after (
		.din(new_net_7810),
		.dout(new_net_7811)
	);

	bfr new_net_7812_bfr_after (
		.din(new_net_7811),
		.dout(new_net_7812)
	);

	bfr new_net_7813_bfr_after (
		.din(new_net_7812),
		.dout(new_net_7813)
	);

	bfr new_net_7814_bfr_after (
		.din(new_net_7813),
		.dout(new_net_7814)
	);

	bfr new_net_7815_bfr_after (
		.din(new_net_7814),
		.dout(new_net_7815)
	);

	bfr new_net_7816_bfr_after (
		.din(new_net_7815),
		.dout(new_net_7816)
	);

	bfr new_net_7817_bfr_after (
		.din(new_net_7816),
		.dout(new_net_7817)
	);

	bfr new_net_7818_bfr_after (
		.din(new_net_7817),
		.dout(new_net_7818)
	);

	bfr new_net_7819_bfr_after (
		.din(new_net_7818),
		.dout(new_net_7819)
	);

	bfr new_net_7820_bfr_after (
		.din(new_net_7819),
		.dout(new_net_7820)
	);

	spl2 _1827__v_fanout (
		.a(new_net_7820),
		.b(new_net_814),
		.c(new_net_815)
	);

	spl2 _1643__v_fanout (
		.a(_1643_),
		.b(new_net_2880),
		.c(new_net_2881)
	);

	bfr new_net_7821_bfr_after (
		.din(_0538_),
		.dout(new_net_7821)
	);

	bfr new_net_7822_bfr_after (
		.din(new_net_7821),
		.dout(new_net_7822)
	);

	bfr new_net_7823_bfr_after (
		.din(new_net_7822),
		.dout(new_net_7823)
	);

	bfr new_net_7824_bfr_after (
		.din(new_net_7823),
		.dout(new_net_7824)
	);

	bfr new_net_7825_bfr_after (
		.din(new_net_7824),
		.dout(new_net_7825)
	);

	bfr new_net_7826_bfr_after (
		.din(new_net_7825),
		.dout(new_net_7826)
	);

	bfr new_net_7827_bfr_after (
		.din(new_net_7826),
		.dout(new_net_7827)
	);

	bfr new_net_7828_bfr_after (
		.din(new_net_7827),
		.dout(new_net_7828)
	);

	bfr new_net_7829_bfr_after (
		.din(new_net_7828),
		.dout(new_net_7829)
	);

	bfr new_net_7830_bfr_after (
		.din(new_net_7829),
		.dout(new_net_7830)
	);

	bfr new_net_7831_bfr_after (
		.din(new_net_7830),
		.dout(new_net_7831)
	);

	bfr new_net_7832_bfr_after (
		.din(new_net_7831),
		.dout(new_net_7832)
	);

	bfr new_net_7833_bfr_after (
		.din(new_net_7832),
		.dout(new_net_7833)
	);

	bfr new_net_7834_bfr_after (
		.din(new_net_7833),
		.dout(new_net_7834)
	);

	bfr new_net_7835_bfr_after (
		.din(new_net_7834),
		.dout(new_net_7835)
	);

	bfr new_net_7836_bfr_after (
		.din(new_net_7835),
		.dout(new_net_7836)
	);

	bfr new_net_7837_bfr_after (
		.din(new_net_7836),
		.dout(new_net_7837)
	);

	bfr new_net_7838_bfr_after (
		.din(new_net_7837),
		.dout(new_net_7838)
	);

	bfr new_net_7839_bfr_after (
		.din(new_net_7838),
		.dout(new_net_7839)
	);

	bfr new_net_7840_bfr_after (
		.din(new_net_7839),
		.dout(new_net_7840)
	);

	bfr new_net_7841_bfr_after (
		.din(new_net_7840),
		.dout(new_net_7841)
	);

	bfr new_net_7842_bfr_after (
		.din(new_net_7841),
		.dout(new_net_7842)
	);

	bfr new_net_7843_bfr_after (
		.din(new_net_7842),
		.dout(new_net_7843)
	);

	bfr new_net_7844_bfr_after (
		.din(new_net_7843),
		.dout(new_net_7844)
	);

	bfr new_net_7845_bfr_after (
		.din(new_net_7844),
		.dout(new_net_7845)
	);

	bfr new_net_7846_bfr_after (
		.din(new_net_7845),
		.dout(new_net_7846)
	);

	bfr new_net_7847_bfr_after (
		.din(new_net_7846),
		.dout(new_net_7847)
	);

	bfr new_net_7848_bfr_after (
		.din(new_net_7847),
		.dout(new_net_7848)
	);

	bfr new_net_7849_bfr_after (
		.din(new_net_7848),
		.dout(new_net_7849)
	);

	bfr new_net_7850_bfr_after (
		.din(new_net_7849),
		.dout(new_net_7850)
	);

	bfr new_net_7851_bfr_after (
		.din(new_net_7850),
		.dout(new_net_7851)
	);

	bfr new_net_7852_bfr_after (
		.din(new_net_7851),
		.dout(new_net_7852)
	);

	bfr new_net_7853_bfr_after (
		.din(new_net_7852),
		.dout(new_net_7853)
	);

	bfr new_net_7854_bfr_after (
		.din(new_net_7853),
		.dout(new_net_7854)
	);

	bfr new_net_7855_bfr_after (
		.din(new_net_7854),
		.dout(new_net_7855)
	);

	bfr new_net_7856_bfr_after (
		.din(new_net_7855),
		.dout(new_net_7856)
	);

	bfr new_net_7857_bfr_after (
		.din(new_net_7856),
		.dout(new_net_7857)
	);

	bfr new_net_7858_bfr_after (
		.din(new_net_7857),
		.dout(new_net_7858)
	);

	bfr new_net_7859_bfr_after (
		.din(new_net_7858),
		.dout(new_net_7859)
	);

	bfr new_net_7860_bfr_after (
		.din(new_net_7859),
		.dout(new_net_7860)
	);

	bfr new_net_7861_bfr_after (
		.din(new_net_7860),
		.dout(new_net_7861)
	);

	bfr new_net_7862_bfr_after (
		.din(new_net_7861),
		.dout(new_net_7862)
	);

	bfr new_net_7863_bfr_after (
		.din(new_net_7862),
		.dout(new_net_7863)
	);

	bfr new_net_7864_bfr_after (
		.din(new_net_7863),
		.dout(new_net_7864)
	);

	bfr new_net_7865_bfr_after (
		.din(new_net_7864),
		.dout(new_net_7865)
	);

	bfr new_net_7866_bfr_after (
		.din(new_net_7865),
		.dout(new_net_7866)
	);

	bfr new_net_7867_bfr_after (
		.din(new_net_7866),
		.dout(new_net_7867)
	);

	bfr new_net_7868_bfr_after (
		.din(new_net_7867),
		.dout(new_net_7868)
	);

	bfr new_net_7869_bfr_after (
		.din(new_net_7868),
		.dout(new_net_7869)
	);

	bfr new_net_7870_bfr_after (
		.din(new_net_7869),
		.dout(new_net_7870)
	);

	bfr new_net_7871_bfr_after (
		.din(new_net_7870),
		.dout(new_net_7871)
	);

	bfr new_net_7872_bfr_after (
		.din(new_net_7871),
		.dout(new_net_7872)
	);

	bfr new_net_7873_bfr_after (
		.din(new_net_7872),
		.dout(new_net_7873)
	);

	bfr new_net_7874_bfr_after (
		.din(new_net_7873),
		.dout(new_net_7874)
	);

	bfr new_net_7875_bfr_after (
		.din(new_net_7874),
		.dout(new_net_7875)
	);

	bfr new_net_7876_bfr_after (
		.din(new_net_7875),
		.dout(new_net_7876)
	);

	bfr new_net_7877_bfr_after (
		.din(new_net_7876),
		.dout(new_net_7877)
	);

	bfr new_net_7878_bfr_after (
		.din(new_net_7877),
		.dout(new_net_7878)
	);

	bfr new_net_7879_bfr_after (
		.din(new_net_7878),
		.dout(new_net_7879)
	);

	bfr new_net_7880_bfr_after (
		.din(new_net_7879),
		.dout(new_net_7880)
	);

	bfr new_net_7881_bfr_after (
		.din(new_net_7880),
		.dout(new_net_7881)
	);

	bfr new_net_7882_bfr_after (
		.din(new_net_7881),
		.dout(new_net_7882)
	);

	bfr new_net_7883_bfr_after (
		.din(new_net_7882),
		.dout(new_net_7883)
	);

	bfr new_net_7884_bfr_after (
		.din(new_net_7883),
		.dout(new_net_7884)
	);

	bfr new_net_7885_bfr_after (
		.din(new_net_7884),
		.dout(new_net_7885)
	);

	bfr new_net_7886_bfr_after (
		.din(new_net_7885),
		.dout(new_net_7886)
	);

	bfr new_net_7887_bfr_after (
		.din(new_net_7886),
		.dout(new_net_7887)
	);

	bfr new_net_7888_bfr_after (
		.din(new_net_7887),
		.dout(new_net_7888)
	);

	bfr new_net_7889_bfr_after (
		.din(new_net_7888),
		.dout(new_net_7889)
	);

	bfr new_net_7890_bfr_after (
		.din(new_net_7889),
		.dout(new_net_7890)
	);

	bfr new_net_7891_bfr_after (
		.din(new_net_7890),
		.dout(new_net_7891)
	);

	bfr new_net_7892_bfr_after (
		.din(new_net_7891),
		.dout(new_net_7892)
	);

	bfr new_net_7893_bfr_after (
		.din(new_net_7892),
		.dout(new_net_7893)
	);

	bfr new_net_7894_bfr_after (
		.din(new_net_7893),
		.dout(new_net_7894)
	);

	bfr new_net_7895_bfr_after (
		.din(new_net_7894),
		.dout(new_net_7895)
	);

	bfr new_net_7896_bfr_after (
		.din(new_net_7895),
		.dout(new_net_7896)
	);

	bfr new_net_7897_bfr_after (
		.din(new_net_7896),
		.dout(new_net_7897)
	);

	bfr new_net_7898_bfr_after (
		.din(new_net_7897),
		.dout(new_net_7898)
	);

	bfr new_net_7899_bfr_after (
		.din(new_net_7898),
		.dout(new_net_7899)
	);

	bfr new_net_7900_bfr_after (
		.din(new_net_7899),
		.dout(new_net_7900)
	);

	spl2 _0538__v_fanout (
		.a(new_net_7900),
		.b(new_net_2359),
		.c(new_net_2360)
	);

	bfr new_net_7901_bfr_after (
		.din(_0634_),
		.dout(new_net_7901)
	);

	bfr new_net_7902_bfr_after (
		.din(new_net_7901),
		.dout(new_net_7902)
	);

	bfr new_net_7903_bfr_after (
		.din(new_net_7902),
		.dout(new_net_7903)
	);

	bfr new_net_7904_bfr_after (
		.din(new_net_7903),
		.dout(new_net_7904)
	);

	bfr new_net_7905_bfr_after (
		.din(new_net_7904),
		.dout(new_net_7905)
	);

	bfr new_net_7906_bfr_after (
		.din(new_net_7905),
		.dout(new_net_7906)
	);

	bfr new_net_7907_bfr_after (
		.din(new_net_7906),
		.dout(new_net_7907)
	);

	bfr new_net_7908_bfr_after (
		.din(new_net_7907),
		.dout(new_net_7908)
	);

	bfr new_net_7909_bfr_after (
		.din(new_net_7908),
		.dout(new_net_7909)
	);

	bfr new_net_7910_bfr_after (
		.din(new_net_7909),
		.dout(new_net_7910)
	);

	bfr new_net_7911_bfr_after (
		.din(new_net_7910),
		.dout(new_net_7911)
	);

	bfr new_net_7912_bfr_after (
		.din(new_net_7911),
		.dout(new_net_7912)
	);

	bfr new_net_7913_bfr_after (
		.din(new_net_7912),
		.dout(new_net_7913)
	);

	bfr new_net_7914_bfr_after (
		.din(new_net_7913),
		.dout(new_net_7914)
	);

	bfr new_net_7915_bfr_after (
		.din(new_net_7914),
		.dout(new_net_7915)
	);

	bfr new_net_7916_bfr_after (
		.din(new_net_7915),
		.dout(new_net_7916)
	);

	bfr new_net_7917_bfr_after (
		.din(new_net_7916),
		.dout(new_net_7917)
	);

	bfr new_net_7918_bfr_after (
		.din(new_net_7917),
		.dout(new_net_7918)
	);

	bfr new_net_7919_bfr_after (
		.din(new_net_7918),
		.dout(new_net_7919)
	);

	bfr new_net_7920_bfr_after (
		.din(new_net_7919),
		.dout(new_net_7920)
	);

	bfr new_net_7921_bfr_after (
		.din(new_net_7920),
		.dout(new_net_7921)
	);

	bfr new_net_7922_bfr_after (
		.din(new_net_7921),
		.dout(new_net_7922)
	);

	bfr new_net_7923_bfr_after (
		.din(new_net_7922),
		.dout(new_net_7923)
	);

	bfr new_net_7924_bfr_after (
		.din(new_net_7923),
		.dout(new_net_7924)
	);

	bfr new_net_7925_bfr_after (
		.din(new_net_7924),
		.dout(new_net_7925)
	);

	bfr new_net_7926_bfr_after (
		.din(new_net_7925),
		.dout(new_net_7926)
	);

	bfr new_net_7927_bfr_after (
		.din(new_net_7926),
		.dout(new_net_7927)
	);

	bfr new_net_7928_bfr_after (
		.din(new_net_7927),
		.dout(new_net_7928)
	);

	bfr new_net_7929_bfr_after (
		.din(new_net_7928),
		.dout(new_net_7929)
	);

	bfr new_net_7930_bfr_after (
		.din(new_net_7929),
		.dout(new_net_7930)
	);

	bfr new_net_7931_bfr_after (
		.din(new_net_7930),
		.dout(new_net_7931)
	);

	bfr new_net_7932_bfr_after (
		.din(new_net_7931),
		.dout(new_net_7932)
	);

	bfr new_net_7933_bfr_after (
		.din(new_net_7932),
		.dout(new_net_7933)
	);

	bfr new_net_7934_bfr_after (
		.din(new_net_7933),
		.dout(new_net_7934)
	);

	bfr new_net_7935_bfr_after (
		.din(new_net_7934),
		.dout(new_net_7935)
	);

	bfr new_net_7936_bfr_after (
		.din(new_net_7935),
		.dout(new_net_7936)
	);

	bfr new_net_7937_bfr_after (
		.din(new_net_7936),
		.dout(new_net_7937)
	);

	bfr new_net_7938_bfr_after (
		.din(new_net_7937),
		.dout(new_net_7938)
	);

	bfr new_net_7939_bfr_after (
		.din(new_net_7938),
		.dout(new_net_7939)
	);

	bfr new_net_7940_bfr_after (
		.din(new_net_7939),
		.dout(new_net_7940)
	);

	bfr new_net_7941_bfr_after (
		.din(new_net_7940),
		.dout(new_net_7941)
	);

	bfr new_net_7942_bfr_after (
		.din(new_net_7941),
		.dout(new_net_7942)
	);

	bfr new_net_7943_bfr_after (
		.din(new_net_7942),
		.dout(new_net_7943)
	);

	bfr new_net_7944_bfr_after (
		.din(new_net_7943),
		.dout(new_net_7944)
	);

	bfr new_net_7945_bfr_after (
		.din(new_net_7944),
		.dout(new_net_7945)
	);

	bfr new_net_7946_bfr_after (
		.din(new_net_7945),
		.dout(new_net_7946)
	);

	spl2 _0634__v_fanout (
		.a(new_net_7946),
		.b(new_net_2311),
		.c(new_net_2312)
	);

	bfr new_net_7947_bfr_after (
		.din(_1832_),
		.dout(new_net_7947)
	);

	bfr new_net_7948_bfr_after (
		.din(new_net_7947),
		.dout(new_net_7948)
	);

	spl2 _1832__v_fanout (
		.a(new_net_7948),
		.b(new_net_2020),
		.c(new_net_2021)
	);

	bfr new_net_7949_bfr_after (
		.din(_1130_),
		.dout(new_net_7949)
	);

	bfr new_net_7950_bfr_after (
		.din(new_net_7949),
		.dout(new_net_7950)
	);

	bfr new_net_7951_bfr_after (
		.din(new_net_7950),
		.dout(new_net_7951)
	);

	bfr new_net_7952_bfr_after (
		.din(new_net_7951),
		.dout(new_net_7952)
	);

	bfr new_net_7953_bfr_after (
		.din(new_net_7952),
		.dout(new_net_7953)
	);

	bfr new_net_7954_bfr_after (
		.din(new_net_7953),
		.dout(new_net_7954)
	);

	bfr new_net_7955_bfr_after (
		.din(new_net_7954),
		.dout(new_net_7955)
	);

	bfr new_net_7956_bfr_after (
		.din(new_net_7955),
		.dout(new_net_7956)
	);

	bfr new_net_7957_bfr_after (
		.din(new_net_7956),
		.dout(new_net_7957)
	);

	bfr new_net_7958_bfr_after (
		.din(new_net_7957),
		.dout(new_net_7958)
	);

	bfr new_net_7959_bfr_after (
		.din(new_net_7958),
		.dout(new_net_7959)
	);

	bfr new_net_7960_bfr_after (
		.din(new_net_7959),
		.dout(new_net_7960)
	);

	bfr new_net_7961_bfr_after (
		.din(new_net_7960),
		.dout(new_net_7961)
	);

	bfr new_net_7962_bfr_after (
		.din(new_net_7961),
		.dout(new_net_7962)
	);

	bfr new_net_7963_bfr_after (
		.din(new_net_7962),
		.dout(new_net_7963)
	);

	bfr new_net_7964_bfr_after (
		.din(new_net_7963),
		.dout(new_net_7964)
	);

	bfr new_net_7965_bfr_after (
		.din(new_net_7964),
		.dout(new_net_7965)
	);

	bfr new_net_7966_bfr_after (
		.din(new_net_7965),
		.dout(new_net_7966)
	);

	bfr new_net_7967_bfr_after (
		.din(new_net_7966),
		.dout(new_net_7967)
	);

	bfr new_net_7968_bfr_after (
		.din(new_net_7967),
		.dout(new_net_7968)
	);

	bfr new_net_7969_bfr_after (
		.din(new_net_7968),
		.dout(new_net_7969)
	);

	bfr new_net_7970_bfr_after (
		.din(new_net_7969),
		.dout(new_net_7970)
	);

	bfr new_net_7971_bfr_after (
		.din(new_net_7970),
		.dout(new_net_7971)
	);

	bfr new_net_7972_bfr_after (
		.din(new_net_7971),
		.dout(new_net_7972)
	);

	bfr new_net_7973_bfr_after (
		.din(new_net_7972),
		.dout(new_net_7973)
	);

	bfr new_net_7974_bfr_after (
		.din(new_net_7973),
		.dout(new_net_7974)
	);

	bfr new_net_7975_bfr_after (
		.din(new_net_7974),
		.dout(new_net_7975)
	);

	bfr new_net_7976_bfr_after (
		.din(new_net_7975),
		.dout(new_net_7976)
	);

	bfr new_net_7977_bfr_after (
		.din(new_net_7976),
		.dout(new_net_7977)
	);

	bfr new_net_7978_bfr_after (
		.din(new_net_7977),
		.dout(new_net_7978)
	);

	bfr new_net_7979_bfr_after (
		.din(new_net_7978),
		.dout(new_net_7979)
	);

	bfr new_net_7980_bfr_after (
		.din(new_net_7979),
		.dout(new_net_7980)
	);

	bfr new_net_7981_bfr_after (
		.din(new_net_7980),
		.dout(new_net_7981)
	);

	bfr new_net_7982_bfr_after (
		.din(new_net_7981),
		.dout(new_net_7982)
	);

	bfr new_net_7983_bfr_after (
		.din(new_net_7982),
		.dout(new_net_7983)
	);

	bfr new_net_7984_bfr_after (
		.din(new_net_7983),
		.dout(new_net_7984)
	);

	bfr new_net_7985_bfr_after (
		.din(new_net_7984),
		.dout(new_net_7985)
	);

	bfr new_net_7986_bfr_after (
		.din(new_net_7985),
		.dout(new_net_7986)
	);

	bfr new_net_7987_bfr_after (
		.din(new_net_7986),
		.dout(new_net_7987)
	);

	bfr new_net_7988_bfr_after (
		.din(new_net_7987),
		.dout(new_net_7988)
	);

	bfr new_net_7989_bfr_after (
		.din(new_net_7988),
		.dout(new_net_7989)
	);

	bfr new_net_7990_bfr_after (
		.din(new_net_7989),
		.dout(new_net_7990)
	);

	bfr new_net_7991_bfr_after (
		.din(new_net_7990),
		.dout(new_net_7991)
	);

	bfr new_net_7992_bfr_after (
		.din(new_net_7991),
		.dout(new_net_7992)
	);

	bfr new_net_7993_bfr_after (
		.din(new_net_7992),
		.dout(new_net_7993)
	);

	bfr new_net_7994_bfr_after (
		.din(new_net_7993),
		.dout(new_net_7994)
	);

	bfr new_net_7995_bfr_after (
		.din(new_net_7994),
		.dout(new_net_7995)
	);

	bfr new_net_7996_bfr_after (
		.din(new_net_7995),
		.dout(new_net_7996)
	);

	bfr new_net_7997_bfr_after (
		.din(new_net_7996),
		.dout(new_net_7997)
	);

	bfr new_net_7998_bfr_after (
		.din(new_net_7997),
		.dout(new_net_7998)
	);

	bfr new_net_7999_bfr_after (
		.din(new_net_7998),
		.dout(new_net_7999)
	);

	bfr new_net_8000_bfr_after (
		.din(new_net_7999),
		.dout(new_net_8000)
	);

	bfr new_net_8001_bfr_after (
		.din(new_net_8000),
		.dout(new_net_8001)
	);

	bfr new_net_8002_bfr_after (
		.din(new_net_8001),
		.dout(new_net_8002)
	);

	bfr new_net_8003_bfr_after (
		.din(new_net_8002),
		.dout(new_net_8003)
	);

	bfr new_net_8004_bfr_after (
		.din(new_net_8003),
		.dout(new_net_8004)
	);

	spl2 _1130__v_fanout (
		.a(new_net_8004),
		.b(new_net_938),
		.c(new_net_939)
	);

	bfr new_net_8005_bfr_after (
		.din(_1691_),
		.dout(new_net_8005)
	);

	bfr new_net_8006_bfr_after (
		.din(new_net_8005),
		.dout(new_net_8006)
	);

	bfr new_net_8007_bfr_after (
		.din(new_net_8006),
		.dout(new_net_8007)
	);

	bfr new_net_8008_bfr_after (
		.din(new_net_8007),
		.dout(new_net_8008)
	);

	bfr new_net_8009_bfr_after (
		.din(new_net_8008),
		.dout(new_net_8009)
	);

	bfr new_net_8010_bfr_after (
		.din(new_net_8009),
		.dout(new_net_8010)
	);

	bfr new_net_8011_bfr_after (
		.din(new_net_8010),
		.dout(new_net_8011)
	);

	bfr new_net_8012_bfr_after (
		.din(new_net_8011),
		.dout(new_net_8012)
	);

	bfr new_net_8013_bfr_after (
		.din(new_net_8012),
		.dout(new_net_8013)
	);

	bfr new_net_8014_bfr_after (
		.din(new_net_8013),
		.dout(new_net_8014)
	);

	bfr new_net_8015_bfr_after (
		.din(new_net_8014),
		.dout(new_net_8015)
	);

	bfr new_net_8016_bfr_after (
		.din(new_net_8015),
		.dout(new_net_8016)
	);

	bfr new_net_8017_bfr_after (
		.din(new_net_8016),
		.dout(new_net_8017)
	);

	bfr new_net_8018_bfr_after (
		.din(new_net_8017),
		.dout(new_net_8018)
	);

	bfr new_net_8019_bfr_after (
		.din(new_net_8018),
		.dout(new_net_8019)
	);

	bfr new_net_8020_bfr_after (
		.din(new_net_8019),
		.dout(new_net_8020)
	);

	bfr new_net_8021_bfr_after (
		.din(new_net_8020),
		.dout(new_net_8021)
	);

	bfr new_net_8022_bfr_after (
		.din(new_net_8021),
		.dout(new_net_8022)
	);

	bfr new_net_8023_bfr_after (
		.din(new_net_8022),
		.dout(new_net_8023)
	);

	bfr new_net_8024_bfr_after (
		.din(new_net_8023),
		.dout(new_net_8024)
	);

	bfr new_net_8025_bfr_after (
		.din(new_net_8024),
		.dout(new_net_8025)
	);

	bfr new_net_8026_bfr_after (
		.din(new_net_8025),
		.dout(new_net_8026)
	);

	bfr new_net_8027_bfr_after (
		.din(new_net_8026),
		.dout(new_net_8027)
	);

	bfr new_net_8028_bfr_after (
		.din(new_net_8027),
		.dout(new_net_8028)
	);

	bfr new_net_8029_bfr_after (
		.din(new_net_8028),
		.dout(new_net_8029)
	);

	bfr new_net_8030_bfr_after (
		.din(new_net_8029),
		.dout(new_net_8030)
	);

	bfr new_net_8031_bfr_after (
		.din(new_net_8030),
		.dout(new_net_8031)
	);

	bfr new_net_8032_bfr_after (
		.din(new_net_8031),
		.dout(new_net_8032)
	);

	bfr new_net_8033_bfr_after (
		.din(new_net_8032),
		.dout(new_net_8033)
	);

	bfr new_net_8034_bfr_after (
		.din(new_net_8033),
		.dout(new_net_8034)
	);

	bfr new_net_8035_bfr_after (
		.din(new_net_8034),
		.dout(new_net_8035)
	);

	bfr new_net_8036_bfr_after (
		.din(new_net_8035),
		.dout(new_net_8036)
	);

	bfr new_net_8037_bfr_after (
		.din(new_net_8036),
		.dout(new_net_8037)
	);

	bfr new_net_8038_bfr_after (
		.din(new_net_8037),
		.dout(new_net_8038)
	);

	bfr new_net_8039_bfr_after (
		.din(new_net_8038),
		.dout(new_net_8039)
	);

	bfr new_net_8040_bfr_after (
		.din(new_net_8039),
		.dout(new_net_8040)
	);

	bfr new_net_8041_bfr_after (
		.din(new_net_8040),
		.dout(new_net_8041)
	);

	bfr new_net_8042_bfr_after (
		.din(new_net_8041),
		.dout(new_net_8042)
	);

	bfr new_net_8043_bfr_after (
		.din(new_net_8042),
		.dout(new_net_8043)
	);

	bfr new_net_8044_bfr_after (
		.din(new_net_8043),
		.dout(new_net_8044)
	);

	bfr new_net_8045_bfr_after (
		.din(new_net_8044),
		.dout(new_net_8045)
	);

	bfr new_net_8046_bfr_after (
		.din(new_net_8045),
		.dout(new_net_8046)
	);

	bfr new_net_8047_bfr_after (
		.din(new_net_8046),
		.dout(new_net_8047)
	);

	bfr new_net_8048_bfr_after (
		.din(new_net_8047),
		.dout(new_net_8048)
	);

	bfr new_net_8049_bfr_after (
		.din(new_net_8048),
		.dout(new_net_8049)
	);

	bfr new_net_8050_bfr_after (
		.din(new_net_8049),
		.dout(new_net_8050)
	);

	bfr new_net_8051_bfr_after (
		.din(new_net_8050),
		.dout(new_net_8051)
	);

	bfr new_net_8052_bfr_after (
		.din(new_net_8051),
		.dout(new_net_8052)
	);

	bfr new_net_8053_bfr_after (
		.din(new_net_8052),
		.dout(new_net_8053)
	);

	bfr new_net_8054_bfr_after (
		.din(new_net_8053),
		.dout(new_net_8054)
	);

	bfr new_net_8055_bfr_after (
		.din(new_net_8054),
		.dout(new_net_8055)
	);

	bfr new_net_8056_bfr_after (
		.din(new_net_8055),
		.dout(new_net_8056)
	);

	bfr new_net_8057_bfr_after (
		.din(new_net_8056),
		.dout(new_net_8057)
	);

	bfr new_net_8058_bfr_after (
		.din(new_net_8057),
		.dout(new_net_8058)
	);

	bfr new_net_8059_bfr_after (
		.din(new_net_8058),
		.dout(new_net_8059)
	);

	bfr new_net_8060_bfr_after (
		.din(new_net_8059),
		.dout(new_net_8060)
	);

	bfr new_net_8061_bfr_after (
		.din(new_net_8060),
		.dout(new_net_8061)
	);

	bfr new_net_8062_bfr_after (
		.din(new_net_8061),
		.dout(new_net_8062)
	);

	bfr new_net_8063_bfr_after (
		.din(new_net_8062),
		.dout(new_net_8063)
	);

	bfr new_net_8064_bfr_after (
		.din(new_net_8063),
		.dout(new_net_8064)
	);

	bfr new_net_8065_bfr_after (
		.din(new_net_8064),
		.dout(new_net_8065)
	);

	bfr new_net_8066_bfr_after (
		.din(new_net_8065),
		.dout(new_net_8066)
	);

	bfr new_net_8067_bfr_after (
		.din(new_net_8066),
		.dout(new_net_8067)
	);

	bfr new_net_8068_bfr_after (
		.din(new_net_8067),
		.dout(new_net_8068)
	);

	spl2 _1691__v_fanout (
		.a(new_net_8068),
		.b(new_net_1465),
		.c(new_net_1466)
	);

	bfr new_net_8069_bfr_after (
		.din(_0627_),
		.dout(new_net_8069)
	);

	bfr new_net_8070_bfr_after (
		.din(new_net_8069),
		.dout(new_net_8070)
	);

	bfr new_net_8071_bfr_after (
		.din(new_net_8070),
		.dout(new_net_8071)
	);

	bfr new_net_8072_bfr_after (
		.din(new_net_8071),
		.dout(new_net_8072)
	);

	bfr new_net_8073_bfr_after (
		.din(new_net_8072),
		.dout(new_net_8073)
	);

	bfr new_net_8074_bfr_after (
		.din(new_net_8073),
		.dout(new_net_8074)
	);

	bfr new_net_8075_bfr_after (
		.din(new_net_8074),
		.dout(new_net_8075)
	);

	bfr new_net_8076_bfr_after (
		.din(new_net_8075),
		.dout(new_net_8076)
	);

	bfr new_net_8077_bfr_after (
		.din(new_net_8076),
		.dout(new_net_8077)
	);

	bfr new_net_8078_bfr_after (
		.din(new_net_8077),
		.dout(new_net_8078)
	);

	bfr new_net_8079_bfr_after (
		.din(new_net_8078),
		.dout(new_net_8079)
	);

	bfr new_net_8080_bfr_after (
		.din(new_net_8079),
		.dout(new_net_8080)
	);

	bfr new_net_8081_bfr_after (
		.din(new_net_8080),
		.dout(new_net_8081)
	);

	bfr new_net_8082_bfr_after (
		.din(new_net_8081),
		.dout(new_net_8082)
	);

	bfr new_net_8083_bfr_after (
		.din(new_net_8082),
		.dout(new_net_8083)
	);

	bfr new_net_8084_bfr_after (
		.din(new_net_8083),
		.dout(new_net_8084)
	);

	bfr new_net_8085_bfr_after (
		.din(new_net_8084),
		.dout(new_net_8085)
	);

	bfr new_net_8086_bfr_after (
		.din(new_net_8085),
		.dout(new_net_8086)
	);

	bfr new_net_8087_bfr_after (
		.din(new_net_8086),
		.dout(new_net_8087)
	);

	bfr new_net_8088_bfr_after (
		.din(new_net_8087),
		.dout(new_net_8088)
	);

	bfr new_net_8089_bfr_after (
		.din(new_net_8088),
		.dout(new_net_8089)
	);

	bfr new_net_8090_bfr_after (
		.din(new_net_8089),
		.dout(new_net_8090)
	);

	bfr new_net_8091_bfr_after (
		.din(new_net_8090),
		.dout(new_net_8091)
	);

	bfr new_net_8092_bfr_after (
		.din(new_net_8091),
		.dout(new_net_8092)
	);

	bfr new_net_8093_bfr_after (
		.din(new_net_8092),
		.dout(new_net_8093)
	);

	bfr new_net_8094_bfr_after (
		.din(new_net_8093),
		.dout(new_net_8094)
	);

	bfr new_net_8095_bfr_after (
		.din(new_net_8094),
		.dout(new_net_8095)
	);

	bfr new_net_8096_bfr_after (
		.din(new_net_8095),
		.dout(new_net_8096)
	);

	bfr new_net_8097_bfr_after (
		.din(new_net_8096),
		.dout(new_net_8097)
	);

	bfr new_net_8098_bfr_after (
		.din(new_net_8097),
		.dout(new_net_8098)
	);

	bfr new_net_8099_bfr_after (
		.din(new_net_8098),
		.dout(new_net_8099)
	);

	bfr new_net_8100_bfr_after (
		.din(new_net_8099),
		.dout(new_net_8100)
	);

	bfr new_net_8101_bfr_after (
		.din(new_net_8100),
		.dout(new_net_8101)
	);

	bfr new_net_8102_bfr_after (
		.din(new_net_8101),
		.dout(new_net_8102)
	);

	bfr new_net_8103_bfr_after (
		.din(new_net_8102),
		.dout(new_net_8103)
	);

	bfr new_net_8104_bfr_after (
		.din(new_net_8103),
		.dout(new_net_8104)
	);

	bfr new_net_8105_bfr_after (
		.din(new_net_8104),
		.dout(new_net_8105)
	);

	bfr new_net_8106_bfr_after (
		.din(new_net_8105),
		.dout(new_net_8106)
	);

	bfr new_net_8107_bfr_after (
		.din(new_net_8106),
		.dout(new_net_8107)
	);

	bfr new_net_8108_bfr_after (
		.din(new_net_8107),
		.dout(new_net_8108)
	);

	bfr new_net_8109_bfr_after (
		.din(new_net_8108),
		.dout(new_net_8109)
	);

	bfr new_net_8110_bfr_after (
		.din(new_net_8109),
		.dout(new_net_8110)
	);

	bfr new_net_8111_bfr_after (
		.din(new_net_8110),
		.dout(new_net_8111)
	);

	bfr new_net_8112_bfr_after (
		.din(new_net_8111),
		.dout(new_net_8112)
	);

	bfr new_net_8113_bfr_after (
		.din(new_net_8112),
		.dout(new_net_8113)
	);

	bfr new_net_8114_bfr_after (
		.din(new_net_8113),
		.dout(new_net_8114)
	);

	bfr new_net_8115_bfr_after (
		.din(new_net_8114),
		.dout(new_net_8115)
	);

	bfr new_net_8116_bfr_after (
		.din(new_net_8115),
		.dout(new_net_8116)
	);

	bfr new_net_8117_bfr_after (
		.din(new_net_8116),
		.dout(new_net_8117)
	);

	bfr new_net_8118_bfr_after (
		.din(new_net_8117),
		.dout(new_net_8118)
	);

	bfr new_net_8119_bfr_after (
		.din(new_net_8118),
		.dout(new_net_8119)
	);

	bfr new_net_8120_bfr_after (
		.din(new_net_8119),
		.dout(new_net_8120)
	);

	bfr new_net_8121_bfr_after (
		.din(new_net_8120),
		.dout(new_net_8121)
	);

	bfr new_net_8122_bfr_after (
		.din(new_net_8121),
		.dout(new_net_8122)
	);

	bfr new_net_8123_bfr_after (
		.din(new_net_8122),
		.dout(new_net_8123)
	);

	bfr new_net_8124_bfr_after (
		.din(new_net_8123),
		.dout(new_net_8124)
	);

	bfr new_net_8125_bfr_after (
		.din(new_net_8124),
		.dout(new_net_8125)
	);

	bfr new_net_8126_bfr_after (
		.din(new_net_8125),
		.dout(new_net_8126)
	);

	bfr new_net_8127_bfr_after (
		.din(new_net_8126),
		.dout(new_net_8127)
	);

	bfr new_net_8128_bfr_after (
		.din(new_net_8127),
		.dout(new_net_8128)
	);

	bfr new_net_8129_bfr_after (
		.din(new_net_8128),
		.dout(new_net_8129)
	);

	bfr new_net_8130_bfr_after (
		.din(new_net_8129),
		.dout(new_net_8130)
	);

	bfr new_net_8131_bfr_after (
		.din(new_net_8130),
		.dout(new_net_8131)
	);

	bfr new_net_8132_bfr_after (
		.din(new_net_8131),
		.dout(new_net_8132)
	);

	bfr new_net_8133_bfr_after (
		.din(new_net_8132),
		.dout(new_net_8133)
	);

	bfr new_net_8134_bfr_after (
		.din(new_net_8133),
		.dout(new_net_8134)
	);

	bfr new_net_8135_bfr_after (
		.din(new_net_8134),
		.dout(new_net_8135)
	);

	bfr new_net_8136_bfr_after (
		.din(new_net_8135),
		.dout(new_net_8136)
	);

	bfr new_net_8137_bfr_after (
		.din(new_net_8136),
		.dout(new_net_8137)
	);

	bfr new_net_8138_bfr_after (
		.din(new_net_8137),
		.dout(new_net_8138)
	);

	bfr new_net_8139_bfr_after (
		.din(new_net_8138),
		.dout(new_net_8139)
	);

	bfr new_net_8140_bfr_after (
		.din(new_net_8139),
		.dout(new_net_8140)
	);

	spl2 _0627__v_fanout (
		.a(new_net_8140),
		.b(new_net_978),
		.c(new_net_979)
	);

	bfr new_net_8141_bfr_after (
		.din(_0344_),
		.dout(new_net_8141)
	);

	bfr new_net_8142_bfr_after (
		.din(new_net_8141),
		.dout(new_net_8142)
	);

	bfr new_net_8143_bfr_after (
		.din(new_net_8142),
		.dout(new_net_8143)
	);

	bfr new_net_8144_bfr_after (
		.din(new_net_8143),
		.dout(new_net_8144)
	);

	bfr new_net_8145_bfr_after (
		.din(new_net_8144),
		.dout(new_net_8145)
	);

	bfr new_net_8146_bfr_after (
		.din(new_net_8145),
		.dout(new_net_8146)
	);

	bfr new_net_8147_bfr_after (
		.din(new_net_8146),
		.dout(new_net_8147)
	);

	bfr new_net_8148_bfr_after (
		.din(new_net_8147),
		.dout(new_net_8148)
	);

	bfr new_net_8149_bfr_after (
		.din(new_net_8148),
		.dout(new_net_8149)
	);

	bfr new_net_8150_bfr_after (
		.din(new_net_8149),
		.dout(new_net_8150)
	);

	bfr new_net_8151_bfr_after (
		.din(new_net_8150),
		.dout(new_net_8151)
	);

	bfr new_net_8152_bfr_after (
		.din(new_net_8151),
		.dout(new_net_8152)
	);

	bfr new_net_8153_bfr_after (
		.din(new_net_8152),
		.dout(new_net_8153)
	);

	bfr new_net_8154_bfr_after (
		.din(new_net_8153),
		.dout(new_net_8154)
	);

	bfr new_net_8155_bfr_after (
		.din(new_net_8154),
		.dout(new_net_8155)
	);

	bfr new_net_8156_bfr_after (
		.din(new_net_8155),
		.dout(new_net_8156)
	);

	bfr new_net_8157_bfr_after (
		.din(new_net_8156),
		.dout(new_net_8157)
	);

	bfr new_net_8158_bfr_after (
		.din(new_net_8157),
		.dout(new_net_8158)
	);

	bfr new_net_8159_bfr_after (
		.din(new_net_8158),
		.dout(new_net_8159)
	);

	bfr new_net_8160_bfr_after (
		.din(new_net_8159),
		.dout(new_net_8160)
	);

	bfr new_net_8161_bfr_after (
		.din(new_net_8160),
		.dout(new_net_8161)
	);

	bfr new_net_8162_bfr_after (
		.din(new_net_8161),
		.dout(new_net_8162)
	);

	bfr new_net_8163_bfr_after (
		.din(new_net_8162),
		.dout(new_net_8163)
	);

	bfr new_net_8164_bfr_after (
		.din(new_net_8163),
		.dout(new_net_8164)
	);

	bfr new_net_8165_bfr_after (
		.din(new_net_8164),
		.dout(new_net_8165)
	);

	bfr new_net_8166_bfr_after (
		.din(new_net_8165),
		.dout(new_net_8166)
	);

	bfr new_net_8167_bfr_after (
		.din(new_net_8166),
		.dout(new_net_8167)
	);

	bfr new_net_8168_bfr_after (
		.din(new_net_8167),
		.dout(new_net_8168)
	);

	bfr new_net_8169_bfr_after (
		.din(new_net_8168),
		.dout(new_net_8169)
	);

	bfr new_net_8170_bfr_after (
		.din(new_net_8169),
		.dout(new_net_8170)
	);

	bfr new_net_8171_bfr_after (
		.din(new_net_8170),
		.dout(new_net_8171)
	);

	bfr new_net_8172_bfr_after (
		.din(new_net_8171),
		.dout(new_net_8172)
	);

	bfr new_net_8173_bfr_after (
		.din(new_net_8172),
		.dout(new_net_8173)
	);

	bfr new_net_8174_bfr_after (
		.din(new_net_8173),
		.dout(new_net_8174)
	);

	bfr new_net_8175_bfr_after (
		.din(new_net_8174),
		.dout(new_net_8175)
	);

	bfr new_net_8176_bfr_after (
		.din(new_net_8175),
		.dout(new_net_8176)
	);

	bfr new_net_8177_bfr_after (
		.din(new_net_8176),
		.dout(new_net_8177)
	);

	bfr new_net_8178_bfr_after (
		.din(new_net_8177),
		.dout(new_net_8178)
	);

	bfr new_net_8179_bfr_after (
		.din(new_net_8178),
		.dout(new_net_8179)
	);

	bfr new_net_8180_bfr_after (
		.din(new_net_8179),
		.dout(new_net_8180)
	);

	bfr new_net_8181_bfr_after (
		.din(new_net_8180),
		.dout(new_net_8181)
	);

	bfr new_net_8182_bfr_after (
		.din(new_net_8181),
		.dout(new_net_8182)
	);

	bfr new_net_8183_bfr_after (
		.din(new_net_8182),
		.dout(new_net_8183)
	);

	bfr new_net_8184_bfr_after (
		.din(new_net_8183),
		.dout(new_net_8184)
	);

	bfr new_net_8185_bfr_after (
		.din(new_net_8184),
		.dout(new_net_8185)
	);

	bfr new_net_8186_bfr_after (
		.din(new_net_8185),
		.dout(new_net_8186)
	);

	bfr new_net_8187_bfr_after (
		.din(new_net_8186),
		.dout(new_net_8187)
	);

	bfr new_net_8188_bfr_after (
		.din(new_net_8187),
		.dout(new_net_8188)
	);

	spl2 _0344__v_fanout (
		.a(new_net_8188),
		.b(new_net_1342),
		.c(new_net_1343)
	);

	bfr new_net_8189_bfr_after (
		.din(_0227_),
		.dout(new_net_8189)
	);

	bfr new_net_8190_bfr_after (
		.din(new_net_8189),
		.dout(new_net_8190)
	);

	bfr new_net_8191_bfr_after (
		.din(new_net_8190),
		.dout(new_net_8191)
	);

	bfr new_net_8192_bfr_after (
		.din(new_net_8191),
		.dout(new_net_8192)
	);

	bfr new_net_8193_bfr_after (
		.din(new_net_8192),
		.dout(new_net_8193)
	);

	bfr new_net_8194_bfr_after (
		.din(new_net_8193),
		.dout(new_net_8194)
	);

	bfr new_net_8195_bfr_after (
		.din(new_net_8194),
		.dout(new_net_8195)
	);

	bfr new_net_8196_bfr_after (
		.din(new_net_8195),
		.dout(new_net_8196)
	);

	bfr new_net_8197_bfr_after (
		.din(new_net_8196),
		.dout(new_net_8197)
	);

	bfr new_net_8198_bfr_after (
		.din(new_net_8197),
		.dout(new_net_8198)
	);

	bfr new_net_8199_bfr_after (
		.din(new_net_8198),
		.dout(new_net_8199)
	);

	bfr new_net_8200_bfr_after (
		.din(new_net_8199),
		.dout(new_net_8200)
	);

	bfr new_net_8201_bfr_after (
		.din(new_net_8200),
		.dout(new_net_8201)
	);

	bfr new_net_8202_bfr_after (
		.din(new_net_8201),
		.dout(new_net_8202)
	);

	bfr new_net_8203_bfr_after (
		.din(new_net_8202),
		.dout(new_net_8203)
	);

	bfr new_net_8204_bfr_after (
		.din(new_net_8203),
		.dout(new_net_8204)
	);

	bfr new_net_8205_bfr_after (
		.din(new_net_8204),
		.dout(new_net_8205)
	);

	bfr new_net_8206_bfr_after (
		.din(new_net_8205),
		.dout(new_net_8206)
	);

	bfr new_net_8207_bfr_after (
		.din(new_net_8206),
		.dout(new_net_8207)
	);

	bfr new_net_8208_bfr_after (
		.din(new_net_8207),
		.dout(new_net_8208)
	);

	bfr new_net_8209_bfr_after (
		.din(new_net_8208),
		.dout(new_net_8209)
	);

	bfr new_net_8210_bfr_after (
		.din(new_net_8209),
		.dout(new_net_8210)
	);

	bfr new_net_8211_bfr_after (
		.din(new_net_8210),
		.dout(new_net_8211)
	);

	bfr new_net_8212_bfr_after (
		.din(new_net_8211),
		.dout(new_net_8212)
	);

	bfr new_net_8213_bfr_after (
		.din(new_net_8212),
		.dout(new_net_8213)
	);

	bfr new_net_8214_bfr_after (
		.din(new_net_8213),
		.dout(new_net_8214)
	);

	bfr new_net_8215_bfr_after (
		.din(new_net_8214),
		.dout(new_net_8215)
	);

	bfr new_net_8216_bfr_after (
		.din(new_net_8215),
		.dout(new_net_8216)
	);

	bfr new_net_8217_bfr_after (
		.din(new_net_8216),
		.dout(new_net_8217)
	);

	bfr new_net_8218_bfr_after (
		.din(new_net_8217),
		.dout(new_net_8218)
	);

	bfr new_net_8219_bfr_after (
		.din(new_net_8218),
		.dout(new_net_8219)
	);

	bfr new_net_8220_bfr_after (
		.din(new_net_8219),
		.dout(new_net_8220)
	);

	bfr new_net_8221_bfr_after (
		.din(new_net_8220),
		.dout(new_net_8221)
	);

	bfr new_net_8222_bfr_after (
		.din(new_net_8221),
		.dout(new_net_8222)
	);

	bfr new_net_8223_bfr_after (
		.din(new_net_8222),
		.dout(new_net_8223)
	);

	bfr new_net_8224_bfr_after (
		.din(new_net_8223),
		.dout(new_net_8224)
	);

	bfr new_net_8225_bfr_after (
		.din(new_net_8224),
		.dout(new_net_8225)
	);

	bfr new_net_8226_bfr_after (
		.din(new_net_8225),
		.dout(new_net_8226)
	);

	bfr new_net_8227_bfr_after (
		.din(new_net_8226),
		.dout(new_net_8227)
	);

	bfr new_net_8228_bfr_after (
		.din(new_net_8227),
		.dout(new_net_8228)
	);

	bfr new_net_8229_bfr_after (
		.din(new_net_8228),
		.dout(new_net_8229)
	);

	bfr new_net_8230_bfr_after (
		.din(new_net_8229),
		.dout(new_net_8230)
	);

	bfr new_net_8231_bfr_after (
		.din(new_net_8230),
		.dout(new_net_8231)
	);

	bfr new_net_8232_bfr_after (
		.din(new_net_8231),
		.dout(new_net_8232)
	);

	bfr new_net_8233_bfr_after (
		.din(new_net_8232),
		.dout(new_net_8233)
	);

	bfr new_net_8234_bfr_after (
		.din(new_net_8233),
		.dout(new_net_8234)
	);

	bfr new_net_8235_bfr_after (
		.din(new_net_8234),
		.dout(new_net_8235)
	);

	bfr new_net_8236_bfr_after (
		.din(new_net_8235),
		.dout(new_net_8236)
	);

	bfr new_net_8237_bfr_after (
		.din(new_net_8236),
		.dout(new_net_8237)
	);

	bfr new_net_8238_bfr_after (
		.din(new_net_8237),
		.dout(new_net_8238)
	);

	bfr new_net_8239_bfr_after (
		.din(new_net_8238),
		.dout(new_net_8239)
	);

	bfr new_net_8240_bfr_after (
		.din(new_net_8239),
		.dout(new_net_8240)
	);

	bfr new_net_8241_bfr_after (
		.din(new_net_8240),
		.dout(new_net_8241)
	);

	bfr new_net_8242_bfr_after (
		.din(new_net_8241),
		.dout(new_net_8242)
	);

	bfr new_net_8243_bfr_after (
		.din(new_net_8242),
		.dout(new_net_8243)
	);

	bfr new_net_8244_bfr_after (
		.din(new_net_8243),
		.dout(new_net_8244)
	);

	spl2 _0227__v_fanout (
		.a(new_net_8244),
		.b(new_net_118),
		.c(new_net_119)
	);

	bfr new_net_8245_bfr_after (
		.din(_0296_),
		.dout(new_net_8245)
	);

	bfr new_net_8246_bfr_after (
		.din(new_net_8245),
		.dout(new_net_8246)
	);

	bfr new_net_8247_bfr_after (
		.din(new_net_8246),
		.dout(new_net_8247)
	);

	bfr new_net_8248_bfr_after (
		.din(new_net_8247),
		.dout(new_net_8248)
	);

	bfr new_net_8249_bfr_after (
		.din(new_net_8248),
		.dout(new_net_8249)
	);

	bfr new_net_8250_bfr_after (
		.din(new_net_8249),
		.dout(new_net_8250)
	);

	bfr new_net_8251_bfr_after (
		.din(new_net_8250),
		.dout(new_net_8251)
	);

	bfr new_net_8252_bfr_after (
		.din(new_net_8251),
		.dout(new_net_8252)
	);

	bfr new_net_8253_bfr_after (
		.din(new_net_8252),
		.dout(new_net_8253)
	);

	bfr new_net_8254_bfr_after (
		.din(new_net_8253),
		.dout(new_net_8254)
	);

	bfr new_net_8255_bfr_after (
		.din(new_net_8254),
		.dout(new_net_8255)
	);

	bfr new_net_8256_bfr_after (
		.din(new_net_8255),
		.dout(new_net_8256)
	);

	bfr new_net_8257_bfr_after (
		.din(new_net_8256),
		.dout(new_net_8257)
	);

	bfr new_net_8258_bfr_after (
		.din(new_net_8257),
		.dout(new_net_8258)
	);

	bfr new_net_8259_bfr_after (
		.din(new_net_8258),
		.dout(new_net_8259)
	);

	bfr new_net_8260_bfr_after (
		.din(new_net_8259),
		.dout(new_net_8260)
	);

	bfr new_net_8261_bfr_after (
		.din(new_net_8260),
		.dout(new_net_8261)
	);

	bfr new_net_8262_bfr_after (
		.din(new_net_8261),
		.dout(new_net_8262)
	);

	bfr new_net_8263_bfr_after (
		.din(new_net_8262),
		.dout(new_net_8263)
	);

	bfr new_net_8264_bfr_after (
		.din(new_net_8263),
		.dout(new_net_8264)
	);

	bfr new_net_8265_bfr_after (
		.din(new_net_8264),
		.dout(new_net_8265)
	);

	bfr new_net_8266_bfr_after (
		.din(new_net_8265),
		.dout(new_net_8266)
	);

	bfr new_net_8267_bfr_after (
		.din(new_net_8266),
		.dout(new_net_8267)
	);

	bfr new_net_8268_bfr_after (
		.din(new_net_8267),
		.dout(new_net_8268)
	);

	spl2 _0296__v_fanout (
		.a(new_net_8268),
		.b(new_net_2759),
		.c(new_net_2760)
	);

	bfr new_net_8269_bfr_after (
		.din(_0234_),
		.dout(new_net_8269)
	);

	bfr new_net_8270_bfr_after (
		.din(new_net_8269),
		.dout(new_net_8270)
	);

	bfr new_net_8271_bfr_after (
		.din(new_net_8270),
		.dout(new_net_8271)
	);

	bfr new_net_8272_bfr_after (
		.din(new_net_8271),
		.dout(new_net_8272)
	);

	bfr new_net_8273_bfr_after (
		.din(new_net_8272),
		.dout(new_net_8273)
	);

	bfr new_net_8274_bfr_after (
		.din(new_net_8273),
		.dout(new_net_8274)
	);

	bfr new_net_8275_bfr_after (
		.din(new_net_8274),
		.dout(new_net_8275)
	);

	bfr new_net_8276_bfr_after (
		.din(new_net_8275),
		.dout(new_net_8276)
	);

	bfr new_net_8277_bfr_after (
		.din(new_net_8276),
		.dout(new_net_8277)
	);

	bfr new_net_8278_bfr_after (
		.din(new_net_8277),
		.dout(new_net_8278)
	);

	bfr new_net_8279_bfr_after (
		.din(new_net_8278),
		.dout(new_net_8279)
	);

	bfr new_net_8280_bfr_after (
		.din(new_net_8279),
		.dout(new_net_8280)
	);

	bfr new_net_8281_bfr_after (
		.din(new_net_8280),
		.dout(new_net_8281)
	);

	bfr new_net_8282_bfr_after (
		.din(new_net_8281),
		.dout(new_net_8282)
	);

	bfr new_net_8283_bfr_after (
		.din(new_net_8282),
		.dout(new_net_8283)
	);

	bfr new_net_8284_bfr_after (
		.din(new_net_8283),
		.dout(new_net_8284)
	);

	bfr new_net_8285_bfr_after (
		.din(new_net_8284),
		.dout(new_net_8285)
	);

	bfr new_net_8286_bfr_after (
		.din(new_net_8285),
		.dout(new_net_8286)
	);

	bfr new_net_8287_bfr_after (
		.din(new_net_8286),
		.dout(new_net_8287)
	);

	bfr new_net_8288_bfr_after (
		.din(new_net_8287),
		.dout(new_net_8288)
	);

	bfr new_net_8289_bfr_after (
		.din(new_net_8288),
		.dout(new_net_8289)
	);

	bfr new_net_8290_bfr_after (
		.din(new_net_8289),
		.dout(new_net_8290)
	);

	bfr new_net_8291_bfr_after (
		.din(new_net_8290),
		.dout(new_net_8291)
	);

	bfr new_net_8292_bfr_after (
		.din(new_net_8291),
		.dout(new_net_8292)
	);

	bfr new_net_8293_bfr_after (
		.din(new_net_8292),
		.dout(new_net_8293)
	);

	bfr new_net_8294_bfr_after (
		.din(new_net_8293),
		.dout(new_net_8294)
	);

	bfr new_net_8295_bfr_after (
		.din(new_net_8294),
		.dout(new_net_8295)
	);

	bfr new_net_8296_bfr_after (
		.din(new_net_8295),
		.dout(new_net_8296)
	);

	bfr new_net_8297_bfr_after (
		.din(new_net_8296),
		.dout(new_net_8297)
	);

	bfr new_net_8298_bfr_after (
		.din(new_net_8297),
		.dout(new_net_8298)
	);

	spl2 _0234__v_fanout (
		.a(new_net_8298),
		.b(new_net_364),
		.c(new_net_365)
	);

	bfr new_net_8299_bfr_after (
		.din(_0212_),
		.dout(new_net_8299)
	);

	bfr new_net_8300_bfr_after (
		.din(new_net_8299),
		.dout(new_net_8300)
	);

	bfr new_net_8301_bfr_after (
		.din(new_net_8300),
		.dout(new_net_8301)
	);

	bfr new_net_8302_bfr_after (
		.din(new_net_8301),
		.dout(new_net_8302)
	);

	bfr new_net_8303_bfr_after (
		.din(new_net_8302),
		.dout(new_net_8303)
	);

	bfr new_net_8304_bfr_after (
		.din(new_net_8303),
		.dout(new_net_8304)
	);

	bfr new_net_8305_bfr_after (
		.din(new_net_8304),
		.dout(new_net_8305)
	);

	bfr new_net_8306_bfr_after (
		.din(new_net_8305),
		.dout(new_net_8306)
	);

	bfr new_net_8307_bfr_after (
		.din(new_net_8306),
		.dout(new_net_8307)
	);

	bfr new_net_8308_bfr_after (
		.din(new_net_8307),
		.dout(new_net_8308)
	);

	bfr new_net_8309_bfr_after (
		.din(new_net_8308),
		.dout(new_net_8309)
	);

	bfr new_net_8310_bfr_after (
		.din(new_net_8309),
		.dout(new_net_8310)
	);

	bfr new_net_8311_bfr_after (
		.din(new_net_8310),
		.dout(new_net_8311)
	);

	bfr new_net_8312_bfr_after (
		.din(new_net_8311),
		.dout(new_net_8312)
	);

	bfr new_net_8313_bfr_after (
		.din(new_net_8312),
		.dout(new_net_8313)
	);

	bfr new_net_8314_bfr_after (
		.din(new_net_8313),
		.dout(new_net_8314)
	);

	bfr new_net_8315_bfr_after (
		.din(new_net_8314),
		.dout(new_net_8315)
	);

	bfr new_net_8316_bfr_after (
		.din(new_net_8315),
		.dout(new_net_8316)
	);

	bfr new_net_8317_bfr_after (
		.din(new_net_8316),
		.dout(new_net_8317)
	);

	bfr new_net_8318_bfr_after (
		.din(new_net_8317),
		.dout(new_net_8318)
	);

	bfr new_net_8319_bfr_after (
		.din(new_net_8318),
		.dout(new_net_8319)
	);

	bfr new_net_8320_bfr_after (
		.din(new_net_8319),
		.dout(new_net_8320)
	);

	bfr new_net_8321_bfr_after (
		.din(new_net_8320),
		.dout(new_net_8321)
	);

	bfr new_net_8322_bfr_after (
		.din(new_net_8321),
		.dout(new_net_8322)
	);

	bfr new_net_8323_bfr_after (
		.din(new_net_8322),
		.dout(new_net_8323)
	);

	bfr new_net_8324_bfr_after (
		.din(new_net_8323),
		.dout(new_net_8324)
	);

	bfr new_net_8325_bfr_after (
		.din(new_net_8324),
		.dout(new_net_8325)
	);

	bfr new_net_8326_bfr_after (
		.din(new_net_8325),
		.dout(new_net_8326)
	);

	bfr new_net_8327_bfr_after (
		.din(new_net_8326),
		.dout(new_net_8327)
	);

	bfr new_net_8328_bfr_after (
		.din(new_net_8327),
		.dout(new_net_8328)
	);

	bfr new_net_8329_bfr_after (
		.din(new_net_8328),
		.dout(new_net_8329)
	);

	bfr new_net_8330_bfr_after (
		.din(new_net_8329),
		.dout(new_net_8330)
	);

	bfr new_net_8331_bfr_after (
		.din(new_net_8330),
		.dout(new_net_8331)
	);

	bfr new_net_8332_bfr_after (
		.din(new_net_8331),
		.dout(new_net_8332)
	);

	bfr new_net_8333_bfr_after (
		.din(new_net_8332),
		.dout(new_net_8333)
	);

	bfr new_net_8334_bfr_after (
		.din(new_net_8333),
		.dout(new_net_8334)
	);

	bfr new_net_8335_bfr_after (
		.din(new_net_8334),
		.dout(new_net_8335)
	);

	bfr new_net_8336_bfr_after (
		.din(new_net_8335),
		.dout(new_net_8336)
	);

	bfr new_net_8337_bfr_after (
		.din(new_net_8336),
		.dout(new_net_8337)
	);

	bfr new_net_8338_bfr_after (
		.din(new_net_8337),
		.dout(new_net_8338)
	);

	bfr new_net_8339_bfr_after (
		.din(new_net_8338),
		.dout(new_net_8339)
	);

	bfr new_net_8340_bfr_after (
		.din(new_net_8339),
		.dout(new_net_8340)
	);

	bfr new_net_8341_bfr_after (
		.din(new_net_8340),
		.dout(new_net_8341)
	);

	bfr new_net_8342_bfr_after (
		.din(new_net_8341),
		.dout(new_net_8342)
	);

	bfr new_net_8343_bfr_after (
		.din(new_net_8342),
		.dout(new_net_8343)
	);

	bfr new_net_8344_bfr_after (
		.din(new_net_8343),
		.dout(new_net_8344)
	);

	bfr new_net_8345_bfr_after (
		.din(new_net_8344),
		.dout(new_net_8345)
	);

	bfr new_net_8346_bfr_after (
		.din(new_net_8345),
		.dout(new_net_8346)
	);

	bfr new_net_8347_bfr_after (
		.din(new_net_8346),
		.dout(new_net_8347)
	);

	bfr new_net_8348_bfr_after (
		.din(new_net_8347),
		.dout(new_net_8348)
	);

	bfr new_net_8349_bfr_after (
		.din(new_net_8348),
		.dout(new_net_8349)
	);

	bfr new_net_8350_bfr_after (
		.din(new_net_8349),
		.dout(new_net_8350)
	);

	bfr new_net_8351_bfr_after (
		.din(new_net_8350),
		.dout(new_net_8351)
	);

	bfr new_net_8352_bfr_after (
		.din(new_net_8351),
		.dout(new_net_8352)
	);

	bfr new_net_8353_bfr_after (
		.din(new_net_8352),
		.dout(new_net_8353)
	);

	bfr new_net_8354_bfr_after (
		.din(new_net_8353),
		.dout(new_net_8354)
	);

	bfr new_net_8355_bfr_after (
		.din(new_net_8354),
		.dout(new_net_8355)
	);

	bfr new_net_8356_bfr_after (
		.din(new_net_8355),
		.dout(new_net_8356)
	);

	bfr new_net_8357_bfr_after (
		.din(new_net_8356),
		.dout(new_net_8357)
	);

	bfr new_net_8358_bfr_after (
		.din(new_net_8357),
		.dout(new_net_8358)
	);

	bfr new_net_8359_bfr_after (
		.din(new_net_8358),
		.dout(new_net_8359)
	);

	bfr new_net_8360_bfr_after (
		.din(new_net_8359),
		.dout(new_net_8360)
	);

	bfr new_net_8361_bfr_after (
		.din(new_net_8360),
		.dout(new_net_8361)
	);

	bfr new_net_8362_bfr_after (
		.din(new_net_8361),
		.dout(new_net_8362)
	);

	bfr new_net_8363_bfr_after (
		.din(new_net_8362),
		.dout(new_net_8363)
	);

	bfr new_net_8364_bfr_after (
		.din(new_net_8363),
		.dout(new_net_8364)
	);

	bfr new_net_8365_bfr_after (
		.din(new_net_8364),
		.dout(new_net_8365)
	);

	bfr new_net_8366_bfr_after (
		.din(new_net_8365),
		.dout(new_net_8366)
	);

	bfr new_net_8367_bfr_after (
		.din(new_net_8366),
		.dout(new_net_8367)
	);

	bfr new_net_8368_bfr_after (
		.din(new_net_8367),
		.dout(new_net_8368)
	);

	bfr new_net_8369_bfr_after (
		.din(new_net_8368),
		.dout(new_net_8369)
	);

	bfr new_net_8370_bfr_after (
		.din(new_net_8369),
		.dout(new_net_8370)
	);

	bfr new_net_8371_bfr_after (
		.din(new_net_8370),
		.dout(new_net_8371)
	);

	bfr new_net_8372_bfr_after (
		.din(new_net_8371),
		.dout(new_net_8372)
	);

	bfr new_net_8373_bfr_after (
		.din(new_net_8372),
		.dout(new_net_8373)
	);

	bfr new_net_8374_bfr_after (
		.din(new_net_8373),
		.dout(new_net_8374)
	);

	bfr new_net_8375_bfr_after (
		.din(new_net_8374),
		.dout(new_net_8375)
	);

	bfr new_net_8376_bfr_after (
		.din(new_net_8375),
		.dout(new_net_8376)
	);

	bfr new_net_8377_bfr_after (
		.din(new_net_8376),
		.dout(new_net_8377)
	);

	bfr new_net_8378_bfr_after (
		.din(new_net_8377),
		.dout(new_net_8378)
	);

	bfr new_net_8379_bfr_after (
		.din(new_net_8378),
		.dout(new_net_8379)
	);

	bfr new_net_8380_bfr_after (
		.din(new_net_8379),
		.dout(new_net_8380)
	);

	bfr new_net_8381_bfr_after (
		.din(new_net_8380),
		.dout(new_net_8381)
	);

	bfr new_net_8382_bfr_after (
		.din(new_net_8381),
		.dout(new_net_8382)
	);

	bfr new_net_8383_bfr_after (
		.din(new_net_8382),
		.dout(new_net_8383)
	);

	bfr new_net_8384_bfr_after (
		.din(new_net_8383),
		.dout(new_net_8384)
	);

	bfr new_net_8385_bfr_after (
		.din(new_net_8384),
		.dout(new_net_8385)
	);

	bfr new_net_8386_bfr_after (
		.din(new_net_8385),
		.dout(new_net_8386)
	);

	bfr new_net_8387_bfr_after (
		.din(new_net_8386),
		.dout(new_net_8387)
	);

	bfr new_net_8388_bfr_after (
		.din(new_net_8387),
		.dout(new_net_8388)
	);

	bfr new_net_8389_bfr_after (
		.din(new_net_8388),
		.dout(new_net_8389)
	);

	bfr new_net_8390_bfr_after (
		.din(new_net_8389),
		.dout(new_net_8390)
	);

	bfr new_net_8391_bfr_after (
		.din(new_net_8390),
		.dout(new_net_8391)
	);

	bfr new_net_8392_bfr_after (
		.din(new_net_8391),
		.dout(new_net_8392)
	);

	bfr new_net_8393_bfr_after (
		.din(new_net_8392),
		.dout(new_net_8393)
	);

	bfr new_net_8394_bfr_after (
		.din(new_net_8393),
		.dout(new_net_8394)
	);

	bfr new_net_8395_bfr_after (
		.din(new_net_8394),
		.dout(new_net_8395)
	);

	bfr new_net_8396_bfr_after (
		.din(new_net_8395),
		.dout(new_net_8396)
	);

	bfr new_net_8397_bfr_after (
		.din(new_net_8396),
		.dout(new_net_8397)
	);

	bfr new_net_8398_bfr_after (
		.din(new_net_8397),
		.dout(new_net_8398)
	);

	bfr new_net_8399_bfr_after (
		.din(new_net_8398),
		.dout(new_net_8399)
	);

	bfr new_net_8400_bfr_after (
		.din(new_net_8399),
		.dout(new_net_8400)
	);

	bfr new_net_8401_bfr_after (
		.din(new_net_8400),
		.dout(new_net_8401)
	);

	bfr new_net_8402_bfr_after (
		.din(new_net_8401),
		.dout(new_net_8402)
	);

	bfr new_net_8403_bfr_after (
		.din(new_net_8402),
		.dout(new_net_8403)
	);

	bfr new_net_8404_bfr_after (
		.din(new_net_8403),
		.dout(new_net_8404)
	);

	bfr new_net_8405_bfr_after (
		.din(new_net_8404),
		.dout(new_net_8405)
	);

	bfr new_net_8406_bfr_after (
		.din(new_net_8405),
		.dout(new_net_8406)
	);

	bfr new_net_8407_bfr_after (
		.din(new_net_8406),
		.dout(new_net_8407)
	);

	bfr new_net_8408_bfr_after (
		.din(new_net_8407),
		.dout(new_net_8408)
	);

	bfr new_net_8409_bfr_after (
		.din(new_net_8408),
		.dout(new_net_8409)
	);

	bfr new_net_8410_bfr_after (
		.din(new_net_8409),
		.dout(new_net_8410)
	);

	spl2 _0212__v_fanout (
		.a(new_net_8410),
		.b(new_net_2752),
		.c(new_net_2753)
	);

	bfr new_net_8411_bfr_after (
		.din(_0625_),
		.dout(new_net_8411)
	);

	bfr new_net_8412_bfr_after (
		.din(new_net_8411),
		.dout(new_net_8412)
	);

	bfr new_net_8413_bfr_after (
		.din(new_net_8412),
		.dout(new_net_8413)
	);

	bfr new_net_8414_bfr_after (
		.din(new_net_8413),
		.dout(new_net_8414)
	);

	bfr new_net_8415_bfr_after (
		.din(new_net_8414),
		.dout(new_net_8415)
	);

	bfr new_net_8416_bfr_after (
		.din(new_net_8415),
		.dout(new_net_8416)
	);

	bfr new_net_8417_bfr_after (
		.din(new_net_8416),
		.dout(new_net_8417)
	);

	bfr new_net_8418_bfr_after (
		.din(new_net_8417),
		.dout(new_net_8418)
	);

	bfr new_net_8419_bfr_after (
		.din(new_net_8418),
		.dout(new_net_8419)
	);

	bfr new_net_8420_bfr_after (
		.din(new_net_8419),
		.dout(new_net_8420)
	);

	bfr new_net_8421_bfr_after (
		.din(new_net_8420),
		.dout(new_net_8421)
	);

	bfr new_net_8422_bfr_after (
		.din(new_net_8421),
		.dout(new_net_8422)
	);

	bfr new_net_8423_bfr_after (
		.din(new_net_8422),
		.dout(new_net_8423)
	);

	bfr new_net_8424_bfr_after (
		.din(new_net_8423),
		.dout(new_net_8424)
	);

	bfr new_net_8425_bfr_after (
		.din(new_net_8424),
		.dout(new_net_8425)
	);

	bfr new_net_8426_bfr_after (
		.din(new_net_8425),
		.dout(new_net_8426)
	);

	bfr new_net_8427_bfr_after (
		.din(new_net_8426),
		.dout(new_net_8427)
	);

	bfr new_net_8428_bfr_after (
		.din(new_net_8427),
		.dout(new_net_8428)
	);

	bfr new_net_8429_bfr_after (
		.din(new_net_8428),
		.dout(new_net_8429)
	);

	bfr new_net_8430_bfr_after (
		.din(new_net_8429),
		.dout(new_net_8430)
	);

	bfr new_net_8431_bfr_after (
		.din(new_net_8430),
		.dout(new_net_8431)
	);

	bfr new_net_8432_bfr_after (
		.din(new_net_8431),
		.dout(new_net_8432)
	);

	bfr new_net_8433_bfr_after (
		.din(new_net_8432),
		.dout(new_net_8433)
	);

	bfr new_net_8434_bfr_after (
		.din(new_net_8433),
		.dout(new_net_8434)
	);

	bfr new_net_8435_bfr_after (
		.din(new_net_8434),
		.dout(new_net_8435)
	);

	bfr new_net_8436_bfr_after (
		.din(new_net_8435),
		.dout(new_net_8436)
	);

	bfr new_net_8437_bfr_after (
		.din(new_net_8436),
		.dout(new_net_8437)
	);

	bfr new_net_8438_bfr_after (
		.din(new_net_8437),
		.dout(new_net_8438)
	);

	bfr new_net_8439_bfr_after (
		.din(new_net_8438),
		.dout(new_net_8439)
	);

	bfr new_net_8440_bfr_after (
		.din(new_net_8439),
		.dout(new_net_8440)
	);

	bfr new_net_8441_bfr_after (
		.din(new_net_8440),
		.dout(new_net_8441)
	);

	bfr new_net_8442_bfr_after (
		.din(new_net_8441),
		.dout(new_net_8442)
	);

	bfr new_net_8443_bfr_after (
		.din(new_net_8442),
		.dout(new_net_8443)
	);

	bfr new_net_8444_bfr_after (
		.din(new_net_8443),
		.dout(new_net_8444)
	);

	bfr new_net_8445_bfr_after (
		.din(new_net_8444),
		.dout(new_net_8445)
	);

	bfr new_net_8446_bfr_after (
		.din(new_net_8445),
		.dout(new_net_8446)
	);

	bfr new_net_8447_bfr_after (
		.din(new_net_8446),
		.dout(new_net_8447)
	);

	bfr new_net_8448_bfr_after (
		.din(new_net_8447),
		.dout(new_net_8448)
	);

	bfr new_net_8449_bfr_after (
		.din(new_net_8448),
		.dout(new_net_8449)
	);

	bfr new_net_8450_bfr_after (
		.din(new_net_8449),
		.dout(new_net_8450)
	);

	bfr new_net_8451_bfr_after (
		.din(new_net_8450),
		.dout(new_net_8451)
	);

	bfr new_net_8452_bfr_after (
		.din(new_net_8451),
		.dout(new_net_8452)
	);

	bfr new_net_8453_bfr_after (
		.din(new_net_8452),
		.dout(new_net_8453)
	);

	bfr new_net_8454_bfr_after (
		.din(new_net_8453),
		.dout(new_net_8454)
	);

	bfr new_net_8455_bfr_after (
		.din(new_net_8454),
		.dout(new_net_8455)
	);

	bfr new_net_8456_bfr_after (
		.din(new_net_8455),
		.dout(new_net_8456)
	);

	bfr new_net_8457_bfr_after (
		.din(new_net_8456),
		.dout(new_net_8457)
	);

	bfr new_net_8458_bfr_after (
		.din(new_net_8457),
		.dout(new_net_8458)
	);

	bfr new_net_8459_bfr_after (
		.din(new_net_8458),
		.dout(new_net_8459)
	);

	bfr new_net_8460_bfr_after (
		.din(new_net_8459),
		.dout(new_net_8460)
	);

	bfr new_net_8461_bfr_after (
		.din(new_net_8460),
		.dout(new_net_8461)
	);

	bfr new_net_8462_bfr_after (
		.din(new_net_8461),
		.dout(new_net_8462)
	);

	bfr new_net_8463_bfr_after (
		.din(new_net_8462),
		.dout(new_net_8463)
	);

	bfr new_net_8464_bfr_after (
		.din(new_net_8463),
		.dout(new_net_8464)
	);

	bfr new_net_8465_bfr_after (
		.din(new_net_8464),
		.dout(new_net_8465)
	);

	bfr new_net_8466_bfr_after (
		.din(new_net_8465),
		.dout(new_net_8466)
	);

	bfr new_net_8467_bfr_after (
		.din(new_net_8466),
		.dout(new_net_8467)
	);

	bfr new_net_8468_bfr_after (
		.din(new_net_8467),
		.dout(new_net_8468)
	);

	bfr new_net_8469_bfr_after (
		.din(new_net_8468),
		.dout(new_net_8469)
	);

	bfr new_net_8470_bfr_after (
		.din(new_net_8469),
		.dout(new_net_8470)
	);

	bfr new_net_8471_bfr_after (
		.din(new_net_8470),
		.dout(new_net_8471)
	);

	bfr new_net_8472_bfr_after (
		.din(new_net_8471),
		.dout(new_net_8472)
	);

	bfr new_net_8473_bfr_after (
		.din(new_net_8472),
		.dout(new_net_8473)
	);

	bfr new_net_8474_bfr_after (
		.din(new_net_8473),
		.dout(new_net_8474)
	);

	bfr new_net_8475_bfr_after (
		.din(new_net_8474),
		.dout(new_net_8475)
	);

	bfr new_net_8476_bfr_after (
		.din(new_net_8475),
		.dout(new_net_8476)
	);

	bfr new_net_8477_bfr_after (
		.din(new_net_8476),
		.dout(new_net_8477)
	);

	bfr new_net_8478_bfr_after (
		.din(new_net_8477),
		.dout(new_net_8478)
	);

	bfr new_net_8479_bfr_after (
		.din(new_net_8478),
		.dout(new_net_8479)
	);

	bfr new_net_8480_bfr_after (
		.din(new_net_8479),
		.dout(new_net_8480)
	);

	bfr new_net_8481_bfr_after (
		.din(new_net_8480),
		.dout(new_net_8481)
	);

	bfr new_net_8482_bfr_after (
		.din(new_net_8481),
		.dout(new_net_8482)
	);

	bfr new_net_8483_bfr_after (
		.din(new_net_8482),
		.dout(new_net_8483)
	);

	bfr new_net_8484_bfr_after (
		.din(new_net_8483),
		.dout(new_net_8484)
	);

	bfr new_net_8485_bfr_after (
		.din(new_net_8484),
		.dout(new_net_8485)
	);

	bfr new_net_8486_bfr_after (
		.din(new_net_8485),
		.dout(new_net_8486)
	);

	bfr new_net_8487_bfr_after (
		.din(new_net_8486),
		.dout(new_net_8487)
	);

	bfr new_net_8488_bfr_after (
		.din(new_net_8487),
		.dout(new_net_8488)
	);

	bfr new_net_8489_bfr_after (
		.din(new_net_8488),
		.dout(new_net_8489)
	);

	bfr new_net_8490_bfr_after (
		.din(new_net_8489),
		.dout(new_net_8490)
	);

	spl2 _0625__v_fanout (
		.a(new_net_8490),
		.b(new_net_637),
		.c(new_net_638)
	);

	bfr new_net_8491_bfr_after (
		.din(_1292_),
		.dout(new_net_8491)
	);

	bfr new_net_8492_bfr_after (
		.din(new_net_8491),
		.dout(new_net_8492)
	);

	bfr new_net_8493_bfr_after (
		.din(new_net_8492),
		.dout(new_net_8493)
	);

	bfr new_net_8494_bfr_after (
		.din(new_net_8493),
		.dout(new_net_8494)
	);

	bfr new_net_8495_bfr_after (
		.din(new_net_8494),
		.dout(new_net_8495)
	);

	bfr new_net_8496_bfr_after (
		.din(new_net_8495),
		.dout(new_net_8496)
	);

	bfr new_net_8497_bfr_after (
		.din(new_net_8496),
		.dout(new_net_8497)
	);

	bfr new_net_8498_bfr_after (
		.din(new_net_8497),
		.dout(new_net_8498)
	);

	bfr new_net_8499_bfr_after (
		.din(new_net_8498),
		.dout(new_net_8499)
	);

	bfr new_net_8500_bfr_after (
		.din(new_net_8499),
		.dout(new_net_8500)
	);

	bfr new_net_8501_bfr_after (
		.din(new_net_8500),
		.dout(new_net_8501)
	);

	bfr new_net_8502_bfr_after (
		.din(new_net_8501),
		.dout(new_net_8502)
	);

	bfr new_net_8503_bfr_after (
		.din(new_net_8502),
		.dout(new_net_8503)
	);

	bfr new_net_8504_bfr_after (
		.din(new_net_8503),
		.dout(new_net_8504)
	);

	bfr new_net_8505_bfr_after (
		.din(new_net_8504),
		.dout(new_net_8505)
	);

	bfr new_net_8506_bfr_after (
		.din(new_net_8505),
		.dout(new_net_8506)
	);

	bfr new_net_8507_bfr_after (
		.din(new_net_8506),
		.dout(new_net_8507)
	);

	bfr new_net_8508_bfr_after (
		.din(new_net_8507),
		.dout(new_net_8508)
	);

	bfr new_net_8509_bfr_after (
		.din(new_net_8508),
		.dout(new_net_8509)
	);

	bfr new_net_8510_bfr_after (
		.din(new_net_8509),
		.dout(new_net_8510)
	);

	bfr new_net_8511_bfr_after (
		.din(new_net_8510),
		.dout(new_net_8511)
	);

	bfr new_net_8512_bfr_after (
		.din(new_net_8511),
		.dout(new_net_8512)
	);

	bfr new_net_8513_bfr_after (
		.din(new_net_8512),
		.dout(new_net_8513)
	);

	bfr new_net_8514_bfr_after (
		.din(new_net_8513),
		.dout(new_net_8514)
	);

	spl2 _1292__v_fanout (
		.a(new_net_8514),
		.b(new_net_699),
		.c(new_net_700)
	);

	bfr new_net_8515_bfr_after (
		.din(_0441_),
		.dout(new_net_8515)
	);

	bfr new_net_8516_bfr_after (
		.din(new_net_8515),
		.dout(new_net_8516)
	);

	bfr new_net_8517_bfr_after (
		.din(new_net_8516),
		.dout(new_net_8517)
	);

	bfr new_net_8518_bfr_after (
		.din(new_net_8517),
		.dout(new_net_8518)
	);

	bfr new_net_8519_bfr_after (
		.din(new_net_8518),
		.dout(new_net_8519)
	);

	bfr new_net_8520_bfr_after (
		.din(new_net_8519),
		.dout(new_net_8520)
	);

	bfr new_net_8521_bfr_after (
		.din(new_net_8520),
		.dout(new_net_8521)
	);

	bfr new_net_8522_bfr_after (
		.din(new_net_8521),
		.dout(new_net_8522)
	);

	bfr new_net_8523_bfr_after (
		.din(new_net_8522),
		.dout(new_net_8523)
	);

	bfr new_net_8524_bfr_after (
		.din(new_net_8523),
		.dout(new_net_8524)
	);

	bfr new_net_8525_bfr_after (
		.din(new_net_8524),
		.dout(new_net_8525)
	);

	bfr new_net_8526_bfr_after (
		.din(new_net_8525),
		.dout(new_net_8526)
	);

	bfr new_net_8527_bfr_after (
		.din(new_net_8526),
		.dout(new_net_8527)
	);

	bfr new_net_8528_bfr_after (
		.din(new_net_8527),
		.dout(new_net_8528)
	);

	bfr new_net_8529_bfr_after (
		.din(new_net_8528),
		.dout(new_net_8529)
	);

	bfr new_net_8530_bfr_after (
		.din(new_net_8529),
		.dout(new_net_8530)
	);

	bfr new_net_8531_bfr_after (
		.din(new_net_8530),
		.dout(new_net_8531)
	);

	bfr new_net_8532_bfr_after (
		.din(new_net_8531),
		.dout(new_net_8532)
	);

	bfr new_net_8533_bfr_after (
		.din(new_net_8532),
		.dout(new_net_8533)
	);

	bfr new_net_8534_bfr_after (
		.din(new_net_8533),
		.dout(new_net_8534)
	);

	bfr new_net_8535_bfr_after (
		.din(new_net_8534),
		.dout(new_net_8535)
	);

	bfr new_net_8536_bfr_after (
		.din(new_net_8535),
		.dout(new_net_8536)
	);

	bfr new_net_8537_bfr_after (
		.din(new_net_8536),
		.dout(new_net_8537)
	);

	bfr new_net_8538_bfr_after (
		.din(new_net_8537),
		.dout(new_net_8538)
	);

	bfr new_net_8539_bfr_after (
		.din(new_net_8538),
		.dout(new_net_8539)
	);

	bfr new_net_8540_bfr_after (
		.din(new_net_8539),
		.dout(new_net_8540)
	);

	bfr new_net_8541_bfr_after (
		.din(new_net_8540),
		.dout(new_net_8541)
	);

	bfr new_net_8542_bfr_after (
		.din(new_net_8541),
		.dout(new_net_8542)
	);

	bfr new_net_8543_bfr_after (
		.din(new_net_8542),
		.dout(new_net_8543)
	);

	bfr new_net_8544_bfr_after (
		.din(new_net_8543),
		.dout(new_net_8544)
	);

	bfr new_net_8545_bfr_after (
		.din(new_net_8544),
		.dout(new_net_8545)
	);

	bfr new_net_8546_bfr_after (
		.din(new_net_8545),
		.dout(new_net_8546)
	);

	bfr new_net_8547_bfr_after (
		.din(new_net_8546),
		.dout(new_net_8547)
	);

	bfr new_net_8548_bfr_after (
		.din(new_net_8547),
		.dout(new_net_8548)
	);

	bfr new_net_8549_bfr_after (
		.din(new_net_8548),
		.dout(new_net_8549)
	);

	bfr new_net_8550_bfr_after (
		.din(new_net_8549),
		.dout(new_net_8550)
	);

	bfr new_net_8551_bfr_after (
		.din(new_net_8550),
		.dout(new_net_8551)
	);

	bfr new_net_8552_bfr_after (
		.din(new_net_8551),
		.dout(new_net_8552)
	);

	bfr new_net_8553_bfr_after (
		.din(new_net_8552),
		.dout(new_net_8553)
	);

	bfr new_net_8554_bfr_after (
		.din(new_net_8553),
		.dout(new_net_8554)
	);

	bfr new_net_8555_bfr_after (
		.din(new_net_8554),
		.dout(new_net_8555)
	);

	bfr new_net_8556_bfr_after (
		.din(new_net_8555),
		.dout(new_net_8556)
	);

	bfr new_net_8557_bfr_after (
		.din(new_net_8556),
		.dout(new_net_8557)
	);

	bfr new_net_8558_bfr_after (
		.din(new_net_8557),
		.dout(new_net_8558)
	);

	bfr new_net_8559_bfr_after (
		.din(new_net_8558),
		.dout(new_net_8559)
	);

	bfr new_net_8560_bfr_after (
		.din(new_net_8559),
		.dout(new_net_8560)
	);

	bfr new_net_8561_bfr_after (
		.din(new_net_8560),
		.dout(new_net_8561)
	);

	bfr new_net_8562_bfr_after (
		.din(new_net_8561),
		.dout(new_net_8562)
	);

	bfr new_net_8563_bfr_after (
		.din(new_net_8562),
		.dout(new_net_8563)
	);

	bfr new_net_8564_bfr_after (
		.din(new_net_8563),
		.dout(new_net_8564)
	);

	bfr new_net_8565_bfr_after (
		.din(new_net_8564),
		.dout(new_net_8565)
	);

	bfr new_net_8566_bfr_after (
		.din(new_net_8565),
		.dout(new_net_8566)
	);

	bfr new_net_8567_bfr_after (
		.din(new_net_8566),
		.dout(new_net_8567)
	);

	bfr new_net_8568_bfr_after (
		.din(new_net_8567),
		.dout(new_net_8568)
	);

	bfr new_net_8569_bfr_after (
		.din(new_net_8568),
		.dout(new_net_8569)
	);

	bfr new_net_8570_bfr_after (
		.din(new_net_8569),
		.dout(new_net_8570)
	);

	bfr new_net_8571_bfr_after (
		.din(new_net_8570),
		.dout(new_net_8571)
	);

	bfr new_net_8572_bfr_after (
		.din(new_net_8571),
		.dout(new_net_8572)
	);

	bfr new_net_8573_bfr_after (
		.din(new_net_8572),
		.dout(new_net_8573)
	);

	bfr new_net_8574_bfr_after (
		.din(new_net_8573),
		.dout(new_net_8574)
	);

	bfr new_net_8575_bfr_after (
		.din(new_net_8574),
		.dout(new_net_8575)
	);

	bfr new_net_8576_bfr_after (
		.din(new_net_8575),
		.dout(new_net_8576)
	);

	bfr new_net_8577_bfr_after (
		.din(new_net_8576),
		.dout(new_net_8577)
	);

	bfr new_net_8578_bfr_after (
		.din(new_net_8577),
		.dout(new_net_8578)
	);

	bfr new_net_8579_bfr_after (
		.din(new_net_8578),
		.dout(new_net_8579)
	);

	bfr new_net_8580_bfr_after (
		.din(new_net_8579),
		.dout(new_net_8580)
	);

	bfr new_net_8581_bfr_after (
		.din(new_net_8580),
		.dout(new_net_8581)
	);

	bfr new_net_8582_bfr_after (
		.din(new_net_8581),
		.dout(new_net_8582)
	);

	bfr new_net_8583_bfr_after (
		.din(new_net_8582),
		.dout(new_net_8583)
	);

	bfr new_net_8584_bfr_after (
		.din(new_net_8583),
		.dout(new_net_8584)
	);

	bfr new_net_8585_bfr_after (
		.din(new_net_8584),
		.dout(new_net_8585)
	);

	bfr new_net_8586_bfr_after (
		.din(new_net_8585),
		.dout(new_net_8586)
	);

	bfr new_net_8587_bfr_after (
		.din(new_net_8586),
		.dout(new_net_8587)
	);

	bfr new_net_8588_bfr_after (
		.din(new_net_8587),
		.dout(new_net_8588)
	);

	bfr new_net_8589_bfr_after (
		.din(new_net_8588),
		.dout(new_net_8589)
	);

	bfr new_net_8590_bfr_after (
		.din(new_net_8589),
		.dout(new_net_8590)
	);

	bfr new_net_8591_bfr_after (
		.din(new_net_8590),
		.dout(new_net_8591)
	);

	bfr new_net_8592_bfr_after (
		.din(new_net_8591),
		.dout(new_net_8592)
	);

	bfr new_net_8593_bfr_after (
		.din(new_net_8592),
		.dout(new_net_8593)
	);

	bfr new_net_8594_bfr_after (
		.din(new_net_8593),
		.dout(new_net_8594)
	);

	spl2 _0441__v_fanout (
		.a(new_net_8594),
		.b(new_net_1302),
		.c(new_net_1303)
	);

	bfr new_net_8595_bfr_after (
		.din(_0112_),
		.dout(new_net_8595)
	);

	bfr new_net_8596_bfr_after (
		.din(new_net_8595),
		.dout(new_net_8596)
	);

	bfr new_net_8597_bfr_after (
		.din(new_net_8596),
		.dout(new_net_8597)
	);

	bfr new_net_8598_bfr_after (
		.din(new_net_8597),
		.dout(new_net_8598)
	);

	bfr new_net_8599_bfr_after (
		.din(new_net_8598),
		.dout(new_net_8599)
	);

	bfr new_net_8600_bfr_after (
		.din(new_net_8599),
		.dout(new_net_8600)
	);

	spl2 _0112__v_fanout (
		.a(new_net_8600),
		.b(new_net_3029),
		.c(new_net_3030)
	);

	bfr new_net_8601_bfr_after (
		.din(_1138_),
		.dout(new_net_8601)
	);

	bfr new_net_8602_bfr_after (
		.din(new_net_8601),
		.dout(new_net_8602)
	);

	bfr new_net_8603_bfr_after (
		.din(new_net_8602),
		.dout(new_net_8603)
	);

	bfr new_net_8604_bfr_after (
		.din(new_net_8603),
		.dout(new_net_8604)
	);

	bfr new_net_8605_bfr_after (
		.din(new_net_8604),
		.dout(new_net_8605)
	);

	bfr new_net_8606_bfr_after (
		.din(new_net_8605),
		.dout(new_net_8606)
	);

	bfr new_net_8607_bfr_after (
		.din(new_net_8606),
		.dout(new_net_8607)
	);

	bfr new_net_8608_bfr_after (
		.din(new_net_8607),
		.dout(new_net_8608)
	);

	bfr new_net_8609_bfr_after (
		.din(new_net_8608),
		.dout(new_net_8609)
	);

	bfr new_net_8610_bfr_after (
		.din(new_net_8609),
		.dout(new_net_8610)
	);

	bfr new_net_8611_bfr_after (
		.din(new_net_8610),
		.dout(new_net_8611)
	);

	bfr new_net_8612_bfr_after (
		.din(new_net_8611),
		.dout(new_net_8612)
	);

	bfr new_net_8613_bfr_after (
		.din(new_net_8612),
		.dout(new_net_8613)
	);

	bfr new_net_8614_bfr_after (
		.din(new_net_8613),
		.dout(new_net_8614)
	);

	bfr new_net_8615_bfr_after (
		.din(new_net_8614),
		.dout(new_net_8615)
	);

	bfr new_net_8616_bfr_after (
		.din(new_net_8615),
		.dout(new_net_8616)
	);

	bfr new_net_8617_bfr_after (
		.din(new_net_8616),
		.dout(new_net_8617)
	);

	bfr new_net_8618_bfr_after (
		.din(new_net_8617),
		.dout(new_net_8618)
	);

	bfr new_net_8619_bfr_after (
		.din(new_net_8618),
		.dout(new_net_8619)
	);

	bfr new_net_8620_bfr_after (
		.din(new_net_8619),
		.dout(new_net_8620)
	);

	bfr new_net_8621_bfr_after (
		.din(new_net_8620),
		.dout(new_net_8621)
	);

	bfr new_net_8622_bfr_after (
		.din(new_net_8621),
		.dout(new_net_8622)
	);

	bfr new_net_8623_bfr_after (
		.din(new_net_8622),
		.dout(new_net_8623)
	);

	bfr new_net_8624_bfr_after (
		.din(new_net_8623),
		.dout(new_net_8624)
	);

	spl2 _1138__v_fanout (
		.a(new_net_8624),
		.b(new_net_1178),
		.c(new_net_1179)
	);

	bfr new_net_8625_bfr_after (
		.din(_1282_),
		.dout(new_net_8625)
	);

	bfr new_net_8626_bfr_after (
		.din(new_net_8625),
		.dout(new_net_8626)
	);

	bfr new_net_8627_bfr_after (
		.din(new_net_8626),
		.dout(new_net_8627)
	);

	bfr new_net_8628_bfr_after (
		.din(new_net_8627),
		.dout(new_net_8628)
	);

	bfr new_net_8629_bfr_after (
		.din(new_net_8628),
		.dout(new_net_8629)
	);

	bfr new_net_8630_bfr_after (
		.din(new_net_8629),
		.dout(new_net_8630)
	);

	bfr new_net_8631_bfr_after (
		.din(new_net_8630),
		.dout(new_net_8631)
	);

	bfr new_net_8632_bfr_after (
		.din(new_net_8631),
		.dout(new_net_8632)
	);

	bfr new_net_8633_bfr_after (
		.din(new_net_8632),
		.dout(new_net_8633)
	);

	bfr new_net_8634_bfr_after (
		.din(new_net_8633),
		.dout(new_net_8634)
	);

	bfr new_net_8635_bfr_after (
		.din(new_net_8634),
		.dout(new_net_8635)
	);

	bfr new_net_8636_bfr_after (
		.din(new_net_8635),
		.dout(new_net_8636)
	);

	bfr new_net_8637_bfr_after (
		.din(new_net_8636),
		.dout(new_net_8637)
	);

	bfr new_net_8638_bfr_after (
		.din(new_net_8637),
		.dout(new_net_8638)
	);

	bfr new_net_8639_bfr_after (
		.din(new_net_8638),
		.dout(new_net_8639)
	);

	bfr new_net_8640_bfr_after (
		.din(new_net_8639),
		.dout(new_net_8640)
	);

	bfr new_net_8641_bfr_after (
		.din(new_net_8640),
		.dout(new_net_8641)
	);

	bfr new_net_8642_bfr_after (
		.din(new_net_8641),
		.dout(new_net_8642)
	);

	bfr new_net_8643_bfr_after (
		.din(new_net_8642),
		.dout(new_net_8643)
	);

	bfr new_net_8644_bfr_after (
		.din(new_net_8643),
		.dout(new_net_8644)
	);

	bfr new_net_8645_bfr_after (
		.din(new_net_8644),
		.dout(new_net_8645)
	);

	bfr new_net_8646_bfr_after (
		.din(new_net_8645),
		.dout(new_net_8646)
	);

	bfr new_net_8647_bfr_after (
		.din(new_net_8646),
		.dout(new_net_8647)
	);

	bfr new_net_8648_bfr_after (
		.din(new_net_8647),
		.dout(new_net_8648)
	);

	bfr new_net_8649_bfr_after (
		.din(new_net_8648),
		.dout(new_net_8649)
	);

	bfr new_net_8650_bfr_after (
		.din(new_net_8649),
		.dout(new_net_8650)
	);

	bfr new_net_8651_bfr_after (
		.din(new_net_8650),
		.dout(new_net_8651)
	);

	bfr new_net_8652_bfr_after (
		.din(new_net_8651),
		.dout(new_net_8652)
	);

	bfr new_net_8653_bfr_after (
		.din(new_net_8652),
		.dout(new_net_8653)
	);

	bfr new_net_8654_bfr_after (
		.din(new_net_8653),
		.dout(new_net_8654)
	);

	bfr new_net_8655_bfr_after (
		.din(new_net_8654),
		.dout(new_net_8655)
	);

	bfr new_net_8656_bfr_after (
		.din(new_net_8655),
		.dout(new_net_8656)
	);

	bfr new_net_8657_bfr_after (
		.din(new_net_8656),
		.dout(new_net_8657)
	);

	bfr new_net_8658_bfr_after (
		.din(new_net_8657),
		.dout(new_net_8658)
	);

	bfr new_net_8659_bfr_after (
		.din(new_net_8658),
		.dout(new_net_8659)
	);

	bfr new_net_8660_bfr_after (
		.din(new_net_8659),
		.dout(new_net_8660)
	);

	bfr new_net_8661_bfr_after (
		.din(new_net_8660),
		.dout(new_net_8661)
	);

	bfr new_net_8662_bfr_after (
		.din(new_net_8661),
		.dout(new_net_8662)
	);

	bfr new_net_8663_bfr_after (
		.din(new_net_8662),
		.dout(new_net_8663)
	);

	bfr new_net_8664_bfr_after (
		.din(new_net_8663),
		.dout(new_net_8664)
	);

	bfr new_net_8665_bfr_after (
		.din(new_net_8664),
		.dout(new_net_8665)
	);

	bfr new_net_8666_bfr_after (
		.din(new_net_8665),
		.dout(new_net_8666)
	);

	bfr new_net_8667_bfr_after (
		.din(new_net_8666),
		.dout(new_net_8667)
	);

	bfr new_net_8668_bfr_after (
		.din(new_net_8667),
		.dout(new_net_8668)
	);

	bfr new_net_8669_bfr_after (
		.din(new_net_8668),
		.dout(new_net_8669)
	);

	bfr new_net_8670_bfr_after (
		.din(new_net_8669),
		.dout(new_net_8670)
	);

	bfr new_net_8671_bfr_after (
		.din(new_net_8670),
		.dout(new_net_8671)
	);

	bfr new_net_8672_bfr_after (
		.din(new_net_8671),
		.dout(new_net_8672)
	);

	bfr new_net_8673_bfr_after (
		.din(new_net_8672),
		.dout(new_net_8673)
	);

	bfr new_net_8674_bfr_after (
		.din(new_net_8673),
		.dout(new_net_8674)
	);

	bfr new_net_8675_bfr_after (
		.din(new_net_8674),
		.dout(new_net_8675)
	);

	bfr new_net_8676_bfr_after (
		.din(new_net_8675),
		.dout(new_net_8676)
	);

	bfr new_net_8677_bfr_after (
		.din(new_net_8676),
		.dout(new_net_8677)
	);

	bfr new_net_8678_bfr_after (
		.din(new_net_8677),
		.dout(new_net_8678)
	);

	bfr new_net_8679_bfr_after (
		.din(new_net_8678),
		.dout(new_net_8679)
	);

	bfr new_net_8680_bfr_after (
		.din(new_net_8679),
		.dout(new_net_8680)
	);

	bfr new_net_8681_bfr_after (
		.din(new_net_8680),
		.dout(new_net_8681)
	);

	bfr new_net_8682_bfr_after (
		.din(new_net_8681),
		.dout(new_net_8682)
	);

	bfr new_net_8683_bfr_after (
		.din(new_net_8682),
		.dout(new_net_8683)
	);

	bfr new_net_8684_bfr_after (
		.din(new_net_8683),
		.dout(new_net_8684)
	);

	bfr new_net_8685_bfr_after (
		.din(new_net_8684),
		.dout(new_net_8685)
	);

	bfr new_net_8686_bfr_after (
		.din(new_net_8685),
		.dout(new_net_8686)
	);

	bfr new_net_8687_bfr_after (
		.din(new_net_8686),
		.dout(new_net_8687)
	);

	bfr new_net_8688_bfr_after (
		.din(new_net_8687),
		.dout(new_net_8688)
	);

	spl2 _1282__v_fanout (
		.a(new_net_8688),
		.b(new_net_842),
		.c(new_net_843)
	);

	bfr new_net_8689_bfr_after (
		.din(_1567_),
		.dout(new_net_8689)
	);

	bfr new_net_8690_bfr_after (
		.din(new_net_8689),
		.dout(new_net_8690)
	);

	bfr new_net_8691_bfr_after (
		.din(new_net_8690),
		.dout(new_net_8691)
	);

	bfr new_net_8692_bfr_after (
		.din(new_net_8691),
		.dout(new_net_8692)
	);

	bfr new_net_8693_bfr_after (
		.din(new_net_8692),
		.dout(new_net_8693)
	);

	bfr new_net_8694_bfr_after (
		.din(new_net_8693),
		.dout(new_net_8694)
	);

	bfr new_net_8695_bfr_after (
		.din(new_net_8694),
		.dout(new_net_8695)
	);

	bfr new_net_8696_bfr_after (
		.din(new_net_8695),
		.dout(new_net_8696)
	);

	bfr new_net_8697_bfr_after (
		.din(new_net_8696),
		.dout(new_net_8697)
	);

	bfr new_net_8698_bfr_after (
		.din(new_net_8697),
		.dout(new_net_8698)
	);

	bfr new_net_8699_bfr_after (
		.din(new_net_8698),
		.dout(new_net_8699)
	);

	bfr new_net_8700_bfr_after (
		.din(new_net_8699),
		.dout(new_net_8700)
	);

	bfr new_net_8701_bfr_after (
		.din(new_net_8700),
		.dout(new_net_8701)
	);

	bfr new_net_8702_bfr_after (
		.din(new_net_8701),
		.dout(new_net_8702)
	);

	bfr new_net_8703_bfr_after (
		.din(new_net_8702),
		.dout(new_net_8703)
	);

	bfr new_net_8704_bfr_after (
		.din(new_net_8703),
		.dout(new_net_8704)
	);

	bfr new_net_8705_bfr_after (
		.din(new_net_8704),
		.dout(new_net_8705)
	);

	bfr new_net_8706_bfr_after (
		.din(new_net_8705),
		.dout(new_net_8706)
	);

	bfr new_net_8707_bfr_after (
		.din(new_net_8706),
		.dout(new_net_8707)
	);

	bfr new_net_8708_bfr_after (
		.din(new_net_8707),
		.dout(new_net_8708)
	);

	bfr new_net_8709_bfr_after (
		.din(new_net_8708),
		.dout(new_net_8709)
	);

	bfr new_net_8710_bfr_after (
		.din(new_net_8709),
		.dout(new_net_8710)
	);

	bfr new_net_8711_bfr_after (
		.din(new_net_8710),
		.dout(new_net_8711)
	);

	bfr new_net_8712_bfr_after (
		.din(new_net_8711),
		.dout(new_net_8712)
	);

	bfr new_net_8713_bfr_after (
		.din(new_net_8712),
		.dout(new_net_8713)
	);

	bfr new_net_8714_bfr_after (
		.din(new_net_8713),
		.dout(new_net_8714)
	);

	bfr new_net_8715_bfr_after (
		.din(new_net_8714),
		.dout(new_net_8715)
	);

	bfr new_net_8716_bfr_after (
		.din(new_net_8715),
		.dout(new_net_8716)
	);

	bfr new_net_8717_bfr_after (
		.din(new_net_8716),
		.dout(new_net_8717)
	);

	bfr new_net_8718_bfr_after (
		.din(new_net_8717),
		.dout(new_net_8718)
	);

	bfr new_net_8719_bfr_after (
		.din(new_net_8718),
		.dout(new_net_8719)
	);

	bfr new_net_8720_bfr_after (
		.din(new_net_8719),
		.dout(new_net_8720)
	);

	bfr new_net_8721_bfr_after (
		.din(new_net_8720),
		.dout(new_net_8721)
	);

	bfr new_net_8722_bfr_after (
		.din(new_net_8721),
		.dout(new_net_8722)
	);

	bfr new_net_8723_bfr_after (
		.din(new_net_8722),
		.dout(new_net_8723)
	);

	bfr new_net_8724_bfr_after (
		.din(new_net_8723),
		.dout(new_net_8724)
	);

	bfr new_net_8725_bfr_after (
		.din(new_net_8724),
		.dout(new_net_8725)
	);

	bfr new_net_8726_bfr_after (
		.din(new_net_8725),
		.dout(new_net_8726)
	);

	bfr new_net_8727_bfr_after (
		.din(new_net_8726),
		.dout(new_net_8727)
	);

	bfr new_net_8728_bfr_after (
		.din(new_net_8727),
		.dout(new_net_8728)
	);

	bfr new_net_8729_bfr_after (
		.din(new_net_8728),
		.dout(new_net_8729)
	);

	bfr new_net_8730_bfr_after (
		.din(new_net_8729),
		.dout(new_net_8730)
	);

	bfr new_net_8731_bfr_after (
		.din(new_net_8730),
		.dout(new_net_8731)
	);

	bfr new_net_8732_bfr_after (
		.din(new_net_8731),
		.dout(new_net_8732)
	);

	bfr new_net_8733_bfr_after (
		.din(new_net_8732),
		.dout(new_net_8733)
	);

	bfr new_net_8734_bfr_after (
		.din(new_net_8733),
		.dout(new_net_8734)
	);

	bfr new_net_8735_bfr_after (
		.din(new_net_8734),
		.dout(new_net_8735)
	);

	bfr new_net_8736_bfr_after (
		.din(new_net_8735),
		.dout(new_net_8736)
	);

	bfr new_net_8737_bfr_after (
		.din(new_net_8736),
		.dout(new_net_8737)
	);

	bfr new_net_8738_bfr_after (
		.din(new_net_8737),
		.dout(new_net_8738)
	);

	bfr new_net_8739_bfr_after (
		.din(new_net_8738),
		.dout(new_net_8739)
	);

	bfr new_net_8740_bfr_after (
		.din(new_net_8739),
		.dout(new_net_8740)
	);

	bfr new_net_8741_bfr_after (
		.din(new_net_8740),
		.dout(new_net_8741)
	);

	bfr new_net_8742_bfr_after (
		.din(new_net_8741),
		.dout(new_net_8742)
	);

	bfr new_net_8743_bfr_after (
		.din(new_net_8742),
		.dout(new_net_8743)
	);

	bfr new_net_8744_bfr_after (
		.din(new_net_8743),
		.dout(new_net_8744)
	);

	bfr new_net_8745_bfr_after (
		.din(new_net_8744),
		.dout(new_net_8745)
	);

	bfr new_net_8746_bfr_after (
		.din(new_net_8745),
		.dout(new_net_8746)
	);

	bfr new_net_8747_bfr_after (
		.din(new_net_8746),
		.dout(new_net_8747)
	);

	bfr new_net_8748_bfr_after (
		.din(new_net_8747),
		.dout(new_net_8748)
	);

	bfr new_net_8749_bfr_after (
		.din(new_net_8748),
		.dout(new_net_8749)
	);

	bfr new_net_8750_bfr_after (
		.din(new_net_8749),
		.dout(new_net_8750)
	);

	bfr new_net_8751_bfr_after (
		.din(new_net_8750),
		.dout(new_net_8751)
	);

	bfr new_net_8752_bfr_after (
		.din(new_net_8751),
		.dout(new_net_8752)
	);

	bfr new_net_8753_bfr_after (
		.din(new_net_8752),
		.dout(new_net_8753)
	);

	bfr new_net_8754_bfr_after (
		.din(new_net_8753),
		.dout(new_net_8754)
	);

	bfr new_net_8755_bfr_after (
		.din(new_net_8754),
		.dout(new_net_8755)
	);

	bfr new_net_8756_bfr_after (
		.din(new_net_8755),
		.dout(new_net_8756)
	);

	bfr new_net_8757_bfr_after (
		.din(new_net_8756),
		.dout(new_net_8757)
	);

	bfr new_net_8758_bfr_after (
		.din(new_net_8757),
		.dout(new_net_8758)
	);

	bfr new_net_8759_bfr_after (
		.din(new_net_8758),
		.dout(new_net_8759)
	);

	bfr new_net_8760_bfr_after (
		.din(new_net_8759),
		.dout(new_net_8760)
	);

	bfr new_net_8761_bfr_after (
		.din(new_net_8760),
		.dout(new_net_8761)
	);

	bfr new_net_8762_bfr_after (
		.din(new_net_8761),
		.dout(new_net_8762)
	);

	bfr new_net_8763_bfr_after (
		.din(new_net_8762),
		.dout(new_net_8763)
	);

	bfr new_net_8764_bfr_after (
		.din(new_net_8763),
		.dout(new_net_8764)
	);

	bfr new_net_8765_bfr_after (
		.din(new_net_8764),
		.dout(new_net_8765)
	);

	bfr new_net_8766_bfr_after (
		.din(new_net_8765),
		.dout(new_net_8766)
	);

	bfr new_net_8767_bfr_after (
		.din(new_net_8766),
		.dout(new_net_8767)
	);

	bfr new_net_8768_bfr_after (
		.din(new_net_8767),
		.dout(new_net_8768)
	);

	spl2 _1567__v_fanout (
		.a(new_net_8768),
		.b(new_net_3250),
		.c(new_net_3251)
	);

	bfr new_net_8769_bfr_after (
		.din(_0631_),
		.dout(new_net_8769)
	);

	bfr new_net_8770_bfr_after (
		.din(new_net_8769),
		.dout(new_net_8770)
	);

	bfr new_net_8771_bfr_after (
		.din(new_net_8770),
		.dout(new_net_8771)
	);

	bfr new_net_8772_bfr_after (
		.din(new_net_8771),
		.dout(new_net_8772)
	);

	bfr new_net_8773_bfr_after (
		.din(new_net_8772),
		.dout(new_net_8773)
	);

	bfr new_net_8774_bfr_after (
		.din(new_net_8773),
		.dout(new_net_8774)
	);

	bfr new_net_8775_bfr_after (
		.din(new_net_8774),
		.dout(new_net_8775)
	);

	bfr new_net_8776_bfr_after (
		.din(new_net_8775),
		.dout(new_net_8776)
	);

	bfr new_net_8777_bfr_after (
		.din(new_net_8776),
		.dout(new_net_8777)
	);

	bfr new_net_8778_bfr_after (
		.din(new_net_8777),
		.dout(new_net_8778)
	);

	bfr new_net_8779_bfr_after (
		.din(new_net_8778),
		.dout(new_net_8779)
	);

	bfr new_net_8780_bfr_after (
		.din(new_net_8779),
		.dout(new_net_8780)
	);

	bfr new_net_8781_bfr_after (
		.din(new_net_8780),
		.dout(new_net_8781)
	);

	bfr new_net_8782_bfr_after (
		.din(new_net_8781),
		.dout(new_net_8782)
	);

	bfr new_net_8783_bfr_after (
		.din(new_net_8782),
		.dout(new_net_8783)
	);

	bfr new_net_8784_bfr_after (
		.din(new_net_8783),
		.dout(new_net_8784)
	);

	bfr new_net_8785_bfr_after (
		.din(new_net_8784),
		.dout(new_net_8785)
	);

	bfr new_net_8786_bfr_after (
		.din(new_net_8785),
		.dout(new_net_8786)
	);

	bfr new_net_8787_bfr_after (
		.din(new_net_8786),
		.dout(new_net_8787)
	);

	bfr new_net_8788_bfr_after (
		.din(new_net_8787),
		.dout(new_net_8788)
	);

	bfr new_net_8789_bfr_after (
		.din(new_net_8788),
		.dout(new_net_8789)
	);

	bfr new_net_8790_bfr_after (
		.din(new_net_8789),
		.dout(new_net_8790)
	);

	bfr new_net_8791_bfr_after (
		.din(new_net_8790),
		.dout(new_net_8791)
	);

	bfr new_net_8792_bfr_after (
		.din(new_net_8791),
		.dout(new_net_8792)
	);

	bfr new_net_8793_bfr_after (
		.din(new_net_8792),
		.dout(new_net_8793)
	);

	bfr new_net_8794_bfr_after (
		.din(new_net_8793),
		.dout(new_net_8794)
	);

	bfr new_net_8795_bfr_after (
		.din(new_net_8794),
		.dout(new_net_8795)
	);

	bfr new_net_8796_bfr_after (
		.din(new_net_8795),
		.dout(new_net_8796)
	);

	bfr new_net_8797_bfr_after (
		.din(new_net_8796),
		.dout(new_net_8797)
	);

	bfr new_net_8798_bfr_after (
		.din(new_net_8797),
		.dout(new_net_8798)
	);

	bfr new_net_8799_bfr_after (
		.din(new_net_8798),
		.dout(new_net_8799)
	);

	bfr new_net_8800_bfr_after (
		.din(new_net_8799),
		.dout(new_net_8800)
	);

	bfr new_net_8801_bfr_after (
		.din(new_net_8800),
		.dout(new_net_8801)
	);

	bfr new_net_8802_bfr_after (
		.din(new_net_8801),
		.dout(new_net_8802)
	);

	bfr new_net_8803_bfr_after (
		.din(new_net_8802),
		.dout(new_net_8803)
	);

	bfr new_net_8804_bfr_after (
		.din(new_net_8803),
		.dout(new_net_8804)
	);

	bfr new_net_8805_bfr_after (
		.din(new_net_8804),
		.dout(new_net_8805)
	);

	bfr new_net_8806_bfr_after (
		.din(new_net_8805),
		.dout(new_net_8806)
	);

	bfr new_net_8807_bfr_after (
		.din(new_net_8806),
		.dout(new_net_8807)
	);

	bfr new_net_8808_bfr_after (
		.din(new_net_8807),
		.dout(new_net_8808)
	);

	bfr new_net_8809_bfr_after (
		.din(new_net_8808),
		.dout(new_net_8809)
	);

	bfr new_net_8810_bfr_after (
		.din(new_net_8809),
		.dout(new_net_8810)
	);

	bfr new_net_8811_bfr_after (
		.din(new_net_8810),
		.dout(new_net_8811)
	);

	bfr new_net_8812_bfr_after (
		.din(new_net_8811),
		.dout(new_net_8812)
	);

	bfr new_net_8813_bfr_after (
		.din(new_net_8812),
		.dout(new_net_8813)
	);

	bfr new_net_8814_bfr_after (
		.din(new_net_8813),
		.dout(new_net_8814)
	);

	bfr new_net_8815_bfr_after (
		.din(new_net_8814),
		.dout(new_net_8815)
	);

	bfr new_net_8816_bfr_after (
		.din(new_net_8815),
		.dout(new_net_8816)
	);

	bfr new_net_8817_bfr_after (
		.din(new_net_8816),
		.dout(new_net_8817)
	);

	bfr new_net_8818_bfr_after (
		.din(new_net_8817),
		.dout(new_net_8818)
	);

	spl2 _0631__v_fanout (
		.a(new_net_8818),
		.b(new_net_1074),
		.c(new_net_1075)
	);

	bfr new_net_8819_bfr_after (
		.din(_1142_),
		.dout(new_net_8819)
	);

	bfr new_net_8820_bfr_after (
		.din(new_net_8819),
		.dout(new_net_8820)
	);

	bfr new_net_8821_bfr_after (
		.din(new_net_8820),
		.dout(new_net_8821)
	);

	bfr new_net_8822_bfr_after (
		.din(new_net_8821),
		.dout(new_net_8822)
	);

	bfr new_net_8823_bfr_after (
		.din(new_net_8822),
		.dout(new_net_8823)
	);

	bfr new_net_8824_bfr_after (
		.din(new_net_8823),
		.dout(new_net_8824)
	);

	bfr new_net_8825_bfr_after (
		.din(new_net_8824),
		.dout(new_net_8825)
	);

	bfr new_net_8826_bfr_after (
		.din(new_net_8825),
		.dout(new_net_8826)
	);

	spl2 _1142__v_fanout (
		.a(new_net_8826),
		.b(new_net_2166),
		.c(new_net_2167)
	);

	bfr new_net_8827_bfr_after (
		.din(_0629_),
		.dout(new_net_8827)
	);

	bfr new_net_8828_bfr_after (
		.din(new_net_8827),
		.dout(new_net_8828)
	);

	bfr new_net_8829_bfr_after (
		.din(new_net_8828),
		.dout(new_net_8829)
	);

	bfr new_net_8830_bfr_after (
		.din(new_net_8829),
		.dout(new_net_8830)
	);

	bfr new_net_8831_bfr_after (
		.din(new_net_8830),
		.dout(new_net_8831)
	);

	bfr new_net_8832_bfr_after (
		.din(new_net_8831),
		.dout(new_net_8832)
	);

	bfr new_net_8833_bfr_after (
		.din(new_net_8832),
		.dout(new_net_8833)
	);

	bfr new_net_8834_bfr_after (
		.din(new_net_8833),
		.dout(new_net_8834)
	);

	bfr new_net_8835_bfr_after (
		.din(new_net_8834),
		.dout(new_net_8835)
	);

	bfr new_net_8836_bfr_after (
		.din(new_net_8835),
		.dout(new_net_8836)
	);

	bfr new_net_8837_bfr_after (
		.din(new_net_8836),
		.dout(new_net_8837)
	);

	bfr new_net_8838_bfr_after (
		.din(new_net_8837),
		.dout(new_net_8838)
	);

	bfr new_net_8839_bfr_after (
		.din(new_net_8838),
		.dout(new_net_8839)
	);

	bfr new_net_8840_bfr_after (
		.din(new_net_8839),
		.dout(new_net_8840)
	);

	bfr new_net_8841_bfr_after (
		.din(new_net_8840),
		.dout(new_net_8841)
	);

	bfr new_net_8842_bfr_after (
		.din(new_net_8841),
		.dout(new_net_8842)
	);

	bfr new_net_8843_bfr_after (
		.din(new_net_8842),
		.dout(new_net_8843)
	);

	bfr new_net_8844_bfr_after (
		.din(new_net_8843),
		.dout(new_net_8844)
	);

	bfr new_net_8845_bfr_after (
		.din(new_net_8844),
		.dout(new_net_8845)
	);

	bfr new_net_8846_bfr_after (
		.din(new_net_8845),
		.dout(new_net_8846)
	);

	bfr new_net_8847_bfr_after (
		.din(new_net_8846),
		.dout(new_net_8847)
	);

	bfr new_net_8848_bfr_after (
		.din(new_net_8847),
		.dout(new_net_8848)
	);

	bfr new_net_8849_bfr_after (
		.din(new_net_8848),
		.dout(new_net_8849)
	);

	bfr new_net_8850_bfr_after (
		.din(new_net_8849),
		.dout(new_net_8850)
	);

	bfr new_net_8851_bfr_after (
		.din(new_net_8850),
		.dout(new_net_8851)
	);

	bfr new_net_8852_bfr_after (
		.din(new_net_8851),
		.dout(new_net_8852)
	);

	bfr new_net_8853_bfr_after (
		.din(new_net_8852),
		.dout(new_net_8853)
	);

	bfr new_net_8854_bfr_after (
		.din(new_net_8853),
		.dout(new_net_8854)
	);

	bfr new_net_8855_bfr_after (
		.din(new_net_8854),
		.dout(new_net_8855)
	);

	bfr new_net_8856_bfr_after (
		.din(new_net_8855),
		.dout(new_net_8856)
	);

	bfr new_net_8857_bfr_after (
		.din(new_net_8856),
		.dout(new_net_8857)
	);

	bfr new_net_8858_bfr_after (
		.din(new_net_8857),
		.dout(new_net_8858)
	);

	bfr new_net_8859_bfr_after (
		.din(new_net_8858),
		.dout(new_net_8859)
	);

	bfr new_net_8860_bfr_after (
		.din(new_net_8859),
		.dout(new_net_8860)
	);

	bfr new_net_8861_bfr_after (
		.din(new_net_8860),
		.dout(new_net_8861)
	);

	bfr new_net_8862_bfr_after (
		.din(new_net_8861),
		.dout(new_net_8862)
	);

	bfr new_net_8863_bfr_after (
		.din(new_net_8862),
		.dout(new_net_8863)
	);

	bfr new_net_8864_bfr_after (
		.din(new_net_8863),
		.dout(new_net_8864)
	);

	bfr new_net_8865_bfr_after (
		.din(new_net_8864),
		.dout(new_net_8865)
	);

	bfr new_net_8866_bfr_after (
		.din(new_net_8865),
		.dout(new_net_8866)
	);

	bfr new_net_8867_bfr_after (
		.din(new_net_8866),
		.dout(new_net_8867)
	);

	bfr new_net_8868_bfr_after (
		.din(new_net_8867),
		.dout(new_net_8868)
	);

	bfr new_net_8869_bfr_after (
		.din(new_net_8868),
		.dout(new_net_8869)
	);

	bfr new_net_8870_bfr_after (
		.din(new_net_8869),
		.dout(new_net_8870)
	);

	bfr new_net_8871_bfr_after (
		.din(new_net_8870),
		.dout(new_net_8871)
	);

	bfr new_net_8872_bfr_after (
		.din(new_net_8871),
		.dout(new_net_8872)
	);

	bfr new_net_8873_bfr_after (
		.din(new_net_8872),
		.dout(new_net_8873)
	);

	bfr new_net_8874_bfr_after (
		.din(new_net_8873),
		.dout(new_net_8874)
	);

	bfr new_net_8875_bfr_after (
		.din(new_net_8874),
		.dout(new_net_8875)
	);

	bfr new_net_8876_bfr_after (
		.din(new_net_8875),
		.dout(new_net_8876)
	);

	bfr new_net_8877_bfr_after (
		.din(new_net_8876),
		.dout(new_net_8877)
	);

	bfr new_net_8878_bfr_after (
		.din(new_net_8877),
		.dout(new_net_8878)
	);

	bfr new_net_8879_bfr_after (
		.din(new_net_8878),
		.dout(new_net_8879)
	);

	bfr new_net_8880_bfr_after (
		.din(new_net_8879),
		.dout(new_net_8880)
	);

	bfr new_net_8881_bfr_after (
		.din(new_net_8880),
		.dout(new_net_8881)
	);

	bfr new_net_8882_bfr_after (
		.din(new_net_8881),
		.dout(new_net_8882)
	);

	bfr new_net_8883_bfr_after (
		.din(new_net_8882),
		.dout(new_net_8883)
	);

	bfr new_net_8884_bfr_after (
		.din(new_net_8883),
		.dout(new_net_8884)
	);

	bfr new_net_8885_bfr_after (
		.din(new_net_8884),
		.dout(new_net_8885)
	);

	bfr new_net_8886_bfr_after (
		.din(new_net_8885),
		.dout(new_net_8886)
	);

	bfr new_net_8887_bfr_after (
		.din(new_net_8886),
		.dout(new_net_8887)
	);

	bfr new_net_8888_bfr_after (
		.din(new_net_8887),
		.dout(new_net_8888)
	);

	spl2 _0629__v_fanout (
		.a(new_net_8888),
		.b(new_net_1360),
		.c(new_net_1361)
	);

	spl2 _1513__v_fanout (
		.a(_1513_),
		.b(new_net_2573),
		.c(new_net_2574)
	);

	bfr new_net_8889_bfr_after (
		.din(_1458_),
		.dout(new_net_8889)
	);

	bfr new_net_8890_bfr_after (
		.din(new_net_8889),
		.dout(new_net_8890)
	);

	bfr new_net_8891_bfr_after (
		.din(new_net_8890),
		.dout(new_net_8891)
	);

	bfr new_net_8892_bfr_after (
		.din(new_net_8891),
		.dout(new_net_8892)
	);

	bfr new_net_8893_bfr_after (
		.din(new_net_8892),
		.dout(new_net_8893)
	);

	bfr new_net_8894_bfr_after (
		.din(new_net_8893),
		.dout(new_net_8894)
	);

	bfr new_net_8895_bfr_after (
		.din(new_net_8894),
		.dout(new_net_8895)
	);

	bfr new_net_8896_bfr_after (
		.din(new_net_8895),
		.dout(new_net_8896)
	);

	bfr new_net_8897_bfr_after (
		.din(new_net_8896),
		.dout(new_net_8897)
	);

	bfr new_net_8898_bfr_after (
		.din(new_net_8897),
		.dout(new_net_8898)
	);

	bfr new_net_8899_bfr_after (
		.din(new_net_8898),
		.dout(new_net_8899)
	);

	bfr new_net_8900_bfr_after (
		.din(new_net_8899),
		.dout(new_net_8900)
	);

	bfr new_net_8901_bfr_after (
		.din(new_net_8900),
		.dout(new_net_8901)
	);

	bfr new_net_8902_bfr_after (
		.din(new_net_8901),
		.dout(new_net_8902)
	);

	bfr new_net_8903_bfr_after (
		.din(new_net_8902),
		.dout(new_net_8903)
	);

	bfr new_net_8904_bfr_after (
		.din(new_net_8903),
		.dout(new_net_8904)
	);

	spl2 _1458__v_fanout (
		.a(new_net_8904),
		.b(new_net_620),
		.c(new_net_621)
	);

	bfr new_net_8905_bfr_after (
		.din(_0701_),
		.dout(new_net_8905)
	);

	bfr new_net_8906_bfr_after (
		.din(new_net_8905),
		.dout(new_net_8906)
	);

	bfr new_net_8907_bfr_after (
		.din(new_net_8906),
		.dout(new_net_8907)
	);

	bfr new_net_8908_bfr_after (
		.din(new_net_8907),
		.dout(new_net_8908)
	);

	bfr new_net_8909_bfr_after (
		.din(new_net_8908),
		.dout(new_net_8909)
	);

	bfr new_net_8910_bfr_after (
		.din(new_net_8909),
		.dout(new_net_8910)
	);

	bfr new_net_8911_bfr_after (
		.din(new_net_8910),
		.dout(new_net_8911)
	);

	bfr new_net_8912_bfr_after (
		.din(new_net_8911),
		.dout(new_net_8912)
	);

	bfr new_net_8913_bfr_after (
		.din(new_net_8912),
		.dout(new_net_8913)
	);

	bfr new_net_8914_bfr_after (
		.din(new_net_8913),
		.dout(new_net_8914)
	);

	bfr new_net_8915_bfr_after (
		.din(new_net_8914),
		.dout(new_net_8915)
	);

	bfr new_net_8916_bfr_after (
		.din(new_net_8915),
		.dout(new_net_8916)
	);

	bfr new_net_8917_bfr_after (
		.din(new_net_8916),
		.dout(new_net_8917)
	);

	bfr new_net_8918_bfr_after (
		.din(new_net_8917),
		.dout(new_net_8918)
	);

	bfr new_net_8919_bfr_after (
		.din(new_net_8918),
		.dout(new_net_8919)
	);

	bfr new_net_8920_bfr_after (
		.din(new_net_8919),
		.dout(new_net_8920)
	);

	bfr new_net_8921_bfr_after (
		.din(new_net_8920),
		.dout(new_net_8921)
	);

	bfr new_net_8922_bfr_after (
		.din(new_net_8921),
		.dout(new_net_8922)
	);

	bfr new_net_8923_bfr_after (
		.din(new_net_8922),
		.dout(new_net_8923)
	);

	bfr new_net_8924_bfr_after (
		.din(new_net_8923),
		.dout(new_net_8924)
	);

	bfr new_net_8925_bfr_after (
		.din(new_net_8924),
		.dout(new_net_8925)
	);

	bfr new_net_8926_bfr_after (
		.din(new_net_8925),
		.dout(new_net_8926)
	);

	bfr new_net_8927_bfr_after (
		.din(new_net_8926),
		.dout(new_net_8927)
	);

	bfr new_net_8928_bfr_after (
		.din(new_net_8927),
		.dout(new_net_8928)
	);

	bfr new_net_8929_bfr_after (
		.din(new_net_8928),
		.dout(new_net_8929)
	);

	bfr new_net_8930_bfr_after (
		.din(new_net_8929),
		.dout(new_net_8930)
	);

	bfr new_net_8931_bfr_after (
		.din(new_net_8930),
		.dout(new_net_8931)
	);

	bfr new_net_8932_bfr_after (
		.din(new_net_8931),
		.dout(new_net_8932)
	);

	bfr new_net_8933_bfr_after (
		.din(new_net_8932),
		.dout(new_net_8933)
	);

	bfr new_net_8934_bfr_after (
		.din(new_net_8933),
		.dout(new_net_8934)
	);

	bfr new_net_8935_bfr_after (
		.din(new_net_8934),
		.dout(new_net_8935)
	);

	bfr new_net_8936_bfr_after (
		.din(new_net_8935),
		.dout(new_net_8936)
	);

	bfr new_net_8937_bfr_after (
		.din(new_net_8936),
		.dout(new_net_8937)
	);

	bfr new_net_8938_bfr_after (
		.din(new_net_8937),
		.dout(new_net_8938)
	);

	bfr new_net_8939_bfr_after (
		.din(new_net_8938),
		.dout(new_net_8939)
	);

	bfr new_net_8940_bfr_after (
		.din(new_net_8939),
		.dout(new_net_8940)
	);

	bfr new_net_8941_bfr_after (
		.din(new_net_8940),
		.dout(new_net_8941)
	);

	bfr new_net_8942_bfr_after (
		.din(new_net_8941),
		.dout(new_net_8942)
	);

	bfr new_net_8943_bfr_after (
		.din(new_net_8942),
		.dout(new_net_8943)
	);

	bfr new_net_8944_bfr_after (
		.din(new_net_8943),
		.dout(new_net_8944)
	);

	bfr new_net_8945_bfr_after (
		.din(new_net_8944),
		.dout(new_net_8945)
	);

	bfr new_net_8946_bfr_after (
		.din(new_net_8945),
		.dout(new_net_8946)
	);

	bfr new_net_8947_bfr_after (
		.din(new_net_8946),
		.dout(new_net_8947)
	);

	bfr new_net_8948_bfr_after (
		.din(new_net_8947),
		.dout(new_net_8948)
	);

	bfr new_net_8949_bfr_after (
		.din(new_net_8948),
		.dout(new_net_8949)
	);

	bfr new_net_8950_bfr_after (
		.din(new_net_8949),
		.dout(new_net_8950)
	);

	bfr new_net_8951_bfr_after (
		.din(new_net_8950),
		.dout(new_net_8951)
	);

	bfr new_net_8952_bfr_after (
		.din(new_net_8951),
		.dout(new_net_8952)
	);

	bfr new_net_8953_bfr_after (
		.din(new_net_8952),
		.dout(new_net_8953)
	);

	bfr new_net_8954_bfr_after (
		.din(new_net_8953),
		.dout(new_net_8954)
	);

	bfr new_net_8955_bfr_after (
		.din(new_net_8954),
		.dout(new_net_8955)
	);

	bfr new_net_8956_bfr_after (
		.din(new_net_8955),
		.dout(new_net_8956)
	);

	bfr new_net_8957_bfr_after (
		.din(new_net_8956),
		.dout(new_net_8957)
	);

	bfr new_net_8958_bfr_after (
		.din(new_net_8957),
		.dout(new_net_8958)
	);

	bfr new_net_8959_bfr_after (
		.din(new_net_8958),
		.dout(new_net_8959)
	);

	bfr new_net_8960_bfr_after (
		.din(new_net_8959),
		.dout(new_net_8960)
	);

	bfr new_net_8961_bfr_after (
		.din(new_net_8960),
		.dout(new_net_8961)
	);

	bfr new_net_8962_bfr_after (
		.din(new_net_8961),
		.dout(new_net_8962)
	);

	bfr new_net_8963_bfr_after (
		.din(new_net_8962),
		.dout(new_net_8963)
	);

	bfr new_net_8964_bfr_after (
		.din(new_net_8963),
		.dout(new_net_8964)
	);

	bfr new_net_8965_bfr_after (
		.din(new_net_8964),
		.dout(new_net_8965)
	);

	bfr new_net_8966_bfr_after (
		.din(new_net_8965),
		.dout(new_net_8966)
	);

	bfr new_net_8967_bfr_after (
		.din(new_net_8966),
		.dout(new_net_8967)
	);

	bfr new_net_8968_bfr_after (
		.din(new_net_8967),
		.dout(new_net_8968)
	);

	bfr new_net_8969_bfr_after (
		.din(new_net_8968),
		.dout(new_net_8969)
	);

	bfr new_net_8970_bfr_after (
		.din(new_net_8969),
		.dout(new_net_8970)
	);

	bfr new_net_8971_bfr_after (
		.din(new_net_8970),
		.dout(new_net_8971)
	);

	bfr new_net_8972_bfr_after (
		.din(new_net_8971),
		.dout(new_net_8972)
	);

	bfr new_net_8973_bfr_after (
		.din(new_net_8972),
		.dout(new_net_8973)
	);

	bfr new_net_8974_bfr_after (
		.din(new_net_8973),
		.dout(new_net_8974)
	);

	bfr new_net_8975_bfr_after (
		.din(new_net_8974),
		.dout(new_net_8975)
	);

	bfr new_net_8976_bfr_after (
		.din(new_net_8975),
		.dout(new_net_8976)
	);

	bfr new_net_8977_bfr_after (
		.din(new_net_8976),
		.dout(new_net_8977)
	);

	bfr new_net_8978_bfr_after (
		.din(new_net_8977),
		.dout(new_net_8978)
	);

	bfr new_net_8979_bfr_after (
		.din(new_net_8978),
		.dout(new_net_8979)
	);

	bfr new_net_8980_bfr_after (
		.din(new_net_8979),
		.dout(new_net_8980)
	);

	bfr new_net_8981_bfr_after (
		.din(new_net_8980),
		.dout(new_net_8981)
	);

	bfr new_net_8982_bfr_after (
		.din(new_net_8981),
		.dout(new_net_8982)
	);

	bfr new_net_8983_bfr_after (
		.din(new_net_8982),
		.dout(new_net_8983)
	);

	bfr new_net_8984_bfr_after (
		.din(new_net_8983),
		.dout(new_net_8984)
	);

	bfr new_net_8985_bfr_after (
		.din(new_net_8984),
		.dout(new_net_8985)
	);

	bfr new_net_8986_bfr_after (
		.din(new_net_8985),
		.dout(new_net_8986)
	);

	bfr new_net_8987_bfr_after (
		.din(new_net_8986),
		.dout(new_net_8987)
	);

	bfr new_net_8988_bfr_after (
		.din(new_net_8987),
		.dout(new_net_8988)
	);

	bfr new_net_8989_bfr_after (
		.din(new_net_8988),
		.dout(new_net_8989)
	);

	bfr new_net_8990_bfr_after (
		.din(new_net_8989),
		.dout(new_net_8990)
	);

	bfr new_net_8991_bfr_after (
		.din(new_net_8990),
		.dout(new_net_8991)
	);

	bfr new_net_8992_bfr_after (
		.din(new_net_8991),
		.dout(new_net_8992)
	);

	bfr new_net_8993_bfr_after (
		.din(new_net_8992),
		.dout(new_net_8993)
	);

	bfr new_net_8994_bfr_after (
		.din(new_net_8993),
		.dout(new_net_8994)
	);

	bfr new_net_8995_bfr_after (
		.din(new_net_8994),
		.dout(new_net_8995)
	);

	bfr new_net_8996_bfr_after (
		.din(new_net_8995),
		.dout(new_net_8996)
	);

	bfr new_net_8997_bfr_after (
		.din(new_net_8996),
		.dout(new_net_8997)
	);

	bfr new_net_8998_bfr_after (
		.din(new_net_8997),
		.dout(new_net_8998)
	);

	bfr new_net_8999_bfr_after (
		.din(new_net_8998),
		.dout(new_net_8999)
	);

	bfr new_net_9000_bfr_after (
		.din(new_net_8999),
		.dout(new_net_9000)
	);

	spl2 _0701__v_fanout (
		.a(new_net_9000),
		.b(new_net_2513),
		.c(new_net_2514)
	);

	spl2 _1665__v_fanout (
		.a(_1665_),
		.b(new_net_2442),
		.c(new_net_2443)
	);

	bfr new_net_9001_bfr_after (
		.din(_1288_),
		.dout(new_net_9001)
	);

	bfr new_net_9002_bfr_after (
		.din(new_net_9001),
		.dout(new_net_9002)
	);

	bfr new_net_9003_bfr_after (
		.din(new_net_9002),
		.dout(new_net_9003)
	);

	bfr new_net_9004_bfr_after (
		.din(new_net_9003),
		.dout(new_net_9004)
	);

	bfr new_net_9005_bfr_after (
		.din(new_net_9004),
		.dout(new_net_9005)
	);

	bfr new_net_9006_bfr_after (
		.din(new_net_9005),
		.dout(new_net_9006)
	);

	bfr new_net_9007_bfr_after (
		.din(new_net_9006),
		.dout(new_net_9007)
	);

	bfr new_net_9008_bfr_after (
		.din(new_net_9007),
		.dout(new_net_9008)
	);

	bfr new_net_9009_bfr_after (
		.din(new_net_9008),
		.dout(new_net_9009)
	);

	bfr new_net_9010_bfr_after (
		.din(new_net_9009),
		.dout(new_net_9010)
	);

	bfr new_net_9011_bfr_after (
		.din(new_net_9010),
		.dout(new_net_9011)
	);

	bfr new_net_9012_bfr_after (
		.din(new_net_9011),
		.dout(new_net_9012)
	);

	bfr new_net_9013_bfr_after (
		.din(new_net_9012),
		.dout(new_net_9013)
	);

	bfr new_net_9014_bfr_after (
		.din(new_net_9013),
		.dout(new_net_9014)
	);

	bfr new_net_9015_bfr_after (
		.din(new_net_9014),
		.dout(new_net_9015)
	);

	bfr new_net_9016_bfr_after (
		.din(new_net_9015),
		.dout(new_net_9016)
	);

	bfr new_net_9017_bfr_after (
		.din(new_net_9016),
		.dout(new_net_9017)
	);

	bfr new_net_9018_bfr_after (
		.din(new_net_9017),
		.dout(new_net_9018)
	);

	bfr new_net_9019_bfr_after (
		.din(new_net_9018),
		.dout(new_net_9019)
	);

	bfr new_net_9020_bfr_after (
		.din(new_net_9019),
		.dout(new_net_9020)
	);

	bfr new_net_9021_bfr_after (
		.din(new_net_9020),
		.dout(new_net_9021)
	);

	bfr new_net_9022_bfr_after (
		.din(new_net_9021),
		.dout(new_net_9022)
	);

	bfr new_net_9023_bfr_after (
		.din(new_net_9022),
		.dout(new_net_9023)
	);

	bfr new_net_9024_bfr_after (
		.din(new_net_9023),
		.dout(new_net_9024)
	);

	bfr new_net_9025_bfr_after (
		.din(new_net_9024),
		.dout(new_net_9025)
	);

	bfr new_net_9026_bfr_after (
		.din(new_net_9025),
		.dout(new_net_9026)
	);

	bfr new_net_9027_bfr_after (
		.din(new_net_9026),
		.dout(new_net_9027)
	);

	bfr new_net_9028_bfr_after (
		.din(new_net_9027),
		.dout(new_net_9028)
	);

	bfr new_net_9029_bfr_after (
		.din(new_net_9028),
		.dout(new_net_9029)
	);

	bfr new_net_9030_bfr_after (
		.din(new_net_9029),
		.dout(new_net_9030)
	);

	bfr new_net_9031_bfr_after (
		.din(new_net_9030),
		.dout(new_net_9031)
	);

	bfr new_net_9032_bfr_after (
		.din(new_net_9031),
		.dout(new_net_9032)
	);

	bfr new_net_9033_bfr_after (
		.din(new_net_9032),
		.dout(new_net_9033)
	);

	bfr new_net_9034_bfr_after (
		.din(new_net_9033),
		.dout(new_net_9034)
	);

	bfr new_net_9035_bfr_after (
		.din(new_net_9034),
		.dout(new_net_9035)
	);

	bfr new_net_9036_bfr_after (
		.din(new_net_9035),
		.dout(new_net_9036)
	);

	bfr new_net_9037_bfr_after (
		.din(new_net_9036),
		.dout(new_net_9037)
	);

	bfr new_net_9038_bfr_after (
		.din(new_net_9037),
		.dout(new_net_9038)
	);

	bfr new_net_9039_bfr_after (
		.din(new_net_9038),
		.dout(new_net_9039)
	);

	bfr new_net_9040_bfr_after (
		.din(new_net_9039),
		.dout(new_net_9040)
	);

	spl2 _1288__v_fanout (
		.a(new_net_9040),
		.b(new_net_1892),
		.c(new_net_1893)
	);

	spl2 _0764__v_fanout (
		.a(_0764_),
		.b(new_net_182),
		.c(new_net_183)
	);

	spl2 _1031__v_fanout (
		.a(_1031_),
		.b(new_net_335),
		.c(new_net_336)
	);

	bfr new_net_9041_bfr_after (
		.din(_1582_),
		.dout(new_net_9041)
	);

	bfr new_net_9042_bfr_after (
		.din(new_net_9041),
		.dout(new_net_9042)
	);

	bfr new_net_9043_bfr_after (
		.din(new_net_9042),
		.dout(new_net_9043)
	);

	bfr new_net_9044_bfr_after (
		.din(new_net_9043),
		.dout(new_net_9044)
	);

	bfr new_net_9045_bfr_after (
		.din(new_net_9044),
		.dout(new_net_9045)
	);

	bfr new_net_9046_bfr_after (
		.din(new_net_9045),
		.dout(new_net_9046)
	);

	bfr new_net_9047_bfr_after (
		.din(new_net_9046),
		.dout(new_net_9047)
	);

	bfr new_net_9048_bfr_after (
		.din(new_net_9047),
		.dout(new_net_9048)
	);

	bfr new_net_9049_bfr_after (
		.din(new_net_9048),
		.dout(new_net_9049)
	);

	bfr new_net_9050_bfr_after (
		.din(new_net_9049),
		.dout(new_net_9050)
	);

	bfr new_net_9051_bfr_after (
		.din(new_net_9050),
		.dout(new_net_9051)
	);

	bfr new_net_9052_bfr_after (
		.din(new_net_9051),
		.dout(new_net_9052)
	);

	bfr new_net_9053_bfr_after (
		.din(new_net_9052),
		.dout(new_net_9053)
	);

	bfr new_net_9054_bfr_after (
		.din(new_net_9053),
		.dout(new_net_9054)
	);

	bfr new_net_9055_bfr_after (
		.din(new_net_9054),
		.dout(new_net_9055)
	);

	bfr new_net_9056_bfr_after (
		.din(new_net_9055),
		.dout(new_net_9056)
	);

	bfr new_net_9057_bfr_after (
		.din(new_net_9056),
		.dout(new_net_9057)
	);

	bfr new_net_9058_bfr_after (
		.din(new_net_9057),
		.dout(new_net_9058)
	);

	bfr new_net_9059_bfr_after (
		.din(new_net_9058),
		.dout(new_net_9059)
	);

	bfr new_net_9060_bfr_after (
		.din(new_net_9059),
		.dout(new_net_9060)
	);

	bfr new_net_9061_bfr_after (
		.din(new_net_9060),
		.dout(new_net_9061)
	);

	bfr new_net_9062_bfr_after (
		.din(new_net_9061),
		.dout(new_net_9062)
	);

	bfr new_net_9063_bfr_after (
		.din(new_net_9062),
		.dout(new_net_9063)
	);

	bfr new_net_9064_bfr_after (
		.din(new_net_9063),
		.dout(new_net_9064)
	);

	spl2 _1582__v_fanout (
		.a(new_net_9064),
		.b(new_net_2114),
		.c(new_net_2115)
	);

	spl2 _1299__v_fanout (
		.a(_1299_),
		.b(new_net_962),
		.c(new_net_963)
	);

	bfr new_net_9065_bfr_after (
		.din(_1076_),
		.dout(new_net_9065)
	);

	bfr new_net_9066_bfr_after (
		.din(new_net_9065),
		.dout(new_net_9066)
	);

	bfr new_net_9067_bfr_after (
		.din(new_net_9066),
		.dout(new_net_9067)
	);

	bfr new_net_9068_bfr_after (
		.din(new_net_9067),
		.dout(new_net_9068)
	);

	bfr new_net_9069_bfr_after (
		.din(new_net_9068),
		.dout(new_net_9069)
	);

	bfr new_net_9070_bfr_after (
		.din(new_net_9069),
		.dout(new_net_9070)
	);

	bfr new_net_9071_bfr_after (
		.din(new_net_9070),
		.dout(new_net_9071)
	);

	bfr new_net_9072_bfr_after (
		.din(new_net_9071),
		.dout(new_net_9072)
	);

	bfr new_net_9073_bfr_after (
		.din(new_net_9072),
		.dout(new_net_9073)
	);

	bfr new_net_9074_bfr_after (
		.din(new_net_9073),
		.dout(new_net_9074)
	);

	bfr new_net_9075_bfr_after (
		.din(new_net_9074),
		.dout(new_net_9075)
	);

	bfr new_net_9076_bfr_after (
		.din(new_net_9075),
		.dout(new_net_9076)
	);

	bfr new_net_9077_bfr_after (
		.din(new_net_9076),
		.dout(new_net_9077)
	);

	bfr new_net_9078_bfr_after (
		.din(new_net_9077),
		.dout(new_net_9078)
	);

	bfr new_net_9079_bfr_after (
		.din(new_net_9078),
		.dout(new_net_9079)
	);

	bfr new_net_9080_bfr_after (
		.din(new_net_9079),
		.dout(new_net_9080)
	);

	bfr new_net_9081_bfr_after (
		.din(new_net_9080),
		.dout(new_net_9081)
	);

	bfr new_net_9082_bfr_after (
		.din(new_net_9081),
		.dout(new_net_9082)
	);

	bfr new_net_9083_bfr_after (
		.din(new_net_9082),
		.dout(new_net_9083)
	);

	bfr new_net_9084_bfr_after (
		.din(new_net_9083),
		.dout(new_net_9084)
	);

	bfr new_net_9085_bfr_after (
		.din(new_net_9084),
		.dout(new_net_9085)
	);

	bfr new_net_9086_bfr_after (
		.din(new_net_9085),
		.dout(new_net_9086)
	);

	bfr new_net_9087_bfr_after (
		.din(new_net_9086),
		.dout(new_net_9087)
	);

	bfr new_net_9088_bfr_after (
		.din(new_net_9087),
		.dout(new_net_9088)
	);

	bfr new_net_9089_bfr_after (
		.din(new_net_9088),
		.dout(new_net_9089)
	);

	bfr new_net_9090_bfr_after (
		.din(new_net_9089),
		.dout(new_net_9090)
	);

	bfr new_net_9091_bfr_after (
		.din(new_net_9090),
		.dout(new_net_9091)
	);

	bfr new_net_9092_bfr_after (
		.din(new_net_9091),
		.dout(new_net_9092)
	);

	bfr new_net_9093_bfr_after (
		.din(new_net_9092),
		.dout(new_net_9093)
	);

	bfr new_net_9094_bfr_after (
		.din(new_net_9093),
		.dout(new_net_9094)
	);

	bfr new_net_9095_bfr_after (
		.din(new_net_9094),
		.dout(new_net_9095)
	);

	bfr new_net_9096_bfr_after (
		.din(new_net_9095),
		.dout(new_net_9096)
	);

	spl2 _1076__v_fanout (
		.a(new_net_9096),
		.b(new_net_2014),
		.c(new_net_2015)
	);

	bfr new_net_9097_bfr_after (
		.din(_0705_),
		.dout(new_net_9097)
	);

	bfr new_net_9098_bfr_after (
		.din(new_net_9097),
		.dout(new_net_9098)
	);

	bfr new_net_9099_bfr_after (
		.din(new_net_9098),
		.dout(new_net_9099)
	);

	bfr new_net_9100_bfr_after (
		.din(new_net_9099),
		.dout(new_net_9100)
	);

	bfr new_net_9101_bfr_after (
		.din(new_net_9100),
		.dout(new_net_9101)
	);

	bfr new_net_9102_bfr_after (
		.din(new_net_9101),
		.dout(new_net_9102)
	);

	bfr new_net_9103_bfr_after (
		.din(new_net_9102),
		.dout(new_net_9103)
	);

	bfr new_net_9104_bfr_after (
		.din(new_net_9103),
		.dout(new_net_9104)
	);

	bfr new_net_9105_bfr_after (
		.din(new_net_9104),
		.dout(new_net_9105)
	);

	bfr new_net_9106_bfr_after (
		.din(new_net_9105),
		.dout(new_net_9106)
	);

	bfr new_net_9107_bfr_after (
		.din(new_net_9106),
		.dout(new_net_9107)
	);

	bfr new_net_9108_bfr_after (
		.din(new_net_9107),
		.dout(new_net_9108)
	);

	bfr new_net_9109_bfr_after (
		.din(new_net_9108),
		.dout(new_net_9109)
	);

	bfr new_net_9110_bfr_after (
		.din(new_net_9109),
		.dout(new_net_9110)
	);

	bfr new_net_9111_bfr_after (
		.din(new_net_9110),
		.dout(new_net_9111)
	);

	bfr new_net_9112_bfr_after (
		.din(new_net_9111),
		.dout(new_net_9112)
	);

	bfr new_net_9113_bfr_after (
		.din(new_net_9112),
		.dout(new_net_9113)
	);

	bfr new_net_9114_bfr_after (
		.din(new_net_9113),
		.dout(new_net_9114)
	);

	bfr new_net_9115_bfr_after (
		.din(new_net_9114),
		.dout(new_net_9115)
	);

	bfr new_net_9116_bfr_after (
		.din(new_net_9115),
		.dout(new_net_9116)
	);

	bfr new_net_9117_bfr_after (
		.din(new_net_9116),
		.dout(new_net_9117)
	);

	bfr new_net_9118_bfr_after (
		.din(new_net_9117),
		.dout(new_net_9118)
	);

	bfr new_net_9119_bfr_after (
		.din(new_net_9118),
		.dout(new_net_9119)
	);

	bfr new_net_9120_bfr_after (
		.din(new_net_9119),
		.dout(new_net_9120)
	);

	bfr new_net_9121_bfr_after (
		.din(new_net_9120),
		.dout(new_net_9121)
	);

	bfr new_net_9122_bfr_after (
		.din(new_net_9121),
		.dout(new_net_9122)
	);

	bfr new_net_9123_bfr_after (
		.din(new_net_9122),
		.dout(new_net_9123)
	);

	bfr new_net_9124_bfr_after (
		.din(new_net_9123),
		.dout(new_net_9124)
	);

	bfr new_net_9125_bfr_after (
		.din(new_net_9124),
		.dout(new_net_9125)
	);

	bfr new_net_9126_bfr_after (
		.din(new_net_9125),
		.dout(new_net_9126)
	);

	bfr new_net_9127_bfr_after (
		.din(new_net_9126),
		.dout(new_net_9127)
	);

	bfr new_net_9128_bfr_after (
		.din(new_net_9127),
		.dout(new_net_9128)
	);

	bfr new_net_9129_bfr_after (
		.din(new_net_9128),
		.dout(new_net_9129)
	);

	bfr new_net_9130_bfr_after (
		.din(new_net_9129),
		.dout(new_net_9130)
	);

	bfr new_net_9131_bfr_after (
		.din(new_net_9130),
		.dout(new_net_9131)
	);

	bfr new_net_9132_bfr_after (
		.din(new_net_9131),
		.dout(new_net_9132)
	);

	bfr new_net_9133_bfr_after (
		.din(new_net_9132),
		.dout(new_net_9133)
	);

	bfr new_net_9134_bfr_after (
		.din(new_net_9133),
		.dout(new_net_9134)
	);

	bfr new_net_9135_bfr_after (
		.din(new_net_9134),
		.dout(new_net_9135)
	);

	bfr new_net_9136_bfr_after (
		.din(new_net_9135),
		.dout(new_net_9136)
	);

	bfr new_net_9137_bfr_after (
		.din(new_net_9136),
		.dout(new_net_9137)
	);

	bfr new_net_9138_bfr_after (
		.din(new_net_9137),
		.dout(new_net_9138)
	);

	bfr new_net_9139_bfr_after (
		.din(new_net_9138),
		.dout(new_net_9139)
	);

	bfr new_net_9140_bfr_after (
		.din(new_net_9139),
		.dout(new_net_9140)
	);

	bfr new_net_9141_bfr_after (
		.din(new_net_9140),
		.dout(new_net_9141)
	);

	bfr new_net_9142_bfr_after (
		.din(new_net_9141),
		.dout(new_net_9142)
	);

	bfr new_net_9143_bfr_after (
		.din(new_net_9142),
		.dout(new_net_9143)
	);

	bfr new_net_9144_bfr_after (
		.din(new_net_9143),
		.dout(new_net_9144)
	);

	bfr new_net_9145_bfr_after (
		.din(new_net_9144),
		.dout(new_net_9145)
	);

	bfr new_net_9146_bfr_after (
		.din(new_net_9145),
		.dout(new_net_9146)
	);

	bfr new_net_9147_bfr_after (
		.din(new_net_9146),
		.dout(new_net_9147)
	);

	bfr new_net_9148_bfr_after (
		.din(new_net_9147),
		.dout(new_net_9148)
	);

	bfr new_net_9149_bfr_after (
		.din(new_net_9148),
		.dout(new_net_9149)
	);

	bfr new_net_9150_bfr_after (
		.din(new_net_9149),
		.dout(new_net_9150)
	);

	bfr new_net_9151_bfr_after (
		.din(new_net_9150),
		.dout(new_net_9151)
	);

	bfr new_net_9152_bfr_after (
		.din(new_net_9151),
		.dout(new_net_9152)
	);

	bfr new_net_9153_bfr_after (
		.din(new_net_9152),
		.dout(new_net_9153)
	);

	bfr new_net_9154_bfr_after (
		.din(new_net_9153),
		.dout(new_net_9154)
	);

	bfr new_net_9155_bfr_after (
		.din(new_net_9154),
		.dout(new_net_9155)
	);

	bfr new_net_9156_bfr_after (
		.din(new_net_9155),
		.dout(new_net_9156)
	);

	bfr new_net_9157_bfr_after (
		.din(new_net_9156),
		.dout(new_net_9157)
	);

	bfr new_net_9158_bfr_after (
		.din(new_net_9157),
		.dout(new_net_9158)
	);

	bfr new_net_9159_bfr_after (
		.din(new_net_9158),
		.dout(new_net_9159)
	);

	bfr new_net_9160_bfr_after (
		.din(new_net_9159),
		.dout(new_net_9160)
	);

	bfr new_net_9161_bfr_after (
		.din(new_net_9160),
		.dout(new_net_9161)
	);

	bfr new_net_9162_bfr_after (
		.din(new_net_9161),
		.dout(new_net_9162)
	);

	bfr new_net_9163_bfr_after (
		.din(new_net_9162),
		.dout(new_net_9163)
	);

	bfr new_net_9164_bfr_after (
		.din(new_net_9163),
		.dout(new_net_9164)
	);

	bfr new_net_9165_bfr_after (
		.din(new_net_9164),
		.dout(new_net_9165)
	);

	bfr new_net_9166_bfr_after (
		.din(new_net_9165),
		.dout(new_net_9166)
	);

	bfr new_net_9167_bfr_after (
		.din(new_net_9166),
		.dout(new_net_9167)
	);

	bfr new_net_9168_bfr_after (
		.din(new_net_9167),
		.dout(new_net_9168)
	);

	bfr new_net_9169_bfr_after (
		.din(new_net_9168),
		.dout(new_net_9169)
	);

	bfr new_net_9170_bfr_after (
		.din(new_net_9169),
		.dout(new_net_9170)
	);

	bfr new_net_9171_bfr_after (
		.din(new_net_9170),
		.dout(new_net_9171)
	);

	bfr new_net_9172_bfr_after (
		.din(new_net_9171),
		.dout(new_net_9172)
	);

	bfr new_net_9173_bfr_after (
		.din(new_net_9172),
		.dout(new_net_9173)
	);

	bfr new_net_9174_bfr_after (
		.din(new_net_9173),
		.dout(new_net_9174)
	);

	bfr new_net_9175_bfr_after (
		.din(new_net_9174),
		.dout(new_net_9175)
	);

	bfr new_net_9176_bfr_after (
		.din(new_net_9175),
		.dout(new_net_9176)
	);

	spl2 _0705__v_fanout (
		.a(new_net_9176),
		.b(new_net_84),
		.c(new_net_85)
	);

	bfr new_net_9177_bfr_after (
		.din(_0837_),
		.dout(new_net_9177)
	);

	bfr new_net_9178_bfr_after (
		.din(new_net_9177),
		.dout(new_net_9178)
	);

	bfr new_net_9179_bfr_after (
		.din(new_net_9178),
		.dout(new_net_9179)
	);

	bfr new_net_9180_bfr_after (
		.din(new_net_9179),
		.dout(new_net_9180)
	);

	bfr new_net_9181_bfr_after (
		.din(new_net_9180),
		.dout(new_net_9181)
	);

	bfr new_net_9182_bfr_after (
		.din(new_net_9181),
		.dout(new_net_9182)
	);

	bfr new_net_9183_bfr_after (
		.din(new_net_9182),
		.dout(new_net_9183)
	);

	bfr new_net_9184_bfr_after (
		.din(new_net_9183),
		.dout(new_net_9184)
	);

	bfr new_net_9185_bfr_after (
		.din(new_net_9184),
		.dout(new_net_9185)
	);

	bfr new_net_9186_bfr_after (
		.din(new_net_9185),
		.dout(new_net_9186)
	);

	bfr new_net_9187_bfr_after (
		.din(new_net_9186),
		.dout(new_net_9187)
	);

	bfr new_net_9188_bfr_after (
		.din(new_net_9187),
		.dout(new_net_9188)
	);

	bfr new_net_9189_bfr_after (
		.din(new_net_9188),
		.dout(new_net_9189)
	);

	bfr new_net_9190_bfr_after (
		.din(new_net_9189),
		.dout(new_net_9190)
	);

	bfr new_net_9191_bfr_after (
		.din(new_net_9190),
		.dout(new_net_9191)
	);

	bfr new_net_9192_bfr_after (
		.din(new_net_9191),
		.dout(new_net_9192)
	);

	bfr new_net_9193_bfr_after (
		.din(new_net_9192),
		.dout(new_net_9193)
	);

	bfr new_net_9194_bfr_after (
		.din(new_net_9193),
		.dout(new_net_9194)
	);

	bfr new_net_9195_bfr_after (
		.din(new_net_9194),
		.dout(new_net_9195)
	);

	bfr new_net_9196_bfr_after (
		.din(new_net_9195),
		.dout(new_net_9196)
	);

	bfr new_net_9197_bfr_after (
		.din(new_net_9196),
		.dout(new_net_9197)
	);

	bfr new_net_9198_bfr_after (
		.din(new_net_9197),
		.dout(new_net_9198)
	);

	bfr new_net_9199_bfr_after (
		.din(new_net_9198),
		.dout(new_net_9199)
	);

	bfr new_net_9200_bfr_after (
		.din(new_net_9199),
		.dout(new_net_9200)
	);

	bfr new_net_9201_bfr_after (
		.din(new_net_9200),
		.dout(new_net_9201)
	);

	bfr new_net_9202_bfr_after (
		.din(new_net_9201),
		.dout(new_net_9202)
	);

	bfr new_net_9203_bfr_after (
		.din(new_net_9202),
		.dout(new_net_9203)
	);

	bfr new_net_9204_bfr_after (
		.din(new_net_9203),
		.dout(new_net_9204)
	);

	bfr new_net_9205_bfr_after (
		.din(new_net_9204),
		.dout(new_net_9205)
	);

	bfr new_net_9206_bfr_after (
		.din(new_net_9205),
		.dout(new_net_9206)
	);

	bfr new_net_9207_bfr_after (
		.din(new_net_9206),
		.dout(new_net_9207)
	);

	bfr new_net_9208_bfr_after (
		.din(new_net_9207),
		.dout(new_net_9208)
	);

	bfr new_net_9209_bfr_after (
		.din(new_net_9208),
		.dout(new_net_9209)
	);

	bfr new_net_9210_bfr_after (
		.din(new_net_9209),
		.dout(new_net_9210)
	);

	bfr new_net_9211_bfr_after (
		.din(new_net_9210),
		.dout(new_net_9211)
	);

	bfr new_net_9212_bfr_after (
		.din(new_net_9211),
		.dout(new_net_9212)
	);

	bfr new_net_9213_bfr_after (
		.din(new_net_9212),
		.dout(new_net_9213)
	);

	bfr new_net_9214_bfr_after (
		.din(new_net_9213),
		.dout(new_net_9214)
	);

	bfr new_net_9215_bfr_after (
		.din(new_net_9214),
		.dout(new_net_9215)
	);

	bfr new_net_9216_bfr_after (
		.din(new_net_9215),
		.dout(new_net_9216)
	);

	bfr new_net_9217_bfr_after (
		.din(new_net_9216),
		.dout(new_net_9217)
	);

	bfr new_net_9218_bfr_after (
		.din(new_net_9217),
		.dout(new_net_9218)
	);

	bfr new_net_9219_bfr_after (
		.din(new_net_9218),
		.dout(new_net_9219)
	);

	bfr new_net_9220_bfr_after (
		.din(new_net_9219),
		.dout(new_net_9220)
	);

	bfr new_net_9221_bfr_after (
		.din(new_net_9220),
		.dout(new_net_9221)
	);

	bfr new_net_9222_bfr_after (
		.din(new_net_9221),
		.dout(new_net_9222)
	);

	bfr new_net_9223_bfr_after (
		.din(new_net_9222),
		.dout(new_net_9223)
	);

	bfr new_net_9224_bfr_after (
		.din(new_net_9223),
		.dout(new_net_9224)
	);

	bfr new_net_9225_bfr_after (
		.din(new_net_9224),
		.dout(new_net_9225)
	);

	bfr new_net_9226_bfr_after (
		.din(new_net_9225),
		.dout(new_net_9226)
	);

	bfr new_net_9227_bfr_after (
		.din(new_net_9226),
		.dout(new_net_9227)
	);

	bfr new_net_9228_bfr_after (
		.din(new_net_9227),
		.dout(new_net_9228)
	);

	bfr new_net_9229_bfr_after (
		.din(new_net_9228),
		.dout(new_net_9229)
	);

	bfr new_net_9230_bfr_after (
		.din(new_net_9229),
		.dout(new_net_9230)
	);

	bfr new_net_9231_bfr_after (
		.din(new_net_9230),
		.dout(new_net_9231)
	);

	bfr new_net_9232_bfr_after (
		.din(new_net_9231),
		.dout(new_net_9232)
	);

	bfr new_net_9233_bfr_after (
		.din(new_net_9232),
		.dout(new_net_9233)
	);

	bfr new_net_9234_bfr_after (
		.din(new_net_9233),
		.dout(new_net_9234)
	);

	bfr new_net_9235_bfr_after (
		.din(new_net_9234),
		.dout(new_net_9235)
	);

	bfr new_net_9236_bfr_after (
		.din(new_net_9235),
		.dout(new_net_9236)
	);

	bfr new_net_9237_bfr_after (
		.din(new_net_9236),
		.dout(new_net_9237)
	);

	bfr new_net_9238_bfr_after (
		.din(new_net_9237),
		.dout(new_net_9238)
	);

	bfr new_net_9239_bfr_after (
		.din(new_net_9238),
		.dout(new_net_9239)
	);

	bfr new_net_9240_bfr_after (
		.din(new_net_9239),
		.dout(new_net_9240)
	);

	bfr new_net_9241_bfr_after (
		.din(new_net_9240),
		.dout(new_net_9241)
	);

	bfr new_net_9242_bfr_after (
		.din(new_net_9241),
		.dout(new_net_9242)
	);

	bfr new_net_9243_bfr_after (
		.din(new_net_9242),
		.dout(new_net_9243)
	);

	bfr new_net_9244_bfr_after (
		.din(new_net_9243),
		.dout(new_net_9244)
	);

	bfr new_net_9245_bfr_after (
		.din(new_net_9244),
		.dout(new_net_9245)
	);

	bfr new_net_9246_bfr_after (
		.din(new_net_9245),
		.dout(new_net_9246)
	);

	bfr new_net_9247_bfr_after (
		.din(new_net_9246),
		.dout(new_net_9247)
	);

	bfr new_net_9248_bfr_after (
		.din(new_net_9247),
		.dout(new_net_9248)
	);

	bfr new_net_9249_bfr_after (
		.din(new_net_9248),
		.dout(new_net_9249)
	);

	bfr new_net_9250_bfr_after (
		.din(new_net_9249),
		.dout(new_net_9250)
	);

	spl2 _0837__v_fanout (
		.a(new_net_9250),
		.b(new_net_2535),
		.c(new_net_2536)
	);

	bfr new_net_9251_bfr_after (
		.din(_1278_),
		.dout(new_net_9251)
	);

	bfr new_net_9252_bfr_after (
		.din(new_net_9251),
		.dout(new_net_9252)
	);

	bfr new_net_9253_bfr_after (
		.din(new_net_9252),
		.dout(new_net_9253)
	);

	bfr new_net_9254_bfr_after (
		.din(new_net_9253),
		.dout(new_net_9254)
	);

	bfr new_net_9255_bfr_after (
		.din(new_net_9254),
		.dout(new_net_9255)
	);

	bfr new_net_9256_bfr_after (
		.din(new_net_9255),
		.dout(new_net_9256)
	);

	bfr new_net_9257_bfr_after (
		.din(new_net_9256),
		.dout(new_net_9257)
	);

	bfr new_net_9258_bfr_after (
		.din(new_net_9257),
		.dout(new_net_9258)
	);

	bfr new_net_9259_bfr_after (
		.din(new_net_9258),
		.dout(new_net_9259)
	);

	bfr new_net_9260_bfr_after (
		.din(new_net_9259),
		.dout(new_net_9260)
	);

	bfr new_net_9261_bfr_after (
		.din(new_net_9260),
		.dout(new_net_9261)
	);

	bfr new_net_9262_bfr_after (
		.din(new_net_9261),
		.dout(new_net_9262)
	);

	bfr new_net_9263_bfr_after (
		.din(new_net_9262),
		.dout(new_net_9263)
	);

	bfr new_net_9264_bfr_after (
		.din(new_net_9263),
		.dout(new_net_9264)
	);

	bfr new_net_9265_bfr_after (
		.din(new_net_9264),
		.dout(new_net_9265)
	);

	bfr new_net_9266_bfr_after (
		.din(new_net_9265),
		.dout(new_net_9266)
	);

	bfr new_net_9267_bfr_after (
		.din(new_net_9266),
		.dout(new_net_9267)
	);

	bfr new_net_9268_bfr_after (
		.din(new_net_9267),
		.dout(new_net_9268)
	);

	bfr new_net_9269_bfr_after (
		.din(new_net_9268),
		.dout(new_net_9269)
	);

	bfr new_net_9270_bfr_after (
		.din(new_net_9269),
		.dout(new_net_9270)
	);

	bfr new_net_9271_bfr_after (
		.din(new_net_9270),
		.dout(new_net_9271)
	);

	bfr new_net_9272_bfr_after (
		.din(new_net_9271),
		.dout(new_net_9272)
	);

	bfr new_net_9273_bfr_after (
		.din(new_net_9272),
		.dout(new_net_9273)
	);

	bfr new_net_9274_bfr_after (
		.din(new_net_9273),
		.dout(new_net_9274)
	);

	bfr new_net_9275_bfr_after (
		.din(new_net_9274),
		.dout(new_net_9275)
	);

	bfr new_net_9276_bfr_after (
		.din(new_net_9275),
		.dout(new_net_9276)
	);

	bfr new_net_9277_bfr_after (
		.din(new_net_9276),
		.dout(new_net_9277)
	);

	bfr new_net_9278_bfr_after (
		.din(new_net_9277),
		.dout(new_net_9278)
	);

	bfr new_net_9279_bfr_after (
		.din(new_net_9278),
		.dout(new_net_9279)
	);

	bfr new_net_9280_bfr_after (
		.din(new_net_9279),
		.dout(new_net_9280)
	);

	bfr new_net_9281_bfr_after (
		.din(new_net_9280),
		.dout(new_net_9281)
	);

	bfr new_net_9282_bfr_after (
		.din(new_net_9281),
		.dout(new_net_9282)
	);

	bfr new_net_9283_bfr_after (
		.din(new_net_9282),
		.dout(new_net_9283)
	);

	bfr new_net_9284_bfr_after (
		.din(new_net_9283),
		.dout(new_net_9284)
	);

	bfr new_net_9285_bfr_after (
		.din(new_net_9284),
		.dout(new_net_9285)
	);

	bfr new_net_9286_bfr_after (
		.din(new_net_9285),
		.dout(new_net_9286)
	);

	bfr new_net_9287_bfr_after (
		.din(new_net_9286),
		.dout(new_net_9287)
	);

	bfr new_net_9288_bfr_after (
		.din(new_net_9287),
		.dout(new_net_9288)
	);

	bfr new_net_9289_bfr_after (
		.din(new_net_9288),
		.dout(new_net_9289)
	);

	bfr new_net_9290_bfr_after (
		.din(new_net_9289),
		.dout(new_net_9290)
	);

	bfr new_net_9291_bfr_after (
		.din(new_net_9290),
		.dout(new_net_9291)
	);

	bfr new_net_9292_bfr_after (
		.din(new_net_9291),
		.dout(new_net_9292)
	);

	bfr new_net_9293_bfr_after (
		.din(new_net_9292),
		.dout(new_net_9293)
	);

	bfr new_net_9294_bfr_after (
		.din(new_net_9293),
		.dout(new_net_9294)
	);

	bfr new_net_9295_bfr_after (
		.din(new_net_9294),
		.dout(new_net_9295)
	);

	bfr new_net_9296_bfr_after (
		.din(new_net_9295),
		.dout(new_net_9296)
	);

	bfr new_net_9297_bfr_after (
		.din(new_net_9296),
		.dout(new_net_9297)
	);

	bfr new_net_9298_bfr_after (
		.din(new_net_9297),
		.dout(new_net_9298)
	);

	bfr new_net_9299_bfr_after (
		.din(new_net_9298),
		.dout(new_net_9299)
	);

	bfr new_net_9300_bfr_after (
		.din(new_net_9299),
		.dout(new_net_9300)
	);

	bfr new_net_9301_bfr_after (
		.din(new_net_9300),
		.dout(new_net_9301)
	);

	bfr new_net_9302_bfr_after (
		.din(new_net_9301),
		.dout(new_net_9302)
	);

	bfr new_net_9303_bfr_after (
		.din(new_net_9302),
		.dout(new_net_9303)
	);

	bfr new_net_9304_bfr_after (
		.din(new_net_9303),
		.dout(new_net_9304)
	);

	bfr new_net_9305_bfr_after (
		.din(new_net_9304),
		.dout(new_net_9305)
	);

	bfr new_net_9306_bfr_after (
		.din(new_net_9305),
		.dout(new_net_9306)
	);

	bfr new_net_9307_bfr_after (
		.din(new_net_9306),
		.dout(new_net_9307)
	);

	bfr new_net_9308_bfr_after (
		.din(new_net_9307),
		.dout(new_net_9308)
	);

	bfr new_net_9309_bfr_after (
		.din(new_net_9308),
		.dout(new_net_9309)
	);

	bfr new_net_9310_bfr_after (
		.din(new_net_9309),
		.dout(new_net_9310)
	);

	bfr new_net_9311_bfr_after (
		.din(new_net_9310),
		.dout(new_net_9311)
	);

	bfr new_net_9312_bfr_after (
		.din(new_net_9311),
		.dout(new_net_9312)
	);

	bfr new_net_9313_bfr_after (
		.din(new_net_9312),
		.dout(new_net_9313)
	);

	bfr new_net_9314_bfr_after (
		.din(new_net_9313),
		.dout(new_net_9314)
	);

	bfr new_net_9315_bfr_after (
		.din(new_net_9314),
		.dout(new_net_9315)
	);

	bfr new_net_9316_bfr_after (
		.din(new_net_9315),
		.dout(new_net_9316)
	);

	bfr new_net_9317_bfr_after (
		.din(new_net_9316),
		.dout(new_net_9317)
	);

	bfr new_net_9318_bfr_after (
		.din(new_net_9317),
		.dout(new_net_9318)
	);

	bfr new_net_9319_bfr_after (
		.din(new_net_9318),
		.dout(new_net_9319)
	);

	bfr new_net_9320_bfr_after (
		.din(new_net_9319),
		.dout(new_net_9320)
	);

	bfr new_net_9321_bfr_after (
		.din(new_net_9320),
		.dout(new_net_9321)
	);

	bfr new_net_9322_bfr_after (
		.din(new_net_9321),
		.dout(new_net_9322)
	);

	bfr new_net_9323_bfr_after (
		.din(new_net_9322),
		.dout(new_net_9323)
	);

	bfr new_net_9324_bfr_after (
		.din(new_net_9323),
		.dout(new_net_9324)
	);

	bfr new_net_9325_bfr_after (
		.din(new_net_9324),
		.dout(new_net_9325)
	);

	bfr new_net_9326_bfr_after (
		.din(new_net_9325),
		.dout(new_net_9326)
	);

	bfr new_net_9327_bfr_after (
		.din(new_net_9326),
		.dout(new_net_9327)
	);

	bfr new_net_9328_bfr_after (
		.din(new_net_9327),
		.dout(new_net_9328)
	);

	bfr new_net_9329_bfr_after (
		.din(new_net_9328),
		.dout(new_net_9329)
	);

	bfr new_net_9330_bfr_after (
		.din(new_net_9329),
		.dout(new_net_9330)
	);

	spl2 _1278__v_fanout (
		.a(new_net_9330),
		.b(new_net_172),
		.c(new_net_173)
	);

	bfr new_net_9331_bfr_after (
		.din(_0232_),
		.dout(new_net_9331)
	);

	bfr new_net_9332_bfr_after (
		.din(new_net_9331),
		.dout(new_net_9332)
	);

	bfr new_net_9333_bfr_after (
		.din(new_net_9332),
		.dout(new_net_9333)
	);

	bfr new_net_9334_bfr_after (
		.din(new_net_9333),
		.dout(new_net_9334)
	);

	bfr new_net_9335_bfr_after (
		.din(new_net_9334),
		.dout(new_net_9335)
	);

	bfr new_net_9336_bfr_after (
		.din(new_net_9335),
		.dout(new_net_9336)
	);

	bfr new_net_9337_bfr_after (
		.din(new_net_9336),
		.dout(new_net_9337)
	);

	bfr new_net_9338_bfr_after (
		.din(new_net_9337),
		.dout(new_net_9338)
	);

	bfr new_net_9339_bfr_after (
		.din(new_net_9338),
		.dout(new_net_9339)
	);

	bfr new_net_9340_bfr_after (
		.din(new_net_9339),
		.dout(new_net_9340)
	);

	bfr new_net_9341_bfr_after (
		.din(new_net_9340),
		.dout(new_net_9341)
	);

	bfr new_net_9342_bfr_after (
		.din(new_net_9341),
		.dout(new_net_9342)
	);

	bfr new_net_9343_bfr_after (
		.din(new_net_9342),
		.dout(new_net_9343)
	);

	bfr new_net_9344_bfr_after (
		.din(new_net_9343),
		.dout(new_net_9344)
	);

	bfr new_net_9345_bfr_after (
		.din(new_net_9344),
		.dout(new_net_9345)
	);

	bfr new_net_9346_bfr_after (
		.din(new_net_9345),
		.dout(new_net_9346)
	);

	bfr new_net_9347_bfr_after (
		.din(new_net_9346),
		.dout(new_net_9347)
	);

	bfr new_net_9348_bfr_after (
		.din(new_net_9347),
		.dout(new_net_9348)
	);

	bfr new_net_9349_bfr_after (
		.din(new_net_9348),
		.dout(new_net_9349)
	);

	bfr new_net_9350_bfr_after (
		.din(new_net_9349),
		.dout(new_net_9350)
	);

	bfr new_net_9351_bfr_after (
		.din(new_net_9350),
		.dout(new_net_9351)
	);

	bfr new_net_9352_bfr_after (
		.din(new_net_9351),
		.dout(new_net_9352)
	);

	bfr new_net_9353_bfr_after (
		.din(new_net_9352),
		.dout(new_net_9353)
	);

	bfr new_net_9354_bfr_after (
		.din(new_net_9353),
		.dout(new_net_9354)
	);

	bfr new_net_9355_bfr_after (
		.din(new_net_9354),
		.dout(new_net_9355)
	);

	bfr new_net_9356_bfr_after (
		.din(new_net_9355),
		.dout(new_net_9356)
	);

	bfr new_net_9357_bfr_after (
		.din(new_net_9356),
		.dout(new_net_9357)
	);

	bfr new_net_9358_bfr_after (
		.din(new_net_9357),
		.dout(new_net_9358)
	);

	bfr new_net_9359_bfr_after (
		.din(new_net_9358),
		.dout(new_net_9359)
	);

	bfr new_net_9360_bfr_after (
		.din(new_net_9359),
		.dout(new_net_9360)
	);

	bfr new_net_9361_bfr_after (
		.din(new_net_9360),
		.dout(new_net_9361)
	);

	bfr new_net_9362_bfr_after (
		.din(new_net_9361),
		.dout(new_net_9362)
	);

	bfr new_net_9363_bfr_after (
		.din(new_net_9362),
		.dout(new_net_9363)
	);

	bfr new_net_9364_bfr_after (
		.din(new_net_9363),
		.dout(new_net_9364)
	);

	bfr new_net_9365_bfr_after (
		.din(new_net_9364),
		.dout(new_net_9365)
	);

	bfr new_net_9366_bfr_after (
		.din(new_net_9365),
		.dout(new_net_9366)
	);

	bfr new_net_9367_bfr_after (
		.din(new_net_9366),
		.dout(new_net_9367)
	);

	bfr new_net_9368_bfr_after (
		.din(new_net_9367),
		.dout(new_net_9368)
	);

	bfr new_net_9369_bfr_after (
		.din(new_net_9368),
		.dout(new_net_9369)
	);

	bfr new_net_9370_bfr_after (
		.din(new_net_9369),
		.dout(new_net_9370)
	);

	spl2 _0232__v_fanout (
		.a(new_net_9370),
		.b(new_net_311),
		.c(new_net_312)
	);

	bfr new_net_9371_bfr_after (
		.din(_0835_),
		.dout(new_net_9371)
	);

	bfr new_net_9372_bfr_after (
		.din(new_net_9371),
		.dout(new_net_9372)
	);

	bfr new_net_9373_bfr_after (
		.din(new_net_9372),
		.dout(new_net_9373)
	);

	bfr new_net_9374_bfr_after (
		.din(new_net_9373),
		.dout(new_net_9374)
	);

	bfr new_net_9375_bfr_after (
		.din(new_net_9374),
		.dout(new_net_9375)
	);

	bfr new_net_9376_bfr_after (
		.din(new_net_9375),
		.dout(new_net_9376)
	);

	bfr new_net_9377_bfr_after (
		.din(new_net_9376),
		.dout(new_net_9377)
	);

	bfr new_net_9378_bfr_after (
		.din(new_net_9377),
		.dout(new_net_9378)
	);

	bfr new_net_9379_bfr_after (
		.din(new_net_9378),
		.dout(new_net_9379)
	);

	bfr new_net_9380_bfr_after (
		.din(new_net_9379),
		.dout(new_net_9380)
	);

	bfr new_net_9381_bfr_after (
		.din(new_net_9380),
		.dout(new_net_9381)
	);

	bfr new_net_9382_bfr_after (
		.din(new_net_9381),
		.dout(new_net_9382)
	);

	bfr new_net_9383_bfr_after (
		.din(new_net_9382),
		.dout(new_net_9383)
	);

	bfr new_net_9384_bfr_after (
		.din(new_net_9383),
		.dout(new_net_9384)
	);

	bfr new_net_9385_bfr_after (
		.din(new_net_9384),
		.dout(new_net_9385)
	);

	bfr new_net_9386_bfr_after (
		.din(new_net_9385),
		.dout(new_net_9386)
	);

	bfr new_net_9387_bfr_after (
		.din(new_net_9386),
		.dout(new_net_9387)
	);

	bfr new_net_9388_bfr_after (
		.din(new_net_9387),
		.dout(new_net_9388)
	);

	bfr new_net_9389_bfr_after (
		.din(new_net_9388),
		.dout(new_net_9389)
	);

	bfr new_net_9390_bfr_after (
		.din(new_net_9389),
		.dout(new_net_9390)
	);

	bfr new_net_9391_bfr_after (
		.din(new_net_9390),
		.dout(new_net_9391)
	);

	bfr new_net_9392_bfr_after (
		.din(new_net_9391),
		.dout(new_net_9392)
	);

	bfr new_net_9393_bfr_after (
		.din(new_net_9392),
		.dout(new_net_9393)
	);

	bfr new_net_9394_bfr_after (
		.din(new_net_9393),
		.dout(new_net_9394)
	);

	bfr new_net_9395_bfr_after (
		.din(new_net_9394),
		.dout(new_net_9395)
	);

	bfr new_net_9396_bfr_after (
		.din(new_net_9395),
		.dout(new_net_9396)
	);

	bfr new_net_9397_bfr_after (
		.din(new_net_9396),
		.dout(new_net_9397)
	);

	bfr new_net_9398_bfr_after (
		.din(new_net_9397),
		.dout(new_net_9398)
	);

	bfr new_net_9399_bfr_after (
		.din(new_net_9398),
		.dout(new_net_9399)
	);

	bfr new_net_9400_bfr_after (
		.din(new_net_9399),
		.dout(new_net_9400)
	);

	bfr new_net_9401_bfr_after (
		.din(new_net_9400),
		.dout(new_net_9401)
	);

	bfr new_net_9402_bfr_after (
		.din(new_net_9401),
		.dout(new_net_9402)
	);

	bfr new_net_9403_bfr_after (
		.din(new_net_9402),
		.dout(new_net_9403)
	);

	bfr new_net_9404_bfr_after (
		.din(new_net_9403),
		.dout(new_net_9404)
	);

	bfr new_net_9405_bfr_after (
		.din(new_net_9404),
		.dout(new_net_9405)
	);

	bfr new_net_9406_bfr_after (
		.din(new_net_9405),
		.dout(new_net_9406)
	);

	bfr new_net_9407_bfr_after (
		.din(new_net_9406),
		.dout(new_net_9407)
	);

	bfr new_net_9408_bfr_after (
		.din(new_net_9407),
		.dout(new_net_9408)
	);

	bfr new_net_9409_bfr_after (
		.din(new_net_9408),
		.dout(new_net_9409)
	);

	bfr new_net_9410_bfr_after (
		.din(new_net_9409),
		.dout(new_net_9410)
	);

	bfr new_net_9411_bfr_after (
		.din(new_net_9410),
		.dout(new_net_9411)
	);

	bfr new_net_9412_bfr_after (
		.din(new_net_9411),
		.dout(new_net_9412)
	);

	bfr new_net_9413_bfr_after (
		.din(new_net_9412),
		.dout(new_net_9413)
	);

	bfr new_net_9414_bfr_after (
		.din(new_net_9413),
		.dout(new_net_9414)
	);

	bfr new_net_9415_bfr_after (
		.din(new_net_9414),
		.dout(new_net_9415)
	);

	bfr new_net_9416_bfr_after (
		.din(new_net_9415),
		.dout(new_net_9416)
	);

	bfr new_net_9417_bfr_after (
		.din(new_net_9416),
		.dout(new_net_9417)
	);

	bfr new_net_9418_bfr_after (
		.din(new_net_9417),
		.dout(new_net_9418)
	);

	bfr new_net_9419_bfr_after (
		.din(new_net_9418),
		.dout(new_net_9419)
	);

	bfr new_net_9420_bfr_after (
		.din(new_net_9419),
		.dout(new_net_9420)
	);

	bfr new_net_9421_bfr_after (
		.din(new_net_9420),
		.dout(new_net_9421)
	);

	bfr new_net_9422_bfr_after (
		.din(new_net_9421),
		.dout(new_net_9422)
	);

	bfr new_net_9423_bfr_after (
		.din(new_net_9422),
		.dout(new_net_9423)
	);

	bfr new_net_9424_bfr_after (
		.din(new_net_9423),
		.dout(new_net_9424)
	);

	bfr new_net_9425_bfr_after (
		.din(new_net_9424),
		.dout(new_net_9425)
	);

	bfr new_net_9426_bfr_after (
		.din(new_net_9425),
		.dout(new_net_9426)
	);

	bfr new_net_9427_bfr_after (
		.din(new_net_9426),
		.dout(new_net_9427)
	);

	bfr new_net_9428_bfr_after (
		.din(new_net_9427),
		.dout(new_net_9428)
	);

	bfr new_net_9429_bfr_after (
		.din(new_net_9428),
		.dout(new_net_9429)
	);

	bfr new_net_9430_bfr_after (
		.din(new_net_9429),
		.dout(new_net_9430)
	);

	bfr new_net_9431_bfr_after (
		.din(new_net_9430),
		.dout(new_net_9431)
	);

	bfr new_net_9432_bfr_after (
		.din(new_net_9431),
		.dout(new_net_9432)
	);

	bfr new_net_9433_bfr_after (
		.din(new_net_9432),
		.dout(new_net_9433)
	);

	bfr new_net_9434_bfr_after (
		.din(new_net_9433),
		.dout(new_net_9434)
	);

	bfr new_net_9435_bfr_after (
		.din(new_net_9434),
		.dout(new_net_9435)
	);

	bfr new_net_9436_bfr_after (
		.din(new_net_9435),
		.dout(new_net_9436)
	);

	bfr new_net_9437_bfr_after (
		.din(new_net_9436),
		.dout(new_net_9437)
	);

	bfr new_net_9438_bfr_after (
		.din(new_net_9437),
		.dout(new_net_9438)
	);

	bfr new_net_9439_bfr_after (
		.din(new_net_9438),
		.dout(new_net_9439)
	);

	bfr new_net_9440_bfr_after (
		.din(new_net_9439),
		.dout(new_net_9440)
	);

	bfr new_net_9441_bfr_after (
		.din(new_net_9440),
		.dout(new_net_9441)
	);

	bfr new_net_9442_bfr_after (
		.din(new_net_9441),
		.dout(new_net_9442)
	);

	bfr new_net_9443_bfr_after (
		.din(new_net_9442),
		.dout(new_net_9443)
	);

	bfr new_net_9444_bfr_after (
		.din(new_net_9443),
		.dout(new_net_9444)
	);

	bfr new_net_9445_bfr_after (
		.din(new_net_9444),
		.dout(new_net_9445)
	);

	bfr new_net_9446_bfr_after (
		.din(new_net_9445),
		.dout(new_net_9446)
	);

	bfr new_net_9447_bfr_after (
		.din(new_net_9446),
		.dout(new_net_9447)
	);

	bfr new_net_9448_bfr_after (
		.din(new_net_9447),
		.dout(new_net_9448)
	);

	bfr new_net_9449_bfr_after (
		.din(new_net_9448),
		.dout(new_net_9449)
	);

	bfr new_net_9450_bfr_after (
		.din(new_net_9449),
		.dout(new_net_9450)
	);

	bfr new_net_9451_bfr_after (
		.din(new_net_9450),
		.dout(new_net_9451)
	);

	bfr new_net_9452_bfr_after (
		.din(new_net_9451),
		.dout(new_net_9452)
	);

	bfr new_net_9453_bfr_after (
		.din(new_net_9452),
		.dout(new_net_9453)
	);

	bfr new_net_9454_bfr_after (
		.din(new_net_9453),
		.dout(new_net_9454)
	);

	bfr new_net_9455_bfr_after (
		.din(new_net_9454),
		.dout(new_net_9455)
	);

	bfr new_net_9456_bfr_after (
		.din(new_net_9455),
		.dout(new_net_9456)
	);

	spl2 _0835__v_fanout (
		.a(new_net_9456),
		.b(new_net_2376),
		.c(new_net_2377)
	);

	bfr new_net_9457_bfr_after (
		.din(_1377_),
		.dout(new_net_9457)
	);

	bfr new_net_9458_bfr_after (
		.din(new_net_9457),
		.dout(new_net_9458)
	);

	bfr new_net_9459_bfr_after (
		.din(new_net_9458),
		.dout(new_net_9459)
	);

	bfr new_net_9460_bfr_after (
		.din(new_net_9459),
		.dout(new_net_9460)
	);

	bfr new_net_9461_bfr_after (
		.din(new_net_9460),
		.dout(new_net_9461)
	);

	bfr new_net_9462_bfr_after (
		.din(new_net_9461),
		.dout(new_net_9462)
	);

	bfr new_net_9463_bfr_after (
		.din(new_net_9462),
		.dout(new_net_9463)
	);

	bfr new_net_9464_bfr_after (
		.din(new_net_9463),
		.dout(new_net_9464)
	);

	bfr new_net_9465_bfr_after (
		.din(new_net_9464),
		.dout(new_net_9465)
	);

	bfr new_net_9466_bfr_after (
		.din(new_net_9465),
		.dout(new_net_9466)
	);

	bfr new_net_9467_bfr_after (
		.din(new_net_9466),
		.dout(new_net_9467)
	);

	bfr new_net_9468_bfr_after (
		.din(new_net_9467),
		.dout(new_net_9468)
	);

	bfr new_net_9469_bfr_after (
		.din(new_net_9468),
		.dout(new_net_9469)
	);

	bfr new_net_9470_bfr_after (
		.din(new_net_9469),
		.dout(new_net_9470)
	);

	bfr new_net_9471_bfr_after (
		.din(new_net_9470),
		.dout(new_net_9471)
	);

	bfr new_net_9472_bfr_after (
		.din(new_net_9471),
		.dout(new_net_9472)
	);

	bfr new_net_9473_bfr_after (
		.din(new_net_9472),
		.dout(new_net_9473)
	);

	bfr new_net_9474_bfr_after (
		.din(new_net_9473),
		.dout(new_net_9474)
	);

	bfr new_net_9475_bfr_after (
		.din(new_net_9474),
		.dout(new_net_9475)
	);

	bfr new_net_9476_bfr_after (
		.din(new_net_9475),
		.dout(new_net_9476)
	);

	bfr new_net_9477_bfr_after (
		.din(new_net_9476),
		.dout(new_net_9477)
	);

	bfr new_net_9478_bfr_after (
		.din(new_net_9477),
		.dout(new_net_9478)
	);

	bfr new_net_9479_bfr_after (
		.din(new_net_9478),
		.dout(new_net_9479)
	);

	bfr new_net_9480_bfr_after (
		.din(new_net_9479),
		.dout(new_net_9480)
	);

	spl2 _1377__v_fanout (
		.a(new_net_9480),
		.b(new_net_2825),
		.c(new_net_2826)
	);

	bfr new_net_9481_bfr_after (
		.din(_1030_),
		.dout(new_net_9481)
	);

	bfr new_net_9482_bfr_after (
		.din(new_net_9481),
		.dout(new_net_9482)
	);

	bfr new_net_9483_bfr_after (
		.din(new_net_9482),
		.dout(new_net_9483)
	);

	bfr new_net_9484_bfr_after (
		.din(new_net_9483),
		.dout(new_net_9484)
	);

	bfr new_net_9485_bfr_after (
		.din(new_net_9484),
		.dout(new_net_9485)
	);

	bfr new_net_9486_bfr_after (
		.din(new_net_9485),
		.dout(new_net_9486)
	);

	bfr new_net_9487_bfr_after (
		.din(new_net_9486),
		.dout(new_net_9487)
	);

	bfr new_net_9488_bfr_after (
		.din(new_net_9487),
		.dout(new_net_9488)
	);

	spl2 _1030__v_fanout (
		.a(new_net_9488),
		.b(new_net_303),
		.c(new_net_304)
	);

	bfr new_net_9489_bfr_after (
		.din(_0229_),
		.dout(new_net_9489)
	);

	bfr new_net_9490_bfr_after (
		.din(new_net_9489),
		.dout(new_net_9490)
	);

	bfr new_net_9491_bfr_after (
		.din(new_net_9490),
		.dout(new_net_9491)
	);

	bfr new_net_9492_bfr_after (
		.din(new_net_9491),
		.dout(new_net_9492)
	);

	bfr new_net_9493_bfr_after (
		.din(new_net_9492),
		.dout(new_net_9493)
	);

	bfr new_net_9494_bfr_after (
		.din(new_net_9493),
		.dout(new_net_9494)
	);

	bfr new_net_9495_bfr_after (
		.din(new_net_9494),
		.dout(new_net_9495)
	);

	bfr new_net_9496_bfr_after (
		.din(new_net_9495),
		.dout(new_net_9496)
	);

	bfr new_net_9497_bfr_after (
		.din(new_net_9496),
		.dout(new_net_9497)
	);

	bfr new_net_9498_bfr_after (
		.din(new_net_9497),
		.dout(new_net_9498)
	);

	bfr new_net_9499_bfr_after (
		.din(new_net_9498),
		.dout(new_net_9499)
	);

	bfr new_net_9500_bfr_after (
		.din(new_net_9499),
		.dout(new_net_9500)
	);

	bfr new_net_9501_bfr_after (
		.din(new_net_9500),
		.dout(new_net_9501)
	);

	bfr new_net_9502_bfr_after (
		.din(new_net_9501),
		.dout(new_net_9502)
	);

	bfr new_net_9503_bfr_after (
		.din(new_net_9502),
		.dout(new_net_9503)
	);

	bfr new_net_9504_bfr_after (
		.din(new_net_9503),
		.dout(new_net_9504)
	);

	bfr new_net_9505_bfr_after (
		.din(new_net_9504),
		.dout(new_net_9505)
	);

	bfr new_net_9506_bfr_after (
		.din(new_net_9505),
		.dout(new_net_9506)
	);

	bfr new_net_9507_bfr_after (
		.din(new_net_9506),
		.dout(new_net_9507)
	);

	bfr new_net_9508_bfr_after (
		.din(new_net_9507),
		.dout(new_net_9508)
	);

	bfr new_net_9509_bfr_after (
		.din(new_net_9508),
		.dout(new_net_9509)
	);

	bfr new_net_9510_bfr_after (
		.din(new_net_9509),
		.dout(new_net_9510)
	);

	bfr new_net_9511_bfr_after (
		.din(new_net_9510),
		.dout(new_net_9511)
	);

	bfr new_net_9512_bfr_after (
		.din(new_net_9511),
		.dout(new_net_9512)
	);

	bfr new_net_9513_bfr_after (
		.din(new_net_9512),
		.dout(new_net_9513)
	);

	bfr new_net_9514_bfr_after (
		.din(new_net_9513),
		.dout(new_net_9514)
	);

	bfr new_net_9515_bfr_after (
		.din(new_net_9514),
		.dout(new_net_9515)
	);

	bfr new_net_9516_bfr_after (
		.din(new_net_9515),
		.dout(new_net_9516)
	);

	bfr new_net_9517_bfr_after (
		.din(new_net_9516),
		.dout(new_net_9517)
	);

	bfr new_net_9518_bfr_after (
		.din(new_net_9517),
		.dout(new_net_9518)
	);

	bfr new_net_9519_bfr_after (
		.din(new_net_9518),
		.dout(new_net_9519)
	);

	bfr new_net_9520_bfr_after (
		.din(new_net_9519),
		.dout(new_net_9520)
	);

	bfr new_net_9521_bfr_after (
		.din(new_net_9520),
		.dout(new_net_9521)
	);

	bfr new_net_9522_bfr_after (
		.din(new_net_9521),
		.dout(new_net_9522)
	);

	bfr new_net_9523_bfr_after (
		.din(new_net_9522),
		.dout(new_net_9523)
	);

	bfr new_net_9524_bfr_after (
		.din(new_net_9523),
		.dout(new_net_9524)
	);

	bfr new_net_9525_bfr_after (
		.din(new_net_9524),
		.dout(new_net_9525)
	);

	bfr new_net_9526_bfr_after (
		.din(new_net_9525),
		.dout(new_net_9526)
	);

	bfr new_net_9527_bfr_after (
		.din(new_net_9526),
		.dout(new_net_9527)
	);

	bfr new_net_9528_bfr_after (
		.din(new_net_9527),
		.dout(new_net_9528)
	);

	bfr new_net_9529_bfr_after (
		.din(new_net_9528),
		.dout(new_net_9529)
	);

	bfr new_net_9530_bfr_after (
		.din(new_net_9529),
		.dout(new_net_9530)
	);

	bfr new_net_9531_bfr_after (
		.din(new_net_9530),
		.dout(new_net_9531)
	);

	bfr new_net_9532_bfr_after (
		.din(new_net_9531),
		.dout(new_net_9532)
	);

	bfr new_net_9533_bfr_after (
		.din(new_net_9532),
		.dout(new_net_9533)
	);

	bfr new_net_9534_bfr_after (
		.din(new_net_9533),
		.dout(new_net_9534)
	);

	bfr new_net_9535_bfr_after (
		.din(new_net_9534),
		.dout(new_net_9535)
	);

	bfr new_net_9536_bfr_after (
		.din(new_net_9535),
		.dout(new_net_9536)
	);

	spl2 _0229__v_fanout (
		.a(new_net_9536),
		.b(new_net_2214),
		.c(new_net_2215)
	);

	bfr new_net_9537_bfr_after (
		.din(_0452_),
		.dout(new_net_9537)
	);

	bfr new_net_9538_bfr_after (
		.din(new_net_9537),
		.dout(new_net_9538)
	);

	bfr new_net_9539_bfr_after (
		.din(new_net_9538),
		.dout(new_net_9539)
	);

	bfr new_net_9540_bfr_after (
		.din(new_net_9539),
		.dout(new_net_9540)
	);

	bfr new_net_9541_bfr_after (
		.din(new_net_9540),
		.dout(new_net_9541)
	);

	bfr new_net_9542_bfr_after (
		.din(new_net_9541),
		.dout(new_net_9542)
	);

	bfr new_net_9543_bfr_after (
		.din(new_net_9542),
		.dout(new_net_9543)
	);

	bfr new_net_9544_bfr_after (
		.din(new_net_9543),
		.dout(new_net_9544)
	);

	bfr new_net_9545_bfr_after (
		.din(new_net_9544),
		.dout(new_net_9545)
	);

	bfr new_net_9546_bfr_after (
		.din(new_net_9545),
		.dout(new_net_9546)
	);

	bfr new_net_9547_bfr_after (
		.din(new_net_9546),
		.dout(new_net_9547)
	);

	bfr new_net_9548_bfr_after (
		.din(new_net_9547),
		.dout(new_net_9548)
	);

	bfr new_net_9549_bfr_after (
		.din(new_net_9548),
		.dout(new_net_9549)
	);

	bfr new_net_9550_bfr_after (
		.din(new_net_9549),
		.dout(new_net_9550)
	);

	bfr new_net_9551_bfr_after (
		.din(new_net_9550),
		.dout(new_net_9551)
	);

	bfr new_net_9552_bfr_after (
		.din(new_net_9551),
		.dout(new_net_9552)
	);

	bfr new_net_9553_bfr_after (
		.din(new_net_9552),
		.dout(new_net_9553)
	);

	bfr new_net_9554_bfr_after (
		.din(new_net_9553),
		.dout(new_net_9554)
	);

	bfr new_net_9555_bfr_after (
		.din(new_net_9554),
		.dout(new_net_9555)
	);

	bfr new_net_9556_bfr_after (
		.din(new_net_9555),
		.dout(new_net_9556)
	);

	bfr new_net_9557_bfr_after (
		.din(new_net_9556),
		.dout(new_net_9557)
	);

	bfr new_net_9558_bfr_after (
		.din(new_net_9557),
		.dout(new_net_9558)
	);

	bfr new_net_9559_bfr_after (
		.din(new_net_9558),
		.dout(new_net_9559)
	);

	bfr new_net_9560_bfr_after (
		.din(new_net_9559),
		.dout(new_net_9560)
	);

	bfr new_net_9561_bfr_after (
		.din(new_net_9560),
		.dout(new_net_9561)
	);

	bfr new_net_9562_bfr_after (
		.din(new_net_9561),
		.dout(new_net_9562)
	);

	bfr new_net_9563_bfr_after (
		.din(new_net_9562),
		.dout(new_net_9563)
	);

	bfr new_net_9564_bfr_after (
		.din(new_net_9563),
		.dout(new_net_9564)
	);

	bfr new_net_9565_bfr_after (
		.din(new_net_9564),
		.dout(new_net_9565)
	);

	bfr new_net_9566_bfr_after (
		.din(new_net_9565),
		.dout(new_net_9566)
	);

	bfr new_net_9567_bfr_after (
		.din(new_net_9566),
		.dout(new_net_9567)
	);

	bfr new_net_9568_bfr_after (
		.din(new_net_9567),
		.dout(new_net_9568)
	);

	bfr new_net_9569_bfr_after (
		.din(new_net_9568),
		.dout(new_net_9569)
	);

	bfr new_net_9570_bfr_after (
		.din(new_net_9569),
		.dout(new_net_9570)
	);

	spl2 _0452__v_fanout (
		.a(new_net_9570),
		.b(new_net_184),
		.c(new_net_185)
	);

	bfr new_net_9571_bfr_after (
		.din(_0086_),
		.dout(new_net_9571)
	);

	bfr new_net_9572_bfr_after (
		.din(new_net_9571),
		.dout(new_net_9572)
	);

	bfr new_net_9573_bfr_after (
		.din(new_net_9572),
		.dout(new_net_9573)
	);

	bfr new_net_9574_bfr_after (
		.din(new_net_9573),
		.dout(new_net_9574)
	);

	bfr new_net_9575_bfr_after (
		.din(new_net_9574),
		.dout(new_net_9575)
	);

	bfr new_net_9576_bfr_after (
		.din(new_net_9575),
		.dout(new_net_9576)
	);

	bfr new_net_9577_bfr_after (
		.din(new_net_9576),
		.dout(new_net_9577)
	);

	bfr new_net_9578_bfr_after (
		.din(new_net_9577),
		.dout(new_net_9578)
	);

	bfr new_net_9579_bfr_after (
		.din(new_net_9578),
		.dout(new_net_9579)
	);

	bfr new_net_9580_bfr_after (
		.din(new_net_9579),
		.dout(new_net_9580)
	);

	bfr new_net_9581_bfr_after (
		.din(new_net_9580),
		.dout(new_net_9581)
	);

	bfr new_net_9582_bfr_after (
		.din(new_net_9581),
		.dout(new_net_9582)
	);

	bfr new_net_9583_bfr_after (
		.din(new_net_9582),
		.dout(new_net_9583)
	);

	bfr new_net_9584_bfr_after (
		.din(new_net_9583),
		.dout(new_net_9584)
	);

	bfr new_net_9585_bfr_after (
		.din(new_net_9584),
		.dout(new_net_9585)
	);

	bfr new_net_9586_bfr_after (
		.din(new_net_9585),
		.dout(new_net_9586)
	);

	bfr new_net_9587_bfr_after (
		.din(new_net_9586),
		.dout(new_net_9587)
	);

	bfr new_net_9588_bfr_after (
		.din(new_net_9587),
		.dout(new_net_9588)
	);

	bfr new_net_9589_bfr_after (
		.din(new_net_9588),
		.dout(new_net_9589)
	);

	bfr new_net_9590_bfr_after (
		.din(new_net_9589),
		.dout(new_net_9590)
	);

	bfr new_net_9591_bfr_after (
		.din(new_net_9590),
		.dout(new_net_9591)
	);

	bfr new_net_9592_bfr_after (
		.din(new_net_9591),
		.dout(new_net_9592)
	);

	bfr new_net_9593_bfr_after (
		.din(new_net_9592),
		.dout(new_net_9593)
	);

	bfr new_net_9594_bfr_after (
		.din(new_net_9593),
		.dout(new_net_9594)
	);

	bfr new_net_9595_bfr_after (
		.din(new_net_9594),
		.dout(new_net_9595)
	);

	bfr new_net_9596_bfr_after (
		.din(new_net_9595),
		.dout(new_net_9596)
	);

	bfr new_net_9597_bfr_after (
		.din(new_net_9596),
		.dout(new_net_9597)
	);

	bfr new_net_9598_bfr_after (
		.din(new_net_9597),
		.dout(new_net_9598)
	);

	bfr new_net_9599_bfr_after (
		.din(new_net_9598),
		.dout(new_net_9599)
	);

	bfr new_net_9600_bfr_after (
		.din(new_net_9599),
		.dout(new_net_9600)
	);

	bfr new_net_9601_bfr_after (
		.din(new_net_9600),
		.dout(new_net_9601)
	);

	bfr new_net_9602_bfr_after (
		.din(new_net_9601),
		.dout(new_net_9602)
	);

	bfr new_net_9603_bfr_after (
		.din(new_net_9602),
		.dout(new_net_9603)
	);

	bfr new_net_9604_bfr_after (
		.din(new_net_9603),
		.dout(new_net_9604)
	);

	bfr new_net_9605_bfr_after (
		.din(new_net_9604),
		.dout(new_net_9605)
	);

	bfr new_net_9606_bfr_after (
		.din(new_net_9605),
		.dout(new_net_9606)
	);

	bfr new_net_9607_bfr_after (
		.din(new_net_9606),
		.dout(new_net_9607)
	);

	bfr new_net_9608_bfr_after (
		.din(new_net_9607),
		.dout(new_net_9608)
	);

	bfr new_net_9609_bfr_after (
		.din(new_net_9608),
		.dout(new_net_9609)
	);

	bfr new_net_9610_bfr_after (
		.din(new_net_9609),
		.dout(new_net_9610)
	);

	bfr new_net_9611_bfr_after (
		.din(new_net_9610),
		.dout(new_net_9611)
	);

	bfr new_net_9612_bfr_after (
		.din(new_net_9611),
		.dout(new_net_9612)
	);

	bfr new_net_9613_bfr_after (
		.din(new_net_9612),
		.dout(new_net_9613)
	);

	bfr new_net_9614_bfr_after (
		.din(new_net_9613),
		.dout(new_net_9614)
	);

	bfr new_net_9615_bfr_after (
		.din(new_net_9614),
		.dout(new_net_9615)
	);

	bfr new_net_9616_bfr_after (
		.din(new_net_9615),
		.dout(new_net_9616)
	);

	bfr new_net_9617_bfr_after (
		.din(new_net_9616),
		.dout(new_net_9617)
	);

	bfr new_net_9618_bfr_after (
		.din(new_net_9617),
		.dout(new_net_9618)
	);

	bfr new_net_9619_bfr_after (
		.din(new_net_9618),
		.dout(new_net_9619)
	);

	bfr new_net_9620_bfr_after (
		.din(new_net_9619),
		.dout(new_net_9620)
	);

	bfr new_net_9621_bfr_after (
		.din(new_net_9620),
		.dout(new_net_9621)
	);

	bfr new_net_9622_bfr_after (
		.din(new_net_9621),
		.dout(new_net_9622)
	);

	bfr new_net_9623_bfr_after (
		.din(new_net_9622),
		.dout(new_net_9623)
	);

	bfr new_net_9624_bfr_after (
		.din(new_net_9623),
		.dout(new_net_9624)
	);

	bfr new_net_9625_bfr_after (
		.din(new_net_9624),
		.dout(new_net_9625)
	);

	bfr new_net_9626_bfr_after (
		.din(new_net_9625),
		.dout(new_net_9626)
	);

	bfr new_net_9627_bfr_after (
		.din(new_net_9626),
		.dout(new_net_9627)
	);

	bfr new_net_9628_bfr_after (
		.din(new_net_9627),
		.dout(new_net_9628)
	);

	bfr new_net_9629_bfr_after (
		.din(new_net_9628),
		.dout(new_net_9629)
	);

	bfr new_net_9630_bfr_after (
		.din(new_net_9629),
		.dout(new_net_9630)
	);

	bfr new_net_9631_bfr_after (
		.din(new_net_9630),
		.dout(new_net_9631)
	);

	bfr new_net_9632_bfr_after (
		.din(new_net_9631),
		.dout(new_net_9632)
	);

	bfr new_net_9633_bfr_after (
		.din(new_net_9632),
		.dout(new_net_9633)
	);

	bfr new_net_9634_bfr_after (
		.din(new_net_9633),
		.dout(new_net_9634)
	);

	bfr new_net_9635_bfr_after (
		.din(new_net_9634),
		.dout(new_net_9635)
	);

	bfr new_net_9636_bfr_after (
		.din(new_net_9635),
		.dout(new_net_9636)
	);

	bfr new_net_9637_bfr_after (
		.din(new_net_9636),
		.dout(new_net_9637)
	);

	bfr new_net_9638_bfr_after (
		.din(new_net_9637),
		.dout(new_net_9638)
	);

	bfr new_net_9639_bfr_after (
		.din(new_net_9638),
		.dout(new_net_9639)
	);

	bfr new_net_9640_bfr_after (
		.din(new_net_9639),
		.dout(new_net_9640)
	);

	bfr new_net_9641_bfr_after (
		.din(new_net_9640),
		.dout(new_net_9641)
	);

	bfr new_net_9642_bfr_after (
		.din(new_net_9641),
		.dout(new_net_9642)
	);

	bfr new_net_9643_bfr_after (
		.din(new_net_9642),
		.dout(new_net_9643)
	);

	bfr new_net_9644_bfr_after (
		.din(new_net_9643),
		.dout(new_net_9644)
	);

	bfr new_net_9645_bfr_after (
		.din(new_net_9644),
		.dout(new_net_9645)
	);

	bfr new_net_9646_bfr_after (
		.din(new_net_9645),
		.dout(new_net_9646)
	);

	bfr new_net_9647_bfr_after (
		.din(new_net_9646),
		.dout(new_net_9647)
	);

	bfr new_net_9648_bfr_after (
		.din(new_net_9647),
		.dout(new_net_9648)
	);

	bfr new_net_9649_bfr_after (
		.din(new_net_9648),
		.dout(new_net_9649)
	);

	bfr new_net_9650_bfr_after (
		.din(new_net_9649),
		.dout(new_net_9650)
	);

	bfr new_net_9651_bfr_after (
		.din(new_net_9650),
		.dout(new_net_9651)
	);

	bfr new_net_9652_bfr_after (
		.din(new_net_9651),
		.dout(new_net_9652)
	);

	bfr new_net_9653_bfr_after (
		.din(new_net_9652),
		.dout(new_net_9653)
	);

	bfr new_net_9654_bfr_after (
		.din(new_net_9653),
		.dout(new_net_9654)
	);

	bfr new_net_9655_bfr_after (
		.din(new_net_9654),
		.dout(new_net_9655)
	);

	bfr new_net_9656_bfr_after (
		.din(new_net_9655),
		.dout(new_net_9656)
	);

	bfr new_net_9657_bfr_after (
		.din(new_net_9656),
		.dout(new_net_9657)
	);

	bfr new_net_9658_bfr_after (
		.din(new_net_9657),
		.dout(new_net_9658)
	);

	bfr new_net_9659_bfr_after (
		.din(new_net_9658),
		.dout(new_net_9659)
	);

	bfr new_net_9660_bfr_after (
		.din(new_net_9659),
		.dout(new_net_9660)
	);

	bfr new_net_9661_bfr_after (
		.din(new_net_9660),
		.dout(new_net_9661)
	);

	bfr new_net_9662_bfr_after (
		.din(new_net_9661),
		.dout(new_net_9662)
	);

	bfr new_net_9663_bfr_after (
		.din(new_net_9662),
		.dout(new_net_9663)
	);

	bfr new_net_9664_bfr_after (
		.din(new_net_9663),
		.dout(new_net_9664)
	);

	bfr new_net_9665_bfr_after (
		.din(new_net_9664),
		.dout(new_net_9665)
	);

	bfr new_net_9666_bfr_after (
		.din(new_net_9665),
		.dout(new_net_9666)
	);

	bfr new_net_9667_bfr_after (
		.din(new_net_9666),
		.dout(new_net_9667)
	);

	bfr new_net_9668_bfr_after (
		.din(new_net_9667),
		.dout(new_net_9668)
	);

	bfr new_net_9669_bfr_after (
		.din(new_net_9668),
		.dout(new_net_9669)
	);

	bfr new_net_9670_bfr_after (
		.din(new_net_9669),
		.dout(new_net_9670)
	);

	bfr new_net_9671_bfr_after (
		.din(new_net_9670),
		.dout(new_net_9671)
	);

	bfr new_net_9672_bfr_after (
		.din(new_net_9671),
		.dout(new_net_9672)
	);

	bfr new_net_9673_bfr_after (
		.din(new_net_9672),
		.dout(new_net_9673)
	);

	bfr new_net_9674_bfr_after (
		.din(new_net_9673),
		.dout(new_net_9674)
	);

	spl2 _0086__v_fanout (
		.a(new_net_9674),
		.b(new_net_2180),
		.c(new_net_2181)
	);

	bfr new_net_9675_bfr_after (
		.din(_1578_),
		.dout(new_net_9675)
	);

	bfr new_net_9676_bfr_after (
		.din(new_net_9675),
		.dout(new_net_9676)
	);

	bfr new_net_9677_bfr_after (
		.din(new_net_9676),
		.dout(new_net_9677)
	);

	bfr new_net_9678_bfr_after (
		.din(new_net_9677),
		.dout(new_net_9678)
	);

	bfr new_net_9679_bfr_after (
		.din(new_net_9678),
		.dout(new_net_9679)
	);

	bfr new_net_9680_bfr_after (
		.din(new_net_9679),
		.dout(new_net_9680)
	);

	bfr new_net_9681_bfr_after (
		.din(new_net_9680),
		.dout(new_net_9681)
	);

	bfr new_net_9682_bfr_after (
		.din(new_net_9681),
		.dout(new_net_9682)
	);

	bfr new_net_9683_bfr_after (
		.din(new_net_9682),
		.dout(new_net_9683)
	);

	bfr new_net_9684_bfr_after (
		.din(new_net_9683),
		.dout(new_net_9684)
	);

	bfr new_net_9685_bfr_after (
		.din(new_net_9684),
		.dout(new_net_9685)
	);

	bfr new_net_9686_bfr_after (
		.din(new_net_9685),
		.dout(new_net_9686)
	);

	bfr new_net_9687_bfr_after (
		.din(new_net_9686),
		.dout(new_net_9687)
	);

	bfr new_net_9688_bfr_after (
		.din(new_net_9687),
		.dout(new_net_9688)
	);

	bfr new_net_9689_bfr_after (
		.din(new_net_9688),
		.dout(new_net_9689)
	);

	bfr new_net_9690_bfr_after (
		.din(new_net_9689),
		.dout(new_net_9690)
	);

	bfr new_net_9691_bfr_after (
		.din(new_net_9690),
		.dout(new_net_9691)
	);

	bfr new_net_9692_bfr_after (
		.din(new_net_9691),
		.dout(new_net_9692)
	);

	bfr new_net_9693_bfr_after (
		.din(new_net_9692),
		.dout(new_net_9693)
	);

	bfr new_net_9694_bfr_after (
		.din(new_net_9693),
		.dout(new_net_9694)
	);

	bfr new_net_9695_bfr_after (
		.din(new_net_9694),
		.dout(new_net_9695)
	);

	bfr new_net_9696_bfr_after (
		.din(new_net_9695),
		.dout(new_net_9696)
	);

	bfr new_net_9697_bfr_after (
		.din(new_net_9696),
		.dout(new_net_9697)
	);

	bfr new_net_9698_bfr_after (
		.din(new_net_9697),
		.dout(new_net_9698)
	);

	bfr new_net_9699_bfr_after (
		.din(new_net_9698),
		.dout(new_net_9699)
	);

	bfr new_net_9700_bfr_after (
		.din(new_net_9699),
		.dout(new_net_9700)
	);

	bfr new_net_9701_bfr_after (
		.din(new_net_9700),
		.dout(new_net_9701)
	);

	bfr new_net_9702_bfr_after (
		.din(new_net_9701),
		.dout(new_net_9702)
	);

	bfr new_net_9703_bfr_after (
		.din(new_net_9702),
		.dout(new_net_9703)
	);

	bfr new_net_9704_bfr_after (
		.din(new_net_9703),
		.dout(new_net_9704)
	);

	bfr new_net_9705_bfr_after (
		.din(new_net_9704),
		.dout(new_net_9705)
	);

	bfr new_net_9706_bfr_after (
		.din(new_net_9705),
		.dout(new_net_9706)
	);

	bfr new_net_9707_bfr_after (
		.din(new_net_9706),
		.dout(new_net_9707)
	);

	bfr new_net_9708_bfr_after (
		.din(new_net_9707),
		.dout(new_net_9708)
	);

	bfr new_net_9709_bfr_after (
		.din(new_net_9708),
		.dout(new_net_9709)
	);

	bfr new_net_9710_bfr_after (
		.din(new_net_9709),
		.dout(new_net_9710)
	);

	bfr new_net_9711_bfr_after (
		.din(new_net_9710),
		.dout(new_net_9711)
	);

	bfr new_net_9712_bfr_after (
		.din(new_net_9711),
		.dout(new_net_9712)
	);

	bfr new_net_9713_bfr_after (
		.din(new_net_9712),
		.dout(new_net_9713)
	);

	bfr new_net_9714_bfr_after (
		.din(new_net_9713),
		.dout(new_net_9714)
	);

	spl2 _1578__v_fanout (
		.a(new_net_9714),
		.b(new_net_1948),
		.c(new_net_1949)
	);

	bfr new_net_9715_bfr_after (
		.din(_0930_),
		.dout(new_net_9715)
	);

	bfr new_net_9716_bfr_after (
		.din(new_net_9715),
		.dout(new_net_9716)
	);

	bfr new_net_9717_bfr_after (
		.din(new_net_9716),
		.dout(new_net_9717)
	);

	bfr new_net_9718_bfr_after (
		.din(new_net_9717),
		.dout(new_net_9718)
	);

	bfr new_net_9719_bfr_after (
		.din(new_net_9718),
		.dout(new_net_9719)
	);

	bfr new_net_9720_bfr_after (
		.din(new_net_9719),
		.dout(new_net_9720)
	);

	bfr new_net_9721_bfr_after (
		.din(new_net_9720),
		.dout(new_net_9721)
	);

	bfr new_net_9722_bfr_after (
		.din(new_net_9721),
		.dout(new_net_9722)
	);

	bfr new_net_9723_bfr_after (
		.din(new_net_9722),
		.dout(new_net_9723)
	);

	bfr new_net_9724_bfr_after (
		.din(new_net_9723),
		.dout(new_net_9724)
	);

	bfr new_net_9725_bfr_after (
		.din(new_net_9724),
		.dout(new_net_9725)
	);

	bfr new_net_9726_bfr_after (
		.din(new_net_9725),
		.dout(new_net_9726)
	);

	bfr new_net_9727_bfr_after (
		.din(new_net_9726),
		.dout(new_net_9727)
	);

	bfr new_net_9728_bfr_after (
		.din(new_net_9727),
		.dout(new_net_9728)
	);

	bfr new_net_9729_bfr_after (
		.din(new_net_9728),
		.dout(new_net_9729)
	);

	bfr new_net_9730_bfr_after (
		.din(new_net_9729),
		.dout(new_net_9730)
	);

	bfr new_net_9731_bfr_after (
		.din(new_net_9730),
		.dout(new_net_9731)
	);

	bfr new_net_9732_bfr_after (
		.din(new_net_9731),
		.dout(new_net_9732)
	);

	bfr new_net_9733_bfr_after (
		.din(new_net_9732),
		.dout(new_net_9733)
	);

	bfr new_net_9734_bfr_after (
		.din(new_net_9733),
		.dout(new_net_9734)
	);

	bfr new_net_9735_bfr_after (
		.din(new_net_9734),
		.dout(new_net_9735)
	);

	bfr new_net_9736_bfr_after (
		.din(new_net_9735),
		.dout(new_net_9736)
	);

	bfr new_net_9737_bfr_after (
		.din(new_net_9736),
		.dout(new_net_9737)
	);

	bfr new_net_9738_bfr_after (
		.din(new_net_9737),
		.dout(new_net_9738)
	);

	bfr new_net_9739_bfr_after (
		.din(new_net_9738),
		.dout(new_net_9739)
	);

	bfr new_net_9740_bfr_after (
		.din(new_net_9739),
		.dout(new_net_9740)
	);

	bfr new_net_9741_bfr_after (
		.din(new_net_9740),
		.dout(new_net_9741)
	);

	bfr new_net_9742_bfr_after (
		.din(new_net_9741),
		.dout(new_net_9742)
	);

	bfr new_net_9743_bfr_after (
		.din(new_net_9742),
		.dout(new_net_9743)
	);

	bfr new_net_9744_bfr_after (
		.din(new_net_9743),
		.dout(new_net_9744)
	);

	bfr new_net_9745_bfr_after (
		.din(new_net_9744),
		.dout(new_net_9745)
	);

	bfr new_net_9746_bfr_after (
		.din(new_net_9745),
		.dout(new_net_9746)
	);

	bfr new_net_9747_bfr_after (
		.din(new_net_9746),
		.dout(new_net_9747)
	);

	bfr new_net_9748_bfr_after (
		.din(new_net_9747),
		.dout(new_net_9748)
	);

	bfr new_net_9749_bfr_after (
		.din(new_net_9748),
		.dout(new_net_9749)
	);

	bfr new_net_9750_bfr_after (
		.din(new_net_9749),
		.dout(new_net_9750)
	);

	bfr new_net_9751_bfr_after (
		.din(new_net_9750),
		.dout(new_net_9751)
	);

	bfr new_net_9752_bfr_after (
		.din(new_net_9751),
		.dout(new_net_9752)
	);

	bfr new_net_9753_bfr_after (
		.din(new_net_9752),
		.dout(new_net_9753)
	);

	bfr new_net_9754_bfr_after (
		.din(new_net_9753),
		.dout(new_net_9754)
	);

	bfr new_net_9755_bfr_after (
		.din(new_net_9754),
		.dout(new_net_9755)
	);

	bfr new_net_9756_bfr_after (
		.din(new_net_9755),
		.dout(new_net_9756)
	);

	bfr new_net_9757_bfr_after (
		.din(new_net_9756),
		.dout(new_net_9757)
	);

	bfr new_net_9758_bfr_after (
		.din(new_net_9757),
		.dout(new_net_9758)
	);

	bfr new_net_9759_bfr_after (
		.din(new_net_9758),
		.dout(new_net_9759)
	);

	bfr new_net_9760_bfr_after (
		.din(new_net_9759),
		.dout(new_net_9760)
	);

	bfr new_net_9761_bfr_after (
		.din(new_net_9760),
		.dout(new_net_9761)
	);

	bfr new_net_9762_bfr_after (
		.din(new_net_9761),
		.dout(new_net_9762)
	);

	bfr new_net_9763_bfr_after (
		.din(new_net_9762),
		.dout(new_net_9763)
	);

	bfr new_net_9764_bfr_after (
		.din(new_net_9763),
		.dout(new_net_9764)
	);

	bfr new_net_9765_bfr_after (
		.din(new_net_9764),
		.dout(new_net_9765)
	);

	bfr new_net_9766_bfr_after (
		.din(new_net_9765),
		.dout(new_net_9766)
	);

	bfr new_net_9767_bfr_after (
		.din(new_net_9766),
		.dout(new_net_9767)
	);

	bfr new_net_9768_bfr_after (
		.din(new_net_9767),
		.dout(new_net_9768)
	);

	bfr new_net_9769_bfr_after (
		.din(new_net_9768),
		.dout(new_net_9769)
	);

	bfr new_net_9770_bfr_after (
		.din(new_net_9769),
		.dout(new_net_9770)
	);

	bfr new_net_9771_bfr_after (
		.din(new_net_9770),
		.dout(new_net_9771)
	);

	bfr new_net_9772_bfr_after (
		.din(new_net_9771),
		.dout(new_net_9772)
	);

	bfr new_net_9773_bfr_after (
		.din(new_net_9772),
		.dout(new_net_9773)
	);

	bfr new_net_9774_bfr_after (
		.din(new_net_9773),
		.dout(new_net_9774)
	);

	bfr new_net_9775_bfr_after (
		.din(new_net_9774),
		.dout(new_net_9775)
	);

	bfr new_net_9776_bfr_after (
		.din(new_net_9775),
		.dout(new_net_9776)
	);

	bfr new_net_9777_bfr_after (
		.din(new_net_9776),
		.dout(new_net_9777)
	);

	bfr new_net_9778_bfr_after (
		.din(new_net_9777),
		.dout(new_net_9778)
	);

	bfr new_net_9779_bfr_after (
		.din(new_net_9778),
		.dout(new_net_9779)
	);

	bfr new_net_9780_bfr_after (
		.din(new_net_9779),
		.dout(new_net_9780)
	);

	bfr new_net_9781_bfr_after (
		.din(new_net_9780),
		.dout(new_net_9781)
	);

	bfr new_net_9782_bfr_after (
		.din(new_net_9781),
		.dout(new_net_9782)
	);

	bfr new_net_9783_bfr_after (
		.din(new_net_9782),
		.dout(new_net_9783)
	);

	bfr new_net_9784_bfr_after (
		.din(new_net_9783),
		.dout(new_net_9784)
	);

	bfr new_net_9785_bfr_after (
		.din(new_net_9784),
		.dout(new_net_9785)
	);

	bfr new_net_9786_bfr_after (
		.din(new_net_9785),
		.dout(new_net_9786)
	);

	bfr new_net_9787_bfr_after (
		.din(new_net_9786),
		.dout(new_net_9787)
	);

	bfr new_net_9788_bfr_after (
		.din(new_net_9787),
		.dout(new_net_9788)
	);

	bfr new_net_9789_bfr_after (
		.din(new_net_9788),
		.dout(new_net_9789)
	);

	bfr new_net_9790_bfr_after (
		.din(new_net_9789),
		.dout(new_net_9790)
	);

	bfr new_net_9791_bfr_after (
		.din(new_net_9790),
		.dout(new_net_9791)
	);

	bfr new_net_9792_bfr_after (
		.din(new_net_9791),
		.dout(new_net_9792)
	);

	bfr new_net_9793_bfr_after (
		.din(new_net_9792),
		.dout(new_net_9793)
	);

	bfr new_net_9794_bfr_after (
		.din(new_net_9793),
		.dout(new_net_9794)
	);

	bfr new_net_9795_bfr_after (
		.din(new_net_9794),
		.dout(new_net_9795)
	);

	bfr new_net_9796_bfr_after (
		.din(new_net_9795),
		.dout(new_net_9796)
	);

	bfr new_net_9797_bfr_after (
		.din(new_net_9796),
		.dout(new_net_9797)
	);

	bfr new_net_9798_bfr_after (
		.din(new_net_9797),
		.dout(new_net_9798)
	);

	bfr new_net_9799_bfr_after (
		.din(new_net_9798),
		.dout(new_net_9799)
	);

	bfr new_net_9800_bfr_after (
		.din(new_net_9799),
		.dout(new_net_9800)
	);

	bfr new_net_9801_bfr_after (
		.din(new_net_9800),
		.dout(new_net_9801)
	);

	bfr new_net_9802_bfr_after (
		.din(new_net_9801),
		.dout(new_net_9802)
	);

	bfr new_net_9803_bfr_after (
		.din(new_net_9802),
		.dout(new_net_9803)
	);

	bfr new_net_9804_bfr_after (
		.din(new_net_9803),
		.dout(new_net_9804)
	);

	spl2 _0930__v_fanout (
		.a(new_net_9804),
		.b(new_net_1291),
		.c(new_net_1292)
	);

	bfr new_net_9805_bfr_after (
		.din(_0617_),
		.dout(new_net_9805)
	);

	bfr new_net_9806_bfr_after (
		.din(new_net_9805),
		.dout(new_net_9806)
	);

	bfr new_net_9807_bfr_after (
		.din(new_net_9806),
		.dout(new_net_9807)
	);

	bfr new_net_9808_bfr_after (
		.din(new_net_9807),
		.dout(new_net_9808)
	);

	bfr new_net_9809_bfr_after (
		.din(new_net_9808),
		.dout(new_net_9809)
	);

	bfr new_net_9810_bfr_after (
		.din(new_net_9809),
		.dout(new_net_9810)
	);

	bfr new_net_9811_bfr_after (
		.din(new_net_9810),
		.dout(new_net_9811)
	);

	bfr new_net_9812_bfr_after (
		.din(new_net_9811),
		.dout(new_net_9812)
	);

	bfr new_net_9813_bfr_after (
		.din(new_net_9812),
		.dout(new_net_9813)
	);

	bfr new_net_9814_bfr_after (
		.din(new_net_9813),
		.dout(new_net_9814)
	);

	bfr new_net_9815_bfr_after (
		.din(new_net_9814),
		.dout(new_net_9815)
	);

	bfr new_net_9816_bfr_after (
		.din(new_net_9815),
		.dout(new_net_9816)
	);

	bfr new_net_9817_bfr_after (
		.din(new_net_9816),
		.dout(new_net_9817)
	);

	bfr new_net_9818_bfr_after (
		.din(new_net_9817),
		.dout(new_net_9818)
	);

	bfr new_net_9819_bfr_after (
		.din(new_net_9818),
		.dout(new_net_9819)
	);

	bfr new_net_9820_bfr_after (
		.din(new_net_9819),
		.dout(new_net_9820)
	);

	bfr new_net_9821_bfr_after (
		.din(new_net_9820),
		.dout(new_net_9821)
	);

	bfr new_net_9822_bfr_after (
		.din(new_net_9821),
		.dout(new_net_9822)
	);

	bfr new_net_9823_bfr_after (
		.din(new_net_9822),
		.dout(new_net_9823)
	);

	bfr new_net_9824_bfr_after (
		.din(new_net_9823),
		.dout(new_net_9824)
	);

	bfr new_net_9825_bfr_after (
		.din(new_net_9824),
		.dout(new_net_9825)
	);

	bfr new_net_9826_bfr_after (
		.din(new_net_9825),
		.dout(new_net_9826)
	);

	bfr new_net_9827_bfr_after (
		.din(new_net_9826),
		.dout(new_net_9827)
	);

	bfr new_net_9828_bfr_after (
		.din(new_net_9827),
		.dout(new_net_9828)
	);

	bfr new_net_9829_bfr_after (
		.din(new_net_9828),
		.dout(new_net_9829)
	);

	bfr new_net_9830_bfr_after (
		.din(new_net_9829),
		.dout(new_net_9830)
	);

	bfr new_net_9831_bfr_after (
		.din(new_net_9830),
		.dout(new_net_9831)
	);

	bfr new_net_9832_bfr_after (
		.din(new_net_9831),
		.dout(new_net_9832)
	);

	bfr new_net_9833_bfr_after (
		.din(new_net_9832),
		.dout(new_net_9833)
	);

	bfr new_net_9834_bfr_after (
		.din(new_net_9833),
		.dout(new_net_9834)
	);

	bfr new_net_9835_bfr_after (
		.din(new_net_9834),
		.dout(new_net_9835)
	);

	bfr new_net_9836_bfr_after (
		.din(new_net_9835),
		.dout(new_net_9836)
	);

	bfr new_net_9837_bfr_after (
		.din(new_net_9836),
		.dout(new_net_9837)
	);

	bfr new_net_9838_bfr_after (
		.din(new_net_9837),
		.dout(new_net_9838)
	);

	bfr new_net_9839_bfr_after (
		.din(new_net_9838),
		.dout(new_net_9839)
	);

	bfr new_net_9840_bfr_after (
		.din(new_net_9839),
		.dout(new_net_9840)
	);

	bfr new_net_9841_bfr_after (
		.din(new_net_9840),
		.dout(new_net_9841)
	);

	bfr new_net_9842_bfr_after (
		.din(new_net_9841),
		.dout(new_net_9842)
	);

	bfr new_net_9843_bfr_after (
		.din(new_net_9842),
		.dout(new_net_9843)
	);

	bfr new_net_9844_bfr_after (
		.din(new_net_9843),
		.dout(new_net_9844)
	);

	bfr new_net_9845_bfr_after (
		.din(new_net_9844),
		.dout(new_net_9845)
	);

	bfr new_net_9846_bfr_after (
		.din(new_net_9845),
		.dout(new_net_9846)
	);

	bfr new_net_9847_bfr_after (
		.din(new_net_9846),
		.dout(new_net_9847)
	);

	bfr new_net_9848_bfr_after (
		.din(new_net_9847),
		.dout(new_net_9848)
	);

	bfr new_net_9849_bfr_after (
		.din(new_net_9848),
		.dout(new_net_9849)
	);

	bfr new_net_9850_bfr_after (
		.din(new_net_9849),
		.dout(new_net_9850)
	);

	bfr new_net_9851_bfr_after (
		.din(new_net_9850),
		.dout(new_net_9851)
	);

	bfr new_net_9852_bfr_after (
		.din(new_net_9851),
		.dout(new_net_9852)
	);

	bfr new_net_9853_bfr_after (
		.din(new_net_9852),
		.dout(new_net_9853)
	);

	bfr new_net_9854_bfr_after (
		.din(new_net_9853),
		.dout(new_net_9854)
	);

	bfr new_net_9855_bfr_after (
		.din(new_net_9854),
		.dout(new_net_9855)
	);

	bfr new_net_9856_bfr_after (
		.din(new_net_9855),
		.dout(new_net_9856)
	);

	bfr new_net_9857_bfr_after (
		.din(new_net_9856),
		.dout(new_net_9857)
	);

	bfr new_net_9858_bfr_after (
		.din(new_net_9857),
		.dout(new_net_9858)
	);

	bfr new_net_9859_bfr_after (
		.din(new_net_9858),
		.dout(new_net_9859)
	);

	bfr new_net_9860_bfr_after (
		.din(new_net_9859),
		.dout(new_net_9860)
	);

	bfr new_net_9861_bfr_after (
		.din(new_net_9860),
		.dout(new_net_9861)
	);

	bfr new_net_9862_bfr_after (
		.din(new_net_9861),
		.dout(new_net_9862)
	);

	bfr new_net_9863_bfr_after (
		.din(new_net_9862),
		.dout(new_net_9863)
	);

	bfr new_net_9864_bfr_after (
		.din(new_net_9863),
		.dout(new_net_9864)
	);

	bfr new_net_9865_bfr_after (
		.din(new_net_9864),
		.dout(new_net_9865)
	);

	bfr new_net_9866_bfr_after (
		.din(new_net_9865),
		.dout(new_net_9866)
	);

	bfr new_net_9867_bfr_after (
		.din(new_net_9866),
		.dout(new_net_9867)
	);

	bfr new_net_9868_bfr_after (
		.din(new_net_9867),
		.dout(new_net_9868)
	);

	bfr new_net_9869_bfr_after (
		.din(new_net_9868),
		.dout(new_net_9869)
	);

	bfr new_net_9870_bfr_after (
		.din(new_net_9869),
		.dout(new_net_9870)
	);

	bfr new_net_9871_bfr_after (
		.din(new_net_9870),
		.dout(new_net_9871)
	);

	bfr new_net_9872_bfr_after (
		.din(new_net_9871),
		.dout(new_net_9872)
	);

	bfr new_net_9873_bfr_after (
		.din(new_net_9872),
		.dout(new_net_9873)
	);

	bfr new_net_9874_bfr_after (
		.din(new_net_9873),
		.dout(new_net_9874)
	);

	bfr new_net_9875_bfr_after (
		.din(new_net_9874),
		.dout(new_net_9875)
	);

	bfr new_net_9876_bfr_after (
		.din(new_net_9875),
		.dout(new_net_9876)
	);

	bfr new_net_9877_bfr_after (
		.din(new_net_9876),
		.dout(new_net_9877)
	);

	bfr new_net_9878_bfr_after (
		.din(new_net_9877),
		.dout(new_net_9878)
	);

	bfr new_net_9879_bfr_after (
		.din(new_net_9878),
		.dout(new_net_9879)
	);

	bfr new_net_9880_bfr_after (
		.din(new_net_9879),
		.dout(new_net_9880)
	);

	bfr new_net_9881_bfr_after (
		.din(new_net_9880),
		.dout(new_net_9881)
	);

	bfr new_net_9882_bfr_after (
		.din(new_net_9881),
		.dout(new_net_9882)
	);

	bfr new_net_9883_bfr_after (
		.din(new_net_9882),
		.dout(new_net_9883)
	);

	bfr new_net_9884_bfr_after (
		.din(new_net_9883),
		.dout(new_net_9884)
	);

	bfr new_net_9885_bfr_after (
		.din(new_net_9884),
		.dout(new_net_9885)
	);

	bfr new_net_9886_bfr_after (
		.din(new_net_9885),
		.dout(new_net_9886)
	);

	bfr new_net_9887_bfr_after (
		.din(new_net_9886),
		.dout(new_net_9887)
	);

	bfr new_net_9888_bfr_after (
		.din(new_net_9887),
		.dout(new_net_9888)
	);

	bfr new_net_9889_bfr_after (
		.din(new_net_9888),
		.dout(new_net_9889)
	);

	bfr new_net_9890_bfr_after (
		.din(new_net_9889),
		.dout(new_net_9890)
	);

	bfr new_net_9891_bfr_after (
		.din(new_net_9890),
		.dout(new_net_9891)
	);

	bfr new_net_9892_bfr_after (
		.din(new_net_9891),
		.dout(new_net_9892)
	);

	bfr new_net_9893_bfr_after (
		.din(new_net_9892),
		.dout(new_net_9893)
	);

	bfr new_net_9894_bfr_after (
		.din(new_net_9893),
		.dout(new_net_9894)
	);

	bfr new_net_9895_bfr_after (
		.din(new_net_9894),
		.dout(new_net_9895)
	);

	bfr new_net_9896_bfr_after (
		.din(new_net_9895),
		.dout(new_net_9896)
	);

	bfr new_net_9897_bfr_after (
		.din(new_net_9896),
		.dout(new_net_9897)
	);

	bfr new_net_9898_bfr_after (
		.din(new_net_9897),
		.dout(new_net_9898)
	);

	bfr new_net_9899_bfr_after (
		.din(new_net_9898),
		.dout(new_net_9899)
	);

	bfr new_net_9900_bfr_after (
		.din(new_net_9899),
		.dout(new_net_9900)
	);

	bfr new_net_9901_bfr_after (
		.din(new_net_9900),
		.dout(new_net_9901)
	);

	bfr new_net_9902_bfr_after (
		.din(new_net_9901),
		.dout(new_net_9902)
	);

	bfr new_net_9903_bfr_after (
		.din(new_net_9902),
		.dout(new_net_9903)
	);

	bfr new_net_9904_bfr_after (
		.din(new_net_9903),
		.dout(new_net_9904)
	);

	bfr new_net_9905_bfr_after (
		.din(new_net_9904),
		.dout(new_net_9905)
	);

	bfr new_net_9906_bfr_after (
		.din(new_net_9905),
		.dout(new_net_9906)
	);

	bfr new_net_9907_bfr_after (
		.din(new_net_9906),
		.dout(new_net_9907)
	);

	bfr new_net_9908_bfr_after (
		.din(new_net_9907),
		.dout(new_net_9908)
	);

	bfr new_net_9909_bfr_after (
		.din(new_net_9908),
		.dout(new_net_9909)
	);

	bfr new_net_9910_bfr_after (
		.din(new_net_9909),
		.dout(new_net_9910)
	);

	bfr new_net_9911_bfr_after (
		.din(new_net_9910),
		.dout(new_net_9911)
	);

	bfr new_net_9912_bfr_after (
		.din(new_net_9911),
		.dout(new_net_9912)
	);

	bfr new_net_9913_bfr_after (
		.din(new_net_9912),
		.dout(new_net_9913)
	);

	bfr new_net_9914_bfr_after (
		.din(new_net_9913),
		.dout(new_net_9914)
	);

	bfr new_net_9915_bfr_after (
		.din(new_net_9914),
		.dout(new_net_9915)
	);

	bfr new_net_9916_bfr_after (
		.din(new_net_9915),
		.dout(new_net_9916)
	);

	spl2 _0617__v_fanout (
		.a(new_net_9916),
		.b(new_net_2284),
		.c(new_net_2285)
	);

	bfr new_net_9917_bfr_after (
		.din(_1476_),
		.dout(new_net_9917)
	);

	bfr new_net_9918_bfr_after (
		.din(new_net_9917),
		.dout(new_net_9918)
	);

	bfr new_net_9919_bfr_after (
		.din(new_net_9918),
		.dout(new_net_9919)
	);

	bfr new_net_9920_bfr_after (
		.din(new_net_9919),
		.dout(new_net_9920)
	);

	bfr new_net_9921_bfr_after (
		.din(new_net_9920),
		.dout(new_net_9921)
	);

	bfr new_net_9922_bfr_after (
		.din(new_net_9921),
		.dout(new_net_9922)
	);

	bfr new_net_9923_bfr_after (
		.din(new_net_9922),
		.dout(new_net_9923)
	);

	bfr new_net_9924_bfr_after (
		.din(new_net_9923),
		.dout(new_net_9924)
	);

	spl2 _1476__v_fanout (
		.a(new_net_9924),
		.b(new_net_1279),
		.c(new_net_1280)
	);

	spl2 _1222__v_fanout (
		.a(_1222_),
		.b(new_net_1174),
		.c(new_net_1175)
	);

	bfr new_net_9925_bfr_after (
		.din(_1825_),
		.dout(new_net_9925)
	);

	bfr new_net_9926_bfr_after (
		.din(new_net_9925),
		.dout(new_net_9926)
	);

	bfr new_net_9927_bfr_after (
		.din(new_net_9926),
		.dout(new_net_9927)
	);

	bfr new_net_9928_bfr_after (
		.din(new_net_9927),
		.dout(new_net_9928)
	);

	bfr new_net_9929_bfr_after (
		.din(new_net_9928),
		.dout(new_net_9929)
	);

	bfr new_net_9930_bfr_after (
		.din(new_net_9929),
		.dout(new_net_9930)
	);

	bfr new_net_9931_bfr_after (
		.din(new_net_9930),
		.dout(new_net_9931)
	);

	bfr new_net_9932_bfr_after (
		.din(new_net_9931),
		.dout(new_net_9932)
	);

	bfr new_net_9933_bfr_after (
		.din(new_net_9932),
		.dout(new_net_9933)
	);

	bfr new_net_9934_bfr_after (
		.din(new_net_9933),
		.dout(new_net_9934)
	);

	bfr new_net_9935_bfr_after (
		.din(new_net_9934),
		.dout(new_net_9935)
	);

	bfr new_net_9936_bfr_after (
		.din(new_net_9935),
		.dout(new_net_9936)
	);

	bfr new_net_9937_bfr_after (
		.din(new_net_9936),
		.dout(new_net_9937)
	);

	bfr new_net_9938_bfr_after (
		.din(new_net_9937),
		.dout(new_net_9938)
	);

	bfr new_net_9939_bfr_after (
		.din(new_net_9938),
		.dout(new_net_9939)
	);

	bfr new_net_9940_bfr_after (
		.din(new_net_9939),
		.dout(new_net_9940)
	);

	bfr new_net_9941_bfr_after (
		.din(new_net_9940),
		.dout(new_net_9941)
	);

	bfr new_net_9942_bfr_after (
		.din(new_net_9941),
		.dout(new_net_9942)
	);

	bfr new_net_9943_bfr_after (
		.din(new_net_9942),
		.dout(new_net_9943)
	);

	bfr new_net_9944_bfr_after (
		.din(new_net_9943),
		.dout(new_net_9944)
	);

	bfr new_net_9945_bfr_after (
		.din(new_net_9944),
		.dout(new_net_9945)
	);

	bfr new_net_9946_bfr_after (
		.din(new_net_9945),
		.dout(new_net_9946)
	);

	bfr new_net_9947_bfr_after (
		.din(new_net_9946),
		.dout(new_net_9947)
	);

	bfr new_net_9948_bfr_after (
		.din(new_net_9947),
		.dout(new_net_9948)
	);

	spl2 _1825__v_fanout (
		.a(new_net_9948),
		.b(new_net_1762),
		.c(new_net_1763)
	);

	bfr new_net_9949_bfr_after (
		.din(_1804_),
		.dout(new_net_9949)
	);

	bfr new_net_9950_bfr_after (
		.din(new_net_9949),
		.dout(new_net_9950)
	);

	bfr new_net_9951_bfr_after (
		.din(new_net_9950),
		.dout(new_net_9951)
	);

	bfr new_net_9952_bfr_after (
		.din(new_net_9951),
		.dout(new_net_9952)
	);

	bfr new_net_9953_bfr_after (
		.din(new_net_9952),
		.dout(new_net_9953)
	);

	bfr new_net_9954_bfr_after (
		.din(new_net_9953),
		.dout(new_net_9954)
	);

	bfr new_net_9955_bfr_after (
		.din(new_net_9954),
		.dout(new_net_9955)
	);

	bfr new_net_9956_bfr_after (
		.din(new_net_9955),
		.dout(new_net_9956)
	);

	bfr new_net_9957_bfr_after (
		.din(new_net_9956),
		.dout(new_net_9957)
	);

	bfr new_net_9958_bfr_after (
		.din(new_net_9957),
		.dout(new_net_9958)
	);

	bfr new_net_9959_bfr_after (
		.din(new_net_9958),
		.dout(new_net_9959)
	);

	bfr new_net_9960_bfr_after (
		.din(new_net_9959),
		.dout(new_net_9960)
	);

	bfr new_net_9961_bfr_after (
		.din(new_net_9960),
		.dout(new_net_9961)
	);

	bfr new_net_9962_bfr_after (
		.din(new_net_9961),
		.dout(new_net_9962)
	);

	bfr new_net_9963_bfr_after (
		.din(new_net_9962),
		.dout(new_net_9963)
	);

	bfr new_net_9964_bfr_after (
		.din(new_net_9963),
		.dout(new_net_9964)
	);

	bfr new_net_9965_bfr_after (
		.din(new_net_9964),
		.dout(new_net_9965)
	);

	bfr new_net_9966_bfr_after (
		.din(new_net_9965),
		.dout(new_net_9966)
	);

	bfr new_net_9967_bfr_after (
		.din(new_net_9966),
		.dout(new_net_9967)
	);

	bfr new_net_9968_bfr_after (
		.din(new_net_9967),
		.dout(new_net_9968)
	);

	bfr new_net_9969_bfr_after (
		.din(new_net_9968),
		.dout(new_net_9969)
	);

	bfr new_net_9970_bfr_after (
		.din(new_net_9969),
		.dout(new_net_9970)
	);

	bfr new_net_9971_bfr_after (
		.din(new_net_9970),
		.dout(new_net_9971)
	);

	bfr new_net_9972_bfr_after (
		.din(new_net_9971),
		.dout(new_net_9972)
	);

	bfr new_net_9973_bfr_after (
		.din(new_net_9972),
		.dout(new_net_9973)
	);

	bfr new_net_9974_bfr_after (
		.din(new_net_9973),
		.dout(new_net_9974)
	);

	bfr new_net_9975_bfr_after (
		.din(new_net_9974),
		.dout(new_net_9975)
	);

	bfr new_net_9976_bfr_after (
		.din(new_net_9975),
		.dout(new_net_9976)
	);

	bfr new_net_9977_bfr_after (
		.din(new_net_9976),
		.dout(new_net_9977)
	);

	bfr new_net_9978_bfr_after (
		.din(new_net_9977),
		.dout(new_net_9978)
	);

	bfr new_net_9979_bfr_after (
		.din(new_net_9978),
		.dout(new_net_9979)
	);

	bfr new_net_9980_bfr_after (
		.din(new_net_9979),
		.dout(new_net_9980)
	);

	bfr new_net_9981_bfr_after (
		.din(new_net_9980),
		.dout(new_net_9981)
	);

	bfr new_net_9982_bfr_after (
		.din(new_net_9981),
		.dout(new_net_9982)
	);

	bfr new_net_9983_bfr_after (
		.din(new_net_9982),
		.dout(new_net_9983)
	);

	bfr new_net_9984_bfr_after (
		.din(new_net_9983),
		.dout(new_net_9984)
	);

	bfr new_net_9985_bfr_after (
		.din(new_net_9984),
		.dout(new_net_9985)
	);

	bfr new_net_9986_bfr_after (
		.din(new_net_9985),
		.dout(new_net_9986)
	);

	bfr new_net_9987_bfr_after (
		.din(new_net_9986),
		.dout(new_net_9987)
	);

	bfr new_net_9988_bfr_after (
		.din(new_net_9987),
		.dout(new_net_9988)
	);

	bfr new_net_9989_bfr_after (
		.din(new_net_9988),
		.dout(new_net_9989)
	);

	bfr new_net_9990_bfr_after (
		.din(new_net_9989),
		.dout(new_net_9990)
	);

	bfr new_net_9991_bfr_after (
		.din(new_net_9990),
		.dout(new_net_9991)
	);

	bfr new_net_9992_bfr_after (
		.din(new_net_9991),
		.dout(new_net_9992)
	);

	bfr new_net_9993_bfr_after (
		.din(new_net_9992),
		.dout(new_net_9993)
	);

	bfr new_net_9994_bfr_after (
		.din(new_net_9993),
		.dout(new_net_9994)
	);

	bfr new_net_9995_bfr_after (
		.din(new_net_9994),
		.dout(new_net_9995)
	);

	bfr new_net_9996_bfr_after (
		.din(new_net_9995),
		.dout(new_net_9996)
	);

	bfr new_net_9997_bfr_after (
		.din(new_net_9996),
		.dout(new_net_9997)
	);

	bfr new_net_9998_bfr_after (
		.din(new_net_9997),
		.dout(new_net_9998)
	);

	bfr new_net_9999_bfr_after (
		.din(new_net_9998),
		.dout(new_net_9999)
	);

	bfr new_net_10000_bfr_after (
		.din(new_net_9999),
		.dout(new_net_10000)
	);

	bfr new_net_10001_bfr_after (
		.din(new_net_10000),
		.dout(new_net_10001)
	);

	bfr new_net_10002_bfr_after (
		.din(new_net_10001),
		.dout(new_net_10002)
	);

	bfr new_net_10003_bfr_after (
		.din(new_net_10002),
		.dout(new_net_10003)
	);

	bfr new_net_10004_bfr_after (
		.din(new_net_10003),
		.dout(new_net_10004)
	);

	bfr new_net_10005_bfr_after (
		.din(new_net_10004),
		.dout(new_net_10005)
	);

	bfr new_net_10006_bfr_after (
		.din(new_net_10005),
		.dout(new_net_10006)
	);

	bfr new_net_10007_bfr_after (
		.din(new_net_10006),
		.dout(new_net_10007)
	);

	bfr new_net_10008_bfr_after (
		.din(new_net_10007),
		.dout(new_net_10008)
	);

	bfr new_net_10009_bfr_after (
		.din(new_net_10008),
		.dout(new_net_10009)
	);

	bfr new_net_10010_bfr_after (
		.din(new_net_10009),
		.dout(new_net_10010)
	);

	bfr new_net_10011_bfr_after (
		.din(new_net_10010),
		.dout(new_net_10011)
	);

	bfr new_net_10012_bfr_after (
		.din(new_net_10011),
		.dout(new_net_10012)
	);

	bfr new_net_10013_bfr_after (
		.din(new_net_10012),
		.dout(new_net_10013)
	);

	bfr new_net_10014_bfr_after (
		.din(new_net_10013),
		.dout(new_net_10014)
	);

	bfr new_net_10015_bfr_after (
		.din(new_net_10014),
		.dout(new_net_10015)
	);

	bfr new_net_10016_bfr_after (
		.din(new_net_10015),
		.dout(new_net_10016)
	);

	bfr new_net_10017_bfr_after (
		.din(new_net_10016),
		.dout(new_net_10017)
	);

	bfr new_net_10018_bfr_after (
		.din(new_net_10017),
		.dout(new_net_10018)
	);

	bfr new_net_10019_bfr_after (
		.din(new_net_10018),
		.dout(new_net_10019)
	);

	bfr new_net_10020_bfr_after (
		.din(new_net_10019),
		.dout(new_net_10020)
	);

	bfr new_net_10021_bfr_after (
		.din(new_net_10020),
		.dout(new_net_10021)
	);

	bfr new_net_10022_bfr_after (
		.din(new_net_10021),
		.dout(new_net_10022)
	);

	bfr new_net_10023_bfr_after (
		.din(new_net_10022),
		.dout(new_net_10023)
	);

	bfr new_net_10024_bfr_after (
		.din(new_net_10023),
		.dout(new_net_10024)
	);

	bfr new_net_10025_bfr_after (
		.din(new_net_10024),
		.dout(new_net_10025)
	);

	bfr new_net_10026_bfr_after (
		.din(new_net_10025),
		.dout(new_net_10026)
	);

	bfr new_net_10027_bfr_after (
		.din(new_net_10026),
		.dout(new_net_10027)
	);

	bfr new_net_10028_bfr_after (
		.din(new_net_10027),
		.dout(new_net_10028)
	);

	bfr new_net_10029_bfr_after (
		.din(new_net_10028),
		.dout(new_net_10029)
	);

	bfr new_net_10030_bfr_after (
		.din(new_net_10029),
		.dout(new_net_10030)
	);

	bfr new_net_10031_bfr_after (
		.din(new_net_10030),
		.dout(new_net_10031)
	);

	bfr new_net_10032_bfr_after (
		.din(new_net_10031),
		.dout(new_net_10032)
	);

	bfr new_net_10033_bfr_after (
		.din(new_net_10032),
		.dout(new_net_10033)
	);

	bfr new_net_10034_bfr_after (
		.din(new_net_10033),
		.dout(new_net_10034)
	);

	bfr new_net_10035_bfr_after (
		.din(new_net_10034),
		.dout(new_net_10035)
	);

	bfr new_net_10036_bfr_after (
		.din(new_net_10035),
		.dout(new_net_10036)
	);

	bfr new_net_10037_bfr_after (
		.din(new_net_10036),
		.dout(new_net_10037)
	);

	bfr new_net_10038_bfr_after (
		.din(new_net_10037),
		.dout(new_net_10038)
	);

	bfr new_net_10039_bfr_after (
		.din(new_net_10038),
		.dout(new_net_10039)
	);

	bfr new_net_10040_bfr_after (
		.din(new_net_10039),
		.dout(new_net_10040)
	);

	bfr new_net_10041_bfr_after (
		.din(new_net_10040),
		.dout(new_net_10041)
	);

	bfr new_net_10042_bfr_after (
		.din(new_net_10041),
		.dout(new_net_10042)
	);

	bfr new_net_10043_bfr_after (
		.din(new_net_10042),
		.dout(new_net_10043)
	);

	bfr new_net_10044_bfr_after (
		.din(new_net_10043),
		.dout(new_net_10044)
	);

	bfr new_net_10045_bfr_after (
		.din(new_net_10044),
		.dout(new_net_10045)
	);

	bfr new_net_10046_bfr_after (
		.din(new_net_10045),
		.dout(new_net_10046)
	);

	bfr new_net_10047_bfr_after (
		.din(new_net_10046),
		.dout(new_net_10047)
	);

	bfr new_net_10048_bfr_after (
		.din(new_net_10047),
		.dout(new_net_10048)
	);

	bfr new_net_10049_bfr_after (
		.din(new_net_10048),
		.dout(new_net_10049)
	);

	bfr new_net_10050_bfr_after (
		.din(new_net_10049),
		.dout(new_net_10050)
	);

	bfr new_net_10051_bfr_after (
		.din(new_net_10050),
		.dout(new_net_10051)
	);

	bfr new_net_10052_bfr_after (
		.din(new_net_10051),
		.dout(new_net_10052)
	);

	spl2 _1804__v_fanout (
		.a(new_net_10052),
		.b(new_net_2058),
		.c(new_net_2059)
	);

	spl2 _1083__v_fanout (
		.a(_1083_),
		.b(new_net_2206),
		.c(new_net_2207)
	);

	bfr new_net_10053_bfr_after (
		.din(_1463_),
		.dout(new_net_10053)
	);

	bfr new_net_10054_bfr_after (
		.din(new_net_10053),
		.dout(new_net_10054)
	);

	bfr new_net_10055_bfr_after (
		.din(new_net_10054),
		.dout(new_net_10055)
	);

	bfr new_net_10056_bfr_after (
		.din(new_net_10055),
		.dout(new_net_10056)
	);

	bfr new_net_10057_bfr_after (
		.din(new_net_10056),
		.dout(new_net_10057)
	);

	bfr new_net_10058_bfr_after (
		.din(new_net_10057),
		.dout(new_net_10058)
	);

	bfr new_net_10059_bfr_after (
		.din(new_net_10058),
		.dout(new_net_10059)
	);

	bfr new_net_10060_bfr_after (
		.din(new_net_10059),
		.dout(new_net_10060)
	);

	bfr new_net_10061_bfr_after (
		.din(new_net_10060),
		.dout(new_net_10061)
	);

	bfr new_net_10062_bfr_after (
		.din(new_net_10061),
		.dout(new_net_10062)
	);

	bfr new_net_10063_bfr_after (
		.din(new_net_10062),
		.dout(new_net_10063)
	);

	bfr new_net_10064_bfr_after (
		.din(new_net_10063),
		.dout(new_net_10064)
	);

	bfr new_net_10065_bfr_after (
		.din(new_net_10064),
		.dout(new_net_10065)
	);

	bfr new_net_10066_bfr_after (
		.din(new_net_10065),
		.dout(new_net_10066)
	);

	bfr new_net_10067_bfr_after (
		.din(new_net_10066),
		.dout(new_net_10067)
	);

	bfr new_net_10068_bfr_after (
		.din(new_net_10067),
		.dout(new_net_10068)
	);

	bfr new_net_10069_bfr_after (
		.din(new_net_10068),
		.dout(new_net_10069)
	);

	bfr new_net_10070_bfr_after (
		.din(new_net_10069),
		.dout(new_net_10070)
	);

	bfr new_net_10071_bfr_after (
		.din(new_net_10070),
		.dout(new_net_10071)
	);

	bfr new_net_10072_bfr_after (
		.din(new_net_10071),
		.dout(new_net_10072)
	);

	bfr new_net_10073_bfr_after (
		.din(new_net_10072),
		.dout(new_net_10073)
	);

	bfr new_net_10074_bfr_after (
		.din(new_net_10073),
		.dout(new_net_10074)
	);

	bfr new_net_10075_bfr_after (
		.din(new_net_10074),
		.dout(new_net_10075)
	);

	bfr new_net_10076_bfr_after (
		.din(new_net_10075),
		.dout(new_net_10076)
	);

	bfr new_net_10077_bfr_after (
		.din(new_net_10076),
		.dout(new_net_10077)
	);

	bfr new_net_10078_bfr_after (
		.din(new_net_10077),
		.dout(new_net_10078)
	);

	bfr new_net_10079_bfr_after (
		.din(new_net_10078),
		.dout(new_net_10079)
	);

	bfr new_net_10080_bfr_after (
		.din(new_net_10079),
		.dout(new_net_10080)
	);

	bfr new_net_10081_bfr_after (
		.din(new_net_10080),
		.dout(new_net_10081)
	);

	bfr new_net_10082_bfr_after (
		.din(new_net_10081),
		.dout(new_net_10082)
	);

	bfr new_net_10083_bfr_after (
		.din(new_net_10082),
		.dout(new_net_10083)
	);

	bfr new_net_10084_bfr_after (
		.din(new_net_10083),
		.dout(new_net_10084)
	);

	bfr new_net_10085_bfr_after (
		.din(new_net_10084),
		.dout(new_net_10085)
	);

	bfr new_net_10086_bfr_after (
		.din(new_net_10085),
		.dout(new_net_10086)
	);

	bfr new_net_10087_bfr_after (
		.din(new_net_10086),
		.dout(new_net_10087)
	);

	bfr new_net_10088_bfr_after (
		.din(new_net_10087),
		.dout(new_net_10088)
	);

	bfr new_net_10089_bfr_after (
		.din(new_net_10088),
		.dout(new_net_10089)
	);

	bfr new_net_10090_bfr_after (
		.din(new_net_10089),
		.dout(new_net_10090)
	);

	bfr new_net_10091_bfr_after (
		.din(new_net_10090),
		.dout(new_net_10091)
	);

	bfr new_net_10092_bfr_after (
		.din(new_net_10091),
		.dout(new_net_10092)
	);

	bfr new_net_10093_bfr_after (
		.din(new_net_10092),
		.dout(new_net_10093)
	);

	bfr new_net_10094_bfr_after (
		.din(new_net_10093),
		.dout(new_net_10094)
	);

	bfr new_net_10095_bfr_after (
		.din(new_net_10094),
		.dout(new_net_10095)
	);

	bfr new_net_10096_bfr_after (
		.din(new_net_10095),
		.dout(new_net_10096)
	);

	bfr new_net_10097_bfr_after (
		.din(new_net_10096),
		.dout(new_net_10097)
	);

	bfr new_net_10098_bfr_after (
		.din(new_net_10097),
		.dout(new_net_10098)
	);

	bfr new_net_10099_bfr_after (
		.din(new_net_10098),
		.dout(new_net_10099)
	);

	bfr new_net_10100_bfr_after (
		.din(new_net_10099),
		.dout(new_net_10100)
	);

	bfr new_net_10101_bfr_after (
		.din(new_net_10100),
		.dout(new_net_10101)
	);

	bfr new_net_10102_bfr_after (
		.din(new_net_10101),
		.dout(new_net_10102)
	);

	bfr new_net_10103_bfr_after (
		.din(new_net_10102),
		.dout(new_net_10103)
	);

	bfr new_net_10104_bfr_after (
		.din(new_net_10103),
		.dout(new_net_10104)
	);

	bfr new_net_10105_bfr_after (
		.din(new_net_10104),
		.dout(new_net_10105)
	);

	bfr new_net_10106_bfr_after (
		.din(new_net_10105),
		.dout(new_net_10106)
	);

	bfr new_net_10107_bfr_after (
		.din(new_net_10106),
		.dout(new_net_10107)
	);

	bfr new_net_10108_bfr_after (
		.din(new_net_10107),
		.dout(new_net_10108)
	);

	spl2 _1463__v_fanout (
		.a(new_net_10108),
		.b(new_net_339),
		.c(new_net_340)
	);

	bfr new_net_10109_bfr_after (
		.din(_0619_),
		.dout(new_net_10109)
	);

	bfr new_net_10110_bfr_after (
		.din(new_net_10109),
		.dout(new_net_10110)
	);

	bfr new_net_10111_bfr_after (
		.din(new_net_10110),
		.dout(new_net_10111)
	);

	bfr new_net_10112_bfr_after (
		.din(new_net_10111),
		.dout(new_net_10112)
	);

	bfr new_net_10113_bfr_after (
		.din(new_net_10112),
		.dout(new_net_10113)
	);

	bfr new_net_10114_bfr_after (
		.din(new_net_10113),
		.dout(new_net_10114)
	);

	bfr new_net_10115_bfr_after (
		.din(new_net_10114),
		.dout(new_net_10115)
	);

	bfr new_net_10116_bfr_after (
		.din(new_net_10115),
		.dout(new_net_10116)
	);

	bfr new_net_10117_bfr_after (
		.din(new_net_10116),
		.dout(new_net_10117)
	);

	bfr new_net_10118_bfr_after (
		.din(new_net_10117),
		.dout(new_net_10118)
	);

	bfr new_net_10119_bfr_after (
		.din(new_net_10118),
		.dout(new_net_10119)
	);

	bfr new_net_10120_bfr_after (
		.din(new_net_10119),
		.dout(new_net_10120)
	);

	bfr new_net_10121_bfr_after (
		.din(new_net_10120),
		.dout(new_net_10121)
	);

	bfr new_net_10122_bfr_after (
		.din(new_net_10121),
		.dout(new_net_10122)
	);

	bfr new_net_10123_bfr_after (
		.din(new_net_10122),
		.dout(new_net_10123)
	);

	bfr new_net_10124_bfr_after (
		.din(new_net_10123),
		.dout(new_net_10124)
	);

	bfr new_net_10125_bfr_after (
		.din(new_net_10124),
		.dout(new_net_10125)
	);

	bfr new_net_10126_bfr_after (
		.din(new_net_10125),
		.dout(new_net_10126)
	);

	bfr new_net_10127_bfr_after (
		.din(new_net_10126),
		.dout(new_net_10127)
	);

	bfr new_net_10128_bfr_after (
		.din(new_net_10127),
		.dout(new_net_10128)
	);

	bfr new_net_10129_bfr_after (
		.din(new_net_10128),
		.dout(new_net_10129)
	);

	bfr new_net_10130_bfr_after (
		.din(new_net_10129),
		.dout(new_net_10130)
	);

	bfr new_net_10131_bfr_after (
		.din(new_net_10130),
		.dout(new_net_10131)
	);

	bfr new_net_10132_bfr_after (
		.din(new_net_10131),
		.dout(new_net_10132)
	);

	bfr new_net_10133_bfr_after (
		.din(new_net_10132),
		.dout(new_net_10133)
	);

	bfr new_net_10134_bfr_after (
		.din(new_net_10133),
		.dout(new_net_10134)
	);

	bfr new_net_10135_bfr_after (
		.din(new_net_10134),
		.dout(new_net_10135)
	);

	bfr new_net_10136_bfr_after (
		.din(new_net_10135),
		.dout(new_net_10136)
	);

	bfr new_net_10137_bfr_after (
		.din(new_net_10136),
		.dout(new_net_10137)
	);

	bfr new_net_10138_bfr_after (
		.din(new_net_10137),
		.dout(new_net_10138)
	);

	bfr new_net_10139_bfr_after (
		.din(new_net_10138),
		.dout(new_net_10139)
	);

	bfr new_net_10140_bfr_after (
		.din(new_net_10139),
		.dout(new_net_10140)
	);

	bfr new_net_10141_bfr_after (
		.din(new_net_10140),
		.dout(new_net_10141)
	);

	bfr new_net_10142_bfr_after (
		.din(new_net_10141),
		.dout(new_net_10142)
	);

	bfr new_net_10143_bfr_after (
		.din(new_net_10142),
		.dout(new_net_10143)
	);

	bfr new_net_10144_bfr_after (
		.din(new_net_10143),
		.dout(new_net_10144)
	);

	bfr new_net_10145_bfr_after (
		.din(new_net_10144),
		.dout(new_net_10145)
	);

	bfr new_net_10146_bfr_after (
		.din(new_net_10145),
		.dout(new_net_10146)
	);

	bfr new_net_10147_bfr_after (
		.din(new_net_10146),
		.dout(new_net_10147)
	);

	bfr new_net_10148_bfr_after (
		.din(new_net_10147),
		.dout(new_net_10148)
	);

	bfr new_net_10149_bfr_after (
		.din(new_net_10148),
		.dout(new_net_10149)
	);

	bfr new_net_10150_bfr_after (
		.din(new_net_10149),
		.dout(new_net_10150)
	);

	bfr new_net_10151_bfr_after (
		.din(new_net_10150),
		.dout(new_net_10151)
	);

	bfr new_net_10152_bfr_after (
		.din(new_net_10151),
		.dout(new_net_10152)
	);

	bfr new_net_10153_bfr_after (
		.din(new_net_10152),
		.dout(new_net_10153)
	);

	bfr new_net_10154_bfr_after (
		.din(new_net_10153),
		.dout(new_net_10154)
	);

	bfr new_net_10155_bfr_after (
		.din(new_net_10154),
		.dout(new_net_10155)
	);

	bfr new_net_10156_bfr_after (
		.din(new_net_10155),
		.dout(new_net_10156)
	);

	bfr new_net_10157_bfr_after (
		.din(new_net_10156),
		.dout(new_net_10157)
	);

	bfr new_net_10158_bfr_after (
		.din(new_net_10157),
		.dout(new_net_10158)
	);

	bfr new_net_10159_bfr_after (
		.din(new_net_10158),
		.dout(new_net_10159)
	);

	bfr new_net_10160_bfr_after (
		.din(new_net_10159),
		.dout(new_net_10160)
	);

	bfr new_net_10161_bfr_after (
		.din(new_net_10160),
		.dout(new_net_10161)
	);

	bfr new_net_10162_bfr_after (
		.din(new_net_10161),
		.dout(new_net_10162)
	);

	bfr new_net_10163_bfr_after (
		.din(new_net_10162),
		.dout(new_net_10163)
	);

	bfr new_net_10164_bfr_after (
		.din(new_net_10163),
		.dout(new_net_10164)
	);

	bfr new_net_10165_bfr_after (
		.din(new_net_10164),
		.dout(new_net_10165)
	);

	bfr new_net_10166_bfr_after (
		.din(new_net_10165),
		.dout(new_net_10166)
	);

	bfr new_net_10167_bfr_after (
		.din(new_net_10166),
		.dout(new_net_10167)
	);

	bfr new_net_10168_bfr_after (
		.din(new_net_10167),
		.dout(new_net_10168)
	);

	bfr new_net_10169_bfr_after (
		.din(new_net_10168),
		.dout(new_net_10169)
	);

	bfr new_net_10170_bfr_after (
		.din(new_net_10169),
		.dout(new_net_10170)
	);

	bfr new_net_10171_bfr_after (
		.din(new_net_10170),
		.dout(new_net_10171)
	);

	bfr new_net_10172_bfr_after (
		.din(new_net_10171),
		.dout(new_net_10172)
	);

	bfr new_net_10173_bfr_after (
		.din(new_net_10172),
		.dout(new_net_10173)
	);

	bfr new_net_10174_bfr_after (
		.din(new_net_10173),
		.dout(new_net_10174)
	);

	bfr new_net_10175_bfr_after (
		.din(new_net_10174),
		.dout(new_net_10175)
	);

	bfr new_net_10176_bfr_after (
		.din(new_net_10175),
		.dout(new_net_10176)
	);

	bfr new_net_10177_bfr_after (
		.din(new_net_10176),
		.dout(new_net_10177)
	);

	bfr new_net_10178_bfr_after (
		.din(new_net_10177),
		.dout(new_net_10178)
	);

	bfr new_net_10179_bfr_after (
		.din(new_net_10178),
		.dout(new_net_10179)
	);

	bfr new_net_10180_bfr_after (
		.din(new_net_10179),
		.dout(new_net_10180)
	);

	bfr new_net_10181_bfr_after (
		.din(new_net_10180),
		.dout(new_net_10181)
	);

	bfr new_net_10182_bfr_after (
		.din(new_net_10181),
		.dout(new_net_10182)
	);

	bfr new_net_10183_bfr_after (
		.din(new_net_10182),
		.dout(new_net_10183)
	);

	bfr new_net_10184_bfr_after (
		.din(new_net_10183),
		.dout(new_net_10184)
	);

	bfr new_net_10185_bfr_after (
		.din(new_net_10184),
		.dout(new_net_10185)
	);

	bfr new_net_10186_bfr_after (
		.din(new_net_10185),
		.dout(new_net_10186)
	);

	bfr new_net_10187_bfr_after (
		.din(new_net_10186),
		.dout(new_net_10187)
	);

	bfr new_net_10188_bfr_after (
		.din(new_net_10187),
		.dout(new_net_10188)
	);

	bfr new_net_10189_bfr_after (
		.din(new_net_10188),
		.dout(new_net_10189)
	);

	bfr new_net_10190_bfr_after (
		.din(new_net_10189),
		.dout(new_net_10190)
	);

	bfr new_net_10191_bfr_after (
		.din(new_net_10190),
		.dout(new_net_10191)
	);

	bfr new_net_10192_bfr_after (
		.din(new_net_10191),
		.dout(new_net_10192)
	);

	bfr new_net_10193_bfr_after (
		.din(new_net_10192),
		.dout(new_net_10193)
	);

	bfr new_net_10194_bfr_after (
		.din(new_net_10193),
		.dout(new_net_10194)
	);

	bfr new_net_10195_bfr_after (
		.din(new_net_10194),
		.dout(new_net_10195)
	);

	bfr new_net_10196_bfr_after (
		.din(new_net_10195),
		.dout(new_net_10196)
	);

	bfr new_net_10197_bfr_after (
		.din(new_net_10196),
		.dout(new_net_10197)
	);

	bfr new_net_10198_bfr_after (
		.din(new_net_10197),
		.dout(new_net_10198)
	);

	bfr new_net_10199_bfr_after (
		.din(new_net_10198),
		.dout(new_net_10199)
	);

	bfr new_net_10200_bfr_after (
		.din(new_net_10199),
		.dout(new_net_10200)
	);

	bfr new_net_10201_bfr_after (
		.din(new_net_10200),
		.dout(new_net_10201)
	);

	bfr new_net_10202_bfr_after (
		.din(new_net_10201),
		.dout(new_net_10202)
	);

	bfr new_net_10203_bfr_after (
		.din(new_net_10202),
		.dout(new_net_10203)
	);

	bfr new_net_10204_bfr_after (
		.din(new_net_10203),
		.dout(new_net_10204)
	);

	bfr new_net_10205_bfr_after (
		.din(new_net_10204),
		.dout(new_net_10205)
	);

	bfr new_net_10206_bfr_after (
		.din(new_net_10205),
		.dout(new_net_10206)
	);

	bfr new_net_10207_bfr_after (
		.din(new_net_10206),
		.dout(new_net_10207)
	);

	bfr new_net_10208_bfr_after (
		.din(new_net_10207),
		.dout(new_net_10208)
	);

	bfr new_net_10209_bfr_after (
		.din(new_net_10208),
		.dout(new_net_10209)
	);

	bfr new_net_10210_bfr_after (
		.din(new_net_10209),
		.dout(new_net_10210)
	);

	bfr new_net_10211_bfr_after (
		.din(new_net_10210),
		.dout(new_net_10211)
	);

	bfr new_net_10212_bfr_after (
		.din(new_net_10211),
		.dout(new_net_10212)
	);

	spl2 _0619__v_fanout (
		.a(new_net_10212),
		.b(new_net_657),
		.c(new_net_658)
	);

	bfr new_net_10213_bfr_after (
		.din(_0331_),
		.dout(new_net_10213)
	);

	bfr new_net_10214_bfr_after (
		.din(new_net_10213),
		.dout(new_net_10214)
	);

	bfr new_net_10215_bfr_after (
		.din(new_net_10214),
		.dout(new_net_10215)
	);

	bfr new_net_10216_bfr_after (
		.din(new_net_10215),
		.dout(new_net_10216)
	);

	bfr new_net_10217_bfr_after (
		.din(new_net_10216),
		.dout(new_net_10217)
	);

	bfr new_net_10218_bfr_after (
		.din(new_net_10217),
		.dout(new_net_10218)
	);

	bfr new_net_10219_bfr_after (
		.din(new_net_10218),
		.dout(new_net_10219)
	);

	bfr new_net_10220_bfr_after (
		.din(new_net_10219),
		.dout(new_net_10220)
	);

	bfr new_net_10221_bfr_after (
		.din(new_net_10220),
		.dout(new_net_10221)
	);

	bfr new_net_10222_bfr_after (
		.din(new_net_10221),
		.dout(new_net_10222)
	);

	bfr new_net_10223_bfr_after (
		.din(new_net_10222),
		.dout(new_net_10223)
	);

	bfr new_net_10224_bfr_after (
		.din(new_net_10223),
		.dout(new_net_10224)
	);

	bfr new_net_10225_bfr_after (
		.din(new_net_10224),
		.dout(new_net_10225)
	);

	bfr new_net_10226_bfr_after (
		.din(new_net_10225),
		.dout(new_net_10226)
	);

	bfr new_net_10227_bfr_after (
		.din(new_net_10226),
		.dout(new_net_10227)
	);

	bfr new_net_10228_bfr_after (
		.din(new_net_10227),
		.dout(new_net_10228)
	);

	bfr new_net_10229_bfr_after (
		.din(new_net_10228),
		.dout(new_net_10229)
	);

	bfr new_net_10230_bfr_after (
		.din(new_net_10229),
		.dout(new_net_10230)
	);

	bfr new_net_10231_bfr_after (
		.din(new_net_10230),
		.dout(new_net_10231)
	);

	bfr new_net_10232_bfr_after (
		.din(new_net_10231),
		.dout(new_net_10232)
	);

	bfr new_net_10233_bfr_after (
		.din(new_net_10232),
		.dout(new_net_10233)
	);

	bfr new_net_10234_bfr_after (
		.din(new_net_10233),
		.dout(new_net_10234)
	);

	bfr new_net_10235_bfr_after (
		.din(new_net_10234),
		.dout(new_net_10235)
	);

	bfr new_net_10236_bfr_after (
		.din(new_net_10235),
		.dout(new_net_10236)
	);

	bfr new_net_10237_bfr_after (
		.din(new_net_10236),
		.dout(new_net_10237)
	);

	bfr new_net_10238_bfr_after (
		.din(new_net_10237),
		.dout(new_net_10238)
	);

	bfr new_net_10239_bfr_after (
		.din(new_net_10238),
		.dout(new_net_10239)
	);

	bfr new_net_10240_bfr_after (
		.din(new_net_10239),
		.dout(new_net_10240)
	);

	bfr new_net_10241_bfr_after (
		.din(new_net_10240),
		.dout(new_net_10241)
	);

	bfr new_net_10242_bfr_after (
		.din(new_net_10241),
		.dout(new_net_10242)
	);

	bfr new_net_10243_bfr_after (
		.din(new_net_10242),
		.dout(new_net_10243)
	);

	bfr new_net_10244_bfr_after (
		.din(new_net_10243),
		.dout(new_net_10244)
	);

	bfr new_net_10245_bfr_after (
		.din(new_net_10244),
		.dout(new_net_10245)
	);

	bfr new_net_10246_bfr_after (
		.din(new_net_10245),
		.dout(new_net_10246)
	);

	bfr new_net_10247_bfr_after (
		.din(new_net_10246),
		.dout(new_net_10247)
	);

	bfr new_net_10248_bfr_after (
		.din(new_net_10247),
		.dout(new_net_10248)
	);

	bfr new_net_10249_bfr_after (
		.din(new_net_10248),
		.dout(new_net_10249)
	);

	bfr new_net_10250_bfr_after (
		.din(new_net_10249),
		.dout(new_net_10250)
	);

	bfr new_net_10251_bfr_after (
		.din(new_net_10250),
		.dout(new_net_10251)
	);

	bfr new_net_10252_bfr_after (
		.din(new_net_10251),
		.dout(new_net_10252)
	);

	bfr new_net_10253_bfr_after (
		.din(new_net_10252),
		.dout(new_net_10253)
	);

	bfr new_net_10254_bfr_after (
		.din(new_net_10253),
		.dout(new_net_10254)
	);

	bfr new_net_10255_bfr_after (
		.din(new_net_10254),
		.dout(new_net_10255)
	);

	bfr new_net_10256_bfr_after (
		.din(new_net_10255),
		.dout(new_net_10256)
	);

	bfr new_net_10257_bfr_after (
		.din(new_net_10256),
		.dout(new_net_10257)
	);

	bfr new_net_10258_bfr_after (
		.din(new_net_10257),
		.dout(new_net_10258)
	);

	bfr new_net_10259_bfr_after (
		.din(new_net_10258),
		.dout(new_net_10259)
	);

	bfr new_net_10260_bfr_after (
		.din(new_net_10259),
		.dout(new_net_10260)
	);

	bfr new_net_10261_bfr_after (
		.din(new_net_10260),
		.dout(new_net_10261)
	);

	bfr new_net_10262_bfr_after (
		.din(new_net_10261),
		.dout(new_net_10262)
	);

	bfr new_net_10263_bfr_after (
		.din(new_net_10262),
		.dout(new_net_10263)
	);

	bfr new_net_10264_bfr_after (
		.din(new_net_10263),
		.dout(new_net_10264)
	);

	bfr new_net_10265_bfr_after (
		.din(new_net_10264),
		.dout(new_net_10265)
	);

	bfr new_net_10266_bfr_after (
		.din(new_net_10265),
		.dout(new_net_10266)
	);

	bfr new_net_10267_bfr_after (
		.din(new_net_10266),
		.dout(new_net_10267)
	);

	bfr new_net_10268_bfr_after (
		.din(new_net_10267),
		.dout(new_net_10268)
	);

	bfr new_net_10269_bfr_after (
		.din(new_net_10268),
		.dout(new_net_10269)
	);

	bfr new_net_10270_bfr_after (
		.din(new_net_10269),
		.dout(new_net_10270)
	);

	bfr new_net_10271_bfr_after (
		.din(new_net_10270),
		.dout(new_net_10271)
	);

	bfr new_net_10272_bfr_after (
		.din(new_net_10271),
		.dout(new_net_10272)
	);

	bfr new_net_10273_bfr_after (
		.din(new_net_10272),
		.dout(new_net_10273)
	);

	bfr new_net_10274_bfr_after (
		.din(new_net_10273),
		.dout(new_net_10274)
	);

	bfr new_net_10275_bfr_after (
		.din(new_net_10274),
		.dout(new_net_10275)
	);

	bfr new_net_10276_bfr_after (
		.din(new_net_10275),
		.dout(new_net_10276)
	);

	bfr new_net_10277_bfr_after (
		.din(new_net_10276),
		.dout(new_net_10277)
	);

	bfr new_net_10278_bfr_after (
		.din(new_net_10277),
		.dout(new_net_10278)
	);

	bfr new_net_10279_bfr_after (
		.din(new_net_10278),
		.dout(new_net_10279)
	);

	bfr new_net_10280_bfr_after (
		.din(new_net_10279),
		.dout(new_net_10280)
	);

	bfr new_net_10281_bfr_after (
		.din(new_net_10280),
		.dout(new_net_10281)
	);

	bfr new_net_10282_bfr_after (
		.din(new_net_10281),
		.dout(new_net_10282)
	);

	bfr new_net_10283_bfr_after (
		.din(new_net_10282),
		.dout(new_net_10283)
	);

	bfr new_net_10284_bfr_after (
		.din(new_net_10283),
		.dout(new_net_10284)
	);

	bfr new_net_10285_bfr_after (
		.din(new_net_10284),
		.dout(new_net_10285)
	);

	bfr new_net_10286_bfr_after (
		.din(new_net_10285),
		.dout(new_net_10286)
	);

	bfr new_net_10287_bfr_after (
		.din(new_net_10286),
		.dout(new_net_10287)
	);

	bfr new_net_10288_bfr_after (
		.din(new_net_10287),
		.dout(new_net_10288)
	);

	bfr new_net_10289_bfr_after (
		.din(new_net_10288),
		.dout(new_net_10289)
	);

	bfr new_net_10290_bfr_after (
		.din(new_net_10289),
		.dout(new_net_10290)
	);

	bfr new_net_10291_bfr_after (
		.din(new_net_10290),
		.dout(new_net_10291)
	);

	bfr new_net_10292_bfr_after (
		.din(new_net_10291),
		.dout(new_net_10292)
	);

	bfr new_net_10293_bfr_after (
		.din(new_net_10292),
		.dout(new_net_10293)
	);

	bfr new_net_10294_bfr_after (
		.din(new_net_10293),
		.dout(new_net_10294)
	);

	bfr new_net_10295_bfr_after (
		.din(new_net_10294),
		.dout(new_net_10295)
	);

	bfr new_net_10296_bfr_after (
		.din(new_net_10295),
		.dout(new_net_10296)
	);

	bfr new_net_10297_bfr_after (
		.din(new_net_10296),
		.dout(new_net_10297)
	);

	bfr new_net_10298_bfr_after (
		.din(new_net_10297),
		.dout(new_net_10298)
	);

	bfr new_net_10299_bfr_after (
		.din(new_net_10298),
		.dout(new_net_10299)
	);

	bfr new_net_10300_bfr_after (
		.din(new_net_10299),
		.dout(new_net_10300)
	);

	bfr new_net_10301_bfr_after (
		.din(new_net_10300),
		.dout(new_net_10301)
	);

	bfr new_net_10302_bfr_after (
		.din(new_net_10301),
		.dout(new_net_10302)
	);

	bfr new_net_10303_bfr_after (
		.din(new_net_10302),
		.dout(new_net_10303)
	);

	bfr new_net_10304_bfr_after (
		.din(new_net_10303),
		.dout(new_net_10304)
	);

	bfr new_net_10305_bfr_after (
		.din(new_net_10304),
		.dout(new_net_10305)
	);

	bfr new_net_10306_bfr_after (
		.din(new_net_10305),
		.dout(new_net_10306)
	);

	bfr new_net_10307_bfr_after (
		.din(new_net_10306),
		.dout(new_net_10307)
	);

	bfr new_net_10308_bfr_after (
		.din(new_net_10307),
		.dout(new_net_10308)
	);

	spl2 _0331__v_fanout (
		.a(new_net_10308),
		.b(new_net_900),
		.c(new_net_901)
	);

	bfr new_net_10309_bfr_after (
		.din(_0699_),
		.dout(new_net_10309)
	);

	bfr new_net_10310_bfr_after (
		.din(new_net_10309),
		.dout(new_net_10310)
	);

	bfr new_net_10311_bfr_after (
		.din(new_net_10310),
		.dout(new_net_10311)
	);

	bfr new_net_10312_bfr_after (
		.din(new_net_10311),
		.dout(new_net_10312)
	);

	bfr new_net_10313_bfr_after (
		.din(new_net_10312),
		.dout(new_net_10313)
	);

	bfr new_net_10314_bfr_after (
		.din(new_net_10313),
		.dout(new_net_10314)
	);

	bfr new_net_10315_bfr_after (
		.din(new_net_10314),
		.dout(new_net_10315)
	);

	bfr new_net_10316_bfr_after (
		.din(new_net_10315),
		.dout(new_net_10316)
	);

	bfr new_net_10317_bfr_after (
		.din(new_net_10316),
		.dout(new_net_10317)
	);

	bfr new_net_10318_bfr_after (
		.din(new_net_10317),
		.dout(new_net_10318)
	);

	bfr new_net_10319_bfr_after (
		.din(new_net_10318),
		.dout(new_net_10319)
	);

	bfr new_net_10320_bfr_after (
		.din(new_net_10319),
		.dout(new_net_10320)
	);

	bfr new_net_10321_bfr_after (
		.din(new_net_10320),
		.dout(new_net_10321)
	);

	bfr new_net_10322_bfr_after (
		.din(new_net_10321),
		.dout(new_net_10322)
	);

	bfr new_net_10323_bfr_after (
		.din(new_net_10322),
		.dout(new_net_10323)
	);

	bfr new_net_10324_bfr_after (
		.din(new_net_10323),
		.dout(new_net_10324)
	);

	bfr new_net_10325_bfr_after (
		.din(new_net_10324),
		.dout(new_net_10325)
	);

	bfr new_net_10326_bfr_after (
		.din(new_net_10325),
		.dout(new_net_10326)
	);

	bfr new_net_10327_bfr_after (
		.din(new_net_10326),
		.dout(new_net_10327)
	);

	bfr new_net_10328_bfr_after (
		.din(new_net_10327),
		.dout(new_net_10328)
	);

	bfr new_net_10329_bfr_after (
		.din(new_net_10328),
		.dout(new_net_10329)
	);

	bfr new_net_10330_bfr_after (
		.din(new_net_10329),
		.dout(new_net_10330)
	);

	bfr new_net_10331_bfr_after (
		.din(new_net_10330),
		.dout(new_net_10331)
	);

	bfr new_net_10332_bfr_after (
		.din(new_net_10331),
		.dout(new_net_10332)
	);

	bfr new_net_10333_bfr_after (
		.din(new_net_10332),
		.dout(new_net_10333)
	);

	bfr new_net_10334_bfr_after (
		.din(new_net_10333),
		.dout(new_net_10334)
	);

	bfr new_net_10335_bfr_after (
		.din(new_net_10334),
		.dout(new_net_10335)
	);

	bfr new_net_10336_bfr_after (
		.din(new_net_10335),
		.dout(new_net_10336)
	);

	bfr new_net_10337_bfr_after (
		.din(new_net_10336),
		.dout(new_net_10337)
	);

	bfr new_net_10338_bfr_after (
		.din(new_net_10337),
		.dout(new_net_10338)
	);

	bfr new_net_10339_bfr_after (
		.din(new_net_10338),
		.dout(new_net_10339)
	);

	bfr new_net_10340_bfr_after (
		.din(new_net_10339),
		.dout(new_net_10340)
	);

	bfr new_net_10341_bfr_after (
		.din(new_net_10340),
		.dout(new_net_10341)
	);

	bfr new_net_10342_bfr_after (
		.din(new_net_10341),
		.dout(new_net_10342)
	);

	bfr new_net_10343_bfr_after (
		.din(new_net_10342),
		.dout(new_net_10343)
	);

	bfr new_net_10344_bfr_after (
		.din(new_net_10343),
		.dout(new_net_10344)
	);

	bfr new_net_10345_bfr_after (
		.din(new_net_10344),
		.dout(new_net_10345)
	);

	bfr new_net_10346_bfr_after (
		.din(new_net_10345),
		.dout(new_net_10346)
	);

	bfr new_net_10347_bfr_after (
		.din(new_net_10346),
		.dout(new_net_10347)
	);

	bfr new_net_10348_bfr_after (
		.din(new_net_10347),
		.dout(new_net_10348)
	);

	bfr new_net_10349_bfr_after (
		.din(new_net_10348),
		.dout(new_net_10349)
	);

	bfr new_net_10350_bfr_after (
		.din(new_net_10349),
		.dout(new_net_10350)
	);

	bfr new_net_10351_bfr_after (
		.din(new_net_10350),
		.dout(new_net_10351)
	);

	bfr new_net_10352_bfr_after (
		.din(new_net_10351),
		.dout(new_net_10352)
	);

	bfr new_net_10353_bfr_after (
		.din(new_net_10352),
		.dout(new_net_10353)
	);

	bfr new_net_10354_bfr_after (
		.din(new_net_10353),
		.dout(new_net_10354)
	);

	bfr new_net_10355_bfr_after (
		.din(new_net_10354),
		.dout(new_net_10355)
	);

	bfr new_net_10356_bfr_after (
		.din(new_net_10355),
		.dout(new_net_10356)
	);

	bfr new_net_10357_bfr_after (
		.din(new_net_10356),
		.dout(new_net_10357)
	);

	bfr new_net_10358_bfr_after (
		.din(new_net_10357),
		.dout(new_net_10358)
	);

	bfr new_net_10359_bfr_after (
		.din(new_net_10358),
		.dout(new_net_10359)
	);

	bfr new_net_10360_bfr_after (
		.din(new_net_10359),
		.dout(new_net_10360)
	);

	bfr new_net_10361_bfr_after (
		.din(new_net_10360),
		.dout(new_net_10361)
	);

	bfr new_net_10362_bfr_after (
		.din(new_net_10361),
		.dout(new_net_10362)
	);

	bfr new_net_10363_bfr_after (
		.din(new_net_10362),
		.dout(new_net_10363)
	);

	bfr new_net_10364_bfr_after (
		.din(new_net_10363),
		.dout(new_net_10364)
	);

	bfr new_net_10365_bfr_after (
		.din(new_net_10364),
		.dout(new_net_10365)
	);

	bfr new_net_10366_bfr_after (
		.din(new_net_10365),
		.dout(new_net_10366)
	);

	bfr new_net_10367_bfr_after (
		.din(new_net_10366),
		.dout(new_net_10367)
	);

	bfr new_net_10368_bfr_after (
		.din(new_net_10367),
		.dout(new_net_10368)
	);

	bfr new_net_10369_bfr_after (
		.din(new_net_10368),
		.dout(new_net_10369)
	);

	bfr new_net_10370_bfr_after (
		.din(new_net_10369),
		.dout(new_net_10370)
	);

	bfr new_net_10371_bfr_after (
		.din(new_net_10370),
		.dout(new_net_10371)
	);

	bfr new_net_10372_bfr_after (
		.din(new_net_10371),
		.dout(new_net_10372)
	);

	bfr new_net_10373_bfr_after (
		.din(new_net_10372),
		.dout(new_net_10373)
	);

	bfr new_net_10374_bfr_after (
		.din(new_net_10373),
		.dout(new_net_10374)
	);

	bfr new_net_10375_bfr_after (
		.din(new_net_10374),
		.dout(new_net_10375)
	);

	bfr new_net_10376_bfr_after (
		.din(new_net_10375),
		.dout(new_net_10376)
	);

	bfr new_net_10377_bfr_after (
		.din(new_net_10376),
		.dout(new_net_10377)
	);

	bfr new_net_10378_bfr_after (
		.din(new_net_10377),
		.dout(new_net_10378)
	);

	bfr new_net_10379_bfr_after (
		.din(new_net_10378),
		.dout(new_net_10379)
	);

	bfr new_net_10380_bfr_after (
		.din(new_net_10379),
		.dout(new_net_10380)
	);

	bfr new_net_10381_bfr_after (
		.din(new_net_10380),
		.dout(new_net_10381)
	);

	bfr new_net_10382_bfr_after (
		.din(new_net_10381),
		.dout(new_net_10382)
	);

	bfr new_net_10383_bfr_after (
		.din(new_net_10382),
		.dout(new_net_10383)
	);

	bfr new_net_10384_bfr_after (
		.din(new_net_10383),
		.dout(new_net_10384)
	);

	bfr new_net_10385_bfr_after (
		.din(new_net_10384),
		.dout(new_net_10385)
	);

	bfr new_net_10386_bfr_after (
		.din(new_net_10385),
		.dout(new_net_10386)
	);

	bfr new_net_10387_bfr_after (
		.din(new_net_10386),
		.dout(new_net_10387)
	);

	bfr new_net_10388_bfr_after (
		.din(new_net_10387),
		.dout(new_net_10388)
	);

	bfr new_net_10389_bfr_after (
		.din(new_net_10388),
		.dout(new_net_10389)
	);

	bfr new_net_10390_bfr_after (
		.din(new_net_10389),
		.dout(new_net_10390)
	);

	bfr new_net_10391_bfr_after (
		.din(new_net_10390),
		.dout(new_net_10391)
	);

	bfr new_net_10392_bfr_after (
		.din(new_net_10391),
		.dout(new_net_10392)
	);

	bfr new_net_10393_bfr_after (
		.din(new_net_10392),
		.dout(new_net_10393)
	);

	bfr new_net_10394_bfr_after (
		.din(new_net_10393),
		.dout(new_net_10394)
	);

	bfr new_net_10395_bfr_after (
		.din(new_net_10394),
		.dout(new_net_10395)
	);

	bfr new_net_10396_bfr_after (
		.din(new_net_10395),
		.dout(new_net_10396)
	);

	bfr new_net_10397_bfr_after (
		.din(new_net_10396),
		.dout(new_net_10397)
	);

	bfr new_net_10398_bfr_after (
		.din(new_net_10397),
		.dout(new_net_10398)
	);

	bfr new_net_10399_bfr_after (
		.din(new_net_10398),
		.dout(new_net_10399)
	);

	bfr new_net_10400_bfr_after (
		.din(new_net_10399),
		.dout(new_net_10400)
	);

	bfr new_net_10401_bfr_after (
		.din(new_net_10400),
		.dout(new_net_10401)
	);

	bfr new_net_10402_bfr_after (
		.din(new_net_10401),
		.dout(new_net_10402)
	);

	bfr new_net_10403_bfr_after (
		.din(new_net_10402),
		.dout(new_net_10403)
	);

	bfr new_net_10404_bfr_after (
		.din(new_net_10403),
		.dout(new_net_10404)
	);

	bfr new_net_10405_bfr_after (
		.din(new_net_10404),
		.dout(new_net_10405)
	);

	bfr new_net_10406_bfr_after (
		.din(new_net_10405),
		.dout(new_net_10406)
	);

	bfr new_net_10407_bfr_after (
		.din(new_net_10406),
		.dout(new_net_10407)
	);

	bfr new_net_10408_bfr_after (
		.din(new_net_10407),
		.dout(new_net_10408)
	);

	bfr new_net_10409_bfr_after (
		.din(new_net_10408),
		.dout(new_net_10409)
	);

	bfr new_net_10410_bfr_after (
		.din(new_net_10409),
		.dout(new_net_10410)
	);

	bfr new_net_10411_bfr_after (
		.din(new_net_10410),
		.dout(new_net_10411)
	);

	bfr new_net_10412_bfr_after (
		.din(new_net_10411),
		.dout(new_net_10412)
	);

	spl2 _0699__v_fanout (
		.a(new_net_10412),
		.b(new_net_2124),
		.c(new_net_2125)
	);

	bfr new_net_10413_bfr_after (
		.din(_0540_),
		.dout(new_net_10413)
	);

	bfr new_net_10414_bfr_after (
		.din(new_net_10413),
		.dout(new_net_10414)
	);

	bfr new_net_10415_bfr_after (
		.din(new_net_10414),
		.dout(new_net_10415)
	);

	bfr new_net_10416_bfr_after (
		.din(new_net_10415),
		.dout(new_net_10416)
	);

	bfr new_net_10417_bfr_after (
		.din(new_net_10416),
		.dout(new_net_10417)
	);

	bfr new_net_10418_bfr_after (
		.din(new_net_10417),
		.dout(new_net_10418)
	);

	bfr new_net_10419_bfr_after (
		.din(new_net_10418),
		.dout(new_net_10419)
	);

	bfr new_net_10420_bfr_after (
		.din(new_net_10419),
		.dout(new_net_10420)
	);

	bfr new_net_10421_bfr_after (
		.din(new_net_10420),
		.dout(new_net_10421)
	);

	bfr new_net_10422_bfr_after (
		.din(new_net_10421),
		.dout(new_net_10422)
	);

	bfr new_net_10423_bfr_after (
		.din(new_net_10422),
		.dout(new_net_10423)
	);

	bfr new_net_10424_bfr_after (
		.din(new_net_10423),
		.dout(new_net_10424)
	);

	bfr new_net_10425_bfr_after (
		.din(new_net_10424),
		.dout(new_net_10425)
	);

	bfr new_net_10426_bfr_after (
		.din(new_net_10425),
		.dout(new_net_10426)
	);

	bfr new_net_10427_bfr_after (
		.din(new_net_10426),
		.dout(new_net_10427)
	);

	bfr new_net_10428_bfr_after (
		.din(new_net_10427),
		.dout(new_net_10428)
	);

	bfr new_net_10429_bfr_after (
		.din(new_net_10428),
		.dout(new_net_10429)
	);

	bfr new_net_10430_bfr_after (
		.din(new_net_10429),
		.dout(new_net_10430)
	);

	bfr new_net_10431_bfr_after (
		.din(new_net_10430),
		.dout(new_net_10431)
	);

	bfr new_net_10432_bfr_after (
		.din(new_net_10431),
		.dout(new_net_10432)
	);

	bfr new_net_10433_bfr_after (
		.din(new_net_10432),
		.dout(new_net_10433)
	);

	bfr new_net_10434_bfr_after (
		.din(new_net_10433),
		.dout(new_net_10434)
	);

	bfr new_net_10435_bfr_after (
		.din(new_net_10434),
		.dout(new_net_10435)
	);

	bfr new_net_10436_bfr_after (
		.din(new_net_10435),
		.dout(new_net_10436)
	);

	bfr new_net_10437_bfr_after (
		.din(new_net_10436),
		.dout(new_net_10437)
	);

	bfr new_net_10438_bfr_after (
		.din(new_net_10437),
		.dout(new_net_10438)
	);

	bfr new_net_10439_bfr_after (
		.din(new_net_10438),
		.dout(new_net_10439)
	);

	bfr new_net_10440_bfr_after (
		.din(new_net_10439),
		.dout(new_net_10440)
	);

	bfr new_net_10441_bfr_after (
		.din(new_net_10440),
		.dout(new_net_10441)
	);

	bfr new_net_10442_bfr_after (
		.din(new_net_10441),
		.dout(new_net_10442)
	);

	bfr new_net_10443_bfr_after (
		.din(new_net_10442),
		.dout(new_net_10443)
	);

	bfr new_net_10444_bfr_after (
		.din(new_net_10443),
		.dout(new_net_10444)
	);

	bfr new_net_10445_bfr_after (
		.din(new_net_10444),
		.dout(new_net_10445)
	);

	bfr new_net_10446_bfr_after (
		.din(new_net_10445),
		.dout(new_net_10446)
	);

	bfr new_net_10447_bfr_after (
		.din(new_net_10446),
		.dout(new_net_10447)
	);

	bfr new_net_10448_bfr_after (
		.din(new_net_10447),
		.dout(new_net_10448)
	);

	bfr new_net_10449_bfr_after (
		.din(new_net_10448),
		.dout(new_net_10449)
	);

	bfr new_net_10450_bfr_after (
		.din(new_net_10449),
		.dout(new_net_10450)
	);

	bfr new_net_10451_bfr_after (
		.din(new_net_10450),
		.dout(new_net_10451)
	);

	bfr new_net_10452_bfr_after (
		.din(new_net_10451),
		.dout(new_net_10452)
	);

	bfr new_net_10453_bfr_after (
		.din(new_net_10452),
		.dout(new_net_10453)
	);

	bfr new_net_10454_bfr_after (
		.din(new_net_10453),
		.dout(new_net_10454)
	);

	bfr new_net_10455_bfr_after (
		.din(new_net_10454),
		.dout(new_net_10455)
	);

	bfr new_net_10456_bfr_after (
		.din(new_net_10455),
		.dout(new_net_10456)
	);

	bfr new_net_10457_bfr_after (
		.din(new_net_10456),
		.dout(new_net_10457)
	);

	bfr new_net_10458_bfr_after (
		.din(new_net_10457),
		.dout(new_net_10458)
	);

	bfr new_net_10459_bfr_after (
		.din(new_net_10458),
		.dout(new_net_10459)
	);

	bfr new_net_10460_bfr_after (
		.din(new_net_10459),
		.dout(new_net_10460)
	);

	bfr new_net_10461_bfr_after (
		.din(new_net_10460),
		.dout(new_net_10461)
	);

	bfr new_net_10462_bfr_after (
		.din(new_net_10461),
		.dout(new_net_10462)
	);

	bfr new_net_10463_bfr_after (
		.din(new_net_10462),
		.dout(new_net_10463)
	);

	bfr new_net_10464_bfr_after (
		.din(new_net_10463),
		.dout(new_net_10464)
	);

	bfr new_net_10465_bfr_after (
		.din(new_net_10464),
		.dout(new_net_10465)
	);

	bfr new_net_10466_bfr_after (
		.din(new_net_10465),
		.dout(new_net_10466)
	);

	bfr new_net_10467_bfr_after (
		.din(new_net_10466),
		.dout(new_net_10467)
	);

	bfr new_net_10468_bfr_after (
		.din(new_net_10467),
		.dout(new_net_10468)
	);

	bfr new_net_10469_bfr_after (
		.din(new_net_10468),
		.dout(new_net_10469)
	);

	bfr new_net_10470_bfr_after (
		.din(new_net_10469),
		.dout(new_net_10470)
	);

	bfr new_net_10471_bfr_after (
		.din(new_net_10470),
		.dout(new_net_10471)
	);

	bfr new_net_10472_bfr_after (
		.din(new_net_10471),
		.dout(new_net_10472)
	);

	bfr new_net_10473_bfr_after (
		.din(new_net_10472),
		.dout(new_net_10473)
	);

	bfr new_net_10474_bfr_after (
		.din(new_net_10473),
		.dout(new_net_10474)
	);

	bfr new_net_10475_bfr_after (
		.din(new_net_10474),
		.dout(new_net_10475)
	);

	bfr new_net_10476_bfr_after (
		.din(new_net_10475),
		.dout(new_net_10476)
	);

	bfr new_net_10477_bfr_after (
		.din(new_net_10476),
		.dout(new_net_10477)
	);

	bfr new_net_10478_bfr_after (
		.din(new_net_10477),
		.dout(new_net_10478)
	);

	bfr new_net_10479_bfr_after (
		.din(new_net_10478),
		.dout(new_net_10479)
	);

	bfr new_net_10480_bfr_after (
		.din(new_net_10479),
		.dout(new_net_10480)
	);

	bfr new_net_10481_bfr_after (
		.din(new_net_10480),
		.dout(new_net_10481)
	);

	bfr new_net_10482_bfr_after (
		.din(new_net_10481),
		.dout(new_net_10482)
	);

	bfr new_net_10483_bfr_after (
		.din(new_net_10482),
		.dout(new_net_10483)
	);

	bfr new_net_10484_bfr_after (
		.din(new_net_10483),
		.dout(new_net_10484)
	);

	spl2 _0540__v_fanout (
		.a(new_net_10484),
		.b(new_net_1696),
		.c(new_net_1697)
	);

	bfr new_net_10485_bfr_after (
		.din(_1580_),
		.dout(new_net_10485)
	);

	bfr new_net_10486_bfr_after (
		.din(new_net_10485),
		.dout(new_net_10486)
	);

	bfr new_net_10487_bfr_after (
		.din(new_net_10486),
		.dout(new_net_10487)
	);

	bfr new_net_10488_bfr_after (
		.din(new_net_10487),
		.dout(new_net_10488)
	);

	bfr new_net_10489_bfr_after (
		.din(new_net_10488),
		.dout(new_net_10489)
	);

	bfr new_net_10490_bfr_after (
		.din(new_net_10489),
		.dout(new_net_10490)
	);

	bfr new_net_10491_bfr_after (
		.din(new_net_10490),
		.dout(new_net_10491)
	);

	bfr new_net_10492_bfr_after (
		.din(new_net_10491),
		.dout(new_net_10492)
	);

	bfr new_net_10493_bfr_after (
		.din(new_net_10492),
		.dout(new_net_10493)
	);

	bfr new_net_10494_bfr_after (
		.din(new_net_10493),
		.dout(new_net_10494)
	);

	bfr new_net_10495_bfr_after (
		.din(new_net_10494),
		.dout(new_net_10495)
	);

	bfr new_net_10496_bfr_after (
		.din(new_net_10495),
		.dout(new_net_10496)
	);

	bfr new_net_10497_bfr_after (
		.din(new_net_10496),
		.dout(new_net_10497)
	);

	bfr new_net_10498_bfr_after (
		.din(new_net_10497),
		.dout(new_net_10498)
	);

	bfr new_net_10499_bfr_after (
		.din(new_net_10498),
		.dout(new_net_10499)
	);

	bfr new_net_10500_bfr_after (
		.din(new_net_10499),
		.dout(new_net_10500)
	);

	bfr new_net_10501_bfr_after (
		.din(new_net_10500),
		.dout(new_net_10501)
	);

	bfr new_net_10502_bfr_after (
		.din(new_net_10501),
		.dout(new_net_10502)
	);

	bfr new_net_10503_bfr_after (
		.din(new_net_10502),
		.dout(new_net_10503)
	);

	bfr new_net_10504_bfr_after (
		.din(new_net_10503),
		.dout(new_net_10504)
	);

	bfr new_net_10505_bfr_after (
		.din(new_net_10504),
		.dout(new_net_10505)
	);

	bfr new_net_10506_bfr_after (
		.din(new_net_10505),
		.dout(new_net_10506)
	);

	bfr new_net_10507_bfr_after (
		.din(new_net_10506),
		.dout(new_net_10507)
	);

	bfr new_net_10508_bfr_after (
		.din(new_net_10507),
		.dout(new_net_10508)
	);

	bfr new_net_10509_bfr_after (
		.din(new_net_10508),
		.dout(new_net_10509)
	);

	bfr new_net_10510_bfr_after (
		.din(new_net_10509),
		.dout(new_net_10510)
	);

	bfr new_net_10511_bfr_after (
		.din(new_net_10510),
		.dout(new_net_10511)
	);

	bfr new_net_10512_bfr_after (
		.din(new_net_10511),
		.dout(new_net_10512)
	);

	bfr new_net_10513_bfr_after (
		.din(new_net_10512),
		.dout(new_net_10513)
	);

	bfr new_net_10514_bfr_after (
		.din(new_net_10513),
		.dout(new_net_10514)
	);

	bfr new_net_10515_bfr_after (
		.din(new_net_10514),
		.dout(new_net_10515)
	);

	bfr new_net_10516_bfr_after (
		.din(new_net_10515),
		.dout(new_net_10516)
	);

	spl2 _1580__v_fanout (
		.a(new_net_10516),
		.b(new_net_2018),
		.c(new_net_2019)
	);

	bfr new_net_10517_bfr_after (
		.din(_0536_),
		.dout(new_net_10517)
	);

	bfr new_net_10518_bfr_after (
		.din(new_net_10517),
		.dout(new_net_10518)
	);

	bfr new_net_10519_bfr_after (
		.din(new_net_10518),
		.dout(new_net_10519)
	);

	bfr new_net_10520_bfr_after (
		.din(new_net_10519),
		.dout(new_net_10520)
	);

	bfr new_net_10521_bfr_after (
		.din(new_net_10520),
		.dout(new_net_10521)
	);

	bfr new_net_10522_bfr_after (
		.din(new_net_10521),
		.dout(new_net_10522)
	);

	bfr new_net_10523_bfr_after (
		.din(new_net_10522),
		.dout(new_net_10523)
	);

	bfr new_net_10524_bfr_after (
		.din(new_net_10523),
		.dout(new_net_10524)
	);

	bfr new_net_10525_bfr_after (
		.din(new_net_10524),
		.dout(new_net_10525)
	);

	bfr new_net_10526_bfr_after (
		.din(new_net_10525),
		.dout(new_net_10526)
	);

	bfr new_net_10527_bfr_after (
		.din(new_net_10526),
		.dout(new_net_10527)
	);

	bfr new_net_10528_bfr_after (
		.din(new_net_10527),
		.dout(new_net_10528)
	);

	bfr new_net_10529_bfr_after (
		.din(new_net_10528),
		.dout(new_net_10529)
	);

	bfr new_net_10530_bfr_after (
		.din(new_net_10529),
		.dout(new_net_10530)
	);

	bfr new_net_10531_bfr_after (
		.din(new_net_10530),
		.dout(new_net_10531)
	);

	bfr new_net_10532_bfr_after (
		.din(new_net_10531),
		.dout(new_net_10532)
	);

	bfr new_net_10533_bfr_after (
		.din(new_net_10532),
		.dout(new_net_10533)
	);

	bfr new_net_10534_bfr_after (
		.din(new_net_10533),
		.dout(new_net_10534)
	);

	bfr new_net_10535_bfr_after (
		.din(new_net_10534),
		.dout(new_net_10535)
	);

	bfr new_net_10536_bfr_after (
		.din(new_net_10535),
		.dout(new_net_10536)
	);

	bfr new_net_10537_bfr_after (
		.din(new_net_10536),
		.dout(new_net_10537)
	);

	bfr new_net_10538_bfr_after (
		.din(new_net_10537),
		.dout(new_net_10538)
	);

	bfr new_net_10539_bfr_after (
		.din(new_net_10538),
		.dout(new_net_10539)
	);

	bfr new_net_10540_bfr_after (
		.din(new_net_10539),
		.dout(new_net_10540)
	);

	bfr new_net_10541_bfr_after (
		.din(new_net_10540),
		.dout(new_net_10541)
	);

	bfr new_net_10542_bfr_after (
		.din(new_net_10541),
		.dout(new_net_10542)
	);

	bfr new_net_10543_bfr_after (
		.din(new_net_10542),
		.dout(new_net_10543)
	);

	bfr new_net_10544_bfr_after (
		.din(new_net_10543),
		.dout(new_net_10544)
	);

	bfr new_net_10545_bfr_after (
		.din(new_net_10544),
		.dout(new_net_10545)
	);

	bfr new_net_10546_bfr_after (
		.din(new_net_10545),
		.dout(new_net_10546)
	);

	bfr new_net_10547_bfr_after (
		.din(new_net_10546),
		.dout(new_net_10547)
	);

	bfr new_net_10548_bfr_after (
		.din(new_net_10547),
		.dout(new_net_10548)
	);

	bfr new_net_10549_bfr_after (
		.din(new_net_10548),
		.dout(new_net_10549)
	);

	bfr new_net_10550_bfr_after (
		.din(new_net_10549),
		.dout(new_net_10550)
	);

	bfr new_net_10551_bfr_after (
		.din(new_net_10550),
		.dout(new_net_10551)
	);

	bfr new_net_10552_bfr_after (
		.din(new_net_10551),
		.dout(new_net_10552)
	);

	bfr new_net_10553_bfr_after (
		.din(new_net_10552),
		.dout(new_net_10553)
	);

	bfr new_net_10554_bfr_after (
		.din(new_net_10553),
		.dout(new_net_10554)
	);

	bfr new_net_10555_bfr_after (
		.din(new_net_10554),
		.dout(new_net_10555)
	);

	bfr new_net_10556_bfr_after (
		.din(new_net_10555),
		.dout(new_net_10556)
	);

	bfr new_net_10557_bfr_after (
		.din(new_net_10556),
		.dout(new_net_10557)
	);

	bfr new_net_10558_bfr_after (
		.din(new_net_10557),
		.dout(new_net_10558)
	);

	bfr new_net_10559_bfr_after (
		.din(new_net_10558),
		.dout(new_net_10559)
	);

	bfr new_net_10560_bfr_after (
		.din(new_net_10559),
		.dout(new_net_10560)
	);

	bfr new_net_10561_bfr_after (
		.din(new_net_10560),
		.dout(new_net_10561)
	);

	bfr new_net_10562_bfr_after (
		.din(new_net_10561),
		.dout(new_net_10562)
	);

	bfr new_net_10563_bfr_after (
		.din(new_net_10562),
		.dout(new_net_10563)
	);

	bfr new_net_10564_bfr_after (
		.din(new_net_10563),
		.dout(new_net_10564)
	);

	bfr new_net_10565_bfr_after (
		.din(new_net_10564),
		.dout(new_net_10565)
	);

	bfr new_net_10566_bfr_after (
		.din(new_net_10565),
		.dout(new_net_10566)
	);

	bfr new_net_10567_bfr_after (
		.din(new_net_10566),
		.dout(new_net_10567)
	);

	bfr new_net_10568_bfr_after (
		.din(new_net_10567),
		.dout(new_net_10568)
	);

	bfr new_net_10569_bfr_after (
		.din(new_net_10568),
		.dout(new_net_10569)
	);

	bfr new_net_10570_bfr_after (
		.din(new_net_10569),
		.dout(new_net_10570)
	);

	bfr new_net_10571_bfr_after (
		.din(new_net_10570),
		.dout(new_net_10571)
	);

	bfr new_net_10572_bfr_after (
		.din(new_net_10571),
		.dout(new_net_10572)
	);

	bfr new_net_10573_bfr_after (
		.din(new_net_10572),
		.dout(new_net_10573)
	);

	bfr new_net_10574_bfr_after (
		.din(new_net_10573),
		.dout(new_net_10574)
	);

	bfr new_net_10575_bfr_after (
		.din(new_net_10574),
		.dout(new_net_10575)
	);

	bfr new_net_10576_bfr_after (
		.din(new_net_10575),
		.dout(new_net_10576)
	);

	bfr new_net_10577_bfr_after (
		.din(new_net_10576),
		.dout(new_net_10577)
	);

	bfr new_net_10578_bfr_after (
		.din(new_net_10577),
		.dout(new_net_10578)
	);

	bfr new_net_10579_bfr_after (
		.din(new_net_10578),
		.dout(new_net_10579)
	);

	bfr new_net_10580_bfr_after (
		.din(new_net_10579),
		.dout(new_net_10580)
	);

	bfr new_net_10581_bfr_after (
		.din(new_net_10580),
		.dout(new_net_10581)
	);

	bfr new_net_10582_bfr_after (
		.din(new_net_10581),
		.dout(new_net_10582)
	);

	bfr new_net_10583_bfr_after (
		.din(new_net_10582),
		.dout(new_net_10583)
	);

	bfr new_net_10584_bfr_after (
		.din(new_net_10583),
		.dout(new_net_10584)
	);

	bfr new_net_10585_bfr_after (
		.din(new_net_10584),
		.dout(new_net_10585)
	);

	bfr new_net_10586_bfr_after (
		.din(new_net_10585),
		.dout(new_net_10586)
	);

	bfr new_net_10587_bfr_after (
		.din(new_net_10586),
		.dout(new_net_10587)
	);

	bfr new_net_10588_bfr_after (
		.din(new_net_10587),
		.dout(new_net_10588)
	);

	bfr new_net_10589_bfr_after (
		.din(new_net_10588),
		.dout(new_net_10589)
	);

	bfr new_net_10590_bfr_after (
		.din(new_net_10589),
		.dout(new_net_10590)
	);

	bfr new_net_10591_bfr_after (
		.din(new_net_10590),
		.dout(new_net_10591)
	);

	bfr new_net_10592_bfr_after (
		.din(new_net_10591),
		.dout(new_net_10592)
	);

	bfr new_net_10593_bfr_after (
		.din(new_net_10592),
		.dout(new_net_10593)
	);

	bfr new_net_10594_bfr_after (
		.din(new_net_10593),
		.dout(new_net_10594)
	);

	bfr new_net_10595_bfr_after (
		.din(new_net_10594),
		.dout(new_net_10595)
	);

	bfr new_net_10596_bfr_after (
		.din(new_net_10595),
		.dout(new_net_10596)
	);

	bfr new_net_10597_bfr_after (
		.din(new_net_10596),
		.dout(new_net_10597)
	);

	bfr new_net_10598_bfr_after (
		.din(new_net_10597),
		.dout(new_net_10598)
	);

	bfr new_net_10599_bfr_after (
		.din(new_net_10598),
		.dout(new_net_10599)
	);

	bfr new_net_10600_bfr_after (
		.din(new_net_10599),
		.dout(new_net_10600)
	);

	bfr new_net_10601_bfr_after (
		.din(new_net_10600),
		.dout(new_net_10601)
	);

	bfr new_net_10602_bfr_after (
		.din(new_net_10601),
		.dout(new_net_10602)
	);

	bfr new_net_10603_bfr_after (
		.din(new_net_10602),
		.dout(new_net_10603)
	);

	bfr new_net_10604_bfr_after (
		.din(new_net_10603),
		.dout(new_net_10604)
	);

	spl2 _0536__v_fanout (
		.a(new_net_10604),
		.b(new_net_2260),
		.c(new_net_2261)
	);

	bfr new_net_10605_bfr_after (
		.din(_0342_),
		.dout(new_net_10605)
	);

	bfr new_net_10606_bfr_after (
		.din(new_net_10605),
		.dout(new_net_10606)
	);

	bfr new_net_10607_bfr_after (
		.din(new_net_10606),
		.dout(new_net_10607)
	);

	bfr new_net_10608_bfr_after (
		.din(new_net_10607),
		.dout(new_net_10608)
	);

	bfr new_net_10609_bfr_after (
		.din(new_net_10608),
		.dout(new_net_10609)
	);

	bfr new_net_10610_bfr_after (
		.din(new_net_10609),
		.dout(new_net_10610)
	);

	bfr new_net_10611_bfr_after (
		.din(new_net_10610),
		.dout(new_net_10611)
	);

	bfr new_net_10612_bfr_after (
		.din(new_net_10611),
		.dout(new_net_10612)
	);

	bfr new_net_10613_bfr_after (
		.din(new_net_10612),
		.dout(new_net_10613)
	);

	bfr new_net_10614_bfr_after (
		.din(new_net_10613),
		.dout(new_net_10614)
	);

	bfr new_net_10615_bfr_after (
		.din(new_net_10614),
		.dout(new_net_10615)
	);

	bfr new_net_10616_bfr_after (
		.din(new_net_10615),
		.dout(new_net_10616)
	);

	bfr new_net_10617_bfr_after (
		.din(new_net_10616),
		.dout(new_net_10617)
	);

	bfr new_net_10618_bfr_after (
		.din(new_net_10617),
		.dout(new_net_10618)
	);

	bfr new_net_10619_bfr_after (
		.din(new_net_10618),
		.dout(new_net_10619)
	);

	bfr new_net_10620_bfr_after (
		.din(new_net_10619),
		.dout(new_net_10620)
	);

	bfr new_net_10621_bfr_after (
		.din(new_net_10620),
		.dout(new_net_10621)
	);

	bfr new_net_10622_bfr_after (
		.din(new_net_10621),
		.dout(new_net_10622)
	);

	bfr new_net_10623_bfr_after (
		.din(new_net_10622),
		.dout(new_net_10623)
	);

	bfr new_net_10624_bfr_after (
		.din(new_net_10623),
		.dout(new_net_10624)
	);

	bfr new_net_10625_bfr_after (
		.din(new_net_10624),
		.dout(new_net_10625)
	);

	bfr new_net_10626_bfr_after (
		.din(new_net_10625),
		.dout(new_net_10626)
	);

	bfr new_net_10627_bfr_after (
		.din(new_net_10626),
		.dout(new_net_10627)
	);

	bfr new_net_10628_bfr_after (
		.din(new_net_10627),
		.dout(new_net_10628)
	);

	bfr new_net_10629_bfr_after (
		.din(new_net_10628),
		.dout(new_net_10629)
	);

	bfr new_net_10630_bfr_after (
		.din(new_net_10629),
		.dout(new_net_10630)
	);

	bfr new_net_10631_bfr_after (
		.din(new_net_10630),
		.dout(new_net_10631)
	);

	bfr new_net_10632_bfr_after (
		.din(new_net_10631),
		.dout(new_net_10632)
	);

	bfr new_net_10633_bfr_after (
		.din(new_net_10632),
		.dout(new_net_10633)
	);

	bfr new_net_10634_bfr_after (
		.din(new_net_10633),
		.dout(new_net_10634)
	);

	bfr new_net_10635_bfr_after (
		.din(new_net_10634),
		.dout(new_net_10635)
	);

	bfr new_net_10636_bfr_after (
		.din(new_net_10635),
		.dout(new_net_10636)
	);

	bfr new_net_10637_bfr_after (
		.din(new_net_10636),
		.dout(new_net_10637)
	);

	bfr new_net_10638_bfr_after (
		.din(new_net_10637),
		.dout(new_net_10638)
	);

	bfr new_net_10639_bfr_after (
		.din(new_net_10638),
		.dout(new_net_10639)
	);

	bfr new_net_10640_bfr_after (
		.din(new_net_10639),
		.dout(new_net_10640)
	);

	bfr new_net_10641_bfr_after (
		.din(new_net_10640),
		.dout(new_net_10641)
	);

	bfr new_net_10642_bfr_after (
		.din(new_net_10641),
		.dout(new_net_10642)
	);

	bfr new_net_10643_bfr_after (
		.din(new_net_10642),
		.dout(new_net_10643)
	);

	bfr new_net_10644_bfr_after (
		.din(new_net_10643),
		.dout(new_net_10644)
	);

	bfr new_net_10645_bfr_after (
		.din(new_net_10644),
		.dout(new_net_10645)
	);

	bfr new_net_10646_bfr_after (
		.din(new_net_10645),
		.dout(new_net_10646)
	);

	bfr new_net_10647_bfr_after (
		.din(new_net_10646),
		.dout(new_net_10647)
	);

	bfr new_net_10648_bfr_after (
		.din(new_net_10647),
		.dout(new_net_10648)
	);

	bfr new_net_10649_bfr_after (
		.din(new_net_10648),
		.dout(new_net_10649)
	);

	bfr new_net_10650_bfr_after (
		.din(new_net_10649),
		.dout(new_net_10650)
	);

	bfr new_net_10651_bfr_after (
		.din(new_net_10650),
		.dout(new_net_10651)
	);

	bfr new_net_10652_bfr_after (
		.din(new_net_10651),
		.dout(new_net_10652)
	);

	bfr new_net_10653_bfr_after (
		.din(new_net_10652),
		.dout(new_net_10653)
	);

	bfr new_net_10654_bfr_after (
		.din(new_net_10653),
		.dout(new_net_10654)
	);

	bfr new_net_10655_bfr_after (
		.din(new_net_10654),
		.dout(new_net_10655)
	);

	bfr new_net_10656_bfr_after (
		.din(new_net_10655),
		.dout(new_net_10656)
	);

	bfr new_net_10657_bfr_after (
		.din(new_net_10656),
		.dout(new_net_10657)
	);

	bfr new_net_10658_bfr_after (
		.din(new_net_10657),
		.dout(new_net_10658)
	);

	bfr new_net_10659_bfr_after (
		.din(new_net_10658),
		.dout(new_net_10659)
	);

	bfr new_net_10660_bfr_after (
		.din(new_net_10659),
		.dout(new_net_10660)
	);

	spl2 _0342__v_fanout (
		.a(new_net_10660),
		.b(new_net_1267),
		.c(new_net_1268)
	);

	bfr new_net_10661_bfr_after (
		.din(_1700_),
		.dout(new_net_10661)
	);

	bfr new_net_10662_bfr_after (
		.din(new_net_10661),
		.dout(new_net_10662)
	);

	bfr new_net_10663_bfr_after (
		.din(new_net_10662),
		.dout(new_net_10663)
	);

	bfr new_net_10664_bfr_after (
		.din(new_net_10663),
		.dout(new_net_10664)
	);

	bfr new_net_10665_bfr_after (
		.din(new_net_10664),
		.dout(new_net_10665)
	);

	bfr new_net_10666_bfr_after (
		.din(new_net_10665),
		.dout(new_net_10666)
	);

	bfr new_net_10667_bfr_after (
		.din(new_net_10666),
		.dout(new_net_10667)
	);

	bfr new_net_10668_bfr_after (
		.din(new_net_10667),
		.dout(new_net_10668)
	);

	bfr new_net_10669_bfr_after (
		.din(new_net_10668),
		.dout(new_net_10669)
	);

	bfr new_net_10670_bfr_after (
		.din(new_net_10669),
		.dout(new_net_10670)
	);

	bfr new_net_10671_bfr_after (
		.din(new_net_10670),
		.dout(new_net_10671)
	);

	bfr new_net_10672_bfr_after (
		.din(new_net_10671),
		.dout(new_net_10672)
	);

	bfr new_net_10673_bfr_after (
		.din(new_net_10672),
		.dout(new_net_10673)
	);

	bfr new_net_10674_bfr_after (
		.din(new_net_10673),
		.dout(new_net_10674)
	);

	bfr new_net_10675_bfr_after (
		.din(new_net_10674),
		.dout(new_net_10675)
	);

	bfr new_net_10676_bfr_after (
		.din(new_net_10675),
		.dout(new_net_10676)
	);

	bfr new_net_10677_bfr_after (
		.din(new_net_10676),
		.dout(new_net_10677)
	);

	bfr new_net_10678_bfr_after (
		.din(new_net_10677),
		.dout(new_net_10678)
	);

	bfr new_net_10679_bfr_after (
		.din(new_net_10678),
		.dout(new_net_10679)
	);

	bfr new_net_10680_bfr_after (
		.din(new_net_10679),
		.dout(new_net_10680)
	);

	bfr new_net_10681_bfr_after (
		.din(new_net_10680),
		.dout(new_net_10681)
	);

	bfr new_net_10682_bfr_after (
		.din(new_net_10681),
		.dout(new_net_10682)
	);

	bfr new_net_10683_bfr_after (
		.din(new_net_10682),
		.dout(new_net_10683)
	);

	bfr new_net_10684_bfr_after (
		.din(new_net_10683),
		.dout(new_net_10684)
	);

	bfr new_net_10685_bfr_after (
		.din(new_net_10684),
		.dout(new_net_10685)
	);

	bfr new_net_10686_bfr_after (
		.din(new_net_10685),
		.dout(new_net_10686)
	);

	bfr new_net_10687_bfr_after (
		.din(new_net_10686),
		.dout(new_net_10687)
	);

	bfr new_net_10688_bfr_after (
		.din(new_net_10687),
		.dout(new_net_10688)
	);

	bfr new_net_10689_bfr_after (
		.din(new_net_10688),
		.dout(new_net_10689)
	);

	bfr new_net_10690_bfr_after (
		.din(new_net_10689),
		.dout(new_net_10690)
	);

	bfr new_net_10691_bfr_after (
		.din(new_net_10690),
		.dout(new_net_10691)
	);

	bfr new_net_10692_bfr_after (
		.din(new_net_10691),
		.dout(new_net_10692)
	);

	spl2 _1700__v_fanout (
		.a(new_net_10692),
		.b(new_net_679),
		.c(new_net_680)
	);

	bfr new_net_10693_bfr_after (
		.din(_0349_),
		.dout(new_net_10693)
	);

	bfr new_net_10694_bfr_after (
		.din(new_net_10693),
		.dout(new_net_10694)
	);

	bfr new_net_10695_bfr_after (
		.din(new_net_10694),
		.dout(new_net_10695)
	);

	bfr new_net_10696_bfr_after (
		.din(new_net_10695),
		.dout(new_net_10696)
	);

	bfr new_net_10697_bfr_after (
		.din(new_net_10696),
		.dout(new_net_10697)
	);

	bfr new_net_10698_bfr_after (
		.din(new_net_10697),
		.dout(new_net_10698)
	);

	bfr new_net_10699_bfr_after (
		.din(new_net_10698),
		.dout(new_net_10699)
	);

	bfr new_net_10700_bfr_after (
		.din(new_net_10699),
		.dout(new_net_10700)
	);

	bfr new_net_10701_bfr_after (
		.din(new_net_10700),
		.dout(new_net_10701)
	);

	bfr new_net_10702_bfr_after (
		.din(new_net_10701),
		.dout(new_net_10702)
	);

	bfr new_net_10703_bfr_after (
		.din(new_net_10702),
		.dout(new_net_10703)
	);

	bfr new_net_10704_bfr_after (
		.din(new_net_10703),
		.dout(new_net_10704)
	);

	bfr new_net_10705_bfr_after (
		.din(new_net_10704),
		.dout(new_net_10705)
	);

	bfr new_net_10706_bfr_after (
		.din(new_net_10705),
		.dout(new_net_10706)
	);

	bfr new_net_10707_bfr_after (
		.din(new_net_10706),
		.dout(new_net_10707)
	);

	bfr new_net_10708_bfr_after (
		.din(new_net_10707),
		.dout(new_net_10708)
	);

	bfr new_net_10709_bfr_after (
		.din(new_net_10708),
		.dout(new_net_10709)
	);

	bfr new_net_10710_bfr_after (
		.din(new_net_10709),
		.dout(new_net_10710)
	);

	bfr new_net_10711_bfr_after (
		.din(new_net_10710),
		.dout(new_net_10711)
	);

	bfr new_net_10712_bfr_after (
		.din(new_net_10711),
		.dout(new_net_10712)
	);

	bfr new_net_10713_bfr_after (
		.din(new_net_10712),
		.dout(new_net_10713)
	);

	bfr new_net_10714_bfr_after (
		.din(new_net_10713),
		.dout(new_net_10714)
	);

	spl2 _0349__v_fanout (
		.a(new_net_10714),
		.b(new_net_1569),
		.c(new_net_1570)
	);

	spl2 _1469__v_fanout (
		.a(_1469_),
		.b(new_net_1020),
		.c(new_net_1021)
	);

	bfr new_net_10715_bfr_after (
		.din(_0100_),
		.dout(new_net_10715)
	);

	bfr new_net_10716_bfr_after (
		.din(new_net_10715),
		.dout(new_net_10716)
	);

	bfr new_net_10717_bfr_after (
		.din(new_net_10716),
		.dout(new_net_10717)
	);

	bfr new_net_10718_bfr_after (
		.din(new_net_10717),
		.dout(new_net_10718)
	);

	bfr new_net_10719_bfr_after (
		.din(new_net_10718),
		.dout(new_net_10719)
	);

	bfr new_net_10720_bfr_after (
		.din(new_net_10719),
		.dout(new_net_10720)
	);

	bfr new_net_10721_bfr_after (
		.din(new_net_10720),
		.dout(new_net_10721)
	);

	bfr new_net_10722_bfr_after (
		.din(new_net_10721),
		.dout(new_net_10722)
	);

	bfr new_net_10723_bfr_after (
		.din(new_net_10722),
		.dout(new_net_10723)
	);

	bfr new_net_10724_bfr_after (
		.din(new_net_10723),
		.dout(new_net_10724)
	);

	bfr new_net_10725_bfr_after (
		.din(new_net_10724),
		.dout(new_net_10725)
	);

	bfr new_net_10726_bfr_after (
		.din(new_net_10725),
		.dout(new_net_10726)
	);

	bfr new_net_10727_bfr_after (
		.din(new_net_10726),
		.dout(new_net_10727)
	);

	bfr new_net_10728_bfr_after (
		.din(new_net_10727),
		.dout(new_net_10728)
	);

	bfr new_net_10729_bfr_after (
		.din(new_net_10728),
		.dout(new_net_10729)
	);

	bfr new_net_10730_bfr_after (
		.din(new_net_10729),
		.dout(new_net_10730)
	);

	bfr new_net_10731_bfr_after (
		.din(new_net_10730),
		.dout(new_net_10731)
	);

	bfr new_net_10732_bfr_after (
		.din(new_net_10731),
		.dout(new_net_10732)
	);

	bfr new_net_10733_bfr_after (
		.din(new_net_10732),
		.dout(new_net_10733)
	);

	bfr new_net_10734_bfr_after (
		.din(new_net_10733),
		.dout(new_net_10734)
	);

	bfr new_net_10735_bfr_after (
		.din(new_net_10734),
		.dout(new_net_10735)
	);

	bfr new_net_10736_bfr_after (
		.din(new_net_10735),
		.dout(new_net_10736)
	);

	bfr new_net_10737_bfr_after (
		.din(new_net_10736),
		.dout(new_net_10737)
	);

	bfr new_net_10738_bfr_after (
		.din(new_net_10737),
		.dout(new_net_10738)
	);

	bfr new_net_10739_bfr_after (
		.din(new_net_10738),
		.dout(new_net_10739)
	);

	bfr new_net_10740_bfr_after (
		.din(new_net_10739),
		.dout(new_net_10740)
	);

	bfr new_net_10741_bfr_after (
		.din(new_net_10740),
		.dout(new_net_10741)
	);

	bfr new_net_10742_bfr_after (
		.din(new_net_10741),
		.dout(new_net_10742)
	);

	bfr new_net_10743_bfr_after (
		.din(new_net_10742),
		.dout(new_net_10743)
	);

	bfr new_net_10744_bfr_after (
		.din(new_net_10743),
		.dout(new_net_10744)
	);

	bfr new_net_10745_bfr_after (
		.din(new_net_10744),
		.dout(new_net_10745)
	);

	bfr new_net_10746_bfr_after (
		.din(new_net_10745),
		.dout(new_net_10746)
	);

	bfr new_net_10747_bfr_after (
		.din(new_net_10746),
		.dout(new_net_10747)
	);

	bfr new_net_10748_bfr_after (
		.din(new_net_10747),
		.dout(new_net_10748)
	);

	bfr new_net_10749_bfr_after (
		.din(new_net_10748),
		.dout(new_net_10749)
	);

	bfr new_net_10750_bfr_after (
		.din(new_net_10749),
		.dout(new_net_10750)
	);

	bfr new_net_10751_bfr_after (
		.din(new_net_10750),
		.dout(new_net_10751)
	);

	bfr new_net_10752_bfr_after (
		.din(new_net_10751),
		.dout(new_net_10752)
	);

	bfr new_net_10753_bfr_after (
		.din(new_net_10752),
		.dout(new_net_10753)
	);

	bfr new_net_10754_bfr_after (
		.din(new_net_10753),
		.dout(new_net_10754)
	);

	bfr new_net_10755_bfr_after (
		.din(new_net_10754),
		.dout(new_net_10755)
	);

	bfr new_net_10756_bfr_after (
		.din(new_net_10755),
		.dout(new_net_10756)
	);

	bfr new_net_10757_bfr_after (
		.din(new_net_10756),
		.dout(new_net_10757)
	);

	bfr new_net_10758_bfr_after (
		.din(new_net_10757),
		.dout(new_net_10758)
	);

	bfr new_net_10759_bfr_after (
		.din(new_net_10758),
		.dout(new_net_10759)
	);

	bfr new_net_10760_bfr_after (
		.din(new_net_10759),
		.dout(new_net_10760)
	);

	bfr new_net_10761_bfr_after (
		.din(new_net_10760),
		.dout(new_net_10761)
	);

	bfr new_net_10762_bfr_after (
		.din(new_net_10761),
		.dout(new_net_10762)
	);

	bfr new_net_10763_bfr_after (
		.din(new_net_10762),
		.dout(new_net_10763)
	);

	bfr new_net_10764_bfr_after (
		.din(new_net_10763),
		.dout(new_net_10764)
	);

	bfr new_net_10765_bfr_after (
		.din(new_net_10764),
		.dout(new_net_10765)
	);

	bfr new_net_10766_bfr_after (
		.din(new_net_10765),
		.dout(new_net_10766)
	);

	bfr new_net_10767_bfr_after (
		.din(new_net_10766),
		.dout(new_net_10767)
	);

	bfr new_net_10768_bfr_after (
		.din(new_net_10767),
		.dout(new_net_10768)
	);

	bfr new_net_10769_bfr_after (
		.din(new_net_10768),
		.dout(new_net_10769)
	);

	bfr new_net_10770_bfr_after (
		.din(new_net_10769),
		.dout(new_net_10770)
	);

	spl2 _0100__v_fanout (
		.a(new_net_10770),
		.b(new_net_735),
		.c(new_net_736)
	);

	bfr new_net_10771_bfr_after (
		.din(_1215_),
		.dout(new_net_10771)
	);

	bfr new_net_10772_bfr_after (
		.din(new_net_10771),
		.dout(new_net_10772)
	);

	bfr new_net_10773_bfr_after (
		.din(new_net_10772),
		.dout(new_net_10773)
	);

	bfr new_net_10774_bfr_after (
		.din(new_net_10773),
		.dout(new_net_10774)
	);

	bfr new_net_10775_bfr_after (
		.din(new_net_10774),
		.dout(new_net_10775)
	);

	bfr new_net_10776_bfr_after (
		.din(new_net_10775),
		.dout(new_net_10776)
	);

	bfr new_net_10777_bfr_after (
		.din(new_net_10776),
		.dout(new_net_10777)
	);

	bfr new_net_10778_bfr_after (
		.din(new_net_10777),
		.dout(new_net_10778)
	);

	bfr new_net_10779_bfr_after (
		.din(new_net_10778),
		.dout(new_net_10779)
	);

	bfr new_net_10780_bfr_after (
		.din(new_net_10779),
		.dout(new_net_10780)
	);

	bfr new_net_10781_bfr_after (
		.din(new_net_10780),
		.dout(new_net_10781)
	);

	bfr new_net_10782_bfr_after (
		.din(new_net_10781),
		.dout(new_net_10782)
	);

	bfr new_net_10783_bfr_after (
		.din(new_net_10782),
		.dout(new_net_10783)
	);

	bfr new_net_10784_bfr_after (
		.din(new_net_10783),
		.dout(new_net_10784)
	);

	bfr new_net_10785_bfr_after (
		.din(new_net_10784),
		.dout(new_net_10785)
	);

	bfr new_net_10786_bfr_after (
		.din(new_net_10785),
		.dout(new_net_10786)
	);

	bfr new_net_10787_bfr_after (
		.din(new_net_10786),
		.dout(new_net_10787)
	);

	bfr new_net_10788_bfr_after (
		.din(new_net_10787),
		.dout(new_net_10788)
	);

	bfr new_net_10789_bfr_after (
		.din(new_net_10788),
		.dout(new_net_10789)
	);

	bfr new_net_10790_bfr_after (
		.din(new_net_10789),
		.dout(new_net_10790)
	);

	bfr new_net_10791_bfr_after (
		.din(new_net_10790),
		.dout(new_net_10791)
	);

	bfr new_net_10792_bfr_after (
		.din(new_net_10791),
		.dout(new_net_10792)
	);

	bfr new_net_10793_bfr_after (
		.din(new_net_10792),
		.dout(new_net_10793)
	);

	bfr new_net_10794_bfr_after (
		.din(new_net_10793),
		.dout(new_net_10794)
	);

	spl2 _1215__v_fanout (
		.a(new_net_10794),
		.b(new_net_1964),
		.c(new_net_1965)
	);

	bfr new_net_10795_bfr_after (
		.din(_1823_),
		.dout(new_net_10795)
	);

	bfr new_net_10796_bfr_after (
		.din(new_net_10795),
		.dout(new_net_10796)
	);

	bfr new_net_10797_bfr_after (
		.din(new_net_10796),
		.dout(new_net_10797)
	);

	bfr new_net_10798_bfr_after (
		.din(new_net_10797),
		.dout(new_net_10798)
	);

	bfr new_net_10799_bfr_after (
		.din(new_net_10798),
		.dout(new_net_10799)
	);

	bfr new_net_10800_bfr_after (
		.din(new_net_10799),
		.dout(new_net_10800)
	);

	bfr new_net_10801_bfr_after (
		.din(new_net_10800),
		.dout(new_net_10801)
	);

	bfr new_net_10802_bfr_after (
		.din(new_net_10801),
		.dout(new_net_10802)
	);

	bfr new_net_10803_bfr_after (
		.din(new_net_10802),
		.dout(new_net_10803)
	);

	bfr new_net_10804_bfr_after (
		.din(new_net_10803),
		.dout(new_net_10804)
	);

	bfr new_net_10805_bfr_after (
		.din(new_net_10804),
		.dout(new_net_10805)
	);

	bfr new_net_10806_bfr_after (
		.din(new_net_10805),
		.dout(new_net_10806)
	);

	bfr new_net_10807_bfr_after (
		.din(new_net_10806),
		.dout(new_net_10807)
	);

	bfr new_net_10808_bfr_after (
		.din(new_net_10807),
		.dout(new_net_10808)
	);

	bfr new_net_10809_bfr_after (
		.din(new_net_10808),
		.dout(new_net_10809)
	);

	bfr new_net_10810_bfr_after (
		.din(new_net_10809),
		.dout(new_net_10810)
	);

	bfr new_net_10811_bfr_after (
		.din(new_net_10810),
		.dout(new_net_10811)
	);

	bfr new_net_10812_bfr_after (
		.din(new_net_10811),
		.dout(new_net_10812)
	);

	bfr new_net_10813_bfr_after (
		.din(new_net_10812),
		.dout(new_net_10813)
	);

	bfr new_net_10814_bfr_after (
		.din(new_net_10813),
		.dout(new_net_10814)
	);

	bfr new_net_10815_bfr_after (
		.din(new_net_10814),
		.dout(new_net_10815)
	);

	bfr new_net_10816_bfr_after (
		.din(new_net_10815),
		.dout(new_net_10816)
	);

	bfr new_net_10817_bfr_after (
		.din(new_net_10816),
		.dout(new_net_10817)
	);

	bfr new_net_10818_bfr_after (
		.din(new_net_10817),
		.dout(new_net_10818)
	);

	bfr new_net_10819_bfr_after (
		.din(new_net_10818),
		.dout(new_net_10819)
	);

	bfr new_net_10820_bfr_after (
		.din(new_net_10819),
		.dout(new_net_10820)
	);

	bfr new_net_10821_bfr_after (
		.din(new_net_10820),
		.dout(new_net_10821)
	);

	bfr new_net_10822_bfr_after (
		.din(new_net_10821),
		.dout(new_net_10822)
	);

	bfr new_net_10823_bfr_after (
		.din(new_net_10822),
		.dout(new_net_10823)
	);

	bfr new_net_10824_bfr_after (
		.din(new_net_10823),
		.dout(new_net_10824)
	);

	bfr new_net_10825_bfr_after (
		.din(new_net_10824),
		.dout(new_net_10825)
	);

	bfr new_net_10826_bfr_after (
		.din(new_net_10825),
		.dout(new_net_10826)
	);

	spl2 _1823__v_fanout (
		.a(new_net_10826),
		.b(new_net_18),
		.c(new_net_19)
	);

	bfr new_net_10827_bfr_after (
		.din(_0011_),
		.dout(new_net_10827)
	);

	bfr new_net_10828_bfr_after (
		.din(new_net_10827),
		.dout(new_net_10828)
	);

	bfr new_net_10829_bfr_after (
		.din(new_net_10828),
		.dout(new_net_10829)
	);

	bfr new_net_10830_bfr_after (
		.din(new_net_10829),
		.dout(new_net_10830)
	);

	bfr new_net_10831_bfr_after (
		.din(new_net_10830),
		.dout(new_net_10831)
	);

	bfr new_net_10832_bfr_after (
		.din(new_net_10831),
		.dout(new_net_10832)
	);

	bfr new_net_10833_bfr_after (
		.din(new_net_10832),
		.dout(new_net_10833)
	);

	bfr new_net_10834_bfr_after (
		.din(new_net_10833),
		.dout(new_net_10834)
	);

	bfr new_net_10835_bfr_after (
		.din(new_net_10834),
		.dout(new_net_10835)
	);

	bfr new_net_10836_bfr_after (
		.din(new_net_10835),
		.dout(new_net_10836)
	);

	bfr new_net_10837_bfr_after (
		.din(new_net_10836),
		.dout(new_net_10837)
	);

	bfr new_net_10838_bfr_after (
		.din(new_net_10837),
		.dout(new_net_10838)
	);

	bfr new_net_10839_bfr_after (
		.din(new_net_10838),
		.dout(new_net_10839)
	);

	bfr new_net_10840_bfr_after (
		.din(new_net_10839),
		.dout(new_net_10840)
	);

	bfr new_net_10841_bfr_after (
		.din(new_net_10840),
		.dout(new_net_10841)
	);

	bfr new_net_10842_bfr_after (
		.din(new_net_10841),
		.dout(new_net_10842)
	);

	spl2 _0011__v_fanout (
		.a(new_net_10842),
		.b(new_net_3226),
		.c(new_net_3227)
	);

	bfr new_net_10843_bfr_after (
		.din(_1811_),
		.dout(new_net_10843)
	);

	bfr new_net_10844_bfr_after (
		.din(new_net_10843),
		.dout(new_net_10844)
	);

	bfr new_net_10845_bfr_after (
		.din(new_net_10844),
		.dout(new_net_10845)
	);

	bfr new_net_10846_bfr_after (
		.din(new_net_10845),
		.dout(new_net_10846)
	);

	bfr new_net_10847_bfr_after (
		.din(new_net_10846),
		.dout(new_net_10847)
	);

	bfr new_net_10848_bfr_after (
		.din(new_net_10847),
		.dout(new_net_10848)
	);

	bfr new_net_10849_bfr_after (
		.din(new_net_10848),
		.dout(new_net_10849)
	);

	bfr new_net_10850_bfr_after (
		.din(new_net_10849),
		.dout(new_net_10850)
	);

	bfr new_net_10851_bfr_after (
		.din(new_net_10850),
		.dout(new_net_10851)
	);

	bfr new_net_10852_bfr_after (
		.din(new_net_10851),
		.dout(new_net_10852)
	);

	bfr new_net_10853_bfr_after (
		.din(new_net_10852),
		.dout(new_net_10853)
	);

	bfr new_net_10854_bfr_after (
		.din(new_net_10853),
		.dout(new_net_10854)
	);

	bfr new_net_10855_bfr_after (
		.din(new_net_10854),
		.dout(new_net_10855)
	);

	bfr new_net_10856_bfr_after (
		.din(new_net_10855),
		.dout(new_net_10856)
	);

	bfr new_net_10857_bfr_after (
		.din(new_net_10856),
		.dout(new_net_10857)
	);

	bfr new_net_10858_bfr_after (
		.din(new_net_10857),
		.dout(new_net_10858)
	);

	bfr new_net_10859_bfr_after (
		.din(new_net_10858),
		.dout(new_net_10859)
	);

	bfr new_net_10860_bfr_after (
		.din(new_net_10859),
		.dout(new_net_10860)
	);

	bfr new_net_10861_bfr_after (
		.din(new_net_10860),
		.dout(new_net_10861)
	);

	bfr new_net_10862_bfr_after (
		.din(new_net_10861),
		.dout(new_net_10862)
	);

	bfr new_net_10863_bfr_after (
		.din(new_net_10862),
		.dout(new_net_10863)
	);

	bfr new_net_10864_bfr_after (
		.din(new_net_10863),
		.dout(new_net_10864)
	);

	bfr new_net_10865_bfr_after (
		.din(new_net_10864),
		.dout(new_net_10865)
	);

	bfr new_net_10866_bfr_after (
		.din(new_net_10865),
		.dout(new_net_10866)
	);

	bfr new_net_10867_bfr_after (
		.din(new_net_10866),
		.dout(new_net_10867)
	);

	bfr new_net_10868_bfr_after (
		.din(new_net_10867),
		.dout(new_net_10868)
	);

	bfr new_net_10869_bfr_after (
		.din(new_net_10868),
		.dout(new_net_10869)
	);

	bfr new_net_10870_bfr_after (
		.din(new_net_10869),
		.dout(new_net_10870)
	);

	bfr new_net_10871_bfr_after (
		.din(new_net_10870),
		.dout(new_net_10871)
	);

	bfr new_net_10872_bfr_after (
		.din(new_net_10871),
		.dout(new_net_10872)
	);

	bfr new_net_10873_bfr_after (
		.din(new_net_10872),
		.dout(new_net_10873)
	);

	bfr new_net_10874_bfr_after (
		.din(new_net_10873),
		.dout(new_net_10874)
	);

	bfr new_net_10875_bfr_after (
		.din(new_net_10874),
		.dout(new_net_10875)
	);

	bfr new_net_10876_bfr_after (
		.din(new_net_10875),
		.dout(new_net_10876)
	);

	bfr new_net_10877_bfr_after (
		.din(new_net_10876),
		.dout(new_net_10877)
	);

	bfr new_net_10878_bfr_after (
		.din(new_net_10877),
		.dout(new_net_10878)
	);

	bfr new_net_10879_bfr_after (
		.din(new_net_10878),
		.dout(new_net_10879)
	);

	bfr new_net_10880_bfr_after (
		.din(new_net_10879),
		.dout(new_net_10880)
	);

	bfr new_net_10881_bfr_after (
		.din(new_net_10880),
		.dout(new_net_10881)
	);

	bfr new_net_10882_bfr_after (
		.din(new_net_10881),
		.dout(new_net_10882)
	);

	bfr new_net_10883_bfr_after (
		.din(new_net_10882),
		.dout(new_net_10883)
	);

	bfr new_net_10884_bfr_after (
		.din(new_net_10883),
		.dout(new_net_10884)
	);

	bfr new_net_10885_bfr_after (
		.din(new_net_10884),
		.dout(new_net_10885)
	);

	bfr new_net_10886_bfr_after (
		.din(new_net_10885),
		.dout(new_net_10886)
	);

	bfr new_net_10887_bfr_after (
		.din(new_net_10886),
		.dout(new_net_10887)
	);

	bfr new_net_10888_bfr_after (
		.din(new_net_10887),
		.dout(new_net_10888)
	);

	bfr new_net_10889_bfr_after (
		.din(new_net_10888),
		.dout(new_net_10889)
	);

	bfr new_net_10890_bfr_after (
		.din(new_net_10889),
		.dout(new_net_10890)
	);

	bfr new_net_10891_bfr_after (
		.din(new_net_10890),
		.dout(new_net_10891)
	);

	bfr new_net_10892_bfr_after (
		.din(new_net_10891),
		.dout(new_net_10892)
	);

	bfr new_net_10893_bfr_after (
		.din(new_net_10892),
		.dout(new_net_10893)
	);

	bfr new_net_10894_bfr_after (
		.din(new_net_10893),
		.dout(new_net_10894)
	);

	bfr new_net_10895_bfr_after (
		.din(new_net_10894),
		.dout(new_net_10895)
	);

	bfr new_net_10896_bfr_after (
		.din(new_net_10895),
		.dout(new_net_10896)
	);

	bfr new_net_10897_bfr_after (
		.din(new_net_10896),
		.dout(new_net_10897)
	);

	bfr new_net_10898_bfr_after (
		.din(new_net_10897),
		.dout(new_net_10898)
	);

	bfr new_net_10899_bfr_after (
		.din(new_net_10898),
		.dout(new_net_10899)
	);

	bfr new_net_10900_bfr_after (
		.din(new_net_10899),
		.dout(new_net_10900)
	);

	bfr new_net_10901_bfr_after (
		.din(new_net_10900),
		.dout(new_net_10901)
	);

	bfr new_net_10902_bfr_after (
		.din(new_net_10901),
		.dout(new_net_10902)
	);

	bfr new_net_10903_bfr_after (
		.din(new_net_10902),
		.dout(new_net_10903)
	);

	bfr new_net_10904_bfr_after (
		.din(new_net_10903),
		.dout(new_net_10904)
	);

	bfr new_net_10905_bfr_after (
		.din(new_net_10904),
		.dout(new_net_10905)
	);

	bfr new_net_10906_bfr_after (
		.din(new_net_10905),
		.dout(new_net_10906)
	);

	bfr new_net_10907_bfr_after (
		.din(new_net_10906),
		.dout(new_net_10907)
	);

	bfr new_net_10908_bfr_after (
		.din(new_net_10907),
		.dout(new_net_10908)
	);

	bfr new_net_10909_bfr_after (
		.din(new_net_10908),
		.dout(new_net_10909)
	);

	bfr new_net_10910_bfr_after (
		.din(new_net_10909),
		.dout(new_net_10910)
	);

	bfr new_net_10911_bfr_after (
		.din(new_net_10910),
		.dout(new_net_10911)
	);

	bfr new_net_10912_bfr_after (
		.din(new_net_10911),
		.dout(new_net_10912)
	);

	bfr new_net_10913_bfr_after (
		.din(new_net_10912),
		.dout(new_net_10913)
	);

	bfr new_net_10914_bfr_after (
		.din(new_net_10913),
		.dout(new_net_10914)
	);

	bfr new_net_10915_bfr_after (
		.din(new_net_10914),
		.dout(new_net_10915)
	);

	bfr new_net_10916_bfr_after (
		.din(new_net_10915),
		.dout(new_net_10916)
	);

	bfr new_net_10917_bfr_after (
		.din(new_net_10916),
		.dout(new_net_10917)
	);

	bfr new_net_10918_bfr_after (
		.din(new_net_10917),
		.dout(new_net_10918)
	);

	bfr new_net_10919_bfr_after (
		.din(new_net_10918),
		.dout(new_net_10919)
	);

	bfr new_net_10920_bfr_after (
		.din(new_net_10919),
		.dout(new_net_10920)
	);

	bfr new_net_10921_bfr_after (
		.din(new_net_10920),
		.dout(new_net_10921)
	);

	bfr new_net_10922_bfr_after (
		.din(new_net_10921),
		.dout(new_net_10922)
	);

	spl2 _1811__v_fanout (
		.a(new_net_10922),
		.b(new_net_218),
		.c(new_net_219)
	);

	bfr new_net_10923_bfr_after (
		.din(_0544_),
		.dout(new_net_10923)
	);

	bfr new_net_10924_bfr_after (
		.din(new_net_10923),
		.dout(new_net_10924)
	);

	bfr new_net_10925_bfr_after (
		.din(new_net_10924),
		.dout(new_net_10925)
	);

	bfr new_net_10926_bfr_after (
		.din(new_net_10925),
		.dout(new_net_10926)
	);

	bfr new_net_10927_bfr_after (
		.din(new_net_10926),
		.dout(new_net_10927)
	);

	bfr new_net_10928_bfr_after (
		.din(new_net_10927),
		.dout(new_net_10928)
	);

	bfr new_net_10929_bfr_after (
		.din(new_net_10928),
		.dout(new_net_10929)
	);

	bfr new_net_10930_bfr_after (
		.din(new_net_10929),
		.dout(new_net_10930)
	);

	bfr new_net_10931_bfr_after (
		.din(new_net_10930),
		.dout(new_net_10931)
	);

	bfr new_net_10932_bfr_after (
		.din(new_net_10931),
		.dout(new_net_10932)
	);

	bfr new_net_10933_bfr_after (
		.din(new_net_10932),
		.dout(new_net_10933)
	);

	bfr new_net_10934_bfr_after (
		.din(new_net_10933),
		.dout(new_net_10934)
	);

	bfr new_net_10935_bfr_after (
		.din(new_net_10934),
		.dout(new_net_10935)
	);

	bfr new_net_10936_bfr_after (
		.din(new_net_10935),
		.dout(new_net_10936)
	);

	bfr new_net_10937_bfr_after (
		.din(new_net_10936),
		.dout(new_net_10937)
	);

	bfr new_net_10938_bfr_after (
		.din(new_net_10937),
		.dout(new_net_10938)
	);

	bfr new_net_10939_bfr_after (
		.din(new_net_10938),
		.dout(new_net_10939)
	);

	bfr new_net_10940_bfr_after (
		.din(new_net_10939),
		.dout(new_net_10940)
	);

	bfr new_net_10941_bfr_after (
		.din(new_net_10940),
		.dout(new_net_10941)
	);

	bfr new_net_10942_bfr_after (
		.din(new_net_10941),
		.dout(new_net_10942)
	);

	bfr new_net_10943_bfr_after (
		.din(new_net_10942),
		.dout(new_net_10943)
	);

	bfr new_net_10944_bfr_after (
		.din(new_net_10943),
		.dout(new_net_10944)
	);

	bfr new_net_10945_bfr_after (
		.din(new_net_10944),
		.dout(new_net_10945)
	);

	bfr new_net_10946_bfr_after (
		.din(new_net_10945),
		.dout(new_net_10946)
	);

	bfr new_net_10947_bfr_after (
		.din(new_net_10946),
		.dout(new_net_10947)
	);

	bfr new_net_10948_bfr_after (
		.din(new_net_10947),
		.dout(new_net_10948)
	);

	bfr new_net_10949_bfr_after (
		.din(new_net_10948),
		.dout(new_net_10949)
	);

	bfr new_net_10950_bfr_after (
		.din(new_net_10949),
		.dout(new_net_10950)
	);

	bfr new_net_10951_bfr_after (
		.din(new_net_10950),
		.dout(new_net_10951)
	);

	bfr new_net_10952_bfr_after (
		.din(new_net_10951),
		.dout(new_net_10952)
	);

	bfr new_net_10953_bfr_after (
		.din(new_net_10952),
		.dout(new_net_10953)
	);

	bfr new_net_10954_bfr_after (
		.din(new_net_10953),
		.dout(new_net_10954)
	);

	bfr new_net_10955_bfr_after (
		.din(new_net_10954),
		.dout(new_net_10955)
	);

	bfr new_net_10956_bfr_after (
		.din(new_net_10955),
		.dout(new_net_10956)
	);

	bfr new_net_10957_bfr_after (
		.din(new_net_10956),
		.dout(new_net_10957)
	);

	bfr new_net_10958_bfr_after (
		.din(new_net_10957),
		.dout(new_net_10958)
	);

	bfr new_net_10959_bfr_after (
		.din(new_net_10958),
		.dout(new_net_10959)
	);

	bfr new_net_10960_bfr_after (
		.din(new_net_10959),
		.dout(new_net_10960)
	);

	bfr new_net_10961_bfr_after (
		.din(new_net_10960),
		.dout(new_net_10961)
	);

	bfr new_net_10962_bfr_after (
		.din(new_net_10961),
		.dout(new_net_10962)
	);

	bfr new_net_10963_bfr_after (
		.din(new_net_10962),
		.dout(new_net_10963)
	);

	bfr new_net_10964_bfr_after (
		.din(new_net_10963),
		.dout(new_net_10964)
	);

	bfr new_net_10965_bfr_after (
		.din(new_net_10964),
		.dout(new_net_10965)
	);

	bfr new_net_10966_bfr_after (
		.din(new_net_10965),
		.dout(new_net_10966)
	);

	bfr new_net_10967_bfr_after (
		.din(new_net_10966),
		.dout(new_net_10967)
	);

	bfr new_net_10968_bfr_after (
		.din(new_net_10967),
		.dout(new_net_10968)
	);

	bfr new_net_10969_bfr_after (
		.din(new_net_10968),
		.dout(new_net_10969)
	);

	bfr new_net_10970_bfr_after (
		.din(new_net_10969),
		.dout(new_net_10970)
	);

	bfr new_net_10971_bfr_after (
		.din(new_net_10970),
		.dout(new_net_10971)
	);

	bfr new_net_10972_bfr_after (
		.din(new_net_10971),
		.dout(new_net_10972)
	);

	bfr new_net_10973_bfr_after (
		.din(new_net_10972),
		.dout(new_net_10973)
	);

	bfr new_net_10974_bfr_after (
		.din(new_net_10973),
		.dout(new_net_10974)
	);

	bfr new_net_10975_bfr_after (
		.din(new_net_10974),
		.dout(new_net_10975)
	);

	bfr new_net_10976_bfr_after (
		.din(new_net_10975),
		.dout(new_net_10976)
	);

	spl2 _0544__v_fanout (
		.a(new_net_10976),
		.b(new_net_2444),
		.c(new_net_2445)
	);

	bfr new_net_10977_bfr_after (
		.din(_0436_),
		.dout(new_net_10977)
	);

	bfr new_net_10978_bfr_after (
		.din(new_net_10977),
		.dout(new_net_10978)
	);

	bfr new_net_10979_bfr_after (
		.din(new_net_10978),
		.dout(new_net_10979)
	);

	bfr new_net_10980_bfr_after (
		.din(new_net_10979),
		.dout(new_net_10980)
	);

	bfr new_net_10981_bfr_after (
		.din(new_net_10980),
		.dout(new_net_10981)
	);

	bfr new_net_10982_bfr_after (
		.din(new_net_10981),
		.dout(new_net_10982)
	);

	bfr new_net_10983_bfr_after (
		.din(new_net_10982),
		.dout(new_net_10983)
	);

	bfr new_net_10984_bfr_after (
		.din(new_net_10983),
		.dout(new_net_10984)
	);

	bfr new_net_10985_bfr_after (
		.din(new_net_10984),
		.dout(new_net_10985)
	);

	bfr new_net_10986_bfr_after (
		.din(new_net_10985),
		.dout(new_net_10986)
	);

	bfr new_net_10987_bfr_after (
		.din(new_net_10986),
		.dout(new_net_10987)
	);

	bfr new_net_10988_bfr_after (
		.din(new_net_10987),
		.dout(new_net_10988)
	);

	bfr new_net_10989_bfr_after (
		.din(new_net_10988),
		.dout(new_net_10989)
	);

	bfr new_net_10990_bfr_after (
		.din(new_net_10989),
		.dout(new_net_10990)
	);

	bfr new_net_10991_bfr_after (
		.din(new_net_10990),
		.dout(new_net_10991)
	);

	bfr new_net_10992_bfr_after (
		.din(new_net_10991),
		.dout(new_net_10992)
	);

	bfr new_net_10993_bfr_after (
		.din(new_net_10992),
		.dout(new_net_10993)
	);

	bfr new_net_10994_bfr_after (
		.din(new_net_10993),
		.dout(new_net_10994)
	);

	bfr new_net_10995_bfr_after (
		.din(new_net_10994),
		.dout(new_net_10995)
	);

	bfr new_net_10996_bfr_after (
		.din(new_net_10995),
		.dout(new_net_10996)
	);

	bfr new_net_10997_bfr_after (
		.din(new_net_10996),
		.dout(new_net_10997)
	);

	bfr new_net_10998_bfr_after (
		.din(new_net_10997),
		.dout(new_net_10998)
	);

	bfr new_net_10999_bfr_after (
		.din(new_net_10998),
		.dout(new_net_10999)
	);

	bfr new_net_11000_bfr_after (
		.din(new_net_10999),
		.dout(new_net_11000)
	);

	bfr new_net_11001_bfr_after (
		.din(new_net_11000),
		.dout(new_net_11001)
	);

	bfr new_net_11002_bfr_after (
		.din(new_net_11001),
		.dout(new_net_11002)
	);

	bfr new_net_11003_bfr_after (
		.din(new_net_11002),
		.dout(new_net_11003)
	);

	bfr new_net_11004_bfr_after (
		.din(new_net_11003),
		.dout(new_net_11004)
	);

	bfr new_net_11005_bfr_after (
		.din(new_net_11004),
		.dout(new_net_11005)
	);

	bfr new_net_11006_bfr_after (
		.din(new_net_11005),
		.dout(new_net_11006)
	);

	bfr new_net_11007_bfr_after (
		.din(new_net_11006),
		.dout(new_net_11007)
	);

	bfr new_net_11008_bfr_after (
		.din(new_net_11007),
		.dout(new_net_11008)
	);

	bfr new_net_11009_bfr_after (
		.din(new_net_11008),
		.dout(new_net_11009)
	);

	bfr new_net_11010_bfr_after (
		.din(new_net_11009),
		.dout(new_net_11010)
	);

	bfr new_net_11011_bfr_after (
		.din(new_net_11010),
		.dout(new_net_11011)
	);

	bfr new_net_11012_bfr_after (
		.din(new_net_11011),
		.dout(new_net_11012)
	);

	bfr new_net_11013_bfr_after (
		.din(new_net_11012),
		.dout(new_net_11013)
	);

	bfr new_net_11014_bfr_after (
		.din(new_net_11013),
		.dout(new_net_11014)
	);

	bfr new_net_11015_bfr_after (
		.din(new_net_11014),
		.dout(new_net_11015)
	);

	bfr new_net_11016_bfr_after (
		.din(new_net_11015),
		.dout(new_net_11016)
	);

	bfr new_net_11017_bfr_after (
		.din(new_net_11016),
		.dout(new_net_11017)
	);

	bfr new_net_11018_bfr_after (
		.din(new_net_11017),
		.dout(new_net_11018)
	);

	bfr new_net_11019_bfr_after (
		.din(new_net_11018),
		.dout(new_net_11019)
	);

	bfr new_net_11020_bfr_after (
		.din(new_net_11019),
		.dout(new_net_11020)
	);

	bfr new_net_11021_bfr_after (
		.din(new_net_11020),
		.dout(new_net_11021)
	);

	bfr new_net_11022_bfr_after (
		.din(new_net_11021),
		.dout(new_net_11022)
	);

	bfr new_net_11023_bfr_after (
		.din(new_net_11022),
		.dout(new_net_11023)
	);

	bfr new_net_11024_bfr_after (
		.din(new_net_11023),
		.dout(new_net_11024)
	);

	bfr new_net_11025_bfr_after (
		.din(new_net_11024),
		.dout(new_net_11025)
	);

	bfr new_net_11026_bfr_after (
		.din(new_net_11025),
		.dout(new_net_11026)
	);

	bfr new_net_11027_bfr_after (
		.din(new_net_11026),
		.dout(new_net_11027)
	);

	bfr new_net_11028_bfr_after (
		.din(new_net_11027),
		.dout(new_net_11028)
	);

	bfr new_net_11029_bfr_after (
		.din(new_net_11028),
		.dout(new_net_11029)
	);

	bfr new_net_11030_bfr_after (
		.din(new_net_11029),
		.dout(new_net_11030)
	);

	bfr new_net_11031_bfr_after (
		.din(new_net_11030),
		.dout(new_net_11031)
	);

	bfr new_net_11032_bfr_after (
		.din(new_net_11031),
		.dout(new_net_11032)
	);

	bfr new_net_11033_bfr_after (
		.din(new_net_11032),
		.dout(new_net_11033)
	);

	bfr new_net_11034_bfr_after (
		.din(new_net_11033),
		.dout(new_net_11034)
	);

	bfr new_net_11035_bfr_after (
		.din(new_net_11034),
		.dout(new_net_11035)
	);

	bfr new_net_11036_bfr_after (
		.din(new_net_11035),
		.dout(new_net_11036)
	);

	bfr new_net_11037_bfr_after (
		.din(new_net_11036),
		.dout(new_net_11037)
	);

	bfr new_net_11038_bfr_after (
		.din(new_net_11037),
		.dout(new_net_11038)
	);

	bfr new_net_11039_bfr_after (
		.din(new_net_11038),
		.dout(new_net_11039)
	);

	bfr new_net_11040_bfr_after (
		.din(new_net_11039),
		.dout(new_net_11040)
	);

	bfr new_net_11041_bfr_after (
		.din(new_net_11040),
		.dout(new_net_11041)
	);

	bfr new_net_11042_bfr_after (
		.din(new_net_11041),
		.dout(new_net_11042)
	);

	bfr new_net_11043_bfr_after (
		.din(new_net_11042),
		.dout(new_net_11043)
	);

	bfr new_net_11044_bfr_after (
		.din(new_net_11043),
		.dout(new_net_11044)
	);

	bfr new_net_11045_bfr_after (
		.din(new_net_11044),
		.dout(new_net_11045)
	);

	bfr new_net_11046_bfr_after (
		.din(new_net_11045),
		.dout(new_net_11046)
	);

	bfr new_net_11047_bfr_after (
		.din(new_net_11046),
		.dout(new_net_11047)
	);

	bfr new_net_11048_bfr_after (
		.din(new_net_11047),
		.dout(new_net_11048)
	);

	bfr new_net_11049_bfr_after (
		.din(new_net_11048),
		.dout(new_net_11049)
	);

	bfr new_net_11050_bfr_after (
		.din(new_net_11049),
		.dout(new_net_11050)
	);

	bfr new_net_11051_bfr_after (
		.din(new_net_11050),
		.dout(new_net_11051)
	);

	bfr new_net_11052_bfr_after (
		.din(new_net_11051),
		.dout(new_net_11052)
	);

	bfr new_net_11053_bfr_after (
		.din(new_net_11052),
		.dout(new_net_11053)
	);

	bfr new_net_11054_bfr_after (
		.din(new_net_11053),
		.dout(new_net_11054)
	);

	bfr new_net_11055_bfr_after (
		.din(new_net_11054),
		.dout(new_net_11055)
	);

	bfr new_net_11056_bfr_after (
		.din(new_net_11055),
		.dout(new_net_11056)
	);

	bfr new_net_11057_bfr_after (
		.din(new_net_11056),
		.dout(new_net_11057)
	);

	bfr new_net_11058_bfr_after (
		.din(new_net_11057),
		.dout(new_net_11058)
	);

	bfr new_net_11059_bfr_after (
		.din(new_net_11058),
		.dout(new_net_11059)
	);

	bfr new_net_11060_bfr_after (
		.din(new_net_11059),
		.dout(new_net_11060)
	);

	bfr new_net_11061_bfr_after (
		.din(new_net_11060),
		.dout(new_net_11061)
	);

	bfr new_net_11062_bfr_after (
		.din(new_net_11061),
		.dout(new_net_11062)
	);

	bfr new_net_11063_bfr_after (
		.din(new_net_11062),
		.dout(new_net_11063)
	);

	bfr new_net_11064_bfr_after (
		.din(new_net_11063),
		.dout(new_net_11064)
	);

	bfr new_net_11065_bfr_after (
		.din(new_net_11064),
		.dout(new_net_11065)
	);

	bfr new_net_11066_bfr_after (
		.din(new_net_11065),
		.dout(new_net_11066)
	);

	bfr new_net_11067_bfr_after (
		.din(new_net_11066),
		.dout(new_net_11067)
	);

	bfr new_net_11068_bfr_after (
		.din(new_net_11067),
		.dout(new_net_11068)
	);

	bfr new_net_11069_bfr_after (
		.din(new_net_11068),
		.dout(new_net_11069)
	);

	bfr new_net_11070_bfr_after (
		.din(new_net_11069),
		.dout(new_net_11070)
	);

	bfr new_net_11071_bfr_after (
		.din(new_net_11070),
		.dout(new_net_11071)
	);

	bfr new_net_11072_bfr_after (
		.din(new_net_11071),
		.dout(new_net_11072)
	);

	spl2 _0436__v_fanout (
		.a(new_net_11072),
		.b(new_net_106),
		.c(new_net_107)
	);

	bfr new_net_11073_bfr_after (
		.din(_0102_),
		.dout(new_net_11073)
	);

	bfr new_net_11074_bfr_after (
		.din(new_net_11073),
		.dout(new_net_11074)
	);

	bfr new_net_11075_bfr_after (
		.din(new_net_11074),
		.dout(new_net_11075)
	);

	bfr new_net_11076_bfr_after (
		.din(new_net_11075),
		.dout(new_net_11076)
	);

	bfr new_net_11077_bfr_after (
		.din(new_net_11076),
		.dout(new_net_11077)
	);

	bfr new_net_11078_bfr_after (
		.din(new_net_11077),
		.dout(new_net_11078)
	);

	bfr new_net_11079_bfr_after (
		.din(new_net_11078),
		.dout(new_net_11079)
	);

	bfr new_net_11080_bfr_after (
		.din(new_net_11079),
		.dout(new_net_11080)
	);

	bfr new_net_11081_bfr_after (
		.din(new_net_11080),
		.dout(new_net_11081)
	);

	bfr new_net_11082_bfr_after (
		.din(new_net_11081),
		.dout(new_net_11082)
	);

	bfr new_net_11083_bfr_after (
		.din(new_net_11082),
		.dout(new_net_11083)
	);

	bfr new_net_11084_bfr_after (
		.din(new_net_11083),
		.dout(new_net_11084)
	);

	bfr new_net_11085_bfr_after (
		.din(new_net_11084),
		.dout(new_net_11085)
	);

	bfr new_net_11086_bfr_after (
		.din(new_net_11085),
		.dout(new_net_11086)
	);

	bfr new_net_11087_bfr_after (
		.din(new_net_11086),
		.dout(new_net_11087)
	);

	bfr new_net_11088_bfr_after (
		.din(new_net_11087),
		.dout(new_net_11088)
	);

	bfr new_net_11089_bfr_after (
		.din(new_net_11088),
		.dout(new_net_11089)
	);

	bfr new_net_11090_bfr_after (
		.din(new_net_11089),
		.dout(new_net_11090)
	);

	bfr new_net_11091_bfr_after (
		.din(new_net_11090),
		.dout(new_net_11091)
	);

	bfr new_net_11092_bfr_after (
		.din(new_net_11091),
		.dout(new_net_11092)
	);

	bfr new_net_11093_bfr_after (
		.din(new_net_11092),
		.dout(new_net_11093)
	);

	bfr new_net_11094_bfr_after (
		.din(new_net_11093),
		.dout(new_net_11094)
	);

	bfr new_net_11095_bfr_after (
		.din(new_net_11094),
		.dout(new_net_11095)
	);

	bfr new_net_11096_bfr_after (
		.din(new_net_11095),
		.dout(new_net_11096)
	);

	bfr new_net_11097_bfr_after (
		.din(new_net_11096),
		.dout(new_net_11097)
	);

	bfr new_net_11098_bfr_after (
		.din(new_net_11097),
		.dout(new_net_11098)
	);

	bfr new_net_11099_bfr_after (
		.din(new_net_11098),
		.dout(new_net_11099)
	);

	bfr new_net_11100_bfr_after (
		.din(new_net_11099),
		.dout(new_net_11100)
	);

	bfr new_net_11101_bfr_after (
		.din(new_net_11100),
		.dout(new_net_11101)
	);

	bfr new_net_11102_bfr_after (
		.din(new_net_11101),
		.dout(new_net_11102)
	);

	bfr new_net_11103_bfr_after (
		.din(new_net_11102),
		.dout(new_net_11103)
	);

	bfr new_net_11104_bfr_after (
		.din(new_net_11103),
		.dout(new_net_11104)
	);

	bfr new_net_11105_bfr_after (
		.din(new_net_11104),
		.dout(new_net_11105)
	);

	bfr new_net_11106_bfr_after (
		.din(new_net_11105),
		.dout(new_net_11106)
	);

	bfr new_net_11107_bfr_after (
		.din(new_net_11106),
		.dout(new_net_11107)
	);

	bfr new_net_11108_bfr_after (
		.din(new_net_11107),
		.dout(new_net_11108)
	);

	bfr new_net_11109_bfr_after (
		.din(new_net_11108),
		.dout(new_net_11109)
	);

	bfr new_net_11110_bfr_after (
		.din(new_net_11109),
		.dout(new_net_11110)
	);

	bfr new_net_11111_bfr_after (
		.din(new_net_11110),
		.dout(new_net_11111)
	);

	bfr new_net_11112_bfr_after (
		.din(new_net_11111),
		.dout(new_net_11112)
	);

	bfr new_net_11113_bfr_after (
		.din(new_net_11112),
		.dout(new_net_11113)
	);

	bfr new_net_11114_bfr_after (
		.din(new_net_11113),
		.dout(new_net_11114)
	);

	bfr new_net_11115_bfr_after (
		.din(new_net_11114),
		.dout(new_net_11115)
	);

	bfr new_net_11116_bfr_after (
		.din(new_net_11115),
		.dout(new_net_11116)
	);

	bfr new_net_11117_bfr_after (
		.din(new_net_11116),
		.dout(new_net_11117)
	);

	bfr new_net_11118_bfr_after (
		.din(new_net_11117),
		.dout(new_net_11118)
	);

	bfr new_net_11119_bfr_after (
		.din(new_net_11118),
		.dout(new_net_11119)
	);

	bfr new_net_11120_bfr_after (
		.din(new_net_11119),
		.dout(new_net_11120)
	);

	spl2 _0102__v_fanout (
		.a(new_net_11120),
		.b(new_net_1736),
		.c(new_net_1737)
	);

	bfr new_net_11121_bfr_after (
		.din(_0542_),
		.dout(new_net_11121)
	);

	bfr new_net_11122_bfr_after (
		.din(new_net_11121),
		.dout(new_net_11122)
	);

	bfr new_net_11123_bfr_after (
		.din(new_net_11122),
		.dout(new_net_11123)
	);

	bfr new_net_11124_bfr_after (
		.din(new_net_11123),
		.dout(new_net_11124)
	);

	bfr new_net_11125_bfr_after (
		.din(new_net_11124),
		.dout(new_net_11125)
	);

	bfr new_net_11126_bfr_after (
		.din(new_net_11125),
		.dout(new_net_11126)
	);

	bfr new_net_11127_bfr_after (
		.din(new_net_11126),
		.dout(new_net_11127)
	);

	bfr new_net_11128_bfr_after (
		.din(new_net_11127),
		.dout(new_net_11128)
	);

	bfr new_net_11129_bfr_after (
		.din(new_net_11128),
		.dout(new_net_11129)
	);

	bfr new_net_11130_bfr_after (
		.din(new_net_11129),
		.dout(new_net_11130)
	);

	bfr new_net_11131_bfr_after (
		.din(new_net_11130),
		.dout(new_net_11131)
	);

	bfr new_net_11132_bfr_after (
		.din(new_net_11131),
		.dout(new_net_11132)
	);

	bfr new_net_11133_bfr_after (
		.din(new_net_11132),
		.dout(new_net_11133)
	);

	bfr new_net_11134_bfr_after (
		.din(new_net_11133),
		.dout(new_net_11134)
	);

	bfr new_net_11135_bfr_after (
		.din(new_net_11134),
		.dout(new_net_11135)
	);

	bfr new_net_11136_bfr_after (
		.din(new_net_11135),
		.dout(new_net_11136)
	);

	bfr new_net_11137_bfr_after (
		.din(new_net_11136),
		.dout(new_net_11137)
	);

	bfr new_net_11138_bfr_after (
		.din(new_net_11137),
		.dout(new_net_11138)
	);

	bfr new_net_11139_bfr_after (
		.din(new_net_11138),
		.dout(new_net_11139)
	);

	bfr new_net_11140_bfr_after (
		.din(new_net_11139),
		.dout(new_net_11140)
	);

	bfr new_net_11141_bfr_after (
		.din(new_net_11140),
		.dout(new_net_11141)
	);

	bfr new_net_11142_bfr_after (
		.din(new_net_11141),
		.dout(new_net_11142)
	);

	bfr new_net_11143_bfr_after (
		.din(new_net_11142),
		.dout(new_net_11143)
	);

	bfr new_net_11144_bfr_after (
		.din(new_net_11143),
		.dout(new_net_11144)
	);

	bfr new_net_11145_bfr_after (
		.din(new_net_11144),
		.dout(new_net_11145)
	);

	bfr new_net_11146_bfr_after (
		.din(new_net_11145),
		.dout(new_net_11146)
	);

	bfr new_net_11147_bfr_after (
		.din(new_net_11146),
		.dout(new_net_11147)
	);

	bfr new_net_11148_bfr_after (
		.din(new_net_11147),
		.dout(new_net_11148)
	);

	bfr new_net_11149_bfr_after (
		.din(new_net_11148),
		.dout(new_net_11149)
	);

	bfr new_net_11150_bfr_after (
		.din(new_net_11149),
		.dout(new_net_11150)
	);

	bfr new_net_11151_bfr_after (
		.din(new_net_11150),
		.dout(new_net_11151)
	);

	bfr new_net_11152_bfr_after (
		.din(new_net_11151),
		.dout(new_net_11152)
	);

	bfr new_net_11153_bfr_after (
		.din(new_net_11152),
		.dout(new_net_11153)
	);

	bfr new_net_11154_bfr_after (
		.din(new_net_11153),
		.dout(new_net_11154)
	);

	bfr new_net_11155_bfr_after (
		.din(new_net_11154),
		.dout(new_net_11155)
	);

	bfr new_net_11156_bfr_after (
		.din(new_net_11155),
		.dout(new_net_11156)
	);

	bfr new_net_11157_bfr_after (
		.din(new_net_11156),
		.dout(new_net_11157)
	);

	bfr new_net_11158_bfr_after (
		.din(new_net_11157),
		.dout(new_net_11158)
	);

	bfr new_net_11159_bfr_after (
		.din(new_net_11158),
		.dout(new_net_11159)
	);

	bfr new_net_11160_bfr_after (
		.din(new_net_11159),
		.dout(new_net_11160)
	);

	bfr new_net_11161_bfr_after (
		.din(new_net_11160),
		.dout(new_net_11161)
	);

	bfr new_net_11162_bfr_after (
		.din(new_net_11161),
		.dout(new_net_11162)
	);

	bfr new_net_11163_bfr_after (
		.din(new_net_11162),
		.dout(new_net_11163)
	);

	bfr new_net_11164_bfr_after (
		.din(new_net_11163),
		.dout(new_net_11164)
	);

	bfr new_net_11165_bfr_after (
		.din(new_net_11164),
		.dout(new_net_11165)
	);

	bfr new_net_11166_bfr_after (
		.din(new_net_11165),
		.dout(new_net_11166)
	);

	bfr new_net_11167_bfr_after (
		.din(new_net_11166),
		.dout(new_net_11167)
	);

	bfr new_net_11168_bfr_after (
		.din(new_net_11167),
		.dout(new_net_11168)
	);

	bfr new_net_11169_bfr_after (
		.din(new_net_11168),
		.dout(new_net_11169)
	);

	bfr new_net_11170_bfr_after (
		.din(new_net_11169),
		.dout(new_net_11170)
	);

	bfr new_net_11171_bfr_after (
		.din(new_net_11170),
		.dout(new_net_11171)
	);

	bfr new_net_11172_bfr_after (
		.din(new_net_11171),
		.dout(new_net_11172)
	);

	bfr new_net_11173_bfr_after (
		.din(new_net_11172),
		.dout(new_net_11173)
	);

	bfr new_net_11174_bfr_after (
		.din(new_net_11173),
		.dout(new_net_11174)
	);

	bfr new_net_11175_bfr_after (
		.din(new_net_11174),
		.dout(new_net_11175)
	);

	bfr new_net_11176_bfr_after (
		.din(new_net_11175),
		.dout(new_net_11176)
	);

	bfr new_net_11177_bfr_after (
		.din(new_net_11176),
		.dout(new_net_11177)
	);

	bfr new_net_11178_bfr_after (
		.din(new_net_11177),
		.dout(new_net_11178)
	);

	bfr new_net_11179_bfr_after (
		.din(new_net_11178),
		.dout(new_net_11179)
	);

	bfr new_net_11180_bfr_after (
		.din(new_net_11179),
		.dout(new_net_11180)
	);

	bfr new_net_11181_bfr_after (
		.din(new_net_11180),
		.dout(new_net_11181)
	);

	bfr new_net_11182_bfr_after (
		.din(new_net_11181),
		.dout(new_net_11182)
	);

	bfr new_net_11183_bfr_after (
		.din(new_net_11182),
		.dout(new_net_11183)
	);

	bfr new_net_11184_bfr_after (
		.din(new_net_11183),
		.dout(new_net_11184)
	);

	spl2 _0542__v_fanout (
		.a(new_net_11184),
		.b(new_net_2486),
		.c(new_net_2487)
	);

	bfr new_net_11185_bfr_after (
		.din(_0612_),
		.dout(new_net_11185)
	);

	bfr new_net_11186_bfr_after (
		.din(new_net_11185),
		.dout(new_net_11186)
	);

	bfr new_net_11187_bfr_after (
		.din(new_net_11186),
		.dout(new_net_11187)
	);

	bfr new_net_11188_bfr_after (
		.din(new_net_11187),
		.dout(new_net_11188)
	);

	bfr new_net_11189_bfr_after (
		.din(new_net_11188),
		.dout(new_net_11189)
	);

	bfr new_net_11190_bfr_after (
		.din(new_net_11189),
		.dout(new_net_11190)
	);

	bfr new_net_11191_bfr_after (
		.din(new_net_11190),
		.dout(new_net_11191)
	);

	bfr new_net_11192_bfr_after (
		.din(new_net_11191),
		.dout(new_net_11192)
	);

	bfr new_net_11193_bfr_after (
		.din(new_net_11192),
		.dout(new_net_11193)
	);

	bfr new_net_11194_bfr_after (
		.din(new_net_11193),
		.dout(new_net_11194)
	);

	bfr new_net_11195_bfr_after (
		.din(new_net_11194),
		.dout(new_net_11195)
	);

	bfr new_net_11196_bfr_after (
		.din(new_net_11195),
		.dout(new_net_11196)
	);

	bfr new_net_11197_bfr_after (
		.din(new_net_11196),
		.dout(new_net_11197)
	);

	bfr new_net_11198_bfr_after (
		.din(new_net_11197),
		.dout(new_net_11198)
	);

	bfr new_net_11199_bfr_after (
		.din(new_net_11198),
		.dout(new_net_11199)
	);

	bfr new_net_11200_bfr_after (
		.din(new_net_11199),
		.dout(new_net_11200)
	);

	bfr new_net_11201_bfr_after (
		.din(new_net_11200),
		.dout(new_net_11201)
	);

	bfr new_net_11202_bfr_after (
		.din(new_net_11201),
		.dout(new_net_11202)
	);

	bfr new_net_11203_bfr_after (
		.din(new_net_11202),
		.dout(new_net_11203)
	);

	bfr new_net_11204_bfr_after (
		.din(new_net_11203),
		.dout(new_net_11204)
	);

	bfr new_net_11205_bfr_after (
		.din(new_net_11204),
		.dout(new_net_11205)
	);

	bfr new_net_11206_bfr_after (
		.din(new_net_11205),
		.dout(new_net_11206)
	);

	bfr new_net_11207_bfr_after (
		.din(new_net_11206),
		.dout(new_net_11207)
	);

	bfr new_net_11208_bfr_after (
		.din(new_net_11207),
		.dout(new_net_11208)
	);

	bfr new_net_11209_bfr_after (
		.din(new_net_11208),
		.dout(new_net_11209)
	);

	bfr new_net_11210_bfr_after (
		.din(new_net_11209),
		.dout(new_net_11210)
	);

	bfr new_net_11211_bfr_after (
		.din(new_net_11210),
		.dout(new_net_11211)
	);

	bfr new_net_11212_bfr_after (
		.din(new_net_11211),
		.dout(new_net_11212)
	);

	bfr new_net_11213_bfr_after (
		.din(new_net_11212),
		.dout(new_net_11213)
	);

	bfr new_net_11214_bfr_after (
		.din(new_net_11213),
		.dout(new_net_11214)
	);

	bfr new_net_11215_bfr_after (
		.din(new_net_11214),
		.dout(new_net_11215)
	);

	bfr new_net_11216_bfr_after (
		.din(new_net_11215),
		.dout(new_net_11216)
	);

	spl2 _0612__v_fanout (
		.a(new_net_11216),
		.b(new_net_1352),
		.c(new_net_1353)
	);

	bfr new_net_11217_bfr_after (
		.din(_0104_),
		.dout(new_net_11217)
	);

	bfr new_net_11218_bfr_after (
		.din(new_net_11217),
		.dout(new_net_11218)
	);

	bfr new_net_11219_bfr_after (
		.din(new_net_11218),
		.dout(new_net_11219)
	);

	bfr new_net_11220_bfr_after (
		.din(new_net_11219),
		.dout(new_net_11220)
	);

	bfr new_net_11221_bfr_after (
		.din(new_net_11220),
		.dout(new_net_11221)
	);

	bfr new_net_11222_bfr_after (
		.din(new_net_11221),
		.dout(new_net_11222)
	);

	bfr new_net_11223_bfr_after (
		.din(new_net_11222),
		.dout(new_net_11223)
	);

	bfr new_net_11224_bfr_after (
		.din(new_net_11223),
		.dout(new_net_11224)
	);

	bfr new_net_11225_bfr_after (
		.din(new_net_11224),
		.dout(new_net_11225)
	);

	bfr new_net_11226_bfr_after (
		.din(new_net_11225),
		.dout(new_net_11226)
	);

	bfr new_net_11227_bfr_after (
		.din(new_net_11226),
		.dout(new_net_11227)
	);

	bfr new_net_11228_bfr_after (
		.din(new_net_11227),
		.dout(new_net_11228)
	);

	bfr new_net_11229_bfr_after (
		.din(new_net_11228),
		.dout(new_net_11229)
	);

	bfr new_net_11230_bfr_after (
		.din(new_net_11229),
		.dout(new_net_11230)
	);

	bfr new_net_11231_bfr_after (
		.din(new_net_11230),
		.dout(new_net_11231)
	);

	bfr new_net_11232_bfr_after (
		.din(new_net_11231),
		.dout(new_net_11232)
	);

	bfr new_net_11233_bfr_after (
		.din(new_net_11232),
		.dout(new_net_11233)
	);

	bfr new_net_11234_bfr_after (
		.din(new_net_11233),
		.dout(new_net_11234)
	);

	bfr new_net_11235_bfr_after (
		.din(new_net_11234),
		.dout(new_net_11235)
	);

	bfr new_net_11236_bfr_after (
		.din(new_net_11235),
		.dout(new_net_11236)
	);

	bfr new_net_11237_bfr_after (
		.din(new_net_11236),
		.dout(new_net_11237)
	);

	bfr new_net_11238_bfr_after (
		.din(new_net_11237),
		.dout(new_net_11238)
	);

	bfr new_net_11239_bfr_after (
		.din(new_net_11238),
		.dout(new_net_11239)
	);

	bfr new_net_11240_bfr_after (
		.din(new_net_11239),
		.dout(new_net_11240)
	);

	bfr new_net_11241_bfr_after (
		.din(new_net_11240),
		.dout(new_net_11241)
	);

	bfr new_net_11242_bfr_after (
		.din(new_net_11241),
		.dout(new_net_11242)
	);

	bfr new_net_11243_bfr_after (
		.din(new_net_11242),
		.dout(new_net_11243)
	);

	bfr new_net_11244_bfr_after (
		.din(new_net_11243),
		.dout(new_net_11244)
	);

	bfr new_net_11245_bfr_after (
		.din(new_net_11244),
		.dout(new_net_11245)
	);

	bfr new_net_11246_bfr_after (
		.din(new_net_11245),
		.dout(new_net_11246)
	);

	bfr new_net_11247_bfr_after (
		.din(new_net_11246),
		.dout(new_net_11247)
	);

	bfr new_net_11248_bfr_after (
		.din(new_net_11247),
		.dout(new_net_11248)
	);

	bfr new_net_11249_bfr_after (
		.din(new_net_11248),
		.dout(new_net_11249)
	);

	bfr new_net_11250_bfr_after (
		.din(new_net_11249),
		.dout(new_net_11250)
	);

	bfr new_net_11251_bfr_after (
		.din(new_net_11250),
		.dout(new_net_11251)
	);

	bfr new_net_11252_bfr_after (
		.din(new_net_11251),
		.dout(new_net_11252)
	);

	bfr new_net_11253_bfr_after (
		.din(new_net_11252),
		.dout(new_net_11253)
	);

	bfr new_net_11254_bfr_after (
		.din(new_net_11253),
		.dout(new_net_11254)
	);

	bfr new_net_11255_bfr_after (
		.din(new_net_11254),
		.dout(new_net_11255)
	);

	bfr new_net_11256_bfr_after (
		.din(new_net_11255),
		.dout(new_net_11256)
	);

	spl2 _0104__v_fanout (
		.a(new_net_11256),
		.b(new_net_1459),
		.c(new_net_1460)
	);

	bfr new_net_11257_bfr_after (
		.din(_0339_),
		.dout(new_net_11257)
	);

	bfr new_net_11258_bfr_after (
		.din(new_net_11257),
		.dout(new_net_11258)
	);

	bfr new_net_11259_bfr_after (
		.din(new_net_11258),
		.dout(new_net_11259)
	);

	bfr new_net_11260_bfr_after (
		.din(new_net_11259),
		.dout(new_net_11260)
	);

	bfr new_net_11261_bfr_after (
		.din(new_net_11260),
		.dout(new_net_11261)
	);

	bfr new_net_11262_bfr_after (
		.din(new_net_11261),
		.dout(new_net_11262)
	);

	bfr new_net_11263_bfr_after (
		.din(new_net_11262),
		.dout(new_net_11263)
	);

	bfr new_net_11264_bfr_after (
		.din(new_net_11263),
		.dout(new_net_11264)
	);

	spl2 _0339__v_fanout (
		.a(new_net_11264),
		.b(new_net_1028),
		.c(new_net_1029)
	);

	bfr new_net_11265_bfr_after (
		.din(_1632_),
		.dout(new_net_11265)
	);

	bfr new_net_11266_bfr_after (
		.din(new_net_11265),
		.dout(new_net_11266)
	);

	bfr new_net_11267_bfr_after (
		.din(new_net_11266),
		.dout(new_net_11267)
	);

	bfr new_net_11268_bfr_after (
		.din(new_net_11267),
		.dout(new_net_11268)
	);

	bfr new_net_11269_bfr_after (
		.din(new_net_11268),
		.dout(new_net_11269)
	);

	bfr new_net_11270_bfr_after (
		.din(new_net_11269),
		.dout(new_net_11270)
	);

	bfr new_net_11271_bfr_after (
		.din(new_net_11270),
		.dout(new_net_11271)
	);

	bfr new_net_11272_bfr_after (
		.din(new_net_11271),
		.dout(new_net_11272)
	);

	spl2 _1632__v_fanout (
		.a(new_net_11272),
		.b(new_net_836),
		.c(new_net_837)
	);

	bfr new_net_11273_bfr_after (
		.din(_0340_),
		.dout(new_net_11273)
	);

	bfr new_net_11274_bfr_after (
		.din(new_net_11273),
		.dout(new_net_11274)
	);

	bfr new_net_11275_bfr_after (
		.din(new_net_11274),
		.dout(new_net_11275)
	);

	bfr new_net_11276_bfr_after (
		.din(new_net_11275),
		.dout(new_net_11276)
	);

	bfr new_net_11277_bfr_after (
		.din(new_net_11276),
		.dout(new_net_11277)
	);

	bfr new_net_11278_bfr_after (
		.din(new_net_11277),
		.dout(new_net_11278)
	);

	bfr new_net_11279_bfr_after (
		.din(new_net_11278),
		.dout(new_net_11279)
	);

	bfr new_net_11280_bfr_after (
		.din(new_net_11279),
		.dout(new_net_11280)
	);

	bfr new_net_11281_bfr_after (
		.din(new_net_11280),
		.dout(new_net_11281)
	);

	bfr new_net_11282_bfr_after (
		.din(new_net_11281),
		.dout(new_net_11282)
	);

	bfr new_net_11283_bfr_after (
		.din(new_net_11282),
		.dout(new_net_11283)
	);

	bfr new_net_11284_bfr_after (
		.din(new_net_11283),
		.dout(new_net_11284)
	);

	bfr new_net_11285_bfr_after (
		.din(new_net_11284),
		.dout(new_net_11285)
	);

	bfr new_net_11286_bfr_after (
		.din(new_net_11285),
		.dout(new_net_11286)
	);

	bfr new_net_11287_bfr_after (
		.din(new_net_11286),
		.dout(new_net_11287)
	);

	bfr new_net_11288_bfr_after (
		.din(new_net_11287),
		.dout(new_net_11288)
	);

	bfr new_net_11289_bfr_after (
		.din(new_net_11288),
		.dout(new_net_11289)
	);

	bfr new_net_11290_bfr_after (
		.din(new_net_11289),
		.dout(new_net_11290)
	);

	bfr new_net_11291_bfr_after (
		.din(new_net_11290),
		.dout(new_net_11291)
	);

	bfr new_net_11292_bfr_after (
		.din(new_net_11291),
		.dout(new_net_11292)
	);

	bfr new_net_11293_bfr_after (
		.din(new_net_11292),
		.dout(new_net_11293)
	);

	bfr new_net_11294_bfr_after (
		.din(new_net_11293),
		.dout(new_net_11294)
	);

	bfr new_net_11295_bfr_after (
		.din(new_net_11294),
		.dout(new_net_11295)
	);

	bfr new_net_11296_bfr_after (
		.din(new_net_11295),
		.dout(new_net_11296)
	);

	bfr new_net_11297_bfr_after (
		.din(new_net_11296),
		.dout(new_net_11297)
	);

	bfr new_net_11298_bfr_after (
		.din(new_net_11297),
		.dout(new_net_11298)
	);

	bfr new_net_11299_bfr_after (
		.din(new_net_11298),
		.dout(new_net_11299)
	);

	bfr new_net_11300_bfr_after (
		.din(new_net_11299),
		.dout(new_net_11300)
	);

	bfr new_net_11301_bfr_after (
		.din(new_net_11300),
		.dout(new_net_11301)
	);

	bfr new_net_11302_bfr_after (
		.din(new_net_11301),
		.dout(new_net_11302)
	);

	bfr new_net_11303_bfr_after (
		.din(new_net_11302),
		.dout(new_net_11303)
	);

	bfr new_net_11304_bfr_after (
		.din(new_net_11303),
		.dout(new_net_11304)
	);

	bfr new_net_11305_bfr_after (
		.din(new_net_11304),
		.dout(new_net_11305)
	);

	bfr new_net_11306_bfr_after (
		.din(new_net_11305),
		.dout(new_net_11306)
	);

	bfr new_net_11307_bfr_after (
		.din(new_net_11306),
		.dout(new_net_11307)
	);

	bfr new_net_11308_bfr_after (
		.din(new_net_11307),
		.dout(new_net_11308)
	);

	bfr new_net_11309_bfr_after (
		.din(new_net_11308),
		.dout(new_net_11309)
	);

	bfr new_net_11310_bfr_after (
		.din(new_net_11309),
		.dout(new_net_11310)
	);

	bfr new_net_11311_bfr_after (
		.din(new_net_11310),
		.dout(new_net_11311)
	);

	bfr new_net_11312_bfr_after (
		.din(new_net_11311),
		.dout(new_net_11312)
	);

	bfr new_net_11313_bfr_after (
		.din(new_net_11312),
		.dout(new_net_11313)
	);

	bfr new_net_11314_bfr_after (
		.din(new_net_11313),
		.dout(new_net_11314)
	);

	bfr new_net_11315_bfr_after (
		.din(new_net_11314),
		.dout(new_net_11315)
	);

	bfr new_net_11316_bfr_after (
		.din(new_net_11315),
		.dout(new_net_11316)
	);

	bfr new_net_11317_bfr_after (
		.din(new_net_11316),
		.dout(new_net_11317)
	);

	bfr new_net_11318_bfr_after (
		.din(new_net_11317),
		.dout(new_net_11318)
	);

	bfr new_net_11319_bfr_after (
		.din(new_net_11318),
		.dout(new_net_11319)
	);

	bfr new_net_11320_bfr_after (
		.din(new_net_11319),
		.dout(new_net_11320)
	);

	bfr new_net_11321_bfr_after (
		.din(new_net_11320),
		.dout(new_net_11321)
	);

	bfr new_net_11322_bfr_after (
		.din(new_net_11321),
		.dout(new_net_11322)
	);

	bfr new_net_11323_bfr_after (
		.din(new_net_11322),
		.dout(new_net_11323)
	);

	bfr new_net_11324_bfr_after (
		.din(new_net_11323),
		.dout(new_net_11324)
	);

	bfr new_net_11325_bfr_after (
		.din(new_net_11324),
		.dout(new_net_11325)
	);

	bfr new_net_11326_bfr_after (
		.din(new_net_11325),
		.dout(new_net_11326)
	);

	bfr new_net_11327_bfr_after (
		.din(new_net_11326),
		.dout(new_net_11327)
	);

	bfr new_net_11328_bfr_after (
		.din(new_net_11327),
		.dout(new_net_11328)
	);

	bfr new_net_11329_bfr_after (
		.din(new_net_11328),
		.dout(new_net_11329)
	);

	bfr new_net_11330_bfr_after (
		.din(new_net_11329),
		.dout(new_net_11330)
	);

	bfr new_net_11331_bfr_after (
		.din(new_net_11330),
		.dout(new_net_11331)
	);

	bfr new_net_11332_bfr_after (
		.din(new_net_11331),
		.dout(new_net_11332)
	);

	bfr new_net_11333_bfr_after (
		.din(new_net_11332),
		.dout(new_net_11333)
	);

	bfr new_net_11334_bfr_after (
		.din(new_net_11333),
		.dout(new_net_11334)
	);

	bfr new_net_11335_bfr_after (
		.din(new_net_11334),
		.dout(new_net_11335)
	);

	bfr new_net_11336_bfr_after (
		.din(new_net_11335),
		.dout(new_net_11336)
	);

	spl2 _0340__v_fanout (
		.a(new_net_11336),
		.b(new_net_1186),
		.c(new_net_1187)
	);

	spl2 _1033__v_fanout (
		.a(_1033_),
		.b(new_net_422),
		.c(new_net_423)
	);

	bfr new_net_11337_bfr_after (
		.din(_0236_),
		.dout(new_net_11337)
	);

	bfr new_net_11338_bfr_after (
		.din(new_net_11337),
		.dout(new_net_11338)
	);

	bfr new_net_11339_bfr_after (
		.din(new_net_11338),
		.dout(new_net_11339)
	);

	bfr new_net_11340_bfr_after (
		.din(new_net_11339),
		.dout(new_net_11340)
	);

	bfr new_net_11341_bfr_after (
		.din(new_net_11340),
		.dout(new_net_11341)
	);

	bfr new_net_11342_bfr_after (
		.din(new_net_11341),
		.dout(new_net_11342)
	);

	bfr new_net_11343_bfr_after (
		.din(new_net_11342),
		.dout(new_net_11343)
	);

	bfr new_net_11344_bfr_after (
		.din(new_net_11343),
		.dout(new_net_11344)
	);

	bfr new_net_11345_bfr_after (
		.din(new_net_11344),
		.dout(new_net_11345)
	);

	bfr new_net_11346_bfr_after (
		.din(new_net_11345),
		.dout(new_net_11346)
	);

	bfr new_net_11347_bfr_after (
		.din(new_net_11346),
		.dout(new_net_11347)
	);

	bfr new_net_11348_bfr_after (
		.din(new_net_11347),
		.dout(new_net_11348)
	);

	bfr new_net_11349_bfr_after (
		.din(new_net_11348),
		.dout(new_net_11349)
	);

	bfr new_net_11350_bfr_after (
		.din(new_net_11349),
		.dout(new_net_11350)
	);

	bfr new_net_11351_bfr_after (
		.din(new_net_11350),
		.dout(new_net_11351)
	);

	bfr new_net_11352_bfr_after (
		.din(new_net_11351),
		.dout(new_net_11352)
	);

	bfr new_net_11353_bfr_after (
		.din(new_net_11352),
		.dout(new_net_11353)
	);

	bfr new_net_11354_bfr_after (
		.din(new_net_11353),
		.dout(new_net_11354)
	);

	spl2 _0236__v_fanout (
		.a(new_net_11354),
		.b(new_net_466),
		.c(new_net_467)
	);

	bfr new_net_11355_bfr_after (
		.din(_1381_),
		.dout(new_net_11355)
	);

	bfr new_net_11356_bfr_after (
		.din(new_net_11355),
		.dout(new_net_11356)
	);

	bfr new_net_11357_bfr_after (
		.din(new_net_11356),
		.dout(new_net_11357)
	);

	bfr new_net_11358_bfr_after (
		.din(new_net_11357),
		.dout(new_net_11358)
	);

	bfr new_net_11359_bfr_after (
		.din(new_net_11358),
		.dout(new_net_11359)
	);

	bfr new_net_11360_bfr_after (
		.din(new_net_11359),
		.dout(new_net_11360)
	);

	bfr new_net_11361_bfr_after (
		.din(new_net_11360),
		.dout(new_net_11361)
	);

	bfr new_net_11362_bfr_after (
		.din(new_net_11361),
		.dout(new_net_11362)
	);

	spl2 _1381__v_fanout (
		.a(new_net_11362),
		.b(new_net_352),
		.c(new_net_353)
	);

	bfr new_net_11363_bfr_after (
		.din(_1067_),
		.dout(new_net_11363)
	);

	bfr new_net_11364_bfr_after (
		.din(new_net_11363),
		.dout(new_net_11364)
	);

	bfr new_net_11365_bfr_after (
		.din(new_net_11364),
		.dout(new_net_11365)
	);

	bfr new_net_11366_bfr_after (
		.din(new_net_11365),
		.dout(new_net_11366)
	);

	bfr new_net_11367_bfr_after (
		.din(new_net_11366),
		.dout(new_net_11367)
	);

	bfr new_net_11368_bfr_after (
		.din(new_net_11367),
		.dout(new_net_11368)
	);

	bfr new_net_11369_bfr_after (
		.din(new_net_11368),
		.dout(new_net_11369)
	);

	bfr new_net_11370_bfr_after (
		.din(new_net_11369),
		.dout(new_net_11370)
	);

	bfr new_net_11371_bfr_after (
		.din(new_net_11370),
		.dout(new_net_11371)
	);

	bfr new_net_11372_bfr_after (
		.din(new_net_11371),
		.dout(new_net_11372)
	);

	bfr new_net_11373_bfr_after (
		.din(new_net_11372),
		.dout(new_net_11373)
	);

	bfr new_net_11374_bfr_after (
		.din(new_net_11373),
		.dout(new_net_11374)
	);

	bfr new_net_11375_bfr_after (
		.din(new_net_11374),
		.dout(new_net_11375)
	);

	bfr new_net_11376_bfr_after (
		.din(new_net_11375),
		.dout(new_net_11376)
	);

	bfr new_net_11377_bfr_after (
		.din(new_net_11376),
		.dout(new_net_11377)
	);

	bfr new_net_11378_bfr_after (
		.din(new_net_11377),
		.dout(new_net_11378)
	);

	bfr new_net_11379_bfr_after (
		.din(new_net_11378),
		.dout(new_net_11379)
	);

	bfr new_net_11380_bfr_after (
		.din(new_net_11379),
		.dout(new_net_11380)
	);

	bfr new_net_11381_bfr_after (
		.din(new_net_11380),
		.dout(new_net_11381)
	);

	bfr new_net_11382_bfr_after (
		.din(new_net_11381),
		.dout(new_net_11382)
	);

	bfr new_net_11383_bfr_after (
		.din(new_net_11382),
		.dout(new_net_11383)
	);

	bfr new_net_11384_bfr_after (
		.din(new_net_11383),
		.dout(new_net_11384)
	);

	bfr new_net_11385_bfr_after (
		.din(new_net_11384),
		.dout(new_net_11385)
	);

	bfr new_net_11386_bfr_after (
		.din(new_net_11385),
		.dout(new_net_11386)
	);

	bfr new_net_11387_bfr_after (
		.din(new_net_11386),
		.dout(new_net_11387)
	);

	bfr new_net_11388_bfr_after (
		.din(new_net_11387),
		.dout(new_net_11388)
	);

	bfr new_net_11389_bfr_after (
		.din(new_net_11388),
		.dout(new_net_11389)
	);

	bfr new_net_11390_bfr_after (
		.din(new_net_11389),
		.dout(new_net_11390)
	);

	bfr new_net_11391_bfr_after (
		.din(new_net_11390),
		.dout(new_net_11391)
	);

	bfr new_net_11392_bfr_after (
		.din(new_net_11391),
		.dout(new_net_11392)
	);

	bfr new_net_11393_bfr_after (
		.din(new_net_11392),
		.dout(new_net_11393)
	);

	bfr new_net_11394_bfr_after (
		.din(new_net_11393),
		.dout(new_net_11394)
	);

	bfr new_net_11395_bfr_after (
		.din(new_net_11394),
		.dout(new_net_11395)
	);

	bfr new_net_11396_bfr_after (
		.din(new_net_11395),
		.dout(new_net_11396)
	);

	bfr new_net_11397_bfr_after (
		.din(new_net_11396),
		.dout(new_net_11397)
	);

	bfr new_net_11398_bfr_after (
		.din(new_net_11397),
		.dout(new_net_11398)
	);

	bfr new_net_11399_bfr_after (
		.din(new_net_11398),
		.dout(new_net_11399)
	);

	bfr new_net_11400_bfr_after (
		.din(new_net_11399),
		.dout(new_net_11400)
	);

	bfr new_net_11401_bfr_after (
		.din(new_net_11400),
		.dout(new_net_11401)
	);

	bfr new_net_11402_bfr_after (
		.din(new_net_11401),
		.dout(new_net_11402)
	);

	bfr new_net_11403_bfr_after (
		.din(new_net_11402),
		.dout(new_net_11403)
	);

	bfr new_net_11404_bfr_after (
		.din(new_net_11403),
		.dout(new_net_11404)
	);

	bfr new_net_11405_bfr_after (
		.din(new_net_11404),
		.dout(new_net_11405)
	);

	bfr new_net_11406_bfr_after (
		.din(new_net_11405),
		.dout(new_net_11406)
	);

	bfr new_net_11407_bfr_after (
		.din(new_net_11406),
		.dout(new_net_11407)
	);

	bfr new_net_11408_bfr_after (
		.din(new_net_11407),
		.dout(new_net_11408)
	);

	bfr new_net_11409_bfr_after (
		.din(new_net_11408),
		.dout(new_net_11409)
	);

	bfr new_net_11410_bfr_after (
		.din(new_net_11409),
		.dout(new_net_11410)
	);

	spl2 _1067__v_fanout (
		.a(new_net_11410),
		.b(new_net_1702),
		.c(new_net_1703)
	);

	bfr new_net_11411_bfr_after (
		.din(_1365_),
		.dout(new_net_11411)
	);

	bfr new_net_11412_bfr_after (
		.din(new_net_11411),
		.dout(new_net_11412)
	);

	bfr new_net_11413_bfr_after (
		.din(new_net_11412),
		.dout(new_net_11413)
	);

	bfr new_net_11414_bfr_after (
		.din(new_net_11413),
		.dout(new_net_11414)
	);

	bfr new_net_11415_bfr_after (
		.din(new_net_11414),
		.dout(new_net_11415)
	);

	bfr new_net_11416_bfr_after (
		.din(new_net_11415),
		.dout(new_net_11416)
	);

	bfr new_net_11417_bfr_after (
		.din(new_net_11416),
		.dout(new_net_11417)
	);

	bfr new_net_11418_bfr_after (
		.din(new_net_11417),
		.dout(new_net_11418)
	);

	bfr new_net_11419_bfr_after (
		.din(new_net_11418),
		.dout(new_net_11419)
	);

	bfr new_net_11420_bfr_after (
		.din(new_net_11419),
		.dout(new_net_11420)
	);

	bfr new_net_11421_bfr_after (
		.din(new_net_11420),
		.dout(new_net_11421)
	);

	bfr new_net_11422_bfr_after (
		.din(new_net_11421),
		.dout(new_net_11422)
	);

	bfr new_net_11423_bfr_after (
		.din(new_net_11422),
		.dout(new_net_11423)
	);

	bfr new_net_11424_bfr_after (
		.din(new_net_11423),
		.dout(new_net_11424)
	);

	bfr new_net_11425_bfr_after (
		.din(new_net_11424),
		.dout(new_net_11425)
	);

	bfr new_net_11426_bfr_after (
		.din(new_net_11425),
		.dout(new_net_11426)
	);

	bfr new_net_11427_bfr_after (
		.din(new_net_11426),
		.dout(new_net_11427)
	);

	bfr new_net_11428_bfr_after (
		.din(new_net_11427),
		.dout(new_net_11428)
	);

	bfr new_net_11429_bfr_after (
		.din(new_net_11428),
		.dout(new_net_11429)
	);

	bfr new_net_11430_bfr_after (
		.din(new_net_11429),
		.dout(new_net_11430)
	);

	bfr new_net_11431_bfr_after (
		.din(new_net_11430),
		.dout(new_net_11431)
	);

	bfr new_net_11432_bfr_after (
		.din(new_net_11431),
		.dout(new_net_11432)
	);

	bfr new_net_11433_bfr_after (
		.din(new_net_11432),
		.dout(new_net_11433)
	);

	bfr new_net_11434_bfr_after (
		.din(new_net_11433),
		.dout(new_net_11434)
	);

	bfr new_net_11435_bfr_after (
		.din(new_net_11434),
		.dout(new_net_11435)
	);

	bfr new_net_11436_bfr_after (
		.din(new_net_11435),
		.dout(new_net_11436)
	);

	bfr new_net_11437_bfr_after (
		.din(new_net_11436),
		.dout(new_net_11437)
	);

	bfr new_net_11438_bfr_after (
		.din(new_net_11437),
		.dout(new_net_11438)
	);

	bfr new_net_11439_bfr_after (
		.din(new_net_11438),
		.dout(new_net_11439)
	);

	bfr new_net_11440_bfr_after (
		.din(new_net_11439),
		.dout(new_net_11440)
	);

	bfr new_net_11441_bfr_after (
		.din(new_net_11440),
		.dout(new_net_11441)
	);

	bfr new_net_11442_bfr_after (
		.din(new_net_11441),
		.dout(new_net_11442)
	);

	bfr new_net_11443_bfr_after (
		.din(new_net_11442),
		.dout(new_net_11443)
	);

	bfr new_net_11444_bfr_after (
		.din(new_net_11443),
		.dout(new_net_11444)
	);

	bfr new_net_11445_bfr_after (
		.din(new_net_11444),
		.dout(new_net_11445)
	);

	bfr new_net_11446_bfr_after (
		.din(new_net_11445),
		.dout(new_net_11446)
	);

	bfr new_net_11447_bfr_after (
		.din(new_net_11446),
		.dout(new_net_11447)
	);

	bfr new_net_11448_bfr_after (
		.din(new_net_11447),
		.dout(new_net_11448)
	);

	bfr new_net_11449_bfr_after (
		.din(new_net_11448),
		.dout(new_net_11449)
	);

	bfr new_net_11450_bfr_after (
		.din(new_net_11449),
		.dout(new_net_11450)
	);

	bfr new_net_11451_bfr_after (
		.din(new_net_11450),
		.dout(new_net_11451)
	);

	bfr new_net_11452_bfr_after (
		.din(new_net_11451),
		.dout(new_net_11452)
	);

	bfr new_net_11453_bfr_after (
		.din(new_net_11452),
		.dout(new_net_11453)
	);

	bfr new_net_11454_bfr_after (
		.din(new_net_11453),
		.dout(new_net_11454)
	);

	bfr new_net_11455_bfr_after (
		.din(new_net_11454),
		.dout(new_net_11455)
	);

	bfr new_net_11456_bfr_after (
		.din(new_net_11455),
		.dout(new_net_11456)
	);

	bfr new_net_11457_bfr_after (
		.din(new_net_11456),
		.dout(new_net_11457)
	);

	bfr new_net_11458_bfr_after (
		.din(new_net_11457),
		.dout(new_net_11458)
	);

	bfr new_net_11459_bfr_after (
		.din(new_net_11458),
		.dout(new_net_11459)
	);

	bfr new_net_11460_bfr_after (
		.din(new_net_11459),
		.dout(new_net_11460)
	);

	bfr new_net_11461_bfr_after (
		.din(new_net_11460),
		.dout(new_net_11461)
	);

	bfr new_net_11462_bfr_after (
		.din(new_net_11461),
		.dout(new_net_11462)
	);

	bfr new_net_11463_bfr_after (
		.din(new_net_11462),
		.dout(new_net_11463)
	);

	bfr new_net_11464_bfr_after (
		.din(new_net_11463),
		.dout(new_net_11464)
	);

	bfr new_net_11465_bfr_after (
		.din(new_net_11464),
		.dout(new_net_11465)
	);

	bfr new_net_11466_bfr_after (
		.din(new_net_11465),
		.dout(new_net_11466)
	);

	bfr new_net_11467_bfr_after (
		.din(new_net_11466),
		.dout(new_net_11467)
	);

	bfr new_net_11468_bfr_after (
		.din(new_net_11467),
		.dout(new_net_11468)
	);

	bfr new_net_11469_bfr_after (
		.din(new_net_11468),
		.dout(new_net_11469)
	);

	bfr new_net_11470_bfr_after (
		.din(new_net_11469),
		.dout(new_net_11470)
	);

	bfr new_net_11471_bfr_after (
		.din(new_net_11470),
		.dout(new_net_11471)
	);

	bfr new_net_11472_bfr_after (
		.din(new_net_11471),
		.dout(new_net_11472)
	);

	bfr new_net_11473_bfr_after (
		.din(new_net_11472),
		.dout(new_net_11473)
	);

	bfr new_net_11474_bfr_after (
		.din(new_net_11473),
		.dout(new_net_11474)
	);

	bfr new_net_11475_bfr_after (
		.din(new_net_11474),
		.dout(new_net_11475)
	);

	bfr new_net_11476_bfr_after (
		.din(new_net_11475),
		.dout(new_net_11476)
	);

	bfr new_net_11477_bfr_after (
		.din(new_net_11476),
		.dout(new_net_11477)
	);

	bfr new_net_11478_bfr_after (
		.din(new_net_11477),
		.dout(new_net_11478)
	);

	bfr new_net_11479_bfr_after (
		.din(new_net_11478),
		.dout(new_net_11479)
	);

	bfr new_net_11480_bfr_after (
		.din(new_net_11479),
		.dout(new_net_11480)
	);

	bfr new_net_11481_bfr_after (
		.din(new_net_11480),
		.dout(new_net_11481)
	);

	bfr new_net_11482_bfr_after (
		.din(new_net_11481),
		.dout(new_net_11482)
	);

	spl2 _1365__v_fanout (
		.a(new_net_11482),
		.b(new_net_1836),
		.c(new_net_1837)
	);

	bfr new_net_11483_bfr_after (
		.din(_1367_),
		.dout(new_net_11483)
	);

	bfr new_net_11484_bfr_after (
		.din(new_net_11483),
		.dout(new_net_11484)
	);

	bfr new_net_11485_bfr_after (
		.din(new_net_11484),
		.dout(new_net_11485)
	);

	bfr new_net_11486_bfr_after (
		.din(new_net_11485),
		.dout(new_net_11486)
	);

	bfr new_net_11487_bfr_after (
		.din(new_net_11486),
		.dout(new_net_11487)
	);

	bfr new_net_11488_bfr_after (
		.din(new_net_11487),
		.dout(new_net_11488)
	);

	bfr new_net_11489_bfr_after (
		.din(new_net_11488),
		.dout(new_net_11489)
	);

	bfr new_net_11490_bfr_after (
		.din(new_net_11489),
		.dout(new_net_11490)
	);

	bfr new_net_11491_bfr_after (
		.din(new_net_11490),
		.dout(new_net_11491)
	);

	bfr new_net_11492_bfr_after (
		.din(new_net_11491),
		.dout(new_net_11492)
	);

	bfr new_net_11493_bfr_after (
		.din(new_net_11492),
		.dout(new_net_11493)
	);

	bfr new_net_11494_bfr_after (
		.din(new_net_11493),
		.dout(new_net_11494)
	);

	bfr new_net_11495_bfr_after (
		.din(new_net_11494),
		.dout(new_net_11495)
	);

	bfr new_net_11496_bfr_after (
		.din(new_net_11495),
		.dout(new_net_11496)
	);

	bfr new_net_11497_bfr_after (
		.din(new_net_11496),
		.dout(new_net_11497)
	);

	bfr new_net_11498_bfr_after (
		.din(new_net_11497),
		.dout(new_net_11498)
	);

	bfr new_net_11499_bfr_after (
		.din(new_net_11498),
		.dout(new_net_11499)
	);

	bfr new_net_11500_bfr_after (
		.din(new_net_11499),
		.dout(new_net_11500)
	);

	bfr new_net_11501_bfr_after (
		.din(new_net_11500),
		.dout(new_net_11501)
	);

	bfr new_net_11502_bfr_after (
		.din(new_net_11501),
		.dout(new_net_11502)
	);

	bfr new_net_11503_bfr_after (
		.din(new_net_11502),
		.dout(new_net_11503)
	);

	bfr new_net_11504_bfr_after (
		.din(new_net_11503),
		.dout(new_net_11504)
	);

	bfr new_net_11505_bfr_after (
		.din(new_net_11504),
		.dout(new_net_11505)
	);

	bfr new_net_11506_bfr_after (
		.din(new_net_11505),
		.dout(new_net_11506)
	);

	bfr new_net_11507_bfr_after (
		.din(new_net_11506),
		.dout(new_net_11507)
	);

	bfr new_net_11508_bfr_after (
		.din(new_net_11507),
		.dout(new_net_11508)
	);

	bfr new_net_11509_bfr_after (
		.din(new_net_11508),
		.dout(new_net_11509)
	);

	bfr new_net_11510_bfr_after (
		.din(new_net_11509),
		.dout(new_net_11510)
	);

	bfr new_net_11511_bfr_after (
		.din(new_net_11510),
		.dout(new_net_11511)
	);

	bfr new_net_11512_bfr_after (
		.din(new_net_11511),
		.dout(new_net_11512)
	);

	bfr new_net_11513_bfr_after (
		.din(new_net_11512),
		.dout(new_net_11513)
	);

	bfr new_net_11514_bfr_after (
		.din(new_net_11513),
		.dout(new_net_11514)
	);

	bfr new_net_11515_bfr_after (
		.din(new_net_11514),
		.dout(new_net_11515)
	);

	bfr new_net_11516_bfr_after (
		.din(new_net_11515),
		.dout(new_net_11516)
	);

	bfr new_net_11517_bfr_after (
		.din(new_net_11516),
		.dout(new_net_11517)
	);

	bfr new_net_11518_bfr_after (
		.din(new_net_11517),
		.dout(new_net_11518)
	);

	bfr new_net_11519_bfr_after (
		.din(new_net_11518),
		.dout(new_net_11519)
	);

	bfr new_net_11520_bfr_after (
		.din(new_net_11519),
		.dout(new_net_11520)
	);

	bfr new_net_11521_bfr_after (
		.din(new_net_11520),
		.dout(new_net_11521)
	);

	bfr new_net_11522_bfr_after (
		.din(new_net_11521),
		.dout(new_net_11522)
	);

	bfr new_net_11523_bfr_after (
		.din(new_net_11522),
		.dout(new_net_11523)
	);

	bfr new_net_11524_bfr_after (
		.din(new_net_11523),
		.dout(new_net_11524)
	);

	bfr new_net_11525_bfr_after (
		.din(new_net_11524),
		.dout(new_net_11525)
	);

	bfr new_net_11526_bfr_after (
		.din(new_net_11525),
		.dout(new_net_11526)
	);

	bfr new_net_11527_bfr_after (
		.din(new_net_11526),
		.dout(new_net_11527)
	);

	bfr new_net_11528_bfr_after (
		.din(new_net_11527),
		.dout(new_net_11528)
	);

	bfr new_net_11529_bfr_after (
		.din(new_net_11528),
		.dout(new_net_11529)
	);

	bfr new_net_11530_bfr_after (
		.din(new_net_11529),
		.dout(new_net_11530)
	);

	bfr new_net_11531_bfr_after (
		.din(new_net_11530),
		.dout(new_net_11531)
	);

	bfr new_net_11532_bfr_after (
		.din(new_net_11531),
		.dout(new_net_11532)
	);

	bfr new_net_11533_bfr_after (
		.din(new_net_11532),
		.dout(new_net_11533)
	);

	bfr new_net_11534_bfr_after (
		.din(new_net_11533),
		.dout(new_net_11534)
	);

	bfr new_net_11535_bfr_after (
		.din(new_net_11534),
		.dout(new_net_11535)
	);

	bfr new_net_11536_bfr_after (
		.din(new_net_11535),
		.dout(new_net_11536)
	);

	bfr new_net_11537_bfr_after (
		.din(new_net_11536),
		.dout(new_net_11537)
	);

	bfr new_net_11538_bfr_after (
		.din(new_net_11537),
		.dout(new_net_11538)
	);

	bfr new_net_11539_bfr_after (
		.din(new_net_11538),
		.dout(new_net_11539)
	);

	bfr new_net_11540_bfr_after (
		.din(new_net_11539),
		.dout(new_net_11540)
	);

	bfr new_net_11541_bfr_after (
		.din(new_net_11540),
		.dout(new_net_11541)
	);

	bfr new_net_11542_bfr_after (
		.din(new_net_11541),
		.dout(new_net_11542)
	);

	bfr new_net_11543_bfr_after (
		.din(new_net_11542),
		.dout(new_net_11543)
	);

	bfr new_net_11544_bfr_after (
		.din(new_net_11543),
		.dout(new_net_11544)
	);

	bfr new_net_11545_bfr_after (
		.din(new_net_11544),
		.dout(new_net_11545)
	);

	bfr new_net_11546_bfr_after (
		.din(new_net_11545),
		.dout(new_net_11546)
	);

	spl2 _1367__v_fanout (
		.a(new_net_11546),
		.b(new_net_1912),
		.c(new_net_1913)
	);

	bfr new_net_11547_bfr_before (
		.din(new_net_11547),
		.dout(new_net_2375)
	);

	spl2 _1709__v_fanout (
		.a(_1709_),
		.b(new_net_2374),
		.c(new_net_11547)
	);

	bfr new_net_11548_bfr_after (
		.din(_1024_),
		.dout(new_net_11548)
	);

	bfr new_net_11549_bfr_after (
		.din(new_net_11548),
		.dout(new_net_11549)
	);

	bfr new_net_11550_bfr_after (
		.din(new_net_11549),
		.dout(new_net_11550)
	);

	bfr new_net_11551_bfr_after (
		.din(new_net_11550),
		.dout(new_net_11551)
	);

	bfr new_net_11552_bfr_after (
		.din(new_net_11551),
		.dout(new_net_11552)
	);

	bfr new_net_11553_bfr_after (
		.din(new_net_11552),
		.dout(new_net_11553)
	);

	bfr new_net_11554_bfr_after (
		.din(new_net_11553),
		.dout(new_net_11554)
	);

	bfr new_net_11555_bfr_after (
		.din(new_net_11554),
		.dout(new_net_11555)
	);

	bfr new_net_11556_bfr_after (
		.din(new_net_11555),
		.dout(new_net_11556)
	);

	bfr new_net_11557_bfr_after (
		.din(new_net_11556),
		.dout(new_net_11557)
	);

	bfr new_net_11558_bfr_after (
		.din(new_net_11557),
		.dout(new_net_11558)
	);

	bfr new_net_11559_bfr_after (
		.din(new_net_11558),
		.dout(new_net_11559)
	);

	bfr new_net_11560_bfr_after (
		.din(new_net_11559),
		.dout(new_net_11560)
	);

	bfr new_net_11561_bfr_after (
		.din(new_net_11560),
		.dout(new_net_11561)
	);

	bfr new_net_11562_bfr_after (
		.din(new_net_11561),
		.dout(new_net_11562)
	);

	bfr new_net_11563_bfr_after (
		.din(new_net_11562),
		.dout(new_net_11563)
	);

	bfr new_net_11564_bfr_after (
		.din(new_net_11563),
		.dout(new_net_11564)
	);

	bfr new_net_11565_bfr_after (
		.din(new_net_11564),
		.dout(new_net_11565)
	);

	bfr new_net_11566_bfr_after (
		.din(new_net_11565),
		.dout(new_net_11566)
	);

	bfr new_net_11567_bfr_after (
		.din(new_net_11566),
		.dout(new_net_11567)
	);

	bfr new_net_11568_bfr_after (
		.din(new_net_11567),
		.dout(new_net_11568)
	);

	bfr new_net_11569_bfr_after (
		.din(new_net_11568),
		.dout(new_net_11569)
	);

	bfr new_net_11570_bfr_after (
		.din(new_net_11569),
		.dout(new_net_11570)
	);

	bfr new_net_11571_bfr_after (
		.din(new_net_11570),
		.dout(new_net_11571)
	);

	bfr new_net_11572_bfr_after (
		.din(new_net_11571),
		.dout(new_net_11572)
	);

	bfr new_net_11573_bfr_after (
		.din(new_net_11572),
		.dout(new_net_11573)
	);

	bfr new_net_11574_bfr_after (
		.din(new_net_11573),
		.dout(new_net_11574)
	);

	bfr new_net_11575_bfr_after (
		.din(new_net_11574),
		.dout(new_net_11575)
	);

	bfr new_net_11576_bfr_after (
		.din(new_net_11575),
		.dout(new_net_11576)
	);

	bfr new_net_11577_bfr_after (
		.din(new_net_11576),
		.dout(new_net_11577)
	);

	bfr new_net_11578_bfr_after (
		.din(new_net_11577),
		.dout(new_net_11578)
	);

	bfr new_net_11579_bfr_after (
		.din(new_net_11578),
		.dout(new_net_11579)
	);

	spl2 _1024__v_fanout (
		.a(new_net_11579),
		.b(new_net_96),
		.c(new_net_97)
	);

	bfr new_net_11580_bfr_after (
		.din(_0453_),
		.dout(new_net_11580)
	);

	bfr new_net_11581_bfr_after (
		.din(new_net_11580),
		.dout(new_net_11581)
	);

	bfr new_net_11582_bfr_after (
		.din(new_net_11581),
		.dout(new_net_11582)
	);

	bfr new_net_11583_bfr_after (
		.din(new_net_11582),
		.dout(new_net_11583)
	);

	bfr new_net_11584_bfr_after (
		.din(new_net_11583),
		.dout(new_net_11584)
	);

	bfr new_net_11585_bfr_after (
		.din(new_net_11584),
		.dout(new_net_11585)
	);

	bfr new_net_11586_bfr_after (
		.din(new_net_11585),
		.dout(new_net_11586)
	);

	bfr new_net_11587_bfr_after (
		.din(new_net_11586),
		.dout(new_net_11587)
	);

	bfr new_net_11588_bfr_after (
		.din(new_net_11587),
		.dout(new_net_11588)
	);

	bfr new_net_11589_bfr_after (
		.din(new_net_11588),
		.dout(new_net_11589)
	);

	bfr new_net_11590_bfr_after (
		.din(new_net_11589),
		.dout(new_net_11590)
	);

	bfr new_net_11591_bfr_after (
		.din(new_net_11590),
		.dout(new_net_11591)
	);

	bfr new_net_11592_bfr_after (
		.din(new_net_11591),
		.dout(new_net_11592)
	);

	bfr new_net_11593_bfr_after (
		.din(new_net_11592),
		.dout(new_net_11593)
	);

	bfr new_net_11594_bfr_after (
		.din(new_net_11593),
		.dout(new_net_11594)
	);

	bfr new_net_11595_bfr_after (
		.din(new_net_11594),
		.dout(new_net_11595)
	);

	bfr new_net_11596_bfr_after (
		.din(new_net_11595),
		.dout(new_net_11596)
	);

	bfr new_net_11597_bfr_after (
		.din(new_net_11596),
		.dout(new_net_11597)
	);

	bfr new_net_11598_bfr_after (
		.din(new_net_11597),
		.dout(new_net_11598)
	);

	bfr new_net_11599_bfr_after (
		.din(new_net_11598),
		.dout(new_net_11599)
	);

	bfr new_net_11600_bfr_after (
		.din(new_net_11599),
		.dout(new_net_11600)
	);

	bfr new_net_11601_bfr_after (
		.din(new_net_11600),
		.dout(new_net_11601)
	);

	bfr new_net_11602_bfr_after (
		.din(new_net_11601),
		.dout(new_net_11602)
	);

	bfr new_net_11603_bfr_after (
		.din(new_net_11602),
		.dout(new_net_11603)
	);

	bfr new_net_11604_bfr_after (
		.din(new_net_11603),
		.dout(new_net_11604)
	);

	bfr new_net_11605_bfr_after (
		.din(new_net_11604),
		.dout(new_net_11605)
	);

	bfr new_net_11606_bfr_after (
		.din(new_net_11605),
		.dout(new_net_11606)
	);

	bfr new_net_11607_bfr_after (
		.din(new_net_11606),
		.dout(new_net_11607)
	);

	bfr new_net_11608_bfr_after (
		.din(new_net_11607),
		.dout(new_net_11608)
	);

	bfr new_net_11609_bfr_after (
		.din(new_net_11608),
		.dout(new_net_11609)
	);

	spl2 _0453__v_fanout (
		.a(new_net_11609),
		.b(new_net_350),
		.c(new_net_351)
	);

	spl2 _1220__v_fanout (
		.a(_1220_),
		.b(new_net_2987),
		.c(new_net_2988)
	);

	spl3L _1587__v_fanout (
		.a(_1587_),
		.b(new_net_2304),
		.c(new_net_2305),
		.d(new_net_2306)
	);

	bfr new_net_11610_bfr_after (
		.din(_0337_),
		.dout(new_net_11610)
	);

	bfr new_net_11611_bfr_after (
		.din(new_net_11610),
		.dout(new_net_11611)
	);

	bfr new_net_11612_bfr_after (
		.din(new_net_11611),
		.dout(new_net_11612)
	);

	bfr new_net_11613_bfr_after (
		.din(new_net_11612),
		.dout(new_net_11613)
	);

	bfr new_net_11614_bfr_after (
		.din(new_net_11613),
		.dout(new_net_11614)
	);

	bfr new_net_11615_bfr_after (
		.din(new_net_11614),
		.dout(new_net_11615)
	);

	bfr new_net_11616_bfr_after (
		.din(new_net_11615),
		.dout(new_net_11616)
	);

	bfr new_net_11617_bfr_after (
		.din(new_net_11616),
		.dout(new_net_11617)
	);

	bfr new_net_11618_bfr_after (
		.din(new_net_11617),
		.dout(new_net_11618)
	);

	bfr new_net_11619_bfr_after (
		.din(new_net_11618),
		.dout(new_net_11619)
	);

	bfr new_net_11620_bfr_after (
		.din(new_net_11619),
		.dout(new_net_11620)
	);

	bfr new_net_11621_bfr_after (
		.din(new_net_11620),
		.dout(new_net_11621)
	);

	bfr new_net_11622_bfr_after (
		.din(new_net_11621),
		.dout(new_net_11622)
	);

	bfr new_net_11623_bfr_after (
		.din(new_net_11622),
		.dout(new_net_11623)
	);

	bfr new_net_11624_bfr_after (
		.din(new_net_11623),
		.dout(new_net_11624)
	);

	bfr new_net_11625_bfr_after (
		.din(new_net_11624),
		.dout(new_net_11625)
	);

	bfr new_net_11626_bfr_after (
		.din(new_net_11625),
		.dout(new_net_11626)
	);

	bfr new_net_11627_bfr_after (
		.din(new_net_11626),
		.dout(new_net_11627)
	);

	bfr new_net_11628_bfr_after (
		.din(new_net_11627),
		.dout(new_net_11628)
	);

	bfr new_net_11629_bfr_after (
		.din(new_net_11628),
		.dout(new_net_11629)
	);

	bfr new_net_11630_bfr_after (
		.din(new_net_11629),
		.dout(new_net_11630)
	);

	bfr new_net_11631_bfr_after (
		.din(new_net_11630),
		.dout(new_net_11631)
	);

	bfr new_net_11632_bfr_after (
		.din(new_net_11631),
		.dout(new_net_11632)
	);

	bfr new_net_11633_bfr_after (
		.din(new_net_11632),
		.dout(new_net_11633)
	);

	bfr new_net_11634_bfr_after (
		.din(new_net_11633),
		.dout(new_net_11634)
	);

	bfr new_net_11635_bfr_after (
		.din(new_net_11634),
		.dout(new_net_11635)
	);

	bfr new_net_11636_bfr_after (
		.din(new_net_11635),
		.dout(new_net_11636)
	);

	bfr new_net_11637_bfr_after (
		.din(new_net_11636),
		.dout(new_net_11637)
	);

	bfr new_net_11638_bfr_after (
		.din(new_net_11637),
		.dout(new_net_11638)
	);

	bfr new_net_11639_bfr_after (
		.din(new_net_11638),
		.dout(new_net_11639)
	);

	bfr new_net_11640_bfr_after (
		.din(new_net_11639),
		.dout(new_net_11640)
	);

	bfr new_net_11641_bfr_after (
		.din(new_net_11640),
		.dout(new_net_11641)
	);

	bfr new_net_11642_bfr_after (
		.din(new_net_11641),
		.dout(new_net_11642)
	);

	bfr new_net_11643_bfr_after (
		.din(new_net_11642),
		.dout(new_net_11643)
	);

	bfr new_net_11644_bfr_after (
		.din(new_net_11643),
		.dout(new_net_11644)
	);

	bfr new_net_11645_bfr_after (
		.din(new_net_11644),
		.dout(new_net_11645)
	);

	bfr new_net_11646_bfr_after (
		.din(new_net_11645),
		.dout(new_net_11646)
	);

	bfr new_net_11647_bfr_after (
		.din(new_net_11646),
		.dout(new_net_11647)
	);

	bfr new_net_11648_bfr_after (
		.din(new_net_11647),
		.dout(new_net_11648)
	);

	bfr new_net_11649_bfr_after (
		.din(new_net_11648),
		.dout(new_net_11649)
	);

	bfr new_net_11650_bfr_after (
		.din(new_net_11649),
		.dout(new_net_11650)
	);

	bfr new_net_11651_bfr_after (
		.din(new_net_11650),
		.dout(new_net_11651)
	);

	bfr new_net_11652_bfr_after (
		.din(new_net_11651),
		.dout(new_net_11652)
	);

	bfr new_net_11653_bfr_after (
		.din(new_net_11652),
		.dout(new_net_11653)
	);

	bfr new_net_11654_bfr_after (
		.din(new_net_11653),
		.dout(new_net_11654)
	);

	bfr new_net_11655_bfr_after (
		.din(new_net_11654),
		.dout(new_net_11655)
	);

	bfr new_net_11656_bfr_after (
		.din(new_net_11655),
		.dout(new_net_11656)
	);

	bfr new_net_11657_bfr_after (
		.din(new_net_11656),
		.dout(new_net_11657)
	);

	bfr new_net_11658_bfr_after (
		.din(new_net_11657),
		.dout(new_net_11658)
	);

	bfr new_net_11659_bfr_after (
		.din(new_net_11658),
		.dout(new_net_11659)
	);

	bfr new_net_11660_bfr_after (
		.din(new_net_11659),
		.dout(new_net_11660)
	);

	bfr new_net_11661_bfr_after (
		.din(new_net_11660),
		.dout(new_net_11661)
	);

	bfr new_net_11662_bfr_after (
		.din(new_net_11661),
		.dout(new_net_11662)
	);

	bfr new_net_11663_bfr_after (
		.din(new_net_11662),
		.dout(new_net_11663)
	);

	bfr new_net_11664_bfr_after (
		.din(new_net_11663),
		.dout(new_net_11664)
	);

	bfr new_net_11665_bfr_after (
		.din(new_net_11664),
		.dout(new_net_11665)
	);

	bfr new_net_11666_bfr_after (
		.din(new_net_11665),
		.dout(new_net_11666)
	);

	bfr new_net_11667_bfr_after (
		.din(new_net_11666),
		.dout(new_net_11667)
	);

	bfr new_net_11668_bfr_after (
		.din(new_net_11667),
		.dout(new_net_11668)
	);

	bfr new_net_11669_bfr_after (
		.din(new_net_11668),
		.dout(new_net_11669)
	);

	bfr new_net_11670_bfr_after (
		.din(new_net_11669),
		.dout(new_net_11670)
	);

	bfr new_net_11671_bfr_after (
		.din(new_net_11670),
		.dout(new_net_11671)
	);

	bfr new_net_11672_bfr_after (
		.din(new_net_11671),
		.dout(new_net_11672)
	);

	bfr new_net_11673_bfr_after (
		.din(new_net_11672),
		.dout(new_net_11673)
	);

	bfr new_net_11674_bfr_after (
		.din(new_net_11673),
		.dout(new_net_11674)
	);

	bfr new_net_11675_bfr_after (
		.din(new_net_11674),
		.dout(new_net_11675)
	);

	bfr new_net_11676_bfr_after (
		.din(new_net_11675),
		.dout(new_net_11676)
	);

	bfr new_net_11677_bfr_after (
		.din(new_net_11676),
		.dout(new_net_11677)
	);

	bfr new_net_11678_bfr_after (
		.din(new_net_11677),
		.dout(new_net_11678)
	);

	bfr new_net_11679_bfr_after (
		.din(new_net_11678),
		.dout(new_net_11679)
	);

	bfr new_net_11680_bfr_after (
		.din(new_net_11679),
		.dout(new_net_11680)
	);

	bfr new_net_11681_bfr_after (
		.din(new_net_11680),
		.dout(new_net_11681)
	);

	spl2 _0337__v_fanout (
		.a(new_net_11681),
		.b(new_net_1078),
		.c(new_net_1079)
	);

	bfr new_net_11682_bfr_after (
		.din(_1470_),
		.dout(new_net_11682)
	);

	bfr new_net_11683_bfr_after (
		.din(new_net_11682),
		.dout(new_net_11683)
	);

	bfr new_net_11684_bfr_after (
		.din(new_net_11683),
		.dout(new_net_11684)
	);

	bfr new_net_11685_bfr_after (
		.din(new_net_11684),
		.dout(new_net_11685)
	);

	bfr new_net_11686_bfr_after (
		.din(new_net_11685),
		.dout(new_net_11686)
	);

	bfr new_net_11687_bfr_after (
		.din(new_net_11686),
		.dout(new_net_11687)
	);

	bfr new_net_11688_bfr_after (
		.din(new_net_11687),
		.dout(new_net_11688)
	);

	bfr new_net_11689_bfr_after (
		.din(new_net_11688),
		.dout(new_net_11689)
	);

	bfr new_net_11690_bfr_after (
		.din(new_net_11689),
		.dout(new_net_11690)
	);

	bfr new_net_11691_bfr_after (
		.din(new_net_11690),
		.dout(new_net_11691)
	);

	bfr new_net_11692_bfr_after (
		.din(new_net_11691),
		.dout(new_net_11692)
	);

	bfr new_net_11693_bfr_after (
		.din(new_net_11692),
		.dout(new_net_11693)
	);

	bfr new_net_11694_bfr_after (
		.din(new_net_11693),
		.dout(new_net_11694)
	);

	bfr new_net_11695_bfr_after (
		.din(new_net_11694),
		.dout(new_net_11695)
	);

	bfr new_net_11696_bfr_after (
		.din(new_net_11695),
		.dout(new_net_11696)
	);

	bfr new_net_11697_bfr_after (
		.din(new_net_11696),
		.dout(new_net_11697)
	);

	bfr new_net_11698_bfr_after (
		.din(new_net_11697),
		.dout(new_net_11698)
	);

	bfr new_net_11699_bfr_after (
		.din(new_net_11698),
		.dout(new_net_11699)
	);

	bfr new_net_11700_bfr_after (
		.din(new_net_11699),
		.dout(new_net_11700)
	);

	bfr new_net_11701_bfr_after (
		.din(new_net_11700),
		.dout(new_net_11701)
	);

	bfr new_net_11702_bfr_after (
		.din(new_net_11701),
		.dout(new_net_11702)
	);

	bfr new_net_11703_bfr_after (
		.din(new_net_11702),
		.dout(new_net_11703)
	);

	bfr new_net_11704_bfr_after (
		.din(new_net_11703),
		.dout(new_net_11704)
	);

	bfr new_net_11705_bfr_after (
		.din(new_net_11704),
		.dout(new_net_11705)
	);

	bfr new_net_11706_bfr_after (
		.din(new_net_11705),
		.dout(new_net_11706)
	);

	bfr new_net_11707_bfr_after (
		.din(new_net_11706),
		.dout(new_net_11707)
	);

	bfr new_net_11708_bfr_after (
		.din(new_net_11707),
		.dout(new_net_11708)
	);

	bfr new_net_11709_bfr_after (
		.din(new_net_11708),
		.dout(new_net_11709)
	);

	bfr new_net_11710_bfr_after (
		.din(new_net_11709),
		.dout(new_net_11710)
	);

	bfr new_net_11711_bfr_after (
		.din(new_net_11710),
		.dout(new_net_11711)
	);

	bfr new_net_11712_bfr_after (
		.din(new_net_11711),
		.dout(new_net_11712)
	);

	bfr new_net_11713_bfr_after (
		.din(new_net_11712),
		.dout(new_net_11713)
	);

	spl2 _1470__v_fanout (
		.a(new_net_11713),
		.b(new_net_1046),
		.c(new_net_1047)
	);

	bfr new_net_11714_bfr_after (
		.din(_1072_),
		.dout(new_net_11714)
	);

	bfr new_net_11715_bfr_after (
		.din(new_net_11714),
		.dout(new_net_11715)
	);

	bfr new_net_11716_bfr_after (
		.din(new_net_11715),
		.dout(new_net_11716)
	);

	bfr new_net_11717_bfr_after (
		.din(new_net_11716),
		.dout(new_net_11717)
	);

	bfr new_net_11718_bfr_after (
		.din(new_net_11717),
		.dout(new_net_11718)
	);

	bfr new_net_11719_bfr_after (
		.din(new_net_11718),
		.dout(new_net_11719)
	);

	bfr new_net_11720_bfr_after (
		.din(new_net_11719),
		.dout(new_net_11720)
	);

	bfr new_net_11721_bfr_after (
		.din(new_net_11720),
		.dout(new_net_11721)
	);

	bfr new_net_11722_bfr_after (
		.din(new_net_11721),
		.dout(new_net_11722)
	);

	bfr new_net_11723_bfr_after (
		.din(new_net_11722),
		.dout(new_net_11723)
	);

	bfr new_net_11724_bfr_after (
		.din(new_net_11723),
		.dout(new_net_11724)
	);

	bfr new_net_11725_bfr_after (
		.din(new_net_11724),
		.dout(new_net_11725)
	);

	bfr new_net_11726_bfr_after (
		.din(new_net_11725),
		.dout(new_net_11726)
	);

	bfr new_net_11727_bfr_after (
		.din(new_net_11726),
		.dout(new_net_11727)
	);

	bfr new_net_11728_bfr_after (
		.din(new_net_11727),
		.dout(new_net_11728)
	);

	bfr new_net_11729_bfr_after (
		.din(new_net_11728),
		.dout(new_net_11729)
	);

	bfr new_net_11730_bfr_after (
		.din(new_net_11729),
		.dout(new_net_11730)
	);

	bfr new_net_11731_bfr_after (
		.din(new_net_11730),
		.dout(new_net_11731)
	);

	bfr new_net_11732_bfr_after (
		.din(new_net_11731),
		.dout(new_net_11732)
	);

	bfr new_net_11733_bfr_after (
		.din(new_net_11732),
		.dout(new_net_11733)
	);

	bfr new_net_11734_bfr_after (
		.din(new_net_11733),
		.dout(new_net_11734)
	);

	bfr new_net_11735_bfr_after (
		.din(new_net_11734),
		.dout(new_net_11735)
	);

	bfr new_net_11736_bfr_after (
		.din(new_net_11735),
		.dout(new_net_11736)
	);

	bfr new_net_11737_bfr_after (
		.din(new_net_11736),
		.dout(new_net_11737)
	);

	bfr new_net_11738_bfr_after (
		.din(new_net_11737),
		.dout(new_net_11738)
	);

	bfr new_net_11739_bfr_after (
		.din(new_net_11738),
		.dout(new_net_11739)
	);

	bfr new_net_11740_bfr_after (
		.din(new_net_11739),
		.dout(new_net_11740)
	);

	bfr new_net_11741_bfr_after (
		.din(new_net_11740),
		.dout(new_net_11741)
	);

	bfr new_net_11742_bfr_after (
		.din(new_net_11741),
		.dout(new_net_11742)
	);

	bfr new_net_11743_bfr_after (
		.din(new_net_11742),
		.dout(new_net_11743)
	);

	bfr new_net_11744_bfr_after (
		.din(new_net_11743),
		.dout(new_net_11744)
	);

	bfr new_net_11745_bfr_after (
		.din(new_net_11744),
		.dout(new_net_11745)
	);

	bfr new_net_11746_bfr_after (
		.din(new_net_11745),
		.dout(new_net_11746)
	);

	bfr new_net_11747_bfr_after (
		.din(new_net_11746),
		.dout(new_net_11747)
	);

	bfr new_net_11748_bfr_after (
		.din(new_net_11747),
		.dout(new_net_11748)
	);

	bfr new_net_11749_bfr_after (
		.din(new_net_11748),
		.dout(new_net_11749)
	);

	bfr new_net_11750_bfr_after (
		.din(new_net_11749),
		.dout(new_net_11750)
	);

	bfr new_net_11751_bfr_after (
		.din(new_net_11750),
		.dout(new_net_11751)
	);

	bfr new_net_11752_bfr_after (
		.din(new_net_11751),
		.dout(new_net_11752)
	);

	bfr new_net_11753_bfr_after (
		.din(new_net_11752),
		.dout(new_net_11753)
	);

	bfr new_net_11754_bfr_after (
		.din(new_net_11753),
		.dout(new_net_11754)
	);

	bfr new_net_11755_bfr_after (
		.din(new_net_11754),
		.dout(new_net_11755)
	);

	bfr new_net_11756_bfr_after (
		.din(new_net_11755),
		.dout(new_net_11756)
	);

	bfr new_net_11757_bfr_after (
		.din(new_net_11756),
		.dout(new_net_11757)
	);

	bfr new_net_11758_bfr_after (
		.din(new_net_11757),
		.dout(new_net_11758)
	);

	bfr new_net_11759_bfr_after (
		.din(new_net_11758),
		.dout(new_net_11759)
	);

	bfr new_net_11760_bfr_after (
		.din(new_net_11759),
		.dout(new_net_11760)
	);

	bfr new_net_11761_bfr_after (
		.din(new_net_11760),
		.dout(new_net_11761)
	);

	spl2 _1072__v_fanout (
		.a(new_net_11761),
		.b(new_net_1874),
		.c(new_net_1875)
	);

	bfr new_net_11762_bfr_after (
		.din(_0688_),
		.dout(new_net_11762)
	);

	bfr new_net_11763_bfr_after (
		.din(new_net_11762),
		.dout(new_net_11763)
	);

	bfr new_net_11764_bfr_after (
		.din(new_net_11763),
		.dout(new_net_11764)
	);

	bfr new_net_11765_bfr_after (
		.din(new_net_11764),
		.dout(new_net_11765)
	);

	bfr new_net_11766_bfr_after (
		.din(new_net_11765),
		.dout(new_net_11766)
	);

	bfr new_net_11767_bfr_after (
		.din(new_net_11766),
		.dout(new_net_11767)
	);

	bfr new_net_11768_bfr_after (
		.din(new_net_11767),
		.dout(new_net_11768)
	);

	bfr new_net_11769_bfr_after (
		.din(new_net_11768),
		.dout(new_net_11769)
	);

	bfr new_net_11770_bfr_after (
		.din(new_net_11769),
		.dout(new_net_11770)
	);

	bfr new_net_11771_bfr_after (
		.din(new_net_11770),
		.dout(new_net_11771)
	);

	bfr new_net_11772_bfr_after (
		.din(new_net_11771),
		.dout(new_net_11772)
	);

	bfr new_net_11773_bfr_after (
		.din(new_net_11772),
		.dout(new_net_11773)
	);

	bfr new_net_11774_bfr_after (
		.din(new_net_11773),
		.dout(new_net_11774)
	);

	bfr new_net_11775_bfr_after (
		.din(new_net_11774),
		.dout(new_net_11775)
	);

	bfr new_net_11776_bfr_after (
		.din(new_net_11775),
		.dout(new_net_11776)
	);

	bfr new_net_11777_bfr_after (
		.din(new_net_11776),
		.dout(new_net_11777)
	);

	bfr new_net_11778_bfr_after (
		.din(new_net_11777),
		.dout(new_net_11778)
	);

	bfr new_net_11779_bfr_after (
		.din(new_net_11778),
		.dout(new_net_11779)
	);

	bfr new_net_11780_bfr_after (
		.din(new_net_11779),
		.dout(new_net_11780)
	);

	bfr new_net_11781_bfr_after (
		.din(new_net_11780),
		.dout(new_net_11781)
	);

	bfr new_net_11782_bfr_after (
		.din(new_net_11781),
		.dout(new_net_11782)
	);

	bfr new_net_11783_bfr_after (
		.din(new_net_11782),
		.dout(new_net_11783)
	);

	bfr new_net_11784_bfr_after (
		.din(new_net_11783),
		.dout(new_net_11784)
	);

	bfr new_net_11785_bfr_after (
		.din(new_net_11784),
		.dout(new_net_11785)
	);

	spl2 _0688__v_fanout (
		.a(new_net_11785),
		.b(new_net_102),
		.c(new_net_103)
	);

	bfr new_net_11786_bfr_after (
		.din(_0926_),
		.dout(new_net_11786)
	);

	bfr new_net_11787_bfr_after (
		.din(new_net_11786),
		.dout(new_net_11787)
	);

	bfr new_net_11788_bfr_after (
		.din(new_net_11787),
		.dout(new_net_11788)
	);

	bfr new_net_11789_bfr_after (
		.din(new_net_11788),
		.dout(new_net_11789)
	);

	bfr new_net_11790_bfr_after (
		.din(new_net_11789),
		.dout(new_net_11790)
	);

	bfr new_net_11791_bfr_after (
		.din(new_net_11790),
		.dout(new_net_11791)
	);

	bfr new_net_11792_bfr_after (
		.din(new_net_11791),
		.dout(new_net_11792)
	);

	bfr new_net_11793_bfr_after (
		.din(new_net_11792),
		.dout(new_net_11793)
	);

	bfr new_net_11794_bfr_after (
		.din(new_net_11793),
		.dout(new_net_11794)
	);

	bfr new_net_11795_bfr_after (
		.din(new_net_11794),
		.dout(new_net_11795)
	);

	bfr new_net_11796_bfr_after (
		.din(new_net_11795),
		.dout(new_net_11796)
	);

	bfr new_net_11797_bfr_after (
		.din(new_net_11796),
		.dout(new_net_11797)
	);

	bfr new_net_11798_bfr_after (
		.din(new_net_11797),
		.dout(new_net_11798)
	);

	bfr new_net_11799_bfr_after (
		.din(new_net_11798),
		.dout(new_net_11799)
	);

	bfr new_net_11800_bfr_after (
		.din(new_net_11799),
		.dout(new_net_11800)
	);

	bfr new_net_11801_bfr_after (
		.din(new_net_11800),
		.dout(new_net_11801)
	);

	bfr new_net_11802_bfr_after (
		.din(new_net_11801),
		.dout(new_net_11802)
	);

	bfr new_net_11803_bfr_after (
		.din(new_net_11802),
		.dout(new_net_11803)
	);

	bfr new_net_11804_bfr_after (
		.din(new_net_11803),
		.dout(new_net_11804)
	);

	bfr new_net_11805_bfr_after (
		.din(new_net_11804),
		.dout(new_net_11805)
	);

	bfr new_net_11806_bfr_after (
		.din(new_net_11805),
		.dout(new_net_11806)
	);

	bfr new_net_11807_bfr_after (
		.din(new_net_11806),
		.dout(new_net_11807)
	);

	bfr new_net_11808_bfr_after (
		.din(new_net_11807),
		.dout(new_net_11808)
	);

	bfr new_net_11809_bfr_after (
		.din(new_net_11808),
		.dout(new_net_11809)
	);

	bfr new_net_11810_bfr_after (
		.din(new_net_11809),
		.dout(new_net_11810)
	);

	bfr new_net_11811_bfr_after (
		.din(new_net_11810),
		.dout(new_net_11811)
	);

	bfr new_net_11812_bfr_after (
		.din(new_net_11811),
		.dout(new_net_11812)
	);

	bfr new_net_11813_bfr_after (
		.din(new_net_11812),
		.dout(new_net_11813)
	);

	bfr new_net_11814_bfr_after (
		.din(new_net_11813),
		.dout(new_net_11814)
	);

	bfr new_net_11815_bfr_after (
		.din(new_net_11814),
		.dout(new_net_11815)
	);

	bfr new_net_11816_bfr_after (
		.din(new_net_11815),
		.dout(new_net_11816)
	);

	bfr new_net_11817_bfr_after (
		.din(new_net_11816),
		.dout(new_net_11817)
	);

	bfr new_net_11818_bfr_after (
		.din(new_net_11817),
		.dout(new_net_11818)
	);

	bfr new_net_11819_bfr_after (
		.din(new_net_11818),
		.dout(new_net_11819)
	);

	bfr new_net_11820_bfr_after (
		.din(new_net_11819),
		.dout(new_net_11820)
	);

	bfr new_net_11821_bfr_after (
		.din(new_net_11820),
		.dout(new_net_11821)
	);

	bfr new_net_11822_bfr_after (
		.din(new_net_11821),
		.dout(new_net_11822)
	);

	bfr new_net_11823_bfr_after (
		.din(new_net_11822),
		.dout(new_net_11823)
	);

	bfr new_net_11824_bfr_after (
		.din(new_net_11823),
		.dout(new_net_11824)
	);

	bfr new_net_11825_bfr_after (
		.din(new_net_11824),
		.dout(new_net_11825)
	);

	bfr new_net_11826_bfr_after (
		.din(new_net_11825),
		.dout(new_net_11826)
	);

	bfr new_net_11827_bfr_after (
		.din(new_net_11826),
		.dout(new_net_11827)
	);

	bfr new_net_11828_bfr_after (
		.din(new_net_11827),
		.dout(new_net_11828)
	);

	bfr new_net_11829_bfr_after (
		.din(new_net_11828),
		.dout(new_net_11829)
	);

	bfr new_net_11830_bfr_after (
		.din(new_net_11829),
		.dout(new_net_11830)
	);

	bfr new_net_11831_bfr_after (
		.din(new_net_11830),
		.dout(new_net_11831)
	);

	bfr new_net_11832_bfr_after (
		.din(new_net_11831),
		.dout(new_net_11832)
	);

	bfr new_net_11833_bfr_after (
		.din(new_net_11832),
		.dout(new_net_11833)
	);

	bfr new_net_11834_bfr_after (
		.din(new_net_11833),
		.dout(new_net_11834)
	);

	bfr new_net_11835_bfr_after (
		.din(new_net_11834),
		.dout(new_net_11835)
	);

	bfr new_net_11836_bfr_after (
		.din(new_net_11835),
		.dout(new_net_11836)
	);

	bfr new_net_11837_bfr_after (
		.din(new_net_11836),
		.dout(new_net_11837)
	);

	bfr new_net_11838_bfr_after (
		.din(new_net_11837),
		.dout(new_net_11838)
	);

	bfr new_net_11839_bfr_after (
		.din(new_net_11838),
		.dout(new_net_11839)
	);

	bfr new_net_11840_bfr_after (
		.din(new_net_11839),
		.dout(new_net_11840)
	);

	bfr new_net_11841_bfr_after (
		.din(new_net_11840),
		.dout(new_net_11841)
	);

	bfr new_net_11842_bfr_after (
		.din(new_net_11841),
		.dout(new_net_11842)
	);

	bfr new_net_11843_bfr_after (
		.din(new_net_11842),
		.dout(new_net_11843)
	);

	bfr new_net_11844_bfr_after (
		.din(new_net_11843),
		.dout(new_net_11844)
	);

	bfr new_net_11845_bfr_after (
		.din(new_net_11844),
		.dout(new_net_11845)
	);

	bfr new_net_11846_bfr_after (
		.din(new_net_11845),
		.dout(new_net_11846)
	);

	bfr new_net_11847_bfr_after (
		.din(new_net_11846),
		.dout(new_net_11847)
	);

	bfr new_net_11848_bfr_after (
		.din(new_net_11847),
		.dout(new_net_11848)
	);

	bfr new_net_11849_bfr_after (
		.din(new_net_11848),
		.dout(new_net_11849)
	);

	bfr new_net_11850_bfr_after (
		.din(new_net_11849),
		.dout(new_net_11850)
	);

	bfr new_net_11851_bfr_after (
		.din(new_net_11850),
		.dout(new_net_11851)
	);

	bfr new_net_11852_bfr_after (
		.din(new_net_11851),
		.dout(new_net_11852)
	);

	bfr new_net_11853_bfr_after (
		.din(new_net_11852),
		.dout(new_net_11853)
	);

	bfr new_net_11854_bfr_after (
		.din(new_net_11853),
		.dout(new_net_11854)
	);

	bfr new_net_11855_bfr_after (
		.din(new_net_11854),
		.dout(new_net_11855)
	);

	bfr new_net_11856_bfr_after (
		.din(new_net_11855),
		.dout(new_net_11856)
	);

	bfr new_net_11857_bfr_after (
		.din(new_net_11856),
		.dout(new_net_11857)
	);

	bfr new_net_11858_bfr_after (
		.din(new_net_11857),
		.dout(new_net_11858)
	);

	bfr new_net_11859_bfr_after (
		.din(new_net_11858),
		.dout(new_net_11859)
	);

	bfr new_net_11860_bfr_after (
		.din(new_net_11859),
		.dout(new_net_11860)
	);

	bfr new_net_11861_bfr_after (
		.din(new_net_11860),
		.dout(new_net_11861)
	);

	bfr new_net_11862_bfr_after (
		.din(new_net_11861),
		.dout(new_net_11862)
	);

	bfr new_net_11863_bfr_after (
		.din(new_net_11862),
		.dout(new_net_11863)
	);

	bfr new_net_11864_bfr_after (
		.din(new_net_11863),
		.dout(new_net_11864)
	);

	bfr new_net_11865_bfr_after (
		.din(new_net_11864),
		.dout(new_net_11865)
	);

	bfr new_net_11866_bfr_after (
		.din(new_net_11865),
		.dout(new_net_11866)
	);

	bfr new_net_11867_bfr_after (
		.din(new_net_11866),
		.dout(new_net_11867)
	);

	bfr new_net_11868_bfr_after (
		.din(new_net_11867),
		.dout(new_net_11868)
	);

	bfr new_net_11869_bfr_after (
		.din(new_net_11868),
		.dout(new_net_11869)
	);

	bfr new_net_11870_bfr_after (
		.din(new_net_11869),
		.dout(new_net_11870)
	);

	bfr new_net_11871_bfr_after (
		.din(new_net_11870),
		.dout(new_net_11871)
	);

	bfr new_net_11872_bfr_after (
		.din(new_net_11871),
		.dout(new_net_11872)
	);

	bfr new_net_11873_bfr_after (
		.din(new_net_11872),
		.dout(new_net_11873)
	);

	bfr new_net_11874_bfr_after (
		.din(new_net_11873),
		.dout(new_net_11874)
	);

	bfr new_net_11875_bfr_after (
		.din(new_net_11874),
		.dout(new_net_11875)
	);

	bfr new_net_11876_bfr_after (
		.din(new_net_11875),
		.dout(new_net_11876)
	);

	bfr new_net_11877_bfr_after (
		.din(new_net_11876),
		.dout(new_net_11877)
	);

	bfr new_net_11878_bfr_after (
		.din(new_net_11877),
		.dout(new_net_11878)
	);

	bfr new_net_11879_bfr_after (
		.din(new_net_11878),
		.dout(new_net_11879)
	);

	bfr new_net_11880_bfr_after (
		.din(new_net_11879),
		.dout(new_net_11880)
	);

	bfr new_net_11881_bfr_after (
		.din(new_net_11880),
		.dout(new_net_11881)
	);

	bfr new_net_11882_bfr_after (
		.din(new_net_11881),
		.dout(new_net_11882)
	);

	bfr new_net_11883_bfr_after (
		.din(new_net_11882),
		.dout(new_net_11883)
	);

	bfr new_net_11884_bfr_after (
		.din(new_net_11883),
		.dout(new_net_11884)
	);

	bfr new_net_11885_bfr_after (
		.din(new_net_11884),
		.dout(new_net_11885)
	);

	bfr new_net_11886_bfr_after (
		.din(new_net_11885),
		.dout(new_net_11886)
	);

	bfr new_net_11887_bfr_after (
		.din(new_net_11886),
		.dout(new_net_11887)
	);

	bfr new_net_11888_bfr_after (
		.din(new_net_11887),
		.dout(new_net_11888)
	);

	bfr new_net_11889_bfr_after (
		.din(new_net_11888),
		.dout(new_net_11889)
	);

	bfr new_net_11890_bfr_after (
		.din(new_net_11889),
		.dout(new_net_11890)
	);

	bfr new_net_11891_bfr_after (
		.din(new_net_11890),
		.dout(new_net_11891)
	);

	bfr new_net_11892_bfr_after (
		.din(new_net_11891),
		.dout(new_net_11892)
	);

	bfr new_net_11893_bfr_after (
		.din(new_net_11892),
		.dout(new_net_11893)
	);

	bfr new_net_11894_bfr_after (
		.din(new_net_11893),
		.dout(new_net_11894)
	);

	bfr new_net_11895_bfr_after (
		.din(new_net_11894),
		.dout(new_net_11895)
	);

	bfr new_net_11896_bfr_after (
		.din(new_net_11895),
		.dout(new_net_11896)
	);

	bfr new_net_11897_bfr_after (
		.din(new_net_11896),
		.dout(new_net_11897)
	);

	spl2 _0926__v_fanout (
		.a(new_net_11897),
		.b(new_net_1114),
		.c(new_net_1115)
	);

	bfr new_net_11898_bfr_after (
		.din(_0696_),
		.dout(new_net_11898)
	);

	bfr new_net_11899_bfr_after (
		.din(new_net_11898),
		.dout(new_net_11899)
	);

	bfr new_net_11900_bfr_after (
		.din(new_net_11899),
		.dout(new_net_11900)
	);

	bfr new_net_11901_bfr_after (
		.din(new_net_11900),
		.dout(new_net_11901)
	);

	bfr new_net_11902_bfr_after (
		.din(new_net_11901),
		.dout(new_net_11902)
	);

	bfr new_net_11903_bfr_after (
		.din(new_net_11902),
		.dout(new_net_11903)
	);

	bfr new_net_11904_bfr_after (
		.din(new_net_11903),
		.dout(new_net_11904)
	);

	bfr new_net_11905_bfr_after (
		.din(new_net_11904),
		.dout(new_net_11905)
	);

	bfr new_net_11906_bfr_after (
		.din(new_net_11905),
		.dout(new_net_11906)
	);

	bfr new_net_11907_bfr_after (
		.din(new_net_11906),
		.dout(new_net_11907)
	);

	bfr new_net_11908_bfr_after (
		.din(new_net_11907),
		.dout(new_net_11908)
	);

	bfr new_net_11909_bfr_after (
		.din(new_net_11908),
		.dout(new_net_11909)
	);

	bfr new_net_11910_bfr_after (
		.din(new_net_11909),
		.dout(new_net_11910)
	);

	bfr new_net_11911_bfr_after (
		.din(new_net_11910),
		.dout(new_net_11911)
	);

	bfr new_net_11912_bfr_after (
		.din(new_net_11911),
		.dout(new_net_11912)
	);

	bfr new_net_11913_bfr_after (
		.din(new_net_11912),
		.dout(new_net_11913)
	);

	bfr new_net_11914_bfr_after (
		.din(new_net_11913),
		.dout(new_net_11914)
	);

	bfr new_net_11915_bfr_after (
		.din(new_net_11914),
		.dout(new_net_11915)
	);

	bfr new_net_11916_bfr_after (
		.din(new_net_11915),
		.dout(new_net_11916)
	);

	bfr new_net_11917_bfr_after (
		.din(new_net_11916),
		.dout(new_net_11917)
	);

	bfr new_net_11918_bfr_after (
		.din(new_net_11917),
		.dout(new_net_11918)
	);

	bfr new_net_11919_bfr_after (
		.din(new_net_11918),
		.dout(new_net_11919)
	);

	bfr new_net_11920_bfr_after (
		.din(new_net_11919),
		.dout(new_net_11920)
	);

	bfr new_net_11921_bfr_after (
		.din(new_net_11920),
		.dout(new_net_11921)
	);

	bfr new_net_11922_bfr_after (
		.din(new_net_11921),
		.dout(new_net_11922)
	);

	bfr new_net_11923_bfr_after (
		.din(new_net_11922),
		.dout(new_net_11923)
	);

	bfr new_net_11924_bfr_after (
		.din(new_net_11923),
		.dout(new_net_11924)
	);

	bfr new_net_11925_bfr_after (
		.din(new_net_11924),
		.dout(new_net_11925)
	);

	bfr new_net_11926_bfr_after (
		.din(new_net_11925),
		.dout(new_net_11926)
	);

	bfr new_net_11927_bfr_after (
		.din(new_net_11926),
		.dout(new_net_11927)
	);

	bfr new_net_11928_bfr_after (
		.din(new_net_11927),
		.dout(new_net_11928)
	);

	bfr new_net_11929_bfr_after (
		.din(new_net_11928),
		.dout(new_net_11929)
	);

	bfr new_net_11930_bfr_after (
		.din(new_net_11929),
		.dout(new_net_11930)
	);

	bfr new_net_11931_bfr_after (
		.din(new_net_11930),
		.dout(new_net_11931)
	);

	bfr new_net_11932_bfr_after (
		.din(new_net_11931),
		.dout(new_net_11932)
	);

	bfr new_net_11933_bfr_after (
		.din(new_net_11932),
		.dout(new_net_11933)
	);

	bfr new_net_11934_bfr_after (
		.din(new_net_11933),
		.dout(new_net_11934)
	);

	bfr new_net_11935_bfr_after (
		.din(new_net_11934),
		.dout(new_net_11935)
	);

	bfr new_net_11936_bfr_after (
		.din(new_net_11935),
		.dout(new_net_11936)
	);

	bfr new_net_11937_bfr_after (
		.din(new_net_11936),
		.dout(new_net_11937)
	);

	bfr new_net_11938_bfr_after (
		.din(new_net_11937),
		.dout(new_net_11938)
	);

	bfr new_net_11939_bfr_after (
		.din(new_net_11938),
		.dout(new_net_11939)
	);

	bfr new_net_11940_bfr_after (
		.din(new_net_11939),
		.dout(new_net_11940)
	);

	bfr new_net_11941_bfr_after (
		.din(new_net_11940),
		.dout(new_net_11941)
	);

	bfr new_net_11942_bfr_after (
		.din(new_net_11941),
		.dout(new_net_11942)
	);

	bfr new_net_11943_bfr_after (
		.din(new_net_11942),
		.dout(new_net_11943)
	);

	bfr new_net_11944_bfr_after (
		.din(new_net_11943),
		.dout(new_net_11944)
	);

	bfr new_net_11945_bfr_after (
		.din(new_net_11944),
		.dout(new_net_11945)
	);

	bfr new_net_11946_bfr_after (
		.din(new_net_11945),
		.dout(new_net_11946)
	);

	bfr new_net_11947_bfr_after (
		.din(new_net_11946),
		.dout(new_net_11947)
	);

	bfr new_net_11948_bfr_after (
		.din(new_net_11947),
		.dout(new_net_11948)
	);

	bfr new_net_11949_bfr_after (
		.din(new_net_11948),
		.dout(new_net_11949)
	);

	bfr new_net_11950_bfr_after (
		.din(new_net_11949),
		.dout(new_net_11950)
	);

	bfr new_net_11951_bfr_after (
		.din(new_net_11950),
		.dout(new_net_11951)
	);

	bfr new_net_11952_bfr_after (
		.din(new_net_11951),
		.dout(new_net_11952)
	);

	bfr new_net_11953_bfr_after (
		.din(new_net_11952),
		.dout(new_net_11953)
	);

	bfr new_net_11954_bfr_after (
		.din(new_net_11953),
		.dout(new_net_11954)
	);

	bfr new_net_11955_bfr_after (
		.din(new_net_11954),
		.dout(new_net_11955)
	);

	bfr new_net_11956_bfr_after (
		.din(new_net_11955),
		.dout(new_net_11956)
	);

	bfr new_net_11957_bfr_after (
		.din(new_net_11956),
		.dout(new_net_11957)
	);

	bfr new_net_11958_bfr_after (
		.din(new_net_11957),
		.dout(new_net_11958)
	);

	bfr new_net_11959_bfr_after (
		.din(new_net_11958),
		.dout(new_net_11959)
	);

	bfr new_net_11960_bfr_after (
		.din(new_net_11959),
		.dout(new_net_11960)
	);

	bfr new_net_11961_bfr_after (
		.din(new_net_11960),
		.dout(new_net_11961)
	);

	bfr new_net_11962_bfr_after (
		.din(new_net_11961),
		.dout(new_net_11962)
	);

	bfr new_net_11963_bfr_after (
		.din(new_net_11962),
		.dout(new_net_11963)
	);

	bfr new_net_11964_bfr_after (
		.din(new_net_11963),
		.dout(new_net_11964)
	);

	bfr new_net_11965_bfr_after (
		.din(new_net_11964),
		.dout(new_net_11965)
	);

	bfr new_net_11966_bfr_after (
		.din(new_net_11965),
		.dout(new_net_11966)
	);

	bfr new_net_11967_bfr_after (
		.din(new_net_11966),
		.dout(new_net_11967)
	);

	bfr new_net_11968_bfr_after (
		.din(new_net_11967),
		.dout(new_net_11968)
	);

	bfr new_net_11969_bfr_after (
		.din(new_net_11968),
		.dout(new_net_11969)
	);

	bfr new_net_11970_bfr_after (
		.din(new_net_11969),
		.dout(new_net_11970)
	);

	bfr new_net_11971_bfr_after (
		.din(new_net_11970),
		.dout(new_net_11971)
	);

	bfr new_net_11972_bfr_after (
		.din(new_net_11971),
		.dout(new_net_11972)
	);

	bfr new_net_11973_bfr_after (
		.din(new_net_11972),
		.dout(new_net_11973)
	);

	bfr new_net_11974_bfr_after (
		.din(new_net_11973),
		.dout(new_net_11974)
	);

	bfr new_net_11975_bfr_after (
		.din(new_net_11974),
		.dout(new_net_11975)
	);

	bfr new_net_11976_bfr_after (
		.din(new_net_11975),
		.dout(new_net_11976)
	);

	bfr new_net_11977_bfr_after (
		.din(new_net_11976),
		.dout(new_net_11977)
	);

	bfr new_net_11978_bfr_after (
		.din(new_net_11977),
		.dout(new_net_11978)
	);

	bfr new_net_11979_bfr_after (
		.din(new_net_11978),
		.dout(new_net_11979)
	);

	bfr new_net_11980_bfr_after (
		.din(new_net_11979),
		.dout(new_net_11980)
	);

	bfr new_net_11981_bfr_after (
		.din(new_net_11980),
		.dout(new_net_11981)
	);

	bfr new_net_11982_bfr_after (
		.din(new_net_11981),
		.dout(new_net_11982)
	);

	bfr new_net_11983_bfr_after (
		.din(new_net_11982),
		.dout(new_net_11983)
	);

	bfr new_net_11984_bfr_after (
		.din(new_net_11983),
		.dout(new_net_11984)
	);

	bfr new_net_11985_bfr_after (
		.din(new_net_11984),
		.dout(new_net_11985)
	);

	bfr new_net_11986_bfr_after (
		.din(new_net_11985),
		.dout(new_net_11986)
	);

	bfr new_net_11987_bfr_after (
		.din(new_net_11986),
		.dout(new_net_11987)
	);

	bfr new_net_11988_bfr_after (
		.din(new_net_11987),
		.dout(new_net_11988)
	);

	bfr new_net_11989_bfr_after (
		.din(new_net_11988),
		.dout(new_net_11989)
	);

	bfr new_net_11990_bfr_after (
		.din(new_net_11989),
		.dout(new_net_11990)
	);

	bfr new_net_11991_bfr_after (
		.din(new_net_11990),
		.dout(new_net_11991)
	);

	bfr new_net_11992_bfr_after (
		.din(new_net_11991),
		.dout(new_net_11992)
	);

	bfr new_net_11993_bfr_after (
		.din(new_net_11992),
		.dout(new_net_11993)
	);

	bfr new_net_11994_bfr_after (
		.din(new_net_11993),
		.dout(new_net_11994)
	);

	bfr new_net_11995_bfr_after (
		.din(new_net_11994),
		.dout(new_net_11995)
	);

	bfr new_net_11996_bfr_after (
		.din(new_net_11995),
		.dout(new_net_11996)
	);

	bfr new_net_11997_bfr_after (
		.din(new_net_11996),
		.dout(new_net_11997)
	);

	bfr new_net_11998_bfr_after (
		.din(new_net_11997),
		.dout(new_net_11998)
	);

	bfr new_net_11999_bfr_after (
		.din(new_net_11998),
		.dout(new_net_11999)
	);

	bfr new_net_12000_bfr_after (
		.din(new_net_11999),
		.dout(new_net_12000)
	);

	bfr new_net_12001_bfr_after (
		.din(new_net_12000),
		.dout(new_net_12001)
	);

	bfr new_net_12002_bfr_after (
		.din(new_net_12001),
		.dout(new_net_12002)
	);

	bfr new_net_12003_bfr_after (
		.din(new_net_12002),
		.dout(new_net_12003)
	);

	bfr new_net_12004_bfr_after (
		.din(new_net_12003),
		.dout(new_net_12004)
	);

	bfr new_net_12005_bfr_after (
		.din(new_net_12004),
		.dout(new_net_12005)
	);

	bfr new_net_12006_bfr_after (
		.din(new_net_12005),
		.dout(new_net_12006)
	);

	bfr new_net_12007_bfr_after (
		.din(new_net_12006),
		.dout(new_net_12007)
	);

	bfr new_net_12008_bfr_after (
		.din(new_net_12007),
		.dout(new_net_12008)
	);

	bfr new_net_12009_bfr_after (
		.din(new_net_12008),
		.dout(new_net_12009)
	);

	spl2 _0696__v_fanout (
		.a(new_net_12009),
		.b(new_net_362),
		.c(new_net_363)
	);

	spl2 _1502__v_fanout (
		.a(_1502_),
		.b(new_net_488),
		.c(new_net_489)
	);

	bfr new_net_12010_bfr_after (
		.din(_0241_),
		.dout(new_net_12010)
	);

	bfr new_net_12011_bfr_after (
		.din(new_net_12010),
		.dout(new_net_12011)
	);

	bfr new_net_12012_bfr_after (
		.din(new_net_12011),
		.dout(new_net_12012)
	);

	bfr new_net_12013_bfr_after (
		.din(new_net_12012),
		.dout(new_net_12013)
	);

	bfr new_net_12014_bfr_after (
		.din(new_net_12013),
		.dout(new_net_12014)
	);

	bfr new_net_12015_bfr_after (
		.din(new_net_12014),
		.dout(new_net_12015)
	);

	bfr new_net_12016_bfr_after (
		.din(new_net_12015),
		.dout(new_net_12016)
	);

	bfr new_net_12017_bfr_after (
		.din(new_net_12016),
		.dout(new_net_12017)
	);

	bfr new_net_12018_bfr_after (
		.din(new_net_12017),
		.dout(new_net_12018)
	);

	bfr new_net_12019_bfr_after (
		.din(new_net_12018),
		.dout(new_net_12019)
	);

	bfr new_net_12020_bfr_after (
		.din(new_net_12019),
		.dout(new_net_12020)
	);

	bfr new_net_12021_bfr_after (
		.din(new_net_12020),
		.dout(new_net_12021)
	);

	bfr new_net_12022_bfr_after (
		.din(new_net_12021),
		.dout(new_net_12022)
	);

	bfr new_net_12023_bfr_after (
		.din(new_net_12022),
		.dout(new_net_12023)
	);

	bfr new_net_12024_bfr_after (
		.din(new_net_12023),
		.dout(new_net_12024)
	);

	bfr new_net_12025_bfr_after (
		.din(new_net_12024),
		.dout(new_net_12025)
	);

	bfr new_net_12026_bfr_after (
		.din(new_net_12025),
		.dout(new_net_12026)
	);

	bfr new_net_12027_bfr_after (
		.din(new_net_12026),
		.dout(new_net_12027)
	);

	bfr new_net_12028_bfr_after (
		.din(new_net_12027),
		.dout(new_net_12028)
	);

	bfr new_net_12029_bfr_after (
		.din(new_net_12028),
		.dout(new_net_12029)
	);

	bfr new_net_12030_bfr_after (
		.din(new_net_12029),
		.dout(new_net_12030)
	);

	bfr new_net_12031_bfr_after (
		.din(new_net_12030),
		.dout(new_net_12031)
	);

	bfr new_net_12032_bfr_after (
		.din(new_net_12031),
		.dout(new_net_12032)
	);

	bfr new_net_12033_bfr_after (
		.din(new_net_12032),
		.dout(new_net_12033)
	);

	spl2 _0241__v_fanout (
		.a(new_net_12033),
		.b(new_net_663),
		.c(new_net_664)
	);

	bfr new_net_12034_bfr_after (
		.din(_0097_),
		.dout(new_net_12034)
	);

	bfr new_net_12035_bfr_after (
		.din(new_net_12034),
		.dout(new_net_12035)
	);

	bfr new_net_12036_bfr_after (
		.din(new_net_12035),
		.dout(new_net_12036)
	);

	bfr new_net_12037_bfr_after (
		.din(new_net_12036),
		.dout(new_net_12037)
	);

	bfr new_net_12038_bfr_after (
		.din(new_net_12037),
		.dout(new_net_12038)
	);

	bfr new_net_12039_bfr_after (
		.din(new_net_12038),
		.dout(new_net_12039)
	);

	bfr new_net_12040_bfr_after (
		.din(new_net_12039),
		.dout(new_net_12040)
	);

	bfr new_net_12041_bfr_after (
		.din(new_net_12040),
		.dout(new_net_12041)
	);

	bfr new_net_12042_bfr_after (
		.din(new_net_12041),
		.dout(new_net_12042)
	);

	bfr new_net_12043_bfr_after (
		.din(new_net_12042),
		.dout(new_net_12043)
	);

	bfr new_net_12044_bfr_after (
		.din(new_net_12043),
		.dout(new_net_12044)
	);

	bfr new_net_12045_bfr_after (
		.din(new_net_12044),
		.dout(new_net_12045)
	);

	bfr new_net_12046_bfr_after (
		.din(new_net_12045),
		.dout(new_net_12046)
	);

	bfr new_net_12047_bfr_after (
		.din(new_net_12046),
		.dout(new_net_12047)
	);

	bfr new_net_12048_bfr_after (
		.din(new_net_12047),
		.dout(new_net_12048)
	);

	bfr new_net_12049_bfr_after (
		.din(new_net_12048),
		.dout(new_net_12049)
	);

	bfr new_net_12050_bfr_after (
		.din(new_net_12049),
		.dout(new_net_12050)
	);

	bfr new_net_12051_bfr_after (
		.din(new_net_12050),
		.dout(new_net_12051)
	);

	bfr new_net_12052_bfr_after (
		.din(new_net_12051),
		.dout(new_net_12052)
	);

	bfr new_net_12053_bfr_after (
		.din(new_net_12052),
		.dout(new_net_12053)
	);

	bfr new_net_12054_bfr_after (
		.din(new_net_12053),
		.dout(new_net_12054)
	);

	bfr new_net_12055_bfr_after (
		.din(new_net_12054),
		.dout(new_net_12055)
	);

	bfr new_net_12056_bfr_after (
		.din(new_net_12055),
		.dout(new_net_12056)
	);

	bfr new_net_12057_bfr_after (
		.din(new_net_12056),
		.dout(new_net_12057)
	);

	bfr new_net_12058_bfr_after (
		.din(new_net_12057),
		.dout(new_net_12058)
	);

	bfr new_net_12059_bfr_after (
		.din(new_net_12058),
		.dout(new_net_12059)
	);

	bfr new_net_12060_bfr_after (
		.din(new_net_12059),
		.dout(new_net_12060)
	);

	bfr new_net_12061_bfr_after (
		.din(new_net_12060),
		.dout(new_net_12061)
	);

	bfr new_net_12062_bfr_after (
		.din(new_net_12061),
		.dout(new_net_12062)
	);

	bfr new_net_12063_bfr_after (
		.din(new_net_12062),
		.dout(new_net_12063)
	);

	bfr new_net_12064_bfr_after (
		.din(new_net_12063),
		.dout(new_net_12064)
	);

	bfr new_net_12065_bfr_after (
		.din(new_net_12064),
		.dout(new_net_12065)
	);

	bfr new_net_12066_bfr_after (
		.din(new_net_12065),
		.dout(new_net_12066)
	);

	bfr new_net_12067_bfr_after (
		.din(new_net_12066),
		.dout(new_net_12067)
	);

	bfr new_net_12068_bfr_after (
		.din(new_net_12067),
		.dout(new_net_12068)
	);

	bfr new_net_12069_bfr_after (
		.din(new_net_12068),
		.dout(new_net_12069)
	);

	bfr new_net_12070_bfr_after (
		.din(new_net_12069),
		.dout(new_net_12070)
	);

	bfr new_net_12071_bfr_after (
		.din(new_net_12070),
		.dout(new_net_12071)
	);

	bfr new_net_12072_bfr_after (
		.din(new_net_12071),
		.dout(new_net_12072)
	);

	bfr new_net_12073_bfr_after (
		.din(new_net_12072),
		.dout(new_net_12073)
	);

	bfr new_net_12074_bfr_after (
		.din(new_net_12073),
		.dout(new_net_12074)
	);

	bfr new_net_12075_bfr_after (
		.din(new_net_12074),
		.dout(new_net_12075)
	);

	bfr new_net_12076_bfr_after (
		.din(new_net_12075),
		.dout(new_net_12076)
	);

	bfr new_net_12077_bfr_after (
		.din(new_net_12076),
		.dout(new_net_12077)
	);

	bfr new_net_12078_bfr_after (
		.din(new_net_12077),
		.dout(new_net_12078)
	);

	bfr new_net_12079_bfr_after (
		.din(new_net_12078),
		.dout(new_net_12079)
	);

	bfr new_net_12080_bfr_after (
		.din(new_net_12079),
		.dout(new_net_12080)
	);

	bfr new_net_12081_bfr_after (
		.din(new_net_12080),
		.dout(new_net_12081)
	);

	bfr new_net_12082_bfr_after (
		.din(new_net_12081),
		.dout(new_net_12082)
	);

	bfr new_net_12083_bfr_after (
		.din(new_net_12082),
		.dout(new_net_12083)
	);

	bfr new_net_12084_bfr_after (
		.din(new_net_12083),
		.dout(new_net_12084)
	);

	bfr new_net_12085_bfr_after (
		.din(new_net_12084),
		.dout(new_net_12085)
	);

	bfr new_net_12086_bfr_after (
		.din(new_net_12085),
		.dout(new_net_12086)
	);

	bfr new_net_12087_bfr_after (
		.din(new_net_12086),
		.dout(new_net_12087)
	);

	bfr new_net_12088_bfr_after (
		.din(new_net_12087),
		.dout(new_net_12088)
	);

	bfr new_net_12089_bfr_after (
		.din(new_net_12088),
		.dout(new_net_12089)
	);

	bfr new_net_12090_bfr_after (
		.din(new_net_12089),
		.dout(new_net_12090)
	);

	bfr new_net_12091_bfr_after (
		.din(new_net_12090),
		.dout(new_net_12091)
	);

	bfr new_net_12092_bfr_after (
		.din(new_net_12091),
		.dout(new_net_12092)
	);

	bfr new_net_12093_bfr_after (
		.din(new_net_12092),
		.dout(new_net_12093)
	);

	bfr new_net_12094_bfr_after (
		.din(new_net_12093),
		.dout(new_net_12094)
	);

	bfr new_net_12095_bfr_after (
		.din(new_net_12094),
		.dout(new_net_12095)
	);

	bfr new_net_12096_bfr_after (
		.din(new_net_12095),
		.dout(new_net_12096)
	);

	bfr new_net_12097_bfr_after (
		.din(new_net_12096),
		.dout(new_net_12097)
	);

	spl2 _0097__v_fanout (
		.a(new_net_12097),
		.b(new_net_3256),
		.c(new_net_3257)
	);

	bfr new_net_12098_bfr_after (
		.din(_0225_),
		.dout(new_net_12098)
	);

	bfr new_net_12099_bfr_after (
		.din(new_net_12098),
		.dout(new_net_12099)
	);

	bfr new_net_12100_bfr_after (
		.din(new_net_12099),
		.dout(new_net_12100)
	);

	bfr new_net_12101_bfr_after (
		.din(new_net_12100),
		.dout(new_net_12101)
	);

	bfr new_net_12102_bfr_after (
		.din(new_net_12101),
		.dout(new_net_12102)
	);

	bfr new_net_12103_bfr_after (
		.din(new_net_12102),
		.dout(new_net_12103)
	);

	bfr new_net_12104_bfr_after (
		.din(new_net_12103),
		.dout(new_net_12104)
	);

	bfr new_net_12105_bfr_after (
		.din(new_net_12104),
		.dout(new_net_12105)
	);

	bfr new_net_12106_bfr_after (
		.din(new_net_12105),
		.dout(new_net_12106)
	);

	bfr new_net_12107_bfr_after (
		.din(new_net_12106),
		.dout(new_net_12107)
	);

	bfr new_net_12108_bfr_after (
		.din(new_net_12107),
		.dout(new_net_12108)
	);

	bfr new_net_12109_bfr_after (
		.din(new_net_12108),
		.dout(new_net_12109)
	);

	bfr new_net_12110_bfr_after (
		.din(new_net_12109),
		.dout(new_net_12110)
	);

	bfr new_net_12111_bfr_after (
		.din(new_net_12110),
		.dout(new_net_12111)
	);

	bfr new_net_12112_bfr_after (
		.din(new_net_12111),
		.dout(new_net_12112)
	);

	bfr new_net_12113_bfr_after (
		.din(new_net_12112),
		.dout(new_net_12113)
	);

	bfr new_net_12114_bfr_after (
		.din(new_net_12113),
		.dout(new_net_12114)
	);

	bfr new_net_12115_bfr_after (
		.din(new_net_12114),
		.dout(new_net_12115)
	);

	bfr new_net_12116_bfr_after (
		.din(new_net_12115),
		.dout(new_net_12116)
	);

	bfr new_net_12117_bfr_after (
		.din(new_net_12116),
		.dout(new_net_12117)
	);

	bfr new_net_12118_bfr_after (
		.din(new_net_12117),
		.dout(new_net_12118)
	);

	bfr new_net_12119_bfr_after (
		.din(new_net_12118),
		.dout(new_net_12119)
	);

	bfr new_net_12120_bfr_after (
		.din(new_net_12119),
		.dout(new_net_12120)
	);

	bfr new_net_12121_bfr_after (
		.din(new_net_12120),
		.dout(new_net_12121)
	);

	bfr new_net_12122_bfr_after (
		.din(new_net_12121),
		.dout(new_net_12122)
	);

	bfr new_net_12123_bfr_after (
		.din(new_net_12122),
		.dout(new_net_12123)
	);

	bfr new_net_12124_bfr_after (
		.din(new_net_12123),
		.dout(new_net_12124)
	);

	bfr new_net_12125_bfr_after (
		.din(new_net_12124),
		.dout(new_net_12125)
	);

	bfr new_net_12126_bfr_after (
		.din(new_net_12125),
		.dout(new_net_12126)
	);

	bfr new_net_12127_bfr_after (
		.din(new_net_12126),
		.dout(new_net_12127)
	);

	bfr new_net_12128_bfr_after (
		.din(new_net_12127),
		.dout(new_net_12128)
	);

	bfr new_net_12129_bfr_after (
		.din(new_net_12128),
		.dout(new_net_12129)
	);

	bfr new_net_12130_bfr_after (
		.din(new_net_12129),
		.dout(new_net_12130)
	);

	bfr new_net_12131_bfr_after (
		.din(new_net_12130),
		.dout(new_net_12131)
	);

	bfr new_net_12132_bfr_after (
		.din(new_net_12131),
		.dout(new_net_12132)
	);

	bfr new_net_12133_bfr_after (
		.din(new_net_12132),
		.dout(new_net_12133)
	);

	bfr new_net_12134_bfr_after (
		.din(new_net_12133),
		.dout(new_net_12134)
	);

	bfr new_net_12135_bfr_after (
		.din(new_net_12134),
		.dout(new_net_12135)
	);

	bfr new_net_12136_bfr_after (
		.din(new_net_12135),
		.dout(new_net_12136)
	);

	bfr new_net_12137_bfr_after (
		.din(new_net_12136),
		.dout(new_net_12137)
	);

	bfr new_net_12138_bfr_after (
		.din(new_net_12137),
		.dout(new_net_12138)
	);

	bfr new_net_12139_bfr_after (
		.din(new_net_12138),
		.dout(new_net_12139)
	);

	bfr new_net_12140_bfr_after (
		.din(new_net_12139),
		.dout(new_net_12140)
	);

	bfr new_net_12141_bfr_after (
		.din(new_net_12140),
		.dout(new_net_12141)
	);

	bfr new_net_12142_bfr_after (
		.din(new_net_12141),
		.dout(new_net_12142)
	);

	bfr new_net_12143_bfr_after (
		.din(new_net_12142),
		.dout(new_net_12143)
	);

	bfr new_net_12144_bfr_after (
		.din(new_net_12143),
		.dout(new_net_12144)
	);

	bfr new_net_12145_bfr_after (
		.din(new_net_12144),
		.dout(new_net_12145)
	);

	bfr new_net_12146_bfr_after (
		.din(new_net_12145),
		.dout(new_net_12146)
	);

	bfr new_net_12147_bfr_after (
		.din(new_net_12146),
		.dout(new_net_12147)
	);

	bfr new_net_12148_bfr_after (
		.din(new_net_12147),
		.dout(new_net_12148)
	);

	bfr new_net_12149_bfr_after (
		.din(new_net_12148),
		.dout(new_net_12149)
	);

	bfr new_net_12150_bfr_after (
		.din(new_net_12149),
		.dout(new_net_12150)
	);

	bfr new_net_12151_bfr_after (
		.din(new_net_12150),
		.dout(new_net_12151)
	);

	bfr new_net_12152_bfr_after (
		.din(new_net_12151),
		.dout(new_net_12152)
	);

	bfr new_net_12153_bfr_after (
		.din(new_net_12152),
		.dout(new_net_12153)
	);

	bfr new_net_12154_bfr_after (
		.din(new_net_12153),
		.dout(new_net_12154)
	);

	bfr new_net_12155_bfr_after (
		.din(new_net_12154),
		.dout(new_net_12155)
	);

	bfr new_net_12156_bfr_after (
		.din(new_net_12155),
		.dout(new_net_12156)
	);

	bfr new_net_12157_bfr_after (
		.din(new_net_12156),
		.dout(new_net_12157)
	);

	bfr new_net_12158_bfr_after (
		.din(new_net_12157),
		.dout(new_net_12158)
	);

	bfr new_net_12159_bfr_after (
		.din(new_net_12158),
		.dout(new_net_12159)
	);

	bfr new_net_12160_bfr_after (
		.din(new_net_12159),
		.dout(new_net_12160)
	);

	bfr new_net_12161_bfr_after (
		.din(new_net_12160),
		.dout(new_net_12161)
	);

	spl2 _0225__v_fanout (
		.a(new_net_12161),
		.b(new_net_1491),
		.c(new_net_1492)
	);

	bfr new_net_12162_bfr_after (
		.din(_1575_),
		.dout(new_net_12162)
	);

	bfr new_net_12163_bfr_after (
		.din(new_net_12162),
		.dout(new_net_12163)
	);

	bfr new_net_12164_bfr_after (
		.din(new_net_12163),
		.dout(new_net_12164)
	);

	bfr new_net_12165_bfr_after (
		.din(new_net_12164),
		.dout(new_net_12165)
	);

	bfr new_net_12166_bfr_after (
		.din(new_net_12165),
		.dout(new_net_12166)
	);

	bfr new_net_12167_bfr_after (
		.din(new_net_12166),
		.dout(new_net_12167)
	);

	bfr new_net_12168_bfr_after (
		.din(new_net_12167),
		.dout(new_net_12168)
	);

	bfr new_net_12169_bfr_after (
		.din(new_net_12168),
		.dout(new_net_12169)
	);

	bfr new_net_12170_bfr_after (
		.din(new_net_12169),
		.dout(new_net_12170)
	);

	bfr new_net_12171_bfr_after (
		.din(new_net_12170),
		.dout(new_net_12171)
	);

	bfr new_net_12172_bfr_after (
		.din(new_net_12171),
		.dout(new_net_12172)
	);

	bfr new_net_12173_bfr_after (
		.din(new_net_12172),
		.dout(new_net_12173)
	);

	bfr new_net_12174_bfr_after (
		.din(new_net_12173),
		.dout(new_net_12174)
	);

	bfr new_net_12175_bfr_after (
		.din(new_net_12174),
		.dout(new_net_12175)
	);

	bfr new_net_12176_bfr_after (
		.din(new_net_12175),
		.dout(new_net_12176)
	);

	bfr new_net_12177_bfr_after (
		.din(new_net_12176),
		.dout(new_net_12177)
	);

	bfr new_net_12178_bfr_after (
		.din(new_net_12177),
		.dout(new_net_12178)
	);

	bfr new_net_12179_bfr_after (
		.din(new_net_12178),
		.dout(new_net_12179)
	);

	bfr new_net_12180_bfr_after (
		.din(new_net_12179),
		.dout(new_net_12180)
	);

	bfr new_net_12181_bfr_after (
		.din(new_net_12180),
		.dout(new_net_12181)
	);

	bfr new_net_12182_bfr_after (
		.din(new_net_12181),
		.dout(new_net_12182)
	);

	bfr new_net_12183_bfr_after (
		.din(new_net_12182),
		.dout(new_net_12183)
	);

	bfr new_net_12184_bfr_after (
		.din(new_net_12183),
		.dout(new_net_12184)
	);

	bfr new_net_12185_bfr_after (
		.din(new_net_12184),
		.dout(new_net_12185)
	);

	bfr new_net_12186_bfr_after (
		.din(new_net_12185),
		.dout(new_net_12186)
	);

	bfr new_net_12187_bfr_after (
		.din(new_net_12186),
		.dout(new_net_12187)
	);

	bfr new_net_12188_bfr_after (
		.din(new_net_12187),
		.dout(new_net_12188)
	);

	bfr new_net_12189_bfr_after (
		.din(new_net_12188),
		.dout(new_net_12189)
	);

	bfr new_net_12190_bfr_after (
		.din(new_net_12189),
		.dout(new_net_12190)
	);

	bfr new_net_12191_bfr_after (
		.din(new_net_12190),
		.dout(new_net_12191)
	);

	bfr new_net_12192_bfr_after (
		.din(new_net_12191),
		.dout(new_net_12192)
	);

	bfr new_net_12193_bfr_after (
		.din(new_net_12192),
		.dout(new_net_12193)
	);

	bfr new_net_12194_bfr_after (
		.din(new_net_12193),
		.dout(new_net_12194)
	);

	bfr new_net_12195_bfr_after (
		.din(new_net_12194),
		.dout(new_net_12195)
	);

	bfr new_net_12196_bfr_after (
		.din(new_net_12195),
		.dout(new_net_12196)
	);

	bfr new_net_12197_bfr_after (
		.din(new_net_12196),
		.dout(new_net_12197)
	);

	bfr new_net_12198_bfr_after (
		.din(new_net_12197),
		.dout(new_net_12198)
	);

	bfr new_net_12199_bfr_after (
		.din(new_net_12198),
		.dout(new_net_12199)
	);

	bfr new_net_12200_bfr_after (
		.din(new_net_12199),
		.dout(new_net_12200)
	);

	bfr new_net_12201_bfr_after (
		.din(new_net_12200),
		.dout(new_net_12201)
	);

	bfr new_net_12202_bfr_after (
		.din(new_net_12201),
		.dout(new_net_12202)
	);

	bfr new_net_12203_bfr_after (
		.din(new_net_12202),
		.dout(new_net_12203)
	);

	bfr new_net_12204_bfr_after (
		.din(new_net_12203),
		.dout(new_net_12204)
	);

	bfr new_net_12205_bfr_after (
		.din(new_net_12204),
		.dout(new_net_12205)
	);

	bfr new_net_12206_bfr_after (
		.din(new_net_12205),
		.dout(new_net_12206)
	);

	bfr new_net_12207_bfr_after (
		.din(new_net_12206),
		.dout(new_net_12207)
	);

	bfr new_net_12208_bfr_after (
		.din(new_net_12207),
		.dout(new_net_12208)
	);

	bfr new_net_12209_bfr_after (
		.din(new_net_12208),
		.dout(new_net_12209)
	);

	spl2 _1575__v_fanout (
		.a(new_net_12209),
		.b(new_net_2132),
		.c(new_net_2133)
	);

	bfr new_net_12210_bfr_after (
		.din(_0889_),
		.dout(new_net_12210)
	);

	bfr new_net_12211_bfr_after (
		.din(new_net_12210),
		.dout(new_net_12211)
	);

	bfr new_net_12212_bfr_after (
		.din(new_net_12211),
		.dout(new_net_12212)
	);

	bfr new_net_12213_bfr_after (
		.din(new_net_12212),
		.dout(new_net_12213)
	);

	bfr new_net_12214_bfr_after (
		.din(new_net_12213),
		.dout(new_net_12214)
	);

	bfr new_net_12215_bfr_after (
		.din(new_net_12214),
		.dout(new_net_12215)
	);

	bfr new_net_12216_bfr_after (
		.din(new_net_12215),
		.dout(new_net_12216)
	);

	bfr new_net_12217_bfr_after (
		.din(new_net_12216),
		.dout(new_net_12217)
	);

	bfr new_net_12218_bfr_after (
		.din(new_net_12217),
		.dout(new_net_12218)
	);

	bfr new_net_12219_bfr_after (
		.din(new_net_12218),
		.dout(new_net_12219)
	);

	bfr new_net_12220_bfr_after (
		.din(new_net_12219),
		.dout(new_net_12220)
	);

	bfr new_net_12221_bfr_after (
		.din(new_net_12220),
		.dout(new_net_12221)
	);

	bfr new_net_12222_bfr_after (
		.din(new_net_12221),
		.dout(new_net_12222)
	);

	bfr new_net_12223_bfr_after (
		.din(new_net_12222),
		.dout(new_net_12223)
	);

	bfr new_net_12224_bfr_after (
		.din(new_net_12223),
		.dout(new_net_12224)
	);

	bfr new_net_12225_bfr_after (
		.din(new_net_12224),
		.dout(new_net_12225)
	);

	bfr new_net_12226_bfr_after (
		.din(new_net_12225),
		.dout(new_net_12226)
	);

	bfr new_net_12227_bfr_after (
		.din(new_net_12226),
		.dout(new_net_12227)
	);

	bfr new_net_12228_bfr_after (
		.din(new_net_12227),
		.dout(new_net_12228)
	);

	bfr new_net_12229_bfr_after (
		.din(new_net_12228),
		.dout(new_net_12229)
	);

	bfr new_net_12230_bfr_after (
		.din(new_net_12229),
		.dout(new_net_12230)
	);

	bfr new_net_12231_bfr_after (
		.din(new_net_12230),
		.dout(new_net_12231)
	);

	bfr new_net_12232_bfr_after (
		.din(new_net_12231),
		.dout(new_net_12232)
	);

	bfr new_net_12233_bfr_after (
		.din(new_net_12232),
		.dout(new_net_12233)
	);

	bfr new_net_12234_bfr_after (
		.din(new_net_12233),
		.dout(new_net_12234)
	);

	bfr new_net_12235_bfr_after (
		.din(new_net_12234),
		.dout(new_net_12235)
	);

	bfr new_net_12236_bfr_after (
		.din(new_net_12235),
		.dout(new_net_12236)
	);

	bfr new_net_12237_bfr_after (
		.din(new_net_12236),
		.dout(new_net_12237)
	);

	bfr new_net_12238_bfr_after (
		.din(new_net_12237),
		.dout(new_net_12238)
	);

	bfr new_net_12239_bfr_after (
		.din(new_net_12238),
		.dout(new_net_12239)
	);

	bfr new_net_12240_bfr_after (
		.din(new_net_12239),
		.dout(new_net_12240)
	);

	bfr new_net_12241_bfr_after (
		.din(new_net_12240),
		.dout(new_net_12241)
	);

	bfr new_net_12242_bfr_after (
		.din(new_net_12241),
		.dout(new_net_12242)
	);

	bfr new_net_12243_bfr_after (
		.din(new_net_12242),
		.dout(new_net_12243)
	);

	bfr new_net_12244_bfr_after (
		.din(new_net_12243),
		.dout(new_net_12244)
	);

	bfr new_net_12245_bfr_after (
		.din(new_net_12244),
		.dout(new_net_12245)
	);

	bfr new_net_12246_bfr_after (
		.din(new_net_12245),
		.dout(new_net_12246)
	);

	bfr new_net_12247_bfr_after (
		.din(new_net_12246),
		.dout(new_net_12247)
	);

	bfr new_net_12248_bfr_after (
		.din(new_net_12247),
		.dout(new_net_12248)
	);

	bfr new_net_12249_bfr_after (
		.din(new_net_12248),
		.dout(new_net_12249)
	);

	bfr new_net_12250_bfr_after (
		.din(new_net_12249),
		.dout(new_net_12250)
	);

	bfr new_net_12251_bfr_after (
		.din(new_net_12250),
		.dout(new_net_12251)
	);

	bfr new_net_12252_bfr_after (
		.din(new_net_12251),
		.dout(new_net_12252)
	);

	bfr new_net_12253_bfr_after (
		.din(new_net_12252),
		.dout(new_net_12253)
	);

	bfr new_net_12254_bfr_after (
		.din(new_net_12253),
		.dout(new_net_12254)
	);

	bfr new_net_12255_bfr_after (
		.din(new_net_12254),
		.dout(new_net_12255)
	);

	bfr new_net_12256_bfr_after (
		.din(new_net_12255),
		.dout(new_net_12256)
	);

	bfr new_net_12257_bfr_after (
		.din(new_net_12256),
		.dout(new_net_12257)
	);

	bfr new_net_12258_bfr_after (
		.din(new_net_12257),
		.dout(new_net_12258)
	);

	bfr new_net_12259_bfr_after (
		.din(new_net_12258),
		.dout(new_net_12259)
	);

	bfr new_net_12260_bfr_after (
		.din(new_net_12259),
		.dout(new_net_12260)
	);

	bfr new_net_12261_bfr_after (
		.din(new_net_12260),
		.dout(new_net_12261)
	);

	bfr new_net_12262_bfr_after (
		.din(new_net_12261),
		.dout(new_net_12262)
	);

	bfr new_net_12263_bfr_after (
		.din(new_net_12262),
		.dout(new_net_12263)
	);

	bfr new_net_12264_bfr_after (
		.din(new_net_12263),
		.dout(new_net_12264)
	);

	bfr new_net_12265_bfr_after (
		.din(new_net_12264),
		.dout(new_net_12265)
	);

	bfr new_net_12266_bfr_after (
		.din(new_net_12265),
		.dout(new_net_12266)
	);

	bfr new_net_12267_bfr_after (
		.din(new_net_12266),
		.dout(new_net_12267)
	);

	bfr new_net_12268_bfr_after (
		.din(new_net_12267),
		.dout(new_net_12268)
	);

	bfr new_net_12269_bfr_after (
		.din(new_net_12268),
		.dout(new_net_12269)
	);

	bfr new_net_12270_bfr_after (
		.din(new_net_12269),
		.dout(new_net_12270)
	);

	bfr new_net_12271_bfr_after (
		.din(new_net_12270),
		.dout(new_net_12271)
	);

	bfr new_net_12272_bfr_after (
		.din(new_net_12271),
		.dout(new_net_12272)
	);

	bfr new_net_12273_bfr_after (
		.din(new_net_12272),
		.dout(new_net_12273)
	);

	bfr new_net_12274_bfr_after (
		.din(new_net_12273),
		.dout(new_net_12274)
	);

	bfr new_net_12275_bfr_after (
		.din(new_net_12274),
		.dout(new_net_12275)
	);

	bfr new_net_12276_bfr_after (
		.din(new_net_12275),
		.dout(new_net_12276)
	);

	bfr new_net_12277_bfr_after (
		.din(new_net_12276),
		.dout(new_net_12277)
	);

	bfr new_net_12278_bfr_after (
		.din(new_net_12277),
		.dout(new_net_12278)
	);

	bfr new_net_12279_bfr_after (
		.din(new_net_12278),
		.dout(new_net_12279)
	);

	bfr new_net_12280_bfr_after (
		.din(new_net_12279),
		.dout(new_net_12280)
	);

	bfr new_net_12281_bfr_after (
		.din(new_net_12280),
		.dout(new_net_12281)
	);

	bfr new_net_12282_bfr_after (
		.din(new_net_12281),
		.dout(new_net_12282)
	);

	bfr new_net_12283_bfr_after (
		.din(new_net_12282),
		.dout(new_net_12283)
	);

	bfr new_net_12284_bfr_after (
		.din(new_net_12283),
		.dout(new_net_12284)
	);

	bfr new_net_12285_bfr_after (
		.din(new_net_12284),
		.dout(new_net_12285)
	);

	bfr new_net_12286_bfr_after (
		.din(new_net_12285),
		.dout(new_net_12286)
	);

	bfr new_net_12287_bfr_after (
		.din(new_net_12286),
		.dout(new_net_12287)
	);

	spl2 _0889__v_fanout (
		.a(new_net_12287),
		.b(new_net_1714),
		.c(new_net_1715)
	);

	bfr new_net_12288_bfr_after (
		.din(_1689_),
		.dout(new_net_12288)
	);

	bfr new_net_12289_bfr_after (
		.din(new_net_12288),
		.dout(new_net_12289)
	);

	bfr new_net_12290_bfr_after (
		.din(new_net_12289),
		.dout(new_net_12290)
	);

	bfr new_net_12291_bfr_after (
		.din(new_net_12290),
		.dout(new_net_12291)
	);

	bfr new_net_12292_bfr_after (
		.din(new_net_12291),
		.dout(new_net_12292)
	);

	bfr new_net_12293_bfr_after (
		.din(new_net_12292),
		.dout(new_net_12293)
	);

	bfr new_net_12294_bfr_after (
		.din(new_net_12293),
		.dout(new_net_12294)
	);

	bfr new_net_12295_bfr_after (
		.din(new_net_12294),
		.dout(new_net_12295)
	);

	bfr new_net_12296_bfr_after (
		.din(new_net_12295),
		.dout(new_net_12296)
	);

	bfr new_net_12297_bfr_after (
		.din(new_net_12296),
		.dout(new_net_12297)
	);

	bfr new_net_12298_bfr_after (
		.din(new_net_12297),
		.dout(new_net_12298)
	);

	bfr new_net_12299_bfr_after (
		.din(new_net_12298),
		.dout(new_net_12299)
	);

	bfr new_net_12300_bfr_after (
		.din(new_net_12299),
		.dout(new_net_12300)
	);

	bfr new_net_12301_bfr_after (
		.din(new_net_12300),
		.dout(new_net_12301)
	);

	bfr new_net_12302_bfr_after (
		.din(new_net_12301),
		.dout(new_net_12302)
	);

	bfr new_net_12303_bfr_after (
		.din(new_net_12302),
		.dout(new_net_12303)
	);

	bfr new_net_12304_bfr_after (
		.din(new_net_12303),
		.dout(new_net_12304)
	);

	bfr new_net_12305_bfr_after (
		.din(new_net_12304),
		.dout(new_net_12305)
	);

	bfr new_net_12306_bfr_after (
		.din(new_net_12305),
		.dout(new_net_12306)
	);

	bfr new_net_12307_bfr_after (
		.din(new_net_12306),
		.dout(new_net_12307)
	);

	bfr new_net_12308_bfr_after (
		.din(new_net_12307),
		.dout(new_net_12308)
	);

	bfr new_net_12309_bfr_after (
		.din(new_net_12308),
		.dout(new_net_12309)
	);

	bfr new_net_12310_bfr_after (
		.din(new_net_12309),
		.dout(new_net_12310)
	);

	bfr new_net_12311_bfr_after (
		.din(new_net_12310),
		.dout(new_net_12311)
	);

	bfr new_net_12312_bfr_after (
		.din(new_net_12311),
		.dout(new_net_12312)
	);

	bfr new_net_12313_bfr_after (
		.din(new_net_12312),
		.dout(new_net_12313)
	);

	bfr new_net_12314_bfr_after (
		.din(new_net_12313),
		.dout(new_net_12314)
	);

	bfr new_net_12315_bfr_after (
		.din(new_net_12314),
		.dout(new_net_12315)
	);

	bfr new_net_12316_bfr_after (
		.din(new_net_12315),
		.dout(new_net_12316)
	);

	bfr new_net_12317_bfr_after (
		.din(new_net_12316),
		.dout(new_net_12317)
	);

	bfr new_net_12318_bfr_after (
		.din(new_net_12317),
		.dout(new_net_12318)
	);

	bfr new_net_12319_bfr_after (
		.din(new_net_12318),
		.dout(new_net_12319)
	);

	bfr new_net_12320_bfr_after (
		.din(new_net_12319),
		.dout(new_net_12320)
	);

	bfr new_net_12321_bfr_after (
		.din(new_net_12320),
		.dout(new_net_12321)
	);

	bfr new_net_12322_bfr_after (
		.din(new_net_12321),
		.dout(new_net_12322)
	);

	bfr new_net_12323_bfr_after (
		.din(new_net_12322),
		.dout(new_net_12323)
	);

	bfr new_net_12324_bfr_after (
		.din(new_net_12323),
		.dout(new_net_12324)
	);

	bfr new_net_12325_bfr_after (
		.din(new_net_12324),
		.dout(new_net_12325)
	);

	bfr new_net_12326_bfr_after (
		.din(new_net_12325),
		.dout(new_net_12326)
	);

	bfr new_net_12327_bfr_after (
		.din(new_net_12326),
		.dout(new_net_12327)
	);

	bfr new_net_12328_bfr_after (
		.din(new_net_12327),
		.dout(new_net_12328)
	);

	bfr new_net_12329_bfr_after (
		.din(new_net_12328),
		.dout(new_net_12329)
	);

	bfr new_net_12330_bfr_after (
		.din(new_net_12329),
		.dout(new_net_12330)
	);

	bfr new_net_12331_bfr_after (
		.din(new_net_12330),
		.dout(new_net_12331)
	);

	bfr new_net_12332_bfr_after (
		.din(new_net_12331),
		.dout(new_net_12332)
	);

	bfr new_net_12333_bfr_after (
		.din(new_net_12332),
		.dout(new_net_12333)
	);

	bfr new_net_12334_bfr_after (
		.din(new_net_12333),
		.dout(new_net_12334)
	);

	bfr new_net_12335_bfr_after (
		.din(new_net_12334),
		.dout(new_net_12335)
	);

	bfr new_net_12336_bfr_after (
		.din(new_net_12335),
		.dout(new_net_12336)
	);

	bfr new_net_12337_bfr_after (
		.din(new_net_12336),
		.dout(new_net_12337)
	);

	bfr new_net_12338_bfr_after (
		.din(new_net_12337),
		.dout(new_net_12338)
	);

	bfr new_net_12339_bfr_after (
		.din(new_net_12338),
		.dout(new_net_12339)
	);

	bfr new_net_12340_bfr_after (
		.din(new_net_12339),
		.dout(new_net_12340)
	);

	bfr new_net_12341_bfr_after (
		.din(new_net_12340),
		.dout(new_net_12341)
	);

	bfr new_net_12342_bfr_after (
		.din(new_net_12341),
		.dout(new_net_12342)
	);

	bfr new_net_12343_bfr_after (
		.din(new_net_12342),
		.dout(new_net_12343)
	);

	bfr new_net_12344_bfr_after (
		.din(new_net_12343),
		.dout(new_net_12344)
	);

	bfr new_net_12345_bfr_after (
		.din(new_net_12344),
		.dout(new_net_12345)
	);

	bfr new_net_12346_bfr_after (
		.din(new_net_12345),
		.dout(new_net_12346)
	);

	bfr new_net_12347_bfr_after (
		.din(new_net_12346),
		.dout(new_net_12347)
	);

	bfr new_net_12348_bfr_after (
		.din(new_net_12347),
		.dout(new_net_12348)
	);

	bfr new_net_12349_bfr_after (
		.din(new_net_12348),
		.dout(new_net_12349)
	);

	bfr new_net_12350_bfr_after (
		.din(new_net_12349),
		.dout(new_net_12350)
	);

	bfr new_net_12351_bfr_after (
		.din(new_net_12350),
		.dout(new_net_12351)
	);

	bfr new_net_12352_bfr_after (
		.din(new_net_12351),
		.dout(new_net_12352)
	);

	bfr new_net_12353_bfr_after (
		.din(new_net_12352),
		.dout(new_net_12353)
	);

	bfr new_net_12354_bfr_after (
		.din(new_net_12353),
		.dout(new_net_12354)
	);

	bfr new_net_12355_bfr_after (
		.din(new_net_12354),
		.dout(new_net_12355)
	);

	bfr new_net_12356_bfr_after (
		.din(new_net_12355),
		.dout(new_net_12356)
	);

	bfr new_net_12357_bfr_after (
		.din(new_net_12356),
		.dout(new_net_12357)
	);

	bfr new_net_12358_bfr_after (
		.din(new_net_12357),
		.dout(new_net_12358)
	);

	bfr new_net_12359_bfr_after (
		.din(new_net_12358),
		.dout(new_net_12359)
	);

	spl2 _1689__v_fanout (
		.a(new_net_12359),
		.b(new_net_584),
		.c(new_net_585)
	);

	spl2 _1384__v_fanout (
		.a(_1384_),
		.b(new_net_958),
		.c(new_net_959)
	);

	bfr new_net_12360_bfr_after (
		.din(_0881_),
		.dout(new_net_12360)
	);

	bfr new_net_12361_bfr_after (
		.din(new_net_12360),
		.dout(new_net_12361)
	);

	bfr new_net_12362_bfr_after (
		.din(new_net_12361),
		.dout(new_net_12362)
	);

	bfr new_net_12363_bfr_after (
		.din(new_net_12362),
		.dout(new_net_12363)
	);

	bfr new_net_12364_bfr_after (
		.din(new_net_12363),
		.dout(new_net_12364)
	);

	bfr new_net_12365_bfr_after (
		.din(new_net_12364),
		.dout(new_net_12365)
	);

	bfr new_net_12366_bfr_after (
		.din(new_net_12365),
		.dout(new_net_12366)
	);

	bfr new_net_12367_bfr_after (
		.din(new_net_12366),
		.dout(new_net_12367)
	);

	bfr new_net_12368_bfr_after (
		.din(new_net_12367),
		.dout(new_net_12368)
	);

	bfr new_net_12369_bfr_after (
		.din(new_net_12368),
		.dout(new_net_12369)
	);

	bfr new_net_12370_bfr_after (
		.din(new_net_12369),
		.dout(new_net_12370)
	);

	bfr new_net_12371_bfr_after (
		.din(new_net_12370),
		.dout(new_net_12371)
	);

	bfr new_net_12372_bfr_after (
		.din(new_net_12371),
		.dout(new_net_12372)
	);

	bfr new_net_12373_bfr_after (
		.din(new_net_12372),
		.dout(new_net_12373)
	);

	bfr new_net_12374_bfr_after (
		.din(new_net_12373),
		.dout(new_net_12374)
	);

	bfr new_net_12375_bfr_after (
		.din(new_net_12374),
		.dout(new_net_12375)
	);

	bfr new_net_12376_bfr_after (
		.din(new_net_12375),
		.dout(new_net_12376)
	);

	bfr new_net_12377_bfr_after (
		.din(new_net_12376),
		.dout(new_net_12377)
	);

	bfr new_net_12378_bfr_after (
		.din(new_net_12377),
		.dout(new_net_12378)
	);

	bfr new_net_12379_bfr_after (
		.din(new_net_12378),
		.dout(new_net_12379)
	);

	bfr new_net_12380_bfr_after (
		.din(new_net_12379),
		.dout(new_net_12380)
	);

	bfr new_net_12381_bfr_after (
		.din(new_net_12380),
		.dout(new_net_12381)
	);

	bfr new_net_12382_bfr_after (
		.din(new_net_12381),
		.dout(new_net_12382)
	);

	bfr new_net_12383_bfr_after (
		.din(new_net_12382),
		.dout(new_net_12383)
	);

	bfr new_net_12384_bfr_after (
		.din(new_net_12383),
		.dout(new_net_12384)
	);

	bfr new_net_12385_bfr_after (
		.din(new_net_12384),
		.dout(new_net_12385)
	);

	bfr new_net_12386_bfr_after (
		.din(new_net_12385),
		.dout(new_net_12386)
	);

	bfr new_net_12387_bfr_after (
		.din(new_net_12386),
		.dout(new_net_12387)
	);

	bfr new_net_12388_bfr_after (
		.din(new_net_12387),
		.dout(new_net_12388)
	);

	bfr new_net_12389_bfr_after (
		.din(new_net_12388),
		.dout(new_net_12389)
	);

	bfr new_net_12390_bfr_after (
		.din(new_net_12389),
		.dout(new_net_12390)
	);

	bfr new_net_12391_bfr_after (
		.din(new_net_12390),
		.dout(new_net_12391)
	);

	bfr new_net_12392_bfr_after (
		.din(new_net_12391),
		.dout(new_net_12392)
	);

	bfr new_net_12393_bfr_after (
		.din(new_net_12392),
		.dout(new_net_12393)
	);

	bfr new_net_12394_bfr_after (
		.din(new_net_12393),
		.dout(new_net_12394)
	);

	bfr new_net_12395_bfr_after (
		.din(new_net_12394),
		.dout(new_net_12395)
	);

	bfr new_net_12396_bfr_after (
		.din(new_net_12395),
		.dout(new_net_12396)
	);

	bfr new_net_12397_bfr_after (
		.din(new_net_12396),
		.dout(new_net_12397)
	);

	bfr new_net_12398_bfr_after (
		.din(new_net_12397),
		.dout(new_net_12398)
	);

	bfr new_net_12399_bfr_after (
		.din(new_net_12398),
		.dout(new_net_12399)
	);

	bfr new_net_12400_bfr_after (
		.din(new_net_12399),
		.dout(new_net_12400)
	);

	bfr new_net_12401_bfr_after (
		.din(new_net_12400),
		.dout(new_net_12401)
	);

	bfr new_net_12402_bfr_after (
		.din(new_net_12401),
		.dout(new_net_12402)
	);

	bfr new_net_12403_bfr_after (
		.din(new_net_12402),
		.dout(new_net_12403)
	);

	bfr new_net_12404_bfr_after (
		.din(new_net_12403),
		.dout(new_net_12404)
	);

	bfr new_net_12405_bfr_after (
		.din(new_net_12404),
		.dout(new_net_12405)
	);

	bfr new_net_12406_bfr_after (
		.din(new_net_12405),
		.dout(new_net_12406)
	);

	bfr new_net_12407_bfr_after (
		.din(new_net_12406),
		.dout(new_net_12407)
	);

	bfr new_net_12408_bfr_after (
		.din(new_net_12407),
		.dout(new_net_12408)
	);

	bfr new_net_12409_bfr_after (
		.din(new_net_12408),
		.dout(new_net_12409)
	);

	bfr new_net_12410_bfr_after (
		.din(new_net_12409),
		.dout(new_net_12410)
	);

	bfr new_net_12411_bfr_after (
		.din(new_net_12410),
		.dout(new_net_12411)
	);

	bfr new_net_12412_bfr_after (
		.din(new_net_12411),
		.dout(new_net_12412)
	);

	bfr new_net_12413_bfr_after (
		.din(new_net_12412),
		.dout(new_net_12413)
	);

	bfr new_net_12414_bfr_after (
		.din(new_net_12413),
		.dout(new_net_12414)
	);

	bfr new_net_12415_bfr_after (
		.din(new_net_12414),
		.dout(new_net_12415)
	);

	bfr new_net_12416_bfr_after (
		.din(new_net_12415),
		.dout(new_net_12416)
	);

	bfr new_net_12417_bfr_after (
		.din(new_net_12416),
		.dout(new_net_12417)
	);

	bfr new_net_12418_bfr_after (
		.din(new_net_12417),
		.dout(new_net_12418)
	);

	bfr new_net_12419_bfr_after (
		.din(new_net_12418),
		.dout(new_net_12419)
	);

	bfr new_net_12420_bfr_after (
		.din(new_net_12419),
		.dout(new_net_12420)
	);

	bfr new_net_12421_bfr_after (
		.din(new_net_12420),
		.dout(new_net_12421)
	);

	bfr new_net_12422_bfr_after (
		.din(new_net_12421),
		.dout(new_net_12422)
	);

	bfr new_net_12423_bfr_after (
		.din(new_net_12422),
		.dout(new_net_12423)
	);

	bfr new_net_12424_bfr_after (
		.din(new_net_12423),
		.dout(new_net_12424)
	);

	bfr new_net_12425_bfr_after (
		.din(new_net_12424),
		.dout(new_net_12425)
	);

	bfr new_net_12426_bfr_after (
		.din(new_net_12425),
		.dout(new_net_12426)
	);

	bfr new_net_12427_bfr_after (
		.din(new_net_12426),
		.dout(new_net_12427)
	);

	bfr new_net_12428_bfr_after (
		.din(new_net_12427),
		.dout(new_net_12428)
	);

	bfr new_net_12429_bfr_after (
		.din(new_net_12428),
		.dout(new_net_12429)
	);

	bfr new_net_12430_bfr_after (
		.din(new_net_12429),
		.dout(new_net_12430)
	);

	bfr new_net_12431_bfr_after (
		.din(new_net_12430),
		.dout(new_net_12431)
	);

	bfr new_net_12432_bfr_after (
		.din(new_net_12431),
		.dout(new_net_12432)
	);

	bfr new_net_12433_bfr_after (
		.din(new_net_12432),
		.dout(new_net_12433)
	);

	bfr new_net_12434_bfr_after (
		.din(new_net_12433),
		.dout(new_net_12434)
	);

	bfr new_net_12435_bfr_after (
		.din(new_net_12434),
		.dout(new_net_12435)
	);

	bfr new_net_12436_bfr_after (
		.din(new_net_12435),
		.dout(new_net_12436)
	);

	bfr new_net_12437_bfr_after (
		.din(new_net_12436),
		.dout(new_net_12437)
	);

	bfr new_net_12438_bfr_after (
		.din(new_net_12437),
		.dout(new_net_12438)
	);

	bfr new_net_12439_bfr_after (
		.din(new_net_12438),
		.dout(new_net_12439)
	);

	bfr new_net_12440_bfr_after (
		.din(new_net_12439),
		.dout(new_net_12440)
	);

	bfr new_net_12441_bfr_after (
		.din(new_net_12440),
		.dout(new_net_12441)
	);

	bfr new_net_12442_bfr_after (
		.din(new_net_12441),
		.dout(new_net_12442)
	);

	bfr new_net_12443_bfr_after (
		.din(new_net_12442),
		.dout(new_net_12443)
	);

	bfr new_net_12444_bfr_after (
		.din(new_net_12443),
		.dout(new_net_12444)
	);

	bfr new_net_12445_bfr_after (
		.din(new_net_12444),
		.dout(new_net_12445)
	);

	bfr new_net_12446_bfr_after (
		.din(new_net_12445),
		.dout(new_net_12446)
	);

	bfr new_net_12447_bfr_after (
		.din(new_net_12446),
		.dout(new_net_12447)
	);

	bfr new_net_12448_bfr_after (
		.din(new_net_12447),
		.dout(new_net_12448)
	);

	bfr new_net_12449_bfr_after (
		.din(new_net_12448),
		.dout(new_net_12449)
	);

	bfr new_net_12450_bfr_after (
		.din(new_net_12449),
		.dout(new_net_12450)
	);

	bfr new_net_12451_bfr_after (
		.din(new_net_12450),
		.dout(new_net_12451)
	);

	bfr new_net_12452_bfr_after (
		.din(new_net_12451),
		.dout(new_net_12452)
	);

	bfr new_net_12453_bfr_after (
		.din(new_net_12452),
		.dout(new_net_12453)
	);

	bfr new_net_12454_bfr_after (
		.din(new_net_12453),
		.dout(new_net_12454)
	);

	bfr new_net_12455_bfr_after (
		.din(new_net_12454),
		.dout(new_net_12455)
	);

	bfr new_net_12456_bfr_after (
		.din(new_net_12455),
		.dout(new_net_12456)
	);

	bfr new_net_12457_bfr_after (
		.din(new_net_12456),
		.dout(new_net_12457)
	);

	bfr new_net_12458_bfr_after (
		.din(new_net_12457),
		.dout(new_net_12458)
	);

	bfr new_net_12459_bfr_after (
		.din(new_net_12458),
		.dout(new_net_12459)
	);

	bfr new_net_12460_bfr_after (
		.din(new_net_12459),
		.dout(new_net_12460)
	);

	bfr new_net_12461_bfr_after (
		.din(new_net_12460),
		.dout(new_net_12461)
	);

	bfr new_net_12462_bfr_after (
		.din(new_net_12461),
		.dout(new_net_12462)
	);

	bfr new_net_12463_bfr_after (
		.din(new_net_12462),
		.dout(new_net_12463)
	);

	bfr new_net_12464_bfr_after (
		.din(new_net_12463),
		.dout(new_net_12464)
	);

	bfr new_net_12465_bfr_after (
		.din(new_net_12464),
		.dout(new_net_12465)
	);

	bfr new_net_12466_bfr_after (
		.din(new_net_12465),
		.dout(new_net_12466)
	);

	bfr new_net_12467_bfr_after (
		.din(new_net_12466),
		.dout(new_net_12467)
	);

	bfr new_net_12468_bfr_after (
		.din(new_net_12467),
		.dout(new_net_12468)
	);

	bfr new_net_12469_bfr_after (
		.din(new_net_12468),
		.dout(new_net_12469)
	);

	bfr new_net_12470_bfr_after (
		.din(new_net_12469),
		.dout(new_net_12470)
	);

	bfr new_net_12471_bfr_after (
		.din(new_net_12470),
		.dout(new_net_12471)
	);

	spl2 _0881__v_fanout (
		.a(new_net_12471),
		.b(new_net_2643),
		.c(new_net_2644)
	);

	bfr new_net_12472_bfr_after (
		.din(_1682_),
		.dout(new_net_12472)
	);

	bfr new_net_12473_bfr_after (
		.din(new_net_12472),
		.dout(new_net_12473)
	);

	bfr new_net_12474_bfr_after (
		.din(new_net_12473),
		.dout(new_net_12474)
	);

	bfr new_net_12475_bfr_after (
		.din(new_net_12474),
		.dout(new_net_12475)
	);

	bfr new_net_12476_bfr_after (
		.din(new_net_12475),
		.dout(new_net_12476)
	);

	bfr new_net_12477_bfr_after (
		.din(new_net_12476),
		.dout(new_net_12477)
	);

	bfr new_net_12478_bfr_after (
		.din(new_net_12477),
		.dout(new_net_12478)
	);

	bfr new_net_12479_bfr_after (
		.din(new_net_12478),
		.dout(new_net_12479)
	);

	bfr new_net_12480_bfr_after (
		.din(new_net_12479),
		.dout(new_net_12480)
	);

	bfr new_net_12481_bfr_after (
		.din(new_net_12480),
		.dout(new_net_12481)
	);

	bfr new_net_12482_bfr_after (
		.din(new_net_12481),
		.dout(new_net_12482)
	);

	bfr new_net_12483_bfr_after (
		.din(new_net_12482),
		.dout(new_net_12483)
	);

	bfr new_net_12484_bfr_after (
		.din(new_net_12483),
		.dout(new_net_12484)
	);

	bfr new_net_12485_bfr_after (
		.din(new_net_12484),
		.dout(new_net_12485)
	);

	bfr new_net_12486_bfr_after (
		.din(new_net_12485),
		.dout(new_net_12486)
	);

	bfr new_net_12487_bfr_after (
		.din(new_net_12486),
		.dout(new_net_12487)
	);

	bfr new_net_12488_bfr_after (
		.din(new_net_12487),
		.dout(new_net_12488)
	);

	bfr new_net_12489_bfr_after (
		.din(new_net_12488),
		.dout(new_net_12489)
	);

	bfr new_net_12490_bfr_after (
		.din(new_net_12489),
		.dout(new_net_12490)
	);

	bfr new_net_12491_bfr_after (
		.din(new_net_12490),
		.dout(new_net_12491)
	);

	bfr new_net_12492_bfr_after (
		.din(new_net_12491),
		.dout(new_net_12492)
	);

	bfr new_net_12493_bfr_after (
		.din(new_net_12492),
		.dout(new_net_12493)
	);

	bfr new_net_12494_bfr_after (
		.din(new_net_12493),
		.dout(new_net_12494)
	);

	bfr new_net_12495_bfr_after (
		.din(new_net_12494),
		.dout(new_net_12495)
	);

	bfr new_net_12496_bfr_after (
		.din(new_net_12495),
		.dout(new_net_12496)
	);

	bfr new_net_12497_bfr_after (
		.din(new_net_12496),
		.dout(new_net_12497)
	);

	bfr new_net_12498_bfr_after (
		.din(new_net_12497),
		.dout(new_net_12498)
	);

	bfr new_net_12499_bfr_after (
		.din(new_net_12498),
		.dout(new_net_12499)
	);

	bfr new_net_12500_bfr_after (
		.din(new_net_12499),
		.dout(new_net_12500)
	);

	bfr new_net_12501_bfr_after (
		.din(new_net_12500),
		.dout(new_net_12501)
	);

	bfr new_net_12502_bfr_after (
		.din(new_net_12501),
		.dout(new_net_12502)
	);

	bfr new_net_12503_bfr_after (
		.din(new_net_12502),
		.dout(new_net_12503)
	);

	bfr new_net_12504_bfr_after (
		.din(new_net_12503),
		.dout(new_net_12504)
	);

	bfr new_net_12505_bfr_after (
		.din(new_net_12504),
		.dout(new_net_12505)
	);

	bfr new_net_12506_bfr_after (
		.din(new_net_12505),
		.dout(new_net_12506)
	);

	bfr new_net_12507_bfr_after (
		.din(new_net_12506),
		.dout(new_net_12507)
	);

	bfr new_net_12508_bfr_after (
		.din(new_net_12507),
		.dout(new_net_12508)
	);

	bfr new_net_12509_bfr_after (
		.din(new_net_12508),
		.dout(new_net_12509)
	);

	bfr new_net_12510_bfr_after (
		.din(new_net_12509),
		.dout(new_net_12510)
	);

	bfr new_net_12511_bfr_after (
		.din(new_net_12510),
		.dout(new_net_12511)
	);

	bfr new_net_12512_bfr_after (
		.din(new_net_12511),
		.dout(new_net_12512)
	);

	bfr new_net_12513_bfr_after (
		.din(new_net_12512),
		.dout(new_net_12513)
	);

	bfr new_net_12514_bfr_after (
		.din(new_net_12513),
		.dout(new_net_12514)
	);

	bfr new_net_12515_bfr_after (
		.din(new_net_12514),
		.dout(new_net_12515)
	);

	bfr new_net_12516_bfr_after (
		.din(new_net_12515),
		.dout(new_net_12516)
	);

	bfr new_net_12517_bfr_after (
		.din(new_net_12516),
		.dout(new_net_12517)
	);

	bfr new_net_12518_bfr_after (
		.din(new_net_12517),
		.dout(new_net_12518)
	);

	bfr new_net_12519_bfr_after (
		.din(new_net_12518),
		.dout(new_net_12519)
	);

	bfr new_net_12520_bfr_after (
		.din(new_net_12519),
		.dout(new_net_12520)
	);

	bfr new_net_12521_bfr_after (
		.din(new_net_12520),
		.dout(new_net_12521)
	);

	bfr new_net_12522_bfr_after (
		.din(new_net_12521),
		.dout(new_net_12522)
	);

	bfr new_net_12523_bfr_after (
		.din(new_net_12522),
		.dout(new_net_12523)
	);

	bfr new_net_12524_bfr_after (
		.din(new_net_12523),
		.dout(new_net_12524)
	);

	bfr new_net_12525_bfr_after (
		.din(new_net_12524),
		.dout(new_net_12525)
	);

	bfr new_net_12526_bfr_after (
		.din(new_net_12525),
		.dout(new_net_12526)
	);

	bfr new_net_12527_bfr_after (
		.din(new_net_12526),
		.dout(new_net_12527)
	);

	bfr new_net_12528_bfr_after (
		.din(new_net_12527),
		.dout(new_net_12528)
	);

	bfr new_net_12529_bfr_after (
		.din(new_net_12528),
		.dout(new_net_12529)
	);

	bfr new_net_12530_bfr_after (
		.din(new_net_12529),
		.dout(new_net_12530)
	);

	bfr new_net_12531_bfr_after (
		.din(new_net_12530),
		.dout(new_net_12531)
	);

	bfr new_net_12532_bfr_after (
		.din(new_net_12531),
		.dout(new_net_12532)
	);

	bfr new_net_12533_bfr_after (
		.din(new_net_12532),
		.dout(new_net_12533)
	);

	bfr new_net_12534_bfr_after (
		.din(new_net_12533),
		.dout(new_net_12534)
	);

	bfr new_net_12535_bfr_after (
		.din(new_net_12534),
		.dout(new_net_12535)
	);

	bfr new_net_12536_bfr_after (
		.din(new_net_12535),
		.dout(new_net_12536)
	);

	bfr new_net_12537_bfr_after (
		.din(new_net_12536),
		.dout(new_net_12537)
	);

	bfr new_net_12538_bfr_after (
		.din(new_net_12537),
		.dout(new_net_12538)
	);

	bfr new_net_12539_bfr_after (
		.din(new_net_12538),
		.dout(new_net_12539)
	);

	bfr new_net_12540_bfr_after (
		.din(new_net_12539),
		.dout(new_net_12540)
	);

	bfr new_net_12541_bfr_after (
		.din(new_net_12540),
		.dout(new_net_12541)
	);

	bfr new_net_12542_bfr_after (
		.din(new_net_12541),
		.dout(new_net_12542)
	);

	bfr new_net_12543_bfr_after (
		.din(new_net_12542),
		.dout(new_net_12543)
	);

	bfr new_net_12544_bfr_after (
		.din(new_net_12543),
		.dout(new_net_12544)
	);

	bfr new_net_12545_bfr_after (
		.din(new_net_12544),
		.dout(new_net_12545)
	);

	bfr new_net_12546_bfr_after (
		.din(new_net_12545),
		.dout(new_net_12546)
	);

	bfr new_net_12547_bfr_after (
		.din(new_net_12546),
		.dout(new_net_12547)
	);

	bfr new_net_12548_bfr_after (
		.din(new_net_12547),
		.dout(new_net_12548)
	);

	bfr new_net_12549_bfr_after (
		.din(new_net_12548),
		.dout(new_net_12549)
	);

	bfr new_net_12550_bfr_after (
		.din(new_net_12549),
		.dout(new_net_12550)
	);

	bfr new_net_12551_bfr_after (
		.din(new_net_12550),
		.dout(new_net_12551)
	);

	bfr new_net_12552_bfr_after (
		.din(new_net_12551),
		.dout(new_net_12552)
	);

	bfr new_net_12553_bfr_after (
		.din(new_net_12552),
		.dout(new_net_12553)
	);

	bfr new_net_12554_bfr_after (
		.din(new_net_12553),
		.dout(new_net_12554)
	);

	bfr new_net_12555_bfr_after (
		.din(new_net_12554),
		.dout(new_net_12555)
	);

	bfr new_net_12556_bfr_after (
		.din(new_net_12555),
		.dout(new_net_12556)
	);

	bfr new_net_12557_bfr_after (
		.din(new_net_12556),
		.dout(new_net_12557)
	);

	bfr new_net_12558_bfr_after (
		.din(new_net_12557),
		.dout(new_net_12558)
	);

	bfr new_net_12559_bfr_after (
		.din(new_net_12558),
		.dout(new_net_12559)
	);

	bfr new_net_12560_bfr_after (
		.din(new_net_12559),
		.dout(new_net_12560)
	);

	bfr new_net_12561_bfr_after (
		.din(new_net_12560),
		.dout(new_net_12561)
	);

	bfr new_net_12562_bfr_after (
		.din(new_net_12561),
		.dout(new_net_12562)
	);

	bfr new_net_12563_bfr_after (
		.din(new_net_12562),
		.dout(new_net_12563)
	);

	bfr new_net_12564_bfr_after (
		.din(new_net_12563),
		.dout(new_net_12564)
	);

	bfr new_net_12565_bfr_after (
		.din(new_net_12564),
		.dout(new_net_12565)
	);

	bfr new_net_12566_bfr_after (
		.din(new_net_12565),
		.dout(new_net_12566)
	);

	bfr new_net_12567_bfr_after (
		.din(new_net_12566),
		.dout(new_net_12567)
	);

	spl2 _1682__v_fanout (
		.a(new_net_12567),
		.b(new_net_1106),
		.c(new_net_1107)
	);

	bfr new_net_12568_bfr_after (
		.din(_1807_),
		.dout(new_net_12568)
	);

	bfr new_net_12569_bfr_after (
		.din(new_net_12568),
		.dout(new_net_12569)
	);

	bfr new_net_12570_bfr_after (
		.din(new_net_12569),
		.dout(new_net_12570)
	);

	bfr new_net_12571_bfr_after (
		.din(new_net_12570),
		.dout(new_net_12571)
	);

	bfr new_net_12572_bfr_after (
		.din(new_net_12571),
		.dout(new_net_12572)
	);

	bfr new_net_12573_bfr_after (
		.din(new_net_12572),
		.dout(new_net_12573)
	);

	bfr new_net_12574_bfr_after (
		.din(new_net_12573),
		.dout(new_net_12574)
	);

	bfr new_net_12575_bfr_after (
		.din(new_net_12574),
		.dout(new_net_12575)
	);

	bfr new_net_12576_bfr_after (
		.din(new_net_12575),
		.dout(new_net_12576)
	);

	bfr new_net_12577_bfr_after (
		.din(new_net_12576),
		.dout(new_net_12577)
	);

	bfr new_net_12578_bfr_after (
		.din(new_net_12577),
		.dout(new_net_12578)
	);

	bfr new_net_12579_bfr_after (
		.din(new_net_12578),
		.dout(new_net_12579)
	);

	bfr new_net_12580_bfr_after (
		.din(new_net_12579),
		.dout(new_net_12580)
	);

	bfr new_net_12581_bfr_after (
		.din(new_net_12580),
		.dout(new_net_12581)
	);

	bfr new_net_12582_bfr_after (
		.din(new_net_12581),
		.dout(new_net_12582)
	);

	bfr new_net_12583_bfr_after (
		.din(new_net_12582),
		.dout(new_net_12583)
	);

	bfr new_net_12584_bfr_after (
		.din(new_net_12583),
		.dout(new_net_12584)
	);

	bfr new_net_12585_bfr_after (
		.din(new_net_12584),
		.dout(new_net_12585)
	);

	bfr new_net_12586_bfr_after (
		.din(new_net_12585),
		.dout(new_net_12586)
	);

	bfr new_net_12587_bfr_after (
		.din(new_net_12586),
		.dout(new_net_12587)
	);

	bfr new_net_12588_bfr_after (
		.din(new_net_12587),
		.dout(new_net_12588)
	);

	bfr new_net_12589_bfr_after (
		.din(new_net_12588),
		.dout(new_net_12589)
	);

	bfr new_net_12590_bfr_after (
		.din(new_net_12589),
		.dout(new_net_12590)
	);

	bfr new_net_12591_bfr_after (
		.din(new_net_12590),
		.dout(new_net_12591)
	);

	bfr new_net_12592_bfr_after (
		.din(new_net_12591),
		.dout(new_net_12592)
	);

	bfr new_net_12593_bfr_after (
		.din(new_net_12592),
		.dout(new_net_12593)
	);

	bfr new_net_12594_bfr_after (
		.din(new_net_12593),
		.dout(new_net_12594)
	);

	bfr new_net_12595_bfr_after (
		.din(new_net_12594),
		.dout(new_net_12595)
	);

	bfr new_net_12596_bfr_after (
		.din(new_net_12595),
		.dout(new_net_12596)
	);

	bfr new_net_12597_bfr_after (
		.din(new_net_12596),
		.dout(new_net_12597)
	);

	bfr new_net_12598_bfr_after (
		.din(new_net_12597),
		.dout(new_net_12598)
	);

	bfr new_net_12599_bfr_after (
		.din(new_net_12598),
		.dout(new_net_12599)
	);

	bfr new_net_12600_bfr_after (
		.din(new_net_12599),
		.dout(new_net_12600)
	);

	bfr new_net_12601_bfr_after (
		.din(new_net_12600),
		.dout(new_net_12601)
	);

	bfr new_net_12602_bfr_after (
		.din(new_net_12601),
		.dout(new_net_12602)
	);

	bfr new_net_12603_bfr_after (
		.din(new_net_12602),
		.dout(new_net_12603)
	);

	bfr new_net_12604_bfr_after (
		.din(new_net_12603),
		.dout(new_net_12604)
	);

	bfr new_net_12605_bfr_after (
		.din(new_net_12604),
		.dout(new_net_12605)
	);

	bfr new_net_12606_bfr_after (
		.din(new_net_12605),
		.dout(new_net_12606)
	);

	bfr new_net_12607_bfr_after (
		.din(new_net_12606),
		.dout(new_net_12607)
	);

	bfr new_net_12608_bfr_after (
		.din(new_net_12607),
		.dout(new_net_12608)
	);

	bfr new_net_12609_bfr_after (
		.din(new_net_12608),
		.dout(new_net_12609)
	);

	bfr new_net_12610_bfr_after (
		.din(new_net_12609),
		.dout(new_net_12610)
	);

	bfr new_net_12611_bfr_after (
		.din(new_net_12610),
		.dout(new_net_12611)
	);

	bfr new_net_12612_bfr_after (
		.din(new_net_12611),
		.dout(new_net_12612)
	);

	bfr new_net_12613_bfr_after (
		.din(new_net_12612),
		.dout(new_net_12613)
	);

	bfr new_net_12614_bfr_after (
		.din(new_net_12613),
		.dout(new_net_12614)
	);

	bfr new_net_12615_bfr_after (
		.din(new_net_12614),
		.dout(new_net_12615)
	);

	bfr new_net_12616_bfr_after (
		.din(new_net_12615),
		.dout(new_net_12616)
	);

	bfr new_net_12617_bfr_after (
		.din(new_net_12616),
		.dout(new_net_12617)
	);

	bfr new_net_12618_bfr_after (
		.din(new_net_12617),
		.dout(new_net_12618)
	);

	bfr new_net_12619_bfr_after (
		.din(new_net_12618),
		.dout(new_net_12619)
	);

	bfr new_net_12620_bfr_after (
		.din(new_net_12619),
		.dout(new_net_12620)
	);

	bfr new_net_12621_bfr_after (
		.din(new_net_12620),
		.dout(new_net_12621)
	);

	bfr new_net_12622_bfr_after (
		.din(new_net_12621),
		.dout(new_net_12622)
	);

	bfr new_net_12623_bfr_after (
		.din(new_net_12622),
		.dout(new_net_12623)
	);

	bfr new_net_12624_bfr_after (
		.din(new_net_12623),
		.dout(new_net_12624)
	);

	bfr new_net_12625_bfr_after (
		.din(new_net_12624),
		.dout(new_net_12625)
	);

	bfr new_net_12626_bfr_after (
		.din(new_net_12625),
		.dout(new_net_12626)
	);

	bfr new_net_12627_bfr_after (
		.din(new_net_12626),
		.dout(new_net_12627)
	);

	bfr new_net_12628_bfr_after (
		.din(new_net_12627),
		.dout(new_net_12628)
	);

	bfr new_net_12629_bfr_after (
		.din(new_net_12628),
		.dout(new_net_12629)
	);

	bfr new_net_12630_bfr_after (
		.din(new_net_12629),
		.dout(new_net_12630)
	);

	bfr new_net_12631_bfr_after (
		.din(new_net_12630),
		.dout(new_net_12631)
	);

	bfr new_net_12632_bfr_after (
		.din(new_net_12631),
		.dout(new_net_12632)
	);

	bfr new_net_12633_bfr_after (
		.din(new_net_12632),
		.dout(new_net_12633)
	);

	bfr new_net_12634_bfr_after (
		.din(new_net_12633),
		.dout(new_net_12634)
	);

	bfr new_net_12635_bfr_after (
		.din(new_net_12634),
		.dout(new_net_12635)
	);

	bfr new_net_12636_bfr_after (
		.din(new_net_12635),
		.dout(new_net_12636)
	);

	bfr new_net_12637_bfr_after (
		.din(new_net_12636),
		.dout(new_net_12637)
	);

	bfr new_net_12638_bfr_after (
		.din(new_net_12637),
		.dout(new_net_12638)
	);

	bfr new_net_12639_bfr_after (
		.din(new_net_12638),
		.dout(new_net_12639)
	);

	bfr new_net_12640_bfr_after (
		.din(new_net_12639),
		.dout(new_net_12640)
	);

	bfr new_net_12641_bfr_after (
		.din(new_net_12640),
		.dout(new_net_12641)
	);

	bfr new_net_12642_bfr_after (
		.din(new_net_12641),
		.dout(new_net_12642)
	);

	bfr new_net_12643_bfr_after (
		.din(new_net_12642),
		.dout(new_net_12643)
	);

	bfr new_net_12644_bfr_after (
		.din(new_net_12643),
		.dout(new_net_12644)
	);

	bfr new_net_12645_bfr_after (
		.din(new_net_12644),
		.dout(new_net_12645)
	);

	bfr new_net_12646_bfr_after (
		.din(new_net_12645),
		.dout(new_net_12646)
	);

	bfr new_net_12647_bfr_after (
		.din(new_net_12646),
		.dout(new_net_12647)
	);

	bfr new_net_12648_bfr_after (
		.din(new_net_12647),
		.dout(new_net_12648)
	);

	bfr new_net_12649_bfr_after (
		.din(new_net_12648),
		.dout(new_net_12649)
	);

	bfr new_net_12650_bfr_after (
		.din(new_net_12649),
		.dout(new_net_12650)
	);

	bfr new_net_12651_bfr_after (
		.din(new_net_12650),
		.dout(new_net_12651)
	);

	bfr new_net_12652_bfr_after (
		.din(new_net_12651),
		.dout(new_net_12652)
	);

	bfr new_net_12653_bfr_after (
		.din(new_net_12652),
		.dout(new_net_12653)
	);

	bfr new_net_12654_bfr_after (
		.din(new_net_12653),
		.dout(new_net_12654)
	);

	bfr new_net_12655_bfr_after (
		.din(new_net_12654),
		.dout(new_net_12655)
	);

	bfr new_net_12656_bfr_after (
		.din(new_net_12655),
		.dout(new_net_12656)
	);

	bfr new_net_12657_bfr_after (
		.din(new_net_12656),
		.dout(new_net_12657)
	);

	bfr new_net_12658_bfr_after (
		.din(new_net_12657),
		.dout(new_net_12658)
	);

	bfr new_net_12659_bfr_after (
		.din(new_net_12658),
		.dout(new_net_12659)
	);

	bfr new_net_12660_bfr_after (
		.din(new_net_12659),
		.dout(new_net_12660)
	);

	bfr new_net_12661_bfr_after (
		.din(new_net_12660),
		.dout(new_net_12661)
	);

	bfr new_net_12662_bfr_after (
		.din(new_net_12661),
		.dout(new_net_12662)
	);

	bfr new_net_12663_bfr_after (
		.din(new_net_12662),
		.dout(new_net_12663)
	);

	spl2 _1807__v_fanout (
		.a(new_net_12663),
		.b(new_net_2663),
		.c(new_net_2664)
	);

	bfr new_net_12664_bfr_after (
		.din(_0218_),
		.dout(new_net_12664)
	);

	bfr new_net_12665_bfr_after (
		.din(new_net_12664),
		.dout(new_net_12665)
	);

	bfr new_net_12666_bfr_after (
		.din(new_net_12665),
		.dout(new_net_12666)
	);

	bfr new_net_12667_bfr_after (
		.din(new_net_12666),
		.dout(new_net_12667)
	);

	bfr new_net_12668_bfr_after (
		.din(new_net_12667),
		.dout(new_net_12668)
	);

	bfr new_net_12669_bfr_after (
		.din(new_net_12668),
		.dout(new_net_12669)
	);

	bfr new_net_12670_bfr_after (
		.din(new_net_12669),
		.dout(new_net_12670)
	);

	bfr new_net_12671_bfr_after (
		.din(new_net_12670),
		.dout(new_net_12671)
	);

	bfr new_net_12672_bfr_after (
		.din(new_net_12671),
		.dout(new_net_12672)
	);

	bfr new_net_12673_bfr_after (
		.din(new_net_12672),
		.dout(new_net_12673)
	);

	bfr new_net_12674_bfr_after (
		.din(new_net_12673),
		.dout(new_net_12674)
	);

	bfr new_net_12675_bfr_after (
		.din(new_net_12674),
		.dout(new_net_12675)
	);

	bfr new_net_12676_bfr_after (
		.din(new_net_12675),
		.dout(new_net_12676)
	);

	bfr new_net_12677_bfr_after (
		.din(new_net_12676),
		.dout(new_net_12677)
	);

	bfr new_net_12678_bfr_after (
		.din(new_net_12677),
		.dout(new_net_12678)
	);

	bfr new_net_12679_bfr_after (
		.din(new_net_12678),
		.dout(new_net_12679)
	);

	bfr new_net_12680_bfr_after (
		.din(new_net_12679),
		.dout(new_net_12680)
	);

	bfr new_net_12681_bfr_after (
		.din(new_net_12680),
		.dout(new_net_12681)
	);

	bfr new_net_12682_bfr_after (
		.din(new_net_12681),
		.dout(new_net_12682)
	);

	bfr new_net_12683_bfr_after (
		.din(new_net_12682),
		.dout(new_net_12683)
	);

	bfr new_net_12684_bfr_after (
		.din(new_net_12683),
		.dout(new_net_12684)
	);

	bfr new_net_12685_bfr_after (
		.din(new_net_12684),
		.dout(new_net_12685)
	);

	bfr new_net_12686_bfr_after (
		.din(new_net_12685),
		.dout(new_net_12686)
	);

	bfr new_net_12687_bfr_after (
		.din(new_net_12686),
		.dout(new_net_12687)
	);

	bfr new_net_12688_bfr_after (
		.din(new_net_12687),
		.dout(new_net_12688)
	);

	bfr new_net_12689_bfr_after (
		.din(new_net_12688),
		.dout(new_net_12689)
	);

	bfr new_net_12690_bfr_after (
		.din(new_net_12689),
		.dout(new_net_12690)
	);

	bfr new_net_12691_bfr_after (
		.din(new_net_12690),
		.dout(new_net_12691)
	);

	bfr new_net_12692_bfr_after (
		.din(new_net_12691),
		.dout(new_net_12692)
	);

	bfr new_net_12693_bfr_after (
		.din(new_net_12692),
		.dout(new_net_12693)
	);

	bfr new_net_12694_bfr_after (
		.din(new_net_12693),
		.dout(new_net_12694)
	);

	bfr new_net_12695_bfr_after (
		.din(new_net_12694),
		.dout(new_net_12695)
	);

	bfr new_net_12696_bfr_after (
		.din(new_net_12695),
		.dout(new_net_12696)
	);

	bfr new_net_12697_bfr_after (
		.din(new_net_12696),
		.dout(new_net_12697)
	);

	bfr new_net_12698_bfr_after (
		.din(new_net_12697),
		.dout(new_net_12698)
	);

	bfr new_net_12699_bfr_after (
		.din(new_net_12698),
		.dout(new_net_12699)
	);

	bfr new_net_12700_bfr_after (
		.din(new_net_12699),
		.dout(new_net_12700)
	);

	bfr new_net_12701_bfr_after (
		.din(new_net_12700),
		.dout(new_net_12701)
	);

	bfr new_net_12702_bfr_after (
		.din(new_net_12701),
		.dout(new_net_12702)
	);

	bfr new_net_12703_bfr_after (
		.din(new_net_12702),
		.dout(new_net_12703)
	);

	bfr new_net_12704_bfr_after (
		.din(new_net_12703),
		.dout(new_net_12704)
	);

	bfr new_net_12705_bfr_after (
		.din(new_net_12704),
		.dout(new_net_12705)
	);

	bfr new_net_12706_bfr_after (
		.din(new_net_12705),
		.dout(new_net_12706)
	);

	bfr new_net_12707_bfr_after (
		.din(new_net_12706),
		.dout(new_net_12707)
	);

	bfr new_net_12708_bfr_after (
		.din(new_net_12707),
		.dout(new_net_12708)
	);

	bfr new_net_12709_bfr_after (
		.din(new_net_12708),
		.dout(new_net_12709)
	);

	bfr new_net_12710_bfr_after (
		.din(new_net_12709),
		.dout(new_net_12710)
	);

	bfr new_net_12711_bfr_after (
		.din(new_net_12710),
		.dout(new_net_12711)
	);

	bfr new_net_12712_bfr_after (
		.din(new_net_12711),
		.dout(new_net_12712)
	);

	bfr new_net_12713_bfr_after (
		.din(new_net_12712),
		.dout(new_net_12713)
	);

	bfr new_net_12714_bfr_after (
		.din(new_net_12713),
		.dout(new_net_12714)
	);

	bfr new_net_12715_bfr_after (
		.din(new_net_12714),
		.dout(new_net_12715)
	);

	bfr new_net_12716_bfr_after (
		.din(new_net_12715),
		.dout(new_net_12716)
	);

	bfr new_net_12717_bfr_after (
		.din(new_net_12716),
		.dout(new_net_12717)
	);

	bfr new_net_12718_bfr_after (
		.din(new_net_12717),
		.dout(new_net_12718)
	);

	bfr new_net_12719_bfr_after (
		.din(new_net_12718),
		.dout(new_net_12719)
	);

	bfr new_net_12720_bfr_after (
		.din(new_net_12719),
		.dout(new_net_12720)
	);

	bfr new_net_12721_bfr_after (
		.din(new_net_12720),
		.dout(new_net_12721)
	);

	bfr new_net_12722_bfr_after (
		.din(new_net_12721),
		.dout(new_net_12722)
	);

	bfr new_net_12723_bfr_after (
		.din(new_net_12722),
		.dout(new_net_12723)
	);

	bfr new_net_12724_bfr_after (
		.din(new_net_12723),
		.dout(new_net_12724)
	);

	bfr new_net_12725_bfr_after (
		.din(new_net_12724),
		.dout(new_net_12725)
	);

	bfr new_net_12726_bfr_after (
		.din(new_net_12725),
		.dout(new_net_12726)
	);

	bfr new_net_12727_bfr_after (
		.din(new_net_12726),
		.dout(new_net_12727)
	);

	bfr new_net_12728_bfr_after (
		.din(new_net_12727),
		.dout(new_net_12728)
	);

	bfr new_net_12729_bfr_after (
		.din(new_net_12728),
		.dout(new_net_12729)
	);

	bfr new_net_12730_bfr_after (
		.din(new_net_12729),
		.dout(new_net_12730)
	);

	bfr new_net_12731_bfr_after (
		.din(new_net_12730),
		.dout(new_net_12731)
	);

	bfr new_net_12732_bfr_after (
		.din(new_net_12731),
		.dout(new_net_12732)
	);

	bfr new_net_12733_bfr_after (
		.din(new_net_12732),
		.dout(new_net_12733)
	);

	bfr new_net_12734_bfr_after (
		.din(new_net_12733),
		.dout(new_net_12734)
	);

	bfr new_net_12735_bfr_after (
		.din(new_net_12734),
		.dout(new_net_12735)
	);

	bfr new_net_12736_bfr_after (
		.din(new_net_12735),
		.dout(new_net_12736)
	);

	bfr new_net_12737_bfr_after (
		.din(new_net_12736),
		.dout(new_net_12737)
	);

	bfr new_net_12738_bfr_after (
		.din(new_net_12737),
		.dout(new_net_12738)
	);

	bfr new_net_12739_bfr_after (
		.din(new_net_12738),
		.dout(new_net_12739)
	);

	bfr new_net_12740_bfr_after (
		.din(new_net_12739),
		.dout(new_net_12740)
	);

	bfr new_net_12741_bfr_after (
		.din(new_net_12740),
		.dout(new_net_12741)
	);

	bfr new_net_12742_bfr_after (
		.din(new_net_12741),
		.dout(new_net_12742)
	);

	bfr new_net_12743_bfr_after (
		.din(new_net_12742),
		.dout(new_net_12743)
	);

	bfr new_net_12744_bfr_after (
		.din(new_net_12743),
		.dout(new_net_12744)
	);

	bfr new_net_12745_bfr_after (
		.din(new_net_12744),
		.dout(new_net_12745)
	);

	bfr new_net_12746_bfr_after (
		.din(new_net_12745),
		.dout(new_net_12746)
	);

	bfr new_net_12747_bfr_after (
		.din(new_net_12746),
		.dout(new_net_12747)
	);

	bfr new_net_12748_bfr_after (
		.din(new_net_12747),
		.dout(new_net_12748)
	);

	bfr new_net_12749_bfr_after (
		.din(new_net_12748),
		.dout(new_net_12749)
	);

	bfr new_net_12750_bfr_after (
		.din(new_net_12749),
		.dout(new_net_12750)
	);

	bfr new_net_12751_bfr_after (
		.din(new_net_12750),
		.dout(new_net_12751)
	);

	spl2 _0218__v_fanout (
		.a(new_net_12751),
		.b(new_net_2740),
		.c(new_net_2741)
	);

	bfr new_net_12752_bfr_after (
		.din(_1454_),
		.dout(new_net_12752)
	);

	bfr new_net_12753_bfr_after (
		.din(new_net_12752),
		.dout(new_net_12753)
	);

	bfr new_net_12754_bfr_after (
		.din(new_net_12753),
		.dout(new_net_12754)
	);

	bfr new_net_12755_bfr_after (
		.din(new_net_12754),
		.dout(new_net_12755)
	);

	bfr new_net_12756_bfr_after (
		.din(new_net_12755),
		.dout(new_net_12756)
	);

	bfr new_net_12757_bfr_after (
		.din(new_net_12756),
		.dout(new_net_12757)
	);

	bfr new_net_12758_bfr_after (
		.din(new_net_12757),
		.dout(new_net_12758)
	);

	bfr new_net_12759_bfr_after (
		.din(new_net_12758),
		.dout(new_net_12759)
	);

	bfr new_net_12760_bfr_after (
		.din(new_net_12759),
		.dout(new_net_12760)
	);

	bfr new_net_12761_bfr_after (
		.din(new_net_12760),
		.dout(new_net_12761)
	);

	bfr new_net_12762_bfr_after (
		.din(new_net_12761),
		.dout(new_net_12762)
	);

	bfr new_net_12763_bfr_after (
		.din(new_net_12762),
		.dout(new_net_12763)
	);

	bfr new_net_12764_bfr_after (
		.din(new_net_12763),
		.dout(new_net_12764)
	);

	bfr new_net_12765_bfr_after (
		.din(new_net_12764),
		.dout(new_net_12765)
	);

	bfr new_net_12766_bfr_after (
		.din(new_net_12765),
		.dout(new_net_12766)
	);

	bfr new_net_12767_bfr_after (
		.din(new_net_12766),
		.dout(new_net_12767)
	);

	bfr new_net_12768_bfr_after (
		.din(new_net_12767),
		.dout(new_net_12768)
	);

	bfr new_net_12769_bfr_after (
		.din(new_net_12768),
		.dout(new_net_12769)
	);

	bfr new_net_12770_bfr_after (
		.din(new_net_12769),
		.dout(new_net_12770)
	);

	bfr new_net_12771_bfr_after (
		.din(new_net_12770),
		.dout(new_net_12771)
	);

	bfr new_net_12772_bfr_after (
		.din(new_net_12771),
		.dout(new_net_12772)
	);

	bfr new_net_12773_bfr_after (
		.din(new_net_12772),
		.dout(new_net_12773)
	);

	bfr new_net_12774_bfr_after (
		.din(new_net_12773),
		.dout(new_net_12774)
	);

	bfr new_net_12775_bfr_after (
		.din(new_net_12774),
		.dout(new_net_12775)
	);

	bfr new_net_12776_bfr_after (
		.din(new_net_12775),
		.dout(new_net_12776)
	);

	bfr new_net_12777_bfr_after (
		.din(new_net_12776),
		.dout(new_net_12777)
	);

	bfr new_net_12778_bfr_after (
		.din(new_net_12777),
		.dout(new_net_12778)
	);

	bfr new_net_12779_bfr_after (
		.din(new_net_12778),
		.dout(new_net_12779)
	);

	bfr new_net_12780_bfr_after (
		.din(new_net_12779),
		.dout(new_net_12780)
	);

	bfr new_net_12781_bfr_after (
		.din(new_net_12780),
		.dout(new_net_12781)
	);

	bfr new_net_12782_bfr_after (
		.din(new_net_12781),
		.dout(new_net_12782)
	);

	bfr new_net_12783_bfr_after (
		.din(new_net_12782),
		.dout(new_net_12783)
	);

	bfr new_net_12784_bfr_after (
		.din(new_net_12783),
		.dout(new_net_12784)
	);

	bfr new_net_12785_bfr_after (
		.din(new_net_12784),
		.dout(new_net_12785)
	);

	bfr new_net_12786_bfr_after (
		.din(new_net_12785),
		.dout(new_net_12786)
	);

	bfr new_net_12787_bfr_after (
		.din(new_net_12786),
		.dout(new_net_12787)
	);

	bfr new_net_12788_bfr_after (
		.din(new_net_12787),
		.dout(new_net_12788)
	);

	bfr new_net_12789_bfr_after (
		.din(new_net_12788),
		.dout(new_net_12789)
	);

	bfr new_net_12790_bfr_after (
		.din(new_net_12789),
		.dout(new_net_12790)
	);

	bfr new_net_12791_bfr_after (
		.din(new_net_12790),
		.dout(new_net_12791)
	);

	bfr new_net_12792_bfr_after (
		.din(new_net_12791),
		.dout(new_net_12792)
	);

	bfr new_net_12793_bfr_after (
		.din(new_net_12792),
		.dout(new_net_12793)
	);

	bfr new_net_12794_bfr_after (
		.din(new_net_12793),
		.dout(new_net_12794)
	);

	bfr new_net_12795_bfr_after (
		.din(new_net_12794),
		.dout(new_net_12795)
	);

	bfr new_net_12796_bfr_after (
		.din(new_net_12795),
		.dout(new_net_12796)
	);

	bfr new_net_12797_bfr_after (
		.din(new_net_12796),
		.dout(new_net_12797)
	);

	bfr new_net_12798_bfr_after (
		.din(new_net_12797),
		.dout(new_net_12798)
	);

	bfr new_net_12799_bfr_after (
		.din(new_net_12798),
		.dout(new_net_12799)
	);

	bfr new_net_12800_bfr_after (
		.din(new_net_12799),
		.dout(new_net_12800)
	);

	bfr new_net_12801_bfr_after (
		.din(new_net_12800),
		.dout(new_net_12801)
	);

	bfr new_net_12802_bfr_after (
		.din(new_net_12801),
		.dout(new_net_12802)
	);

	bfr new_net_12803_bfr_after (
		.din(new_net_12802),
		.dout(new_net_12803)
	);

	bfr new_net_12804_bfr_after (
		.din(new_net_12803),
		.dout(new_net_12804)
	);

	bfr new_net_12805_bfr_after (
		.din(new_net_12804),
		.dout(new_net_12805)
	);

	bfr new_net_12806_bfr_after (
		.din(new_net_12805),
		.dout(new_net_12806)
	);

	bfr new_net_12807_bfr_after (
		.din(new_net_12806),
		.dout(new_net_12807)
	);

	bfr new_net_12808_bfr_after (
		.din(new_net_12807),
		.dout(new_net_12808)
	);

	bfr new_net_12809_bfr_after (
		.din(new_net_12808),
		.dout(new_net_12809)
	);

	bfr new_net_12810_bfr_after (
		.din(new_net_12809),
		.dout(new_net_12810)
	);

	bfr new_net_12811_bfr_after (
		.din(new_net_12810),
		.dout(new_net_12811)
	);

	bfr new_net_12812_bfr_after (
		.din(new_net_12811),
		.dout(new_net_12812)
	);

	bfr new_net_12813_bfr_after (
		.din(new_net_12812),
		.dout(new_net_12813)
	);

	bfr new_net_12814_bfr_after (
		.din(new_net_12813),
		.dout(new_net_12814)
	);

	bfr new_net_12815_bfr_after (
		.din(new_net_12814),
		.dout(new_net_12815)
	);

	bfr new_net_12816_bfr_after (
		.din(new_net_12815),
		.dout(new_net_12816)
	);

	bfr new_net_12817_bfr_after (
		.din(new_net_12816),
		.dout(new_net_12817)
	);

	bfr new_net_12818_bfr_after (
		.din(new_net_12817),
		.dout(new_net_12818)
	);

	bfr new_net_12819_bfr_after (
		.din(new_net_12818),
		.dout(new_net_12819)
	);

	bfr new_net_12820_bfr_after (
		.din(new_net_12819),
		.dout(new_net_12820)
	);

	bfr new_net_12821_bfr_after (
		.din(new_net_12820),
		.dout(new_net_12821)
	);

	bfr new_net_12822_bfr_after (
		.din(new_net_12821),
		.dout(new_net_12822)
	);

	bfr new_net_12823_bfr_after (
		.din(new_net_12822),
		.dout(new_net_12823)
	);

	bfr new_net_12824_bfr_after (
		.din(new_net_12823),
		.dout(new_net_12824)
	);

	bfr new_net_12825_bfr_after (
		.din(new_net_12824),
		.dout(new_net_12825)
	);

	bfr new_net_12826_bfr_after (
		.din(new_net_12825),
		.dout(new_net_12826)
	);

	bfr new_net_12827_bfr_after (
		.din(new_net_12826),
		.dout(new_net_12827)
	);

	bfr new_net_12828_bfr_after (
		.din(new_net_12827),
		.dout(new_net_12828)
	);

	bfr new_net_12829_bfr_after (
		.din(new_net_12828),
		.dout(new_net_12829)
	);

	bfr new_net_12830_bfr_after (
		.din(new_net_12829),
		.dout(new_net_12830)
	);

	bfr new_net_12831_bfr_after (
		.din(new_net_12830),
		.dout(new_net_12831)
	);

	bfr new_net_12832_bfr_after (
		.din(new_net_12831),
		.dout(new_net_12832)
	);

	bfr new_net_12833_bfr_after (
		.din(new_net_12832),
		.dout(new_net_12833)
	);

	bfr new_net_12834_bfr_after (
		.din(new_net_12833),
		.dout(new_net_12834)
	);

	bfr new_net_12835_bfr_after (
		.din(new_net_12834),
		.dout(new_net_12835)
	);

	bfr new_net_12836_bfr_after (
		.din(new_net_12835),
		.dout(new_net_12836)
	);

	bfr new_net_12837_bfr_after (
		.din(new_net_12836),
		.dout(new_net_12837)
	);

	bfr new_net_12838_bfr_after (
		.din(new_net_12837),
		.dout(new_net_12838)
	);

	bfr new_net_12839_bfr_after (
		.din(new_net_12838),
		.dout(new_net_12839)
	);

	spl2 _1454__v_fanout (
		.a(new_net_12839),
		.b(new_net_1812),
		.c(new_net_1813)
	);

	bfr new_net_12840_bfr_after (
		.din(_1363_),
		.dout(new_net_12840)
	);

	bfr new_net_12841_bfr_after (
		.din(new_net_12840),
		.dout(new_net_12841)
	);

	bfr new_net_12842_bfr_after (
		.din(new_net_12841),
		.dout(new_net_12842)
	);

	bfr new_net_12843_bfr_after (
		.din(new_net_12842),
		.dout(new_net_12843)
	);

	bfr new_net_12844_bfr_after (
		.din(new_net_12843),
		.dout(new_net_12844)
	);

	bfr new_net_12845_bfr_after (
		.din(new_net_12844),
		.dout(new_net_12845)
	);

	bfr new_net_12846_bfr_after (
		.din(new_net_12845),
		.dout(new_net_12846)
	);

	bfr new_net_12847_bfr_after (
		.din(new_net_12846),
		.dout(new_net_12847)
	);

	bfr new_net_12848_bfr_after (
		.din(new_net_12847),
		.dout(new_net_12848)
	);

	bfr new_net_12849_bfr_after (
		.din(new_net_12848),
		.dout(new_net_12849)
	);

	bfr new_net_12850_bfr_after (
		.din(new_net_12849),
		.dout(new_net_12850)
	);

	bfr new_net_12851_bfr_after (
		.din(new_net_12850),
		.dout(new_net_12851)
	);

	bfr new_net_12852_bfr_after (
		.din(new_net_12851),
		.dout(new_net_12852)
	);

	bfr new_net_12853_bfr_after (
		.din(new_net_12852),
		.dout(new_net_12853)
	);

	bfr new_net_12854_bfr_after (
		.din(new_net_12853),
		.dout(new_net_12854)
	);

	bfr new_net_12855_bfr_after (
		.din(new_net_12854),
		.dout(new_net_12855)
	);

	bfr new_net_12856_bfr_after (
		.din(new_net_12855),
		.dout(new_net_12856)
	);

	bfr new_net_12857_bfr_after (
		.din(new_net_12856),
		.dout(new_net_12857)
	);

	bfr new_net_12858_bfr_after (
		.din(new_net_12857),
		.dout(new_net_12858)
	);

	bfr new_net_12859_bfr_after (
		.din(new_net_12858),
		.dout(new_net_12859)
	);

	bfr new_net_12860_bfr_after (
		.din(new_net_12859),
		.dout(new_net_12860)
	);

	bfr new_net_12861_bfr_after (
		.din(new_net_12860),
		.dout(new_net_12861)
	);

	bfr new_net_12862_bfr_after (
		.din(new_net_12861),
		.dout(new_net_12862)
	);

	bfr new_net_12863_bfr_after (
		.din(new_net_12862),
		.dout(new_net_12863)
	);

	bfr new_net_12864_bfr_after (
		.din(new_net_12863),
		.dout(new_net_12864)
	);

	bfr new_net_12865_bfr_after (
		.din(new_net_12864),
		.dout(new_net_12865)
	);

	bfr new_net_12866_bfr_after (
		.din(new_net_12865),
		.dout(new_net_12866)
	);

	bfr new_net_12867_bfr_after (
		.din(new_net_12866),
		.dout(new_net_12867)
	);

	bfr new_net_12868_bfr_after (
		.din(new_net_12867),
		.dout(new_net_12868)
	);

	bfr new_net_12869_bfr_after (
		.din(new_net_12868),
		.dout(new_net_12869)
	);

	bfr new_net_12870_bfr_after (
		.din(new_net_12869),
		.dout(new_net_12870)
	);

	bfr new_net_12871_bfr_after (
		.din(new_net_12870),
		.dout(new_net_12871)
	);

	bfr new_net_12872_bfr_after (
		.din(new_net_12871),
		.dout(new_net_12872)
	);

	bfr new_net_12873_bfr_after (
		.din(new_net_12872),
		.dout(new_net_12873)
	);

	bfr new_net_12874_bfr_after (
		.din(new_net_12873),
		.dout(new_net_12874)
	);

	bfr new_net_12875_bfr_after (
		.din(new_net_12874),
		.dout(new_net_12875)
	);

	bfr new_net_12876_bfr_after (
		.din(new_net_12875),
		.dout(new_net_12876)
	);

	bfr new_net_12877_bfr_after (
		.din(new_net_12876),
		.dout(new_net_12877)
	);

	bfr new_net_12878_bfr_after (
		.din(new_net_12877),
		.dout(new_net_12878)
	);

	bfr new_net_12879_bfr_after (
		.din(new_net_12878),
		.dout(new_net_12879)
	);

	bfr new_net_12880_bfr_after (
		.din(new_net_12879),
		.dout(new_net_12880)
	);

	bfr new_net_12881_bfr_after (
		.din(new_net_12880),
		.dout(new_net_12881)
	);

	bfr new_net_12882_bfr_after (
		.din(new_net_12881),
		.dout(new_net_12882)
	);

	bfr new_net_12883_bfr_after (
		.din(new_net_12882),
		.dout(new_net_12883)
	);

	bfr new_net_12884_bfr_after (
		.din(new_net_12883),
		.dout(new_net_12884)
	);

	bfr new_net_12885_bfr_after (
		.din(new_net_12884),
		.dout(new_net_12885)
	);

	bfr new_net_12886_bfr_after (
		.din(new_net_12885),
		.dout(new_net_12886)
	);

	bfr new_net_12887_bfr_after (
		.din(new_net_12886),
		.dout(new_net_12887)
	);

	bfr new_net_12888_bfr_after (
		.din(new_net_12887),
		.dout(new_net_12888)
	);

	bfr new_net_12889_bfr_after (
		.din(new_net_12888),
		.dout(new_net_12889)
	);

	bfr new_net_12890_bfr_after (
		.din(new_net_12889),
		.dout(new_net_12890)
	);

	bfr new_net_12891_bfr_after (
		.din(new_net_12890),
		.dout(new_net_12891)
	);

	bfr new_net_12892_bfr_after (
		.din(new_net_12891),
		.dout(new_net_12892)
	);

	bfr new_net_12893_bfr_after (
		.din(new_net_12892),
		.dout(new_net_12893)
	);

	bfr new_net_12894_bfr_after (
		.din(new_net_12893),
		.dout(new_net_12894)
	);

	bfr new_net_12895_bfr_after (
		.din(new_net_12894),
		.dout(new_net_12895)
	);

	bfr new_net_12896_bfr_after (
		.din(new_net_12895),
		.dout(new_net_12896)
	);

	bfr new_net_12897_bfr_after (
		.din(new_net_12896),
		.dout(new_net_12897)
	);

	bfr new_net_12898_bfr_after (
		.din(new_net_12897),
		.dout(new_net_12898)
	);

	bfr new_net_12899_bfr_after (
		.din(new_net_12898),
		.dout(new_net_12899)
	);

	bfr new_net_12900_bfr_after (
		.din(new_net_12899),
		.dout(new_net_12900)
	);

	bfr new_net_12901_bfr_after (
		.din(new_net_12900),
		.dout(new_net_12901)
	);

	bfr new_net_12902_bfr_after (
		.din(new_net_12901),
		.dout(new_net_12902)
	);

	bfr new_net_12903_bfr_after (
		.din(new_net_12902),
		.dout(new_net_12903)
	);

	bfr new_net_12904_bfr_after (
		.din(new_net_12903),
		.dout(new_net_12904)
	);

	bfr new_net_12905_bfr_after (
		.din(new_net_12904),
		.dout(new_net_12905)
	);

	bfr new_net_12906_bfr_after (
		.din(new_net_12905),
		.dout(new_net_12906)
	);

	bfr new_net_12907_bfr_after (
		.din(new_net_12906),
		.dout(new_net_12907)
	);

	bfr new_net_12908_bfr_after (
		.din(new_net_12907),
		.dout(new_net_12908)
	);

	bfr new_net_12909_bfr_after (
		.din(new_net_12908),
		.dout(new_net_12909)
	);

	bfr new_net_12910_bfr_after (
		.din(new_net_12909),
		.dout(new_net_12910)
	);

	bfr new_net_12911_bfr_after (
		.din(new_net_12910),
		.dout(new_net_12911)
	);

	bfr new_net_12912_bfr_after (
		.din(new_net_12911),
		.dout(new_net_12912)
	);

	bfr new_net_12913_bfr_after (
		.din(new_net_12912),
		.dout(new_net_12913)
	);

	bfr new_net_12914_bfr_after (
		.din(new_net_12913),
		.dout(new_net_12914)
	);

	bfr new_net_12915_bfr_after (
		.din(new_net_12914),
		.dout(new_net_12915)
	);

	bfr new_net_12916_bfr_after (
		.din(new_net_12915),
		.dout(new_net_12916)
	);

	bfr new_net_12917_bfr_after (
		.din(new_net_12916),
		.dout(new_net_12917)
	);

	bfr new_net_12918_bfr_after (
		.din(new_net_12917),
		.dout(new_net_12918)
	);

	bfr new_net_12919_bfr_after (
		.din(new_net_12918),
		.dout(new_net_12919)
	);

	spl2 _1363__v_fanout (
		.a(new_net_12919),
		.b(new_net_1754),
		.c(new_net_1755)
	);

	bfr new_net_12920_bfr_after (
		.din(_1280_),
		.dout(new_net_12920)
	);

	bfr new_net_12921_bfr_after (
		.din(new_net_12920),
		.dout(new_net_12921)
	);

	bfr new_net_12922_bfr_after (
		.din(new_net_12921),
		.dout(new_net_12922)
	);

	bfr new_net_12923_bfr_after (
		.din(new_net_12922),
		.dout(new_net_12923)
	);

	bfr new_net_12924_bfr_after (
		.din(new_net_12923),
		.dout(new_net_12924)
	);

	bfr new_net_12925_bfr_after (
		.din(new_net_12924),
		.dout(new_net_12925)
	);

	bfr new_net_12926_bfr_after (
		.din(new_net_12925),
		.dout(new_net_12926)
	);

	bfr new_net_12927_bfr_after (
		.din(new_net_12926),
		.dout(new_net_12927)
	);

	bfr new_net_12928_bfr_after (
		.din(new_net_12927),
		.dout(new_net_12928)
	);

	bfr new_net_12929_bfr_after (
		.din(new_net_12928),
		.dout(new_net_12929)
	);

	bfr new_net_12930_bfr_after (
		.din(new_net_12929),
		.dout(new_net_12930)
	);

	bfr new_net_12931_bfr_after (
		.din(new_net_12930),
		.dout(new_net_12931)
	);

	bfr new_net_12932_bfr_after (
		.din(new_net_12931),
		.dout(new_net_12932)
	);

	bfr new_net_12933_bfr_after (
		.din(new_net_12932),
		.dout(new_net_12933)
	);

	bfr new_net_12934_bfr_after (
		.din(new_net_12933),
		.dout(new_net_12934)
	);

	bfr new_net_12935_bfr_after (
		.din(new_net_12934),
		.dout(new_net_12935)
	);

	bfr new_net_12936_bfr_after (
		.din(new_net_12935),
		.dout(new_net_12936)
	);

	bfr new_net_12937_bfr_after (
		.din(new_net_12936),
		.dout(new_net_12937)
	);

	bfr new_net_12938_bfr_after (
		.din(new_net_12937),
		.dout(new_net_12938)
	);

	bfr new_net_12939_bfr_after (
		.din(new_net_12938),
		.dout(new_net_12939)
	);

	bfr new_net_12940_bfr_after (
		.din(new_net_12939),
		.dout(new_net_12940)
	);

	bfr new_net_12941_bfr_after (
		.din(new_net_12940),
		.dout(new_net_12941)
	);

	bfr new_net_12942_bfr_after (
		.din(new_net_12941),
		.dout(new_net_12942)
	);

	bfr new_net_12943_bfr_after (
		.din(new_net_12942),
		.dout(new_net_12943)
	);

	bfr new_net_12944_bfr_after (
		.din(new_net_12943),
		.dout(new_net_12944)
	);

	bfr new_net_12945_bfr_after (
		.din(new_net_12944),
		.dout(new_net_12945)
	);

	bfr new_net_12946_bfr_after (
		.din(new_net_12945),
		.dout(new_net_12946)
	);

	bfr new_net_12947_bfr_after (
		.din(new_net_12946),
		.dout(new_net_12947)
	);

	bfr new_net_12948_bfr_after (
		.din(new_net_12947),
		.dout(new_net_12948)
	);

	bfr new_net_12949_bfr_after (
		.din(new_net_12948),
		.dout(new_net_12949)
	);

	bfr new_net_12950_bfr_after (
		.din(new_net_12949),
		.dout(new_net_12950)
	);

	bfr new_net_12951_bfr_after (
		.din(new_net_12950),
		.dout(new_net_12951)
	);

	bfr new_net_12952_bfr_after (
		.din(new_net_12951),
		.dout(new_net_12952)
	);

	bfr new_net_12953_bfr_after (
		.din(new_net_12952),
		.dout(new_net_12953)
	);

	bfr new_net_12954_bfr_after (
		.din(new_net_12953),
		.dout(new_net_12954)
	);

	bfr new_net_12955_bfr_after (
		.din(new_net_12954),
		.dout(new_net_12955)
	);

	bfr new_net_12956_bfr_after (
		.din(new_net_12955),
		.dout(new_net_12956)
	);

	bfr new_net_12957_bfr_after (
		.din(new_net_12956),
		.dout(new_net_12957)
	);

	bfr new_net_12958_bfr_after (
		.din(new_net_12957),
		.dout(new_net_12958)
	);

	bfr new_net_12959_bfr_after (
		.din(new_net_12958),
		.dout(new_net_12959)
	);

	bfr new_net_12960_bfr_after (
		.din(new_net_12959),
		.dout(new_net_12960)
	);

	bfr new_net_12961_bfr_after (
		.din(new_net_12960),
		.dout(new_net_12961)
	);

	bfr new_net_12962_bfr_after (
		.din(new_net_12961),
		.dout(new_net_12962)
	);

	bfr new_net_12963_bfr_after (
		.din(new_net_12962),
		.dout(new_net_12963)
	);

	bfr new_net_12964_bfr_after (
		.din(new_net_12963),
		.dout(new_net_12964)
	);

	bfr new_net_12965_bfr_after (
		.din(new_net_12964),
		.dout(new_net_12965)
	);

	bfr new_net_12966_bfr_after (
		.din(new_net_12965),
		.dout(new_net_12966)
	);

	bfr new_net_12967_bfr_after (
		.din(new_net_12966),
		.dout(new_net_12967)
	);

	bfr new_net_12968_bfr_after (
		.din(new_net_12967),
		.dout(new_net_12968)
	);

	bfr new_net_12969_bfr_after (
		.din(new_net_12968),
		.dout(new_net_12969)
	);

	bfr new_net_12970_bfr_after (
		.din(new_net_12969),
		.dout(new_net_12970)
	);

	bfr new_net_12971_bfr_after (
		.din(new_net_12970),
		.dout(new_net_12971)
	);

	bfr new_net_12972_bfr_after (
		.din(new_net_12971),
		.dout(new_net_12972)
	);

	bfr new_net_12973_bfr_after (
		.din(new_net_12972),
		.dout(new_net_12973)
	);

	bfr new_net_12974_bfr_after (
		.din(new_net_12973),
		.dout(new_net_12974)
	);

	bfr new_net_12975_bfr_after (
		.din(new_net_12974),
		.dout(new_net_12975)
	);

	bfr new_net_12976_bfr_after (
		.din(new_net_12975),
		.dout(new_net_12976)
	);

	bfr new_net_12977_bfr_after (
		.din(new_net_12976),
		.dout(new_net_12977)
	);

	bfr new_net_12978_bfr_after (
		.din(new_net_12977),
		.dout(new_net_12978)
	);

	bfr new_net_12979_bfr_after (
		.din(new_net_12978),
		.dout(new_net_12979)
	);

	bfr new_net_12980_bfr_after (
		.din(new_net_12979),
		.dout(new_net_12980)
	);

	bfr new_net_12981_bfr_after (
		.din(new_net_12980),
		.dout(new_net_12981)
	);

	bfr new_net_12982_bfr_after (
		.din(new_net_12981),
		.dout(new_net_12982)
	);

	bfr new_net_12983_bfr_after (
		.din(new_net_12982),
		.dout(new_net_12983)
	);

	bfr new_net_12984_bfr_after (
		.din(new_net_12983),
		.dout(new_net_12984)
	);

	bfr new_net_12985_bfr_after (
		.din(new_net_12984),
		.dout(new_net_12985)
	);

	bfr new_net_12986_bfr_after (
		.din(new_net_12985),
		.dout(new_net_12986)
	);

	bfr new_net_12987_bfr_after (
		.din(new_net_12986),
		.dout(new_net_12987)
	);

	bfr new_net_12988_bfr_after (
		.din(new_net_12987),
		.dout(new_net_12988)
	);

	bfr new_net_12989_bfr_after (
		.din(new_net_12988),
		.dout(new_net_12989)
	);

	bfr new_net_12990_bfr_after (
		.din(new_net_12989),
		.dout(new_net_12990)
	);

	bfr new_net_12991_bfr_after (
		.din(new_net_12990),
		.dout(new_net_12991)
	);

	spl2 _1280__v_fanout (
		.a(new_net_12991),
		.b(new_net_238),
		.c(new_net_239)
	);

	bfr new_net_12992_bfr_after (
		.din(_0445_),
		.dout(new_net_12992)
	);

	bfr new_net_12993_bfr_after (
		.din(new_net_12992),
		.dout(new_net_12993)
	);

	bfr new_net_12994_bfr_after (
		.din(new_net_12993),
		.dout(new_net_12994)
	);

	bfr new_net_12995_bfr_after (
		.din(new_net_12994),
		.dout(new_net_12995)
	);

	bfr new_net_12996_bfr_after (
		.din(new_net_12995),
		.dout(new_net_12996)
	);

	bfr new_net_12997_bfr_after (
		.din(new_net_12996),
		.dout(new_net_12997)
	);

	bfr new_net_12998_bfr_after (
		.din(new_net_12997),
		.dout(new_net_12998)
	);

	bfr new_net_12999_bfr_after (
		.din(new_net_12998),
		.dout(new_net_12999)
	);

	bfr new_net_13000_bfr_after (
		.din(new_net_12999),
		.dout(new_net_13000)
	);

	bfr new_net_13001_bfr_after (
		.din(new_net_13000),
		.dout(new_net_13001)
	);

	bfr new_net_13002_bfr_after (
		.din(new_net_13001),
		.dout(new_net_13002)
	);

	bfr new_net_13003_bfr_after (
		.din(new_net_13002),
		.dout(new_net_13003)
	);

	bfr new_net_13004_bfr_after (
		.din(new_net_13003),
		.dout(new_net_13004)
	);

	bfr new_net_13005_bfr_after (
		.din(new_net_13004),
		.dout(new_net_13005)
	);

	bfr new_net_13006_bfr_after (
		.din(new_net_13005),
		.dout(new_net_13006)
	);

	bfr new_net_13007_bfr_after (
		.din(new_net_13006),
		.dout(new_net_13007)
	);

	bfr new_net_13008_bfr_after (
		.din(new_net_13007),
		.dout(new_net_13008)
	);

	bfr new_net_13009_bfr_after (
		.din(new_net_13008),
		.dout(new_net_13009)
	);

	bfr new_net_13010_bfr_after (
		.din(new_net_13009),
		.dout(new_net_13010)
	);

	bfr new_net_13011_bfr_after (
		.din(new_net_13010),
		.dout(new_net_13011)
	);

	bfr new_net_13012_bfr_after (
		.din(new_net_13011),
		.dout(new_net_13012)
	);

	bfr new_net_13013_bfr_after (
		.din(new_net_13012),
		.dout(new_net_13013)
	);

	bfr new_net_13014_bfr_after (
		.din(new_net_13013),
		.dout(new_net_13014)
	);

	bfr new_net_13015_bfr_after (
		.din(new_net_13014),
		.dout(new_net_13015)
	);

	bfr new_net_13016_bfr_after (
		.din(new_net_13015),
		.dout(new_net_13016)
	);

	bfr new_net_13017_bfr_after (
		.din(new_net_13016),
		.dout(new_net_13017)
	);

	bfr new_net_13018_bfr_after (
		.din(new_net_13017),
		.dout(new_net_13018)
	);

	bfr new_net_13019_bfr_after (
		.din(new_net_13018),
		.dout(new_net_13019)
	);

	bfr new_net_13020_bfr_after (
		.din(new_net_13019),
		.dout(new_net_13020)
	);

	bfr new_net_13021_bfr_after (
		.din(new_net_13020),
		.dout(new_net_13021)
	);

	bfr new_net_13022_bfr_after (
		.din(new_net_13021),
		.dout(new_net_13022)
	);

	bfr new_net_13023_bfr_after (
		.din(new_net_13022),
		.dout(new_net_13023)
	);

	bfr new_net_13024_bfr_after (
		.din(new_net_13023),
		.dout(new_net_13024)
	);

	bfr new_net_13025_bfr_after (
		.din(new_net_13024),
		.dout(new_net_13025)
	);

	bfr new_net_13026_bfr_after (
		.din(new_net_13025),
		.dout(new_net_13026)
	);

	bfr new_net_13027_bfr_after (
		.din(new_net_13026),
		.dout(new_net_13027)
	);

	bfr new_net_13028_bfr_after (
		.din(new_net_13027),
		.dout(new_net_13028)
	);

	bfr new_net_13029_bfr_after (
		.din(new_net_13028),
		.dout(new_net_13029)
	);

	bfr new_net_13030_bfr_after (
		.din(new_net_13029),
		.dout(new_net_13030)
	);

	bfr new_net_13031_bfr_after (
		.din(new_net_13030),
		.dout(new_net_13031)
	);

	bfr new_net_13032_bfr_after (
		.din(new_net_13031),
		.dout(new_net_13032)
	);

	bfr new_net_13033_bfr_after (
		.din(new_net_13032),
		.dout(new_net_13033)
	);

	bfr new_net_13034_bfr_after (
		.din(new_net_13033),
		.dout(new_net_13034)
	);

	bfr new_net_13035_bfr_after (
		.din(new_net_13034),
		.dout(new_net_13035)
	);

	bfr new_net_13036_bfr_after (
		.din(new_net_13035),
		.dout(new_net_13036)
	);

	bfr new_net_13037_bfr_after (
		.din(new_net_13036),
		.dout(new_net_13037)
	);

	bfr new_net_13038_bfr_after (
		.din(new_net_13037),
		.dout(new_net_13038)
	);

	bfr new_net_13039_bfr_after (
		.din(new_net_13038),
		.dout(new_net_13039)
	);

	bfr new_net_13040_bfr_after (
		.din(new_net_13039),
		.dout(new_net_13040)
	);

	bfr new_net_13041_bfr_after (
		.din(new_net_13040),
		.dout(new_net_13041)
	);

	bfr new_net_13042_bfr_after (
		.din(new_net_13041),
		.dout(new_net_13042)
	);

	bfr new_net_13043_bfr_after (
		.din(new_net_13042),
		.dout(new_net_13043)
	);

	bfr new_net_13044_bfr_after (
		.din(new_net_13043),
		.dout(new_net_13044)
	);

	bfr new_net_13045_bfr_after (
		.din(new_net_13044),
		.dout(new_net_13045)
	);

	bfr new_net_13046_bfr_after (
		.din(new_net_13045),
		.dout(new_net_13046)
	);

	bfr new_net_13047_bfr_after (
		.din(new_net_13046),
		.dout(new_net_13047)
	);

	bfr new_net_13048_bfr_after (
		.din(new_net_13047),
		.dout(new_net_13048)
	);

	bfr new_net_13049_bfr_after (
		.din(new_net_13048),
		.dout(new_net_13049)
	);

	bfr new_net_13050_bfr_after (
		.din(new_net_13049),
		.dout(new_net_13050)
	);

	bfr new_net_13051_bfr_after (
		.din(new_net_13050),
		.dout(new_net_13051)
	);

	bfr new_net_13052_bfr_after (
		.din(new_net_13051),
		.dout(new_net_13052)
	);

	bfr new_net_13053_bfr_after (
		.din(new_net_13052),
		.dout(new_net_13053)
	);

	bfr new_net_13054_bfr_after (
		.din(new_net_13053),
		.dout(new_net_13054)
	);

	bfr new_net_13055_bfr_after (
		.din(new_net_13054),
		.dout(new_net_13055)
	);

	spl2 _0445__v_fanout (
		.a(new_net_13055),
		.b(new_net_2026),
		.c(new_net_2027)
	);

	spl2 _1480__v_fanout (
		.a(_1480_),
		.b(new_net_1425),
		.c(new_net_1426)
	);

	bfr new_net_13056_bfr_after (
		.din(_0108_),
		.dout(new_net_13056)
	);

	bfr new_net_13057_bfr_after (
		.din(new_net_13056),
		.dout(new_net_13057)
	);

	bfr new_net_13058_bfr_after (
		.din(new_net_13057),
		.dout(new_net_13058)
	);

	bfr new_net_13059_bfr_after (
		.din(new_net_13058),
		.dout(new_net_13059)
	);

	bfr new_net_13060_bfr_after (
		.din(new_net_13059),
		.dout(new_net_13060)
	);

	bfr new_net_13061_bfr_after (
		.din(new_net_13060),
		.dout(new_net_13061)
	);

	bfr new_net_13062_bfr_after (
		.din(new_net_13061),
		.dout(new_net_13062)
	);

	bfr new_net_13063_bfr_after (
		.din(new_net_13062),
		.dout(new_net_13063)
	);

	bfr new_net_13064_bfr_after (
		.din(new_net_13063),
		.dout(new_net_13064)
	);

	bfr new_net_13065_bfr_after (
		.din(new_net_13064),
		.dout(new_net_13065)
	);

	bfr new_net_13066_bfr_after (
		.din(new_net_13065),
		.dout(new_net_13066)
	);

	bfr new_net_13067_bfr_after (
		.din(new_net_13066),
		.dout(new_net_13067)
	);

	bfr new_net_13068_bfr_after (
		.din(new_net_13067),
		.dout(new_net_13068)
	);

	bfr new_net_13069_bfr_after (
		.din(new_net_13068),
		.dout(new_net_13069)
	);

	bfr new_net_13070_bfr_after (
		.din(new_net_13069),
		.dout(new_net_13070)
	);

	bfr new_net_13071_bfr_after (
		.din(new_net_13070),
		.dout(new_net_13071)
	);

	bfr new_net_13072_bfr_after (
		.din(new_net_13071),
		.dout(new_net_13072)
	);

	bfr new_net_13073_bfr_after (
		.din(new_net_13072),
		.dout(new_net_13073)
	);

	bfr new_net_13074_bfr_after (
		.din(new_net_13073),
		.dout(new_net_13074)
	);

	bfr new_net_13075_bfr_after (
		.din(new_net_13074),
		.dout(new_net_13075)
	);

	bfr new_net_13076_bfr_after (
		.din(new_net_13075),
		.dout(new_net_13076)
	);

	bfr new_net_13077_bfr_after (
		.din(new_net_13076),
		.dout(new_net_13077)
	);

	spl2 _0108__v_fanout (
		.a(new_net_13077),
		.b(new_net_2208),
		.c(new_net_2209)
	);

	bfr new_net_13078_bfr_after (
		.din(_1203_),
		.dout(new_net_13078)
	);

	bfr new_net_13079_bfr_after (
		.din(new_net_13078),
		.dout(new_net_13079)
	);

	bfr new_net_13080_bfr_after (
		.din(new_net_13079),
		.dout(new_net_13080)
	);

	bfr new_net_13081_bfr_after (
		.din(new_net_13080),
		.dout(new_net_13081)
	);

	bfr new_net_13082_bfr_after (
		.din(new_net_13081),
		.dout(new_net_13082)
	);

	bfr new_net_13083_bfr_after (
		.din(new_net_13082),
		.dout(new_net_13083)
	);

	bfr new_net_13084_bfr_after (
		.din(new_net_13083),
		.dout(new_net_13084)
	);

	bfr new_net_13085_bfr_after (
		.din(new_net_13084),
		.dout(new_net_13085)
	);

	bfr new_net_13086_bfr_after (
		.din(new_net_13085),
		.dout(new_net_13086)
	);

	bfr new_net_13087_bfr_after (
		.din(new_net_13086),
		.dout(new_net_13087)
	);

	bfr new_net_13088_bfr_after (
		.din(new_net_13087),
		.dout(new_net_13088)
	);

	bfr new_net_13089_bfr_after (
		.din(new_net_13088),
		.dout(new_net_13089)
	);

	bfr new_net_13090_bfr_after (
		.din(new_net_13089),
		.dout(new_net_13090)
	);

	bfr new_net_13091_bfr_after (
		.din(new_net_13090),
		.dout(new_net_13091)
	);

	bfr new_net_13092_bfr_after (
		.din(new_net_13091),
		.dout(new_net_13092)
	);

	bfr new_net_13093_bfr_after (
		.din(new_net_13092),
		.dout(new_net_13093)
	);

	bfr new_net_13094_bfr_after (
		.din(new_net_13093),
		.dout(new_net_13094)
	);

	bfr new_net_13095_bfr_after (
		.din(new_net_13094),
		.dout(new_net_13095)
	);

	bfr new_net_13096_bfr_after (
		.din(new_net_13095),
		.dout(new_net_13096)
	);

	bfr new_net_13097_bfr_after (
		.din(new_net_13096),
		.dout(new_net_13097)
	);

	bfr new_net_13098_bfr_after (
		.din(new_net_13097),
		.dout(new_net_13098)
	);

	bfr new_net_13099_bfr_after (
		.din(new_net_13098),
		.dout(new_net_13099)
	);

	bfr new_net_13100_bfr_after (
		.din(new_net_13099),
		.dout(new_net_13100)
	);

	bfr new_net_13101_bfr_after (
		.din(new_net_13100),
		.dout(new_net_13101)
	);

	bfr new_net_13102_bfr_after (
		.din(new_net_13101),
		.dout(new_net_13102)
	);

	bfr new_net_13103_bfr_after (
		.din(new_net_13102),
		.dout(new_net_13103)
	);

	bfr new_net_13104_bfr_after (
		.din(new_net_13103),
		.dout(new_net_13104)
	);

	bfr new_net_13105_bfr_after (
		.din(new_net_13104),
		.dout(new_net_13105)
	);

	bfr new_net_13106_bfr_after (
		.din(new_net_13105),
		.dout(new_net_13106)
	);

	bfr new_net_13107_bfr_after (
		.din(new_net_13106),
		.dout(new_net_13107)
	);

	bfr new_net_13108_bfr_after (
		.din(new_net_13107),
		.dout(new_net_13108)
	);

	bfr new_net_13109_bfr_after (
		.din(new_net_13108),
		.dout(new_net_13109)
	);

	bfr new_net_13110_bfr_after (
		.din(new_net_13109),
		.dout(new_net_13110)
	);

	bfr new_net_13111_bfr_after (
		.din(new_net_13110),
		.dout(new_net_13111)
	);

	bfr new_net_13112_bfr_after (
		.din(new_net_13111),
		.dout(new_net_13112)
	);

	bfr new_net_13113_bfr_after (
		.din(new_net_13112),
		.dout(new_net_13113)
	);

	bfr new_net_13114_bfr_after (
		.din(new_net_13113),
		.dout(new_net_13114)
	);

	bfr new_net_13115_bfr_after (
		.din(new_net_13114),
		.dout(new_net_13115)
	);

	bfr new_net_13116_bfr_after (
		.din(new_net_13115),
		.dout(new_net_13116)
	);

	bfr new_net_13117_bfr_after (
		.din(new_net_13116),
		.dout(new_net_13117)
	);

	bfr new_net_13118_bfr_after (
		.din(new_net_13117),
		.dout(new_net_13118)
	);

	bfr new_net_13119_bfr_after (
		.din(new_net_13118),
		.dout(new_net_13119)
	);

	bfr new_net_13120_bfr_after (
		.din(new_net_13119),
		.dout(new_net_13120)
	);

	bfr new_net_13121_bfr_after (
		.din(new_net_13120),
		.dout(new_net_13121)
	);

	bfr new_net_13122_bfr_after (
		.din(new_net_13121),
		.dout(new_net_13122)
	);

	bfr new_net_13123_bfr_after (
		.din(new_net_13122),
		.dout(new_net_13123)
	);

	bfr new_net_13124_bfr_after (
		.din(new_net_13123),
		.dout(new_net_13124)
	);

	bfr new_net_13125_bfr_after (
		.din(new_net_13124),
		.dout(new_net_13125)
	);

	bfr new_net_13126_bfr_after (
		.din(new_net_13125),
		.dout(new_net_13126)
	);

	bfr new_net_13127_bfr_after (
		.din(new_net_13126),
		.dout(new_net_13127)
	);

	bfr new_net_13128_bfr_after (
		.din(new_net_13127),
		.dout(new_net_13128)
	);

	bfr new_net_13129_bfr_after (
		.din(new_net_13128),
		.dout(new_net_13129)
	);

	bfr new_net_13130_bfr_after (
		.din(new_net_13129),
		.dout(new_net_13130)
	);

	bfr new_net_13131_bfr_after (
		.din(new_net_13130),
		.dout(new_net_13131)
	);

	bfr new_net_13132_bfr_after (
		.din(new_net_13131),
		.dout(new_net_13132)
	);

	bfr new_net_13133_bfr_after (
		.din(new_net_13132),
		.dout(new_net_13133)
	);

	bfr new_net_13134_bfr_after (
		.din(new_net_13133),
		.dout(new_net_13134)
	);

	bfr new_net_13135_bfr_after (
		.din(new_net_13134),
		.dout(new_net_13135)
	);

	bfr new_net_13136_bfr_after (
		.din(new_net_13135),
		.dout(new_net_13136)
	);

	bfr new_net_13137_bfr_after (
		.din(new_net_13136),
		.dout(new_net_13137)
	);

	bfr new_net_13138_bfr_after (
		.din(new_net_13137),
		.dout(new_net_13138)
	);

	bfr new_net_13139_bfr_after (
		.din(new_net_13138),
		.dout(new_net_13139)
	);

	bfr new_net_13140_bfr_after (
		.din(new_net_13139),
		.dout(new_net_13140)
	);

	bfr new_net_13141_bfr_after (
		.din(new_net_13140),
		.dout(new_net_13141)
	);

	bfr new_net_13142_bfr_after (
		.din(new_net_13141),
		.dout(new_net_13142)
	);

	bfr new_net_13143_bfr_after (
		.din(new_net_13142),
		.dout(new_net_13143)
	);

	bfr new_net_13144_bfr_after (
		.din(new_net_13143),
		.dout(new_net_13144)
	);

	bfr new_net_13145_bfr_after (
		.din(new_net_13144),
		.dout(new_net_13145)
	);

	bfr new_net_13146_bfr_after (
		.din(new_net_13145),
		.dout(new_net_13146)
	);

	bfr new_net_13147_bfr_after (
		.din(new_net_13146),
		.dout(new_net_13147)
	);

	bfr new_net_13148_bfr_after (
		.din(new_net_13147),
		.dout(new_net_13148)
	);

	bfr new_net_13149_bfr_after (
		.din(new_net_13148),
		.dout(new_net_13149)
	);

	spl2 _1203__v_fanout (
		.a(new_net_13149),
		.b(new_net_2981),
		.c(new_net_2982)
	);

	bfr new_net_13150_bfr_after (
		.din(_0434_),
		.dout(new_net_13150)
	);

	bfr new_net_13151_bfr_after (
		.din(new_net_13150),
		.dout(new_net_13151)
	);

	bfr new_net_13152_bfr_after (
		.din(new_net_13151),
		.dout(new_net_13152)
	);

	bfr new_net_13153_bfr_after (
		.din(new_net_13152),
		.dout(new_net_13153)
	);

	bfr new_net_13154_bfr_after (
		.din(new_net_13153),
		.dout(new_net_13154)
	);

	bfr new_net_13155_bfr_after (
		.din(new_net_13154),
		.dout(new_net_13155)
	);

	bfr new_net_13156_bfr_after (
		.din(new_net_13155),
		.dout(new_net_13156)
	);

	bfr new_net_13157_bfr_after (
		.din(new_net_13156),
		.dout(new_net_13157)
	);

	bfr new_net_13158_bfr_after (
		.din(new_net_13157),
		.dout(new_net_13158)
	);

	bfr new_net_13159_bfr_after (
		.din(new_net_13158),
		.dout(new_net_13159)
	);

	bfr new_net_13160_bfr_after (
		.din(new_net_13159),
		.dout(new_net_13160)
	);

	bfr new_net_13161_bfr_after (
		.din(new_net_13160),
		.dout(new_net_13161)
	);

	bfr new_net_13162_bfr_after (
		.din(new_net_13161),
		.dout(new_net_13162)
	);

	bfr new_net_13163_bfr_after (
		.din(new_net_13162),
		.dout(new_net_13163)
	);

	bfr new_net_13164_bfr_after (
		.din(new_net_13163),
		.dout(new_net_13164)
	);

	bfr new_net_13165_bfr_after (
		.din(new_net_13164),
		.dout(new_net_13165)
	);

	bfr new_net_13166_bfr_after (
		.din(new_net_13165),
		.dout(new_net_13166)
	);

	bfr new_net_13167_bfr_after (
		.din(new_net_13166),
		.dout(new_net_13167)
	);

	bfr new_net_13168_bfr_after (
		.din(new_net_13167),
		.dout(new_net_13168)
	);

	bfr new_net_13169_bfr_after (
		.din(new_net_13168),
		.dout(new_net_13169)
	);

	bfr new_net_13170_bfr_after (
		.din(new_net_13169),
		.dout(new_net_13170)
	);

	bfr new_net_13171_bfr_after (
		.din(new_net_13170),
		.dout(new_net_13171)
	);

	bfr new_net_13172_bfr_after (
		.din(new_net_13171),
		.dout(new_net_13172)
	);

	bfr new_net_13173_bfr_after (
		.din(new_net_13172),
		.dout(new_net_13173)
	);

	bfr new_net_13174_bfr_after (
		.din(new_net_13173),
		.dout(new_net_13174)
	);

	bfr new_net_13175_bfr_after (
		.din(new_net_13174),
		.dout(new_net_13175)
	);

	bfr new_net_13176_bfr_after (
		.din(new_net_13175),
		.dout(new_net_13176)
	);

	bfr new_net_13177_bfr_after (
		.din(new_net_13176),
		.dout(new_net_13177)
	);

	bfr new_net_13178_bfr_after (
		.din(new_net_13177),
		.dout(new_net_13178)
	);

	bfr new_net_13179_bfr_after (
		.din(new_net_13178),
		.dout(new_net_13179)
	);

	bfr new_net_13180_bfr_after (
		.din(new_net_13179),
		.dout(new_net_13180)
	);

	bfr new_net_13181_bfr_after (
		.din(new_net_13180),
		.dout(new_net_13181)
	);

	bfr new_net_13182_bfr_after (
		.din(new_net_13181),
		.dout(new_net_13182)
	);

	bfr new_net_13183_bfr_after (
		.din(new_net_13182),
		.dout(new_net_13183)
	);

	bfr new_net_13184_bfr_after (
		.din(new_net_13183),
		.dout(new_net_13184)
	);

	bfr new_net_13185_bfr_after (
		.din(new_net_13184),
		.dout(new_net_13185)
	);

	bfr new_net_13186_bfr_after (
		.din(new_net_13185),
		.dout(new_net_13186)
	);

	bfr new_net_13187_bfr_after (
		.din(new_net_13186),
		.dout(new_net_13187)
	);

	bfr new_net_13188_bfr_after (
		.din(new_net_13187),
		.dout(new_net_13188)
	);

	bfr new_net_13189_bfr_after (
		.din(new_net_13188),
		.dout(new_net_13189)
	);

	bfr new_net_13190_bfr_after (
		.din(new_net_13189),
		.dout(new_net_13190)
	);

	bfr new_net_13191_bfr_after (
		.din(new_net_13190),
		.dout(new_net_13191)
	);

	bfr new_net_13192_bfr_after (
		.din(new_net_13191),
		.dout(new_net_13192)
	);

	bfr new_net_13193_bfr_after (
		.din(new_net_13192),
		.dout(new_net_13193)
	);

	bfr new_net_13194_bfr_after (
		.din(new_net_13193),
		.dout(new_net_13194)
	);

	bfr new_net_13195_bfr_after (
		.din(new_net_13194),
		.dout(new_net_13195)
	);

	bfr new_net_13196_bfr_after (
		.din(new_net_13195),
		.dout(new_net_13196)
	);

	bfr new_net_13197_bfr_after (
		.din(new_net_13196),
		.dout(new_net_13197)
	);

	bfr new_net_13198_bfr_after (
		.din(new_net_13197),
		.dout(new_net_13198)
	);

	bfr new_net_13199_bfr_after (
		.din(new_net_13198),
		.dout(new_net_13199)
	);

	bfr new_net_13200_bfr_after (
		.din(new_net_13199),
		.dout(new_net_13200)
	);

	bfr new_net_13201_bfr_after (
		.din(new_net_13200),
		.dout(new_net_13201)
	);

	bfr new_net_13202_bfr_after (
		.din(new_net_13201),
		.dout(new_net_13202)
	);

	bfr new_net_13203_bfr_after (
		.din(new_net_13202),
		.dout(new_net_13203)
	);

	bfr new_net_13204_bfr_after (
		.din(new_net_13203),
		.dout(new_net_13204)
	);

	bfr new_net_13205_bfr_after (
		.din(new_net_13204),
		.dout(new_net_13205)
	);

	bfr new_net_13206_bfr_after (
		.din(new_net_13205),
		.dout(new_net_13206)
	);

	bfr new_net_13207_bfr_after (
		.din(new_net_13206),
		.dout(new_net_13207)
	);

	bfr new_net_13208_bfr_after (
		.din(new_net_13207),
		.dout(new_net_13208)
	);

	bfr new_net_13209_bfr_after (
		.din(new_net_13208),
		.dout(new_net_13209)
	);

	bfr new_net_13210_bfr_after (
		.din(new_net_13209),
		.dout(new_net_13210)
	);

	bfr new_net_13211_bfr_after (
		.din(new_net_13210),
		.dout(new_net_13211)
	);

	bfr new_net_13212_bfr_after (
		.din(new_net_13211),
		.dout(new_net_13212)
	);

	bfr new_net_13213_bfr_after (
		.din(new_net_13212),
		.dout(new_net_13213)
	);

	bfr new_net_13214_bfr_after (
		.din(new_net_13213),
		.dout(new_net_13214)
	);

	bfr new_net_13215_bfr_after (
		.din(new_net_13214),
		.dout(new_net_13215)
	);

	bfr new_net_13216_bfr_after (
		.din(new_net_13215),
		.dout(new_net_13216)
	);

	bfr new_net_13217_bfr_after (
		.din(new_net_13216),
		.dout(new_net_13217)
	);

	bfr new_net_13218_bfr_after (
		.din(new_net_13217),
		.dout(new_net_13218)
	);

	bfr new_net_13219_bfr_after (
		.din(new_net_13218),
		.dout(new_net_13219)
	);

	bfr new_net_13220_bfr_after (
		.din(new_net_13219),
		.dout(new_net_13220)
	);

	bfr new_net_13221_bfr_after (
		.din(new_net_13220),
		.dout(new_net_13221)
	);

	bfr new_net_13222_bfr_after (
		.din(new_net_13221),
		.dout(new_net_13222)
	);

	bfr new_net_13223_bfr_after (
		.din(new_net_13222),
		.dout(new_net_13223)
	);

	bfr new_net_13224_bfr_after (
		.din(new_net_13223),
		.dout(new_net_13224)
	);

	bfr new_net_13225_bfr_after (
		.din(new_net_13224),
		.dout(new_net_13225)
	);

	bfr new_net_13226_bfr_after (
		.din(new_net_13225),
		.dout(new_net_13226)
	);

	bfr new_net_13227_bfr_after (
		.din(new_net_13226),
		.dout(new_net_13227)
	);

	bfr new_net_13228_bfr_after (
		.din(new_net_13227),
		.dout(new_net_13228)
	);

	bfr new_net_13229_bfr_after (
		.din(new_net_13228),
		.dout(new_net_13229)
	);

	bfr new_net_13230_bfr_after (
		.din(new_net_13229),
		.dout(new_net_13230)
	);

	bfr new_net_13231_bfr_after (
		.din(new_net_13230),
		.dout(new_net_13231)
	);

	bfr new_net_13232_bfr_after (
		.din(new_net_13231),
		.dout(new_net_13232)
	);

	bfr new_net_13233_bfr_after (
		.din(new_net_13232),
		.dout(new_net_13233)
	);

	bfr new_net_13234_bfr_after (
		.din(new_net_13233),
		.dout(new_net_13234)
	);

	bfr new_net_13235_bfr_after (
		.din(new_net_13234),
		.dout(new_net_13235)
	);

	bfr new_net_13236_bfr_after (
		.din(new_net_13235),
		.dout(new_net_13236)
	);

	bfr new_net_13237_bfr_after (
		.din(new_net_13236),
		.dout(new_net_13237)
	);

	bfr new_net_13238_bfr_after (
		.din(new_net_13237),
		.dout(new_net_13238)
	);

	bfr new_net_13239_bfr_after (
		.din(new_net_13238),
		.dout(new_net_13239)
	);

	bfr new_net_13240_bfr_after (
		.din(new_net_13239),
		.dout(new_net_13240)
	);

	bfr new_net_13241_bfr_after (
		.din(new_net_13240),
		.dout(new_net_13241)
	);

	bfr new_net_13242_bfr_after (
		.din(new_net_13241),
		.dout(new_net_13242)
	);

	bfr new_net_13243_bfr_after (
		.din(new_net_13242),
		.dout(new_net_13243)
	);

	bfr new_net_13244_bfr_after (
		.din(new_net_13243),
		.dout(new_net_13244)
	);

	bfr new_net_13245_bfr_after (
		.din(new_net_13244),
		.dout(new_net_13245)
	);

	bfr new_net_13246_bfr_after (
		.din(new_net_13245),
		.dout(new_net_13246)
	);

	bfr new_net_13247_bfr_after (
		.din(new_net_13246),
		.dout(new_net_13247)
	);

	bfr new_net_13248_bfr_after (
		.din(new_net_13247),
		.dout(new_net_13248)
	);

	bfr new_net_13249_bfr_after (
		.din(new_net_13248),
		.dout(new_net_13249)
	);

	bfr new_net_13250_bfr_after (
		.din(new_net_13249),
		.dout(new_net_13250)
	);

	bfr new_net_13251_bfr_after (
		.din(new_net_13250),
		.dout(new_net_13251)
	);

	bfr new_net_13252_bfr_after (
		.din(new_net_13251),
		.dout(new_net_13252)
	);

	bfr new_net_13253_bfr_after (
		.din(new_net_13252),
		.dout(new_net_13253)
	);

	spl2 _0434__v_fanout (
		.a(new_net_13253),
		.b(new_net_26),
		.c(new_net_27)
	);

	bfr new_net_13254_bfr_after (
		.din(_1819_),
		.dout(new_net_13254)
	);

	bfr new_net_13255_bfr_after (
		.din(new_net_13254),
		.dout(new_net_13255)
	);

	bfr new_net_13256_bfr_after (
		.din(new_net_13255),
		.dout(new_net_13256)
	);

	bfr new_net_13257_bfr_after (
		.din(new_net_13256),
		.dout(new_net_13257)
	);

	bfr new_net_13258_bfr_after (
		.din(new_net_13257),
		.dout(new_net_13258)
	);

	bfr new_net_13259_bfr_after (
		.din(new_net_13258),
		.dout(new_net_13259)
	);

	bfr new_net_13260_bfr_after (
		.din(new_net_13259),
		.dout(new_net_13260)
	);

	bfr new_net_13261_bfr_after (
		.din(new_net_13260),
		.dout(new_net_13261)
	);

	bfr new_net_13262_bfr_after (
		.din(new_net_13261),
		.dout(new_net_13262)
	);

	bfr new_net_13263_bfr_after (
		.din(new_net_13262),
		.dout(new_net_13263)
	);

	bfr new_net_13264_bfr_after (
		.din(new_net_13263),
		.dout(new_net_13264)
	);

	bfr new_net_13265_bfr_after (
		.din(new_net_13264),
		.dout(new_net_13265)
	);

	bfr new_net_13266_bfr_after (
		.din(new_net_13265),
		.dout(new_net_13266)
	);

	bfr new_net_13267_bfr_after (
		.din(new_net_13266),
		.dout(new_net_13267)
	);

	bfr new_net_13268_bfr_after (
		.din(new_net_13267),
		.dout(new_net_13268)
	);

	bfr new_net_13269_bfr_after (
		.din(new_net_13268),
		.dout(new_net_13269)
	);

	bfr new_net_13270_bfr_after (
		.din(new_net_13269),
		.dout(new_net_13270)
	);

	bfr new_net_13271_bfr_after (
		.din(new_net_13270),
		.dout(new_net_13271)
	);

	bfr new_net_13272_bfr_after (
		.din(new_net_13271),
		.dout(new_net_13272)
	);

	bfr new_net_13273_bfr_after (
		.din(new_net_13272),
		.dout(new_net_13273)
	);

	bfr new_net_13274_bfr_after (
		.din(new_net_13273),
		.dout(new_net_13274)
	);

	bfr new_net_13275_bfr_after (
		.din(new_net_13274),
		.dout(new_net_13275)
	);

	bfr new_net_13276_bfr_after (
		.din(new_net_13275),
		.dout(new_net_13276)
	);

	bfr new_net_13277_bfr_after (
		.din(new_net_13276),
		.dout(new_net_13277)
	);

	bfr new_net_13278_bfr_after (
		.din(new_net_13277),
		.dout(new_net_13278)
	);

	bfr new_net_13279_bfr_after (
		.din(new_net_13278),
		.dout(new_net_13279)
	);

	bfr new_net_13280_bfr_after (
		.din(new_net_13279),
		.dout(new_net_13280)
	);

	bfr new_net_13281_bfr_after (
		.din(new_net_13280),
		.dout(new_net_13281)
	);

	bfr new_net_13282_bfr_after (
		.din(new_net_13281),
		.dout(new_net_13282)
	);

	bfr new_net_13283_bfr_after (
		.din(new_net_13282),
		.dout(new_net_13283)
	);

	bfr new_net_13284_bfr_after (
		.din(new_net_13283),
		.dout(new_net_13284)
	);

	bfr new_net_13285_bfr_after (
		.din(new_net_13284),
		.dout(new_net_13285)
	);

	bfr new_net_13286_bfr_after (
		.din(new_net_13285),
		.dout(new_net_13286)
	);

	bfr new_net_13287_bfr_after (
		.din(new_net_13286),
		.dout(new_net_13287)
	);

	bfr new_net_13288_bfr_after (
		.din(new_net_13287),
		.dout(new_net_13288)
	);

	bfr new_net_13289_bfr_after (
		.din(new_net_13288),
		.dout(new_net_13289)
	);

	bfr new_net_13290_bfr_after (
		.din(new_net_13289),
		.dout(new_net_13290)
	);

	bfr new_net_13291_bfr_after (
		.din(new_net_13290),
		.dout(new_net_13291)
	);

	bfr new_net_13292_bfr_after (
		.din(new_net_13291),
		.dout(new_net_13292)
	);

	bfr new_net_13293_bfr_after (
		.din(new_net_13292),
		.dout(new_net_13293)
	);

	bfr new_net_13294_bfr_after (
		.din(new_net_13293),
		.dout(new_net_13294)
	);

	bfr new_net_13295_bfr_after (
		.din(new_net_13294),
		.dout(new_net_13295)
	);

	bfr new_net_13296_bfr_after (
		.din(new_net_13295),
		.dout(new_net_13296)
	);

	bfr new_net_13297_bfr_after (
		.din(new_net_13296),
		.dout(new_net_13297)
	);

	bfr new_net_13298_bfr_after (
		.din(new_net_13297),
		.dout(new_net_13298)
	);

	bfr new_net_13299_bfr_after (
		.din(new_net_13298),
		.dout(new_net_13299)
	);

	bfr new_net_13300_bfr_after (
		.din(new_net_13299),
		.dout(new_net_13300)
	);

	bfr new_net_13301_bfr_after (
		.din(new_net_13300),
		.dout(new_net_13301)
	);

	spl2 _1819__v_fanout (
		.a(new_net_13301),
		.b(new_net_1698),
		.c(new_net_1699)
	);

	bfr new_net_13302_bfr_after (
		.din(_0838_),
		.dout(new_net_13302)
	);

	bfr new_net_13303_bfr_after (
		.din(new_net_13302),
		.dout(new_net_13303)
	);

	bfr new_net_13304_bfr_after (
		.din(new_net_13303),
		.dout(new_net_13304)
	);

	bfr new_net_13305_bfr_after (
		.din(new_net_13304),
		.dout(new_net_13305)
	);

	bfr new_net_13306_bfr_after (
		.din(new_net_13305),
		.dout(new_net_13306)
	);

	bfr new_net_13307_bfr_after (
		.din(new_net_13306),
		.dout(new_net_13307)
	);

	bfr new_net_13308_bfr_after (
		.din(new_net_13307),
		.dout(new_net_13308)
	);

	bfr new_net_13309_bfr_after (
		.din(new_net_13308),
		.dout(new_net_13309)
	);

	bfr new_net_13310_bfr_after (
		.din(new_net_13309),
		.dout(new_net_13310)
	);

	bfr new_net_13311_bfr_after (
		.din(new_net_13310),
		.dout(new_net_13311)
	);

	bfr new_net_13312_bfr_after (
		.din(new_net_13311),
		.dout(new_net_13312)
	);

	bfr new_net_13313_bfr_after (
		.din(new_net_13312),
		.dout(new_net_13313)
	);

	bfr new_net_13314_bfr_after (
		.din(new_net_13313),
		.dout(new_net_13314)
	);

	bfr new_net_13315_bfr_after (
		.din(new_net_13314),
		.dout(new_net_13315)
	);

	bfr new_net_13316_bfr_after (
		.din(new_net_13315),
		.dout(new_net_13316)
	);

	bfr new_net_13317_bfr_after (
		.din(new_net_13316),
		.dout(new_net_13317)
	);

	bfr new_net_13318_bfr_after (
		.din(new_net_13317),
		.dout(new_net_13318)
	);

	bfr new_net_13319_bfr_after (
		.din(new_net_13318),
		.dout(new_net_13319)
	);

	bfr new_net_13320_bfr_after (
		.din(new_net_13319),
		.dout(new_net_13320)
	);

	bfr new_net_13321_bfr_after (
		.din(new_net_13320),
		.dout(new_net_13321)
	);

	bfr new_net_13322_bfr_after (
		.din(new_net_13321),
		.dout(new_net_13322)
	);

	bfr new_net_13323_bfr_after (
		.din(new_net_13322),
		.dout(new_net_13323)
	);

	bfr new_net_13324_bfr_after (
		.din(new_net_13323),
		.dout(new_net_13324)
	);

	bfr new_net_13325_bfr_after (
		.din(new_net_13324),
		.dout(new_net_13325)
	);

	bfr new_net_13326_bfr_after (
		.din(new_net_13325),
		.dout(new_net_13326)
	);

	bfr new_net_13327_bfr_after (
		.din(new_net_13326),
		.dout(new_net_13327)
	);

	bfr new_net_13328_bfr_after (
		.din(new_net_13327),
		.dout(new_net_13328)
	);

	bfr new_net_13329_bfr_after (
		.din(new_net_13328),
		.dout(new_net_13329)
	);

	bfr new_net_13330_bfr_after (
		.din(new_net_13329),
		.dout(new_net_13330)
	);

	bfr new_net_13331_bfr_after (
		.din(new_net_13330),
		.dout(new_net_13331)
	);

	bfr new_net_13332_bfr_after (
		.din(new_net_13331),
		.dout(new_net_13332)
	);

	bfr new_net_13333_bfr_after (
		.din(new_net_13332),
		.dout(new_net_13333)
	);

	bfr new_net_13334_bfr_after (
		.din(new_net_13333),
		.dout(new_net_13334)
	);

	bfr new_net_13335_bfr_after (
		.din(new_net_13334),
		.dout(new_net_13335)
	);

	bfr new_net_13336_bfr_after (
		.din(new_net_13335),
		.dout(new_net_13336)
	);

	bfr new_net_13337_bfr_after (
		.din(new_net_13336),
		.dout(new_net_13337)
	);

	bfr new_net_13338_bfr_after (
		.din(new_net_13337),
		.dout(new_net_13338)
	);

	bfr new_net_13339_bfr_after (
		.din(new_net_13338),
		.dout(new_net_13339)
	);

	bfr new_net_13340_bfr_after (
		.din(new_net_13339),
		.dout(new_net_13340)
	);

	bfr new_net_13341_bfr_after (
		.din(new_net_13340),
		.dout(new_net_13341)
	);

	bfr new_net_13342_bfr_after (
		.din(new_net_13341),
		.dout(new_net_13342)
	);

	bfr new_net_13343_bfr_after (
		.din(new_net_13342),
		.dout(new_net_13343)
	);

	bfr new_net_13344_bfr_after (
		.din(new_net_13343),
		.dout(new_net_13344)
	);

	bfr new_net_13345_bfr_after (
		.din(new_net_13344),
		.dout(new_net_13345)
	);

	bfr new_net_13346_bfr_after (
		.din(new_net_13345),
		.dout(new_net_13346)
	);

	bfr new_net_13347_bfr_after (
		.din(new_net_13346),
		.dout(new_net_13347)
	);

	bfr new_net_13348_bfr_after (
		.din(new_net_13347),
		.dout(new_net_13348)
	);

	bfr new_net_13349_bfr_after (
		.din(new_net_13348),
		.dout(new_net_13349)
	);

	bfr new_net_13350_bfr_after (
		.din(new_net_13349),
		.dout(new_net_13350)
	);

	bfr new_net_13351_bfr_after (
		.din(new_net_13350),
		.dout(new_net_13351)
	);

	bfr new_net_13352_bfr_after (
		.din(new_net_13351),
		.dout(new_net_13352)
	);

	bfr new_net_13353_bfr_after (
		.din(new_net_13352),
		.dout(new_net_13353)
	);

	bfr new_net_13354_bfr_after (
		.din(new_net_13353),
		.dout(new_net_13354)
	);

	bfr new_net_13355_bfr_after (
		.din(new_net_13354),
		.dout(new_net_13355)
	);

	bfr new_net_13356_bfr_after (
		.din(new_net_13355),
		.dout(new_net_13356)
	);

	bfr new_net_13357_bfr_after (
		.din(new_net_13356),
		.dout(new_net_13357)
	);

	bfr new_net_13358_bfr_after (
		.din(new_net_13357),
		.dout(new_net_13358)
	);

	bfr new_net_13359_bfr_after (
		.din(new_net_13358),
		.dout(new_net_13359)
	);

	bfr new_net_13360_bfr_after (
		.din(new_net_13359),
		.dout(new_net_13360)
	);

	bfr new_net_13361_bfr_after (
		.din(new_net_13360),
		.dout(new_net_13361)
	);

	bfr new_net_13362_bfr_after (
		.din(new_net_13361),
		.dout(new_net_13362)
	);

	bfr new_net_13363_bfr_after (
		.din(new_net_13362),
		.dout(new_net_13363)
	);

	bfr new_net_13364_bfr_after (
		.din(new_net_13363),
		.dout(new_net_13364)
	);

	bfr new_net_13365_bfr_after (
		.din(new_net_13364),
		.dout(new_net_13365)
	);

	bfr new_net_13366_bfr_after (
		.din(new_net_13365),
		.dout(new_net_13366)
	);

	bfr new_net_13367_bfr_after (
		.din(new_net_13366),
		.dout(new_net_13367)
	);

	bfr new_net_13368_bfr_after (
		.din(new_net_13367),
		.dout(new_net_13368)
	);

	bfr new_net_13369_bfr_after (
		.din(new_net_13368),
		.dout(new_net_13369)
	);

	bfr new_net_13370_bfr_after (
		.din(new_net_13369),
		.dout(new_net_13370)
	);

	bfr new_net_13371_bfr_after (
		.din(new_net_13370),
		.dout(new_net_13371)
	);

	spl2 _0838__v_fanout (
		.a(new_net_13371),
		.b(new_net_2593),
		.c(new_net_2594)
	);

	bfr new_net_13372_bfr_after (
		.din(_1026_),
		.dout(new_net_13372)
	);

	bfr new_net_13373_bfr_after (
		.din(new_net_13372),
		.dout(new_net_13373)
	);

	bfr new_net_13374_bfr_after (
		.din(new_net_13373),
		.dout(new_net_13374)
	);

	bfr new_net_13375_bfr_after (
		.din(new_net_13374),
		.dout(new_net_13375)
	);

	bfr new_net_13376_bfr_after (
		.din(new_net_13375),
		.dout(new_net_13376)
	);

	bfr new_net_13377_bfr_after (
		.din(new_net_13376),
		.dout(new_net_13377)
	);

	bfr new_net_13378_bfr_after (
		.din(new_net_13377),
		.dout(new_net_13378)
	);

	bfr new_net_13379_bfr_after (
		.din(new_net_13378),
		.dout(new_net_13379)
	);

	bfr new_net_13380_bfr_after (
		.din(new_net_13379),
		.dout(new_net_13380)
	);

	bfr new_net_13381_bfr_after (
		.din(new_net_13380),
		.dout(new_net_13381)
	);

	bfr new_net_13382_bfr_after (
		.din(new_net_13381),
		.dout(new_net_13382)
	);

	bfr new_net_13383_bfr_after (
		.din(new_net_13382),
		.dout(new_net_13383)
	);

	bfr new_net_13384_bfr_after (
		.din(new_net_13383),
		.dout(new_net_13384)
	);

	bfr new_net_13385_bfr_after (
		.din(new_net_13384),
		.dout(new_net_13385)
	);

	bfr new_net_13386_bfr_after (
		.din(new_net_13385),
		.dout(new_net_13386)
	);

	bfr new_net_13387_bfr_after (
		.din(new_net_13386),
		.dout(new_net_13387)
	);

	bfr new_net_13388_bfr_after (
		.din(new_net_13387),
		.dout(new_net_13388)
	);

	bfr new_net_13389_bfr_after (
		.din(new_net_13388),
		.dout(new_net_13389)
	);

	bfr new_net_13390_bfr_after (
		.din(new_net_13389),
		.dout(new_net_13390)
	);

	bfr new_net_13391_bfr_after (
		.din(new_net_13390),
		.dout(new_net_13391)
	);

	bfr new_net_13392_bfr_after (
		.din(new_net_13391),
		.dout(new_net_13392)
	);

	bfr new_net_13393_bfr_after (
		.din(new_net_13392),
		.dout(new_net_13393)
	);

	bfr new_net_13394_bfr_after (
		.din(new_net_13393),
		.dout(new_net_13394)
	);

	bfr new_net_13395_bfr_after (
		.din(new_net_13394),
		.dout(new_net_13395)
	);

	spl2 _1026__v_fanout (
		.a(new_net_13395),
		.b(new_net_168),
		.c(new_net_169)
	);

	bfr new_net_13396_bfr_after (
		.din(_0450_),
		.dout(new_net_13396)
	);

	bfr new_net_13397_bfr_after (
		.din(new_net_13396),
		.dout(new_net_13397)
	);

	bfr new_net_13398_bfr_after (
		.din(new_net_13397),
		.dout(new_net_13398)
	);

	bfr new_net_13399_bfr_after (
		.din(new_net_13398),
		.dout(new_net_13399)
	);

	bfr new_net_13400_bfr_after (
		.din(new_net_13399),
		.dout(new_net_13400)
	);

	bfr new_net_13401_bfr_after (
		.din(new_net_13400),
		.dout(new_net_13401)
	);

	bfr new_net_13402_bfr_after (
		.din(new_net_13401),
		.dout(new_net_13402)
	);

	bfr new_net_13403_bfr_after (
		.din(new_net_13402),
		.dout(new_net_13403)
	);

	bfr new_net_13404_bfr_after (
		.din(new_net_13403),
		.dout(new_net_13404)
	);

	bfr new_net_13405_bfr_after (
		.din(new_net_13404),
		.dout(new_net_13405)
	);

	bfr new_net_13406_bfr_after (
		.din(new_net_13405),
		.dout(new_net_13406)
	);

	bfr new_net_13407_bfr_after (
		.din(new_net_13406),
		.dout(new_net_13407)
	);

	bfr new_net_13408_bfr_after (
		.din(new_net_13407),
		.dout(new_net_13408)
	);

	bfr new_net_13409_bfr_after (
		.din(new_net_13408),
		.dout(new_net_13409)
	);

	bfr new_net_13410_bfr_after (
		.din(new_net_13409),
		.dout(new_net_13410)
	);

	bfr new_net_13411_bfr_after (
		.din(new_net_13410),
		.dout(new_net_13411)
	);

	bfr new_net_13412_bfr_after (
		.din(new_net_13411),
		.dout(new_net_13412)
	);

	bfr new_net_13413_bfr_after (
		.din(new_net_13412),
		.dout(new_net_13413)
	);

	bfr new_net_13414_bfr_after (
		.din(new_net_13413),
		.dout(new_net_13414)
	);

	bfr new_net_13415_bfr_after (
		.din(new_net_13414),
		.dout(new_net_13415)
	);

	bfr new_net_13416_bfr_after (
		.din(new_net_13415),
		.dout(new_net_13416)
	);

	bfr new_net_13417_bfr_after (
		.din(new_net_13416),
		.dout(new_net_13417)
	);

	bfr new_net_13418_bfr_after (
		.din(new_net_13417),
		.dout(new_net_13418)
	);

	bfr new_net_13419_bfr_after (
		.din(new_net_13418),
		.dout(new_net_13419)
	);

	bfr new_net_13420_bfr_after (
		.din(new_net_13419),
		.dout(new_net_13420)
	);

	bfr new_net_13421_bfr_after (
		.din(new_net_13420),
		.dout(new_net_13421)
	);

	bfr new_net_13422_bfr_after (
		.din(new_net_13421),
		.dout(new_net_13422)
	);

	bfr new_net_13423_bfr_after (
		.din(new_net_13422),
		.dout(new_net_13423)
	);

	bfr new_net_13424_bfr_after (
		.din(new_net_13423),
		.dout(new_net_13424)
	);

	bfr new_net_13425_bfr_after (
		.din(new_net_13424),
		.dout(new_net_13425)
	);

	bfr new_net_13426_bfr_after (
		.din(new_net_13425),
		.dout(new_net_13426)
	);

	bfr new_net_13427_bfr_after (
		.din(new_net_13426),
		.dout(new_net_13427)
	);

	bfr new_net_13428_bfr_after (
		.din(new_net_13427),
		.dout(new_net_13428)
	);

	bfr new_net_13429_bfr_after (
		.din(new_net_13428),
		.dout(new_net_13429)
	);

	bfr new_net_13430_bfr_after (
		.din(new_net_13429),
		.dout(new_net_13430)
	);

	bfr new_net_13431_bfr_after (
		.din(new_net_13430),
		.dout(new_net_13431)
	);

	bfr new_net_13432_bfr_after (
		.din(new_net_13431),
		.dout(new_net_13432)
	);

	bfr new_net_13433_bfr_after (
		.din(new_net_13432),
		.dout(new_net_13433)
	);

	bfr new_net_13434_bfr_after (
		.din(new_net_13433),
		.dout(new_net_13434)
	);

	bfr new_net_13435_bfr_after (
		.din(new_net_13434),
		.dout(new_net_13435)
	);

	bfr new_net_13436_bfr_after (
		.din(new_net_13435),
		.dout(new_net_13436)
	);

	bfr new_net_13437_bfr_after (
		.din(new_net_13436),
		.dout(new_net_13437)
	);

	bfr new_net_13438_bfr_after (
		.din(new_net_13437),
		.dout(new_net_13438)
	);

	bfr new_net_13439_bfr_after (
		.din(new_net_13438),
		.dout(new_net_13439)
	);

	bfr new_net_13440_bfr_after (
		.din(new_net_13439),
		.dout(new_net_13440)
	);

	bfr new_net_13441_bfr_after (
		.din(new_net_13440),
		.dout(new_net_13441)
	);

	spl2 _0450__v_fanout (
		.a(new_net_13441),
		.b(new_net_3061),
		.c(new_net_3062)
	);

	bfr new_net_13442_bfr_after (
		.din(_1074_),
		.dout(new_net_13442)
	);

	bfr new_net_13443_bfr_after (
		.din(new_net_13442),
		.dout(new_net_13443)
	);

	bfr new_net_13444_bfr_after (
		.din(new_net_13443),
		.dout(new_net_13444)
	);

	bfr new_net_13445_bfr_after (
		.din(new_net_13444),
		.dout(new_net_13445)
	);

	bfr new_net_13446_bfr_after (
		.din(new_net_13445),
		.dout(new_net_13446)
	);

	bfr new_net_13447_bfr_after (
		.din(new_net_13446),
		.dout(new_net_13447)
	);

	bfr new_net_13448_bfr_after (
		.din(new_net_13447),
		.dout(new_net_13448)
	);

	bfr new_net_13449_bfr_after (
		.din(new_net_13448),
		.dout(new_net_13449)
	);

	bfr new_net_13450_bfr_after (
		.din(new_net_13449),
		.dout(new_net_13450)
	);

	bfr new_net_13451_bfr_after (
		.din(new_net_13450),
		.dout(new_net_13451)
	);

	bfr new_net_13452_bfr_after (
		.din(new_net_13451),
		.dout(new_net_13452)
	);

	bfr new_net_13453_bfr_after (
		.din(new_net_13452),
		.dout(new_net_13453)
	);

	bfr new_net_13454_bfr_after (
		.din(new_net_13453),
		.dout(new_net_13454)
	);

	bfr new_net_13455_bfr_after (
		.din(new_net_13454),
		.dout(new_net_13455)
	);

	bfr new_net_13456_bfr_after (
		.din(new_net_13455),
		.dout(new_net_13456)
	);

	bfr new_net_13457_bfr_after (
		.din(new_net_13456),
		.dout(new_net_13457)
	);

	bfr new_net_13458_bfr_after (
		.din(new_net_13457),
		.dout(new_net_13458)
	);

	bfr new_net_13459_bfr_after (
		.din(new_net_13458),
		.dout(new_net_13459)
	);

	bfr new_net_13460_bfr_after (
		.din(new_net_13459),
		.dout(new_net_13460)
	);

	bfr new_net_13461_bfr_after (
		.din(new_net_13460),
		.dout(new_net_13461)
	);

	bfr new_net_13462_bfr_after (
		.din(new_net_13461),
		.dout(new_net_13462)
	);

	bfr new_net_13463_bfr_after (
		.din(new_net_13462),
		.dout(new_net_13463)
	);

	bfr new_net_13464_bfr_after (
		.din(new_net_13463),
		.dout(new_net_13464)
	);

	bfr new_net_13465_bfr_after (
		.din(new_net_13464),
		.dout(new_net_13465)
	);

	bfr new_net_13466_bfr_after (
		.din(new_net_13465),
		.dout(new_net_13466)
	);

	bfr new_net_13467_bfr_after (
		.din(new_net_13466),
		.dout(new_net_13467)
	);

	bfr new_net_13468_bfr_after (
		.din(new_net_13467),
		.dout(new_net_13468)
	);

	bfr new_net_13469_bfr_after (
		.din(new_net_13468),
		.dout(new_net_13469)
	);

	bfr new_net_13470_bfr_after (
		.din(new_net_13469),
		.dout(new_net_13470)
	);

	bfr new_net_13471_bfr_after (
		.din(new_net_13470),
		.dout(new_net_13471)
	);

	bfr new_net_13472_bfr_after (
		.din(new_net_13471),
		.dout(new_net_13472)
	);

	bfr new_net_13473_bfr_after (
		.din(new_net_13472),
		.dout(new_net_13473)
	);

	bfr new_net_13474_bfr_after (
		.din(new_net_13473),
		.dout(new_net_13474)
	);

	bfr new_net_13475_bfr_after (
		.din(new_net_13474),
		.dout(new_net_13475)
	);

	bfr new_net_13476_bfr_after (
		.din(new_net_13475),
		.dout(new_net_13476)
	);

	bfr new_net_13477_bfr_after (
		.din(new_net_13476),
		.dout(new_net_13477)
	);

	bfr new_net_13478_bfr_after (
		.din(new_net_13477),
		.dout(new_net_13478)
	);

	bfr new_net_13479_bfr_after (
		.din(new_net_13478),
		.dout(new_net_13479)
	);

	bfr new_net_13480_bfr_after (
		.din(new_net_13479),
		.dout(new_net_13480)
	);

	bfr new_net_13481_bfr_after (
		.din(new_net_13480),
		.dout(new_net_13481)
	);

	spl2 _1074__v_fanout (
		.a(new_net_13481),
		.b(new_net_522),
		.c(new_net_523)
	);

	bfr new_net_13482_bfr_after (
		.din(_1560_),
		.dout(new_net_13482)
	);

	bfr new_net_13483_bfr_after (
		.din(new_net_13482),
		.dout(new_net_13483)
	);

	bfr new_net_13484_bfr_after (
		.din(new_net_13483),
		.dout(new_net_13484)
	);

	bfr new_net_13485_bfr_after (
		.din(new_net_13484),
		.dout(new_net_13485)
	);

	bfr new_net_13486_bfr_after (
		.din(new_net_13485),
		.dout(new_net_13486)
	);

	bfr new_net_13487_bfr_after (
		.din(new_net_13486),
		.dout(new_net_13487)
	);

	bfr new_net_13488_bfr_after (
		.din(new_net_13487),
		.dout(new_net_13488)
	);

	bfr new_net_13489_bfr_after (
		.din(new_net_13488),
		.dout(new_net_13489)
	);

	bfr new_net_13490_bfr_after (
		.din(new_net_13489),
		.dout(new_net_13490)
	);

	bfr new_net_13491_bfr_after (
		.din(new_net_13490),
		.dout(new_net_13491)
	);

	bfr new_net_13492_bfr_after (
		.din(new_net_13491),
		.dout(new_net_13492)
	);

	bfr new_net_13493_bfr_after (
		.din(new_net_13492),
		.dout(new_net_13493)
	);

	bfr new_net_13494_bfr_after (
		.din(new_net_13493),
		.dout(new_net_13494)
	);

	bfr new_net_13495_bfr_after (
		.din(new_net_13494),
		.dout(new_net_13495)
	);

	bfr new_net_13496_bfr_after (
		.din(new_net_13495),
		.dout(new_net_13496)
	);

	bfr new_net_13497_bfr_after (
		.din(new_net_13496),
		.dout(new_net_13497)
	);

	bfr new_net_13498_bfr_after (
		.din(new_net_13497),
		.dout(new_net_13498)
	);

	bfr new_net_13499_bfr_after (
		.din(new_net_13498),
		.dout(new_net_13499)
	);

	bfr new_net_13500_bfr_after (
		.din(new_net_13499),
		.dout(new_net_13500)
	);

	bfr new_net_13501_bfr_after (
		.din(new_net_13500),
		.dout(new_net_13501)
	);

	bfr new_net_13502_bfr_after (
		.din(new_net_13501),
		.dout(new_net_13502)
	);

	bfr new_net_13503_bfr_after (
		.din(new_net_13502),
		.dout(new_net_13503)
	);

	bfr new_net_13504_bfr_after (
		.din(new_net_13503),
		.dout(new_net_13504)
	);

	bfr new_net_13505_bfr_after (
		.din(new_net_13504),
		.dout(new_net_13505)
	);

	bfr new_net_13506_bfr_after (
		.din(new_net_13505),
		.dout(new_net_13506)
	);

	bfr new_net_13507_bfr_after (
		.din(new_net_13506),
		.dout(new_net_13507)
	);

	bfr new_net_13508_bfr_after (
		.din(new_net_13507),
		.dout(new_net_13508)
	);

	bfr new_net_13509_bfr_after (
		.din(new_net_13508),
		.dout(new_net_13509)
	);

	bfr new_net_13510_bfr_after (
		.din(new_net_13509),
		.dout(new_net_13510)
	);

	bfr new_net_13511_bfr_after (
		.din(new_net_13510),
		.dout(new_net_13511)
	);

	bfr new_net_13512_bfr_after (
		.din(new_net_13511),
		.dout(new_net_13512)
	);

	bfr new_net_13513_bfr_after (
		.din(new_net_13512),
		.dout(new_net_13513)
	);

	bfr new_net_13514_bfr_after (
		.din(new_net_13513),
		.dout(new_net_13514)
	);

	bfr new_net_13515_bfr_after (
		.din(new_net_13514),
		.dout(new_net_13515)
	);

	bfr new_net_13516_bfr_after (
		.din(new_net_13515),
		.dout(new_net_13516)
	);

	bfr new_net_13517_bfr_after (
		.din(new_net_13516),
		.dout(new_net_13517)
	);

	bfr new_net_13518_bfr_after (
		.din(new_net_13517),
		.dout(new_net_13518)
	);

	bfr new_net_13519_bfr_after (
		.din(new_net_13518),
		.dout(new_net_13519)
	);

	bfr new_net_13520_bfr_after (
		.din(new_net_13519),
		.dout(new_net_13520)
	);

	bfr new_net_13521_bfr_after (
		.din(new_net_13520),
		.dout(new_net_13521)
	);

	bfr new_net_13522_bfr_after (
		.din(new_net_13521),
		.dout(new_net_13522)
	);

	bfr new_net_13523_bfr_after (
		.din(new_net_13522),
		.dout(new_net_13523)
	);

	bfr new_net_13524_bfr_after (
		.din(new_net_13523),
		.dout(new_net_13524)
	);

	bfr new_net_13525_bfr_after (
		.din(new_net_13524),
		.dout(new_net_13525)
	);

	bfr new_net_13526_bfr_after (
		.din(new_net_13525),
		.dout(new_net_13526)
	);

	bfr new_net_13527_bfr_after (
		.din(new_net_13526),
		.dout(new_net_13527)
	);

	bfr new_net_13528_bfr_after (
		.din(new_net_13527),
		.dout(new_net_13528)
	);

	bfr new_net_13529_bfr_after (
		.din(new_net_13528),
		.dout(new_net_13529)
	);

	bfr new_net_13530_bfr_after (
		.din(new_net_13529),
		.dout(new_net_13530)
	);

	bfr new_net_13531_bfr_after (
		.din(new_net_13530),
		.dout(new_net_13531)
	);

	bfr new_net_13532_bfr_after (
		.din(new_net_13531),
		.dout(new_net_13532)
	);

	bfr new_net_13533_bfr_after (
		.din(new_net_13532),
		.dout(new_net_13533)
	);

	bfr new_net_13534_bfr_after (
		.din(new_net_13533),
		.dout(new_net_13534)
	);

	bfr new_net_13535_bfr_after (
		.din(new_net_13534),
		.dout(new_net_13535)
	);

	bfr new_net_13536_bfr_after (
		.din(new_net_13535),
		.dout(new_net_13536)
	);

	bfr new_net_13537_bfr_after (
		.din(new_net_13536),
		.dout(new_net_13537)
	);

	bfr new_net_13538_bfr_after (
		.din(new_net_13537),
		.dout(new_net_13538)
	);

	bfr new_net_13539_bfr_after (
		.din(new_net_13538),
		.dout(new_net_13539)
	);

	bfr new_net_13540_bfr_after (
		.din(new_net_13539),
		.dout(new_net_13540)
	);

	bfr new_net_13541_bfr_after (
		.din(new_net_13540),
		.dout(new_net_13541)
	);

	bfr new_net_13542_bfr_after (
		.din(new_net_13541),
		.dout(new_net_13542)
	);

	bfr new_net_13543_bfr_after (
		.din(new_net_13542),
		.dout(new_net_13543)
	);

	bfr new_net_13544_bfr_after (
		.din(new_net_13543),
		.dout(new_net_13544)
	);

	bfr new_net_13545_bfr_after (
		.din(new_net_13544),
		.dout(new_net_13545)
	);

	bfr new_net_13546_bfr_after (
		.din(new_net_13545),
		.dout(new_net_13546)
	);

	bfr new_net_13547_bfr_after (
		.din(new_net_13546),
		.dout(new_net_13547)
	);

	bfr new_net_13548_bfr_after (
		.din(new_net_13547),
		.dout(new_net_13548)
	);

	bfr new_net_13549_bfr_after (
		.din(new_net_13548),
		.dout(new_net_13549)
	);

	bfr new_net_13550_bfr_after (
		.din(new_net_13549),
		.dout(new_net_13550)
	);

	bfr new_net_13551_bfr_after (
		.din(new_net_13550),
		.dout(new_net_13551)
	);

	bfr new_net_13552_bfr_after (
		.din(new_net_13551),
		.dout(new_net_13552)
	);

	bfr new_net_13553_bfr_after (
		.din(new_net_13552),
		.dout(new_net_13553)
	);

	bfr new_net_13554_bfr_after (
		.din(new_net_13553),
		.dout(new_net_13554)
	);

	bfr new_net_13555_bfr_after (
		.din(new_net_13554),
		.dout(new_net_13555)
	);

	bfr new_net_13556_bfr_after (
		.din(new_net_13555),
		.dout(new_net_13556)
	);

	bfr new_net_13557_bfr_after (
		.din(new_net_13556),
		.dout(new_net_13557)
	);

	bfr new_net_13558_bfr_after (
		.din(new_net_13557),
		.dout(new_net_13558)
	);

	bfr new_net_13559_bfr_after (
		.din(new_net_13558),
		.dout(new_net_13559)
	);

	bfr new_net_13560_bfr_after (
		.din(new_net_13559),
		.dout(new_net_13560)
	);

	bfr new_net_13561_bfr_after (
		.din(new_net_13560),
		.dout(new_net_13561)
	);

	bfr new_net_13562_bfr_after (
		.din(new_net_13561),
		.dout(new_net_13562)
	);

	bfr new_net_13563_bfr_after (
		.din(new_net_13562),
		.dout(new_net_13563)
	);

	bfr new_net_13564_bfr_after (
		.din(new_net_13563),
		.dout(new_net_13564)
	);

	bfr new_net_13565_bfr_after (
		.din(new_net_13564),
		.dout(new_net_13565)
	);

	bfr new_net_13566_bfr_after (
		.din(new_net_13565),
		.dout(new_net_13566)
	);

	bfr new_net_13567_bfr_after (
		.din(new_net_13566),
		.dout(new_net_13567)
	);

	bfr new_net_13568_bfr_after (
		.din(new_net_13567),
		.dout(new_net_13568)
	);

	bfr new_net_13569_bfr_after (
		.din(new_net_13568),
		.dout(new_net_13569)
	);

	bfr new_net_13570_bfr_after (
		.din(new_net_13569),
		.dout(new_net_13570)
	);

	bfr new_net_13571_bfr_after (
		.din(new_net_13570),
		.dout(new_net_13571)
	);

	bfr new_net_13572_bfr_after (
		.din(new_net_13571),
		.dout(new_net_13572)
	);

	bfr new_net_13573_bfr_after (
		.din(new_net_13572),
		.dout(new_net_13573)
	);

	bfr new_net_13574_bfr_after (
		.din(new_net_13573),
		.dout(new_net_13574)
	);

	bfr new_net_13575_bfr_after (
		.din(new_net_13574),
		.dout(new_net_13575)
	);

	bfr new_net_13576_bfr_after (
		.din(new_net_13575),
		.dout(new_net_13576)
	);

	bfr new_net_13577_bfr_after (
		.din(new_net_13576),
		.dout(new_net_13577)
	);

	bfr new_net_13578_bfr_after (
		.din(new_net_13577),
		.dout(new_net_13578)
	);

	bfr new_net_13579_bfr_after (
		.din(new_net_13578),
		.dout(new_net_13579)
	);

	bfr new_net_13580_bfr_after (
		.din(new_net_13579),
		.dout(new_net_13580)
	);

	bfr new_net_13581_bfr_after (
		.din(new_net_13580),
		.dout(new_net_13581)
	);

	bfr new_net_13582_bfr_after (
		.din(new_net_13581),
		.dout(new_net_13582)
	);

	bfr new_net_13583_bfr_after (
		.din(new_net_13582),
		.dout(new_net_13583)
	);

	bfr new_net_13584_bfr_after (
		.din(new_net_13583),
		.dout(new_net_13584)
	);

	bfr new_net_13585_bfr_after (
		.din(new_net_13584),
		.dout(new_net_13585)
	);

	spl2 _1560__v_fanout (
		.a(new_net_13585),
		.b(new_net_2903),
		.c(new_net_2904)
	);

	bfr new_net_13586_bfr_after (
		.din(_1698_),
		.dout(new_net_13586)
	);

	bfr new_net_13587_bfr_after (
		.din(new_net_13586),
		.dout(new_net_13587)
	);

	bfr new_net_13588_bfr_after (
		.din(new_net_13587),
		.dout(new_net_13588)
	);

	bfr new_net_13589_bfr_after (
		.din(new_net_13588),
		.dout(new_net_13589)
	);

	bfr new_net_13590_bfr_after (
		.din(new_net_13589),
		.dout(new_net_13590)
	);

	bfr new_net_13591_bfr_after (
		.din(new_net_13590),
		.dout(new_net_13591)
	);

	bfr new_net_13592_bfr_after (
		.din(new_net_13591),
		.dout(new_net_13592)
	);

	bfr new_net_13593_bfr_after (
		.din(new_net_13592),
		.dout(new_net_13593)
	);

	bfr new_net_13594_bfr_after (
		.din(new_net_13593),
		.dout(new_net_13594)
	);

	bfr new_net_13595_bfr_after (
		.din(new_net_13594),
		.dout(new_net_13595)
	);

	bfr new_net_13596_bfr_after (
		.din(new_net_13595),
		.dout(new_net_13596)
	);

	bfr new_net_13597_bfr_after (
		.din(new_net_13596),
		.dout(new_net_13597)
	);

	bfr new_net_13598_bfr_after (
		.din(new_net_13597),
		.dout(new_net_13598)
	);

	bfr new_net_13599_bfr_after (
		.din(new_net_13598),
		.dout(new_net_13599)
	);

	bfr new_net_13600_bfr_after (
		.din(new_net_13599),
		.dout(new_net_13600)
	);

	bfr new_net_13601_bfr_after (
		.din(new_net_13600),
		.dout(new_net_13601)
	);

	bfr new_net_13602_bfr_after (
		.din(new_net_13601),
		.dout(new_net_13602)
	);

	bfr new_net_13603_bfr_after (
		.din(new_net_13602),
		.dout(new_net_13603)
	);

	bfr new_net_13604_bfr_after (
		.din(new_net_13603),
		.dout(new_net_13604)
	);

	bfr new_net_13605_bfr_after (
		.din(new_net_13604),
		.dout(new_net_13605)
	);

	bfr new_net_13606_bfr_after (
		.din(new_net_13605),
		.dout(new_net_13606)
	);

	bfr new_net_13607_bfr_after (
		.din(new_net_13606),
		.dout(new_net_13607)
	);

	bfr new_net_13608_bfr_after (
		.din(new_net_13607),
		.dout(new_net_13608)
	);

	bfr new_net_13609_bfr_after (
		.din(new_net_13608),
		.dout(new_net_13609)
	);

	bfr new_net_13610_bfr_after (
		.din(new_net_13609),
		.dout(new_net_13610)
	);

	bfr new_net_13611_bfr_after (
		.din(new_net_13610),
		.dout(new_net_13611)
	);

	bfr new_net_13612_bfr_after (
		.din(new_net_13611),
		.dout(new_net_13612)
	);

	bfr new_net_13613_bfr_after (
		.din(new_net_13612),
		.dout(new_net_13613)
	);

	bfr new_net_13614_bfr_after (
		.din(new_net_13613),
		.dout(new_net_13614)
	);

	bfr new_net_13615_bfr_after (
		.din(new_net_13614),
		.dout(new_net_13615)
	);

	bfr new_net_13616_bfr_after (
		.din(new_net_13615),
		.dout(new_net_13616)
	);

	bfr new_net_13617_bfr_after (
		.din(new_net_13616),
		.dout(new_net_13617)
	);

	bfr new_net_13618_bfr_after (
		.din(new_net_13617),
		.dout(new_net_13618)
	);

	bfr new_net_13619_bfr_after (
		.din(new_net_13618),
		.dout(new_net_13619)
	);

	bfr new_net_13620_bfr_after (
		.din(new_net_13619),
		.dout(new_net_13620)
	);

	bfr new_net_13621_bfr_after (
		.din(new_net_13620),
		.dout(new_net_13621)
	);

	bfr new_net_13622_bfr_after (
		.din(new_net_13621),
		.dout(new_net_13622)
	);

	bfr new_net_13623_bfr_after (
		.din(new_net_13622),
		.dout(new_net_13623)
	);

	bfr new_net_13624_bfr_after (
		.din(new_net_13623),
		.dout(new_net_13624)
	);

	bfr new_net_13625_bfr_after (
		.din(new_net_13624),
		.dout(new_net_13625)
	);

	spl2 _1698__v_fanout (
		.a(new_net_13625),
		.b(new_net_291),
		.c(new_net_292)
	);

	bfr new_net_13626_bfr_after (
		.din(_0084_),
		.dout(new_net_13626)
	);

	bfr new_net_13627_bfr_after (
		.din(new_net_13626),
		.dout(new_net_13627)
	);

	bfr new_net_13628_bfr_after (
		.din(new_net_13627),
		.dout(new_net_13628)
	);

	bfr new_net_13629_bfr_after (
		.din(new_net_13628),
		.dout(new_net_13629)
	);

	bfr new_net_13630_bfr_after (
		.din(new_net_13629),
		.dout(new_net_13630)
	);

	bfr new_net_13631_bfr_after (
		.din(new_net_13630),
		.dout(new_net_13631)
	);

	bfr new_net_13632_bfr_after (
		.din(new_net_13631),
		.dout(new_net_13632)
	);

	bfr new_net_13633_bfr_after (
		.din(new_net_13632),
		.dout(new_net_13633)
	);

	bfr new_net_13634_bfr_after (
		.din(new_net_13633),
		.dout(new_net_13634)
	);

	bfr new_net_13635_bfr_after (
		.din(new_net_13634),
		.dout(new_net_13635)
	);

	bfr new_net_13636_bfr_after (
		.din(new_net_13635),
		.dout(new_net_13636)
	);

	bfr new_net_13637_bfr_after (
		.din(new_net_13636),
		.dout(new_net_13637)
	);

	bfr new_net_13638_bfr_after (
		.din(new_net_13637),
		.dout(new_net_13638)
	);

	bfr new_net_13639_bfr_after (
		.din(new_net_13638),
		.dout(new_net_13639)
	);

	bfr new_net_13640_bfr_after (
		.din(new_net_13639),
		.dout(new_net_13640)
	);

	bfr new_net_13641_bfr_after (
		.din(new_net_13640),
		.dout(new_net_13641)
	);

	bfr new_net_13642_bfr_after (
		.din(new_net_13641),
		.dout(new_net_13642)
	);

	bfr new_net_13643_bfr_after (
		.din(new_net_13642),
		.dout(new_net_13643)
	);

	bfr new_net_13644_bfr_after (
		.din(new_net_13643),
		.dout(new_net_13644)
	);

	bfr new_net_13645_bfr_after (
		.din(new_net_13644),
		.dout(new_net_13645)
	);

	bfr new_net_13646_bfr_after (
		.din(new_net_13645),
		.dout(new_net_13646)
	);

	bfr new_net_13647_bfr_after (
		.din(new_net_13646),
		.dout(new_net_13647)
	);

	bfr new_net_13648_bfr_after (
		.din(new_net_13647),
		.dout(new_net_13648)
	);

	bfr new_net_13649_bfr_after (
		.din(new_net_13648),
		.dout(new_net_13649)
	);

	bfr new_net_13650_bfr_after (
		.din(new_net_13649),
		.dout(new_net_13650)
	);

	bfr new_net_13651_bfr_after (
		.din(new_net_13650),
		.dout(new_net_13651)
	);

	bfr new_net_13652_bfr_after (
		.din(new_net_13651),
		.dout(new_net_13652)
	);

	bfr new_net_13653_bfr_after (
		.din(new_net_13652),
		.dout(new_net_13653)
	);

	bfr new_net_13654_bfr_after (
		.din(new_net_13653),
		.dout(new_net_13654)
	);

	bfr new_net_13655_bfr_after (
		.din(new_net_13654),
		.dout(new_net_13655)
	);

	bfr new_net_13656_bfr_after (
		.din(new_net_13655),
		.dout(new_net_13656)
	);

	bfr new_net_13657_bfr_after (
		.din(new_net_13656),
		.dout(new_net_13657)
	);

	bfr new_net_13658_bfr_after (
		.din(new_net_13657),
		.dout(new_net_13658)
	);

	bfr new_net_13659_bfr_after (
		.din(new_net_13658),
		.dout(new_net_13659)
	);

	bfr new_net_13660_bfr_after (
		.din(new_net_13659),
		.dout(new_net_13660)
	);

	bfr new_net_13661_bfr_after (
		.din(new_net_13660),
		.dout(new_net_13661)
	);

	bfr new_net_13662_bfr_after (
		.din(new_net_13661),
		.dout(new_net_13662)
	);

	bfr new_net_13663_bfr_after (
		.din(new_net_13662),
		.dout(new_net_13663)
	);

	bfr new_net_13664_bfr_after (
		.din(new_net_13663),
		.dout(new_net_13664)
	);

	bfr new_net_13665_bfr_after (
		.din(new_net_13664),
		.dout(new_net_13665)
	);

	bfr new_net_13666_bfr_after (
		.din(new_net_13665),
		.dout(new_net_13666)
	);

	bfr new_net_13667_bfr_after (
		.din(new_net_13666),
		.dout(new_net_13667)
	);

	bfr new_net_13668_bfr_after (
		.din(new_net_13667),
		.dout(new_net_13668)
	);

	bfr new_net_13669_bfr_after (
		.din(new_net_13668),
		.dout(new_net_13669)
	);

	bfr new_net_13670_bfr_after (
		.din(new_net_13669),
		.dout(new_net_13670)
	);

	bfr new_net_13671_bfr_after (
		.din(new_net_13670),
		.dout(new_net_13671)
	);

	bfr new_net_13672_bfr_after (
		.din(new_net_13671),
		.dout(new_net_13672)
	);

	bfr new_net_13673_bfr_after (
		.din(new_net_13672),
		.dout(new_net_13673)
	);

	bfr new_net_13674_bfr_after (
		.din(new_net_13673),
		.dout(new_net_13674)
	);

	bfr new_net_13675_bfr_after (
		.din(new_net_13674),
		.dout(new_net_13675)
	);

	bfr new_net_13676_bfr_after (
		.din(new_net_13675),
		.dout(new_net_13676)
	);

	bfr new_net_13677_bfr_after (
		.din(new_net_13676),
		.dout(new_net_13677)
	);

	bfr new_net_13678_bfr_after (
		.din(new_net_13677),
		.dout(new_net_13678)
	);

	bfr new_net_13679_bfr_after (
		.din(new_net_13678),
		.dout(new_net_13679)
	);

	bfr new_net_13680_bfr_after (
		.din(new_net_13679),
		.dout(new_net_13680)
	);

	bfr new_net_13681_bfr_after (
		.din(new_net_13680),
		.dout(new_net_13681)
	);

	bfr new_net_13682_bfr_after (
		.din(new_net_13681),
		.dout(new_net_13682)
	);

	bfr new_net_13683_bfr_after (
		.din(new_net_13682),
		.dout(new_net_13683)
	);

	bfr new_net_13684_bfr_after (
		.din(new_net_13683),
		.dout(new_net_13684)
	);

	bfr new_net_13685_bfr_after (
		.din(new_net_13684),
		.dout(new_net_13685)
	);

	bfr new_net_13686_bfr_after (
		.din(new_net_13685),
		.dout(new_net_13686)
	);

	bfr new_net_13687_bfr_after (
		.din(new_net_13686),
		.dout(new_net_13687)
	);

	bfr new_net_13688_bfr_after (
		.din(new_net_13687),
		.dout(new_net_13688)
	);

	bfr new_net_13689_bfr_after (
		.din(new_net_13688),
		.dout(new_net_13689)
	);

	bfr new_net_13690_bfr_after (
		.din(new_net_13689),
		.dout(new_net_13690)
	);

	bfr new_net_13691_bfr_after (
		.din(new_net_13690),
		.dout(new_net_13691)
	);

	bfr new_net_13692_bfr_after (
		.din(new_net_13691),
		.dout(new_net_13692)
	);

	bfr new_net_13693_bfr_after (
		.din(new_net_13692),
		.dout(new_net_13693)
	);

	bfr new_net_13694_bfr_after (
		.din(new_net_13693),
		.dout(new_net_13694)
	);

	bfr new_net_13695_bfr_after (
		.din(new_net_13694),
		.dout(new_net_13695)
	);

	bfr new_net_13696_bfr_after (
		.din(new_net_13695),
		.dout(new_net_13696)
	);

	bfr new_net_13697_bfr_after (
		.din(new_net_13696),
		.dout(new_net_13697)
	);

	bfr new_net_13698_bfr_after (
		.din(new_net_13697),
		.dout(new_net_13698)
	);

	bfr new_net_13699_bfr_after (
		.din(new_net_13698),
		.dout(new_net_13699)
	);

	bfr new_net_13700_bfr_after (
		.din(new_net_13699),
		.dout(new_net_13700)
	);

	bfr new_net_13701_bfr_after (
		.din(new_net_13700),
		.dout(new_net_13701)
	);

	bfr new_net_13702_bfr_after (
		.din(new_net_13701),
		.dout(new_net_13702)
	);

	bfr new_net_13703_bfr_after (
		.din(new_net_13702),
		.dout(new_net_13703)
	);

	bfr new_net_13704_bfr_after (
		.din(new_net_13703),
		.dout(new_net_13704)
	);

	bfr new_net_13705_bfr_after (
		.din(new_net_13704),
		.dout(new_net_13705)
	);

	bfr new_net_13706_bfr_after (
		.din(new_net_13705),
		.dout(new_net_13706)
	);

	bfr new_net_13707_bfr_after (
		.din(new_net_13706),
		.dout(new_net_13707)
	);

	bfr new_net_13708_bfr_after (
		.din(new_net_13707),
		.dout(new_net_13708)
	);

	bfr new_net_13709_bfr_after (
		.din(new_net_13708),
		.dout(new_net_13709)
	);

	bfr new_net_13710_bfr_after (
		.din(new_net_13709),
		.dout(new_net_13710)
	);

	bfr new_net_13711_bfr_after (
		.din(new_net_13710),
		.dout(new_net_13711)
	);

	bfr new_net_13712_bfr_after (
		.din(new_net_13711),
		.dout(new_net_13712)
	);

	bfr new_net_13713_bfr_after (
		.din(new_net_13712),
		.dout(new_net_13713)
	);

	bfr new_net_13714_bfr_after (
		.din(new_net_13713),
		.dout(new_net_13714)
	);

	bfr new_net_13715_bfr_after (
		.din(new_net_13714),
		.dout(new_net_13715)
	);

	bfr new_net_13716_bfr_after (
		.din(new_net_13715),
		.dout(new_net_13716)
	);

	bfr new_net_13717_bfr_after (
		.din(new_net_13716),
		.dout(new_net_13717)
	);

	bfr new_net_13718_bfr_after (
		.din(new_net_13717),
		.dout(new_net_13718)
	);

	bfr new_net_13719_bfr_after (
		.din(new_net_13718),
		.dout(new_net_13719)
	);

	bfr new_net_13720_bfr_after (
		.din(new_net_13719),
		.dout(new_net_13720)
	);

	bfr new_net_13721_bfr_after (
		.din(new_net_13720),
		.dout(new_net_13721)
	);

	bfr new_net_13722_bfr_after (
		.din(new_net_13721),
		.dout(new_net_13722)
	);

	bfr new_net_13723_bfr_after (
		.din(new_net_13722),
		.dout(new_net_13723)
	);

	bfr new_net_13724_bfr_after (
		.din(new_net_13723),
		.dout(new_net_13724)
	);

	bfr new_net_13725_bfr_after (
		.din(new_net_13724),
		.dout(new_net_13725)
	);

	bfr new_net_13726_bfr_after (
		.din(new_net_13725),
		.dout(new_net_13726)
	);

	bfr new_net_13727_bfr_after (
		.din(new_net_13726),
		.dout(new_net_13727)
	);

	bfr new_net_13728_bfr_after (
		.din(new_net_13727),
		.dout(new_net_13728)
	);

	bfr new_net_13729_bfr_after (
		.din(new_net_13728),
		.dout(new_net_13729)
	);

	bfr new_net_13730_bfr_after (
		.din(new_net_13729),
		.dout(new_net_13730)
	);

	bfr new_net_13731_bfr_after (
		.din(new_net_13730),
		.dout(new_net_13731)
	);

	bfr new_net_13732_bfr_after (
		.din(new_net_13731),
		.dout(new_net_13732)
	);

	bfr new_net_13733_bfr_after (
		.din(new_net_13732),
		.dout(new_net_13733)
	);

	bfr new_net_13734_bfr_after (
		.din(new_net_13733),
		.dout(new_net_13734)
	);

	bfr new_net_13735_bfr_after (
		.din(new_net_13734),
		.dout(new_net_13735)
	);

	bfr new_net_13736_bfr_after (
		.din(new_net_13735),
		.dout(new_net_13736)
	);

	bfr new_net_13737_bfr_after (
		.din(new_net_13736),
		.dout(new_net_13737)
	);

	spl2 _0084__v_fanout (
		.a(new_net_13737),
		.b(new_net_2667),
		.c(new_net_2668)
	);

	spl2 _0372__v_fanout (
		.a(_0372_),
		.b(new_net_142),
		.c(new_net_143)
	);

	bfr new_net_13738_bfr_after (
		.din(_1209_),
		.dout(new_net_13738)
	);

	bfr new_net_13739_bfr_after (
		.din(new_net_13738),
		.dout(new_net_13739)
	);

	bfr new_net_13740_bfr_after (
		.din(new_net_13739),
		.dout(new_net_13740)
	);

	bfr new_net_13741_bfr_after (
		.din(new_net_13740),
		.dout(new_net_13741)
	);

	bfr new_net_13742_bfr_after (
		.din(new_net_13741),
		.dout(new_net_13742)
	);

	bfr new_net_13743_bfr_after (
		.din(new_net_13742),
		.dout(new_net_13743)
	);

	bfr new_net_13744_bfr_after (
		.din(new_net_13743),
		.dout(new_net_13744)
	);

	bfr new_net_13745_bfr_after (
		.din(new_net_13744),
		.dout(new_net_13745)
	);

	bfr new_net_13746_bfr_after (
		.din(new_net_13745),
		.dout(new_net_13746)
	);

	bfr new_net_13747_bfr_after (
		.din(new_net_13746),
		.dout(new_net_13747)
	);

	bfr new_net_13748_bfr_after (
		.din(new_net_13747),
		.dout(new_net_13748)
	);

	bfr new_net_13749_bfr_after (
		.din(new_net_13748),
		.dout(new_net_13749)
	);

	bfr new_net_13750_bfr_after (
		.din(new_net_13749),
		.dout(new_net_13750)
	);

	bfr new_net_13751_bfr_after (
		.din(new_net_13750),
		.dout(new_net_13751)
	);

	bfr new_net_13752_bfr_after (
		.din(new_net_13751),
		.dout(new_net_13752)
	);

	bfr new_net_13753_bfr_after (
		.din(new_net_13752),
		.dout(new_net_13753)
	);

	bfr new_net_13754_bfr_after (
		.din(new_net_13753),
		.dout(new_net_13754)
	);

	bfr new_net_13755_bfr_after (
		.din(new_net_13754),
		.dout(new_net_13755)
	);

	bfr new_net_13756_bfr_after (
		.din(new_net_13755),
		.dout(new_net_13756)
	);

	bfr new_net_13757_bfr_after (
		.din(new_net_13756),
		.dout(new_net_13757)
	);

	bfr new_net_13758_bfr_after (
		.din(new_net_13757),
		.dout(new_net_13758)
	);

	bfr new_net_13759_bfr_after (
		.din(new_net_13758),
		.dout(new_net_13759)
	);

	bfr new_net_13760_bfr_after (
		.din(new_net_13759),
		.dout(new_net_13760)
	);

	bfr new_net_13761_bfr_after (
		.din(new_net_13760),
		.dout(new_net_13761)
	);

	bfr new_net_13762_bfr_after (
		.din(new_net_13761),
		.dout(new_net_13762)
	);

	bfr new_net_13763_bfr_after (
		.din(new_net_13762),
		.dout(new_net_13763)
	);

	bfr new_net_13764_bfr_after (
		.din(new_net_13763),
		.dout(new_net_13764)
	);

	bfr new_net_13765_bfr_after (
		.din(new_net_13764),
		.dout(new_net_13765)
	);

	bfr new_net_13766_bfr_after (
		.din(new_net_13765),
		.dout(new_net_13766)
	);

	bfr new_net_13767_bfr_after (
		.din(new_net_13766),
		.dout(new_net_13767)
	);

	bfr new_net_13768_bfr_after (
		.din(new_net_13767),
		.dout(new_net_13768)
	);

	bfr new_net_13769_bfr_after (
		.din(new_net_13768),
		.dout(new_net_13769)
	);

	bfr new_net_13770_bfr_after (
		.din(new_net_13769),
		.dout(new_net_13770)
	);

	bfr new_net_13771_bfr_after (
		.din(new_net_13770),
		.dout(new_net_13771)
	);

	bfr new_net_13772_bfr_after (
		.din(new_net_13771),
		.dout(new_net_13772)
	);

	bfr new_net_13773_bfr_after (
		.din(new_net_13772),
		.dout(new_net_13773)
	);

	bfr new_net_13774_bfr_after (
		.din(new_net_13773),
		.dout(new_net_13774)
	);

	bfr new_net_13775_bfr_after (
		.din(new_net_13774),
		.dout(new_net_13775)
	);

	bfr new_net_13776_bfr_after (
		.din(new_net_13775),
		.dout(new_net_13776)
	);

	bfr new_net_13777_bfr_after (
		.din(new_net_13776),
		.dout(new_net_13777)
	);

	bfr new_net_13778_bfr_after (
		.din(new_net_13777),
		.dout(new_net_13778)
	);

	bfr new_net_13779_bfr_after (
		.din(new_net_13778),
		.dout(new_net_13779)
	);

	bfr new_net_13780_bfr_after (
		.din(new_net_13779),
		.dout(new_net_13780)
	);

	bfr new_net_13781_bfr_after (
		.din(new_net_13780),
		.dout(new_net_13781)
	);

	bfr new_net_13782_bfr_after (
		.din(new_net_13781),
		.dout(new_net_13782)
	);

	bfr new_net_13783_bfr_after (
		.din(new_net_13782),
		.dout(new_net_13783)
	);

	bfr new_net_13784_bfr_after (
		.din(new_net_13783),
		.dout(new_net_13784)
	);

	bfr new_net_13785_bfr_after (
		.din(new_net_13784),
		.dout(new_net_13785)
	);

	spl2 _1209__v_fanout (
		.a(new_net_13785),
		.b(new_net_894),
		.c(new_net_895)
	);

	bfr new_net_13786_bfr_after (
		.din(_1586_),
		.dout(new_net_13786)
	);

	bfr new_net_13787_bfr_after (
		.din(new_net_13786),
		.dout(new_net_13787)
	);

	bfr new_net_13788_bfr_after (
		.din(new_net_13787),
		.dout(new_net_13788)
	);

	bfr new_net_13789_bfr_after (
		.din(new_net_13788),
		.dout(new_net_13789)
	);

	bfr new_net_13790_bfr_after (
		.din(new_net_13789),
		.dout(new_net_13790)
	);

	bfr new_net_13791_bfr_after (
		.din(new_net_13790),
		.dout(new_net_13791)
	);

	bfr new_net_13792_bfr_after (
		.din(new_net_13791),
		.dout(new_net_13792)
	);

	bfr new_net_13793_bfr_after (
		.din(new_net_13792),
		.dout(new_net_13793)
	);

	spl2 _1586__v_fanout (
		.a(new_net_13793),
		.b(new_net_2262),
		.c(new_net_2263)
	);

	bfr new_net_13794_bfr_after (
		.din(_0767_),
		.dout(new_net_13794)
	);

	bfr new_net_13795_bfr_after (
		.din(new_net_13794),
		.dout(new_net_13795)
	);

	bfr new_net_13796_bfr_after (
		.din(new_net_13795),
		.dout(new_net_13796)
	);

	bfr new_net_13797_bfr_after (
		.din(new_net_13796),
		.dout(new_net_13797)
	);

	bfr new_net_13798_bfr_after (
		.din(new_net_13797),
		.dout(new_net_13798)
	);

	bfr new_net_13799_bfr_after (
		.din(new_net_13798),
		.dout(new_net_13799)
	);

	bfr new_net_13800_bfr_after (
		.din(new_net_13799),
		.dout(new_net_13800)
	);

	bfr new_net_13801_bfr_after (
		.din(new_net_13800),
		.dout(new_net_13801)
	);

	bfr new_net_13802_bfr_after (
		.din(new_net_13801),
		.dout(new_net_13802)
	);

	bfr new_net_13803_bfr_after (
		.din(new_net_13802),
		.dout(new_net_13803)
	);

	bfr new_net_13804_bfr_after (
		.din(new_net_13803),
		.dout(new_net_13804)
	);

	bfr new_net_13805_bfr_after (
		.din(new_net_13804),
		.dout(new_net_13805)
	);

	bfr new_net_13806_bfr_after (
		.din(new_net_13805),
		.dout(new_net_13806)
	);

	bfr new_net_13807_bfr_after (
		.din(new_net_13806),
		.dout(new_net_13807)
	);

	bfr new_net_13808_bfr_after (
		.din(new_net_13807),
		.dout(new_net_13808)
	);

	bfr new_net_13809_bfr_after (
		.din(new_net_13808),
		.dout(new_net_13809)
	);

	bfr new_net_13810_bfr_after (
		.din(new_net_13809),
		.dout(new_net_13810)
	);

	bfr new_net_13811_bfr_after (
		.din(new_net_13810),
		.dout(new_net_13811)
	);

	bfr new_net_13812_bfr_after (
		.din(new_net_13811),
		.dout(new_net_13812)
	);

	bfr new_net_13813_bfr_after (
		.din(new_net_13812),
		.dout(new_net_13813)
	);

	bfr new_net_13814_bfr_after (
		.din(new_net_13813),
		.dout(new_net_13814)
	);

	bfr new_net_13815_bfr_after (
		.din(new_net_13814),
		.dout(new_net_13815)
	);

	bfr new_net_13816_bfr_after (
		.din(new_net_13815),
		.dout(new_net_13816)
	);

	bfr new_net_13817_bfr_after (
		.din(new_net_13816),
		.dout(new_net_13817)
	);

	bfr new_net_13818_bfr_after (
		.din(new_net_13817),
		.dout(new_net_13818)
	);

	bfr new_net_13819_bfr_after (
		.din(new_net_13818),
		.dout(new_net_13819)
	);

	bfr new_net_13820_bfr_after (
		.din(new_net_13819),
		.dout(new_net_13820)
	);

	bfr new_net_13821_bfr_after (
		.din(new_net_13820),
		.dout(new_net_13821)
	);

	bfr new_net_13822_bfr_after (
		.din(new_net_13821),
		.dout(new_net_13822)
	);

	bfr new_net_13823_bfr_after (
		.din(new_net_13822),
		.dout(new_net_13823)
	);

	bfr new_net_13824_bfr_after (
		.din(new_net_13823),
		.dout(new_net_13824)
	);

	bfr new_net_13825_bfr_after (
		.din(new_net_13824),
		.dout(new_net_13825)
	);

	bfr new_net_13826_bfr_after (
		.din(new_net_13825),
		.dout(new_net_13826)
	);

	bfr new_net_13827_bfr_after (
		.din(new_net_13826),
		.dout(new_net_13827)
	);

	bfr new_net_13828_bfr_after (
		.din(new_net_13827),
		.dout(new_net_13828)
	);

	bfr new_net_13829_bfr_after (
		.din(new_net_13828),
		.dout(new_net_13829)
	);

	bfr new_net_13830_bfr_after (
		.din(new_net_13829),
		.dout(new_net_13830)
	);

	bfr new_net_13831_bfr_after (
		.din(new_net_13830),
		.dout(new_net_13831)
	);

	bfr new_net_13832_bfr_after (
		.din(new_net_13831),
		.dout(new_net_13832)
	);

	bfr new_net_13833_bfr_after (
		.din(new_net_13832),
		.dout(new_net_13833)
	);

	bfr new_net_13834_bfr_after (
		.din(new_net_13833),
		.dout(new_net_13834)
	);

	bfr new_net_13835_bfr_after (
		.din(new_net_13834),
		.dout(new_net_13835)
	);

	bfr new_net_13836_bfr_after (
		.din(new_net_13835),
		.dout(new_net_13836)
	);

	bfr new_net_13837_bfr_after (
		.din(new_net_13836),
		.dout(new_net_13837)
	);

	bfr new_net_13838_bfr_after (
		.din(new_net_13837),
		.dout(new_net_13838)
	);

	bfr new_net_13839_bfr_after (
		.din(new_net_13838),
		.dout(new_net_13839)
	);

	bfr new_net_13840_bfr_after (
		.din(new_net_13839),
		.dout(new_net_13840)
	);

	bfr new_net_13841_bfr_after (
		.din(new_net_13840),
		.dout(new_net_13841)
	);

	bfr new_net_13842_bfr_after (
		.din(new_net_13841),
		.dout(new_net_13842)
	);

	bfr new_net_13843_bfr_after (
		.din(new_net_13842),
		.dout(new_net_13843)
	);

	bfr new_net_13844_bfr_after (
		.din(new_net_13843),
		.dout(new_net_13844)
	);

	bfr new_net_13845_bfr_after (
		.din(new_net_13844),
		.dout(new_net_13845)
	);

	bfr new_net_13846_bfr_after (
		.din(new_net_13845),
		.dout(new_net_13846)
	);

	bfr new_net_13847_bfr_after (
		.din(new_net_13846),
		.dout(new_net_13847)
	);

	bfr new_net_13848_bfr_after (
		.din(new_net_13847),
		.dout(new_net_13848)
	);

	bfr new_net_13849_bfr_after (
		.din(new_net_13848),
		.dout(new_net_13849)
	);

	bfr new_net_13850_bfr_after (
		.din(new_net_13849),
		.dout(new_net_13850)
	);

	bfr new_net_13851_bfr_after (
		.din(new_net_13850),
		.dout(new_net_13851)
	);

	bfr new_net_13852_bfr_after (
		.din(new_net_13851),
		.dout(new_net_13852)
	);

	bfr new_net_13853_bfr_after (
		.din(new_net_13852),
		.dout(new_net_13853)
	);

	bfr new_net_13854_bfr_after (
		.din(new_net_13853),
		.dout(new_net_13854)
	);

	bfr new_net_13855_bfr_after (
		.din(new_net_13854),
		.dout(new_net_13855)
	);

	bfr new_net_13856_bfr_after (
		.din(new_net_13855),
		.dout(new_net_13856)
	);

	bfr new_net_13857_bfr_after (
		.din(new_net_13856),
		.dout(new_net_13857)
	);

	bfr new_net_13858_bfr_after (
		.din(new_net_13857),
		.dout(new_net_13858)
	);

	bfr new_net_13859_bfr_after (
		.din(new_net_13858),
		.dout(new_net_13859)
	);

	bfr new_net_13860_bfr_after (
		.din(new_net_13859),
		.dout(new_net_13860)
	);

	bfr new_net_13861_bfr_after (
		.din(new_net_13860),
		.dout(new_net_13861)
	);

	bfr new_net_13862_bfr_after (
		.din(new_net_13861),
		.dout(new_net_13862)
	);

	bfr new_net_13863_bfr_after (
		.din(new_net_13862),
		.dout(new_net_13863)
	);

	bfr new_net_13864_bfr_after (
		.din(new_net_13863),
		.dout(new_net_13864)
	);

	bfr new_net_13865_bfr_after (
		.din(new_net_13864),
		.dout(new_net_13865)
	);

	bfr new_net_13866_bfr_after (
		.din(new_net_13865),
		.dout(new_net_13866)
	);

	bfr new_net_13867_bfr_after (
		.din(new_net_13866),
		.dout(new_net_13867)
	);

	bfr new_net_13868_bfr_after (
		.din(new_net_13867),
		.dout(new_net_13868)
	);

	bfr new_net_13869_bfr_after (
		.din(new_net_13868),
		.dout(new_net_13869)
	);

	bfr new_net_13870_bfr_after (
		.din(new_net_13869),
		.dout(new_net_13870)
	);

	bfr new_net_13871_bfr_after (
		.din(new_net_13870),
		.dout(new_net_13871)
	);

	bfr new_net_13872_bfr_after (
		.din(new_net_13871),
		.dout(new_net_13872)
	);

	bfr new_net_13873_bfr_after (
		.din(new_net_13872),
		.dout(new_net_13873)
	);

	bfr new_net_13874_bfr_after (
		.din(new_net_13873),
		.dout(new_net_13874)
	);

	bfr new_net_13875_bfr_after (
		.din(new_net_13874),
		.dout(new_net_13875)
	);

	bfr new_net_13876_bfr_after (
		.din(new_net_13875),
		.dout(new_net_13876)
	);

	bfr new_net_13877_bfr_after (
		.din(new_net_13876),
		.dout(new_net_13877)
	);

	bfr new_net_13878_bfr_after (
		.din(new_net_13877),
		.dout(new_net_13878)
	);

	bfr new_net_13879_bfr_after (
		.din(new_net_13878),
		.dout(new_net_13879)
	);

	bfr new_net_13880_bfr_after (
		.din(new_net_13879),
		.dout(new_net_13880)
	);

	bfr new_net_13881_bfr_after (
		.din(new_net_13880),
		.dout(new_net_13881)
	);

	bfr new_net_13882_bfr_after (
		.din(new_net_13881),
		.dout(new_net_13882)
	);

	bfr new_net_13883_bfr_after (
		.din(new_net_13882),
		.dout(new_net_13883)
	);

	bfr new_net_13884_bfr_after (
		.din(new_net_13883),
		.dout(new_net_13884)
	);

	bfr new_net_13885_bfr_after (
		.din(new_net_13884),
		.dout(new_net_13885)
	);

	bfr new_net_13886_bfr_after (
		.din(new_net_13885),
		.dout(new_net_13886)
	);

	bfr new_net_13887_bfr_after (
		.din(new_net_13886),
		.dout(new_net_13887)
	);

	bfr new_net_13888_bfr_after (
		.din(new_net_13887),
		.dout(new_net_13888)
	);

	bfr new_net_13889_bfr_after (
		.din(new_net_13888),
		.dout(new_net_13889)
	);

	bfr new_net_13890_bfr_after (
		.din(new_net_13889),
		.dout(new_net_13890)
	);

	bfr new_net_13891_bfr_after (
		.din(new_net_13890),
		.dout(new_net_13891)
	);

	bfr new_net_13892_bfr_after (
		.din(new_net_13891),
		.dout(new_net_13892)
	);

	bfr new_net_13893_bfr_after (
		.din(new_net_13892),
		.dout(new_net_13893)
	);

	bfr new_net_13894_bfr_after (
		.din(new_net_13893),
		.dout(new_net_13894)
	);

	bfr new_net_13895_bfr_after (
		.din(new_net_13894),
		.dout(new_net_13895)
	);

	bfr new_net_13896_bfr_after (
		.din(new_net_13895),
		.dout(new_net_13896)
	);

	bfr new_net_13897_bfr_after (
		.din(new_net_13896),
		.dout(new_net_13897)
	);

	bfr new_net_13898_bfr_after (
		.din(new_net_13897),
		.dout(new_net_13898)
	);

	bfr new_net_13899_bfr_after (
		.din(new_net_13898),
		.dout(new_net_13899)
	);

	bfr new_net_13900_bfr_after (
		.din(new_net_13899),
		.dout(new_net_13900)
	);

	bfr new_net_13901_bfr_after (
		.din(new_net_13900),
		.dout(new_net_13901)
	);

	bfr new_net_13902_bfr_after (
		.din(new_net_13901),
		.dout(new_net_13902)
	);

	bfr new_net_13903_bfr_after (
		.din(new_net_13902),
		.dout(new_net_13903)
	);

	bfr new_net_13904_bfr_after (
		.din(new_net_13903),
		.dout(new_net_13904)
	);

	bfr new_net_13905_bfr_after (
		.din(new_net_13904),
		.dout(new_net_13905)
	);

	spl2 _0767__v_fanout (
		.a(new_net_13905),
		.b(new_net_797),
		.c(new_net_798)
	);

	bfr new_net_13906_bfr_after (
		.din(_1467_),
		.dout(new_net_13906)
	);

	bfr new_net_13907_bfr_after (
		.din(new_net_13906),
		.dout(new_net_13907)
	);

	bfr new_net_13908_bfr_after (
		.din(new_net_13907),
		.dout(new_net_13908)
	);

	bfr new_net_13909_bfr_after (
		.din(new_net_13908),
		.dout(new_net_13909)
	);

	bfr new_net_13910_bfr_after (
		.din(new_net_13909),
		.dout(new_net_13910)
	);

	bfr new_net_13911_bfr_after (
		.din(new_net_13910),
		.dout(new_net_13911)
	);

	bfr new_net_13912_bfr_after (
		.din(new_net_13911),
		.dout(new_net_13912)
	);

	bfr new_net_13913_bfr_after (
		.din(new_net_13912),
		.dout(new_net_13913)
	);

	bfr new_net_13914_bfr_after (
		.din(new_net_13913),
		.dout(new_net_13914)
	);

	bfr new_net_13915_bfr_after (
		.din(new_net_13914),
		.dout(new_net_13915)
	);

	bfr new_net_13916_bfr_after (
		.din(new_net_13915),
		.dout(new_net_13916)
	);

	bfr new_net_13917_bfr_after (
		.din(new_net_13916),
		.dout(new_net_13917)
	);

	bfr new_net_13918_bfr_after (
		.din(new_net_13917),
		.dout(new_net_13918)
	);

	bfr new_net_13919_bfr_after (
		.din(new_net_13918),
		.dout(new_net_13919)
	);

	bfr new_net_13920_bfr_after (
		.din(new_net_13919),
		.dout(new_net_13920)
	);

	bfr new_net_13921_bfr_after (
		.din(new_net_13920),
		.dout(new_net_13921)
	);

	bfr new_net_13922_bfr_after (
		.din(new_net_13921),
		.dout(new_net_13922)
	);

	bfr new_net_13923_bfr_after (
		.din(new_net_13922),
		.dout(new_net_13923)
	);

	bfr new_net_13924_bfr_after (
		.din(new_net_13923),
		.dout(new_net_13924)
	);

	bfr new_net_13925_bfr_after (
		.din(new_net_13924),
		.dout(new_net_13925)
	);

	bfr new_net_13926_bfr_after (
		.din(new_net_13925),
		.dout(new_net_13926)
	);

	bfr new_net_13927_bfr_after (
		.din(new_net_13926),
		.dout(new_net_13927)
	);

	bfr new_net_13928_bfr_after (
		.din(new_net_13927),
		.dout(new_net_13928)
	);

	bfr new_net_13929_bfr_after (
		.din(new_net_13928),
		.dout(new_net_13929)
	);

	bfr new_net_13930_bfr_after (
		.din(new_net_13929),
		.dout(new_net_13930)
	);

	bfr new_net_13931_bfr_after (
		.din(new_net_13930),
		.dout(new_net_13931)
	);

	bfr new_net_13932_bfr_after (
		.din(new_net_13931),
		.dout(new_net_13932)
	);

	bfr new_net_13933_bfr_after (
		.din(new_net_13932),
		.dout(new_net_13933)
	);

	bfr new_net_13934_bfr_after (
		.din(new_net_13933),
		.dout(new_net_13934)
	);

	bfr new_net_13935_bfr_after (
		.din(new_net_13934),
		.dout(new_net_13935)
	);

	bfr new_net_13936_bfr_after (
		.din(new_net_13935),
		.dout(new_net_13936)
	);

	bfr new_net_13937_bfr_after (
		.din(new_net_13936),
		.dout(new_net_13937)
	);

	bfr new_net_13938_bfr_after (
		.din(new_net_13937),
		.dout(new_net_13938)
	);

	bfr new_net_13939_bfr_after (
		.din(new_net_13938),
		.dout(new_net_13939)
	);

	bfr new_net_13940_bfr_after (
		.din(new_net_13939),
		.dout(new_net_13940)
	);

	bfr new_net_13941_bfr_after (
		.din(new_net_13940),
		.dout(new_net_13941)
	);

	bfr new_net_13942_bfr_after (
		.din(new_net_13941),
		.dout(new_net_13942)
	);

	bfr new_net_13943_bfr_after (
		.din(new_net_13942),
		.dout(new_net_13943)
	);

	bfr new_net_13944_bfr_after (
		.din(new_net_13943),
		.dout(new_net_13944)
	);

	bfr new_net_13945_bfr_after (
		.din(new_net_13944),
		.dout(new_net_13945)
	);

	spl2 _1467__v_fanout (
		.a(new_net_13945),
		.b(new_net_980),
		.c(new_net_981)
	);

	bfr new_net_13946_bfr_after (
		.din(_1132_),
		.dout(new_net_13946)
	);

	bfr new_net_13947_bfr_after (
		.din(new_net_13946),
		.dout(new_net_13947)
	);

	bfr new_net_13948_bfr_after (
		.din(new_net_13947),
		.dout(new_net_13948)
	);

	bfr new_net_13949_bfr_after (
		.din(new_net_13948),
		.dout(new_net_13949)
	);

	bfr new_net_13950_bfr_after (
		.din(new_net_13949),
		.dout(new_net_13950)
	);

	bfr new_net_13951_bfr_after (
		.din(new_net_13950),
		.dout(new_net_13951)
	);

	bfr new_net_13952_bfr_after (
		.din(new_net_13951),
		.dout(new_net_13952)
	);

	bfr new_net_13953_bfr_after (
		.din(new_net_13952),
		.dout(new_net_13953)
	);

	bfr new_net_13954_bfr_after (
		.din(new_net_13953),
		.dout(new_net_13954)
	);

	bfr new_net_13955_bfr_after (
		.din(new_net_13954),
		.dout(new_net_13955)
	);

	bfr new_net_13956_bfr_after (
		.din(new_net_13955),
		.dout(new_net_13956)
	);

	bfr new_net_13957_bfr_after (
		.din(new_net_13956),
		.dout(new_net_13957)
	);

	bfr new_net_13958_bfr_after (
		.din(new_net_13957),
		.dout(new_net_13958)
	);

	bfr new_net_13959_bfr_after (
		.din(new_net_13958),
		.dout(new_net_13959)
	);

	bfr new_net_13960_bfr_after (
		.din(new_net_13959),
		.dout(new_net_13960)
	);

	bfr new_net_13961_bfr_after (
		.din(new_net_13960),
		.dout(new_net_13961)
	);

	bfr new_net_13962_bfr_after (
		.din(new_net_13961),
		.dout(new_net_13962)
	);

	bfr new_net_13963_bfr_after (
		.din(new_net_13962),
		.dout(new_net_13963)
	);

	bfr new_net_13964_bfr_after (
		.din(new_net_13963),
		.dout(new_net_13964)
	);

	bfr new_net_13965_bfr_after (
		.din(new_net_13964),
		.dout(new_net_13965)
	);

	bfr new_net_13966_bfr_after (
		.din(new_net_13965),
		.dout(new_net_13966)
	);

	bfr new_net_13967_bfr_after (
		.din(new_net_13966),
		.dout(new_net_13967)
	);

	bfr new_net_13968_bfr_after (
		.din(new_net_13967),
		.dout(new_net_13968)
	);

	bfr new_net_13969_bfr_after (
		.din(new_net_13968),
		.dout(new_net_13969)
	);

	bfr new_net_13970_bfr_after (
		.din(new_net_13969),
		.dout(new_net_13970)
	);

	bfr new_net_13971_bfr_after (
		.din(new_net_13970),
		.dout(new_net_13971)
	);

	bfr new_net_13972_bfr_after (
		.din(new_net_13971),
		.dout(new_net_13972)
	);

	bfr new_net_13973_bfr_after (
		.din(new_net_13972),
		.dout(new_net_13973)
	);

	bfr new_net_13974_bfr_after (
		.din(new_net_13973),
		.dout(new_net_13974)
	);

	bfr new_net_13975_bfr_after (
		.din(new_net_13974),
		.dout(new_net_13975)
	);

	bfr new_net_13976_bfr_after (
		.din(new_net_13975),
		.dout(new_net_13976)
	);

	bfr new_net_13977_bfr_after (
		.din(new_net_13976),
		.dout(new_net_13977)
	);

	bfr new_net_13978_bfr_after (
		.din(new_net_13977),
		.dout(new_net_13978)
	);

	bfr new_net_13979_bfr_after (
		.din(new_net_13978),
		.dout(new_net_13979)
	);

	bfr new_net_13980_bfr_after (
		.din(new_net_13979),
		.dout(new_net_13980)
	);

	bfr new_net_13981_bfr_after (
		.din(new_net_13980),
		.dout(new_net_13981)
	);

	bfr new_net_13982_bfr_after (
		.din(new_net_13981),
		.dout(new_net_13982)
	);

	bfr new_net_13983_bfr_after (
		.din(new_net_13982),
		.dout(new_net_13983)
	);

	bfr new_net_13984_bfr_after (
		.din(new_net_13983),
		.dout(new_net_13984)
	);

	bfr new_net_13985_bfr_after (
		.din(new_net_13984),
		.dout(new_net_13985)
	);

	bfr new_net_13986_bfr_after (
		.din(new_net_13985),
		.dout(new_net_13986)
	);

	bfr new_net_13987_bfr_after (
		.din(new_net_13986),
		.dout(new_net_13987)
	);

	bfr new_net_13988_bfr_after (
		.din(new_net_13987),
		.dout(new_net_13988)
	);

	bfr new_net_13989_bfr_after (
		.din(new_net_13988),
		.dout(new_net_13989)
	);

	bfr new_net_13990_bfr_after (
		.din(new_net_13989),
		.dout(new_net_13990)
	);

	bfr new_net_13991_bfr_after (
		.din(new_net_13990),
		.dout(new_net_13991)
	);

	bfr new_net_13992_bfr_after (
		.din(new_net_13991),
		.dout(new_net_13992)
	);

	bfr new_net_13993_bfr_after (
		.din(new_net_13992),
		.dout(new_net_13993)
	);

	spl2 _1132__v_fanout (
		.a(new_net_13993),
		.b(new_net_293),
		.c(new_net_294)
	);

	bfr new_net_13994_bfr_after (
		.din(_1817_),
		.dout(new_net_13994)
	);

	bfr new_net_13995_bfr_after (
		.din(new_net_13994),
		.dout(new_net_13995)
	);

	bfr new_net_13996_bfr_after (
		.din(new_net_13995),
		.dout(new_net_13996)
	);

	bfr new_net_13997_bfr_after (
		.din(new_net_13996),
		.dout(new_net_13997)
	);

	bfr new_net_13998_bfr_after (
		.din(new_net_13997),
		.dout(new_net_13998)
	);

	bfr new_net_13999_bfr_after (
		.din(new_net_13998),
		.dout(new_net_13999)
	);

	bfr new_net_14000_bfr_after (
		.din(new_net_13999),
		.dout(new_net_14000)
	);

	bfr new_net_14001_bfr_after (
		.din(new_net_14000),
		.dout(new_net_14001)
	);

	bfr new_net_14002_bfr_after (
		.din(new_net_14001),
		.dout(new_net_14002)
	);

	bfr new_net_14003_bfr_after (
		.din(new_net_14002),
		.dout(new_net_14003)
	);

	bfr new_net_14004_bfr_after (
		.din(new_net_14003),
		.dout(new_net_14004)
	);

	bfr new_net_14005_bfr_after (
		.din(new_net_14004),
		.dout(new_net_14005)
	);

	bfr new_net_14006_bfr_after (
		.din(new_net_14005),
		.dout(new_net_14006)
	);

	bfr new_net_14007_bfr_after (
		.din(new_net_14006),
		.dout(new_net_14007)
	);

	bfr new_net_14008_bfr_after (
		.din(new_net_14007),
		.dout(new_net_14008)
	);

	bfr new_net_14009_bfr_after (
		.din(new_net_14008),
		.dout(new_net_14009)
	);

	bfr new_net_14010_bfr_after (
		.din(new_net_14009),
		.dout(new_net_14010)
	);

	bfr new_net_14011_bfr_after (
		.din(new_net_14010),
		.dout(new_net_14011)
	);

	bfr new_net_14012_bfr_after (
		.din(new_net_14011),
		.dout(new_net_14012)
	);

	bfr new_net_14013_bfr_after (
		.din(new_net_14012),
		.dout(new_net_14013)
	);

	bfr new_net_14014_bfr_after (
		.din(new_net_14013),
		.dout(new_net_14014)
	);

	bfr new_net_14015_bfr_after (
		.din(new_net_14014),
		.dout(new_net_14015)
	);

	bfr new_net_14016_bfr_after (
		.din(new_net_14015),
		.dout(new_net_14016)
	);

	bfr new_net_14017_bfr_after (
		.din(new_net_14016),
		.dout(new_net_14017)
	);

	bfr new_net_14018_bfr_after (
		.din(new_net_14017),
		.dout(new_net_14018)
	);

	bfr new_net_14019_bfr_after (
		.din(new_net_14018),
		.dout(new_net_14019)
	);

	bfr new_net_14020_bfr_after (
		.din(new_net_14019),
		.dout(new_net_14020)
	);

	bfr new_net_14021_bfr_after (
		.din(new_net_14020),
		.dout(new_net_14021)
	);

	bfr new_net_14022_bfr_after (
		.din(new_net_14021),
		.dout(new_net_14022)
	);

	bfr new_net_14023_bfr_after (
		.din(new_net_14022),
		.dout(new_net_14023)
	);

	bfr new_net_14024_bfr_after (
		.din(new_net_14023),
		.dout(new_net_14024)
	);

	bfr new_net_14025_bfr_after (
		.din(new_net_14024),
		.dout(new_net_14025)
	);

	bfr new_net_14026_bfr_after (
		.din(new_net_14025),
		.dout(new_net_14026)
	);

	bfr new_net_14027_bfr_after (
		.din(new_net_14026),
		.dout(new_net_14027)
	);

	bfr new_net_14028_bfr_after (
		.din(new_net_14027),
		.dout(new_net_14028)
	);

	bfr new_net_14029_bfr_after (
		.din(new_net_14028),
		.dout(new_net_14029)
	);

	bfr new_net_14030_bfr_after (
		.din(new_net_14029),
		.dout(new_net_14030)
	);

	bfr new_net_14031_bfr_after (
		.din(new_net_14030),
		.dout(new_net_14031)
	);

	bfr new_net_14032_bfr_after (
		.din(new_net_14031),
		.dout(new_net_14032)
	);

	bfr new_net_14033_bfr_after (
		.din(new_net_14032),
		.dout(new_net_14033)
	);

	bfr new_net_14034_bfr_after (
		.din(new_net_14033),
		.dout(new_net_14034)
	);

	bfr new_net_14035_bfr_after (
		.din(new_net_14034),
		.dout(new_net_14035)
	);

	bfr new_net_14036_bfr_after (
		.din(new_net_14035),
		.dout(new_net_14036)
	);

	bfr new_net_14037_bfr_after (
		.din(new_net_14036),
		.dout(new_net_14037)
	);

	bfr new_net_14038_bfr_after (
		.din(new_net_14037),
		.dout(new_net_14038)
	);

	bfr new_net_14039_bfr_after (
		.din(new_net_14038),
		.dout(new_net_14039)
	);

	bfr new_net_14040_bfr_after (
		.din(new_net_14039),
		.dout(new_net_14040)
	);

	bfr new_net_14041_bfr_after (
		.din(new_net_14040),
		.dout(new_net_14041)
	);

	bfr new_net_14042_bfr_after (
		.din(new_net_14041),
		.dout(new_net_14042)
	);

	bfr new_net_14043_bfr_after (
		.din(new_net_14042),
		.dout(new_net_14043)
	);

	bfr new_net_14044_bfr_after (
		.din(new_net_14043),
		.dout(new_net_14044)
	);

	bfr new_net_14045_bfr_after (
		.din(new_net_14044),
		.dout(new_net_14045)
	);

	bfr new_net_14046_bfr_after (
		.din(new_net_14045),
		.dout(new_net_14046)
	);

	bfr new_net_14047_bfr_after (
		.din(new_net_14046),
		.dout(new_net_14047)
	);

	bfr new_net_14048_bfr_after (
		.din(new_net_14047),
		.dout(new_net_14048)
	);

	bfr new_net_14049_bfr_after (
		.din(new_net_14048),
		.dout(new_net_14049)
	);

	spl2 _1817__v_fanout (
		.a(new_net_14049),
		.b(new_net_1326),
		.c(new_net_1327)
	);

	bfr new_net_14050_bfr_after (
		.din(_1082_),
		.dout(new_net_14050)
	);

	bfr new_net_14051_bfr_after (
		.din(new_net_14050),
		.dout(new_net_14051)
	);

	bfr new_net_14052_bfr_after (
		.din(new_net_14051),
		.dout(new_net_14052)
	);

	bfr new_net_14053_bfr_after (
		.din(new_net_14052),
		.dout(new_net_14053)
	);

	bfr new_net_14054_bfr_after (
		.din(new_net_14053),
		.dout(new_net_14054)
	);

	bfr new_net_14055_bfr_after (
		.din(new_net_14054),
		.dout(new_net_14055)
	);

	bfr new_net_14056_bfr_after (
		.din(new_net_14055),
		.dout(new_net_14056)
	);

	bfr new_net_14057_bfr_after (
		.din(new_net_14056),
		.dout(new_net_14057)
	);

	spl2 _1082__v_fanout (
		.a(new_net_14057),
		.b(new_net_1990),
		.c(new_net_1991)
	);

	bfr new_net_14058_bfr_after (
		.din(_1213_),
		.dout(new_net_14058)
	);

	bfr new_net_14059_bfr_after (
		.din(new_net_14058),
		.dout(new_net_14059)
	);

	bfr new_net_14060_bfr_after (
		.din(new_net_14059),
		.dout(new_net_14060)
	);

	bfr new_net_14061_bfr_after (
		.din(new_net_14060),
		.dout(new_net_14061)
	);

	bfr new_net_14062_bfr_after (
		.din(new_net_14061),
		.dout(new_net_14062)
	);

	bfr new_net_14063_bfr_after (
		.din(new_net_14062),
		.dout(new_net_14063)
	);

	bfr new_net_14064_bfr_after (
		.din(new_net_14063),
		.dout(new_net_14064)
	);

	bfr new_net_14065_bfr_after (
		.din(new_net_14064),
		.dout(new_net_14065)
	);

	bfr new_net_14066_bfr_after (
		.din(new_net_14065),
		.dout(new_net_14066)
	);

	bfr new_net_14067_bfr_after (
		.din(new_net_14066),
		.dout(new_net_14067)
	);

	bfr new_net_14068_bfr_after (
		.din(new_net_14067),
		.dout(new_net_14068)
	);

	bfr new_net_14069_bfr_after (
		.din(new_net_14068),
		.dout(new_net_14069)
	);

	bfr new_net_14070_bfr_after (
		.din(new_net_14069),
		.dout(new_net_14070)
	);

	bfr new_net_14071_bfr_after (
		.din(new_net_14070),
		.dout(new_net_14071)
	);

	bfr new_net_14072_bfr_after (
		.din(new_net_14071),
		.dout(new_net_14072)
	);

	bfr new_net_14073_bfr_after (
		.din(new_net_14072),
		.dout(new_net_14073)
	);

	bfr new_net_14074_bfr_after (
		.din(new_net_14073),
		.dout(new_net_14074)
	);

	bfr new_net_14075_bfr_after (
		.din(new_net_14074),
		.dout(new_net_14075)
	);

	bfr new_net_14076_bfr_after (
		.din(new_net_14075),
		.dout(new_net_14076)
	);

	bfr new_net_14077_bfr_after (
		.din(new_net_14076),
		.dout(new_net_14077)
	);

	bfr new_net_14078_bfr_after (
		.din(new_net_14077),
		.dout(new_net_14078)
	);

	bfr new_net_14079_bfr_after (
		.din(new_net_14078),
		.dout(new_net_14079)
	);

	bfr new_net_14080_bfr_after (
		.din(new_net_14079),
		.dout(new_net_14080)
	);

	bfr new_net_14081_bfr_after (
		.din(new_net_14080),
		.dout(new_net_14081)
	);

	bfr new_net_14082_bfr_after (
		.din(new_net_14081),
		.dout(new_net_14082)
	);

	bfr new_net_14083_bfr_after (
		.din(new_net_14082),
		.dout(new_net_14083)
	);

	bfr new_net_14084_bfr_after (
		.din(new_net_14083),
		.dout(new_net_14084)
	);

	bfr new_net_14085_bfr_after (
		.din(new_net_14084),
		.dout(new_net_14085)
	);

	bfr new_net_14086_bfr_after (
		.din(new_net_14085),
		.dout(new_net_14086)
	);

	bfr new_net_14087_bfr_after (
		.din(new_net_14086),
		.dout(new_net_14087)
	);

	bfr new_net_14088_bfr_after (
		.din(new_net_14087),
		.dout(new_net_14088)
	);

	bfr new_net_14089_bfr_after (
		.din(new_net_14088),
		.dout(new_net_14089)
	);

	spl2 _1213__v_fanout (
		.a(new_net_14089),
		.b(new_net_896),
		.c(new_net_897)
	);

	bfr new_net_14090_bfr_after (
		.din(_1684_),
		.dout(new_net_14090)
	);

	bfr new_net_14091_bfr_after (
		.din(new_net_14090),
		.dout(new_net_14091)
	);

	bfr new_net_14092_bfr_after (
		.din(new_net_14091),
		.dout(new_net_14092)
	);

	bfr new_net_14093_bfr_after (
		.din(new_net_14092),
		.dout(new_net_14093)
	);

	bfr new_net_14094_bfr_after (
		.din(new_net_14093),
		.dout(new_net_14094)
	);

	bfr new_net_14095_bfr_after (
		.din(new_net_14094),
		.dout(new_net_14095)
	);

	bfr new_net_14096_bfr_after (
		.din(new_net_14095),
		.dout(new_net_14096)
	);

	bfr new_net_14097_bfr_after (
		.din(new_net_14096),
		.dout(new_net_14097)
	);

	bfr new_net_14098_bfr_after (
		.din(new_net_14097),
		.dout(new_net_14098)
	);

	bfr new_net_14099_bfr_after (
		.din(new_net_14098),
		.dout(new_net_14099)
	);

	bfr new_net_14100_bfr_after (
		.din(new_net_14099),
		.dout(new_net_14100)
	);

	bfr new_net_14101_bfr_after (
		.din(new_net_14100),
		.dout(new_net_14101)
	);

	bfr new_net_14102_bfr_after (
		.din(new_net_14101),
		.dout(new_net_14102)
	);

	bfr new_net_14103_bfr_after (
		.din(new_net_14102),
		.dout(new_net_14103)
	);

	bfr new_net_14104_bfr_after (
		.din(new_net_14103),
		.dout(new_net_14104)
	);

	bfr new_net_14105_bfr_after (
		.din(new_net_14104),
		.dout(new_net_14105)
	);

	bfr new_net_14106_bfr_after (
		.din(new_net_14105),
		.dout(new_net_14106)
	);

	bfr new_net_14107_bfr_after (
		.din(new_net_14106),
		.dout(new_net_14107)
	);

	bfr new_net_14108_bfr_after (
		.din(new_net_14107),
		.dout(new_net_14108)
	);

	bfr new_net_14109_bfr_after (
		.din(new_net_14108),
		.dout(new_net_14109)
	);

	bfr new_net_14110_bfr_after (
		.din(new_net_14109),
		.dout(new_net_14110)
	);

	bfr new_net_14111_bfr_after (
		.din(new_net_14110),
		.dout(new_net_14111)
	);

	bfr new_net_14112_bfr_after (
		.din(new_net_14111),
		.dout(new_net_14112)
	);

	bfr new_net_14113_bfr_after (
		.din(new_net_14112),
		.dout(new_net_14113)
	);

	bfr new_net_14114_bfr_after (
		.din(new_net_14113),
		.dout(new_net_14114)
	);

	bfr new_net_14115_bfr_after (
		.din(new_net_14114),
		.dout(new_net_14115)
	);

	bfr new_net_14116_bfr_after (
		.din(new_net_14115),
		.dout(new_net_14116)
	);

	bfr new_net_14117_bfr_after (
		.din(new_net_14116),
		.dout(new_net_14117)
	);

	bfr new_net_14118_bfr_after (
		.din(new_net_14117),
		.dout(new_net_14118)
	);

	bfr new_net_14119_bfr_after (
		.din(new_net_14118),
		.dout(new_net_14119)
	);

	bfr new_net_14120_bfr_after (
		.din(new_net_14119),
		.dout(new_net_14120)
	);

	bfr new_net_14121_bfr_after (
		.din(new_net_14120),
		.dout(new_net_14121)
	);

	bfr new_net_14122_bfr_after (
		.din(new_net_14121),
		.dout(new_net_14122)
	);

	bfr new_net_14123_bfr_after (
		.din(new_net_14122),
		.dout(new_net_14123)
	);

	bfr new_net_14124_bfr_after (
		.din(new_net_14123),
		.dout(new_net_14124)
	);

	bfr new_net_14125_bfr_after (
		.din(new_net_14124),
		.dout(new_net_14125)
	);

	bfr new_net_14126_bfr_after (
		.din(new_net_14125),
		.dout(new_net_14126)
	);

	bfr new_net_14127_bfr_after (
		.din(new_net_14126),
		.dout(new_net_14127)
	);

	bfr new_net_14128_bfr_after (
		.din(new_net_14127),
		.dout(new_net_14128)
	);

	bfr new_net_14129_bfr_after (
		.din(new_net_14128),
		.dout(new_net_14129)
	);

	bfr new_net_14130_bfr_after (
		.din(new_net_14129),
		.dout(new_net_14130)
	);

	bfr new_net_14131_bfr_after (
		.din(new_net_14130),
		.dout(new_net_14131)
	);

	bfr new_net_14132_bfr_after (
		.din(new_net_14131),
		.dout(new_net_14132)
	);

	bfr new_net_14133_bfr_after (
		.din(new_net_14132),
		.dout(new_net_14133)
	);

	bfr new_net_14134_bfr_after (
		.din(new_net_14133),
		.dout(new_net_14134)
	);

	bfr new_net_14135_bfr_after (
		.din(new_net_14134),
		.dout(new_net_14135)
	);

	bfr new_net_14136_bfr_after (
		.din(new_net_14135),
		.dout(new_net_14136)
	);

	bfr new_net_14137_bfr_after (
		.din(new_net_14136),
		.dout(new_net_14137)
	);

	bfr new_net_14138_bfr_after (
		.din(new_net_14137),
		.dout(new_net_14138)
	);

	bfr new_net_14139_bfr_after (
		.din(new_net_14138),
		.dout(new_net_14139)
	);

	bfr new_net_14140_bfr_after (
		.din(new_net_14139),
		.dout(new_net_14140)
	);

	bfr new_net_14141_bfr_after (
		.din(new_net_14140),
		.dout(new_net_14141)
	);

	bfr new_net_14142_bfr_after (
		.din(new_net_14141),
		.dout(new_net_14142)
	);

	bfr new_net_14143_bfr_after (
		.din(new_net_14142),
		.dout(new_net_14143)
	);

	bfr new_net_14144_bfr_after (
		.din(new_net_14143),
		.dout(new_net_14144)
	);

	bfr new_net_14145_bfr_after (
		.din(new_net_14144),
		.dout(new_net_14145)
	);

	bfr new_net_14146_bfr_after (
		.din(new_net_14145),
		.dout(new_net_14146)
	);

	bfr new_net_14147_bfr_after (
		.din(new_net_14146),
		.dout(new_net_14147)
	);

	bfr new_net_14148_bfr_after (
		.din(new_net_14147),
		.dout(new_net_14148)
	);

	bfr new_net_14149_bfr_after (
		.din(new_net_14148),
		.dout(new_net_14149)
	);

	bfr new_net_14150_bfr_after (
		.din(new_net_14149),
		.dout(new_net_14150)
	);

	bfr new_net_14151_bfr_after (
		.din(new_net_14150),
		.dout(new_net_14151)
	);

	bfr new_net_14152_bfr_after (
		.din(new_net_14151),
		.dout(new_net_14152)
	);

	bfr new_net_14153_bfr_after (
		.din(new_net_14152),
		.dout(new_net_14153)
	);

	bfr new_net_14154_bfr_after (
		.din(new_net_14153),
		.dout(new_net_14154)
	);

	bfr new_net_14155_bfr_after (
		.din(new_net_14154),
		.dout(new_net_14155)
	);

	bfr new_net_14156_bfr_after (
		.din(new_net_14155),
		.dout(new_net_14156)
	);

	bfr new_net_14157_bfr_after (
		.din(new_net_14156),
		.dout(new_net_14157)
	);

	bfr new_net_14158_bfr_after (
		.din(new_net_14157),
		.dout(new_net_14158)
	);

	bfr new_net_14159_bfr_after (
		.din(new_net_14158),
		.dout(new_net_14159)
	);

	bfr new_net_14160_bfr_after (
		.din(new_net_14159),
		.dout(new_net_14160)
	);

	bfr new_net_14161_bfr_after (
		.din(new_net_14160),
		.dout(new_net_14161)
	);

	bfr new_net_14162_bfr_after (
		.din(new_net_14161),
		.dout(new_net_14162)
	);

	bfr new_net_14163_bfr_after (
		.din(new_net_14162),
		.dout(new_net_14163)
	);

	bfr new_net_14164_bfr_after (
		.din(new_net_14163),
		.dout(new_net_14164)
	);

	bfr new_net_14165_bfr_after (
		.din(new_net_14164),
		.dout(new_net_14165)
	);

	bfr new_net_14166_bfr_after (
		.din(new_net_14165),
		.dout(new_net_14166)
	);

	bfr new_net_14167_bfr_after (
		.din(new_net_14166),
		.dout(new_net_14167)
	);

	bfr new_net_14168_bfr_after (
		.din(new_net_14167),
		.dout(new_net_14168)
	);

	bfr new_net_14169_bfr_after (
		.din(new_net_14168),
		.dout(new_net_14169)
	);

	bfr new_net_14170_bfr_after (
		.din(new_net_14169),
		.dout(new_net_14170)
	);

	bfr new_net_14171_bfr_after (
		.din(new_net_14170),
		.dout(new_net_14171)
	);

	bfr new_net_14172_bfr_after (
		.din(new_net_14171),
		.dout(new_net_14172)
	);

	bfr new_net_14173_bfr_after (
		.din(new_net_14172),
		.dout(new_net_14173)
	);

	bfr new_net_14174_bfr_after (
		.din(new_net_14173),
		.dout(new_net_14174)
	);

	bfr new_net_14175_bfr_after (
		.din(new_net_14174),
		.dout(new_net_14175)
	);

	bfr new_net_14176_bfr_after (
		.din(new_net_14175),
		.dout(new_net_14176)
	);

	bfr new_net_14177_bfr_after (
		.din(new_net_14176),
		.dout(new_net_14177)
	);

	spl2 _1684__v_fanout (
		.a(new_net_14177),
		.b(new_net_2827),
		.c(new_net_2828)
	);

	bfr new_net_14178_bfr_after (
		.din(_1125_),
		.dout(new_net_14178)
	);

	bfr new_net_14179_bfr_after (
		.din(new_net_14178),
		.dout(new_net_14179)
	);

	bfr new_net_14180_bfr_after (
		.din(new_net_14179),
		.dout(new_net_14180)
	);

	bfr new_net_14181_bfr_after (
		.din(new_net_14180),
		.dout(new_net_14181)
	);

	bfr new_net_14182_bfr_after (
		.din(new_net_14181),
		.dout(new_net_14182)
	);

	bfr new_net_14183_bfr_after (
		.din(new_net_14182),
		.dout(new_net_14183)
	);

	bfr new_net_14184_bfr_after (
		.din(new_net_14183),
		.dout(new_net_14184)
	);

	bfr new_net_14185_bfr_after (
		.din(new_net_14184),
		.dout(new_net_14185)
	);

	bfr new_net_14186_bfr_after (
		.din(new_net_14185),
		.dout(new_net_14186)
	);

	bfr new_net_14187_bfr_after (
		.din(new_net_14186),
		.dout(new_net_14187)
	);

	bfr new_net_14188_bfr_after (
		.din(new_net_14187),
		.dout(new_net_14188)
	);

	bfr new_net_14189_bfr_after (
		.din(new_net_14188),
		.dout(new_net_14189)
	);

	bfr new_net_14190_bfr_after (
		.din(new_net_14189),
		.dout(new_net_14190)
	);

	bfr new_net_14191_bfr_after (
		.din(new_net_14190),
		.dout(new_net_14191)
	);

	bfr new_net_14192_bfr_after (
		.din(new_net_14191),
		.dout(new_net_14192)
	);

	bfr new_net_14193_bfr_after (
		.din(new_net_14192),
		.dout(new_net_14193)
	);

	bfr new_net_14194_bfr_after (
		.din(new_net_14193),
		.dout(new_net_14194)
	);

	bfr new_net_14195_bfr_after (
		.din(new_net_14194),
		.dout(new_net_14195)
	);

	bfr new_net_14196_bfr_after (
		.din(new_net_14195),
		.dout(new_net_14196)
	);

	bfr new_net_14197_bfr_after (
		.din(new_net_14196),
		.dout(new_net_14197)
	);

	bfr new_net_14198_bfr_after (
		.din(new_net_14197),
		.dout(new_net_14198)
	);

	bfr new_net_14199_bfr_after (
		.din(new_net_14198),
		.dout(new_net_14199)
	);

	bfr new_net_14200_bfr_after (
		.din(new_net_14199),
		.dout(new_net_14200)
	);

	bfr new_net_14201_bfr_after (
		.din(new_net_14200),
		.dout(new_net_14201)
	);

	bfr new_net_14202_bfr_after (
		.din(new_net_14201),
		.dout(new_net_14202)
	);

	bfr new_net_14203_bfr_after (
		.din(new_net_14202),
		.dout(new_net_14203)
	);

	bfr new_net_14204_bfr_after (
		.din(new_net_14203),
		.dout(new_net_14204)
	);

	bfr new_net_14205_bfr_after (
		.din(new_net_14204),
		.dout(new_net_14205)
	);

	bfr new_net_14206_bfr_after (
		.din(new_net_14205),
		.dout(new_net_14206)
	);

	bfr new_net_14207_bfr_after (
		.din(new_net_14206),
		.dout(new_net_14207)
	);

	bfr new_net_14208_bfr_after (
		.din(new_net_14207),
		.dout(new_net_14208)
	);

	bfr new_net_14209_bfr_after (
		.din(new_net_14208),
		.dout(new_net_14209)
	);

	bfr new_net_14210_bfr_after (
		.din(new_net_14209),
		.dout(new_net_14210)
	);

	bfr new_net_14211_bfr_after (
		.din(new_net_14210),
		.dout(new_net_14211)
	);

	bfr new_net_14212_bfr_after (
		.din(new_net_14211),
		.dout(new_net_14212)
	);

	bfr new_net_14213_bfr_after (
		.din(new_net_14212),
		.dout(new_net_14213)
	);

	bfr new_net_14214_bfr_after (
		.din(new_net_14213),
		.dout(new_net_14214)
	);

	bfr new_net_14215_bfr_after (
		.din(new_net_14214),
		.dout(new_net_14215)
	);

	bfr new_net_14216_bfr_after (
		.din(new_net_14215),
		.dout(new_net_14216)
	);

	bfr new_net_14217_bfr_after (
		.din(new_net_14216),
		.dout(new_net_14217)
	);

	bfr new_net_14218_bfr_after (
		.din(new_net_14217),
		.dout(new_net_14218)
	);

	bfr new_net_14219_bfr_after (
		.din(new_net_14218),
		.dout(new_net_14219)
	);

	bfr new_net_14220_bfr_after (
		.din(new_net_14219),
		.dout(new_net_14220)
	);

	bfr new_net_14221_bfr_after (
		.din(new_net_14220),
		.dout(new_net_14221)
	);

	bfr new_net_14222_bfr_after (
		.din(new_net_14221),
		.dout(new_net_14222)
	);

	bfr new_net_14223_bfr_after (
		.din(new_net_14222),
		.dout(new_net_14223)
	);

	bfr new_net_14224_bfr_after (
		.din(new_net_14223),
		.dout(new_net_14224)
	);

	bfr new_net_14225_bfr_after (
		.din(new_net_14224),
		.dout(new_net_14225)
	);

	bfr new_net_14226_bfr_after (
		.din(new_net_14225),
		.dout(new_net_14226)
	);

	bfr new_net_14227_bfr_after (
		.din(new_net_14226),
		.dout(new_net_14227)
	);

	bfr new_net_14228_bfr_after (
		.din(new_net_14227),
		.dout(new_net_14228)
	);

	bfr new_net_14229_bfr_after (
		.din(new_net_14228),
		.dout(new_net_14229)
	);

	bfr new_net_14230_bfr_after (
		.din(new_net_14229),
		.dout(new_net_14230)
	);

	bfr new_net_14231_bfr_after (
		.din(new_net_14230),
		.dout(new_net_14231)
	);

	bfr new_net_14232_bfr_after (
		.din(new_net_14231),
		.dout(new_net_14232)
	);

	bfr new_net_14233_bfr_after (
		.din(new_net_14232),
		.dout(new_net_14233)
	);

	spl2 _1125__v_fanout (
		.a(new_net_14233),
		.b(new_net_2146),
		.c(new_net_2147)
	);

	bfr new_net_14234_bfr_after (
		.din(_0439_),
		.dout(new_net_14234)
	);

	bfr new_net_14235_bfr_after (
		.din(new_net_14234),
		.dout(new_net_14235)
	);

	bfr new_net_14236_bfr_after (
		.din(new_net_14235),
		.dout(new_net_14236)
	);

	bfr new_net_14237_bfr_after (
		.din(new_net_14236),
		.dout(new_net_14237)
	);

	bfr new_net_14238_bfr_after (
		.din(new_net_14237),
		.dout(new_net_14238)
	);

	bfr new_net_14239_bfr_after (
		.din(new_net_14238),
		.dout(new_net_14239)
	);

	bfr new_net_14240_bfr_after (
		.din(new_net_14239),
		.dout(new_net_14240)
	);

	bfr new_net_14241_bfr_after (
		.din(new_net_14240),
		.dout(new_net_14241)
	);

	bfr new_net_14242_bfr_after (
		.din(new_net_14241),
		.dout(new_net_14242)
	);

	bfr new_net_14243_bfr_after (
		.din(new_net_14242),
		.dout(new_net_14243)
	);

	bfr new_net_14244_bfr_after (
		.din(new_net_14243),
		.dout(new_net_14244)
	);

	bfr new_net_14245_bfr_after (
		.din(new_net_14244),
		.dout(new_net_14245)
	);

	bfr new_net_14246_bfr_after (
		.din(new_net_14245),
		.dout(new_net_14246)
	);

	bfr new_net_14247_bfr_after (
		.din(new_net_14246),
		.dout(new_net_14247)
	);

	bfr new_net_14248_bfr_after (
		.din(new_net_14247),
		.dout(new_net_14248)
	);

	bfr new_net_14249_bfr_after (
		.din(new_net_14248),
		.dout(new_net_14249)
	);

	bfr new_net_14250_bfr_after (
		.din(new_net_14249),
		.dout(new_net_14250)
	);

	bfr new_net_14251_bfr_after (
		.din(new_net_14250),
		.dout(new_net_14251)
	);

	bfr new_net_14252_bfr_after (
		.din(new_net_14251),
		.dout(new_net_14252)
	);

	bfr new_net_14253_bfr_after (
		.din(new_net_14252),
		.dout(new_net_14253)
	);

	bfr new_net_14254_bfr_after (
		.din(new_net_14253),
		.dout(new_net_14254)
	);

	bfr new_net_14255_bfr_after (
		.din(new_net_14254),
		.dout(new_net_14255)
	);

	bfr new_net_14256_bfr_after (
		.din(new_net_14255),
		.dout(new_net_14256)
	);

	bfr new_net_14257_bfr_after (
		.din(new_net_14256),
		.dout(new_net_14257)
	);

	bfr new_net_14258_bfr_after (
		.din(new_net_14257),
		.dout(new_net_14258)
	);

	bfr new_net_14259_bfr_after (
		.din(new_net_14258),
		.dout(new_net_14259)
	);

	bfr new_net_14260_bfr_after (
		.din(new_net_14259),
		.dout(new_net_14260)
	);

	bfr new_net_14261_bfr_after (
		.din(new_net_14260),
		.dout(new_net_14261)
	);

	bfr new_net_14262_bfr_after (
		.din(new_net_14261),
		.dout(new_net_14262)
	);

	bfr new_net_14263_bfr_after (
		.din(new_net_14262),
		.dout(new_net_14263)
	);

	bfr new_net_14264_bfr_after (
		.din(new_net_14263),
		.dout(new_net_14264)
	);

	bfr new_net_14265_bfr_after (
		.din(new_net_14264),
		.dout(new_net_14265)
	);

	bfr new_net_14266_bfr_after (
		.din(new_net_14265),
		.dout(new_net_14266)
	);

	bfr new_net_14267_bfr_after (
		.din(new_net_14266),
		.dout(new_net_14267)
	);

	bfr new_net_14268_bfr_after (
		.din(new_net_14267),
		.dout(new_net_14268)
	);

	bfr new_net_14269_bfr_after (
		.din(new_net_14268),
		.dout(new_net_14269)
	);

	bfr new_net_14270_bfr_after (
		.din(new_net_14269),
		.dout(new_net_14270)
	);

	bfr new_net_14271_bfr_after (
		.din(new_net_14270),
		.dout(new_net_14271)
	);

	bfr new_net_14272_bfr_after (
		.din(new_net_14271),
		.dout(new_net_14272)
	);

	bfr new_net_14273_bfr_after (
		.din(new_net_14272),
		.dout(new_net_14273)
	);

	bfr new_net_14274_bfr_after (
		.din(new_net_14273),
		.dout(new_net_14274)
	);

	bfr new_net_14275_bfr_after (
		.din(new_net_14274),
		.dout(new_net_14275)
	);

	bfr new_net_14276_bfr_after (
		.din(new_net_14275),
		.dout(new_net_14276)
	);

	bfr new_net_14277_bfr_after (
		.din(new_net_14276),
		.dout(new_net_14277)
	);

	bfr new_net_14278_bfr_after (
		.din(new_net_14277),
		.dout(new_net_14278)
	);

	bfr new_net_14279_bfr_after (
		.din(new_net_14278),
		.dout(new_net_14279)
	);

	bfr new_net_14280_bfr_after (
		.din(new_net_14279),
		.dout(new_net_14280)
	);

	bfr new_net_14281_bfr_after (
		.din(new_net_14280),
		.dout(new_net_14281)
	);

	bfr new_net_14282_bfr_after (
		.din(new_net_14281),
		.dout(new_net_14282)
	);

	bfr new_net_14283_bfr_after (
		.din(new_net_14282),
		.dout(new_net_14283)
	);

	bfr new_net_14284_bfr_after (
		.din(new_net_14283),
		.dout(new_net_14284)
	);

	bfr new_net_14285_bfr_after (
		.din(new_net_14284),
		.dout(new_net_14285)
	);

	bfr new_net_14286_bfr_after (
		.din(new_net_14285),
		.dout(new_net_14286)
	);

	bfr new_net_14287_bfr_after (
		.din(new_net_14286),
		.dout(new_net_14287)
	);

	bfr new_net_14288_bfr_after (
		.din(new_net_14287),
		.dout(new_net_14288)
	);

	bfr new_net_14289_bfr_after (
		.din(new_net_14288),
		.dout(new_net_14289)
	);

	bfr new_net_14290_bfr_after (
		.din(new_net_14289),
		.dout(new_net_14290)
	);

	bfr new_net_14291_bfr_after (
		.din(new_net_14290),
		.dout(new_net_14291)
	);

	bfr new_net_14292_bfr_after (
		.din(new_net_14291),
		.dout(new_net_14292)
	);

	bfr new_net_14293_bfr_after (
		.din(new_net_14292),
		.dout(new_net_14293)
	);

	bfr new_net_14294_bfr_after (
		.din(new_net_14293),
		.dout(new_net_14294)
	);

	bfr new_net_14295_bfr_after (
		.din(new_net_14294),
		.dout(new_net_14295)
	);

	bfr new_net_14296_bfr_after (
		.din(new_net_14295),
		.dout(new_net_14296)
	);

	bfr new_net_14297_bfr_after (
		.din(new_net_14296),
		.dout(new_net_14297)
	);

	bfr new_net_14298_bfr_after (
		.din(new_net_14297),
		.dout(new_net_14298)
	);

	bfr new_net_14299_bfr_after (
		.din(new_net_14298),
		.dout(new_net_14299)
	);

	bfr new_net_14300_bfr_after (
		.din(new_net_14299),
		.dout(new_net_14300)
	);

	bfr new_net_14301_bfr_after (
		.din(new_net_14300),
		.dout(new_net_14301)
	);

	bfr new_net_14302_bfr_after (
		.din(new_net_14301),
		.dout(new_net_14302)
	);

	bfr new_net_14303_bfr_after (
		.din(new_net_14302),
		.dout(new_net_14303)
	);

	bfr new_net_14304_bfr_after (
		.din(new_net_14303),
		.dout(new_net_14304)
	);

	bfr new_net_14305_bfr_after (
		.din(new_net_14304),
		.dout(new_net_14305)
	);

	bfr new_net_14306_bfr_after (
		.din(new_net_14305),
		.dout(new_net_14306)
	);

	bfr new_net_14307_bfr_after (
		.din(new_net_14306),
		.dout(new_net_14307)
	);

	bfr new_net_14308_bfr_after (
		.din(new_net_14307),
		.dout(new_net_14308)
	);

	bfr new_net_14309_bfr_after (
		.din(new_net_14308),
		.dout(new_net_14309)
	);

	bfr new_net_14310_bfr_after (
		.din(new_net_14309),
		.dout(new_net_14310)
	);

	bfr new_net_14311_bfr_after (
		.din(new_net_14310),
		.dout(new_net_14311)
	);

	bfr new_net_14312_bfr_after (
		.din(new_net_14311),
		.dout(new_net_14312)
	);

	bfr new_net_14313_bfr_after (
		.din(new_net_14312),
		.dout(new_net_14313)
	);

	bfr new_net_14314_bfr_after (
		.din(new_net_14313),
		.dout(new_net_14314)
	);

	bfr new_net_14315_bfr_after (
		.din(new_net_14314),
		.dout(new_net_14315)
	);

	bfr new_net_14316_bfr_after (
		.din(new_net_14315),
		.dout(new_net_14316)
	);

	bfr new_net_14317_bfr_after (
		.din(new_net_14316),
		.dout(new_net_14317)
	);

	bfr new_net_14318_bfr_after (
		.din(new_net_14317),
		.dout(new_net_14318)
	);

	bfr new_net_14319_bfr_after (
		.din(new_net_14318),
		.dout(new_net_14319)
	);

	bfr new_net_14320_bfr_after (
		.din(new_net_14319),
		.dout(new_net_14320)
	);

	bfr new_net_14321_bfr_after (
		.din(new_net_14320),
		.dout(new_net_14321)
	);

	spl2 _0439__v_fanout (
		.a(new_net_14321),
		.b(new_net_194),
		.c(new_net_195)
	);

	spl2 _1477__v_fanout (
		.a(_1477_),
		.b(new_net_3037),
		.c(new_net_3038)
	);

	bfr new_net_14322_bfr_after (
		.din(_1080_),
		.dout(new_net_14322)
	);

	bfr new_net_14323_bfr_after (
		.din(new_net_14322),
		.dout(new_net_14323)
	);

	bfr new_net_14324_bfr_after (
		.din(new_net_14323),
		.dout(new_net_14324)
	);

	bfr new_net_14325_bfr_after (
		.din(new_net_14324),
		.dout(new_net_14325)
	);

	bfr new_net_14326_bfr_after (
		.din(new_net_14325),
		.dout(new_net_14326)
	);

	bfr new_net_14327_bfr_after (
		.din(new_net_14326),
		.dout(new_net_14327)
	);

	bfr new_net_14328_bfr_after (
		.din(new_net_14327),
		.dout(new_net_14328)
	);

	bfr new_net_14329_bfr_after (
		.din(new_net_14328),
		.dout(new_net_14329)
	);

	bfr new_net_14330_bfr_after (
		.din(new_net_14329),
		.dout(new_net_14330)
	);

	bfr new_net_14331_bfr_after (
		.din(new_net_14330),
		.dout(new_net_14331)
	);

	bfr new_net_14332_bfr_after (
		.din(new_net_14331),
		.dout(new_net_14332)
	);

	bfr new_net_14333_bfr_after (
		.din(new_net_14332),
		.dout(new_net_14333)
	);

	bfr new_net_14334_bfr_after (
		.din(new_net_14333),
		.dout(new_net_14334)
	);

	bfr new_net_14335_bfr_after (
		.din(new_net_14334),
		.dout(new_net_14335)
	);

	bfr new_net_14336_bfr_after (
		.din(new_net_14335),
		.dout(new_net_14336)
	);

	bfr new_net_14337_bfr_after (
		.din(new_net_14336),
		.dout(new_net_14337)
	);

	spl2 _1080__v_fanout (
		.a(new_net_14337),
		.b(new_net_1656),
		.c(new_net_1657)
	);

	spl2 _0350__v_fanout (
		.a(_0350_),
		.b(new_net_20),
		.c(new_net_21)
	);

	bfr new_net_14338_bfr_after (
		.din(_0710_),
		.dout(new_net_14338)
	);

	bfr new_net_14339_bfr_after (
		.din(new_net_14338),
		.dout(new_net_14339)
	);

	bfr new_net_14340_bfr_after (
		.din(new_net_14339),
		.dout(new_net_14340)
	);

	bfr new_net_14341_bfr_after (
		.din(new_net_14340),
		.dout(new_net_14341)
	);

	bfr new_net_14342_bfr_after (
		.din(new_net_14341),
		.dout(new_net_14342)
	);

	bfr new_net_14343_bfr_after (
		.din(new_net_14342),
		.dout(new_net_14343)
	);

	bfr new_net_14344_bfr_after (
		.din(new_net_14343),
		.dout(new_net_14344)
	);

	bfr new_net_14345_bfr_after (
		.din(new_net_14344),
		.dout(new_net_14345)
	);

	bfr new_net_14346_bfr_after (
		.din(new_net_14345),
		.dout(new_net_14346)
	);

	bfr new_net_14347_bfr_after (
		.din(new_net_14346),
		.dout(new_net_14347)
	);

	bfr new_net_14348_bfr_after (
		.din(new_net_14347),
		.dout(new_net_14348)
	);

	bfr new_net_14349_bfr_after (
		.din(new_net_14348),
		.dout(new_net_14349)
	);

	bfr new_net_14350_bfr_after (
		.din(new_net_14349),
		.dout(new_net_14350)
	);

	bfr new_net_14351_bfr_after (
		.din(new_net_14350),
		.dout(new_net_14351)
	);

	bfr new_net_14352_bfr_after (
		.din(new_net_14351),
		.dout(new_net_14352)
	);

	bfr new_net_14353_bfr_after (
		.din(new_net_14352),
		.dout(new_net_14353)
	);

	bfr new_net_14354_bfr_after (
		.din(new_net_14353),
		.dout(new_net_14354)
	);

	bfr new_net_14355_bfr_after (
		.din(new_net_14354),
		.dout(new_net_14355)
	);

	bfr new_net_14356_bfr_after (
		.din(new_net_14355),
		.dout(new_net_14356)
	);

	bfr new_net_14357_bfr_after (
		.din(new_net_14356),
		.dout(new_net_14357)
	);

	bfr new_net_14358_bfr_after (
		.din(new_net_14357),
		.dout(new_net_14358)
	);

	bfr new_net_14359_bfr_after (
		.din(new_net_14358),
		.dout(new_net_14359)
	);

	bfr new_net_14360_bfr_after (
		.din(new_net_14359),
		.dout(new_net_14360)
	);

	bfr new_net_14361_bfr_after (
		.din(new_net_14360),
		.dout(new_net_14361)
	);

	bfr new_net_14362_bfr_after (
		.din(new_net_14361),
		.dout(new_net_14362)
	);

	bfr new_net_14363_bfr_after (
		.din(new_net_14362),
		.dout(new_net_14363)
	);

	bfr new_net_14364_bfr_after (
		.din(new_net_14363),
		.dout(new_net_14364)
	);

	bfr new_net_14365_bfr_after (
		.din(new_net_14364),
		.dout(new_net_14365)
	);

	bfr new_net_14366_bfr_after (
		.din(new_net_14365),
		.dout(new_net_14366)
	);

	bfr new_net_14367_bfr_after (
		.din(new_net_14366),
		.dout(new_net_14367)
	);

	bfr new_net_14368_bfr_after (
		.din(new_net_14367),
		.dout(new_net_14368)
	);

	bfr new_net_14369_bfr_after (
		.din(new_net_14368),
		.dout(new_net_14369)
	);

	bfr new_net_14370_bfr_after (
		.din(new_net_14369),
		.dout(new_net_14370)
	);

	bfr new_net_14371_bfr_after (
		.din(new_net_14370),
		.dout(new_net_14371)
	);

	bfr new_net_14372_bfr_after (
		.din(new_net_14371),
		.dout(new_net_14372)
	);

	bfr new_net_14373_bfr_after (
		.din(new_net_14372),
		.dout(new_net_14373)
	);

	bfr new_net_14374_bfr_after (
		.din(new_net_14373),
		.dout(new_net_14374)
	);

	bfr new_net_14375_bfr_after (
		.din(new_net_14374),
		.dout(new_net_14375)
	);

	bfr new_net_14376_bfr_after (
		.din(new_net_14375),
		.dout(new_net_14376)
	);

	bfr new_net_14377_bfr_after (
		.din(new_net_14376),
		.dout(new_net_14377)
	);

	bfr new_net_14378_bfr_after (
		.din(new_net_14377),
		.dout(new_net_14378)
	);

	bfr new_net_14379_bfr_after (
		.din(new_net_14378),
		.dout(new_net_14379)
	);

	bfr new_net_14380_bfr_after (
		.din(new_net_14379),
		.dout(new_net_14380)
	);

	bfr new_net_14381_bfr_after (
		.din(new_net_14380),
		.dout(new_net_14381)
	);

	bfr new_net_14382_bfr_after (
		.din(new_net_14381),
		.dout(new_net_14382)
	);

	bfr new_net_14383_bfr_after (
		.din(new_net_14382),
		.dout(new_net_14383)
	);

	bfr new_net_14384_bfr_after (
		.din(new_net_14383),
		.dout(new_net_14384)
	);

	bfr new_net_14385_bfr_after (
		.din(new_net_14384),
		.dout(new_net_14385)
	);

	bfr new_net_14386_bfr_after (
		.din(new_net_14385),
		.dout(new_net_14386)
	);

	bfr new_net_14387_bfr_after (
		.din(new_net_14386),
		.dout(new_net_14387)
	);

	bfr new_net_14388_bfr_after (
		.din(new_net_14387),
		.dout(new_net_14388)
	);

	bfr new_net_14389_bfr_after (
		.din(new_net_14388),
		.dout(new_net_14389)
	);

	bfr new_net_14390_bfr_after (
		.din(new_net_14389),
		.dout(new_net_14390)
	);

	bfr new_net_14391_bfr_after (
		.din(new_net_14390),
		.dout(new_net_14391)
	);

	bfr new_net_14392_bfr_after (
		.din(new_net_14391),
		.dout(new_net_14392)
	);

	bfr new_net_14393_bfr_after (
		.din(new_net_14392),
		.dout(new_net_14393)
	);

	bfr new_net_14394_bfr_after (
		.din(new_net_14393),
		.dout(new_net_14394)
	);

	bfr new_net_14395_bfr_after (
		.din(new_net_14394),
		.dout(new_net_14395)
	);

	spl2 _0710__v_fanout (
		.a(new_net_14395),
		.b(new_net_1008),
		.c(new_net_1009)
	);

	bfr new_net_14396_bfr_after (
		.din(_0987_),
		.dout(new_net_14396)
	);

	bfr new_net_14397_bfr_after (
		.din(new_net_14396),
		.dout(new_net_14397)
	);

	bfr new_net_14398_bfr_after (
		.din(new_net_14397),
		.dout(new_net_14398)
	);

	bfr new_net_14399_bfr_after (
		.din(new_net_14398),
		.dout(new_net_14399)
	);

	bfr new_net_14400_bfr_after (
		.din(new_net_14399),
		.dout(new_net_14400)
	);

	bfr new_net_14401_bfr_after (
		.din(new_net_14400),
		.dout(new_net_14401)
	);

	bfr new_net_14402_bfr_after (
		.din(new_net_14401),
		.dout(new_net_14402)
	);

	bfr new_net_14403_bfr_after (
		.din(new_net_14402),
		.dout(new_net_14403)
	);

	bfr new_net_14404_bfr_after (
		.din(new_net_14403),
		.dout(new_net_14404)
	);

	bfr new_net_14405_bfr_after (
		.din(new_net_14404),
		.dout(new_net_14405)
	);

	bfr new_net_14406_bfr_after (
		.din(new_net_14405),
		.dout(new_net_14406)
	);

	bfr new_net_14407_bfr_after (
		.din(new_net_14406),
		.dout(new_net_14407)
	);

	bfr new_net_14408_bfr_after (
		.din(new_net_14407),
		.dout(new_net_14408)
	);

	bfr new_net_14409_bfr_after (
		.din(new_net_14408),
		.dout(new_net_14409)
	);

	bfr new_net_14410_bfr_after (
		.din(new_net_14409),
		.dout(new_net_14410)
	);

	bfr new_net_14411_bfr_after (
		.din(new_net_14410),
		.dout(new_net_14411)
	);

	bfr new_net_14412_bfr_after (
		.din(new_net_14411),
		.dout(new_net_14412)
	);

	bfr new_net_14413_bfr_after (
		.din(new_net_14412),
		.dout(new_net_14413)
	);

	bfr new_net_14414_bfr_after (
		.din(new_net_14413),
		.dout(new_net_14414)
	);

	bfr new_net_14415_bfr_after (
		.din(new_net_14414),
		.dout(new_net_14415)
	);

	bfr new_net_14416_bfr_after (
		.din(new_net_14415),
		.dout(new_net_14416)
	);

	bfr new_net_14417_bfr_after (
		.din(new_net_14416),
		.dout(new_net_14417)
	);

	bfr new_net_14418_bfr_after (
		.din(new_net_14417),
		.dout(new_net_14418)
	);

	bfr new_net_14419_bfr_after (
		.din(new_net_14418),
		.dout(new_net_14419)
	);

	bfr new_net_14420_bfr_after (
		.din(new_net_14419),
		.dout(new_net_14420)
	);

	bfr new_net_14421_bfr_after (
		.din(new_net_14420),
		.dout(new_net_14421)
	);

	bfr new_net_14422_bfr_after (
		.din(new_net_14421),
		.dout(new_net_14422)
	);

	bfr new_net_14423_bfr_after (
		.din(new_net_14422),
		.dout(new_net_14423)
	);

	bfr new_net_14424_bfr_after (
		.din(new_net_14423),
		.dout(new_net_14424)
	);

	bfr new_net_14425_bfr_after (
		.din(new_net_14424),
		.dout(new_net_14425)
	);

	bfr new_net_14426_bfr_after (
		.din(new_net_14425),
		.dout(new_net_14426)
	);

	bfr new_net_14427_bfr_after (
		.din(new_net_14426),
		.dout(new_net_14427)
	);

	bfr new_net_14428_bfr_after (
		.din(new_net_14427),
		.dout(new_net_14428)
	);

	bfr new_net_14429_bfr_after (
		.din(new_net_14428),
		.dout(new_net_14429)
	);

	bfr new_net_14430_bfr_after (
		.din(new_net_14429),
		.dout(new_net_14430)
	);

	bfr new_net_14431_bfr_after (
		.din(new_net_14430),
		.dout(new_net_14431)
	);

	bfr new_net_14432_bfr_after (
		.din(new_net_14431),
		.dout(new_net_14432)
	);

	bfr new_net_14433_bfr_after (
		.din(new_net_14432),
		.dout(new_net_14433)
	);

	bfr new_net_14434_bfr_after (
		.din(new_net_14433),
		.dout(new_net_14434)
	);

	bfr new_net_14435_bfr_after (
		.din(new_net_14434),
		.dout(new_net_14435)
	);

	bfr new_net_14436_bfr_after (
		.din(new_net_14435),
		.dout(new_net_14436)
	);

	bfr new_net_14437_bfr_after (
		.din(new_net_14436),
		.dout(new_net_14437)
	);

	bfr new_net_14438_bfr_after (
		.din(new_net_14437),
		.dout(new_net_14438)
	);

	bfr new_net_14439_bfr_after (
		.din(new_net_14438),
		.dout(new_net_14439)
	);

	bfr new_net_14440_bfr_after (
		.din(new_net_14439),
		.dout(new_net_14440)
	);

	bfr new_net_14441_bfr_after (
		.din(new_net_14440),
		.dout(new_net_14441)
	);

	bfr new_net_14442_bfr_after (
		.din(new_net_14441),
		.dout(new_net_14442)
	);

	bfr new_net_14443_bfr_after (
		.din(new_net_14442),
		.dout(new_net_14443)
	);

	bfr new_net_14444_bfr_after (
		.din(new_net_14443),
		.dout(new_net_14444)
	);

	bfr new_net_14445_bfr_after (
		.din(new_net_14444),
		.dout(new_net_14445)
	);

	bfr new_net_14446_bfr_after (
		.din(new_net_14445),
		.dout(new_net_14446)
	);

	bfr new_net_14447_bfr_after (
		.din(new_net_14446),
		.dout(new_net_14447)
	);

	bfr new_net_14448_bfr_after (
		.din(new_net_14447),
		.dout(new_net_14448)
	);

	bfr new_net_14449_bfr_after (
		.din(new_net_14448),
		.dout(new_net_14449)
	);

	bfr new_net_14450_bfr_after (
		.din(new_net_14449),
		.dout(new_net_14450)
	);

	bfr new_net_14451_bfr_after (
		.din(new_net_14450),
		.dout(new_net_14451)
	);

	bfr new_net_14452_bfr_after (
		.din(new_net_14451),
		.dout(new_net_14452)
	);

	bfr new_net_14453_bfr_after (
		.din(new_net_14452),
		.dout(new_net_14453)
	);

	bfr new_net_14454_bfr_after (
		.din(new_net_14453),
		.dout(new_net_14454)
	);

	bfr new_net_14455_bfr_after (
		.din(new_net_14454),
		.dout(new_net_14455)
	);

	bfr new_net_14456_bfr_after (
		.din(new_net_14455),
		.dout(new_net_14456)
	);

	bfr new_net_14457_bfr_after (
		.din(new_net_14456),
		.dout(new_net_14457)
	);

	bfr new_net_14458_bfr_after (
		.din(new_net_14457),
		.dout(new_net_14458)
	);

	bfr new_net_14459_bfr_after (
		.din(new_net_14458),
		.dout(new_net_14459)
	);

	bfr new_net_14460_bfr_after (
		.din(new_net_14459),
		.dout(new_net_14460)
	);

	bfr new_net_14461_bfr_after (
		.din(new_net_14460),
		.dout(new_net_14461)
	);

	bfr new_net_14462_bfr_after (
		.din(new_net_14461),
		.dout(new_net_14462)
	);

	bfr new_net_14463_bfr_after (
		.din(new_net_14462),
		.dout(new_net_14463)
	);

	bfr new_net_14464_bfr_after (
		.din(new_net_14463),
		.dout(new_net_14464)
	);

	bfr new_net_14465_bfr_after (
		.din(new_net_14464),
		.dout(new_net_14465)
	);

	bfr new_net_14466_bfr_after (
		.din(new_net_14465),
		.dout(new_net_14466)
	);

	bfr new_net_14467_bfr_after (
		.din(new_net_14466),
		.dout(new_net_14467)
	);

	bfr new_net_14468_bfr_after (
		.din(new_net_14467),
		.dout(new_net_14468)
	);

	bfr new_net_14469_bfr_after (
		.din(new_net_14468),
		.dout(new_net_14469)
	);

	bfr new_net_14470_bfr_after (
		.din(new_net_14469),
		.dout(new_net_14470)
	);

	bfr new_net_14471_bfr_after (
		.din(new_net_14470),
		.dout(new_net_14471)
	);

	bfr new_net_14472_bfr_after (
		.din(new_net_14471),
		.dout(new_net_14472)
	);

	bfr new_net_14473_bfr_after (
		.din(new_net_14472),
		.dout(new_net_14473)
	);

	bfr new_net_14474_bfr_after (
		.din(new_net_14473),
		.dout(new_net_14474)
	);

	bfr new_net_14475_bfr_after (
		.din(new_net_14474),
		.dout(new_net_14475)
	);

	bfr new_net_14476_bfr_after (
		.din(new_net_14475),
		.dout(new_net_14476)
	);

	bfr new_net_14477_bfr_after (
		.din(new_net_14476),
		.dout(new_net_14477)
	);

	bfr new_net_14478_bfr_after (
		.din(new_net_14477),
		.dout(new_net_14478)
	);

	bfr new_net_14479_bfr_after (
		.din(new_net_14478),
		.dout(new_net_14479)
	);

	bfr new_net_14480_bfr_after (
		.din(new_net_14479),
		.dout(new_net_14480)
	);

	bfr new_net_14481_bfr_after (
		.din(new_net_14480),
		.dout(new_net_14481)
	);

	bfr new_net_14482_bfr_after (
		.din(new_net_14481),
		.dout(new_net_14482)
	);

	bfr new_net_14483_bfr_after (
		.din(new_net_14482),
		.dout(new_net_14483)
	);

	bfr new_net_14484_bfr_after (
		.din(new_net_14483),
		.dout(new_net_14484)
	);

	bfr new_net_14485_bfr_after (
		.din(new_net_14484),
		.dout(new_net_14485)
	);

	bfr new_net_14486_bfr_after (
		.din(new_net_14485),
		.dout(new_net_14486)
	);

	bfr new_net_14487_bfr_after (
		.din(new_net_14486),
		.dout(new_net_14487)
	);

	bfr new_net_14488_bfr_after (
		.din(new_net_14487),
		.dout(new_net_14488)
	);

	bfr new_net_14489_bfr_after (
		.din(new_net_14488),
		.dout(new_net_14489)
	);

	bfr new_net_14490_bfr_after (
		.din(new_net_14489),
		.dout(new_net_14490)
	);

	bfr new_net_14491_bfr_after (
		.din(new_net_14490),
		.dout(new_net_14491)
	);

	bfr new_net_14492_bfr_after (
		.din(new_net_14491),
		.dout(new_net_14492)
	);

	bfr new_net_14493_bfr_after (
		.din(new_net_14492),
		.dout(new_net_14493)
	);

	bfr new_net_14494_bfr_after (
		.din(new_net_14493),
		.dout(new_net_14494)
	);

	bfr new_net_14495_bfr_after (
		.din(new_net_14494),
		.dout(new_net_14495)
	);

	bfr new_net_14496_bfr_after (
		.din(new_net_14495),
		.dout(new_net_14496)
	);

	bfr new_net_14497_bfr_after (
		.din(new_net_14496),
		.dout(new_net_14497)
	);

	bfr new_net_14498_bfr_after (
		.din(new_net_14497),
		.dout(new_net_14498)
	);

	bfr new_net_14499_bfr_after (
		.din(new_net_14498),
		.dout(new_net_14499)
	);

	bfr new_net_14500_bfr_after (
		.din(new_net_14499),
		.dout(new_net_14500)
	);

	bfr new_net_14501_bfr_after (
		.din(new_net_14500),
		.dout(new_net_14501)
	);

	spl2 _0987__v_fanout (
		.a(new_net_14501),
		.b(new_net_1816),
		.c(new_net_1817)
	);

	bfr new_net_14502_bfr_after (
		.din(_0335_),
		.dout(new_net_14502)
	);

	bfr new_net_14503_bfr_after (
		.din(new_net_14502),
		.dout(new_net_14503)
	);

	bfr new_net_14504_bfr_after (
		.din(new_net_14503),
		.dout(new_net_14504)
	);

	bfr new_net_14505_bfr_after (
		.din(new_net_14504),
		.dout(new_net_14505)
	);

	bfr new_net_14506_bfr_after (
		.din(new_net_14505),
		.dout(new_net_14506)
	);

	bfr new_net_14507_bfr_after (
		.din(new_net_14506),
		.dout(new_net_14507)
	);

	bfr new_net_14508_bfr_after (
		.din(new_net_14507),
		.dout(new_net_14508)
	);

	bfr new_net_14509_bfr_after (
		.din(new_net_14508),
		.dout(new_net_14509)
	);

	bfr new_net_14510_bfr_after (
		.din(new_net_14509),
		.dout(new_net_14510)
	);

	bfr new_net_14511_bfr_after (
		.din(new_net_14510),
		.dout(new_net_14511)
	);

	bfr new_net_14512_bfr_after (
		.din(new_net_14511),
		.dout(new_net_14512)
	);

	bfr new_net_14513_bfr_after (
		.din(new_net_14512),
		.dout(new_net_14513)
	);

	bfr new_net_14514_bfr_after (
		.din(new_net_14513),
		.dout(new_net_14514)
	);

	bfr new_net_14515_bfr_after (
		.din(new_net_14514),
		.dout(new_net_14515)
	);

	bfr new_net_14516_bfr_after (
		.din(new_net_14515),
		.dout(new_net_14516)
	);

	bfr new_net_14517_bfr_after (
		.din(new_net_14516),
		.dout(new_net_14517)
	);

	bfr new_net_14518_bfr_after (
		.din(new_net_14517),
		.dout(new_net_14518)
	);

	bfr new_net_14519_bfr_after (
		.din(new_net_14518),
		.dout(new_net_14519)
	);

	bfr new_net_14520_bfr_after (
		.din(new_net_14519),
		.dout(new_net_14520)
	);

	bfr new_net_14521_bfr_after (
		.din(new_net_14520),
		.dout(new_net_14521)
	);

	bfr new_net_14522_bfr_after (
		.din(new_net_14521),
		.dout(new_net_14522)
	);

	bfr new_net_14523_bfr_after (
		.din(new_net_14522),
		.dout(new_net_14523)
	);

	bfr new_net_14524_bfr_after (
		.din(new_net_14523),
		.dout(new_net_14524)
	);

	bfr new_net_14525_bfr_after (
		.din(new_net_14524),
		.dout(new_net_14525)
	);

	bfr new_net_14526_bfr_after (
		.din(new_net_14525),
		.dout(new_net_14526)
	);

	bfr new_net_14527_bfr_after (
		.din(new_net_14526),
		.dout(new_net_14527)
	);

	bfr new_net_14528_bfr_after (
		.din(new_net_14527),
		.dout(new_net_14528)
	);

	bfr new_net_14529_bfr_after (
		.din(new_net_14528),
		.dout(new_net_14529)
	);

	bfr new_net_14530_bfr_after (
		.din(new_net_14529),
		.dout(new_net_14530)
	);

	bfr new_net_14531_bfr_after (
		.din(new_net_14530),
		.dout(new_net_14531)
	);

	bfr new_net_14532_bfr_after (
		.din(new_net_14531),
		.dout(new_net_14532)
	);

	bfr new_net_14533_bfr_after (
		.din(new_net_14532),
		.dout(new_net_14533)
	);

	bfr new_net_14534_bfr_after (
		.din(new_net_14533),
		.dout(new_net_14534)
	);

	bfr new_net_14535_bfr_after (
		.din(new_net_14534),
		.dout(new_net_14535)
	);

	bfr new_net_14536_bfr_after (
		.din(new_net_14535),
		.dout(new_net_14536)
	);

	bfr new_net_14537_bfr_after (
		.din(new_net_14536),
		.dout(new_net_14537)
	);

	bfr new_net_14538_bfr_after (
		.din(new_net_14537),
		.dout(new_net_14538)
	);

	bfr new_net_14539_bfr_after (
		.din(new_net_14538),
		.dout(new_net_14539)
	);

	bfr new_net_14540_bfr_after (
		.din(new_net_14539),
		.dout(new_net_14540)
	);

	bfr new_net_14541_bfr_after (
		.din(new_net_14540),
		.dout(new_net_14541)
	);

	bfr new_net_14542_bfr_after (
		.din(new_net_14541),
		.dout(new_net_14542)
	);

	bfr new_net_14543_bfr_after (
		.din(new_net_14542),
		.dout(new_net_14543)
	);

	bfr new_net_14544_bfr_after (
		.din(new_net_14543),
		.dout(new_net_14544)
	);

	bfr new_net_14545_bfr_after (
		.din(new_net_14544),
		.dout(new_net_14545)
	);

	bfr new_net_14546_bfr_after (
		.din(new_net_14545),
		.dout(new_net_14546)
	);

	bfr new_net_14547_bfr_after (
		.din(new_net_14546),
		.dout(new_net_14547)
	);

	bfr new_net_14548_bfr_after (
		.din(new_net_14547),
		.dout(new_net_14548)
	);

	bfr new_net_14549_bfr_after (
		.din(new_net_14548),
		.dout(new_net_14549)
	);

	bfr new_net_14550_bfr_after (
		.din(new_net_14549),
		.dout(new_net_14550)
	);

	bfr new_net_14551_bfr_after (
		.din(new_net_14550),
		.dout(new_net_14551)
	);

	bfr new_net_14552_bfr_after (
		.din(new_net_14551),
		.dout(new_net_14552)
	);

	bfr new_net_14553_bfr_after (
		.din(new_net_14552),
		.dout(new_net_14553)
	);

	bfr new_net_14554_bfr_after (
		.din(new_net_14553),
		.dout(new_net_14554)
	);

	bfr new_net_14555_bfr_after (
		.din(new_net_14554),
		.dout(new_net_14555)
	);

	bfr new_net_14556_bfr_after (
		.din(new_net_14555),
		.dout(new_net_14556)
	);

	bfr new_net_14557_bfr_after (
		.din(new_net_14556),
		.dout(new_net_14557)
	);

	bfr new_net_14558_bfr_after (
		.din(new_net_14557),
		.dout(new_net_14558)
	);

	bfr new_net_14559_bfr_after (
		.din(new_net_14558),
		.dout(new_net_14559)
	);

	bfr new_net_14560_bfr_after (
		.din(new_net_14559),
		.dout(new_net_14560)
	);

	bfr new_net_14561_bfr_after (
		.din(new_net_14560),
		.dout(new_net_14561)
	);

	bfr new_net_14562_bfr_after (
		.din(new_net_14561),
		.dout(new_net_14562)
	);

	bfr new_net_14563_bfr_after (
		.din(new_net_14562),
		.dout(new_net_14563)
	);

	bfr new_net_14564_bfr_after (
		.din(new_net_14563),
		.dout(new_net_14564)
	);

	bfr new_net_14565_bfr_after (
		.din(new_net_14564),
		.dout(new_net_14565)
	);

	bfr new_net_14566_bfr_after (
		.din(new_net_14565),
		.dout(new_net_14566)
	);

	bfr new_net_14567_bfr_after (
		.din(new_net_14566),
		.dout(new_net_14567)
	);

	bfr new_net_14568_bfr_after (
		.din(new_net_14567),
		.dout(new_net_14568)
	);

	bfr new_net_14569_bfr_after (
		.din(new_net_14568),
		.dout(new_net_14569)
	);

	bfr new_net_14570_bfr_after (
		.din(new_net_14569),
		.dout(new_net_14570)
	);

	bfr new_net_14571_bfr_after (
		.din(new_net_14570),
		.dout(new_net_14571)
	);

	bfr new_net_14572_bfr_after (
		.din(new_net_14571),
		.dout(new_net_14572)
	);

	bfr new_net_14573_bfr_after (
		.din(new_net_14572),
		.dout(new_net_14573)
	);

	bfr new_net_14574_bfr_after (
		.din(new_net_14573),
		.dout(new_net_14574)
	);

	bfr new_net_14575_bfr_after (
		.din(new_net_14574),
		.dout(new_net_14575)
	);

	bfr new_net_14576_bfr_after (
		.din(new_net_14575),
		.dout(new_net_14576)
	);

	bfr new_net_14577_bfr_after (
		.din(new_net_14576),
		.dout(new_net_14577)
	);

	bfr new_net_14578_bfr_after (
		.din(new_net_14577),
		.dout(new_net_14578)
	);

	bfr new_net_14579_bfr_after (
		.din(new_net_14578),
		.dout(new_net_14579)
	);

	bfr new_net_14580_bfr_after (
		.din(new_net_14579),
		.dout(new_net_14580)
	);

	bfr new_net_14581_bfr_after (
		.din(new_net_14580),
		.dout(new_net_14581)
	);

	spl2 _0335__v_fanout (
		.a(new_net_14581),
		.b(new_net_1024),
		.c(new_net_1025)
	);

	bfr new_net_14582_bfr_after (
		.din(_1375_),
		.dout(new_net_14582)
	);

	bfr new_net_14583_bfr_after (
		.din(new_net_14582),
		.dout(new_net_14583)
	);

	bfr new_net_14584_bfr_after (
		.din(new_net_14583),
		.dout(new_net_14584)
	);

	bfr new_net_14585_bfr_after (
		.din(new_net_14584),
		.dout(new_net_14585)
	);

	bfr new_net_14586_bfr_after (
		.din(new_net_14585),
		.dout(new_net_14586)
	);

	bfr new_net_14587_bfr_after (
		.din(new_net_14586),
		.dout(new_net_14587)
	);

	bfr new_net_14588_bfr_after (
		.din(new_net_14587),
		.dout(new_net_14588)
	);

	bfr new_net_14589_bfr_after (
		.din(new_net_14588),
		.dout(new_net_14589)
	);

	bfr new_net_14590_bfr_after (
		.din(new_net_14589),
		.dout(new_net_14590)
	);

	bfr new_net_14591_bfr_after (
		.din(new_net_14590),
		.dout(new_net_14591)
	);

	bfr new_net_14592_bfr_after (
		.din(new_net_14591),
		.dout(new_net_14592)
	);

	bfr new_net_14593_bfr_after (
		.din(new_net_14592),
		.dout(new_net_14593)
	);

	bfr new_net_14594_bfr_after (
		.din(new_net_14593),
		.dout(new_net_14594)
	);

	bfr new_net_14595_bfr_after (
		.din(new_net_14594),
		.dout(new_net_14595)
	);

	bfr new_net_14596_bfr_after (
		.din(new_net_14595),
		.dout(new_net_14596)
	);

	bfr new_net_14597_bfr_after (
		.din(new_net_14596),
		.dout(new_net_14597)
	);

	bfr new_net_14598_bfr_after (
		.din(new_net_14597),
		.dout(new_net_14598)
	);

	bfr new_net_14599_bfr_after (
		.din(new_net_14598),
		.dout(new_net_14599)
	);

	bfr new_net_14600_bfr_after (
		.din(new_net_14599),
		.dout(new_net_14600)
	);

	bfr new_net_14601_bfr_after (
		.din(new_net_14600),
		.dout(new_net_14601)
	);

	bfr new_net_14602_bfr_after (
		.din(new_net_14601),
		.dout(new_net_14602)
	);

	bfr new_net_14603_bfr_after (
		.din(new_net_14602),
		.dout(new_net_14603)
	);

	bfr new_net_14604_bfr_after (
		.din(new_net_14603),
		.dout(new_net_14604)
	);

	bfr new_net_14605_bfr_after (
		.din(new_net_14604),
		.dout(new_net_14605)
	);

	bfr new_net_14606_bfr_after (
		.din(new_net_14605),
		.dout(new_net_14606)
	);

	bfr new_net_14607_bfr_after (
		.din(new_net_14606),
		.dout(new_net_14607)
	);

	bfr new_net_14608_bfr_after (
		.din(new_net_14607),
		.dout(new_net_14608)
	);

	bfr new_net_14609_bfr_after (
		.din(new_net_14608),
		.dout(new_net_14609)
	);

	bfr new_net_14610_bfr_after (
		.din(new_net_14609),
		.dout(new_net_14610)
	);

	bfr new_net_14611_bfr_after (
		.din(new_net_14610),
		.dout(new_net_14611)
	);

	bfr new_net_14612_bfr_after (
		.din(new_net_14611),
		.dout(new_net_14612)
	);

	bfr new_net_14613_bfr_after (
		.din(new_net_14612),
		.dout(new_net_14613)
	);

	spl2 _1375__v_fanout (
		.a(new_net_14613),
		.b(new_net_2228),
		.c(new_net_2229)
	);

	spl2 _1479__v_fanout (
		.a(_1479_),
		.b(new_net_1372),
		.c(new_net_1373)
	);

	bfr new_net_14614_bfr_after (
		.din(_0348_),
		.dout(new_net_14614)
	);

	bfr new_net_14615_bfr_after (
		.din(new_net_14614),
		.dout(new_net_14615)
	);

	bfr new_net_14616_bfr_after (
		.din(new_net_14615),
		.dout(new_net_14616)
	);

	bfr new_net_14617_bfr_after (
		.din(new_net_14616),
		.dout(new_net_14617)
	);

	bfr new_net_14618_bfr_after (
		.din(new_net_14617),
		.dout(new_net_14618)
	);

	bfr new_net_14619_bfr_after (
		.din(new_net_14618),
		.dout(new_net_14619)
	);

	bfr new_net_14620_bfr_after (
		.din(new_net_14619),
		.dout(new_net_14620)
	);

	bfr new_net_14621_bfr_after (
		.din(new_net_14620),
		.dout(new_net_14621)
	);

	bfr new_net_14622_bfr_after (
		.din(new_net_14621),
		.dout(new_net_14622)
	);

	bfr new_net_14623_bfr_after (
		.din(new_net_14622),
		.dout(new_net_14623)
	);

	bfr new_net_14624_bfr_after (
		.din(new_net_14623),
		.dout(new_net_14624)
	);

	bfr new_net_14625_bfr_after (
		.din(new_net_14624),
		.dout(new_net_14625)
	);

	bfr new_net_14626_bfr_after (
		.din(new_net_14625),
		.dout(new_net_14626)
	);

	bfr new_net_14627_bfr_after (
		.din(new_net_14626),
		.dout(new_net_14627)
	);

	bfr new_net_14628_bfr_after (
		.din(new_net_14627),
		.dout(new_net_14628)
	);

	bfr new_net_14629_bfr_after (
		.din(new_net_14628),
		.dout(new_net_14629)
	);

	bfr new_net_14630_bfr_after (
		.din(new_net_14629),
		.dout(new_net_14630)
	);

	bfr new_net_14631_bfr_after (
		.din(new_net_14630),
		.dout(new_net_14631)
	);

	bfr new_net_14632_bfr_after (
		.din(new_net_14631),
		.dout(new_net_14632)
	);

	bfr new_net_14633_bfr_after (
		.din(new_net_14632),
		.dout(new_net_14633)
	);

	bfr new_net_14634_bfr_after (
		.din(new_net_14633),
		.dout(new_net_14634)
	);

	bfr new_net_14635_bfr_after (
		.din(new_net_14634),
		.dout(new_net_14635)
	);

	bfr new_net_14636_bfr_after (
		.din(new_net_14635),
		.dout(new_net_14636)
	);

	bfr new_net_14637_bfr_after (
		.din(new_net_14636),
		.dout(new_net_14637)
	);

	bfr new_net_14638_bfr_after (
		.din(new_net_14637),
		.dout(new_net_14638)
	);

	bfr new_net_14639_bfr_after (
		.din(new_net_14638),
		.dout(new_net_14639)
	);

	spl2 _0348__v_fanout (
		.a(new_net_14639),
		.b(new_net_2746),
		.c(new_net_2747)
	);

	bfr new_net_14640_bfr_after (
		.din(_0771_),
		.dout(new_net_14640)
	);

	bfr new_net_14641_bfr_after (
		.din(new_net_14640),
		.dout(new_net_14641)
	);

	bfr new_net_14642_bfr_after (
		.din(new_net_14641),
		.dout(new_net_14642)
	);

	bfr new_net_14643_bfr_after (
		.din(new_net_14642),
		.dout(new_net_14643)
	);

	bfr new_net_14644_bfr_after (
		.din(new_net_14643),
		.dout(new_net_14644)
	);

	bfr new_net_14645_bfr_after (
		.din(new_net_14644),
		.dout(new_net_14645)
	);

	bfr new_net_14646_bfr_after (
		.din(new_net_14645),
		.dout(new_net_14646)
	);

	bfr new_net_14647_bfr_after (
		.din(new_net_14646),
		.dout(new_net_14647)
	);

	bfr new_net_14648_bfr_after (
		.din(new_net_14647),
		.dout(new_net_14648)
	);

	bfr new_net_14649_bfr_after (
		.din(new_net_14648),
		.dout(new_net_14649)
	);

	bfr new_net_14650_bfr_after (
		.din(new_net_14649),
		.dout(new_net_14650)
	);

	bfr new_net_14651_bfr_after (
		.din(new_net_14650),
		.dout(new_net_14651)
	);

	bfr new_net_14652_bfr_after (
		.din(new_net_14651),
		.dout(new_net_14652)
	);

	bfr new_net_14653_bfr_after (
		.din(new_net_14652),
		.dout(new_net_14653)
	);

	bfr new_net_14654_bfr_after (
		.din(new_net_14653),
		.dout(new_net_14654)
	);

	bfr new_net_14655_bfr_after (
		.din(new_net_14654),
		.dout(new_net_14655)
	);

	bfr new_net_14656_bfr_after (
		.din(new_net_14655),
		.dout(new_net_14656)
	);

	bfr new_net_14657_bfr_after (
		.din(new_net_14656),
		.dout(new_net_14657)
	);

	bfr new_net_14658_bfr_after (
		.din(new_net_14657),
		.dout(new_net_14658)
	);

	bfr new_net_14659_bfr_after (
		.din(new_net_14658),
		.dout(new_net_14659)
	);

	bfr new_net_14660_bfr_after (
		.din(new_net_14659),
		.dout(new_net_14660)
	);

	bfr new_net_14661_bfr_after (
		.din(new_net_14660),
		.dout(new_net_14661)
	);

	bfr new_net_14662_bfr_after (
		.din(new_net_14661),
		.dout(new_net_14662)
	);

	bfr new_net_14663_bfr_after (
		.din(new_net_14662),
		.dout(new_net_14663)
	);

	bfr new_net_14664_bfr_after (
		.din(new_net_14663),
		.dout(new_net_14664)
	);

	bfr new_net_14665_bfr_after (
		.din(new_net_14664),
		.dout(new_net_14665)
	);

	bfr new_net_14666_bfr_after (
		.din(new_net_14665),
		.dout(new_net_14666)
	);

	bfr new_net_14667_bfr_after (
		.din(new_net_14666),
		.dout(new_net_14667)
	);

	bfr new_net_14668_bfr_after (
		.din(new_net_14667),
		.dout(new_net_14668)
	);

	bfr new_net_14669_bfr_after (
		.din(new_net_14668),
		.dout(new_net_14669)
	);

	bfr new_net_14670_bfr_after (
		.din(new_net_14669),
		.dout(new_net_14670)
	);

	bfr new_net_14671_bfr_after (
		.din(new_net_14670),
		.dout(new_net_14671)
	);

	bfr new_net_14672_bfr_after (
		.din(new_net_14671),
		.dout(new_net_14672)
	);

	bfr new_net_14673_bfr_after (
		.din(new_net_14672),
		.dout(new_net_14673)
	);

	bfr new_net_14674_bfr_after (
		.din(new_net_14673),
		.dout(new_net_14674)
	);

	bfr new_net_14675_bfr_after (
		.din(new_net_14674),
		.dout(new_net_14675)
	);

	bfr new_net_14676_bfr_after (
		.din(new_net_14675),
		.dout(new_net_14676)
	);

	bfr new_net_14677_bfr_after (
		.din(new_net_14676),
		.dout(new_net_14677)
	);

	bfr new_net_14678_bfr_after (
		.din(new_net_14677),
		.dout(new_net_14678)
	);

	bfr new_net_14679_bfr_after (
		.din(new_net_14678),
		.dout(new_net_14679)
	);

	bfr new_net_14680_bfr_after (
		.din(new_net_14679),
		.dout(new_net_14680)
	);

	bfr new_net_14681_bfr_after (
		.din(new_net_14680),
		.dout(new_net_14681)
	);

	bfr new_net_14682_bfr_after (
		.din(new_net_14681),
		.dout(new_net_14682)
	);

	bfr new_net_14683_bfr_after (
		.din(new_net_14682),
		.dout(new_net_14683)
	);

	bfr new_net_14684_bfr_after (
		.din(new_net_14683),
		.dout(new_net_14684)
	);

	bfr new_net_14685_bfr_after (
		.din(new_net_14684),
		.dout(new_net_14685)
	);

	bfr new_net_14686_bfr_after (
		.din(new_net_14685),
		.dout(new_net_14686)
	);

	bfr new_net_14687_bfr_after (
		.din(new_net_14686),
		.dout(new_net_14687)
	);

	bfr new_net_14688_bfr_after (
		.din(new_net_14687),
		.dout(new_net_14688)
	);

	bfr new_net_14689_bfr_after (
		.din(new_net_14688),
		.dout(new_net_14689)
	);

	bfr new_net_14690_bfr_after (
		.din(new_net_14689),
		.dout(new_net_14690)
	);

	bfr new_net_14691_bfr_after (
		.din(new_net_14690),
		.dout(new_net_14691)
	);

	bfr new_net_14692_bfr_after (
		.din(new_net_14691),
		.dout(new_net_14692)
	);

	bfr new_net_14693_bfr_after (
		.din(new_net_14692),
		.dout(new_net_14693)
	);

	bfr new_net_14694_bfr_after (
		.din(new_net_14693),
		.dout(new_net_14694)
	);

	bfr new_net_14695_bfr_after (
		.din(new_net_14694),
		.dout(new_net_14695)
	);

	bfr new_net_14696_bfr_after (
		.din(new_net_14695),
		.dout(new_net_14696)
	);

	bfr new_net_14697_bfr_after (
		.din(new_net_14696),
		.dout(new_net_14697)
	);

	bfr new_net_14698_bfr_after (
		.din(new_net_14697),
		.dout(new_net_14698)
	);

	bfr new_net_14699_bfr_after (
		.din(new_net_14698),
		.dout(new_net_14699)
	);

	bfr new_net_14700_bfr_after (
		.din(new_net_14699),
		.dout(new_net_14700)
	);

	bfr new_net_14701_bfr_after (
		.din(new_net_14700),
		.dout(new_net_14701)
	);

	bfr new_net_14702_bfr_after (
		.din(new_net_14701),
		.dout(new_net_14702)
	);

	bfr new_net_14703_bfr_after (
		.din(new_net_14702),
		.dout(new_net_14703)
	);

	bfr new_net_14704_bfr_after (
		.din(new_net_14703),
		.dout(new_net_14704)
	);

	bfr new_net_14705_bfr_after (
		.din(new_net_14704),
		.dout(new_net_14705)
	);

	bfr new_net_14706_bfr_after (
		.din(new_net_14705),
		.dout(new_net_14706)
	);

	bfr new_net_14707_bfr_after (
		.din(new_net_14706),
		.dout(new_net_14707)
	);

	bfr new_net_14708_bfr_after (
		.din(new_net_14707),
		.dout(new_net_14708)
	);

	bfr new_net_14709_bfr_after (
		.din(new_net_14708),
		.dout(new_net_14709)
	);

	bfr new_net_14710_bfr_after (
		.din(new_net_14709),
		.dout(new_net_14710)
	);

	bfr new_net_14711_bfr_after (
		.din(new_net_14710),
		.dout(new_net_14711)
	);

	bfr new_net_14712_bfr_after (
		.din(new_net_14711),
		.dout(new_net_14712)
	);

	bfr new_net_14713_bfr_after (
		.din(new_net_14712),
		.dout(new_net_14713)
	);

	bfr new_net_14714_bfr_after (
		.din(new_net_14713),
		.dout(new_net_14714)
	);

	bfr new_net_14715_bfr_after (
		.din(new_net_14714),
		.dout(new_net_14715)
	);

	bfr new_net_14716_bfr_after (
		.din(new_net_14715),
		.dout(new_net_14716)
	);

	bfr new_net_14717_bfr_after (
		.din(new_net_14716),
		.dout(new_net_14717)
	);

	bfr new_net_14718_bfr_after (
		.din(new_net_14717),
		.dout(new_net_14718)
	);

	bfr new_net_14719_bfr_after (
		.din(new_net_14718),
		.dout(new_net_14719)
	);

	bfr new_net_14720_bfr_after (
		.din(new_net_14719),
		.dout(new_net_14720)
	);

	bfr new_net_14721_bfr_after (
		.din(new_net_14720),
		.dout(new_net_14721)
	);

	bfr new_net_14722_bfr_after (
		.din(new_net_14721),
		.dout(new_net_14722)
	);

	bfr new_net_14723_bfr_after (
		.din(new_net_14722),
		.dout(new_net_14723)
	);

	bfr new_net_14724_bfr_after (
		.din(new_net_14723),
		.dout(new_net_14724)
	);

	bfr new_net_14725_bfr_after (
		.din(new_net_14724),
		.dout(new_net_14725)
	);

	bfr new_net_14726_bfr_after (
		.din(new_net_14725),
		.dout(new_net_14726)
	);

	bfr new_net_14727_bfr_after (
		.din(new_net_14726),
		.dout(new_net_14727)
	);

	bfr new_net_14728_bfr_after (
		.din(new_net_14727),
		.dout(new_net_14728)
	);

	bfr new_net_14729_bfr_after (
		.din(new_net_14728),
		.dout(new_net_14729)
	);

	bfr new_net_14730_bfr_after (
		.din(new_net_14729),
		.dout(new_net_14730)
	);

	bfr new_net_14731_bfr_after (
		.din(new_net_14730),
		.dout(new_net_14731)
	);

	bfr new_net_14732_bfr_after (
		.din(new_net_14731),
		.dout(new_net_14732)
	);

	bfr new_net_14733_bfr_after (
		.din(new_net_14732),
		.dout(new_net_14733)
	);

	bfr new_net_14734_bfr_after (
		.din(new_net_14733),
		.dout(new_net_14734)
	);

	bfr new_net_14735_bfr_after (
		.din(new_net_14734),
		.dout(new_net_14735)
	);

	spl2 _0771__v_fanout (
		.a(new_net_14735),
		.b(new_net_984),
		.c(new_net_985)
	);

	bfr new_net_14736_bfr_after (
		.din(_1695_),
		.dout(new_net_14736)
	);

	bfr new_net_14737_bfr_after (
		.din(new_net_14736),
		.dout(new_net_14737)
	);

	bfr new_net_14738_bfr_after (
		.din(new_net_14737),
		.dout(new_net_14738)
	);

	bfr new_net_14739_bfr_after (
		.din(new_net_14738),
		.dout(new_net_14739)
	);

	bfr new_net_14740_bfr_after (
		.din(new_net_14739),
		.dout(new_net_14740)
	);

	bfr new_net_14741_bfr_after (
		.din(new_net_14740),
		.dout(new_net_14741)
	);

	bfr new_net_14742_bfr_after (
		.din(new_net_14741),
		.dout(new_net_14742)
	);

	bfr new_net_14743_bfr_after (
		.din(new_net_14742),
		.dout(new_net_14743)
	);

	bfr new_net_14744_bfr_after (
		.din(new_net_14743),
		.dout(new_net_14744)
	);

	bfr new_net_14745_bfr_after (
		.din(new_net_14744),
		.dout(new_net_14745)
	);

	bfr new_net_14746_bfr_after (
		.din(new_net_14745),
		.dout(new_net_14746)
	);

	bfr new_net_14747_bfr_after (
		.din(new_net_14746),
		.dout(new_net_14747)
	);

	bfr new_net_14748_bfr_after (
		.din(new_net_14747),
		.dout(new_net_14748)
	);

	bfr new_net_14749_bfr_after (
		.din(new_net_14748),
		.dout(new_net_14749)
	);

	bfr new_net_14750_bfr_after (
		.din(new_net_14749),
		.dout(new_net_14750)
	);

	bfr new_net_14751_bfr_after (
		.din(new_net_14750),
		.dout(new_net_14751)
	);

	bfr new_net_14752_bfr_after (
		.din(new_net_14751),
		.dout(new_net_14752)
	);

	bfr new_net_14753_bfr_after (
		.din(new_net_14752),
		.dout(new_net_14753)
	);

	bfr new_net_14754_bfr_after (
		.din(new_net_14753),
		.dout(new_net_14754)
	);

	bfr new_net_14755_bfr_after (
		.din(new_net_14754),
		.dout(new_net_14755)
	);

	bfr new_net_14756_bfr_after (
		.din(new_net_14755),
		.dout(new_net_14756)
	);

	bfr new_net_14757_bfr_after (
		.din(new_net_14756),
		.dout(new_net_14757)
	);

	bfr new_net_14758_bfr_after (
		.din(new_net_14757),
		.dout(new_net_14758)
	);

	bfr new_net_14759_bfr_after (
		.din(new_net_14758),
		.dout(new_net_14759)
	);

	bfr new_net_14760_bfr_after (
		.din(new_net_14759),
		.dout(new_net_14760)
	);

	bfr new_net_14761_bfr_after (
		.din(new_net_14760),
		.dout(new_net_14761)
	);

	bfr new_net_14762_bfr_after (
		.din(new_net_14761),
		.dout(new_net_14762)
	);

	bfr new_net_14763_bfr_after (
		.din(new_net_14762),
		.dout(new_net_14763)
	);

	bfr new_net_14764_bfr_after (
		.din(new_net_14763),
		.dout(new_net_14764)
	);

	bfr new_net_14765_bfr_after (
		.din(new_net_14764),
		.dout(new_net_14765)
	);

	bfr new_net_14766_bfr_after (
		.din(new_net_14765),
		.dout(new_net_14766)
	);

	bfr new_net_14767_bfr_after (
		.din(new_net_14766),
		.dout(new_net_14767)
	);

	bfr new_net_14768_bfr_after (
		.din(new_net_14767),
		.dout(new_net_14768)
	);

	bfr new_net_14769_bfr_after (
		.din(new_net_14768),
		.dout(new_net_14769)
	);

	bfr new_net_14770_bfr_after (
		.din(new_net_14769),
		.dout(new_net_14770)
	);

	bfr new_net_14771_bfr_after (
		.din(new_net_14770),
		.dout(new_net_14771)
	);

	bfr new_net_14772_bfr_after (
		.din(new_net_14771),
		.dout(new_net_14772)
	);

	bfr new_net_14773_bfr_after (
		.din(new_net_14772),
		.dout(new_net_14773)
	);

	bfr new_net_14774_bfr_after (
		.din(new_net_14773),
		.dout(new_net_14774)
	);

	bfr new_net_14775_bfr_after (
		.din(new_net_14774),
		.dout(new_net_14775)
	);

	bfr new_net_14776_bfr_after (
		.din(new_net_14775),
		.dout(new_net_14776)
	);

	bfr new_net_14777_bfr_after (
		.din(new_net_14776),
		.dout(new_net_14777)
	);

	bfr new_net_14778_bfr_after (
		.din(new_net_14777),
		.dout(new_net_14778)
	);

	bfr new_net_14779_bfr_after (
		.din(new_net_14778),
		.dout(new_net_14779)
	);

	bfr new_net_14780_bfr_after (
		.din(new_net_14779),
		.dout(new_net_14780)
	);

	bfr new_net_14781_bfr_after (
		.din(new_net_14780),
		.dout(new_net_14781)
	);

	bfr new_net_14782_bfr_after (
		.din(new_net_14781),
		.dout(new_net_14782)
	);

	bfr new_net_14783_bfr_after (
		.din(new_net_14782),
		.dout(new_net_14783)
	);

	spl2 _1695__v_fanout (
		.a(new_net_14783),
		.b(new_net_2975),
		.c(new_net_2976)
	);

	bfr new_net_14784_bfr_after (
		.din(_0709_),
		.dout(new_net_14784)
	);

	bfr new_net_14785_bfr_after (
		.din(new_net_14784),
		.dout(new_net_14785)
	);

	bfr new_net_14786_bfr_after (
		.din(new_net_14785),
		.dout(new_net_14786)
	);

	bfr new_net_14787_bfr_after (
		.din(new_net_14786),
		.dout(new_net_14787)
	);

	bfr new_net_14788_bfr_after (
		.din(new_net_14787),
		.dout(new_net_14788)
	);

	bfr new_net_14789_bfr_after (
		.din(new_net_14788),
		.dout(new_net_14789)
	);

	bfr new_net_14790_bfr_after (
		.din(new_net_14789),
		.dout(new_net_14790)
	);

	bfr new_net_14791_bfr_after (
		.din(new_net_14790),
		.dout(new_net_14791)
	);

	bfr new_net_14792_bfr_after (
		.din(new_net_14791),
		.dout(new_net_14792)
	);

	bfr new_net_14793_bfr_after (
		.din(new_net_14792),
		.dout(new_net_14793)
	);

	bfr new_net_14794_bfr_after (
		.din(new_net_14793),
		.dout(new_net_14794)
	);

	bfr new_net_14795_bfr_after (
		.din(new_net_14794),
		.dout(new_net_14795)
	);

	bfr new_net_14796_bfr_after (
		.din(new_net_14795),
		.dout(new_net_14796)
	);

	bfr new_net_14797_bfr_after (
		.din(new_net_14796),
		.dout(new_net_14797)
	);

	bfr new_net_14798_bfr_after (
		.din(new_net_14797),
		.dout(new_net_14798)
	);

	bfr new_net_14799_bfr_after (
		.din(new_net_14798),
		.dout(new_net_14799)
	);

	spl2 _0709__v_fanout (
		.a(new_net_14799),
		.b(new_net_868),
		.c(new_net_869)
	);

	bfr new_net_14800_bfr_after (
		.din(_1219_),
		.dout(new_net_14800)
	);

	bfr new_net_14801_bfr_after (
		.din(new_net_14800),
		.dout(new_net_14801)
	);

	bfr new_net_14802_bfr_after (
		.din(new_net_14801),
		.dout(new_net_14802)
	);

	bfr new_net_14803_bfr_after (
		.din(new_net_14802),
		.dout(new_net_14803)
	);

	bfr new_net_14804_bfr_after (
		.din(new_net_14803),
		.dout(new_net_14804)
	);

	bfr new_net_14805_bfr_after (
		.din(new_net_14804),
		.dout(new_net_14805)
	);

	bfr new_net_14806_bfr_after (
		.din(new_net_14805),
		.dout(new_net_14806)
	);

	bfr new_net_14807_bfr_after (
		.din(new_net_14806),
		.dout(new_net_14807)
	);

	spl2 _1219__v_fanout (
		.a(new_net_14807),
		.b(new_net_1082),
		.c(new_net_1083)
	);

	bfr new_net_14808_bfr_before (
		.din(new_net_14808),
		.dout(N545)
	);

	bfr new_net_14809_bfr_before (
		.din(new_net_14809),
		.dout(new_net_14808)
	);

	bfr new_net_14810_bfr_before (
		.din(new_net_14810),
		.dout(new_net_14809)
	);

	bfr new_net_14811_bfr_before (
		.din(new_net_14811),
		.dout(new_net_14810)
	);

	bfr new_net_14812_bfr_before (
		.din(new_net_14812),
		.dout(new_net_14811)
	);

	bfr new_net_14813_bfr_before (
		.din(new_net_14813),
		.dout(new_net_14812)
	);

	bfr new_net_14814_bfr_before (
		.din(new_net_14814),
		.dout(new_net_14813)
	);

	bfr new_net_14815_bfr_before (
		.din(new_net_14815),
		.dout(new_net_14814)
	);

	bfr new_net_14816_bfr_before (
		.din(new_net_14816),
		.dout(new_net_14815)
	);

	bfr new_net_14817_bfr_before (
		.din(new_net_14817),
		.dout(new_net_14816)
	);

	bfr new_net_14818_bfr_before (
		.din(new_net_14818),
		.dout(new_net_14817)
	);

	bfr new_net_14819_bfr_before (
		.din(new_net_14819),
		.dout(new_net_14818)
	);

	bfr new_net_14820_bfr_before (
		.din(new_net_14820),
		.dout(new_net_14819)
	);

	bfr new_net_14821_bfr_before (
		.din(new_net_14821),
		.dout(new_net_14820)
	);

	bfr new_net_14822_bfr_before (
		.din(new_net_14822),
		.dout(new_net_14821)
	);

	bfr new_net_14823_bfr_before (
		.din(new_net_14823),
		.dout(new_net_14822)
	);

	bfr new_net_14824_bfr_before (
		.din(new_net_14824),
		.dout(new_net_14823)
	);

	bfr new_net_14825_bfr_before (
		.din(new_net_14825),
		.dout(new_net_14824)
	);

	bfr new_net_14826_bfr_before (
		.din(new_net_14826),
		.dout(new_net_14825)
	);

	bfr new_net_14827_bfr_before (
		.din(new_net_14827),
		.dout(new_net_14826)
	);

	bfr new_net_14828_bfr_before (
		.din(new_net_14828),
		.dout(new_net_14827)
	);

	bfr new_net_14829_bfr_before (
		.din(new_net_14829),
		.dout(new_net_14828)
	);

	bfr new_net_14830_bfr_before (
		.din(new_net_14830),
		.dout(new_net_14829)
	);

	bfr new_net_14831_bfr_before (
		.din(new_net_14831),
		.dout(new_net_14830)
	);

	bfr new_net_14832_bfr_before (
		.din(new_net_14832),
		.dout(new_net_14831)
	);

	bfr new_net_14833_bfr_before (
		.din(new_net_14833),
		.dout(new_net_14832)
	);

	bfr new_net_14834_bfr_before (
		.din(new_net_14834),
		.dout(new_net_14833)
	);

	bfr new_net_14835_bfr_before (
		.din(new_net_14835),
		.dout(new_net_14834)
	);

	bfr new_net_14836_bfr_before (
		.din(new_net_14836),
		.dout(new_net_14835)
	);

	bfr new_net_14837_bfr_before (
		.din(new_net_14837),
		.dout(new_net_14836)
	);

	bfr new_net_14838_bfr_before (
		.din(new_net_14838),
		.dout(new_net_14837)
	);

	bfr new_net_14839_bfr_before (
		.din(new_net_14839),
		.dout(new_net_14838)
	);

	bfr new_net_14840_bfr_before (
		.din(new_net_14840),
		.dout(new_net_14839)
	);

	bfr new_net_14841_bfr_before (
		.din(new_net_14841),
		.dout(new_net_14840)
	);

	bfr new_net_14842_bfr_before (
		.din(new_net_14842),
		.dout(new_net_14841)
	);

	bfr new_net_14843_bfr_before (
		.din(new_net_14843),
		.dout(new_net_14842)
	);

	bfr new_net_14844_bfr_before (
		.din(new_net_14844),
		.dout(new_net_14843)
	);

	bfr new_net_14845_bfr_before (
		.din(new_net_14845),
		.dout(new_net_14844)
	);

	bfr new_net_14846_bfr_before (
		.din(new_net_14846),
		.dout(new_net_14845)
	);

	bfr new_net_14847_bfr_before (
		.din(new_net_14847),
		.dout(new_net_14846)
	);

	bfr new_net_14848_bfr_before (
		.din(new_net_14848),
		.dout(new_net_14847)
	);

	bfr new_net_14849_bfr_before (
		.din(new_net_14849),
		.dout(new_net_14848)
	);

	bfr new_net_14850_bfr_before (
		.din(new_net_14850),
		.dout(new_net_14849)
	);

	bfr new_net_14851_bfr_before (
		.din(new_net_14851),
		.dout(new_net_14850)
	);

	bfr new_net_14852_bfr_before (
		.din(new_net_14852),
		.dout(new_net_14851)
	);

	bfr new_net_14853_bfr_before (
		.din(new_net_14853),
		.dout(new_net_14852)
	);

	bfr new_net_14854_bfr_before (
		.din(new_net_14854),
		.dout(new_net_14853)
	);

	bfr new_net_14855_bfr_before (
		.din(new_net_14855),
		.dout(new_net_14854)
	);

	bfr new_net_14856_bfr_before (
		.din(new_net_14856),
		.dout(new_net_14855)
	);

	bfr new_net_14857_bfr_before (
		.din(new_net_14857),
		.dout(new_net_14856)
	);

	bfr new_net_14858_bfr_before (
		.din(new_net_14858),
		.dout(new_net_14857)
	);

	bfr new_net_14859_bfr_before (
		.din(new_net_14859),
		.dout(new_net_14858)
	);

	bfr new_net_14860_bfr_before (
		.din(new_net_14860),
		.dout(new_net_14859)
	);

	bfr new_net_14861_bfr_before (
		.din(new_net_14861),
		.dout(new_net_14860)
	);

	bfr new_net_14862_bfr_before (
		.din(new_net_14862),
		.dout(new_net_14861)
	);

	bfr new_net_14863_bfr_before (
		.din(new_net_14863),
		.dout(new_net_14862)
	);

	bfr new_net_14864_bfr_before (
		.din(new_net_14864),
		.dout(new_net_14863)
	);

	bfr new_net_14865_bfr_before (
		.din(new_net_14865),
		.dout(new_net_14864)
	);

	bfr new_net_14866_bfr_before (
		.din(new_net_14866),
		.dout(new_net_14865)
	);

	bfr new_net_14867_bfr_before (
		.din(new_net_14867),
		.dout(new_net_14866)
	);

	bfr new_net_14868_bfr_before (
		.din(new_net_14868),
		.dout(new_net_14867)
	);

	bfr new_net_14869_bfr_before (
		.din(new_net_14869),
		.dout(new_net_14868)
	);

	bfr new_net_14870_bfr_before (
		.din(new_net_14870),
		.dout(new_net_14869)
	);

	bfr new_net_14871_bfr_before (
		.din(new_net_14871),
		.dout(new_net_14870)
	);

	bfr new_net_14872_bfr_before (
		.din(new_net_14872),
		.dout(new_net_14871)
	);

	bfr new_net_14873_bfr_before (
		.din(new_net_14873),
		.dout(new_net_14872)
	);

	bfr new_net_14874_bfr_before (
		.din(new_net_14874),
		.dout(new_net_14873)
	);

	bfr new_net_14875_bfr_before (
		.din(new_net_14875),
		.dout(new_net_14874)
	);

	bfr new_net_14876_bfr_before (
		.din(new_net_14876),
		.dout(new_net_14875)
	);

	bfr new_net_14877_bfr_before (
		.din(new_net_14877),
		.dout(new_net_14876)
	);

	bfr new_net_14878_bfr_before (
		.din(new_net_14878),
		.dout(new_net_14877)
	);

	bfr new_net_14879_bfr_before (
		.din(new_net_14879),
		.dout(new_net_14878)
	);

	bfr new_net_14880_bfr_before (
		.din(new_net_14880),
		.dout(new_net_14879)
	);

	bfr new_net_14881_bfr_before (
		.din(new_net_14881),
		.dout(new_net_14880)
	);

	bfr new_net_14882_bfr_before (
		.din(new_net_14882),
		.dout(new_net_14881)
	);

	bfr new_net_14883_bfr_before (
		.din(new_net_14883),
		.dout(new_net_14882)
	);

	bfr new_net_14884_bfr_before (
		.din(new_net_14884),
		.dout(new_net_14883)
	);

	bfr new_net_14885_bfr_before (
		.din(new_net_14885),
		.dout(new_net_14884)
	);

	bfr new_net_14886_bfr_before (
		.din(new_net_14886),
		.dout(new_net_14885)
	);

	bfr new_net_14887_bfr_before (
		.din(new_net_14887),
		.dout(new_net_14886)
	);

	bfr new_net_14888_bfr_before (
		.din(new_net_14888),
		.dout(new_net_14887)
	);

	bfr new_net_14889_bfr_before (
		.din(new_net_14889),
		.dout(new_net_14888)
	);

	bfr new_net_14890_bfr_before (
		.din(new_net_14890),
		.dout(new_net_14889)
	);

	bfr new_net_14891_bfr_before (
		.din(new_net_14891),
		.dout(new_net_14890)
	);

	bfr new_net_14892_bfr_before (
		.din(new_net_14892),
		.dout(new_net_14891)
	);

	bfr new_net_14893_bfr_before (
		.din(new_net_14893),
		.dout(new_net_14892)
	);

	bfr new_net_14894_bfr_before (
		.din(new_net_14894),
		.dout(new_net_14893)
	);

	bfr new_net_14895_bfr_before (
		.din(new_net_14895),
		.dout(new_net_14894)
	);

	bfr new_net_14896_bfr_before (
		.din(new_net_14896),
		.dout(new_net_14895)
	);

	bfr new_net_14897_bfr_before (
		.din(new_net_14897),
		.dout(new_net_14896)
	);

	bfr new_net_14898_bfr_before (
		.din(new_net_14898),
		.dout(new_net_14897)
	);

	bfr new_net_14899_bfr_before (
		.din(new_net_14899),
		.dout(new_net_14898)
	);

	bfr new_net_14900_bfr_before (
		.din(new_net_14900),
		.dout(new_net_14899)
	);

	bfr new_net_14901_bfr_before (
		.din(new_net_14901),
		.dout(new_net_14900)
	);

	bfr new_net_14902_bfr_before (
		.din(new_net_14902),
		.dout(new_net_14901)
	);

	bfr new_net_14903_bfr_before (
		.din(new_net_14903),
		.dout(new_net_14902)
	);

	bfr new_net_14904_bfr_before (
		.din(new_net_14904),
		.dout(new_net_14903)
	);

	bfr new_net_14905_bfr_before (
		.din(new_net_14905),
		.dout(new_net_14904)
	);

	bfr new_net_14906_bfr_before (
		.din(new_net_14906),
		.dout(new_net_14905)
	);

	bfr new_net_14907_bfr_before (
		.din(new_net_14907),
		.dout(new_net_14906)
	);

	bfr new_net_14908_bfr_before (
		.din(new_net_14908),
		.dout(new_net_14907)
	);

	bfr new_net_14909_bfr_before (
		.din(new_net_14909),
		.dout(new_net_14908)
	);

	bfr new_net_14910_bfr_before (
		.din(new_net_14910),
		.dout(new_net_14909)
	);

	bfr new_net_14911_bfr_before (
		.din(new_net_14911),
		.dout(new_net_14910)
	);

	bfr new_net_14912_bfr_before (
		.din(new_net_14912),
		.dout(new_net_14911)
	);

	bfr new_net_14913_bfr_before (
		.din(new_net_14913),
		.dout(new_net_14912)
	);

	bfr new_net_14914_bfr_before (
		.din(new_net_14914),
		.dout(new_net_14913)
	);

	bfr new_net_14915_bfr_before (
		.din(new_net_14915),
		.dout(new_net_14914)
	);

	bfr new_net_14916_bfr_before (
		.din(new_net_14916),
		.dout(new_net_14915)
	);

	bfr new_net_14917_bfr_before (
		.din(new_net_14917),
		.dout(new_net_14916)
	);

	bfr new_net_14918_bfr_before (
		.din(new_net_14918),
		.dout(new_net_14917)
	);

	bfr new_net_14919_bfr_before (
		.din(new_net_14919),
		.dout(new_net_14918)
	);

	bfr new_net_14920_bfr_before (
		.din(new_net_14920),
		.dout(new_net_14919)
	);

	bfr new_net_14921_bfr_before (
		.din(new_net_14921),
		.dout(new_net_14920)
	);

	bfr new_net_14922_bfr_before (
		.din(new_net_14922),
		.dout(new_net_14921)
	);

	bfr new_net_14923_bfr_before (
		.din(new_net_14923),
		.dout(new_net_14922)
	);

	bfr new_net_14924_bfr_before (
		.din(new_net_14924),
		.dout(new_net_14923)
	);

	bfr new_net_14925_bfr_before (
		.din(new_net_14925),
		.dout(new_net_14924)
	);

	bfr new_net_14926_bfr_before (
		.din(new_net_14926),
		.dout(new_net_14925)
	);

	bfr new_net_14927_bfr_before (
		.din(new_net_14927),
		.dout(new_net_14926)
	);

	bfr new_net_14928_bfr_before (
		.din(new_net_14928),
		.dout(new_net_14927)
	);

	bfr new_net_14929_bfr_before (
		.din(new_net_14929),
		.dout(new_net_14928)
	);

	bfr new_net_14930_bfr_before (
		.din(new_net_14930),
		.dout(new_net_14929)
	);

	bfr new_net_14931_bfr_before (
		.din(new_net_14931),
		.dout(new_net_14930)
	);

	bfr new_net_14932_bfr_before (
		.din(new_net_14932),
		.dout(new_net_14931)
	);

	bfr new_net_14933_bfr_before (
		.din(new_net_14933),
		.dout(new_net_14932)
	);

	bfr new_net_14934_bfr_before (
		.din(new_net_14934),
		.dout(new_net_14933)
	);

	bfr new_net_14935_bfr_before (
		.din(new_net_14935),
		.dout(new_net_14934)
	);

	bfr new_net_14936_bfr_before (
		.din(new_net_14936),
		.dout(new_net_14935)
	);

	bfr new_net_14937_bfr_before (
		.din(new_net_14937),
		.dout(new_net_14936)
	);

	bfr new_net_14938_bfr_before (
		.din(new_net_14938),
		.dout(new_net_14937)
	);

	bfr new_net_14939_bfr_before (
		.din(new_net_14939),
		.dout(new_net_14938)
	);

	bfr new_net_14940_bfr_before (
		.din(new_net_14940),
		.dout(new_net_14939)
	);

	bfr new_net_14941_bfr_before (
		.din(new_net_14941),
		.dout(new_net_14940)
	);

	bfr new_net_14942_bfr_before (
		.din(new_net_14942),
		.dout(new_net_14941)
	);

	bfr new_net_14943_bfr_before (
		.din(new_net_14943),
		.dout(new_net_14942)
	);

	bfr new_net_14944_bfr_before (
		.din(new_net_14944),
		.dout(new_net_14943)
	);

	bfr new_net_14945_bfr_before (
		.din(new_net_14945),
		.dout(new_net_14944)
	);

	bfr new_net_14946_bfr_before (
		.din(new_net_14946),
		.dout(new_net_14945)
	);

	bfr new_net_14947_bfr_before (
		.din(new_net_14947),
		.dout(new_net_14946)
	);

	bfr new_net_14948_bfr_before (
		.din(new_net_14948),
		.dout(new_net_14947)
	);

	bfr new_net_14949_bfr_before (
		.din(new_net_14949),
		.dout(new_net_14948)
	);

	bfr new_net_14950_bfr_before (
		.din(new_net_14950),
		.dout(new_net_14949)
	);

	bfr new_net_14951_bfr_before (
		.din(new_net_14951),
		.dout(new_net_14950)
	);

	bfr new_net_14952_bfr_before (
		.din(new_net_14952),
		.dout(new_net_14951)
	);

	bfr new_net_14953_bfr_before (
		.din(new_net_14953),
		.dout(new_net_14952)
	);

	bfr new_net_14954_bfr_before (
		.din(new_net_14954),
		.dout(new_net_14953)
	);

	bfr new_net_14955_bfr_before (
		.din(new_net_14955),
		.dout(new_net_14954)
	);

	bfr new_net_14956_bfr_before (
		.din(new_net_14956),
		.dout(new_net_14955)
	);

	bfr new_net_14957_bfr_before (
		.din(new_net_14957),
		.dout(new_net_14956)
	);

	bfr new_net_14958_bfr_before (
		.din(new_net_14958),
		.dout(new_net_14957)
	);

	bfr new_net_14959_bfr_before (
		.din(new_net_14959),
		.dout(new_net_14958)
	);

	bfr new_net_14960_bfr_before (
		.din(new_net_14960),
		.dout(new_net_14959)
	);

	bfr new_net_14961_bfr_before (
		.din(new_net_14961),
		.dout(new_net_14960)
	);

	bfr new_net_14962_bfr_before (
		.din(new_net_14962),
		.dout(new_net_14961)
	);

	bfr new_net_14963_bfr_before (
		.din(new_net_14963),
		.dout(new_net_14962)
	);

	bfr new_net_14964_bfr_before (
		.din(new_net_14964),
		.dout(new_net_14963)
	);

	bfr new_net_14965_bfr_before (
		.din(new_net_14965),
		.dout(new_net_14964)
	);

	bfr new_net_14966_bfr_before (
		.din(new_net_14966),
		.dout(new_net_14965)
	);

	bfr new_net_14967_bfr_before (
		.din(new_net_14967),
		.dout(new_net_14966)
	);

	bfr new_net_14968_bfr_before (
		.din(new_net_14968),
		.dout(new_net_14967)
	);

	bfr new_net_14969_bfr_before (
		.din(new_net_14969),
		.dout(new_net_14968)
	);

	bfr new_net_14970_bfr_before (
		.din(new_net_14970),
		.dout(new_net_14969)
	);

	bfr new_net_14971_bfr_before (
		.din(new_net_14971),
		.dout(new_net_14970)
	);

	bfr new_net_14972_bfr_before (
		.din(new_net_14972),
		.dout(new_net_14971)
	);

	bfr new_net_14973_bfr_before (
		.din(new_net_14973),
		.dout(new_net_14972)
	);

	bfr new_net_14974_bfr_before (
		.din(new_net_14974),
		.dout(new_net_14973)
	);

	bfr new_net_14975_bfr_before (
		.din(new_net_14975),
		.dout(new_net_14974)
	);

	bfr new_net_14976_bfr_before (
		.din(new_net_14976),
		.dout(new_net_14975)
	);

	bfr new_net_14977_bfr_before (
		.din(new_net_14977),
		.dout(new_net_14976)
	);

	bfr new_net_14978_bfr_before (
		.din(new_net_14978),
		.dout(new_net_14977)
	);

	bfr new_net_14979_bfr_before (
		.din(new_net_14979),
		.dout(new_net_14978)
	);

	bfr new_net_14980_bfr_before (
		.din(new_net_14980),
		.dout(new_net_14979)
	);

	bfr new_net_14981_bfr_before (
		.din(new_net_14981),
		.dout(new_net_14980)
	);

	bfr new_net_14982_bfr_before (
		.din(new_net_14982),
		.dout(new_net_14981)
	);

	spl2 new_net_0_v_fanout (
		.a(new_net_0),
		.b(new_net_14982),
		.c(new_net_1195)
	);

	spl2 _1085__v_fanout (
		.a(_1085_),
		.b(new_net_2621),
		.c(new_net_2622)
	);

	bfr new_net_14983_bfr_after (
		.din(_1296_),
		.dout(new_net_14983)
	);

	bfr new_net_14984_bfr_after (
		.din(new_net_14983),
		.dout(new_net_14984)
	);

	bfr new_net_14985_bfr_after (
		.din(new_net_14984),
		.dout(new_net_14985)
	);

	bfr new_net_14986_bfr_after (
		.din(new_net_14985),
		.dout(new_net_14986)
	);

	bfr new_net_14987_bfr_after (
		.din(new_net_14986),
		.dout(new_net_14987)
	);

	bfr new_net_14988_bfr_after (
		.din(new_net_14987),
		.dout(new_net_14988)
	);

	bfr new_net_14989_bfr_after (
		.din(new_net_14988),
		.dout(new_net_14989)
	);

	bfr new_net_14990_bfr_after (
		.din(new_net_14989),
		.dout(new_net_14990)
	);

	spl2 _1296__v_fanout (
		.a(new_net_14990),
		.b(new_net_874),
		.c(new_net_875)
	);

	bfr new_net_14991_bfr_after (
		.din(_0318_),
		.dout(new_net_14991)
	);

	bfr new_net_14992_bfr_after (
		.din(new_net_14991),
		.dout(new_net_14992)
	);

	bfr new_net_14993_bfr_after (
		.din(new_net_14992),
		.dout(new_net_14993)
	);

	bfr new_net_14994_bfr_after (
		.din(new_net_14993),
		.dout(new_net_14994)
	);

	bfr new_net_14995_bfr_after (
		.din(new_net_14994),
		.dout(new_net_14995)
	);

	bfr new_net_14996_bfr_after (
		.din(new_net_14995),
		.dout(new_net_14996)
	);

	bfr new_net_14997_bfr_after (
		.din(new_net_14996),
		.dout(new_net_14997)
	);

	bfr new_net_14998_bfr_after (
		.din(new_net_14997),
		.dout(new_net_14998)
	);

	bfr new_net_14999_bfr_after (
		.din(new_net_14998),
		.dout(new_net_14999)
	);

	bfr new_net_15000_bfr_after (
		.din(new_net_14999),
		.dout(new_net_15000)
	);

	bfr new_net_15001_bfr_after (
		.din(new_net_15000),
		.dout(new_net_15001)
	);

	bfr new_net_15002_bfr_after (
		.din(new_net_15001),
		.dout(new_net_15002)
	);

	bfr new_net_15003_bfr_after (
		.din(new_net_15002),
		.dout(new_net_15003)
	);

	bfr new_net_15004_bfr_after (
		.din(new_net_15003),
		.dout(new_net_15004)
	);

	bfr new_net_15005_bfr_after (
		.din(new_net_15004),
		.dout(new_net_15005)
	);

	bfr new_net_15006_bfr_after (
		.din(new_net_15005),
		.dout(new_net_15006)
	);

	spl2 _0318__v_fanout (
		.a(new_net_15006),
		.b(new_net_287),
		.c(new_net_288)
	);

	bfr new_net_15007_bfr_after (
		.din(_0666_),
		.dout(new_net_15007)
	);

	bfr new_net_15008_bfr_after (
		.din(new_net_15007),
		.dout(new_net_15008)
	);

	bfr new_net_15009_bfr_after (
		.din(new_net_15008),
		.dout(new_net_15009)
	);

	bfr new_net_15010_bfr_after (
		.din(new_net_15009),
		.dout(new_net_15010)
	);

	bfr new_net_15011_bfr_after (
		.din(new_net_15010),
		.dout(new_net_15011)
	);

	bfr new_net_15012_bfr_after (
		.din(new_net_15011),
		.dout(new_net_15012)
	);

	bfr new_net_15013_bfr_after (
		.din(new_net_15012),
		.dout(new_net_15013)
	);

	bfr new_net_15014_bfr_after (
		.din(new_net_15013),
		.dout(new_net_15014)
	);

	bfr new_net_15015_bfr_after (
		.din(new_net_15014),
		.dout(new_net_15015)
	);

	bfr new_net_15016_bfr_after (
		.din(new_net_15015),
		.dout(new_net_15016)
	);

	bfr new_net_15017_bfr_after (
		.din(new_net_15016),
		.dout(new_net_15017)
	);

	bfr new_net_15018_bfr_after (
		.din(new_net_15017),
		.dout(new_net_15018)
	);

	bfr new_net_15019_bfr_after (
		.din(new_net_15018),
		.dout(new_net_15019)
	);

	bfr new_net_15020_bfr_after (
		.din(new_net_15019),
		.dout(new_net_15020)
	);

	bfr new_net_15021_bfr_after (
		.din(new_net_15020),
		.dout(new_net_15021)
	);

	bfr new_net_15022_bfr_after (
		.din(new_net_15021),
		.dout(new_net_15022)
	);

	bfr new_net_15023_bfr_after (
		.din(new_net_15022),
		.dout(new_net_15023)
	);

	bfr new_net_15024_bfr_after (
		.din(new_net_15023),
		.dout(new_net_15024)
	);

	bfr new_net_15025_bfr_after (
		.din(new_net_15024),
		.dout(new_net_15025)
	);

	bfr new_net_15026_bfr_after (
		.din(new_net_15025),
		.dout(new_net_15026)
	);

	bfr new_net_15027_bfr_after (
		.din(new_net_15026),
		.dout(new_net_15027)
	);

	bfr new_net_15028_bfr_after (
		.din(new_net_15027),
		.dout(new_net_15028)
	);

	bfr new_net_15029_bfr_after (
		.din(new_net_15028),
		.dout(new_net_15029)
	);

	bfr new_net_15030_bfr_after (
		.din(new_net_15029),
		.dout(new_net_15030)
	);

	bfr new_net_15031_bfr_after (
		.din(new_net_15030),
		.dout(new_net_15031)
	);

	bfr new_net_15032_bfr_after (
		.din(new_net_15031),
		.dout(new_net_15032)
	);

	bfr new_net_15033_bfr_after (
		.din(new_net_15032),
		.dout(new_net_15033)
	);

	bfr new_net_15034_bfr_after (
		.din(new_net_15033),
		.dout(new_net_15034)
	);

	bfr new_net_15035_bfr_after (
		.din(new_net_15034),
		.dout(new_net_15035)
	);

	bfr new_net_15036_bfr_after (
		.din(new_net_15035),
		.dout(new_net_15036)
	);

	bfr new_net_15037_bfr_after (
		.din(new_net_15036),
		.dout(new_net_15037)
	);

	bfr new_net_15038_bfr_after (
		.din(new_net_15037),
		.dout(new_net_15038)
	);

	spl2 _0666__v_fanout (
		.a(new_net_15038),
		.b(new_net_327),
		.c(new_net_328)
	);

	bfr new_net_15039_bfr_after (
		.din(_1821_),
		.dout(new_net_15039)
	);

	bfr new_net_15040_bfr_after (
		.din(new_net_15039),
		.dout(new_net_15040)
	);

	bfr new_net_15041_bfr_after (
		.din(new_net_15040),
		.dout(new_net_15041)
	);

	bfr new_net_15042_bfr_after (
		.din(new_net_15041),
		.dout(new_net_15042)
	);

	bfr new_net_15043_bfr_after (
		.din(new_net_15042),
		.dout(new_net_15043)
	);

	bfr new_net_15044_bfr_after (
		.din(new_net_15043),
		.dout(new_net_15044)
	);

	bfr new_net_15045_bfr_after (
		.din(new_net_15044),
		.dout(new_net_15045)
	);

	bfr new_net_15046_bfr_after (
		.din(new_net_15045),
		.dout(new_net_15046)
	);

	bfr new_net_15047_bfr_after (
		.din(new_net_15046),
		.dout(new_net_15047)
	);

	bfr new_net_15048_bfr_after (
		.din(new_net_15047),
		.dout(new_net_15048)
	);

	bfr new_net_15049_bfr_after (
		.din(new_net_15048),
		.dout(new_net_15049)
	);

	bfr new_net_15050_bfr_after (
		.din(new_net_15049),
		.dout(new_net_15050)
	);

	bfr new_net_15051_bfr_after (
		.din(new_net_15050),
		.dout(new_net_15051)
	);

	bfr new_net_15052_bfr_after (
		.din(new_net_15051),
		.dout(new_net_15052)
	);

	bfr new_net_15053_bfr_after (
		.din(new_net_15052),
		.dout(new_net_15053)
	);

	bfr new_net_15054_bfr_after (
		.din(new_net_15053),
		.dout(new_net_15054)
	);

	bfr new_net_15055_bfr_after (
		.din(new_net_15054),
		.dout(new_net_15055)
	);

	bfr new_net_15056_bfr_after (
		.din(new_net_15055),
		.dout(new_net_15056)
	);

	bfr new_net_15057_bfr_after (
		.din(new_net_15056),
		.dout(new_net_15057)
	);

	bfr new_net_15058_bfr_after (
		.din(new_net_15057),
		.dout(new_net_15058)
	);

	bfr new_net_15059_bfr_after (
		.din(new_net_15058),
		.dout(new_net_15059)
	);

	bfr new_net_15060_bfr_after (
		.din(new_net_15059),
		.dout(new_net_15060)
	);

	bfr new_net_15061_bfr_after (
		.din(new_net_15060),
		.dout(new_net_15061)
	);

	bfr new_net_15062_bfr_after (
		.din(new_net_15061),
		.dout(new_net_15062)
	);

	bfr new_net_15063_bfr_after (
		.din(new_net_15062),
		.dout(new_net_15063)
	);

	bfr new_net_15064_bfr_after (
		.din(new_net_15063),
		.dout(new_net_15064)
	);

	bfr new_net_15065_bfr_after (
		.din(new_net_15064),
		.dout(new_net_15065)
	);

	bfr new_net_15066_bfr_after (
		.din(new_net_15065),
		.dout(new_net_15066)
	);

	bfr new_net_15067_bfr_after (
		.din(new_net_15066),
		.dout(new_net_15067)
	);

	bfr new_net_15068_bfr_after (
		.din(new_net_15067),
		.dout(new_net_15068)
	);

	bfr new_net_15069_bfr_after (
		.din(new_net_15068),
		.dout(new_net_15069)
	);

	bfr new_net_15070_bfr_after (
		.din(new_net_15069),
		.dout(new_net_15070)
	);

	bfr new_net_15071_bfr_after (
		.din(new_net_15070),
		.dout(new_net_15071)
	);

	bfr new_net_15072_bfr_after (
		.din(new_net_15071),
		.dout(new_net_15072)
	);

	bfr new_net_15073_bfr_after (
		.din(new_net_15072),
		.dout(new_net_15073)
	);

	bfr new_net_15074_bfr_after (
		.din(new_net_15073),
		.dout(new_net_15074)
	);

	bfr new_net_15075_bfr_after (
		.din(new_net_15074),
		.dout(new_net_15075)
	);

	bfr new_net_15076_bfr_after (
		.din(new_net_15075),
		.dout(new_net_15076)
	);

	bfr new_net_15077_bfr_after (
		.din(new_net_15076),
		.dout(new_net_15077)
	);

	bfr new_net_15078_bfr_after (
		.din(new_net_15077),
		.dout(new_net_15078)
	);

	spl2 _1821__v_fanout (
		.a(new_net_15078),
		.b(new_net_1646),
		.c(new_net_1647)
	);

	bfr new_net_15079_bfr_after (
		.din(_1290_),
		.dout(new_net_15079)
	);

	bfr new_net_15080_bfr_after (
		.din(new_net_15079),
		.dout(new_net_15080)
	);

	bfr new_net_15081_bfr_after (
		.din(new_net_15080),
		.dout(new_net_15081)
	);

	bfr new_net_15082_bfr_after (
		.din(new_net_15081),
		.dout(new_net_15082)
	);

	bfr new_net_15083_bfr_after (
		.din(new_net_15082),
		.dout(new_net_15083)
	);

	bfr new_net_15084_bfr_after (
		.din(new_net_15083),
		.dout(new_net_15084)
	);

	bfr new_net_15085_bfr_after (
		.din(new_net_15084),
		.dout(new_net_15085)
	);

	bfr new_net_15086_bfr_after (
		.din(new_net_15085),
		.dout(new_net_15086)
	);

	bfr new_net_15087_bfr_after (
		.din(new_net_15086),
		.dout(new_net_15087)
	);

	bfr new_net_15088_bfr_after (
		.din(new_net_15087),
		.dout(new_net_15088)
	);

	bfr new_net_15089_bfr_after (
		.din(new_net_15088),
		.dout(new_net_15089)
	);

	bfr new_net_15090_bfr_after (
		.din(new_net_15089),
		.dout(new_net_15090)
	);

	bfr new_net_15091_bfr_after (
		.din(new_net_15090),
		.dout(new_net_15091)
	);

	bfr new_net_15092_bfr_after (
		.din(new_net_15091),
		.dout(new_net_15092)
	);

	bfr new_net_15093_bfr_after (
		.din(new_net_15092),
		.dout(new_net_15093)
	);

	bfr new_net_15094_bfr_after (
		.din(new_net_15093),
		.dout(new_net_15094)
	);

	bfr new_net_15095_bfr_after (
		.din(new_net_15094),
		.dout(new_net_15095)
	);

	bfr new_net_15096_bfr_after (
		.din(new_net_15095),
		.dout(new_net_15096)
	);

	bfr new_net_15097_bfr_after (
		.din(new_net_15096),
		.dout(new_net_15097)
	);

	bfr new_net_15098_bfr_after (
		.din(new_net_15097),
		.dout(new_net_15098)
	);

	bfr new_net_15099_bfr_after (
		.din(new_net_15098),
		.dout(new_net_15099)
	);

	bfr new_net_15100_bfr_after (
		.din(new_net_15099),
		.dout(new_net_15100)
	);

	bfr new_net_15101_bfr_after (
		.din(new_net_15100),
		.dout(new_net_15101)
	);

	bfr new_net_15102_bfr_after (
		.din(new_net_15101),
		.dout(new_net_15102)
	);

	bfr new_net_15103_bfr_after (
		.din(new_net_15102),
		.dout(new_net_15103)
	);

	bfr new_net_15104_bfr_after (
		.din(new_net_15103),
		.dout(new_net_15104)
	);

	bfr new_net_15105_bfr_after (
		.din(new_net_15104),
		.dout(new_net_15105)
	);

	bfr new_net_15106_bfr_after (
		.din(new_net_15105),
		.dout(new_net_15106)
	);

	bfr new_net_15107_bfr_after (
		.din(new_net_15106),
		.dout(new_net_15107)
	);

	bfr new_net_15108_bfr_after (
		.din(new_net_15107),
		.dout(new_net_15108)
	);

	bfr new_net_15109_bfr_after (
		.din(new_net_15108),
		.dout(new_net_15109)
	);

	bfr new_net_15110_bfr_after (
		.din(new_net_15109),
		.dout(new_net_15110)
	);

	spl2 _1290__v_fanout (
		.a(new_net_15110),
		.b(new_net_2274),
		.c(new_net_2275)
	);

	bfr new_net_15111_bfr_after (
		.din(_0773_),
		.dout(new_net_15111)
	);

	bfr new_net_15112_bfr_after (
		.din(new_net_15111),
		.dout(new_net_15112)
	);

	bfr new_net_15113_bfr_after (
		.din(new_net_15112),
		.dout(new_net_15113)
	);

	bfr new_net_15114_bfr_after (
		.din(new_net_15113),
		.dout(new_net_15114)
	);

	bfr new_net_15115_bfr_after (
		.din(new_net_15114),
		.dout(new_net_15115)
	);

	bfr new_net_15116_bfr_after (
		.din(new_net_15115),
		.dout(new_net_15116)
	);

	bfr new_net_15117_bfr_after (
		.din(new_net_15116),
		.dout(new_net_15117)
	);

	bfr new_net_15118_bfr_after (
		.din(new_net_15117),
		.dout(new_net_15118)
	);

	bfr new_net_15119_bfr_after (
		.din(new_net_15118),
		.dout(new_net_15119)
	);

	bfr new_net_15120_bfr_after (
		.din(new_net_15119),
		.dout(new_net_15120)
	);

	bfr new_net_15121_bfr_after (
		.din(new_net_15120),
		.dout(new_net_15121)
	);

	bfr new_net_15122_bfr_after (
		.din(new_net_15121),
		.dout(new_net_15122)
	);

	bfr new_net_15123_bfr_after (
		.din(new_net_15122),
		.dout(new_net_15123)
	);

	bfr new_net_15124_bfr_after (
		.din(new_net_15123),
		.dout(new_net_15124)
	);

	bfr new_net_15125_bfr_after (
		.din(new_net_15124),
		.dout(new_net_15125)
	);

	bfr new_net_15126_bfr_after (
		.din(new_net_15125),
		.dout(new_net_15126)
	);

	bfr new_net_15127_bfr_after (
		.din(new_net_15126),
		.dout(new_net_15127)
	);

	bfr new_net_15128_bfr_after (
		.din(new_net_15127),
		.dout(new_net_15128)
	);

	bfr new_net_15129_bfr_after (
		.din(new_net_15128),
		.dout(new_net_15129)
	);

	bfr new_net_15130_bfr_after (
		.din(new_net_15129),
		.dout(new_net_15130)
	);

	bfr new_net_15131_bfr_after (
		.din(new_net_15130),
		.dout(new_net_15131)
	);

	bfr new_net_15132_bfr_after (
		.din(new_net_15131),
		.dout(new_net_15132)
	);

	bfr new_net_15133_bfr_after (
		.din(new_net_15132),
		.dout(new_net_15133)
	);

	bfr new_net_15134_bfr_after (
		.din(new_net_15133),
		.dout(new_net_15134)
	);

	bfr new_net_15135_bfr_after (
		.din(new_net_15134),
		.dout(new_net_15135)
	);

	bfr new_net_15136_bfr_after (
		.din(new_net_15135),
		.dout(new_net_15136)
	);

	bfr new_net_15137_bfr_after (
		.din(new_net_15136),
		.dout(new_net_15137)
	);

	bfr new_net_15138_bfr_after (
		.din(new_net_15137),
		.dout(new_net_15138)
	);

	bfr new_net_15139_bfr_after (
		.din(new_net_15138),
		.dout(new_net_15139)
	);

	bfr new_net_15140_bfr_after (
		.din(new_net_15139),
		.dout(new_net_15140)
	);

	bfr new_net_15141_bfr_after (
		.din(new_net_15140),
		.dout(new_net_15141)
	);

	bfr new_net_15142_bfr_after (
		.din(new_net_15141),
		.dout(new_net_15142)
	);

	bfr new_net_15143_bfr_after (
		.din(new_net_15142),
		.dout(new_net_15143)
	);

	bfr new_net_15144_bfr_after (
		.din(new_net_15143),
		.dout(new_net_15144)
	);

	bfr new_net_15145_bfr_after (
		.din(new_net_15144),
		.dout(new_net_15145)
	);

	bfr new_net_15146_bfr_after (
		.din(new_net_15145),
		.dout(new_net_15146)
	);

	bfr new_net_15147_bfr_after (
		.din(new_net_15146),
		.dout(new_net_15147)
	);

	bfr new_net_15148_bfr_after (
		.din(new_net_15147),
		.dout(new_net_15148)
	);

	bfr new_net_15149_bfr_after (
		.din(new_net_15148),
		.dout(new_net_15149)
	);

	bfr new_net_15150_bfr_after (
		.din(new_net_15149),
		.dout(new_net_15150)
	);

	bfr new_net_15151_bfr_after (
		.din(new_net_15150),
		.dout(new_net_15151)
	);

	bfr new_net_15152_bfr_after (
		.din(new_net_15151),
		.dout(new_net_15152)
	);

	bfr new_net_15153_bfr_after (
		.din(new_net_15152),
		.dout(new_net_15153)
	);

	bfr new_net_15154_bfr_after (
		.din(new_net_15153),
		.dout(new_net_15154)
	);

	bfr new_net_15155_bfr_after (
		.din(new_net_15154),
		.dout(new_net_15155)
	);

	bfr new_net_15156_bfr_after (
		.din(new_net_15155),
		.dout(new_net_15156)
	);

	bfr new_net_15157_bfr_after (
		.din(new_net_15156),
		.dout(new_net_15157)
	);

	bfr new_net_15158_bfr_after (
		.din(new_net_15157),
		.dout(new_net_15158)
	);

	bfr new_net_15159_bfr_after (
		.din(new_net_15158),
		.dout(new_net_15159)
	);

	bfr new_net_15160_bfr_after (
		.din(new_net_15159),
		.dout(new_net_15160)
	);

	bfr new_net_15161_bfr_after (
		.din(new_net_15160),
		.dout(new_net_15161)
	);

	bfr new_net_15162_bfr_after (
		.din(new_net_15161),
		.dout(new_net_15162)
	);

	bfr new_net_15163_bfr_after (
		.din(new_net_15162),
		.dout(new_net_15163)
	);

	bfr new_net_15164_bfr_after (
		.din(new_net_15163),
		.dout(new_net_15164)
	);

	bfr new_net_15165_bfr_after (
		.din(new_net_15164),
		.dout(new_net_15165)
	);

	bfr new_net_15166_bfr_after (
		.din(new_net_15165),
		.dout(new_net_15166)
	);

	bfr new_net_15167_bfr_after (
		.din(new_net_15166),
		.dout(new_net_15167)
	);

	bfr new_net_15168_bfr_after (
		.din(new_net_15167),
		.dout(new_net_15168)
	);

	bfr new_net_15169_bfr_after (
		.din(new_net_15168),
		.dout(new_net_15169)
	);

	bfr new_net_15170_bfr_after (
		.din(new_net_15169),
		.dout(new_net_15170)
	);

	bfr new_net_15171_bfr_after (
		.din(new_net_15170),
		.dout(new_net_15171)
	);

	bfr new_net_15172_bfr_after (
		.din(new_net_15171),
		.dout(new_net_15172)
	);

	bfr new_net_15173_bfr_after (
		.din(new_net_15172),
		.dout(new_net_15173)
	);

	bfr new_net_15174_bfr_after (
		.din(new_net_15173),
		.dout(new_net_15174)
	);

	bfr new_net_15175_bfr_after (
		.din(new_net_15174),
		.dout(new_net_15175)
	);

	bfr new_net_15176_bfr_after (
		.din(new_net_15175),
		.dout(new_net_15176)
	);

	bfr new_net_15177_bfr_after (
		.din(new_net_15176),
		.dout(new_net_15177)
	);

	bfr new_net_15178_bfr_after (
		.din(new_net_15177),
		.dout(new_net_15178)
	);

	bfr new_net_15179_bfr_after (
		.din(new_net_15178),
		.dout(new_net_15179)
	);

	bfr new_net_15180_bfr_after (
		.din(new_net_15179),
		.dout(new_net_15180)
	);

	bfr new_net_15181_bfr_after (
		.din(new_net_15180),
		.dout(new_net_15181)
	);

	bfr new_net_15182_bfr_after (
		.din(new_net_15181),
		.dout(new_net_15182)
	);

	bfr new_net_15183_bfr_after (
		.din(new_net_15182),
		.dout(new_net_15183)
	);

	bfr new_net_15184_bfr_after (
		.din(new_net_15183),
		.dout(new_net_15184)
	);

	bfr new_net_15185_bfr_after (
		.din(new_net_15184),
		.dout(new_net_15185)
	);

	bfr new_net_15186_bfr_after (
		.din(new_net_15185),
		.dout(new_net_15186)
	);

	bfr new_net_15187_bfr_after (
		.din(new_net_15186),
		.dout(new_net_15187)
	);

	bfr new_net_15188_bfr_after (
		.din(new_net_15187),
		.dout(new_net_15188)
	);

	bfr new_net_15189_bfr_after (
		.din(new_net_15188),
		.dout(new_net_15189)
	);

	bfr new_net_15190_bfr_after (
		.din(new_net_15189),
		.dout(new_net_15190)
	);

	bfr new_net_15191_bfr_after (
		.din(new_net_15190),
		.dout(new_net_15191)
	);

	bfr new_net_15192_bfr_after (
		.din(new_net_15191),
		.dout(new_net_15192)
	);

	bfr new_net_15193_bfr_after (
		.din(new_net_15192),
		.dout(new_net_15193)
	);

	bfr new_net_15194_bfr_after (
		.din(new_net_15193),
		.dout(new_net_15194)
	);

	bfr new_net_15195_bfr_after (
		.din(new_net_15194),
		.dout(new_net_15195)
	);

	bfr new_net_15196_bfr_after (
		.din(new_net_15195),
		.dout(new_net_15196)
	);

	bfr new_net_15197_bfr_after (
		.din(new_net_15196),
		.dout(new_net_15197)
	);

	bfr new_net_15198_bfr_after (
		.din(new_net_15197),
		.dout(new_net_15198)
	);

	spl2 _0773__v_fanout (
		.a(new_net_15198),
		.b(new_net_1330),
		.c(new_net_1331)
	);

	bfr new_net_15199_bfr_after (
		.din(_1459_),
		.dout(new_net_15199)
	);

	bfr new_net_15200_bfr_after (
		.din(new_net_15199),
		.dout(new_net_15200)
	);

	bfr new_net_15201_bfr_after (
		.din(new_net_15200),
		.dout(new_net_15201)
	);

	bfr new_net_15202_bfr_after (
		.din(new_net_15201),
		.dout(new_net_15202)
	);

	bfr new_net_15203_bfr_after (
		.din(new_net_15202),
		.dout(new_net_15203)
	);

	bfr new_net_15204_bfr_after (
		.din(new_net_15203),
		.dout(new_net_15204)
	);

	bfr new_net_15205_bfr_after (
		.din(new_net_15204),
		.dout(new_net_15205)
	);

	bfr new_net_15206_bfr_after (
		.din(new_net_15205),
		.dout(new_net_15206)
	);

	bfr new_net_15207_bfr_after (
		.din(new_net_15206),
		.dout(new_net_15207)
	);

	bfr new_net_15208_bfr_after (
		.din(new_net_15207),
		.dout(new_net_15208)
	);

	bfr new_net_15209_bfr_after (
		.din(new_net_15208),
		.dout(new_net_15209)
	);

	bfr new_net_15210_bfr_after (
		.din(new_net_15209),
		.dout(new_net_15210)
	);

	bfr new_net_15211_bfr_after (
		.din(new_net_15210),
		.dout(new_net_15211)
	);

	bfr new_net_15212_bfr_after (
		.din(new_net_15211),
		.dout(new_net_15212)
	);

	bfr new_net_15213_bfr_after (
		.din(new_net_15212),
		.dout(new_net_15213)
	);

	bfr new_net_15214_bfr_after (
		.din(new_net_15213),
		.dout(new_net_15214)
	);

	bfr new_net_15215_bfr_after (
		.din(new_net_15214),
		.dout(new_net_15215)
	);

	bfr new_net_15216_bfr_after (
		.din(new_net_15215),
		.dout(new_net_15216)
	);

	bfr new_net_15217_bfr_after (
		.din(new_net_15216),
		.dout(new_net_15217)
	);

	bfr new_net_15218_bfr_after (
		.din(new_net_15217),
		.dout(new_net_15218)
	);

	bfr new_net_15219_bfr_after (
		.din(new_net_15218),
		.dout(new_net_15219)
	);

	bfr new_net_15220_bfr_after (
		.din(new_net_15219),
		.dout(new_net_15220)
	);

	bfr new_net_15221_bfr_after (
		.din(new_net_15220),
		.dout(new_net_15221)
	);

	bfr new_net_15222_bfr_after (
		.din(new_net_15221),
		.dout(new_net_15222)
	);

	bfr new_net_15223_bfr_after (
		.din(new_net_15222),
		.dout(new_net_15223)
	);

	bfr new_net_15224_bfr_after (
		.din(new_net_15223),
		.dout(new_net_15224)
	);

	bfr new_net_15225_bfr_after (
		.din(new_net_15224),
		.dout(new_net_15225)
	);

	bfr new_net_15226_bfr_after (
		.din(new_net_15225),
		.dout(new_net_15226)
	);

	bfr new_net_15227_bfr_after (
		.din(new_net_15226),
		.dout(new_net_15227)
	);

	bfr new_net_15228_bfr_after (
		.din(new_net_15227),
		.dout(new_net_15228)
	);

	bfr new_net_15229_bfr_after (
		.din(new_net_15228),
		.dout(new_net_15229)
	);

	bfr new_net_15230_bfr_after (
		.din(new_net_15229),
		.dout(new_net_15230)
	);

	bfr new_net_15231_bfr_after (
		.din(new_net_15230),
		.dout(new_net_15231)
	);

	bfr new_net_15232_bfr_after (
		.din(new_net_15231),
		.dout(new_net_15232)
	);

	bfr new_net_15233_bfr_after (
		.din(new_net_15232),
		.dout(new_net_15233)
	);

	bfr new_net_15234_bfr_after (
		.din(new_net_15233),
		.dout(new_net_15234)
	);

	bfr new_net_15235_bfr_after (
		.din(new_net_15234),
		.dout(new_net_15235)
	);

	bfr new_net_15236_bfr_after (
		.din(new_net_15235),
		.dout(new_net_15236)
	);

	bfr new_net_15237_bfr_after (
		.din(new_net_15236),
		.dout(new_net_15237)
	);

	bfr new_net_15238_bfr_after (
		.din(new_net_15237),
		.dout(new_net_15238)
	);

	bfr new_net_15239_bfr_after (
		.din(new_net_15238),
		.dout(new_net_15239)
	);

	bfr new_net_15240_bfr_after (
		.din(new_net_15239),
		.dout(new_net_15240)
	);

	bfr new_net_15241_bfr_after (
		.din(new_net_15240),
		.dout(new_net_15241)
	);

	bfr new_net_15242_bfr_after (
		.din(new_net_15241),
		.dout(new_net_15242)
	);

	bfr new_net_15243_bfr_after (
		.din(new_net_15242),
		.dout(new_net_15243)
	);

	bfr new_net_15244_bfr_after (
		.din(new_net_15243),
		.dout(new_net_15244)
	);

	bfr new_net_15245_bfr_after (
		.din(new_net_15244),
		.dout(new_net_15245)
	);

	bfr new_net_15246_bfr_after (
		.din(new_net_15245),
		.dout(new_net_15246)
	);

	bfr new_net_15247_bfr_after (
		.din(new_net_15246),
		.dout(new_net_15247)
	);

	bfr new_net_15248_bfr_after (
		.din(new_net_15247),
		.dout(new_net_15248)
	);

	bfr new_net_15249_bfr_after (
		.din(new_net_15248),
		.dout(new_net_15249)
	);

	bfr new_net_15250_bfr_after (
		.din(new_net_15249),
		.dout(new_net_15250)
	);

	bfr new_net_15251_bfr_after (
		.din(new_net_15250),
		.dout(new_net_15251)
	);

	bfr new_net_15252_bfr_after (
		.din(new_net_15251),
		.dout(new_net_15252)
	);

	bfr new_net_15253_bfr_after (
		.din(new_net_15252),
		.dout(new_net_15253)
	);

	bfr new_net_15254_bfr_after (
		.din(new_net_15253),
		.dout(new_net_15254)
	);

	bfr new_net_15255_bfr_after (
		.din(new_net_15254),
		.dout(new_net_15255)
	);

	bfr new_net_15256_bfr_after (
		.din(new_net_15255),
		.dout(new_net_15256)
	);

	bfr new_net_15257_bfr_after (
		.din(new_net_15256),
		.dout(new_net_15257)
	);

	bfr new_net_15258_bfr_after (
		.din(new_net_15257),
		.dout(new_net_15258)
	);

	bfr new_net_15259_bfr_after (
		.din(new_net_15258),
		.dout(new_net_15259)
	);

	bfr new_net_15260_bfr_after (
		.din(new_net_15259),
		.dout(new_net_15260)
	);

	bfr new_net_15261_bfr_after (
		.din(new_net_15260),
		.dout(new_net_15261)
	);

	bfr new_net_15262_bfr_after (
		.din(new_net_15261),
		.dout(new_net_15262)
	);

	bfr new_net_15263_bfr_after (
		.din(new_net_15262),
		.dout(new_net_15263)
	);

	bfr new_net_15264_bfr_after (
		.din(new_net_15263),
		.dout(new_net_15264)
	);

	bfr new_net_15265_bfr_after (
		.din(new_net_15264),
		.dout(new_net_15265)
	);

	bfr new_net_15266_bfr_after (
		.din(new_net_15265),
		.dout(new_net_15266)
	);

	bfr new_net_15267_bfr_after (
		.din(new_net_15266),
		.dout(new_net_15267)
	);

	bfr new_net_15268_bfr_after (
		.din(new_net_15267),
		.dout(new_net_15268)
	);

	bfr new_net_15269_bfr_after (
		.din(new_net_15268),
		.dout(new_net_15269)
	);

	bfr new_net_15270_bfr_after (
		.din(new_net_15269),
		.dout(new_net_15270)
	);

	spl2 _1459__v_fanout (
		.a(new_net_15270),
		.b(new_net_2795),
		.c(new_net_2796)
	);

	bfr new_net_15271_bfr_after (
		.din(_0529_),
		.dout(new_net_15271)
	);

	bfr new_net_15272_bfr_after (
		.din(new_net_15271),
		.dout(new_net_15272)
	);

	bfr new_net_15273_bfr_after (
		.din(new_net_15272),
		.dout(new_net_15273)
	);

	bfr new_net_15274_bfr_after (
		.din(new_net_15273),
		.dout(new_net_15274)
	);

	bfr new_net_15275_bfr_after (
		.din(new_net_15274),
		.dout(new_net_15275)
	);

	bfr new_net_15276_bfr_after (
		.din(new_net_15275),
		.dout(new_net_15276)
	);

	bfr new_net_15277_bfr_after (
		.din(new_net_15276),
		.dout(new_net_15277)
	);

	bfr new_net_15278_bfr_after (
		.din(new_net_15277),
		.dout(new_net_15278)
	);

	bfr new_net_15279_bfr_after (
		.din(new_net_15278),
		.dout(new_net_15279)
	);

	bfr new_net_15280_bfr_after (
		.din(new_net_15279),
		.dout(new_net_15280)
	);

	bfr new_net_15281_bfr_after (
		.din(new_net_15280),
		.dout(new_net_15281)
	);

	bfr new_net_15282_bfr_after (
		.din(new_net_15281),
		.dout(new_net_15282)
	);

	bfr new_net_15283_bfr_after (
		.din(new_net_15282),
		.dout(new_net_15283)
	);

	bfr new_net_15284_bfr_after (
		.din(new_net_15283),
		.dout(new_net_15284)
	);

	bfr new_net_15285_bfr_after (
		.din(new_net_15284),
		.dout(new_net_15285)
	);

	bfr new_net_15286_bfr_after (
		.din(new_net_15285),
		.dout(new_net_15286)
	);

	bfr new_net_15287_bfr_after (
		.din(new_net_15286),
		.dout(new_net_15287)
	);

	bfr new_net_15288_bfr_after (
		.din(new_net_15287),
		.dout(new_net_15288)
	);

	bfr new_net_15289_bfr_after (
		.din(new_net_15288),
		.dout(new_net_15289)
	);

	bfr new_net_15290_bfr_after (
		.din(new_net_15289),
		.dout(new_net_15290)
	);

	bfr new_net_15291_bfr_after (
		.din(new_net_15290),
		.dout(new_net_15291)
	);

	bfr new_net_15292_bfr_after (
		.din(new_net_15291),
		.dout(new_net_15292)
	);

	bfr new_net_15293_bfr_after (
		.din(new_net_15292),
		.dout(new_net_15293)
	);

	bfr new_net_15294_bfr_after (
		.din(new_net_15293),
		.dout(new_net_15294)
	);

	bfr new_net_15295_bfr_after (
		.din(new_net_15294),
		.dout(new_net_15295)
	);

	bfr new_net_15296_bfr_after (
		.din(new_net_15295),
		.dout(new_net_15296)
	);

	bfr new_net_15297_bfr_after (
		.din(new_net_15296),
		.dout(new_net_15297)
	);

	bfr new_net_15298_bfr_after (
		.din(new_net_15297),
		.dout(new_net_15298)
	);

	bfr new_net_15299_bfr_after (
		.din(new_net_15298),
		.dout(new_net_15299)
	);

	bfr new_net_15300_bfr_after (
		.din(new_net_15299),
		.dout(new_net_15300)
	);

	bfr new_net_15301_bfr_after (
		.din(new_net_15300),
		.dout(new_net_15301)
	);

	bfr new_net_15302_bfr_after (
		.din(new_net_15301),
		.dout(new_net_15302)
	);

	bfr new_net_15303_bfr_after (
		.din(new_net_15302),
		.dout(new_net_15303)
	);

	bfr new_net_15304_bfr_after (
		.din(new_net_15303),
		.dout(new_net_15304)
	);

	bfr new_net_15305_bfr_after (
		.din(new_net_15304),
		.dout(new_net_15305)
	);

	bfr new_net_15306_bfr_after (
		.din(new_net_15305),
		.dout(new_net_15306)
	);

	bfr new_net_15307_bfr_after (
		.din(new_net_15306),
		.dout(new_net_15307)
	);

	bfr new_net_15308_bfr_after (
		.din(new_net_15307),
		.dout(new_net_15308)
	);

	bfr new_net_15309_bfr_after (
		.din(new_net_15308),
		.dout(new_net_15309)
	);

	bfr new_net_15310_bfr_after (
		.din(new_net_15309),
		.dout(new_net_15310)
	);

	bfr new_net_15311_bfr_after (
		.din(new_net_15310),
		.dout(new_net_15311)
	);

	bfr new_net_15312_bfr_after (
		.din(new_net_15311),
		.dout(new_net_15312)
	);

	bfr new_net_15313_bfr_after (
		.din(new_net_15312),
		.dout(new_net_15313)
	);

	bfr new_net_15314_bfr_after (
		.din(new_net_15313),
		.dout(new_net_15314)
	);

	bfr new_net_15315_bfr_after (
		.din(new_net_15314),
		.dout(new_net_15315)
	);

	bfr new_net_15316_bfr_after (
		.din(new_net_15315),
		.dout(new_net_15316)
	);

	bfr new_net_15317_bfr_after (
		.din(new_net_15316),
		.dout(new_net_15317)
	);

	bfr new_net_15318_bfr_after (
		.din(new_net_15317),
		.dout(new_net_15318)
	);

	bfr new_net_15319_bfr_after (
		.din(new_net_15318),
		.dout(new_net_15319)
	);

	bfr new_net_15320_bfr_after (
		.din(new_net_15319),
		.dout(new_net_15320)
	);

	bfr new_net_15321_bfr_after (
		.din(new_net_15320),
		.dout(new_net_15321)
	);

	bfr new_net_15322_bfr_after (
		.din(new_net_15321),
		.dout(new_net_15322)
	);

	bfr new_net_15323_bfr_after (
		.din(new_net_15322),
		.dout(new_net_15323)
	);

	bfr new_net_15324_bfr_after (
		.din(new_net_15323),
		.dout(new_net_15324)
	);

	bfr new_net_15325_bfr_after (
		.din(new_net_15324),
		.dout(new_net_15325)
	);

	bfr new_net_15326_bfr_after (
		.din(new_net_15325),
		.dout(new_net_15326)
	);

	bfr new_net_15327_bfr_after (
		.din(new_net_15326),
		.dout(new_net_15327)
	);

	bfr new_net_15328_bfr_after (
		.din(new_net_15327),
		.dout(new_net_15328)
	);

	bfr new_net_15329_bfr_after (
		.din(new_net_15328),
		.dout(new_net_15329)
	);

	bfr new_net_15330_bfr_after (
		.din(new_net_15329),
		.dout(new_net_15330)
	);

	bfr new_net_15331_bfr_after (
		.din(new_net_15330),
		.dout(new_net_15331)
	);

	bfr new_net_15332_bfr_after (
		.din(new_net_15331),
		.dout(new_net_15332)
	);

	bfr new_net_15333_bfr_after (
		.din(new_net_15332),
		.dout(new_net_15333)
	);

	bfr new_net_15334_bfr_after (
		.din(new_net_15333),
		.dout(new_net_15334)
	);

	bfr new_net_15335_bfr_after (
		.din(new_net_15334),
		.dout(new_net_15335)
	);

	bfr new_net_15336_bfr_after (
		.din(new_net_15335),
		.dout(new_net_15336)
	);

	bfr new_net_15337_bfr_after (
		.din(new_net_15336),
		.dout(new_net_15337)
	);

	bfr new_net_15338_bfr_after (
		.din(new_net_15337),
		.dout(new_net_15338)
	);

	bfr new_net_15339_bfr_after (
		.din(new_net_15338),
		.dout(new_net_15339)
	);

	bfr new_net_15340_bfr_after (
		.din(new_net_15339),
		.dout(new_net_15340)
	);

	bfr new_net_15341_bfr_after (
		.din(new_net_15340),
		.dout(new_net_15341)
	);

	bfr new_net_15342_bfr_after (
		.din(new_net_15341),
		.dout(new_net_15342)
	);

	bfr new_net_15343_bfr_after (
		.din(new_net_15342),
		.dout(new_net_15343)
	);

	bfr new_net_15344_bfr_after (
		.din(new_net_15343),
		.dout(new_net_15344)
	);

	bfr new_net_15345_bfr_after (
		.din(new_net_15344),
		.dout(new_net_15345)
	);

	bfr new_net_15346_bfr_after (
		.din(new_net_15345),
		.dout(new_net_15346)
	);

	bfr new_net_15347_bfr_after (
		.din(new_net_15346),
		.dout(new_net_15347)
	);

	bfr new_net_15348_bfr_after (
		.din(new_net_15347),
		.dout(new_net_15348)
	);

	bfr new_net_15349_bfr_after (
		.din(new_net_15348),
		.dout(new_net_15349)
	);

	bfr new_net_15350_bfr_after (
		.din(new_net_15349),
		.dout(new_net_15350)
	);

	bfr new_net_15351_bfr_after (
		.din(new_net_15350),
		.dout(new_net_15351)
	);

	bfr new_net_15352_bfr_after (
		.din(new_net_15351),
		.dout(new_net_15352)
	);

	bfr new_net_15353_bfr_after (
		.din(new_net_15352),
		.dout(new_net_15353)
	);

	bfr new_net_15354_bfr_after (
		.din(new_net_15353),
		.dout(new_net_15354)
	);

	bfr new_net_15355_bfr_after (
		.din(new_net_15354),
		.dout(new_net_15355)
	);

	bfr new_net_15356_bfr_after (
		.din(new_net_15355),
		.dout(new_net_15356)
	);

	bfr new_net_15357_bfr_after (
		.din(new_net_15356),
		.dout(new_net_15357)
	);

	bfr new_net_15358_bfr_after (
		.din(new_net_15357),
		.dout(new_net_15358)
	);

	bfr new_net_15359_bfr_after (
		.din(new_net_15358),
		.dout(new_net_15359)
	);

	bfr new_net_15360_bfr_after (
		.din(new_net_15359),
		.dout(new_net_15360)
	);

	bfr new_net_15361_bfr_after (
		.din(new_net_15360),
		.dout(new_net_15361)
	);

	bfr new_net_15362_bfr_after (
		.din(new_net_15361),
		.dout(new_net_15362)
	);

	bfr new_net_15363_bfr_after (
		.din(new_net_15362),
		.dout(new_net_15363)
	);

	bfr new_net_15364_bfr_after (
		.din(new_net_15363),
		.dout(new_net_15364)
	);

	bfr new_net_15365_bfr_after (
		.din(new_net_15364),
		.dout(new_net_15365)
	);

	bfr new_net_15366_bfr_after (
		.din(new_net_15365),
		.dout(new_net_15366)
	);

	bfr new_net_15367_bfr_after (
		.din(new_net_15366),
		.dout(new_net_15367)
	);

	bfr new_net_15368_bfr_after (
		.din(new_net_15367),
		.dout(new_net_15368)
	);

	bfr new_net_15369_bfr_after (
		.din(new_net_15368),
		.dout(new_net_15369)
	);

	bfr new_net_15370_bfr_after (
		.din(new_net_15369),
		.dout(new_net_15370)
	);

	bfr new_net_15371_bfr_after (
		.din(new_net_15370),
		.dout(new_net_15371)
	);

	bfr new_net_15372_bfr_after (
		.din(new_net_15371),
		.dout(new_net_15372)
	);

	bfr new_net_15373_bfr_after (
		.din(new_net_15372),
		.dout(new_net_15373)
	);

	bfr new_net_15374_bfr_after (
		.din(new_net_15373),
		.dout(new_net_15374)
	);

	bfr new_net_15375_bfr_after (
		.din(new_net_15374),
		.dout(new_net_15375)
	);

	bfr new_net_15376_bfr_after (
		.din(new_net_15375),
		.dout(new_net_15376)
	);

	bfr new_net_15377_bfr_after (
		.din(new_net_15376),
		.dout(new_net_15377)
	);

	bfr new_net_15378_bfr_after (
		.din(new_net_15377),
		.dout(new_net_15378)
	);

	bfr new_net_15379_bfr_after (
		.din(new_net_15378),
		.dout(new_net_15379)
	);

	bfr new_net_15380_bfr_after (
		.din(new_net_15379),
		.dout(new_net_15380)
	);

	bfr new_net_15381_bfr_after (
		.din(new_net_15380),
		.dout(new_net_15381)
	);

	bfr new_net_15382_bfr_after (
		.din(new_net_15381),
		.dout(new_net_15382)
	);

	spl2 _0529__v_fanout (
		.a(new_net_15382),
		.b(new_net_1980),
		.c(new_net_1981)
	);

	bfr new_net_15383_bfr_after (
		.din(_1017_),
		.dout(new_net_15383)
	);

	bfr new_net_15384_bfr_after (
		.din(new_net_15383),
		.dout(new_net_15384)
	);

	bfr new_net_15385_bfr_after (
		.din(new_net_15384),
		.dout(new_net_15385)
	);

	bfr new_net_15386_bfr_after (
		.din(new_net_15385),
		.dout(new_net_15386)
	);

	bfr new_net_15387_bfr_after (
		.din(new_net_15386),
		.dout(new_net_15387)
	);

	bfr new_net_15388_bfr_after (
		.din(new_net_15387),
		.dout(new_net_15388)
	);

	bfr new_net_15389_bfr_after (
		.din(new_net_15388),
		.dout(new_net_15389)
	);

	bfr new_net_15390_bfr_after (
		.din(new_net_15389),
		.dout(new_net_15390)
	);

	bfr new_net_15391_bfr_after (
		.din(new_net_15390),
		.dout(new_net_15391)
	);

	bfr new_net_15392_bfr_after (
		.din(new_net_15391),
		.dout(new_net_15392)
	);

	bfr new_net_15393_bfr_after (
		.din(new_net_15392),
		.dout(new_net_15393)
	);

	bfr new_net_15394_bfr_after (
		.din(new_net_15393),
		.dout(new_net_15394)
	);

	bfr new_net_15395_bfr_after (
		.din(new_net_15394),
		.dout(new_net_15395)
	);

	bfr new_net_15396_bfr_after (
		.din(new_net_15395),
		.dout(new_net_15396)
	);

	bfr new_net_15397_bfr_after (
		.din(new_net_15396),
		.dout(new_net_15397)
	);

	bfr new_net_15398_bfr_after (
		.din(new_net_15397),
		.dout(new_net_15398)
	);

	bfr new_net_15399_bfr_after (
		.din(new_net_15398),
		.dout(new_net_15399)
	);

	bfr new_net_15400_bfr_after (
		.din(new_net_15399),
		.dout(new_net_15400)
	);

	bfr new_net_15401_bfr_after (
		.din(new_net_15400),
		.dout(new_net_15401)
	);

	bfr new_net_15402_bfr_after (
		.din(new_net_15401),
		.dout(new_net_15402)
	);

	bfr new_net_15403_bfr_after (
		.din(new_net_15402),
		.dout(new_net_15403)
	);

	bfr new_net_15404_bfr_after (
		.din(new_net_15403),
		.dout(new_net_15404)
	);

	bfr new_net_15405_bfr_after (
		.din(new_net_15404),
		.dout(new_net_15405)
	);

	bfr new_net_15406_bfr_after (
		.din(new_net_15405),
		.dout(new_net_15406)
	);

	bfr new_net_15407_bfr_after (
		.din(new_net_15406),
		.dout(new_net_15407)
	);

	bfr new_net_15408_bfr_after (
		.din(new_net_15407),
		.dout(new_net_15408)
	);

	bfr new_net_15409_bfr_after (
		.din(new_net_15408),
		.dout(new_net_15409)
	);

	bfr new_net_15410_bfr_after (
		.din(new_net_15409),
		.dout(new_net_15410)
	);

	bfr new_net_15411_bfr_after (
		.din(new_net_15410),
		.dout(new_net_15411)
	);

	bfr new_net_15412_bfr_after (
		.din(new_net_15411),
		.dout(new_net_15412)
	);

	bfr new_net_15413_bfr_after (
		.din(new_net_15412),
		.dout(new_net_15413)
	);

	bfr new_net_15414_bfr_after (
		.din(new_net_15413),
		.dout(new_net_15414)
	);

	bfr new_net_15415_bfr_after (
		.din(new_net_15414),
		.dout(new_net_15415)
	);

	bfr new_net_15416_bfr_after (
		.din(new_net_15415),
		.dout(new_net_15416)
	);

	bfr new_net_15417_bfr_after (
		.din(new_net_15416),
		.dout(new_net_15417)
	);

	bfr new_net_15418_bfr_after (
		.din(new_net_15417),
		.dout(new_net_15418)
	);

	bfr new_net_15419_bfr_after (
		.din(new_net_15418),
		.dout(new_net_15419)
	);

	bfr new_net_15420_bfr_after (
		.din(new_net_15419),
		.dout(new_net_15420)
	);

	bfr new_net_15421_bfr_after (
		.din(new_net_15420),
		.dout(new_net_15421)
	);

	bfr new_net_15422_bfr_after (
		.din(new_net_15421),
		.dout(new_net_15422)
	);

	spl2 _1017__v_fanout (
		.a(new_net_15422),
		.b(new_net_1092),
		.c(new_net_1093)
	);

	bfr new_net_15423_bfr_after (
		.din(_1584_),
		.dout(new_net_15423)
	);

	bfr new_net_15424_bfr_after (
		.din(new_net_15423),
		.dout(new_net_15424)
	);

	bfr new_net_15425_bfr_after (
		.din(new_net_15424),
		.dout(new_net_15425)
	);

	bfr new_net_15426_bfr_after (
		.din(new_net_15425),
		.dout(new_net_15426)
	);

	bfr new_net_15427_bfr_after (
		.din(new_net_15426),
		.dout(new_net_15427)
	);

	bfr new_net_15428_bfr_after (
		.din(new_net_15427),
		.dout(new_net_15428)
	);

	bfr new_net_15429_bfr_after (
		.din(new_net_15428),
		.dout(new_net_15429)
	);

	bfr new_net_15430_bfr_after (
		.din(new_net_15429),
		.dout(new_net_15430)
	);

	bfr new_net_15431_bfr_after (
		.din(new_net_15430),
		.dout(new_net_15431)
	);

	bfr new_net_15432_bfr_after (
		.din(new_net_15431),
		.dout(new_net_15432)
	);

	bfr new_net_15433_bfr_after (
		.din(new_net_15432),
		.dout(new_net_15433)
	);

	bfr new_net_15434_bfr_after (
		.din(new_net_15433),
		.dout(new_net_15434)
	);

	bfr new_net_15435_bfr_after (
		.din(new_net_15434),
		.dout(new_net_15435)
	);

	bfr new_net_15436_bfr_after (
		.din(new_net_15435),
		.dout(new_net_15436)
	);

	bfr new_net_15437_bfr_after (
		.din(new_net_15436),
		.dout(new_net_15437)
	);

	bfr new_net_15438_bfr_after (
		.din(new_net_15437),
		.dout(new_net_15438)
	);

	spl2 _1584__v_fanout (
		.a(new_net_15438),
		.b(new_net_671),
		.c(new_net_672)
	);

	bfr new_net_15439_bfr_after (
		.din(_0432_),
		.dout(new_net_15439)
	);

	bfr new_net_15440_bfr_after (
		.din(new_net_15439),
		.dout(new_net_15440)
	);

	bfr new_net_15441_bfr_after (
		.din(new_net_15440),
		.dout(new_net_15441)
	);

	bfr new_net_15442_bfr_after (
		.din(new_net_15441),
		.dout(new_net_15442)
	);

	bfr new_net_15443_bfr_after (
		.din(new_net_15442),
		.dout(new_net_15443)
	);

	bfr new_net_15444_bfr_after (
		.din(new_net_15443),
		.dout(new_net_15444)
	);

	bfr new_net_15445_bfr_after (
		.din(new_net_15444),
		.dout(new_net_15445)
	);

	bfr new_net_15446_bfr_after (
		.din(new_net_15445),
		.dout(new_net_15446)
	);

	bfr new_net_15447_bfr_after (
		.din(new_net_15446),
		.dout(new_net_15447)
	);

	bfr new_net_15448_bfr_after (
		.din(new_net_15447),
		.dout(new_net_15448)
	);

	bfr new_net_15449_bfr_after (
		.din(new_net_15448),
		.dout(new_net_15449)
	);

	bfr new_net_15450_bfr_after (
		.din(new_net_15449),
		.dout(new_net_15450)
	);

	bfr new_net_15451_bfr_after (
		.din(new_net_15450),
		.dout(new_net_15451)
	);

	bfr new_net_15452_bfr_after (
		.din(new_net_15451),
		.dout(new_net_15452)
	);

	bfr new_net_15453_bfr_after (
		.din(new_net_15452),
		.dout(new_net_15453)
	);

	bfr new_net_15454_bfr_after (
		.din(new_net_15453),
		.dout(new_net_15454)
	);

	bfr new_net_15455_bfr_after (
		.din(new_net_15454),
		.dout(new_net_15455)
	);

	bfr new_net_15456_bfr_after (
		.din(new_net_15455),
		.dout(new_net_15456)
	);

	bfr new_net_15457_bfr_after (
		.din(new_net_15456),
		.dout(new_net_15457)
	);

	bfr new_net_15458_bfr_after (
		.din(new_net_15457),
		.dout(new_net_15458)
	);

	bfr new_net_15459_bfr_after (
		.din(new_net_15458),
		.dout(new_net_15459)
	);

	bfr new_net_15460_bfr_after (
		.din(new_net_15459),
		.dout(new_net_15460)
	);

	bfr new_net_15461_bfr_after (
		.din(new_net_15460),
		.dout(new_net_15461)
	);

	bfr new_net_15462_bfr_after (
		.din(new_net_15461),
		.dout(new_net_15462)
	);

	bfr new_net_15463_bfr_after (
		.din(new_net_15462),
		.dout(new_net_15463)
	);

	bfr new_net_15464_bfr_after (
		.din(new_net_15463),
		.dout(new_net_15464)
	);

	bfr new_net_15465_bfr_after (
		.din(new_net_15464),
		.dout(new_net_15465)
	);

	bfr new_net_15466_bfr_after (
		.din(new_net_15465),
		.dout(new_net_15466)
	);

	bfr new_net_15467_bfr_after (
		.din(new_net_15466),
		.dout(new_net_15467)
	);

	bfr new_net_15468_bfr_after (
		.din(new_net_15467),
		.dout(new_net_15468)
	);

	bfr new_net_15469_bfr_after (
		.din(new_net_15468),
		.dout(new_net_15469)
	);

	bfr new_net_15470_bfr_after (
		.din(new_net_15469),
		.dout(new_net_15470)
	);

	bfr new_net_15471_bfr_after (
		.din(new_net_15470),
		.dout(new_net_15471)
	);

	bfr new_net_15472_bfr_after (
		.din(new_net_15471),
		.dout(new_net_15472)
	);

	bfr new_net_15473_bfr_after (
		.din(new_net_15472),
		.dout(new_net_15473)
	);

	bfr new_net_15474_bfr_after (
		.din(new_net_15473),
		.dout(new_net_15474)
	);

	bfr new_net_15475_bfr_after (
		.din(new_net_15474),
		.dout(new_net_15475)
	);

	bfr new_net_15476_bfr_after (
		.din(new_net_15475),
		.dout(new_net_15476)
	);

	bfr new_net_15477_bfr_after (
		.din(new_net_15476),
		.dout(new_net_15477)
	);

	bfr new_net_15478_bfr_after (
		.din(new_net_15477),
		.dout(new_net_15478)
	);

	bfr new_net_15479_bfr_after (
		.din(new_net_15478),
		.dout(new_net_15479)
	);

	bfr new_net_15480_bfr_after (
		.din(new_net_15479),
		.dout(new_net_15480)
	);

	bfr new_net_15481_bfr_after (
		.din(new_net_15480),
		.dout(new_net_15481)
	);

	bfr new_net_15482_bfr_after (
		.din(new_net_15481),
		.dout(new_net_15482)
	);

	bfr new_net_15483_bfr_after (
		.din(new_net_15482),
		.dout(new_net_15483)
	);

	bfr new_net_15484_bfr_after (
		.din(new_net_15483),
		.dout(new_net_15484)
	);

	bfr new_net_15485_bfr_after (
		.din(new_net_15484),
		.dout(new_net_15485)
	);

	bfr new_net_15486_bfr_after (
		.din(new_net_15485),
		.dout(new_net_15486)
	);

	bfr new_net_15487_bfr_after (
		.din(new_net_15486),
		.dout(new_net_15487)
	);

	bfr new_net_15488_bfr_after (
		.din(new_net_15487),
		.dout(new_net_15488)
	);

	bfr new_net_15489_bfr_after (
		.din(new_net_15488),
		.dout(new_net_15489)
	);

	bfr new_net_15490_bfr_after (
		.din(new_net_15489),
		.dout(new_net_15490)
	);

	bfr new_net_15491_bfr_after (
		.din(new_net_15490),
		.dout(new_net_15491)
	);

	bfr new_net_15492_bfr_after (
		.din(new_net_15491),
		.dout(new_net_15492)
	);

	bfr new_net_15493_bfr_after (
		.din(new_net_15492),
		.dout(new_net_15493)
	);

	bfr new_net_15494_bfr_after (
		.din(new_net_15493),
		.dout(new_net_15494)
	);

	bfr new_net_15495_bfr_after (
		.din(new_net_15494),
		.dout(new_net_15495)
	);

	bfr new_net_15496_bfr_after (
		.din(new_net_15495),
		.dout(new_net_15496)
	);

	bfr new_net_15497_bfr_after (
		.din(new_net_15496),
		.dout(new_net_15497)
	);

	bfr new_net_15498_bfr_after (
		.din(new_net_15497),
		.dout(new_net_15498)
	);

	bfr new_net_15499_bfr_after (
		.din(new_net_15498),
		.dout(new_net_15499)
	);

	bfr new_net_15500_bfr_after (
		.din(new_net_15499),
		.dout(new_net_15500)
	);

	bfr new_net_15501_bfr_after (
		.din(new_net_15500),
		.dout(new_net_15501)
	);

	bfr new_net_15502_bfr_after (
		.din(new_net_15501),
		.dout(new_net_15502)
	);

	bfr new_net_15503_bfr_after (
		.din(new_net_15502),
		.dout(new_net_15503)
	);

	bfr new_net_15504_bfr_after (
		.din(new_net_15503),
		.dout(new_net_15504)
	);

	bfr new_net_15505_bfr_after (
		.din(new_net_15504),
		.dout(new_net_15505)
	);

	bfr new_net_15506_bfr_after (
		.din(new_net_15505),
		.dout(new_net_15506)
	);

	bfr new_net_15507_bfr_after (
		.din(new_net_15506),
		.dout(new_net_15507)
	);

	bfr new_net_15508_bfr_after (
		.din(new_net_15507),
		.dout(new_net_15508)
	);

	bfr new_net_15509_bfr_after (
		.din(new_net_15508),
		.dout(new_net_15509)
	);

	bfr new_net_15510_bfr_after (
		.din(new_net_15509),
		.dout(new_net_15510)
	);

	bfr new_net_15511_bfr_after (
		.din(new_net_15510),
		.dout(new_net_15511)
	);

	bfr new_net_15512_bfr_after (
		.din(new_net_15511),
		.dout(new_net_15512)
	);

	bfr new_net_15513_bfr_after (
		.din(new_net_15512),
		.dout(new_net_15513)
	);

	bfr new_net_15514_bfr_after (
		.din(new_net_15513),
		.dout(new_net_15514)
	);

	bfr new_net_15515_bfr_after (
		.din(new_net_15514),
		.dout(new_net_15515)
	);

	bfr new_net_15516_bfr_after (
		.din(new_net_15515),
		.dout(new_net_15516)
	);

	bfr new_net_15517_bfr_after (
		.din(new_net_15516),
		.dout(new_net_15517)
	);

	bfr new_net_15518_bfr_after (
		.din(new_net_15517),
		.dout(new_net_15518)
	);

	bfr new_net_15519_bfr_after (
		.din(new_net_15518),
		.dout(new_net_15519)
	);

	bfr new_net_15520_bfr_after (
		.din(new_net_15519),
		.dout(new_net_15520)
	);

	bfr new_net_15521_bfr_after (
		.din(new_net_15520),
		.dout(new_net_15521)
	);

	bfr new_net_15522_bfr_after (
		.din(new_net_15521),
		.dout(new_net_15522)
	);

	bfr new_net_15523_bfr_after (
		.din(new_net_15522),
		.dout(new_net_15523)
	);

	bfr new_net_15524_bfr_after (
		.din(new_net_15523),
		.dout(new_net_15524)
	);

	bfr new_net_15525_bfr_after (
		.din(new_net_15524),
		.dout(new_net_15525)
	);

	bfr new_net_15526_bfr_after (
		.din(new_net_15525),
		.dout(new_net_15526)
	);

	bfr new_net_15527_bfr_after (
		.din(new_net_15526),
		.dout(new_net_15527)
	);

	bfr new_net_15528_bfr_after (
		.din(new_net_15527),
		.dout(new_net_15528)
	);

	bfr new_net_15529_bfr_after (
		.din(new_net_15528),
		.dout(new_net_15529)
	);

	bfr new_net_15530_bfr_after (
		.din(new_net_15529),
		.dout(new_net_15530)
	);

	bfr new_net_15531_bfr_after (
		.din(new_net_15530),
		.dout(new_net_15531)
	);

	bfr new_net_15532_bfr_after (
		.din(new_net_15531),
		.dout(new_net_15532)
	);

	bfr new_net_15533_bfr_after (
		.din(new_net_15532),
		.dout(new_net_15533)
	);

	bfr new_net_15534_bfr_after (
		.din(new_net_15533),
		.dout(new_net_15534)
	);

	bfr new_net_15535_bfr_after (
		.din(new_net_15534),
		.dout(new_net_15535)
	);

	bfr new_net_15536_bfr_after (
		.din(new_net_15535),
		.dout(new_net_15536)
	);

	bfr new_net_15537_bfr_after (
		.din(new_net_15536),
		.dout(new_net_15537)
	);

	bfr new_net_15538_bfr_after (
		.din(new_net_15537),
		.dout(new_net_15538)
	);

	bfr new_net_15539_bfr_after (
		.din(new_net_15538),
		.dout(new_net_15539)
	);

	bfr new_net_15540_bfr_after (
		.din(new_net_15539),
		.dout(new_net_15540)
	);

	bfr new_net_15541_bfr_after (
		.din(new_net_15540),
		.dout(new_net_15541)
	);

	bfr new_net_15542_bfr_after (
		.din(new_net_15541),
		.dout(new_net_15542)
	);

	bfr new_net_15543_bfr_after (
		.din(new_net_15542),
		.dout(new_net_15543)
	);

	bfr new_net_15544_bfr_after (
		.din(new_net_15543),
		.dout(new_net_15544)
	);

	bfr new_net_15545_bfr_after (
		.din(new_net_15544),
		.dout(new_net_15545)
	);

	bfr new_net_15546_bfr_after (
		.din(new_net_15545),
		.dout(new_net_15546)
	);

	bfr new_net_15547_bfr_after (
		.din(new_net_15546),
		.dout(new_net_15547)
	);

	bfr new_net_15548_bfr_after (
		.din(new_net_15547),
		.dout(new_net_15548)
	);

	bfr new_net_15549_bfr_after (
		.din(new_net_15548),
		.dout(new_net_15549)
	);

	bfr new_net_15550_bfr_after (
		.din(new_net_15549),
		.dout(new_net_15550)
	);

	spl2 _0432__v_fanout (
		.a(new_net_15550),
		.b(new_net_1778),
		.c(new_net_1779)
	);

	bfr new_net_15551_bfr_after (
		.din(_1284_),
		.dout(new_net_15551)
	);

	bfr new_net_15552_bfr_after (
		.din(new_net_15551),
		.dout(new_net_15552)
	);

	bfr new_net_15553_bfr_after (
		.din(new_net_15552),
		.dout(new_net_15553)
	);

	bfr new_net_15554_bfr_after (
		.din(new_net_15553),
		.dout(new_net_15554)
	);

	bfr new_net_15555_bfr_after (
		.din(new_net_15554),
		.dout(new_net_15555)
	);

	bfr new_net_15556_bfr_after (
		.din(new_net_15555),
		.dout(new_net_15556)
	);

	bfr new_net_15557_bfr_after (
		.din(new_net_15556),
		.dout(new_net_15557)
	);

	bfr new_net_15558_bfr_after (
		.din(new_net_15557),
		.dout(new_net_15558)
	);

	bfr new_net_15559_bfr_after (
		.din(new_net_15558),
		.dout(new_net_15559)
	);

	bfr new_net_15560_bfr_after (
		.din(new_net_15559),
		.dout(new_net_15560)
	);

	bfr new_net_15561_bfr_after (
		.din(new_net_15560),
		.dout(new_net_15561)
	);

	bfr new_net_15562_bfr_after (
		.din(new_net_15561),
		.dout(new_net_15562)
	);

	bfr new_net_15563_bfr_after (
		.din(new_net_15562),
		.dout(new_net_15563)
	);

	bfr new_net_15564_bfr_after (
		.din(new_net_15563),
		.dout(new_net_15564)
	);

	bfr new_net_15565_bfr_after (
		.din(new_net_15564),
		.dout(new_net_15565)
	);

	bfr new_net_15566_bfr_after (
		.din(new_net_15565),
		.dout(new_net_15566)
	);

	bfr new_net_15567_bfr_after (
		.din(new_net_15566),
		.dout(new_net_15567)
	);

	bfr new_net_15568_bfr_after (
		.din(new_net_15567),
		.dout(new_net_15568)
	);

	bfr new_net_15569_bfr_after (
		.din(new_net_15568),
		.dout(new_net_15569)
	);

	bfr new_net_15570_bfr_after (
		.din(new_net_15569),
		.dout(new_net_15570)
	);

	bfr new_net_15571_bfr_after (
		.din(new_net_15570),
		.dout(new_net_15571)
	);

	bfr new_net_15572_bfr_after (
		.din(new_net_15571),
		.dout(new_net_15572)
	);

	bfr new_net_15573_bfr_after (
		.din(new_net_15572),
		.dout(new_net_15573)
	);

	bfr new_net_15574_bfr_after (
		.din(new_net_15573),
		.dout(new_net_15574)
	);

	bfr new_net_15575_bfr_after (
		.din(new_net_15574),
		.dout(new_net_15575)
	);

	bfr new_net_15576_bfr_after (
		.din(new_net_15575),
		.dout(new_net_15576)
	);

	bfr new_net_15577_bfr_after (
		.din(new_net_15576),
		.dout(new_net_15577)
	);

	bfr new_net_15578_bfr_after (
		.din(new_net_15577),
		.dout(new_net_15578)
	);

	bfr new_net_15579_bfr_after (
		.din(new_net_15578),
		.dout(new_net_15579)
	);

	bfr new_net_15580_bfr_after (
		.din(new_net_15579),
		.dout(new_net_15580)
	);

	bfr new_net_15581_bfr_after (
		.din(new_net_15580),
		.dout(new_net_15581)
	);

	bfr new_net_15582_bfr_after (
		.din(new_net_15581),
		.dout(new_net_15582)
	);

	bfr new_net_15583_bfr_after (
		.din(new_net_15582),
		.dout(new_net_15583)
	);

	bfr new_net_15584_bfr_after (
		.din(new_net_15583),
		.dout(new_net_15584)
	);

	bfr new_net_15585_bfr_after (
		.din(new_net_15584),
		.dout(new_net_15585)
	);

	bfr new_net_15586_bfr_after (
		.din(new_net_15585),
		.dout(new_net_15586)
	);

	bfr new_net_15587_bfr_after (
		.din(new_net_15586),
		.dout(new_net_15587)
	);

	bfr new_net_15588_bfr_after (
		.din(new_net_15587),
		.dout(new_net_15588)
	);

	bfr new_net_15589_bfr_after (
		.din(new_net_15588),
		.dout(new_net_15589)
	);

	bfr new_net_15590_bfr_after (
		.din(new_net_15589),
		.dout(new_net_15590)
	);

	bfr new_net_15591_bfr_after (
		.din(new_net_15590),
		.dout(new_net_15591)
	);

	bfr new_net_15592_bfr_after (
		.din(new_net_15591),
		.dout(new_net_15592)
	);

	bfr new_net_15593_bfr_after (
		.din(new_net_15592),
		.dout(new_net_15593)
	);

	bfr new_net_15594_bfr_after (
		.din(new_net_15593),
		.dout(new_net_15594)
	);

	bfr new_net_15595_bfr_after (
		.din(new_net_15594),
		.dout(new_net_15595)
	);

	bfr new_net_15596_bfr_after (
		.din(new_net_15595),
		.dout(new_net_15596)
	);

	bfr new_net_15597_bfr_after (
		.din(new_net_15596),
		.dout(new_net_15597)
	);

	bfr new_net_15598_bfr_after (
		.din(new_net_15597),
		.dout(new_net_15598)
	);

	bfr new_net_15599_bfr_after (
		.din(new_net_15598),
		.dout(new_net_15599)
	);

	bfr new_net_15600_bfr_after (
		.din(new_net_15599),
		.dout(new_net_15600)
	);

	bfr new_net_15601_bfr_after (
		.din(new_net_15600),
		.dout(new_net_15601)
	);

	bfr new_net_15602_bfr_after (
		.din(new_net_15601),
		.dout(new_net_15602)
	);

	bfr new_net_15603_bfr_after (
		.din(new_net_15602),
		.dout(new_net_15603)
	);

	bfr new_net_15604_bfr_after (
		.din(new_net_15603),
		.dout(new_net_15604)
	);

	bfr new_net_15605_bfr_after (
		.din(new_net_15604),
		.dout(new_net_15605)
	);

	bfr new_net_15606_bfr_after (
		.din(new_net_15605),
		.dout(new_net_15606)
	);

	spl2 _1284__v_fanout (
		.a(new_net_15606),
		.b(new_net_366),
		.c(new_net_367)
	);

	bfr new_net_15607_bfr_after (
		.din(_0221_),
		.dout(new_net_15607)
	);

	bfr new_net_15608_bfr_after (
		.din(new_net_15607),
		.dout(new_net_15608)
	);

	bfr new_net_15609_bfr_after (
		.din(new_net_15608),
		.dout(new_net_15609)
	);

	bfr new_net_15610_bfr_after (
		.din(new_net_15609),
		.dout(new_net_15610)
	);

	bfr new_net_15611_bfr_after (
		.din(new_net_15610),
		.dout(new_net_15611)
	);

	bfr new_net_15612_bfr_after (
		.din(new_net_15611),
		.dout(new_net_15612)
	);

	bfr new_net_15613_bfr_after (
		.din(new_net_15612),
		.dout(new_net_15613)
	);

	bfr new_net_15614_bfr_after (
		.din(new_net_15613),
		.dout(new_net_15614)
	);

	bfr new_net_15615_bfr_after (
		.din(new_net_15614),
		.dout(new_net_15615)
	);

	bfr new_net_15616_bfr_after (
		.din(new_net_15615),
		.dout(new_net_15616)
	);

	bfr new_net_15617_bfr_after (
		.din(new_net_15616),
		.dout(new_net_15617)
	);

	bfr new_net_15618_bfr_after (
		.din(new_net_15617),
		.dout(new_net_15618)
	);

	bfr new_net_15619_bfr_after (
		.din(new_net_15618),
		.dout(new_net_15619)
	);

	bfr new_net_15620_bfr_after (
		.din(new_net_15619),
		.dout(new_net_15620)
	);

	bfr new_net_15621_bfr_after (
		.din(new_net_15620),
		.dout(new_net_15621)
	);

	bfr new_net_15622_bfr_after (
		.din(new_net_15621),
		.dout(new_net_15622)
	);

	bfr new_net_15623_bfr_after (
		.din(new_net_15622),
		.dout(new_net_15623)
	);

	bfr new_net_15624_bfr_after (
		.din(new_net_15623),
		.dout(new_net_15624)
	);

	bfr new_net_15625_bfr_after (
		.din(new_net_15624),
		.dout(new_net_15625)
	);

	bfr new_net_15626_bfr_after (
		.din(new_net_15625),
		.dout(new_net_15626)
	);

	bfr new_net_15627_bfr_after (
		.din(new_net_15626),
		.dout(new_net_15627)
	);

	bfr new_net_15628_bfr_after (
		.din(new_net_15627),
		.dout(new_net_15628)
	);

	bfr new_net_15629_bfr_after (
		.din(new_net_15628),
		.dout(new_net_15629)
	);

	bfr new_net_15630_bfr_after (
		.din(new_net_15629),
		.dout(new_net_15630)
	);

	bfr new_net_15631_bfr_after (
		.din(new_net_15630),
		.dout(new_net_15631)
	);

	bfr new_net_15632_bfr_after (
		.din(new_net_15631),
		.dout(new_net_15632)
	);

	bfr new_net_15633_bfr_after (
		.din(new_net_15632),
		.dout(new_net_15633)
	);

	bfr new_net_15634_bfr_after (
		.din(new_net_15633),
		.dout(new_net_15634)
	);

	bfr new_net_15635_bfr_after (
		.din(new_net_15634),
		.dout(new_net_15635)
	);

	bfr new_net_15636_bfr_after (
		.din(new_net_15635),
		.dout(new_net_15636)
	);

	bfr new_net_15637_bfr_after (
		.din(new_net_15636),
		.dout(new_net_15637)
	);

	bfr new_net_15638_bfr_after (
		.din(new_net_15637),
		.dout(new_net_15638)
	);

	bfr new_net_15639_bfr_after (
		.din(new_net_15638),
		.dout(new_net_15639)
	);

	bfr new_net_15640_bfr_after (
		.din(new_net_15639),
		.dout(new_net_15640)
	);

	bfr new_net_15641_bfr_after (
		.din(new_net_15640),
		.dout(new_net_15641)
	);

	bfr new_net_15642_bfr_after (
		.din(new_net_15641),
		.dout(new_net_15642)
	);

	bfr new_net_15643_bfr_after (
		.din(new_net_15642),
		.dout(new_net_15643)
	);

	bfr new_net_15644_bfr_after (
		.din(new_net_15643),
		.dout(new_net_15644)
	);

	bfr new_net_15645_bfr_after (
		.din(new_net_15644),
		.dout(new_net_15645)
	);

	bfr new_net_15646_bfr_after (
		.din(new_net_15645),
		.dout(new_net_15646)
	);

	bfr new_net_15647_bfr_after (
		.din(new_net_15646),
		.dout(new_net_15647)
	);

	bfr new_net_15648_bfr_after (
		.din(new_net_15647),
		.dout(new_net_15648)
	);

	bfr new_net_15649_bfr_after (
		.din(new_net_15648),
		.dout(new_net_15649)
	);

	bfr new_net_15650_bfr_after (
		.din(new_net_15649),
		.dout(new_net_15650)
	);

	bfr new_net_15651_bfr_after (
		.din(new_net_15650),
		.dout(new_net_15651)
	);

	bfr new_net_15652_bfr_after (
		.din(new_net_15651),
		.dout(new_net_15652)
	);

	bfr new_net_15653_bfr_after (
		.din(new_net_15652),
		.dout(new_net_15653)
	);

	bfr new_net_15654_bfr_after (
		.din(new_net_15653),
		.dout(new_net_15654)
	);

	bfr new_net_15655_bfr_after (
		.din(new_net_15654),
		.dout(new_net_15655)
	);

	bfr new_net_15656_bfr_after (
		.din(new_net_15655),
		.dout(new_net_15656)
	);

	bfr new_net_15657_bfr_after (
		.din(new_net_15656),
		.dout(new_net_15657)
	);

	bfr new_net_15658_bfr_after (
		.din(new_net_15657),
		.dout(new_net_15658)
	);

	bfr new_net_15659_bfr_after (
		.din(new_net_15658),
		.dout(new_net_15659)
	);

	bfr new_net_15660_bfr_after (
		.din(new_net_15659),
		.dout(new_net_15660)
	);

	bfr new_net_15661_bfr_after (
		.din(new_net_15660),
		.dout(new_net_15661)
	);

	bfr new_net_15662_bfr_after (
		.din(new_net_15661),
		.dout(new_net_15662)
	);

	bfr new_net_15663_bfr_after (
		.din(new_net_15662),
		.dout(new_net_15663)
	);

	bfr new_net_15664_bfr_after (
		.din(new_net_15663),
		.dout(new_net_15664)
	);

	bfr new_net_15665_bfr_after (
		.din(new_net_15664),
		.dout(new_net_15665)
	);

	bfr new_net_15666_bfr_after (
		.din(new_net_15665),
		.dout(new_net_15666)
	);

	bfr new_net_15667_bfr_after (
		.din(new_net_15666),
		.dout(new_net_15667)
	);

	bfr new_net_15668_bfr_after (
		.din(new_net_15667),
		.dout(new_net_15668)
	);

	bfr new_net_15669_bfr_after (
		.din(new_net_15668),
		.dout(new_net_15669)
	);

	bfr new_net_15670_bfr_after (
		.din(new_net_15669),
		.dout(new_net_15670)
	);

	bfr new_net_15671_bfr_after (
		.din(new_net_15670),
		.dout(new_net_15671)
	);

	bfr new_net_15672_bfr_after (
		.din(new_net_15671),
		.dout(new_net_15672)
	);

	bfr new_net_15673_bfr_after (
		.din(new_net_15672),
		.dout(new_net_15673)
	);

	bfr new_net_15674_bfr_after (
		.din(new_net_15673),
		.dout(new_net_15674)
	);

	bfr new_net_15675_bfr_after (
		.din(new_net_15674),
		.dout(new_net_15675)
	);

	bfr new_net_15676_bfr_after (
		.din(new_net_15675),
		.dout(new_net_15676)
	);

	bfr new_net_15677_bfr_after (
		.din(new_net_15676),
		.dout(new_net_15677)
	);

	bfr new_net_15678_bfr_after (
		.din(new_net_15677),
		.dout(new_net_15678)
	);

	bfr new_net_15679_bfr_after (
		.din(new_net_15678),
		.dout(new_net_15679)
	);

	bfr new_net_15680_bfr_after (
		.din(new_net_15679),
		.dout(new_net_15680)
	);

	bfr new_net_15681_bfr_after (
		.din(new_net_15680),
		.dout(new_net_15681)
	);

	bfr new_net_15682_bfr_after (
		.din(new_net_15681),
		.dout(new_net_15682)
	);

	bfr new_net_15683_bfr_after (
		.din(new_net_15682),
		.dout(new_net_15683)
	);

	bfr new_net_15684_bfr_after (
		.din(new_net_15683),
		.dout(new_net_15684)
	);

	bfr new_net_15685_bfr_after (
		.din(new_net_15684),
		.dout(new_net_15685)
	);

	bfr new_net_15686_bfr_after (
		.din(new_net_15685),
		.dout(new_net_15686)
	);

	spl2 _0221__v_fanout (
		.a(new_net_15686),
		.b(new_net_110),
		.c(new_net_111)
	);

	bfr new_net_15687_bfr_after (
		.din(_0531_),
		.dout(new_net_15687)
	);

	bfr new_net_15688_bfr_after (
		.din(new_net_15687),
		.dout(new_net_15688)
	);

	bfr new_net_15689_bfr_after (
		.din(new_net_15688),
		.dout(new_net_15689)
	);

	bfr new_net_15690_bfr_after (
		.din(new_net_15689),
		.dout(new_net_15690)
	);

	bfr new_net_15691_bfr_after (
		.din(new_net_15690),
		.dout(new_net_15691)
	);

	bfr new_net_15692_bfr_after (
		.din(new_net_15691),
		.dout(new_net_15692)
	);

	bfr new_net_15693_bfr_after (
		.din(new_net_15692),
		.dout(new_net_15693)
	);

	bfr new_net_15694_bfr_after (
		.din(new_net_15693),
		.dout(new_net_15694)
	);

	bfr new_net_15695_bfr_after (
		.din(new_net_15694),
		.dout(new_net_15695)
	);

	bfr new_net_15696_bfr_after (
		.din(new_net_15695),
		.dout(new_net_15696)
	);

	bfr new_net_15697_bfr_after (
		.din(new_net_15696),
		.dout(new_net_15697)
	);

	bfr new_net_15698_bfr_after (
		.din(new_net_15697),
		.dout(new_net_15698)
	);

	bfr new_net_15699_bfr_after (
		.din(new_net_15698),
		.dout(new_net_15699)
	);

	bfr new_net_15700_bfr_after (
		.din(new_net_15699),
		.dout(new_net_15700)
	);

	bfr new_net_15701_bfr_after (
		.din(new_net_15700),
		.dout(new_net_15701)
	);

	bfr new_net_15702_bfr_after (
		.din(new_net_15701),
		.dout(new_net_15702)
	);

	bfr new_net_15703_bfr_after (
		.din(new_net_15702),
		.dout(new_net_15703)
	);

	bfr new_net_15704_bfr_after (
		.din(new_net_15703),
		.dout(new_net_15704)
	);

	bfr new_net_15705_bfr_after (
		.din(new_net_15704),
		.dout(new_net_15705)
	);

	bfr new_net_15706_bfr_after (
		.din(new_net_15705),
		.dout(new_net_15706)
	);

	bfr new_net_15707_bfr_after (
		.din(new_net_15706),
		.dout(new_net_15707)
	);

	bfr new_net_15708_bfr_after (
		.din(new_net_15707),
		.dout(new_net_15708)
	);

	bfr new_net_15709_bfr_after (
		.din(new_net_15708),
		.dout(new_net_15709)
	);

	bfr new_net_15710_bfr_after (
		.din(new_net_15709),
		.dout(new_net_15710)
	);

	bfr new_net_15711_bfr_after (
		.din(new_net_15710),
		.dout(new_net_15711)
	);

	bfr new_net_15712_bfr_after (
		.din(new_net_15711),
		.dout(new_net_15712)
	);

	bfr new_net_15713_bfr_after (
		.din(new_net_15712),
		.dout(new_net_15713)
	);

	bfr new_net_15714_bfr_after (
		.din(new_net_15713),
		.dout(new_net_15714)
	);

	bfr new_net_15715_bfr_after (
		.din(new_net_15714),
		.dout(new_net_15715)
	);

	bfr new_net_15716_bfr_after (
		.din(new_net_15715),
		.dout(new_net_15716)
	);

	bfr new_net_15717_bfr_after (
		.din(new_net_15716),
		.dout(new_net_15717)
	);

	bfr new_net_15718_bfr_after (
		.din(new_net_15717),
		.dout(new_net_15718)
	);

	bfr new_net_15719_bfr_after (
		.din(new_net_15718),
		.dout(new_net_15719)
	);

	bfr new_net_15720_bfr_after (
		.din(new_net_15719),
		.dout(new_net_15720)
	);

	bfr new_net_15721_bfr_after (
		.din(new_net_15720),
		.dout(new_net_15721)
	);

	bfr new_net_15722_bfr_after (
		.din(new_net_15721),
		.dout(new_net_15722)
	);

	bfr new_net_15723_bfr_after (
		.din(new_net_15722),
		.dout(new_net_15723)
	);

	bfr new_net_15724_bfr_after (
		.din(new_net_15723),
		.dout(new_net_15724)
	);

	bfr new_net_15725_bfr_after (
		.din(new_net_15724),
		.dout(new_net_15725)
	);

	bfr new_net_15726_bfr_after (
		.din(new_net_15725),
		.dout(new_net_15726)
	);

	bfr new_net_15727_bfr_after (
		.din(new_net_15726),
		.dout(new_net_15727)
	);

	bfr new_net_15728_bfr_after (
		.din(new_net_15727),
		.dout(new_net_15728)
	);

	bfr new_net_15729_bfr_after (
		.din(new_net_15728),
		.dout(new_net_15729)
	);

	bfr new_net_15730_bfr_after (
		.din(new_net_15729),
		.dout(new_net_15730)
	);

	bfr new_net_15731_bfr_after (
		.din(new_net_15730),
		.dout(new_net_15731)
	);

	bfr new_net_15732_bfr_after (
		.din(new_net_15731),
		.dout(new_net_15732)
	);

	bfr new_net_15733_bfr_after (
		.din(new_net_15732),
		.dout(new_net_15733)
	);

	bfr new_net_15734_bfr_after (
		.din(new_net_15733),
		.dout(new_net_15734)
	);

	bfr new_net_15735_bfr_after (
		.din(new_net_15734),
		.dout(new_net_15735)
	);

	bfr new_net_15736_bfr_after (
		.din(new_net_15735),
		.dout(new_net_15736)
	);

	bfr new_net_15737_bfr_after (
		.din(new_net_15736),
		.dout(new_net_15737)
	);

	bfr new_net_15738_bfr_after (
		.din(new_net_15737),
		.dout(new_net_15738)
	);

	bfr new_net_15739_bfr_after (
		.din(new_net_15738),
		.dout(new_net_15739)
	);

	bfr new_net_15740_bfr_after (
		.din(new_net_15739),
		.dout(new_net_15740)
	);

	bfr new_net_15741_bfr_after (
		.din(new_net_15740),
		.dout(new_net_15741)
	);

	bfr new_net_15742_bfr_after (
		.din(new_net_15741),
		.dout(new_net_15742)
	);

	bfr new_net_15743_bfr_after (
		.din(new_net_15742),
		.dout(new_net_15743)
	);

	bfr new_net_15744_bfr_after (
		.din(new_net_15743),
		.dout(new_net_15744)
	);

	bfr new_net_15745_bfr_after (
		.din(new_net_15744),
		.dout(new_net_15745)
	);

	bfr new_net_15746_bfr_after (
		.din(new_net_15745),
		.dout(new_net_15746)
	);

	bfr new_net_15747_bfr_after (
		.din(new_net_15746),
		.dout(new_net_15747)
	);

	bfr new_net_15748_bfr_after (
		.din(new_net_15747),
		.dout(new_net_15748)
	);

	bfr new_net_15749_bfr_after (
		.din(new_net_15748),
		.dout(new_net_15749)
	);

	bfr new_net_15750_bfr_after (
		.din(new_net_15749),
		.dout(new_net_15750)
	);

	bfr new_net_15751_bfr_after (
		.din(new_net_15750),
		.dout(new_net_15751)
	);

	bfr new_net_15752_bfr_after (
		.din(new_net_15751),
		.dout(new_net_15752)
	);

	bfr new_net_15753_bfr_after (
		.din(new_net_15752),
		.dout(new_net_15753)
	);

	bfr new_net_15754_bfr_after (
		.din(new_net_15753),
		.dout(new_net_15754)
	);

	bfr new_net_15755_bfr_after (
		.din(new_net_15754),
		.dout(new_net_15755)
	);

	bfr new_net_15756_bfr_after (
		.din(new_net_15755),
		.dout(new_net_15756)
	);

	bfr new_net_15757_bfr_after (
		.din(new_net_15756),
		.dout(new_net_15757)
	);

	bfr new_net_15758_bfr_after (
		.din(new_net_15757),
		.dout(new_net_15758)
	);

	bfr new_net_15759_bfr_after (
		.din(new_net_15758),
		.dout(new_net_15759)
	);

	bfr new_net_15760_bfr_after (
		.din(new_net_15759),
		.dout(new_net_15760)
	);

	bfr new_net_15761_bfr_after (
		.din(new_net_15760),
		.dout(new_net_15761)
	);

	bfr new_net_15762_bfr_after (
		.din(new_net_15761),
		.dout(new_net_15762)
	);

	bfr new_net_15763_bfr_after (
		.din(new_net_15762),
		.dout(new_net_15763)
	);

	bfr new_net_15764_bfr_after (
		.din(new_net_15763),
		.dout(new_net_15764)
	);

	bfr new_net_15765_bfr_after (
		.din(new_net_15764),
		.dout(new_net_15765)
	);

	bfr new_net_15766_bfr_after (
		.din(new_net_15765),
		.dout(new_net_15766)
	);

	bfr new_net_15767_bfr_after (
		.din(new_net_15766),
		.dout(new_net_15767)
	);

	bfr new_net_15768_bfr_after (
		.din(new_net_15767),
		.dout(new_net_15768)
	);

	bfr new_net_15769_bfr_after (
		.din(new_net_15768),
		.dout(new_net_15769)
	);

	bfr new_net_15770_bfr_after (
		.din(new_net_15769),
		.dout(new_net_15770)
	);

	bfr new_net_15771_bfr_after (
		.din(new_net_15770),
		.dout(new_net_15771)
	);

	bfr new_net_15772_bfr_after (
		.din(new_net_15771),
		.dout(new_net_15772)
	);

	bfr new_net_15773_bfr_after (
		.din(new_net_15772),
		.dout(new_net_15773)
	);

	bfr new_net_15774_bfr_after (
		.din(new_net_15773),
		.dout(new_net_15774)
	);

	bfr new_net_15775_bfr_after (
		.din(new_net_15774),
		.dout(new_net_15775)
	);

	bfr new_net_15776_bfr_after (
		.din(new_net_15775),
		.dout(new_net_15776)
	);

	bfr new_net_15777_bfr_after (
		.din(new_net_15776),
		.dout(new_net_15777)
	);

	bfr new_net_15778_bfr_after (
		.din(new_net_15777),
		.dout(new_net_15778)
	);

	bfr new_net_15779_bfr_after (
		.din(new_net_15778),
		.dout(new_net_15779)
	);

	bfr new_net_15780_bfr_after (
		.din(new_net_15779),
		.dout(new_net_15780)
	);

	bfr new_net_15781_bfr_after (
		.din(new_net_15780),
		.dout(new_net_15781)
	);

	bfr new_net_15782_bfr_after (
		.din(new_net_15781),
		.dout(new_net_15782)
	);

	bfr new_net_15783_bfr_after (
		.din(new_net_15782),
		.dout(new_net_15783)
	);

	bfr new_net_15784_bfr_after (
		.din(new_net_15783),
		.dout(new_net_15784)
	);

	bfr new_net_15785_bfr_after (
		.din(new_net_15784),
		.dout(new_net_15785)
	);

	bfr new_net_15786_bfr_after (
		.din(new_net_15785),
		.dout(new_net_15786)
	);

	bfr new_net_15787_bfr_after (
		.din(new_net_15786),
		.dout(new_net_15787)
	);

	bfr new_net_15788_bfr_after (
		.din(new_net_15787),
		.dout(new_net_15788)
	);

	bfr new_net_15789_bfr_after (
		.din(new_net_15788),
		.dout(new_net_15789)
	);

	bfr new_net_15790_bfr_after (
		.din(new_net_15789),
		.dout(new_net_15790)
	);

	spl2 _0531__v_fanout (
		.a(new_net_15790),
		.b(new_net_2060),
		.c(new_net_2061)
	);

	bfr new_net_15791_bfr_after (
		.din(_0533_),
		.dout(new_net_15791)
	);

	bfr new_net_15792_bfr_after (
		.din(new_net_15791),
		.dout(new_net_15792)
	);

	bfr new_net_15793_bfr_after (
		.din(new_net_15792),
		.dout(new_net_15793)
	);

	bfr new_net_15794_bfr_after (
		.din(new_net_15793),
		.dout(new_net_15794)
	);

	bfr new_net_15795_bfr_after (
		.din(new_net_15794),
		.dout(new_net_15795)
	);

	bfr new_net_15796_bfr_after (
		.din(new_net_15795),
		.dout(new_net_15796)
	);

	bfr new_net_15797_bfr_after (
		.din(new_net_15796),
		.dout(new_net_15797)
	);

	bfr new_net_15798_bfr_after (
		.din(new_net_15797),
		.dout(new_net_15798)
	);

	bfr new_net_15799_bfr_after (
		.din(new_net_15798),
		.dout(new_net_15799)
	);

	bfr new_net_15800_bfr_after (
		.din(new_net_15799),
		.dout(new_net_15800)
	);

	bfr new_net_15801_bfr_after (
		.din(new_net_15800),
		.dout(new_net_15801)
	);

	bfr new_net_15802_bfr_after (
		.din(new_net_15801),
		.dout(new_net_15802)
	);

	bfr new_net_15803_bfr_after (
		.din(new_net_15802),
		.dout(new_net_15803)
	);

	bfr new_net_15804_bfr_after (
		.din(new_net_15803),
		.dout(new_net_15804)
	);

	bfr new_net_15805_bfr_after (
		.din(new_net_15804),
		.dout(new_net_15805)
	);

	bfr new_net_15806_bfr_after (
		.din(new_net_15805),
		.dout(new_net_15806)
	);

	bfr new_net_15807_bfr_after (
		.din(new_net_15806),
		.dout(new_net_15807)
	);

	bfr new_net_15808_bfr_after (
		.din(new_net_15807),
		.dout(new_net_15808)
	);

	bfr new_net_15809_bfr_after (
		.din(new_net_15808),
		.dout(new_net_15809)
	);

	bfr new_net_15810_bfr_after (
		.din(new_net_15809),
		.dout(new_net_15810)
	);

	bfr new_net_15811_bfr_after (
		.din(new_net_15810),
		.dout(new_net_15811)
	);

	bfr new_net_15812_bfr_after (
		.din(new_net_15811),
		.dout(new_net_15812)
	);

	bfr new_net_15813_bfr_after (
		.din(new_net_15812),
		.dout(new_net_15813)
	);

	bfr new_net_15814_bfr_after (
		.din(new_net_15813),
		.dout(new_net_15814)
	);

	bfr new_net_15815_bfr_after (
		.din(new_net_15814),
		.dout(new_net_15815)
	);

	bfr new_net_15816_bfr_after (
		.din(new_net_15815),
		.dout(new_net_15816)
	);

	bfr new_net_15817_bfr_after (
		.din(new_net_15816),
		.dout(new_net_15817)
	);

	bfr new_net_15818_bfr_after (
		.din(new_net_15817),
		.dout(new_net_15818)
	);

	bfr new_net_15819_bfr_after (
		.din(new_net_15818),
		.dout(new_net_15819)
	);

	bfr new_net_15820_bfr_after (
		.din(new_net_15819),
		.dout(new_net_15820)
	);

	bfr new_net_15821_bfr_after (
		.din(new_net_15820),
		.dout(new_net_15821)
	);

	bfr new_net_15822_bfr_after (
		.din(new_net_15821),
		.dout(new_net_15822)
	);

	bfr new_net_15823_bfr_after (
		.din(new_net_15822),
		.dout(new_net_15823)
	);

	bfr new_net_15824_bfr_after (
		.din(new_net_15823),
		.dout(new_net_15824)
	);

	bfr new_net_15825_bfr_after (
		.din(new_net_15824),
		.dout(new_net_15825)
	);

	bfr new_net_15826_bfr_after (
		.din(new_net_15825),
		.dout(new_net_15826)
	);

	bfr new_net_15827_bfr_after (
		.din(new_net_15826),
		.dout(new_net_15827)
	);

	bfr new_net_15828_bfr_after (
		.din(new_net_15827),
		.dout(new_net_15828)
	);

	bfr new_net_15829_bfr_after (
		.din(new_net_15828),
		.dout(new_net_15829)
	);

	bfr new_net_15830_bfr_after (
		.din(new_net_15829),
		.dout(new_net_15830)
	);

	bfr new_net_15831_bfr_after (
		.din(new_net_15830),
		.dout(new_net_15831)
	);

	bfr new_net_15832_bfr_after (
		.din(new_net_15831),
		.dout(new_net_15832)
	);

	bfr new_net_15833_bfr_after (
		.din(new_net_15832),
		.dout(new_net_15833)
	);

	bfr new_net_15834_bfr_after (
		.din(new_net_15833),
		.dout(new_net_15834)
	);

	bfr new_net_15835_bfr_after (
		.din(new_net_15834),
		.dout(new_net_15835)
	);

	bfr new_net_15836_bfr_after (
		.din(new_net_15835),
		.dout(new_net_15836)
	);

	bfr new_net_15837_bfr_after (
		.din(new_net_15836),
		.dout(new_net_15837)
	);

	bfr new_net_15838_bfr_after (
		.din(new_net_15837),
		.dout(new_net_15838)
	);

	bfr new_net_15839_bfr_after (
		.din(new_net_15838),
		.dout(new_net_15839)
	);

	bfr new_net_15840_bfr_after (
		.din(new_net_15839),
		.dout(new_net_15840)
	);

	bfr new_net_15841_bfr_after (
		.din(new_net_15840),
		.dout(new_net_15841)
	);

	bfr new_net_15842_bfr_after (
		.din(new_net_15841),
		.dout(new_net_15842)
	);

	bfr new_net_15843_bfr_after (
		.din(new_net_15842),
		.dout(new_net_15843)
	);

	bfr new_net_15844_bfr_after (
		.din(new_net_15843),
		.dout(new_net_15844)
	);

	bfr new_net_15845_bfr_after (
		.din(new_net_15844),
		.dout(new_net_15845)
	);

	bfr new_net_15846_bfr_after (
		.din(new_net_15845),
		.dout(new_net_15846)
	);

	bfr new_net_15847_bfr_after (
		.din(new_net_15846),
		.dout(new_net_15847)
	);

	bfr new_net_15848_bfr_after (
		.din(new_net_15847),
		.dout(new_net_15848)
	);

	bfr new_net_15849_bfr_after (
		.din(new_net_15848),
		.dout(new_net_15849)
	);

	bfr new_net_15850_bfr_after (
		.din(new_net_15849),
		.dout(new_net_15850)
	);

	bfr new_net_15851_bfr_after (
		.din(new_net_15850),
		.dout(new_net_15851)
	);

	bfr new_net_15852_bfr_after (
		.din(new_net_15851),
		.dout(new_net_15852)
	);

	bfr new_net_15853_bfr_after (
		.din(new_net_15852),
		.dout(new_net_15853)
	);

	bfr new_net_15854_bfr_after (
		.din(new_net_15853),
		.dout(new_net_15854)
	);

	bfr new_net_15855_bfr_after (
		.din(new_net_15854),
		.dout(new_net_15855)
	);

	bfr new_net_15856_bfr_after (
		.din(new_net_15855),
		.dout(new_net_15856)
	);

	bfr new_net_15857_bfr_after (
		.din(new_net_15856),
		.dout(new_net_15857)
	);

	bfr new_net_15858_bfr_after (
		.din(new_net_15857),
		.dout(new_net_15858)
	);

	bfr new_net_15859_bfr_after (
		.din(new_net_15858),
		.dout(new_net_15859)
	);

	bfr new_net_15860_bfr_after (
		.din(new_net_15859),
		.dout(new_net_15860)
	);

	bfr new_net_15861_bfr_after (
		.din(new_net_15860),
		.dout(new_net_15861)
	);

	bfr new_net_15862_bfr_after (
		.din(new_net_15861),
		.dout(new_net_15862)
	);

	bfr new_net_15863_bfr_after (
		.din(new_net_15862),
		.dout(new_net_15863)
	);

	bfr new_net_15864_bfr_after (
		.din(new_net_15863),
		.dout(new_net_15864)
	);

	bfr new_net_15865_bfr_after (
		.din(new_net_15864),
		.dout(new_net_15865)
	);

	bfr new_net_15866_bfr_after (
		.din(new_net_15865),
		.dout(new_net_15866)
	);

	bfr new_net_15867_bfr_after (
		.din(new_net_15866),
		.dout(new_net_15867)
	);

	bfr new_net_15868_bfr_after (
		.din(new_net_15867),
		.dout(new_net_15868)
	);

	bfr new_net_15869_bfr_after (
		.din(new_net_15868),
		.dout(new_net_15869)
	);

	bfr new_net_15870_bfr_after (
		.din(new_net_15869),
		.dout(new_net_15870)
	);

	bfr new_net_15871_bfr_after (
		.din(new_net_15870),
		.dout(new_net_15871)
	);

	bfr new_net_15872_bfr_after (
		.din(new_net_15871),
		.dout(new_net_15872)
	);

	bfr new_net_15873_bfr_after (
		.din(new_net_15872),
		.dout(new_net_15873)
	);

	bfr new_net_15874_bfr_after (
		.din(new_net_15873),
		.dout(new_net_15874)
	);

	bfr new_net_15875_bfr_after (
		.din(new_net_15874),
		.dout(new_net_15875)
	);

	bfr new_net_15876_bfr_after (
		.din(new_net_15875),
		.dout(new_net_15876)
	);

	bfr new_net_15877_bfr_after (
		.din(new_net_15876),
		.dout(new_net_15877)
	);

	bfr new_net_15878_bfr_after (
		.din(new_net_15877),
		.dout(new_net_15878)
	);

	bfr new_net_15879_bfr_after (
		.din(new_net_15878),
		.dout(new_net_15879)
	);

	bfr new_net_15880_bfr_after (
		.din(new_net_15879),
		.dout(new_net_15880)
	);

	bfr new_net_15881_bfr_after (
		.din(new_net_15880),
		.dout(new_net_15881)
	);

	bfr new_net_15882_bfr_after (
		.din(new_net_15881),
		.dout(new_net_15882)
	);

	bfr new_net_15883_bfr_after (
		.din(new_net_15882),
		.dout(new_net_15883)
	);

	bfr new_net_15884_bfr_after (
		.din(new_net_15883),
		.dout(new_net_15884)
	);

	bfr new_net_15885_bfr_after (
		.din(new_net_15884),
		.dout(new_net_15885)
	);

	bfr new_net_15886_bfr_after (
		.din(new_net_15885),
		.dout(new_net_15886)
	);

	spl2 _0533__v_fanout (
		.a(new_net_15886),
		.b(new_net_2160),
		.c(new_net_2161)
	);

	bfr new_net_15887_bfr_before (
		.din(new_net_15887),
		.dout(new_net_1321)
	);

	bfr new_net_15888_bfr_before (
		.din(new_net_15888),
		.dout(new_net_15887)
	);

	bfr new_net_15889_bfr_before (
		.din(new_net_15889),
		.dout(new_net_15888)
	);

	bfr new_net_15890_bfr_before (
		.din(new_net_15890),
		.dout(new_net_15889)
	);

	spl2 _1830__v_fanout (
		.a(_1830_),
		.b(new_net_1320),
		.c(new_net_15890)
	);

	bfr new_net_15891_bfr_after (
		.din(_0928_),
		.dout(new_net_15891)
	);

	bfr new_net_15892_bfr_after (
		.din(new_net_15891),
		.dout(new_net_15892)
	);

	bfr new_net_15893_bfr_after (
		.din(new_net_15892),
		.dout(new_net_15893)
	);

	bfr new_net_15894_bfr_after (
		.din(new_net_15893),
		.dout(new_net_15894)
	);

	bfr new_net_15895_bfr_after (
		.din(new_net_15894),
		.dout(new_net_15895)
	);

	bfr new_net_15896_bfr_after (
		.din(new_net_15895),
		.dout(new_net_15896)
	);

	bfr new_net_15897_bfr_after (
		.din(new_net_15896),
		.dout(new_net_15897)
	);

	bfr new_net_15898_bfr_after (
		.din(new_net_15897),
		.dout(new_net_15898)
	);

	bfr new_net_15899_bfr_after (
		.din(new_net_15898),
		.dout(new_net_15899)
	);

	bfr new_net_15900_bfr_after (
		.din(new_net_15899),
		.dout(new_net_15900)
	);

	bfr new_net_15901_bfr_after (
		.din(new_net_15900),
		.dout(new_net_15901)
	);

	bfr new_net_15902_bfr_after (
		.din(new_net_15901),
		.dout(new_net_15902)
	);

	bfr new_net_15903_bfr_after (
		.din(new_net_15902),
		.dout(new_net_15903)
	);

	bfr new_net_15904_bfr_after (
		.din(new_net_15903),
		.dout(new_net_15904)
	);

	bfr new_net_15905_bfr_after (
		.din(new_net_15904),
		.dout(new_net_15905)
	);

	bfr new_net_15906_bfr_after (
		.din(new_net_15905),
		.dout(new_net_15906)
	);

	bfr new_net_15907_bfr_after (
		.din(new_net_15906),
		.dout(new_net_15907)
	);

	bfr new_net_15908_bfr_after (
		.din(new_net_15907),
		.dout(new_net_15908)
	);

	bfr new_net_15909_bfr_after (
		.din(new_net_15908),
		.dout(new_net_15909)
	);

	bfr new_net_15910_bfr_after (
		.din(new_net_15909),
		.dout(new_net_15910)
	);

	bfr new_net_15911_bfr_after (
		.din(new_net_15910),
		.dout(new_net_15911)
	);

	bfr new_net_15912_bfr_after (
		.din(new_net_15911),
		.dout(new_net_15912)
	);

	bfr new_net_15913_bfr_after (
		.din(new_net_15912),
		.dout(new_net_15913)
	);

	bfr new_net_15914_bfr_after (
		.din(new_net_15913),
		.dout(new_net_15914)
	);

	bfr new_net_15915_bfr_after (
		.din(new_net_15914),
		.dout(new_net_15915)
	);

	bfr new_net_15916_bfr_after (
		.din(new_net_15915),
		.dout(new_net_15916)
	);

	bfr new_net_15917_bfr_after (
		.din(new_net_15916),
		.dout(new_net_15917)
	);

	bfr new_net_15918_bfr_after (
		.din(new_net_15917),
		.dout(new_net_15918)
	);

	bfr new_net_15919_bfr_after (
		.din(new_net_15918),
		.dout(new_net_15919)
	);

	bfr new_net_15920_bfr_after (
		.din(new_net_15919),
		.dout(new_net_15920)
	);

	bfr new_net_15921_bfr_after (
		.din(new_net_15920),
		.dout(new_net_15921)
	);

	bfr new_net_15922_bfr_after (
		.din(new_net_15921),
		.dout(new_net_15922)
	);

	bfr new_net_15923_bfr_after (
		.din(new_net_15922),
		.dout(new_net_15923)
	);

	bfr new_net_15924_bfr_after (
		.din(new_net_15923),
		.dout(new_net_15924)
	);

	bfr new_net_15925_bfr_after (
		.din(new_net_15924),
		.dout(new_net_15925)
	);

	bfr new_net_15926_bfr_after (
		.din(new_net_15925),
		.dout(new_net_15926)
	);

	bfr new_net_15927_bfr_after (
		.din(new_net_15926),
		.dout(new_net_15927)
	);

	bfr new_net_15928_bfr_after (
		.din(new_net_15927),
		.dout(new_net_15928)
	);

	bfr new_net_15929_bfr_after (
		.din(new_net_15928),
		.dout(new_net_15929)
	);

	bfr new_net_15930_bfr_after (
		.din(new_net_15929),
		.dout(new_net_15930)
	);

	bfr new_net_15931_bfr_after (
		.din(new_net_15930),
		.dout(new_net_15931)
	);

	bfr new_net_15932_bfr_after (
		.din(new_net_15931),
		.dout(new_net_15932)
	);

	bfr new_net_15933_bfr_after (
		.din(new_net_15932),
		.dout(new_net_15933)
	);

	bfr new_net_15934_bfr_after (
		.din(new_net_15933),
		.dout(new_net_15934)
	);

	bfr new_net_15935_bfr_after (
		.din(new_net_15934),
		.dout(new_net_15935)
	);

	bfr new_net_15936_bfr_after (
		.din(new_net_15935),
		.dout(new_net_15936)
	);

	bfr new_net_15937_bfr_after (
		.din(new_net_15936),
		.dout(new_net_15937)
	);

	bfr new_net_15938_bfr_after (
		.din(new_net_15937),
		.dout(new_net_15938)
	);

	bfr new_net_15939_bfr_after (
		.din(new_net_15938),
		.dout(new_net_15939)
	);

	bfr new_net_15940_bfr_after (
		.din(new_net_15939),
		.dout(new_net_15940)
	);

	bfr new_net_15941_bfr_after (
		.din(new_net_15940),
		.dout(new_net_15941)
	);

	bfr new_net_15942_bfr_after (
		.din(new_net_15941),
		.dout(new_net_15942)
	);

	bfr new_net_15943_bfr_after (
		.din(new_net_15942),
		.dout(new_net_15943)
	);

	bfr new_net_15944_bfr_after (
		.din(new_net_15943),
		.dout(new_net_15944)
	);

	bfr new_net_15945_bfr_after (
		.din(new_net_15944),
		.dout(new_net_15945)
	);

	bfr new_net_15946_bfr_after (
		.din(new_net_15945),
		.dout(new_net_15946)
	);

	bfr new_net_15947_bfr_after (
		.din(new_net_15946),
		.dout(new_net_15947)
	);

	bfr new_net_15948_bfr_after (
		.din(new_net_15947),
		.dout(new_net_15948)
	);

	bfr new_net_15949_bfr_after (
		.din(new_net_15948),
		.dout(new_net_15949)
	);

	bfr new_net_15950_bfr_after (
		.din(new_net_15949),
		.dout(new_net_15950)
	);

	bfr new_net_15951_bfr_after (
		.din(new_net_15950),
		.dout(new_net_15951)
	);

	bfr new_net_15952_bfr_after (
		.din(new_net_15951),
		.dout(new_net_15952)
	);

	bfr new_net_15953_bfr_after (
		.din(new_net_15952),
		.dout(new_net_15953)
	);

	bfr new_net_15954_bfr_after (
		.din(new_net_15953),
		.dout(new_net_15954)
	);

	bfr new_net_15955_bfr_after (
		.din(new_net_15954),
		.dout(new_net_15955)
	);

	bfr new_net_15956_bfr_after (
		.din(new_net_15955),
		.dout(new_net_15956)
	);

	bfr new_net_15957_bfr_after (
		.din(new_net_15956),
		.dout(new_net_15957)
	);

	bfr new_net_15958_bfr_after (
		.din(new_net_15957),
		.dout(new_net_15958)
	);

	bfr new_net_15959_bfr_after (
		.din(new_net_15958),
		.dout(new_net_15959)
	);

	bfr new_net_15960_bfr_after (
		.din(new_net_15959),
		.dout(new_net_15960)
	);

	bfr new_net_15961_bfr_after (
		.din(new_net_15960),
		.dout(new_net_15961)
	);

	bfr new_net_15962_bfr_after (
		.din(new_net_15961),
		.dout(new_net_15962)
	);

	bfr new_net_15963_bfr_after (
		.din(new_net_15962),
		.dout(new_net_15963)
	);

	bfr new_net_15964_bfr_after (
		.din(new_net_15963),
		.dout(new_net_15964)
	);

	bfr new_net_15965_bfr_after (
		.din(new_net_15964),
		.dout(new_net_15965)
	);

	bfr new_net_15966_bfr_after (
		.din(new_net_15965),
		.dout(new_net_15966)
	);

	bfr new_net_15967_bfr_after (
		.din(new_net_15966),
		.dout(new_net_15967)
	);

	bfr new_net_15968_bfr_after (
		.din(new_net_15967),
		.dout(new_net_15968)
	);

	bfr new_net_15969_bfr_after (
		.din(new_net_15968),
		.dout(new_net_15969)
	);

	bfr new_net_15970_bfr_after (
		.din(new_net_15969),
		.dout(new_net_15970)
	);

	bfr new_net_15971_bfr_after (
		.din(new_net_15970),
		.dout(new_net_15971)
	);

	bfr new_net_15972_bfr_after (
		.din(new_net_15971),
		.dout(new_net_15972)
	);

	bfr new_net_15973_bfr_after (
		.din(new_net_15972),
		.dout(new_net_15973)
	);

	bfr new_net_15974_bfr_after (
		.din(new_net_15973),
		.dout(new_net_15974)
	);

	bfr new_net_15975_bfr_after (
		.din(new_net_15974),
		.dout(new_net_15975)
	);

	bfr new_net_15976_bfr_after (
		.din(new_net_15975),
		.dout(new_net_15976)
	);

	bfr new_net_15977_bfr_after (
		.din(new_net_15976),
		.dout(new_net_15977)
	);

	bfr new_net_15978_bfr_after (
		.din(new_net_15977),
		.dout(new_net_15978)
	);

	bfr new_net_15979_bfr_after (
		.din(new_net_15978),
		.dout(new_net_15979)
	);

	bfr new_net_15980_bfr_after (
		.din(new_net_15979),
		.dout(new_net_15980)
	);

	bfr new_net_15981_bfr_after (
		.din(new_net_15980),
		.dout(new_net_15981)
	);

	bfr new_net_15982_bfr_after (
		.din(new_net_15981),
		.dout(new_net_15982)
	);

	bfr new_net_15983_bfr_after (
		.din(new_net_15982),
		.dout(new_net_15983)
	);

	bfr new_net_15984_bfr_after (
		.din(new_net_15983),
		.dout(new_net_15984)
	);

	bfr new_net_15985_bfr_after (
		.din(new_net_15984),
		.dout(new_net_15985)
	);

	bfr new_net_15986_bfr_after (
		.din(new_net_15985),
		.dout(new_net_15986)
	);

	bfr new_net_15987_bfr_after (
		.din(new_net_15986),
		.dout(new_net_15987)
	);

	bfr new_net_15988_bfr_after (
		.din(new_net_15987),
		.dout(new_net_15988)
	);

	bfr new_net_15989_bfr_after (
		.din(new_net_15988),
		.dout(new_net_15989)
	);

	bfr new_net_15990_bfr_after (
		.din(new_net_15989),
		.dout(new_net_15990)
	);

	bfr new_net_15991_bfr_after (
		.din(new_net_15990),
		.dout(new_net_15991)
	);

	bfr new_net_15992_bfr_after (
		.din(new_net_15991),
		.dout(new_net_15992)
	);

	spl2 _0928__v_fanout (
		.a(new_net_15992),
		.b(new_net_1176),
		.c(new_net_1177)
	);

	bfr new_net_15993_bfr_after (
		.din(_1564_),
		.dout(new_net_15993)
	);

	bfr new_net_15994_bfr_after (
		.din(new_net_15993),
		.dout(new_net_15994)
	);

	bfr new_net_15995_bfr_after (
		.din(new_net_15994),
		.dout(new_net_15995)
	);

	bfr new_net_15996_bfr_after (
		.din(new_net_15995),
		.dout(new_net_15996)
	);

	bfr new_net_15997_bfr_after (
		.din(new_net_15996),
		.dout(new_net_15997)
	);

	bfr new_net_15998_bfr_after (
		.din(new_net_15997),
		.dout(new_net_15998)
	);

	bfr new_net_15999_bfr_after (
		.din(new_net_15998),
		.dout(new_net_15999)
	);

	bfr new_net_16000_bfr_after (
		.din(new_net_15999),
		.dout(new_net_16000)
	);

	bfr new_net_16001_bfr_after (
		.din(new_net_16000),
		.dout(new_net_16001)
	);

	bfr new_net_16002_bfr_after (
		.din(new_net_16001),
		.dout(new_net_16002)
	);

	bfr new_net_16003_bfr_after (
		.din(new_net_16002),
		.dout(new_net_16003)
	);

	bfr new_net_16004_bfr_after (
		.din(new_net_16003),
		.dout(new_net_16004)
	);

	bfr new_net_16005_bfr_after (
		.din(new_net_16004),
		.dout(new_net_16005)
	);

	bfr new_net_16006_bfr_after (
		.din(new_net_16005),
		.dout(new_net_16006)
	);

	bfr new_net_16007_bfr_after (
		.din(new_net_16006),
		.dout(new_net_16007)
	);

	bfr new_net_16008_bfr_after (
		.din(new_net_16007),
		.dout(new_net_16008)
	);

	bfr new_net_16009_bfr_after (
		.din(new_net_16008),
		.dout(new_net_16009)
	);

	bfr new_net_16010_bfr_after (
		.din(new_net_16009),
		.dout(new_net_16010)
	);

	bfr new_net_16011_bfr_after (
		.din(new_net_16010),
		.dout(new_net_16011)
	);

	bfr new_net_16012_bfr_after (
		.din(new_net_16011),
		.dout(new_net_16012)
	);

	bfr new_net_16013_bfr_after (
		.din(new_net_16012),
		.dout(new_net_16013)
	);

	bfr new_net_16014_bfr_after (
		.din(new_net_16013),
		.dout(new_net_16014)
	);

	bfr new_net_16015_bfr_after (
		.din(new_net_16014),
		.dout(new_net_16015)
	);

	bfr new_net_16016_bfr_after (
		.din(new_net_16015),
		.dout(new_net_16016)
	);

	bfr new_net_16017_bfr_after (
		.din(new_net_16016),
		.dout(new_net_16017)
	);

	bfr new_net_16018_bfr_after (
		.din(new_net_16017),
		.dout(new_net_16018)
	);

	bfr new_net_16019_bfr_after (
		.din(new_net_16018),
		.dout(new_net_16019)
	);

	bfr new_net_16020_bfr_after (
		.din(new_net_16019),
		.dout(new_net_16020)
	);

	bfr new_net_16021_bfr_after (
		.din(new_net_16020),
		.dout(new_net_16021)
	);

	bfr new_net_16022_bfr_after (
		.din(new_net_16021),
		.dout(new_net_16022)
	);

	bfr new_net_16023_bfr_after (
		.din(new_net_16022),
		.dout(new_net_16023)
	);

	bfr new_net_16024_bfr_after (
		.din(new_net_16023),
		.dout(new_net_16024)
	);

	bfr new_net_16025_bfr_after (
		.din(new_net_16024),
		.dout(new_net_16025)
	);

	bfr new_net_16026_bfr_after (
		.din(new_net_16025),
		.dout(new_net_16026)
	);

	bfr new_net_16027_bfr_after (
		.din(new_net_16026),
		.dout(new_net_16027)
	);

	bfr new_net_16028_bfr_after (
		.din(new_net_16027),
		.dout(new_net_16028)
	);

	bfr new_net_16029_bfr_after (
		.din(new_net_16028),
		.dout(new_net_16029)
	);

	bfr new_net_16030_bfr_after (
		.din(new_net_16029),
		.dout(new_net_16030)
	);

	bfr new_net_16031_bfr_after (
		.din(new_net_16030),
		.dout(new_net_16031)
	);

	bfr new_net_16032_bfr_after (
		.din(new_net_16031),
		.dout(new_net_16032)
	);

	bfr new_net_16033_bfr_after (
		.din(new_net_16032),
		.dout(new_net_16033)
	);

	bfr new_net_16034_bfr_after (
		.din(new_net_16033),
		.dout(new_net_16034)
	);

	bfr new_net_16035_bfr_after (
		.din(new_net_16034),
		.dout(new_net_16035)
	);

	bfr new_net_16036_bfr_after (
		.din(new_net_16035),
		.dout(new_net_16036)
	);

	bfr new_net_16037_bfr_after (
		.din(new_net_16036),
		.dout(new_net_16037)
	);

	bfr new_net_16038_bfr_after (
		.din(new_net_16037),
		.dout(new_net_16038)
	);

	bfr new_net_16039_bfr_after (
		.din(new_net_16038),
		.dout(new_net_16039)
	);

	bfr new_net_16040_bfr_after (
		.din(new_net_16039),
		.dout(new_net_16040)
	);

	bfr new_net_16041_bfr_after (
		.din(new_net_16040),
		.dout(new_net_16041)
	);

	bfr new_net_16042_bfr_after (
		.din(new_net_16041),
		.dout(new_net_16042)
	);

	bfr new_net_16043_bfr_after (
		.din(new_net_16042),
		.dout(new_net_16043)
	);

	bfr new_net_16044_bfr_after (
		.din(new_net_16043),
		.dout(new_net_16044)
	);

	bfr new_net_16045_bfr_after (
		.din(new_net_16044),
		.dout(new_net_16045)
	);

	bfr new_net_16046_bfr_after (
		.din(new_net_16045),
		.dout(new_net_16046)
	);

	bfr new_net_16047_bfr_after (
		.din(new_net_16046),
		.dout(new_net_16047)
	);

	bfr new_net_16048_bfr_after (
		.din(new_net_16047),
		.dout(new_net_16048)
	);

	bfr new_net_16049_bfr_after (
		.din(new_net_16048),
		.dout(new_net_16049)
	);

	bfr new_net_16050_bfr_after (
		.din(new_net_16049),
		.dout(new_net_16050)
	);

	bfr new_net_16051_bfr_after (
		.din(new_net_16050),
		.dout(new_net_16051)
	);

	bfr new_net_16052_bfr_after (
		.din(new_net_16051),
		.dout(new_net_16052)
	);

	bfr new_net_16053_bfr_after (
		.din(new_net_16052),
		.dout(new_net_16053)
	);

	bfr new_net_16054_bfr_after (
		.din(new_net_16053),
		.dout(new_net_16054)
	);

	bfr new_net_16055_bfr_after (
		.din(new_net_16054),
		.dout(new_net_16055)
	);

	bfr new_net_16056_bfr_after (
		.din(new_net_16055),
		.dout(new_net_16056)
	);

	bfr new_net_16057_bfr_after (
		.din(new_net_16056),
		.dout(new_net_16057)
	);

	bfr new_net_16058_bfr_after (
		.din(new_net_16057),
		.dout(new_net_16058)
	);

	bfr new_net_16059_bfr_after (
		.din(new_net_16058),
		.dout(new_net_16059)
	);

	bfr new_net_16060_bfr_after (
		.din(new_net_16059),
		.dout(new_net_16060)
	);

	bfr new_net_16061_bfr_after (
		.din(new_net_16060),
		.dout(new_net_16061)
	);

	bfr new_net_16062_bfr_after (
		.din(new_net_16061),
		.dout(new_net_16062)
	);

	bfr new_net_16063_bfr_after (
		.din(new_net_16062),
		.dout(new_net_16063)
	);

	bfr new_net_16064_bfr_after (
		.din(new_net_16063),
		.dout(new_net_16064)
	);

	bfr new_net_16065_bfr_after (
		.din(new_net_16064),
		.dout(new_net_16065)
	);

	bfr new_net_16066_bfr_after (
		.din(new_net_16065),
		.dout(new_net_16066)
	);

	bfr new_net_16067_bfr_after (
		.din(new_net_16066),
		.dout(new_net_16067)
	);

	bfr new_net_16068_bfr_after (
		.din(new_net_16067),
		.dout(new_net_16068)
	);

	bfr new_net_16069_bfr_after (
		.din(new_net_16068),
		.dout(new_net_16069)
	);

	bfr new_net_16070_bfr_after (
		.din(new_net_16069),
		.dout(new_net_16070)
	);

	bfr new_net_16071_bfr_after (
		.din(new_net_16070),
		.dout(new_net_16071)
	);

	bfr new_net_16072_bfr_after (
		.din(new_net_16071),
		.dout(new_net_16072)
	);

	bfr new_net_16073_bfr_after (
		.din(new_net_16072),
		.dout(new_net_16073)
	);

	bfr new_net_16074_bfr_after (
		.din(new_net_16073),
		.dout(new_net_16074)
	);

	bfr new_net_16075_bfr_after (
		.din(new_net_16074),
		.dout(new_net_16075)
	);

	bfr new_net_16076_bfr_after (
		.din(new_net_16075),
		.dout(new_net_16076)
	);

	bfr new_net_16077_bfr_after (
		.din(new_net_16076),
		.dout(new_net_16077)
	);

	bfr new_net_16078_bfr_after (
		.din(new_net_16077),
		.dout(new_net_16078)
	);

	bfr new_net_16079_bfr_after (
		.din(new_net_16078),
		.dout(new_net_16079)
	);

	bfr new_net_16080_bfr_after (
		.din(new_net_16079),
		.dout(new_net_16080)
	);

	spl2 _1564__v_fanout (
		.a(new_net_16080),
		.b(new_net_3119),
		.c(new_net_3120)
	);

	spl2 _1590__v_fanout (
		.a(_1590_),
		.b(new_net_1744),
		.c(new_net_1745)
	);

	bfr new_net_16081_bfr_after (
		.din(_1140_),
		.dout(new_net_16081)
	);

	bfr new_net_16082_bfr_after (
		.din(new_net_16081),
		.dout(new_net_16082)
	);

	bfr new_net_16083_bfr_after (
		.din(new_net_16082),
		.dout(new_net_16083)
	);

	bfr new_net_16084_bfr_after (
		.din(new_net_16083),
		.dout(new_net_16084)
	);

	bfr new_net_16085_bfr_after (
		.din(new_net_16084),
		.dout(new_net_16085)
	);

	bfr new_net_16086_bfr_after (
		.din(new_net_16085),
		.dout(new_net_16086)
	);

	bfr new_net_16087_bfr_after (
		.din(new_net_16086),
		.dout(new_net_16087)
	);

	bfr new_net_16088_bfr_after (
		.din(new_net_16087),
		.dout(new_net_16088)
	);

	bfr new_net_16089_bfr_after (
		.din(new_net_16088),
		.dout(new_net_16089)
	);

	bfr new_net_16090_bfr_after (
		.din(new_net_16089),
		.dout(new_net_16090)
	);

	bfr new_net_16091_bfr_after (
		.din(new_net_16090),
		.dout(new_net_16091)
	);

	bfr new_net_16092_bfr_after (
		.din(new_net_16091),
		.dout(new_net_16092)
	);

	bfr new_net_16093_bfr_after (
		.din(new_net_16092),
		.dout(new_net_16093)
	);

	bfr new_net_16094_bfr_after (
		.din(new_net_16093),
		.dout(new_net_16094)
	);

	bfr new_net_16095_bfr_after (
		.din(new_net_16094),
		.dout(new_net_16095)
	);

	bfr new_net_16096_bfr_after (
		.din(new_net_16095),
		.dout(new_net_16096)
	);

	spl2 _1140__v_fanout (
		.a(new_net_16096),
		.b(new_net_1275),
		.c(new_net_1276)
	);

	bfr new_net_16097_bfr_after (
		.din(_1294_),
		.dout(new_net_16097)
	);

	bfr new_net_16098_bfr_after (
		.din(new_net_16097),
		.dout(new_net_16098)
	);

	bfr new_net_16099_bfr_after (
		.din(new_net_16098),
		.dout(new_net_16099)
	);

	bfr new_net_16100_bfr_after (
		.din(new_net_16099),
		.dout(new_net_16100)
	);

	bfr new_net_16101_bfr_after (
		.din(new_net_16100),
		.dout(new_net_16101)
	);

	bfr new_net_16102_bfr_after (
		.din(new_net_16101),
		.dout(new_net_16102)
	);

	bfr new_net_16103_bfr_after (
		.din(new_net_16102),
		.dout(new_net_16103)
	);

	bfr new_net_16104_bfr_after (
		.din(new_net_16103),
		.dout(new_net_16104)
	);

	bfr new_net_16105_bfr_after (
		.din(new_net_16104),
		.dout(new_net_16105)
	);

	bfr new_net_16106_bfr_after (
		.din(new_net_16105),
		.dout(new_net_16106)
	);

	bfr new_net_16107_bfr_after (
		.din(new_net_16106),
		.dout(new_net_16107)
	);

	bfr new_net_16108_bfr_after (
		.din(new_net_16107),
		.dout(new_net_16108)
	);

	bfr new_net_16109_bfr_after (
		.din(new_net_16108),
		.dout(new_net_16109)
	);

	bfr new_net_16110_bfr_after (
		.din(new_net_16109),
		.dout(new_net_16110)
	);

	bfr new_net_16111_bfr_after (
		.din(new_net_16110),
		.dout(new_net_16111)
	);

	bfr new_net_16112_bfr_after (
		.din(new_net_16111),
		.dout(new_net_16112)
	);

	spl2 _1294__v_fanout (
		.a(new_net_16112),
		.b(new_net_3129),
		.c(new_net_3130)
	);

	bfr new_net_16113_bfr_after (
		.din(_0964_),
		.dout(new_net_16113)
	);

	bfr new_net_16114_bfr_after (
		.din(new_net_16113),
		.dout(new_net_16114)
	);

	bfr new_net_16115_bfr_after (
		.din(new_net_16114),
		.dout(new_net_16115)
	);

	bfr new_net_16116_bfr_after (
		.din(new_net_16115),
		.dout(new_net_16116)
	);

	bfr new_net_16117_bfr_after (
		.din(new_net_16116),
		.dout(new_net_16117)
	);

	bfr new_net_16118_bfr_after (
		.din(new_net_16117),
		.dout(new_net_16118)
	);

	bfr new_net_16119_bfr_after (
		.din(new_net_16118),
		.dout(new_net_16119)
	);

	bfr new_net_16120_bfr_after (
		.din(new_net_16119),
		.dout(new_net_16120)
	);

	bfr new_net_16121_bfr_after (
		.din(new_net_16120),
		.dout(new_net_16121)
	);

	bfr new_net_16122_bfr_after (
		.din(new_net_16121),
		.dout(new_net_16122)
	);

	bfr new_net_16123_bfr_after (
		.din(new_net_16122),
		.dout(new_net_16123)
	);

	bfr new_net_16124_bfr_after (
		.din(new_net_16123),
		.dout(new_net_16124)
	);

	bfr new_net_16125_bfr_after (
		.din(new_net_16124),
		.dout(new_net_16125)
	);

	bfr new_net_16126_bfr_after (
		.din(new_net_16125),
		.dout(new_net_16126)
	);

	bfr new_net_16127_bfr_after (
		.din(new_net_16126),
		.dout(new_net_16127)
	);

	bfr new_net_16128_bfr_after (
		.din(new_net_16127),
		.dout(new_net_16128)
	);

	bfr new_net_16129_bfr_after (
		.din(new_net_16128),
		.dout(new_net_16129)
	);

	bfr new_net_16130_bfr_after (
		.din(new_net_16129),
		.dout(new_net_16130)
	);

	bfr new_net_16131_bfr_after (
		.din(new_net_16130),
		.dout(new_net_16131)
	);

	bfr new_net_16132_bfr_after (
		.din(new_net_16131),
		.dout(new_net_16132)
	);

	bfr new_net_16133_bfr_after (
		.din(new_net_16132),
		.dout(new_net_16133)
	);

	bfr new_net_16134_bfr_after (
		.din(new_net_16133),
		.dout(new_net_16134)
	);

	bfr new_net_16135_bfr_after (
		.din(new_net_16134),
		.dout(new_net_16135)
	);

	bfr new_net_16136_bfr_after (
		.din(new_net_16135),
		.dout(new_net_16136)
	);

	bfr new_net_16137_bfr_after (
		.din(new_net_16136),
		.dout(new_net_16137)
	);

	bfr new_net_16138_bfr_after (
		.din(new_net_16137),
		.dout(new_net_16138)
	);

	bfr new_net_16139_bfr_after (
		.din(new_net_16138),
		.dout(new_net_16139)
	);

	bfr new_net_16140_bfr_after (
		.din(new_net_16139),
		.dout(new_net_16140)
	);

	bfr new_net_16141_bfr_after (
		.din(new_net_16140),
		.dout(new_net_16141)
	);

	bfr new_net_16142_bfr_after (
		.din(new_net_16141),
		.dout(new_net_16142)
	);

	bfr new_net_16143_bfr_after (
		.din(new_net_16142),
		.dout(new_net_16143)
	);

	bfr new_net_16144_bfr_after (
		.din(new_net_16143),
		.dout(new_net_16144)
	);

	bfr new_net_16145_bfr_after (
		.din(new_net_16144),
		.dout(new_net_16145)
	);

	bfr new_net_16146_bfr_after (
		.din(new_net_16145),
		.dout(new_net_16146)
	);

	bfr new_net_16147_bfr_after (
		.din(new_net_16146),
		.dout(new_net_16147)
	);

	bfr new_net_16148_bfr_after (
		.din(new_net_16147),
		.dout(new_net_16148)
	);

	bfr new_net_16149_bfr_after (
		.din(new_net_16148),
		.dout(new_net_16149)
	);

	bfr new_net_16150_bfr_after (
		.din(new_net_16149),
		.dout(new_net_16150)
	);

	bfr new_net_16151_bfr_after (
		.din(new_net_16150),
		.dout(new_net_16151)
	);

	bfr new_net_16152_bfr_after (
		.din(new_net_16151),
		.dout(new_net_16152)
	);

	bfr new_net_16153_bfr_after (
		.din(new_net_16152),
		.dout(new_net_16153)
	);

	bfr new_net_16154_bfr_after (
		.din(new_net_16153),
		.dout(new_net_16154)
	);

	bfr new_net_16155_bfr_after (
		.din(new_net_16154),
		.dout(new_net_16155)
	);

	bfr new_net_16156_bfr_after (
		.din(new_net_16155),
		.dout(new_net_16156)
	);

	bfr new_net_16157_bfr_after (
		.din(new_net_16156),
		.dout(new_net_16157)
	);

	bfr new_net_16158_bfr_after (
		.din(new_net_16157),
		.dout(new_net_16158)
	);

	bfr new_net_16159_bfr_after (
		.din(new_net_16158),
		.dout(new_net_16159)
	);

	bfr new_net_16160_bfr_after (
		.din(new_net_16159),
		.dout(new_net_16160)
	);

	bfr new_net_16161_bfr_after (
		.din(new_net_16160),
		.dout(new_net_16161)
	);

	bfr new_net_16162_bfr_after (
		.din(new_net_16161),
		.dout(new_net_16162)
	);

	bfr new_net_16163_bfr_after (
		.din(new_net_16162),
		.dout(new_net_16163)
	);

	bfr new_net_16164_bfr_after (
		.din(new_net_16163),
		.dout(new_net_16164)
	);

	bfr new_net_16165_bfr_after (
		.din(new_net_16164),
		.dout(new_net_16165)
	);

	bfr new_net_16166_bfr_after (
		.din(new_net_16165),
		.dout(new_net_16166)
	);

	bfr new_net_16167_bfr_after (
		.din(new_net_16166),
		.dout(new_net_16167)
	);

	bfr new_net_16168_bfr_after (
		.din(new_net_16167),
		.dout(new_net_16168)
	);

	bfr new_net_16169_bfr_after (
		.din(new_net_16168),
		.dout(new_net_16169)
	);

	bfr new_net_16170_bfr_after (
		.din(new_net_16169),
		.dout(new_net_16170)
	);

	bfr new_net_16171_bfr_after (
		.din(new_net_16170),
		.dout(new_net_16171)
	);

	bfr new_net_16172_bfr_after (
		.din(new_net_16171),
		.dout(new_net_16172)
	);

	bfr new_net_16173_bfr_after (
		.din(new_net_16172),
		.dout(new_net_16173)
	);

	bfr new_net_16174_bfr_after (
		.din(new_net_16173),
		.dout(new_net_16174)
	);

	bfr new_net_16175_bfr_after (
		.din(new_net_16174),
		.dout(new_net_16175)
	);

	bfr new_net_16176_bfr_after (
		.din(new_net_16175),
		.dout(new_net_16176)
	);

	bfr new_net_16177_bfr_after (
		.din(new_net_16176),
		.dout(new_net_16177)
	);

	bfr new_net_16178_bfr_after (
		.din(new_net_16177),
		.dout(new_net_16178)
	);

	bfr new_net_16179_bfr_after (
		.din(new_net_16178),
		.dout(new_net_16179)
	);

	bfr new_net_16180_bfr_after (
		.din(new_net_16179),
		.dout(new_net_16180)
	);

	bfr new_net_16181_bfr_after (
		.din(new_net_16180),
		.dout(new_net_16181)
	);

	bfr new_net_16182_bfr_after (
		.din(new_net_16181),
		.dout(new_net_16182)
	);

	bfr new_net_16183_bfr_after (
		.din(new_net_16182),
		.dout(new_net_16183)
	);

	bfr new_net_16184_bfr_after (
		.din(new_net_16183),
		.dout(new_net_16184)
	);

	bfr new_net_16185_bfr_after (
		.din(new_net_16184),
		.dout(new_net_16185)
	);

	bfr new_net_16186_bfr_after (
		.din(new_net_16185),
		.dout(new_net_16186)
	);

	bfr new_net_16187_bfr_after (
		.din(new_net_16186),
		.dout(new_net_16187)
	);

	bfr new_net_16188_bfr_after (
		.din(new_net_16187),
		.dout(new_net_16188)
	);

	bfr new_net_16189_bfr_after (
		.din(new_net_16188),
		.dout(new_net_16189)
	);

	bfr new_net_16190_bfr_after (
		.din(new_net_16189),
		.dout(new_net_16190)
	);

	bfr new_net_16191_bfr_after (
		.din(new_net_16190),
		.dout(new_net_16191)
	);

	bfr new_net_16192_bfr_after (
		.din(new_net_16191),
		.dout(new_net_16192)
	);

	bfr new_net_16193_bfr_after (
		.din(new_net_16192),
		.dout(new_net_16193)
	);

	bfr new_net_16194_bfr_after (
		.din(new_net_16193),
		.dout(new_net_16194)
	);

	bfr new_net_16195_bfr_after (
		.din(new_net_16194),
		.dout(new_net_16195)
	);

	bfr new_net_16196_bfr_after (
		.din(new_net_16195),
		.dout(new_net_16196)
	);

	bfr new_net_16197_bfr_after (
		.din(new_net_16196),
		.dout(new_net_16197)
	);

	bfr new_net_16198_bfr_after (
		.din(new_net_16197),
		.dout(new_net_16198)
	);

	bfr new_net_16199_bfr_after (
		.din(new_net_16198),
		.dout(new_net_16199)
	);

	bfr new_net_16200_bfr_after (
		.din(new_net_16199),
		.dout(new_net_16200)
	);

	bfr new_net_16201_bfr_after (
		.din(new_net_16200),
		.dout(new_net_16201)
	);

	bfr new_net_16202_bfr_after (
		.din(new_net_16201),
		.dout(new_net_16202)
	);

	bfr new_net_16203_bfr_after (
		.din(new_net_16202),
		.dout(new_net_16203)
	);

	bfr new_net_16204_bfr_after (
		.din(new_net_16203),
		.dout(new_net_16204)
	);

	bfr new_net_16205_bfr_after (
		.din(new_net_16204),
		.dout(new_net_16205)
	);

	bfr new_net_16206_bfr_after (
		.din(new_net_16205),
		.dout(new_net_16206)
	);

	spl2 _0964__v_fanout (
		.a(new_net_16206),
		.b(new_net_2585),
		.c(new_net_2586)
	);

	bfr new_net_16207_bfr_after (
		.din(_0961_),
		.dout(new_net_16207)
	);

	bfr new_net_16208_bfr_after (
		.din(new_net_16207),
		.dout(new_net_16208)
	);

	bfr new_net_16209_bfr_after (
		.din(new_net_16208),
		.dout(new_net_16209)
	);

	bfr new_net_16210_bfr_after (
		.din(new_net_16209),
		.dout(new_net_16210)
	);

	bfr new_net_16211_bfr_after (
		.din(new_net_16210),
		.dout(new_net_16211)
	);

	bfr new_net_16212_bfr_after (
		.din(new_net_16211),
		.dout(new_net_16212)
	);

	bfr new_net_16213_bfr_after (
		.din(new_net_16212),
		.dout(new_net_16213)
	);

	bfr new_net_16214_bfr_after (
		.din(new_net_16213),
		.dout(new_net_16214)
	);

	bfr new_net_16215_bfr_after (
		.din(new_net_16214),
		.dout(new_net_16215)
	);

	bfr new_net_16216_bfr_after (
		.din(new_net_16215),
		.dout(new_net_16216)
	);

	bfr new_net_16217_bfr_after (
		.din(new_net_16216),
		.dout(new_net_16217)
	);

	bfr new_net_16218_bfr_after (
		.din(new_net_16217),
		.dout(new_net_16218)
	);

	bfr new_net_16219_bfr_after (
		.din(new_net_16218),
		.dout(new_net_16219)
	);

	bfr new_net_16220_bfr_after (
		.din(new_net_16219),
		.dout(new_net_16220)
	);

	bfr new_net_16221_bfr_after (
		.din(new_net_16220),
		.dout(new_net_16221)
	);

	bfr new_net_16222_bfr_after (
		.din(new_net_16221),
		.dout(new_net_16222)
	);

	bfr new_net_16223_bfr_after (
		.din(new_net_16222),
		.dout(new_net_16223)
	);

	bfr new_net_16224_bfr_after (
		.din(new_net_16223),
		.dout(new_net_16224)
	);

	bfr new_net_16225_bfr_after (
		.din(new_net_16224),
		.dout(new_net_16225)
	);

	bfr new_net_16226_bfr_after (
		.din(new_net_16225),
		.dout(new_net_16226)
	);

	bfr new_net_16227_bfr_after (
		.din(new_net_16226),
		.dout(new_net_16227)
	);

	bfr new_net_16228_bfr_after (
		.din(new_net_16227),
		.dout(new_net_16228)
	);

	bfr new_net_16229_bfr_after (
		.din(new_net_16228),
		.dout(new_net_16229)
	);

	bfr new_net_16230_bfr_after (
		.din(new_net_16229),
		.dout(new_net_16230)
	);

	bfr new_net_16231_bfr_after (
		.din(new_net_16230),
		.dout(new_net_16231)
	);

	bfr new_net_16232_bfr_after (
		.din(new_net_16231),
		.dout(new_net_16232)
	);

	bfr new_net_16233_bfr_after (
		.din(new_net_16232),
		.dout(new_net_16233)
	);

	bfr new_net_16234_bfr_after (
		.din(new_net_16233),
		.dout(new_net_16234)
	);

	bfr new_net_16235_bfr_after (
		.din(new_net_16234),
		.dout(new_net_16235)
	);

	bfr new_net_16236_bfr_after (
		.din(new_net_16235),
		.dout(new_net_16236)
	);

	bfr new_net_16237_bfr_after (
		.din(new_net_16236),
		.dout(new_net_16237)
	);

	bfr new_net_16238_bfr_after (
		.din(new_net_16237),
		.dout(new_net_16238)
	);

	bfr new_net_16239_bfr_after (
		.din(new_net_16238),
		.dout(new_net_16239)
	);

	bfr new_net_16240_bfr_after (
		.din(new_net_16239),
		.dout(new_net_16240)
	);

	bfr new_net_16241_bfr_after (
		.din(new_net_16240),
		.dout(new_net_16241)
	);

	bfr new_net_16242_bfr_after (
		.din(new_net_16241),
		.dout(new_net_16242)
	);

	bfr new_net_16243_bfr_after (
		.din(new_net_16242),
		.dout(new_net_16243)
	);

	bfr new_net_16244_bfr_after (
		.din(new_net_16243),
		.dout(new_net_16244)
	);

	bfr new_net_16245_bfr_after (
		.din(new_net_16244),
		.dout(new_net_16245)
	);

	bfr new_net_16246_bfr_after (
		.din(new_net_16245),
		.dout(new_net_16246)
	);

	bfr new_net_16247_bfr_after (
		.din(new_net_16246),
		.dout(new_net_16247)
	);

	bfr new_net_16248_bfr_after (
		.din(new_net_16247),
		.dout(new_net_16248)
	);

	bfr new_net_16249_bfr_after (
		.din(new_net_16248),
		.dout(new_net_16249)
	);

	bfr new_net_16250_bfr_after (
		.din(new_net_16249),
		.dout(new_net_16250)
	);

	bfr new_net_16251_bfr_after (
		.din(new_net_16250),
		.dout(new_net_16251)
	);

	bfr new_net_16252_bfr_after (
		.din(new_net_16251),
		.dout(new_net_16252)
	);

	bfr new_net_16253_bfr_after (
		.din(new_net_16252),
		.dout(new_net_16253)
	);

	bfr new_net_16254_bfr_after (
		.din(new_net_16253),
		.dout(new_net_16254)
	);

	bfr new_net_16255_bfr_after (
		.din(new_net_16254),
		.dout(new_net_16255)
	);

	bfr new_net_16256_bfr_after (
		.din(new_net_16255),
		.dout(new_net_16256)
	);

	bfr new_net_16257_bfr_after (
		.din(new_net_16256),
		.dout(new_net_16257)
	);

	bfr new_net_16258_bfr_after (
		.din(new_net_16257),
		.dout(new_net_16258)
	);

	bfr new_net_16259_bfr_after (
		.din(new_net_16258),
		.dout(new_net_16259)
	);

	bfr new_net_16260_bfr_after (
		.din(new_net_16259),
		.dout(new_net_16260)
	);

	bfr new_net_16261_bfr_after (
		.din(new_net_16260),
		.dout(new_net_16261)
	);

	bfr new_net_16262_bfr_after (
		.din(new_net_16261),
		.dout(new_net_16262)
	);

	bfr new_net_16263_bfr_after (
		.din(new_net_16262),
		.dout(new_net_16263)
	);

	bfr new_net_16264_bfr_after (
		.din(new_net_16263),
		.dout(new_net_16264)
	);

	bfr new_net_16265_bfr_after (
		.din(new_net_16264),
		.dout(new_net_16265)
	);

	bfr new_net_16266_bfr_after (
		.din(new_net_16265),
		.dout(new_net_16266)
	);

	bfr new_net_16267_bfr_after (
		.din(new_net_16266),
		.dout(new_net_16267)
	);

	bfr new_net_16268_bfr_after (
		.din(new_net_16267),
		.dout(new_net_16268)
	);

	bfr new_net_16269_bfr_after (
		.din(new_net_16268),
		.dout(new_net_16269)
	);

	bfr new_net_16270_bfr_after (
		.din(new_net_16269),
		.dout(new_net_16270)
	);

	bfr new_net_16271_bfr_after (
		.din(new_net_16270),
		.dout(new_net_16271)
	);

	bfr new_net_16272_bfr_after (
		.din(new_net_16271),
		.dout(new_net_16272)
	);

	bfr new_net_16273_bfr_after (
		.din(new_net_16272),
		.dout(new_net_16273)
	);

	bfr new_net_16274_bfr_after (
		.din(new_net_16273),
		.dout(new_net_16274)
	);

	bfr new_net_16275_bfr_after (
		.din(new_net_16274),
		.dout(new_net_16275)
	);

	bfr new_net_16276_bfr_after (
		.din(new_net_16275),
		.dout(new_net_16276)
	);

	bfr new_net_16277_bfr_after (
		.din(new_net_16276),
		.dout(new_net_16277)
	);

	bfr new_net_16278_bfr_after (
		.din(new_net_16277),
		.dout(new_net_16278)
	);

	bfr new_net_16279_bfr_after (
		.din(new_net_16278),
		.dout(new_net_16279)
	);

	bfr new_net_16280_bfr_after (
		.din(new_net_16279),
		.dout(new_net_16280)
	);

	bfr new_net_16281_bfr_after (
		.din(new_net_16280),
		.dout(new_net_16281)
	);

	bfr new_net_16282_bfr_after (
		.din(new_net_16281),
		.dout(new_net_16282)
	);

	bfr new_net_16283_bfr_after (
		.din(new_net_16282),
		.dout(new_net_16283)
	);

	bfr new_net_16284_bfr_after (
		.din(new_net_16283),
		.dout(new_net_16284)
	);

	bfr new_net_16285_bfr_after (
		.din(new_net_16284),
		.dout(new_net_16285)
	);

	bfr new_net_16286_bfr_after (
		.din(new_net_16285),
		.dout(new_net_16286)
	);

	bfr new_net_16287_bfr_after (
		.din(new_net_16286),
		.dout(new_net_16287)
	);

	bfr new_net_16288_bfr_after (
		.din(new_net_16287),
		.dout(new_net_16288)
	);

	bfr new_net_16289_bfr_after (
		.din(new_net_16288),
		.dout(new_net_16289)
	);

	bfr new_net_16290_bfr_after (
		.din(new_net_16289),
		.dout(new_net_16290)
	);

	bfr new_net_16291_bfr_after (
		.din(new_net_16290),
		.dout(new_net_16291)
	);

	bfr new_net_16292_bfr_after (
		.din(new_net_16291),
		.dout(new_net_16292)
	);

	bfr new_net_16293_bfr_after (
		.din(new_net_16292),
		.dout(new_net_16293)
	);

	bfr new_net_16294_bfr_after (
		.din(new_net_16293),
		.dout(new_net_16294)
	);

	bfr new_net_16295_bfr_after (
		.din(new_net_16294),
		.dout(new_net_16295)
	);

	bfr new_net_16296_bfr_after (
		.din(new_net_16295),
		.dout(new_net_16296)
	);

	bfr new_net_16297_bfr_after (
		.din(new_net_16296),
		.dout(new_net_16297)
	);

	bfr new_net_16298_bfr_after (
		.din(new_net_16297),
		.dout(new_net_16298)
	);

	bfr new_net_16299_bfr_after (
		.din(new_net_16298),
		.dout(new_net_16299)
	);

	bfr new_net_16300_bfr_after (
		.din(new_net_16299),
		.dout(new_net_16300)
	);

	bfr new_net_16301_bfr_after (
		.din(new_net_16300),
		.dout(new_net_16301)
	);

	bfr new_net_16302_bfr_after (
		.din(new_net_16301),
		.dout(new_net_16302)
	);

	bfr new_net_16303_bfr_after (
		.din(new_net_16302),
		.dout(new_net_16303)
	);

	bfr new_net_16304_bfr_after (
		.din(new_net_16303),
		.dout(new_net_16304)
	);

	bfr new_net_16305_bfr_after (
		.din(new_net_16304),
		.dout(new_net_16305)
	);

	bfr new_net_16306_bfr_after (
		.din(new_net_16305),
		.dout(new_net_16306)
	);

	bfr new_net_16307_bfr_after (
		.din(new_net_16306),
		.dout(new_net_16307)
	);

	bfr new_net_16308_bfr_after (
		.din(new_net_16307),
		.dout(new_net_16308)
	);

	bfr new_net_16309_bfr_after (
		.din(new_net_16308),
		.dout(new_net_16309)
	);

	bfr new_net_16310_bfr_after (
		.din(new_net_16309),
		.dout(new_net_16310)
	);

	bfr new_net_16311_bfr_after (
		.din(new_net_16310),
		.dout(new_net_16311)
	);

	bfr new_net_16312_bfr_after (
		.din(new_net_16311),
		.dout(new_net_16312)
	);

	bfr new_net_16313_bfr_after (
		.din(new_net_16312),
		.dout(new_net_16313)
	);

	bfr new_net_16314_bfr_after (
		.din(new_net_16313),
		.dout(new_net_16314)
	);

	bfr new_net_16315_bfr_after (
		.din(new_net_16314),
		.dout(new_net_16315)
	);

	bfr new_net_16316_bfr_after (
		.din(new_net_16315),
		.dout(new_net_16316)
	);

	spl2 _0961__v_fanout (
		.a(new_net_16316),
		.b(new_net_2785),
		.c(new_net_2786)
	);

	bfr new_net_16317_bfr_after (
		.din(_0769_),
		.dout(new_net_16317)
	);

	bfr new_net_16318_bfr_after (
		.din(new_net_16317),
		.dout(new_net_16318)
	);

	bfr new_net_16319_bfr_after (
		.din(new_net_16318),
		.dout(new_net_16319)
	);

	bfr new_net_16320_bfr_after (
		.din(new_net_16319),
		.dout(new_net_16320)
	);

	bfr new_net_16321_bfr_after (
		.din(new_net_16320),
		.dout(new_net_16321)
	);

	bfr new_net_16322_bfr_after (
		.din(new_net_16321),
		.dout(new_net_16322)
	);

	bfr new_net_16323_bfr_after (
		.din(new_net_16322),
		.dout(new_net_16323)
	);

	bfr new_net_16324_bfr_after (
		.din(new_net_16323),
		.dout(new_net_16324)
	);

	bfr new_net_16325_bfr_after (
		.din(new_net_16324),
		.dout(new_net_16325)
	);

	bfr new_net_16326_bfr_after (
		.din(new_net_16325),
		.dout(new_net_16326)
	);

	bfr new_net_16327_bfr_after (
		.din(new_net_16326),
		.dout(new_net_16327)
	);

	bfr new_net_16328_bfr_after (
		.din(new_net_16327),
		.dout(new_net_16328)
	);

	bfr new_net_16329_bfr_after (
		.din(new_net_16328),
		.dout(new_net_16329)
	);

	bfr new_net_16330_bfr_after (
		.din(new_net_16329),
		.dout(new_net_16330)
	);

	bfr new_net_16331_bfr_after (
		.din(new_net_16330),
		.dout(new_net_16331)
	);

	bfr new_net_16332_bfr_after (
		.din(new_net_16331),
		.dout(new_net_16332)
	);

	bfr new_net_16333_bfr_after (
		.din(new_net_16332),
		.dout(new_net_16333)
	);

	bfr new_net_16334_bfr_after (
		.din(new_net_16333),
		.dout(new_net_16334)
	);

	bfr new_net_16335_bfr_after (
		.din(new_net_16334),
		.dout(new_net_16335)
	);

	bfr new_net_16336_bfr_after (
		.din(new_net_16335),
		.dout(new_net_16336)
	);

	bfr new_net_16337_bfr_after (
		.din(new_net_16336),
		.dout(new_net_16337)
	);

	bfr new_net_16338_bfr_after (
		.din(new_net_16337),
		.dout(new_net_16338)
	);

	bfr new_net_16339_bfr_after (
		.din(new_net_16338),
		.dout(new_net_16339)
	);

	bfr new_net_16340_bfr_after (
		.din(new_net_16339),
		.dout(new_net_16340)
	);

	bfr new_net_16341_bfr_after (
		.din(new_net_16340),
		.dout(new_net_16341)
	);

	bfr new_net_16342_bfr_after (
		.din(new_net_16341),
		.dout(new_net_16342)
	);

	bfr new_net_16343_bfr_after (
		.din(new_net_16342),
		.dout(new_net_16343)
	);

	bfr new_net_16344_bfr_after (
		.din(new_net_16343),
		.dout(new_net_16344)
	);

	bfr new_net_16345_bfr_after (
		.din(new_net_16344),
		.dout(new_net_16345)
	);

	bfr new_net_16346_bfr_after (
		.din(new_net_16345),
		.dout(new_net_16346)
	);

	bfr new_net_16347_bfr_after (
		.din(new_net_16346),
		.dout(new_net_16347)
	);

	bfr new_net_16348_bfr_after (
		.din(new_net_16347),
		.dout(new_net_16348)
	);

	bfr new_net_16349_bfr_after (
		.din(new_net_16348),
		.dout(new_net_16349)
	);

	bfr new_net_16350_bfr_after (
		.din(new_net_16349),
		.dout(new_net_16350)
	);

	bfr new_net_16351_bfr_after (
		.din(new_net_16350),
		.dout(new_net_16351)
	);

	bfr new_net_16352_bfr_after (
		.din(new_net_16351),
		.dout(new_net_16352)
	);

	bfr new_net_16353_bfr_after (
		.din(new_net_16352),
		.dout(new_net_16353)
	);

	bfr new_net_16354_bfr_after (
		.din(new_net_16353),
		.dout(new_net_16354)
	);

	bfr new_net_16355_bfr_after (
		.din(new_net_16354),
		.dout(new_net_16355)
	);

	bfr new_net_16356_bfr_after (
		.din(new_net_16355),
		.dout(new_net_16356)
	);

	bfr new_net_16357_bfr_after (
		.din(new_net_16356),
		.dout(new_net_16357)
	);

	bfr new_net_16358_bfr_after (
		.din(new_net_16357),
		.dout(new_net_16358)
	);

	bfr new_net_16359_bfr_after (
		.din(new_net_16358),
		.dout(new_net_16359)
	);

	bfr new_net_16360_bfr_after (
		.din(new_net_16359),
		.dout(new_net_16360)
	);

	bfr new_net_16361_bfr_after (
		.din(new_net_16360),
		.dout(new_net_16361)
	);

	bfr new_net_16362_bfr_after (
		.din(new_net_16361),
		.dout(new_net_16362)
	);

	bfr new_net_16363_bfr_after (
		.din(new_net_16362),
		.dout(new_net_16363)
	);

	bfr new_net_16364_bfr_after (
		.din(new_net_16363),
		.dout(new_net_16364)
	);

	bfr new_net_16365_bfr_after (
		.din(new_net_16364),
		.dout(new_net_16365)
	);

	bfr new_net_16366_bfr_after (
		.din(new_net_16365),
		.dout(new_net_16366)
	);

	bfr new_net_16367_bfr_after (
		.din(new_net_16366),
		.dout(new_net_16367)
	);

	bfr new_net_16368_bfr_after (
		.din(new_net_16367),
		.dout(new_net_16368)
	);

	bfr new_net_16369_bfr_after (
		.din(new_net_16368),
		.dout(new_net_16369)
	);

	bfr new_net_16370_bfr_after (
		.din(new_net_16369),
		.dout(new_net_16370)
	);

	bfr new_net_16371_bfr_after (
		.din(new_net_16370),
		.dout(new_net_16371)
	);

	bfr new_net_16372_bfr_after (
		.din(new_net_16371),
		.dout(new_net_16372)
	);

	bfr new_net_16373_bfr_after (
		.din(new_net_16372),
		.dout(new_net_16373)
	);

	bfr new_net_16374_bfr_after (
		.din(new_net_16373),
		.dout(new_net_16374)
	);

	bfr new_net_16375_bfr_after (
		.din(new_net_16374),
		.dout(new_net_16375)
	);

	bfr new_net_16376_bfr_after (
		.din(new_net_16375),
		.dout(new_net_16376)
	);

	bfr new_net_16377_bfr_after (
		.din(new_net_16376),
		.dout(new_net_16377)
	);

	bfr new_net_16378_bfr_after (
		.din(new_net_16377),
		.dout(new_net_16378)
	);

	bfr new_net_16379_bfr_after (
		.din(new_net_16378),
		.dout(new_net_16379)
	);

	bfr new_net_16380_bfr_after (
		.din(new_net_16379),
		.dout(new_net_16380)
	);

	bfr new_net_16381_bfr_after (
		.din(new_net_16380),
		.dout(new_net_16381)
	);

	bfr new_net_16382_bfr_after (
		.din(new_net_16381),
		.dout(new_net_16382)
	);

	bfr new_net_16383_bfr_after (
		.din(new_net_16382),
		.dout(new_net_16383)
	);

	bfr new_net_16384_bfr_after (
		.din(new_net_16383),
		.dout(new_net_16384)
	);

	bfr new_net_16385_bfr_after (
		.din(new_net_16384),
		.dout(new_net_16385)
	);

	bfr new_net_16386_bfr_after (
		.din(new_net_16385),
		.dout(new_net_16386)
	);

	bfr new_net_16387_bfr_after (
		.din(new_net_16386),
		.dout(new_net_16387)
	);

	bfr new_net_16388_bfr_after (
		.din(new_net_16387),
		.dout(new_net_16388)
	);

	bfr new_net_16389_bfr_after (
		.din(new_net_16388),
		.dout(new_net_16389)
	);

	bfr new_net_16390_bfr_after (
		.din(new_net_16389),
		.dout(new_net_16390)
	);

	bfr new_net_16391_bfr_after (
		.din(new_net_16390),
		.dout(new_net_16391)
	);

	bfr new_net_16392_bfr_after (
		.din(new_net_16391),
		.dout(new_net_16392)
	);

	bfr new_net_16393_bfr_after (
		.din(new_net_16392),
		.dout(new_net_16393)
	);

	bfr new_net_16394_bfr_after (
		.din(new_net_16393),
		.dout(new_net_16394)
	);

	bfr new_net_16395_bfr_after (
		.din(new_net_16394),
		.dout(new_net_16395)
	);

	bfr new_net_16396_bfr_after (
		.din(new_net_16395),
		.dout(new_net_16396)
	);

	bfr new_net_16397_bfr_after (
		.din(new_net_16396),
		.dout(new_net_16397)
	);

	bfr new_net_16398_bfr_after (
		.din(new_net_16397),
		.dout(new_net_16398)
	);

	bfr new_net_16399_bfr_after (
		.din(new_net_16398),
		.dout(new_net_16399)
	);

	bfr new_net_16400_bfr_after (
		.din(new_net_16399),
		.dout(new_net_16400)
	);

	bfr new_net_16401_bfr_after (
		.din(new_net_16400),
		.dout(new_net_16401)
	);

	bfr new_net_16402_bfr_after (
		.din(new_net_16401),
		.dout(new_net_16402)
	);

	bfr new_net_16403_bfr_after (
		.din(new_net_16402),
		.dout(new_net_16403)
	);

	bfr new_net_16404_bfr_after (
		.din(new_net_16403),
		.dout(new_net_16404)
	);

	bfr new_net_16405_bfr_after (
		.din(new_net_16404),
		.dout(new_net_16405)
	);

	bfr new_net_16406_bfr_after (
		.din(new_net_16405),
		.dout(new_net_16406)
	);

	bfr new_net_16407_bfr_after (
		.din(new_net_16406),
		.dout(new_net_16407)
	);

	bfr new_net_16408_bfr_after (
		.din(new_net_16407),
		.dout(new_net_16408)
	);

	bfr new_net_16409_bfr_after (
		.din(new_net_16408),
		.dout(new_net_16409)
	);

	bfr new_net_16410_bfr_after (
		.din(new_net_16409),
		.dout(new_net_16410)
	);

	bfr new_net_16411_bfr_after (
		.din(new_net_16410),
		.dout(new_net_16411)
	);

	bfr new_net_16412_bfr_after (
		.din(new_net_16411),
		.dout(new_net_16412)
	);

	bfr new_net_16413_bfr_after (
		.din(new_net_16412),
		.dout(new_net_16413)
	);

	bfr new_net_16414_bfr_after (
		.din(new_net_16413),
		.dout(new_net_16414)
	);

	bfr new_net_16415_bfr_after (
		.din(new_net_16414),
		.dout(new_net_16415)
	);

	bfr new_net_16416_bfr_after (
		.din(new_net_16415),
		.dout(new_net_16416)
	);

	bfr new_net_16417_bfr_after (
		.din(new_net_16416),
		.dout(new_net_16417)
	);

	bfr new_net_16418_bfr_after (
		.din(new_net_16417),
		.dout(new_net_16418)
	);

	bfr new_net_16419_bfr_after (
		.din(new_net_16418),
		.dout(new_net_16419)
	);

	bfr new_net_16420_bfr_after (
		.din(new_net_16419),
		.dout(new_net_16420)
	);

	spl2 _0769__v_fanout (
		.a(new_net_16420),
		.b(new_net_1096),
		.c(new_net_1097)
	);

	bfr new_net_16421_bfr_after (
		.din(_0888_),
		.dout(new_net_16421)
	);

	bfr new_net_16422_bfr_after (
		.din(new_net_16421),
		.dout(new_net_16422)
	);

	bfr new_net_16423_bfr_after (
		.din(new_net_16422),
		.dout(new_net_16423)
	);

	bfr new_net_16424_bfr_after (
		.din(new_net_16423),
		.dout(new_net_16424)
	);

	bfr new_net_16425_bfr_after (
		.din(new_net_16424),
		.dout(new_net_16425)
	);

	bfr new_net_16426_bfr_after (
		.din(new_net_16425),
		.dout(new_net_16426)
	);

	bfr new_net_16427_bfr_after (
		.din(new_net_16426),
		.dout(new_net_16427)
	);

	bfr new_net_16428_bfr_after (
		.din(new_net_16427),
		.dout(new_net_16428)
	);

	bfr new_net_16429_bfr_after (
		.din(new_net_16428),
		.dout(new_net_16429)
	);

	bfr new_net_16430_bfr_after (
		.din(new_net_16429),
		.dout(new_net_16430)
	);

	bfr new_net_16431_bfr_after (
		.din(new_net_16430),
		.dout(new_net_16431)
	);

	bfr new_net_16432_bfr_after (
		.din(new_net_16431),
		.dout(new_net_16432)
	);

	bfr new_net_16433_bfr_after (
		.din(new_net_16432),
		.dout(new_net_16433)
	);

	bfr new_net_16434_bfr_after (
		.din(new_net_16433),
		.dout(new_net_16434)
	);

	bfr new_net_16435_bfr_after (
		.din(new_net_16434),
		.dout(new_net_16435)
	);

	bfr new_net_16436_bfr_after (
		.din(new_net_16435),
		.dout(new_net_16436)
	);

	bfr new_net_16437_bfr_after (
		.din(new_net_16436),
		.dout(new_net_16437)
	);

	bfr new_net_16438_bfr_after (
		.din(new_net_16437),
		.dout(new_net_16438)
	);

	bfr new_net_16439_bfr_after (
		.din(new_net_16438),
		.dout(new_net_16439)
	);

	bfr new_net_16440_bfr_after (
		.din(new_net_16439),
		.dout(new_net_16440)
	);

	bfr new_net_16441_bfr_after (
		.din(new_net_16440),
		.dout(new_net_16441)
	);

	bfr new_net_16442_bfr_after (
		.din(new_net_16441),
		.dout(new_net_16442)
	);

	bfr new_net_16443_bfr_after (
		.din(new_net_16442),
		.dout(new_net_16443)
	);

	bfr new_net_16444_bfr_after (
		.din(new_net_16443),
		.dout(new_net_16444)
	);

	bfr new_net_16445_bfr_after (
		.din(new_net_16444),
		.dout(new_net_16445)
	);

	bfr new_net_16446_bfr_after (
		.din(new_net_16445),
		.dout(new_net_16446)
	);

	bfr new_net_16447_bfr_after (
		.din(new_net_16446),
		.dout(new_net_16447)
	);

	bfr new_net_16448_bfr_after (
		.din(new_net_16447),
		.dout(new_net_16448)
	);

	bfr new_net_16449_bfr_after (
		.din(new_net_16448),
		.dout(new_net_16449)
	);

	bfr new_net_16450_bfr_after (
		.din(new_net_16449),
		.dout(new_net_16450)
	);

	bfr new_net_16451_bfr_after (
		.din(new_net_16450),
		.dout(new_net_16451)
	);

	bfr new_net_16452_bfr_after (
		.din(new_net_16451),
		.dout(new_net_16452)
	);

	bfr new_net_16453_bfr_after (
		.din(new_net_16452),
		.dout(new_net_16453)
	);

	bfr new_net_16454_bfr_after (
		.din(new_net_16453),
		.dout(new_net_16454)
	);

	bfr new_net_16455_bfr_after (
		.din(new_net_16454),
		.dout(new_net_16455)
	);

	bfr new_net_16456_bfr_after (
		.din(new_net_16455),
		.dout(new_net_16456)
	);

	bfr new_net_16457_bfr_after (
		.din(new_net_16456),
		.dout(new_net_16457)
	);

	bfr new_net_16458_bfr_after (
		.din(new_net_16457),
		.dout(new_net_16458)
	);

	bfr new_net_16459_bfr_after (
		.din(new_net_16458),
		.dout(new_net_16459)
	);

	bfr new_net_16460_bfr_after (
		.din(new_net_16459),
		.dout(new_net_16460)
	);

	bfr new_net_16461_bfr_after (
		.din(new_net_16460),
		.dout(new_net_16461)
	);

	bfr new_net_16462_bfr_after (
		.din(new_net_16461),
		.dout(new_net_16462)
	);

	bfr new_net_16463_bfr_after (
		.din(new_net_16462),
		.dout(new_net_16463)
	);

	bfr new_net_16464_bfr_after (
		.din(new_net_16463),
		.dout(new_net_16464)
	);

	bfr new_net_16465_bfr_after (
		.din(new_net_16464),
		.dout(new_net_16465)
	);

	bfr new_net_16466_bfr_after (
		.din(new_net_16465),
		.dout(new_net_16466)
	);

	bfr new_net_16467_bfr_after (
		.din(new_net_16466),
		.dout(new_net_16467)
	);

	bfr new_net_16468_bfr_after (
		.din(new_net_16467),
		.dout(new_net_16468)
	);

	bfr new_net_16469_bfr_after (
		.din(new_net_16468),
		.dout(new_net_16469)
	);

	bfr new_net_16470_bfr_after (
		.din(new_net_16469),
		.dout(new_net_16470)
	);

	bfr new_net_16471_bfr_after (
		.din(new_net_16470),
		.dout(new_net_16471)
	);

	bfr new_net_16472_bfr_after (
		.din(new_net_16471),
		.dout(new_net_16472)
	);

	bfr new_net_16473_bfr_after (
		.din(new_net_16472),
		.dout(new_net_16473)
	);

	bfr new_net_16474_bfr_after (
		.din(new_net_16473),
		.dout(new_net_16474)
	);

	bfr new_net_16475_bfr_after (
		.din(new_net_16474),
		.dout(new_net_16475)
	);

	bfr new_net_16476_bfr_after (
		.din(new_net_16475),
		.dout(new_net_16476)
	);

	bfr new_net_16477_bfr_after (
		.din(new_net_16476),
		.dout(new_net_16477)
	);

	bfr new_net_16478_bfr_after (
		.din(new_net_16477),
		.dout(new_net_16478)
	);

	bfr new_net_16479_bfr_after (
		.din(new_net_16478),
		.dout(new_net_16479)
	);

	bfr new_net_16480_bfr_after (
		.din(new_net_16479),
		.dout(new_net_16480)
	);

	bfr new_net_16481_bfr_after (
		.din(new_net_16480),
		.dout(new_net_16481)
	);

	bfr new_net_16482_bfr_after (
		.din(new_net_16481),
		.dout(new_net_16482)
	);

	bfr new_net_16483_bfr_after (
		.din(new_net_16482),
		.dout(new_net_16483)
	);

	bfr new_net_16484_bfr_after (
		.din(new_net_16483),
		.dout(new_net_16484)
	);

	bfr new_net_16485_bfr_after (
		.din(new_net_16484),
		.dout(new_net_16485)
	);

	bfr new_net_16486_bfr_after (
		.din(new_net_16485),
		.dout(new_net_16486)
	);

	bfr new_net_16487_bfr_after (
		.din(new_net_16486),
		.dout(new_net_16487)
	);

	bfr new_net_16488_bfr_after (
		.din(new_net_16487),
		.dout(new_net_16488)
	);

	bfr new_net_16489_bfr_after (
		.din(new_net_16488),
		.dout(new_net_16489)
	);

	bfr new_net_16490_bfr_after (
		.din(new_net_16489),
		.dout(new_net_16490)
	);

	bfr new_net_16491_bfr_after (
		.din(new_net_16490),
		.dout(new_net_16491)
	);

	bfr new_net_16492_bfr_after (
		.din(new_net_16491),
		.dout(new_net_16492)
	);

	bfr new_net_16493_bfr_after (
		.din(new_net_16492),
		.dout(new_net_16493)
	);

	bfr new_net_16494_bfr_after (
		.din(new_net_16493),
		.dout(new_net_16494)
	);

	bfr new_net_16495_bfr_after (
		.din(new_net_16494),
		.dout(new_net_16495)
	);

	bfr new_net_16496_bfr_after (
		.din(new_net_16495),
		.dout(new_net_16496)
	);

	bfr new_net_16497_bfr_after (
		.din(new_net_16496),
		.dout(new_net_16497)
	);

	bfr new_net_16498_bfr_after (
		.din(new_net_16497),
		.dout(new_net_16498)
	);

	bfr new_net_16499_bfr_after (
		.din(new_net_16498),
		.dout(new_net_16499)
	);

	bfr new_net_16500_bfr_after (
		.din(new_net_16499),
		.dout(new_net_16500)
	);

	bfr new_net_16501_bfr_after (
		.din(new_net_16500),
		.dout(new_net_16501)
	);

	bfr new_net_16502_bfr_after (
		.din(new_net_16501),
		.dout(new_net_16502)
	);

	spl2 _0888__v_fanout (
		.a(new_net_16502),
		.b(new_net_1582),
		.c(new_net_1583)
	);

	bfr new_net_16503_bfr_after (
		.din(_0623_),
		.dout(new_net_16503)
	);

	bfr new_net_16504_bfr_after (
		.din(new_net_16503),
		.dout(new_net_16504)
	);

	bfr new_net_16505_bfr_after (
		.din(new_net_16504),
		.dout(new_net_16505)
	);

	bfr new_net_16506_bfr_after (
		.din(new_net_16505),
		.dout(new_net_16506)
	);

	bfr new_net_16507_bfr_after (
		.din(new_net_16506),
		.dout(new_net_16507)
	);

	bfr new_net_16508_bfr_after (
		.din(new_net_16507),
		.dout(new_net_16508)
	);

	bfr new_net_16509_bfr_after (
		.din(new_net_16508),
		.dout(new_net_16509)
	);

	bfr new_net_16510_bfr_after (
		.din(new_net_16509),
		.dout(new_net_16510)
	);

	bfr new_net_16511_bfr_after (
		.din(new_net_16510),
		.dout(new_net_16511)
	);

	bfr new_net_16512_bfr_after (
		.din(new_net_16511),
		.dout(new_net_16512)
	);

	bfr new_net_16513_bfr_after (
		.din(new_net_16512),
		.dout(new_net_16513)
	);

	bfr new_net_16514_bfr_after (
		.din(new_net_16513),
		.dout(new_net_16514)
	);

	bfr new_net_16515_bfr_after (
		.din(new_net_16514),
		.dout(new_net_16515)
	);

	bfr new_net_16516_bfr_after (
		.din(new_net_16515),
		.dout(new_net_16516)
	);

	bfr new_net_16517_bfr_after (
		.din(new_net_16516),
		.dout(new_net_16517)
	);

	bfr new_net_16518_bfr_after (
		.din(new_net_16517),
		.dout(new_net_16518)
	);

	bfr new_net_16519_bfr_after (
		.din(new_net_16518),
		.dout(new_net_16519)
	);

	bfr new_net_16520_bfr_after (
		.din(new_net_16519),
		.dout(new_net_16520)
	);

	bfr new_net_16521_bfr_after (
		.din(new_net_16520),
		.dout(new_net_16521)
	);

	bfr new_net_16522_bfr_after (
		.din(new_net_16521),
		.dout(new_net_16522)
	);

	bfr new_net_16523_bfr_after (
		.din(new_net_16522),
		.dout(new_net_16523)
	);

	bfr new_net_16524_bfr_after (
		.din(new_net_16523),
		.dout(new_net_16524)
	);

	bfr new_net_16525_bfr_after (
		.din(new_net_16524),
		.dout(new_net_16525)
	);

	bfr new_net_16526_bfr_after (
		.din(new_net_16525),
		.dout(new_net_16526)
	);

	bfr new_net_16527_bfr_after (
		.din(new_net_16526),
		.dout(new_net_16527)
	);

	bfr new_net_16528_bfr_after (
		.din(new_net_16527),
		.dout(new_net_16528)
	);

	bfr new_net_16529_bfr_after (
		.din(new_net_16528),
		.dout(new_net_16529)
	);

	bfr new_net_16530_bfr_after (
		.din(new_net_16529),
		.dout(new_net_16530)
	);

	bfr new_net_16531_bfr_after (
		.din(new_net_16530),
		.dout(new_net_16531)
	);

	bfr new_net_16532_bfr_after (
		.din(new_net_16531),
		.dout(new_net_16532)
	);

	bfr new_net_16533_bfr_after (
		.din(new_net_16532),
		.dout(new_net_16533)
	);

	bfr new_net_16534_bfr_after (
		.din(new_net_16533),
		.dout(new_net_16534)
	);

	bfr new_net_16535_bfr_after (
		.din(new_net_16534),
		.dout(new_net_16535)
	);

	bfr new_net_16536_bfr_after (
		.din(new_net_16535),
		.dout(new_net_16536)
	);

	bfr new_net_16537_bfr_after (
		.din(new_net_16536),
		.dout(new_net_16537)
	);

	bfr new_net_16538_bfr_after (
		.din(new_net_16537),
		.dout(new_net_16538)
	);

	bfr new_net_16539_bfr_after (
		.din(new_net_16538),
		.dout(new_net_16539)
	);

	bfr new_net_16540_bfr_after (
		.din(new_net_16539),
		.dout(new_net_16540)
	);

	bfr new_net_16541_bfr_after (
		.din(new_net_16540),
		.dout(new_net_16541)
	);

	bfr new_net_16542_bfr_after (
		.din(new_net_16541),
		.dout(new_net_16542)
	);

	bfr new_net_16543_bfr_after (
		.din(new_net_16542),
		.dout(new_net_16543)
	);

	bfr new_net_16544_bfr_after (
		.din(new_net_16543),
		.dout(new_net_16544)
	);

	bfr new_net_16545_bfr_after (
		.din(new_net_16544),
		.dout(new_net_16545)
	);

	bfr new_net_16546_bfr_after (
		.din(new_net_16545),
		.dout(new_net_16546)
	);

	bfr new_net_16547_bfr_after (
		.din(new_net_16546),
		.dout(new_net_16547)
	);

	bfr new_net_16548_bfr_after (
		.din(new_net_16547),
		.dout(new_net_16548)
	);

	bfr new_net_16549_bfr_after (
		.din(new_net_16548),
		.dout(new_net_16549)
	);

	bfr new_net_16550_bfr_after (
		.din(new_net_16549),
		.dout(new_net_16550)
	);

	bfr new_net_16551_bfr_after (
		.din(new_net_16550),
		.dout(new_net_16551)
	);

	bfr new_net_16552_bfr_after (
		.din(new_net_16551),
		.dout(new_net_16552)
	);

	bfr new_net_16553_bfr_after (
		.din(new_net_16552),
		.dout(new_net_16553)
	);

	bfr new_net_16554_bfr_after (
		.din(new_net_16553),
		.dout(new_net_16554)
	);

	bfr new_net_16555_bfr_after (
		.din(new_net_16554),
		.dout(new_net_16555)
	);

	bfr new_net_16556_bfr_after (
		.din(new_net_16555),
		.dout(new_net_16556)
	);

	bfr new_net_16557_bfr_after (
		.din(new_net_16556),
		.dout(new_net_16557)
	);

	bfr new_net_16558_bfr_after (
		.din(new_net_16557),
		.dout(new_net_16558)
	);

	bfr new_net_16559_bfr_after (
		.din(new_net_16558),
		.dout(new_net_16559)
	);

	bfr new_net_16560_bfr_after (
		.din(new_net_16559),
		.dout(new_net_16560)
	);

	bfr new_net_16561_bfr_after (
		.din(new_net_16560),
		.dout(new_net_16561)
	);

	bfr new_net_16562_bfr_after (
		.din(new_net_16561),
		.dout(new_net_16562)
	);

	bfr new_net_16563_bfr_after (
		.din(new_net_16562),
		.dout(new_net_16563)
	);

	bfr new_net_16564_bfr_after (
		.din(new_net_16563),
		.dout(new_net_16564)
	);

	bfr new_net_16565_bfr_after (
		.din(new_net_16564),
		.dout(new_net_16565)
	);

	bfr new_net_16566_bfr_after (
		.din(new_net_16565),
		.dout(new_net_16566)
	);

	bfr new_net_16567_bfr_after (
		.din(new_net_16566),
		.dout(new_net_16567)
	);

	bfr new_net_16568_bfr_after (
		.din(new_net_16567),
		.dout(new_net_16568)
	);

	bfr new_net_16569_bfr_after (
		.din(new_net_16568),
		.dout(new_net_16569)
	);

	bfr new_net_16570_bfr_after (
		.din(new_net_16569),
		.dout(new_net_16570)
	);

	bfr new_net_16571_bfr_after (
		.din(new_net_16570),
		.dout(new_net_16571)
	);

	bfr new_net_16572_bfr_after (
		.din(new_net_16571),
		.dout(new_net_16572)
	);

	bfr new_net_16573_bfr_after (
		.din(new_net_16572),
		.dout(new_net_16573)
	);

	bfr new_net_16574_bfr_after (
		.din(new_net_16573),
		.dout(new_net_16574)
	);

	bfr new_net_16575_bfr_after (
		.din(new_net_16574),
		.dout(new_net_16575)
	);

	bfr new_net_16576_bfr_after (
		.din(new_net_16575),
		.dout(new_net_16576)
	);

	bfr new_net_16577_bfr_after (
		.din(new_net_16576),
		.dout(new_net_16577)
	);

	bfr new_net_16578_bfr_after (
		.din(new_net_16577),
		.dout(new_net_16578)
	);

	bfr new_net_16579_bfr_after (
		.din(new_net_16578),
		.dout(new_net_16579)
	);

	bfr new_net_16580_bfr_after (
		.din(new_net_16579),
		.dout(new_net_16580)
	);

	bfr new_net_16581_bfr_after (
		.din(new_net_16580),
		.dout(new_net_16581)
	);

	bfr new_net_16582_bfr_after (
		.din(new_net_16581),
		.dout(new_net_16582)
	);

	bfr new_net_16583_bfr_after (
		.din(new_net_16582),
		.dout(new_net_16583)
	);

	bfr new_net_16584_bfr_after (
		.din(new_net_16583),
		.dout(new_net_16584)
	);

	bfr new_net_16585_bfr_after (
		.din(new_net_16584),
		.dout(new_net_16585)
	);

	bfr new_net_16586_bfr_after (
		.din(new_net_16585),
		.dout(new_net_16586)
	);

	bfr new_net_16587_bfr_after (
		.din(new_net_16586),
		.dout(new_net_16587)
	);

	bfr new_net_16588_bfr_after (
		.din(new_net_16587),
		.dout(new_net_16588)
	);

	bfr new_net_16589_bfr_after (
		.din(new_net_16588),
		.dout(new_net_16589)
	);

	bfr new_net_16590_bfr_after (
		.din(new_net_16589),
		.dout(new_net_16590)
	);

	spl2 _0623__v_fanout (
		.a(new_net_16590),
		.b(new_net_246),
		.c(new_net_247)
	);

	bfr new_net_16591_bfr_after (
		.din(_0548_),
		.dout(new_net_16591)
	);

	bfr new_net_16592_bfr_after (
		.din(new_net_16591),
		.dout(new_net_16592)
	);

	bfr new_net_16593_bfr_after (
		.din(new_net_16592),
		.dout(new_net_16593)
	);

	bfr new_net_16594_bfr_after (
		.din(new_net_16593),
		.dout(new_net_16594)
	);

	bfr new_net_16595_bfr_after (
		.din(new_net_16594),
		.dout(new_net_16595)
	);

	bfr new_net_16596_bfr_after (
		.din(new_net_16595),
		.dout(new_net_16596)
	);

	bfr new_net_16597_bfr_after (
		.din(new_net_16596),
		.dout(new_net_16597)
	);

	bfr new_net_16598_bfr_after (
		.din(new_net_16597),
		.dout(new_net_16598)
	);

	bfr new_net_16599_bfr_after (
		.din(new_net_16598),
		.dout(new_net_16599)
	);

	bfr new_net_16600_bfr_after (
		.din(new_net_16599),
		.dout(new_net_16600)
	);

	bfr new_net_16601_bfr_after (
		.din(new_net_16600),
		.dout(new_net_16601)
	);

	bfr new_net_16602_bfr_after (
		.din(new_net_16601),
		.dout(new_net_16602)
	);

	bfr new_net_16603_bfr_after (
		.din(new_net_16602),
		.dout(new_net_16603)
	);

	bfr new_net_16604_bfr_after (
		.din(new_net_16603),
		.dout(new_net_16604)
	);

	bfr new_net_16605_bfr_after (
		.din(new_net_16604),
		.dout(new_net_16605)
	);

	bfr new_net_16606_bfr_after (
		.din(new_net_16605),
		.dout(new_net_16606)
	);

	bfr new_net_16607_bfr_after (
		.din(new_net_16606),
		.dout(new_net_16607)
	);

	bfr new_net_16608_bfr_after (
		.din(new_net_16607),
		.dout(new_net_16608)
	);

	bfr new_net_16609_bfr_after (
		.din(new_net_16608),
		.dout(new_net_16609)
	);

	bfr new_net_16610_bfr_after (
		.din(new_net_16609),
		.dout(new_net_16610)
	);

	bfr new_net_16611_bfr_after (
		.din(new_net_16610),
		.dout(new_net_16611)
	);

	bfr new_net_16612_bfr_after (
		.din(new_net_16611),
		.dout(new_net_16612)
	);

	bfr new_net_16613_bfr_after (
		.din(new_net_16612),
		.dout(new_net_16613)
	);

	bfr new_net_16614_bfr_after (
		.din(new_net_16613),
		.dout(new_net_16614)
	);

	bfr new_net_16615_bfr_after (
		.din(new_net_16614),
		.dout(new_net_16615)
	);

	bfr new_net_16616_bfr_after (
		.din(new_net_16615),
		.dout(new_net_16616)
	);

	bfr new_net_16617_bfr_after (
		.din(new_net_16616),
		.dout(new_net_16617)
	);

	bfr new_net_16618_bfr_after (
		.din(new_net_16617),
		.dout(new_net_16618)
	);

	bfr new_net_16619_bfr_after (
		.din(new_net_16618),
		.dout(new_net_16619)
	);

	bfr new_net_16620_bfr_after (
		.din(new_net_16619),
		.dout(new_net_16620)
	);

	bfr new_net_16621_bfr_after (
		.din(new_net_16620),
		.dout(new_net_16621)
	);

	bfr new_net_16622_bfr_after (
		.din(new_net_16621),
		.dout(new_net_16622)
	);

	bfr new_net_16623_bfr_after (
		.din(new_net_16622),
		.dout(new_net_16623)
	);

	bfr new_net_16624_bfr_after (
		.din(new_net_16623),
		.dout(new_net_16624)
	);

	bfr new_net_16625_bfr_after (
		.din(new_net_16624),
		.dout(new_net_16625)
	);

	bfr new_net_16626_bfr_after (
		.din(new_net_16625),
		.dout(new_net_16626)
	);

	bfr new_net_16627_bfr_after (
		.din(new_net_16626),
		.dout(new_net_16627)
	);

	bfr new_net_16628_bfr_after (
		.din(new_net_16627),
		.dout(new_net_16628)
	);

	spl2 _0548__v_fanout (
		.a(new_net_16628),
		.b(new_net_12),
		.c(new_net_13)
	);

	bfr new_net_16629_bfr_after (
		.din(_1373_),
		.dout(new_net_16629)
	);

	bfr new_net_16630_bfr_after (
		.din(new_net_16629),
		.dout(new_net_16630)
	);

	bfr new_net_16631_bfr_after (
		.din(new_net_16630),
		.dout(new_net_16631)
	);

	bfr new_net_16632_bfr_after (
		.din(new_net_16631),
		.dout(new_net_16632)
	);

	bfr new_net_16633_bfr_after (
		.din(new_net_16632),
		.dout(new_net_16633)
	);

	bfr new_net_16634_bfr_after (
		.din(new_net_16633),
		.dout(new_net_16634)
	);

	bfr new_net_16635_bfr_after (
		.din(new_net_16634),
		.dout(new_net_16635)
	);

	bfr new_net_16636_bfr_after (
		.din(new_net_16635),
		.dout(new_net_16636)
	);

	bfr new_net_16637_bfr_after (
		.din(new_net_16636),
		.dout(new_net_16637)
	);

	bfr new_net_16638_bfr_after (
		.din(new_net_16637),
		.dout(new_net_16638)
	);

	bfr new_net_16639_bfr_after (
		.din(new_net_16638),
		.dout(new_net_16639)
	);

	bfr new_net_16640_bfr_after (
		.din(new_net_16639),
		.dout(new_net_16640)
	);

	bfr new_net_16641_bfr_after (
		.din(new_net_16640),
		.dout(new_net_16641)
	);

	bfr new_net_16642_bfr_after (
		.din(new_net_16641),
		.dout(new_net_16642)
	);

	bfr new_net_16643_bfr_after (
		.din(new_net_16642),
		.dout(new_net_16643)
	);

	bfr new_net_16644_bfr_after (
		.din(new_net_16643),
		.dout(new_net_16644)
	);

	bfr new_net_16645_bfr_after (
		.din(new_net_16644),
		.dout(new_net_16645)
	);

	bfr new_net_16646_bfr_after (
		.din(new_net_16645),
		.dout(new_net_16646)
	);

	bfr new_net_16647_bfr_after (
		.din(new_net_16646),
		.dout(new_net_16647)
	);

	bfr new_net_16648_bfr_after (
		.din(new_net_16647),
		.dout(new_net_16648)
	);

	bfr new_net_16649_bfr_after (
		.din(new_net_16648),
		.dout(new_net_16649)
	);

	bfr new_net_16650_bfr_after (
		.din(new_net_16649),
		.dout(new_net_16650)
	);

	bfr new_net_16651_bfr_after (
		.din(new_net_16650),
		.dout(new_net_16651)
	);

	bfr new_net_16652_bfr_after (
		.din(new_net_16651),
		.dout(new_net_16652)
	);

	bfr new_net_16653_bfr_after (
		.din(new_net_16652),
		.dout(new_net_16653)
	);

	bfr new_net_16654_bfr_after (
		.din(new_net_16653),
		.dout(new_net_16654)
	);

	bfr new_net_16655_bfr_after (
		.din(new_net_16654),
		.dout(new_net_16655)
	);

	bfr new_net_16656_bfr_after (
		.din(new_net_16655),
		.dout(new_net_16656)
	);

	bfr new_net_16657_bfr_after (
		.din(new_net_16656),
		.dout(new_net_16657)
	);

	bfr new_net_16658_bfr_after (
		.din(new_net_16657),
		.dout(new_net_16658)
	);

	bfr new_net_16659_bfr_after (
		.din(new_net_16658),
		.dout(new_net_16659)
	);

	bfr new_net_16660_bfr_after (
		.din(new_net_16659),
		.dout(new_net_16660)
	);

	bfr new_net_16661_bfr_after (
		.din(new_net_16660),
		.dout(new_net_16661)
	);

	bfr new_net_16662_bfr_after (
		.din(new_net_16661),
		.dout(new_net_16662)
	);

	bfr new_net_16663_bfr_after (
		.din(new_net_16662),
		.dout(new_net_16663)
	);

	bfr new_net_16664_bfr_after (
		.din(new_net_16663),
		.dout(new_net_16664)
	);

	bfr new_net_16665_bfr_after (
		.din(new_net_16664),
		.dout(new_net_16665)
	);

	bfr new_net_16666_bfr_after (
		.din(new_net_16665),
		.dout(new_net_16666)
	);

	bfr new_net_16667_bfr_after (
		.din(new_net_16666),
		.dout(new_net_16667)
	);

	bfr new_net_16668_bfr_after (
		.din(new_net_16667),
		.dout(new_net_16668)
	);

	spl2 _1373__v_fanout (
		.a(new_net_16668),
		.b(new_net_2028),
		.c(new_net_2029)
	);

	bfr new_net_16669_bfr_after (
		.din(_1361_),
		.dout(new_net_16669)
	);

	bfr new_net_16670_bfr_after (
		.din(new_net_16669),
		.dout(new_net_16670)
	);

	bfr new_net_16671_bfr_after (
		.din(new_net_16670),
		.dout(new_net_16671)
	);

	bfr new_net_16672_bfr_after (
		.din(new_net_16671),
		.dout(new_net_16672)
	);

	bfr new_net_16673_bfr_after (
		.din(new_net_16672),
		.dout(new_net_16673)
	);

	bfr new_net_16674_bfr_after (
		.din(new_net_16673),
		.dout(new_net_16674)
	);

	bfr new_net_16675_bfr_after (
		.din(new_net_16674),
		.dout(new_net_16675)
	);

	bfr new_net_16676_bfr_after (
		.din(new_net_16675),
		.dout(new_net_16676)
	);

	bfr new_net_16677_bfr_after (
		.din(new_net_16676),
		.dout(new_net_16677)
	);

	bfr new_net_16678_bfr_after (
		.din(new_net_16677),
		.dout(new_net_16678)
	);

	bfr new_net_16679_bfr_after (
		.din(new_net_16678),
		.dout(new_net_16679)
	);

	bfr new_net_16680_bfr_after (
		.din(new_net_16679),
		.dout(new_net_16680)
	);

	bfr new_net_16681_bfr_after (
		.din(new_net_16680),
		.dout(new_net_16681)
	);

	bfr new_net_16682_bfr_after (
		.din(new_net_16681),
		.dout(new_net_16682)
	);

	bfr new_net_16683_bfr_after (
		.din(new_net_16682),
		.dout(new_net_16683)
	);

	bfr new_net_16684_bfr_after (
		.din(new_net_16683),
		.dout(new_net_16684)
	);

	bfr new_net_16685_bfr_after (
		.din(new_net_16684),
		.dout(new_net_16685)
	);

	bfr new_net_16686_bfr_after (
		.din(new_net_16685),
		.dout(new_net_16686)
	);

	bfr new_net_16687_bfr_after (
		.din(new_net_16686),
		.dout(new_net_16687)
	);

	bfr new_net_16688_bfr_after (
		.din(new_net_16687),
		.dout(new_net_16688)
	);

	bfr new_net_16689_bfr_after (
		.din(new_net_16688),
		.dout(new_net_16689)
	);

	bfr new_net_16690_bfr_after (
		.din(new_net_16689),
		.dout(new_net_16690)
	);

	bfr new_net_16691_bfr_after (
		.din(new_net_16690),
		.dout(new_net_16691)
	);

	bfr new_net_16692_bfr_after (
		.din(new_net_16691),
		.dout(new_net_16692)
	);

	bfr new_net_16693_bfr_after (
		.din(new_net_16692),
		.dout(new_net_16693)
	);

	bfr new_net_16694_bfr_after (
		.din(new_net_16693),
		.dout(new_net_16694)
	);

	bfr new_net_16695_bfr_after (
		.din(new_net_16694),
		.dout(new_net_16695)
	);

	bfr new_net_16696_bfr_after (
		.din(new_net_16695),
		.dout(new_net_16696)
	);

	bfr new_net_16697_bfr_after (
		.din(new_net_16696),
		.dout(new_net_16697)
	);

	bfr new_net_16698_bfr_after (
		.din(new_net_16697),
		.dout(new_net_16698)
	);

	bfr new_net_16699_bfr_after (
		.din(new_net_16698),
		.dout(new_net_16699)
	);

	bfr new_net_16700_bfr_after (
		.din(new_net_16699),
		.dout(new_net_16700)
	);

	bfr new_net_16701_bfr_after (
		.din(new_net_16700),
		.dout(new_net_16701)
	);

	bfr new_net_16702_bfr_after (
		.din(new_net_16701),
		.dout(new_net_16702)
	);

	bfr new_net_16703_bfr_after (
		.din(new_net_16702),
		.dout(new_net_16703)
	);

	bfr new_net_16704_bfr_after (
		.din(new_net_16703),
		.dout(new_net_16704)
	);

	bfr new_net_16705_bfr_after (
		.din(new_net_16704),
		.dout(new_net_16705)
	);

	bfr new_net_16706_bfr_after (
		.din(new_net_16705),
		.dout(new_net_16706)
	);

	bfr new_net_16707_bfr_after (
		.din(new_net_16706),
		.dout(new_net_16707)
	);

	bfr new_net_16708_bfr_after (
		.din(new_net_16707),
		.dout(new_net_16708)
	);

	bfr new_net_16709_bfr_after (
		.din(new_net_16708),
		.dout(new_net_16709)
	);

	bfr new_net_16710_bfr_after (
		.din(new_net_16709),
		.dout(new_net_16710)
	);

	bfr new_net_16711_bfr_after (
		.din(new_net_16710),
		.dout(new_net_16711)
	);

	bfr new_net_16712_bfr_after (
		.din(new_net_16711),
		.dout(new_net_16712)
	);

	bfr new_net_16713_bfr_after (
		.din(new_net_16712),
		.dout(new_net_16713)
	);

	bfr new_net_16714_bfr_after (
		.din(new_net_16713),
		.dout(new_net_16714)
	);

	bfr new_net_16715_bfr_after (
		.din(new_net_16714),
		.dout(new_net_16715)
	);

	bfr new_net_16716_bfr_after (
		.din(new_net_16715),
		.dout(new_net_16716)
	);

	bfr new_net_16717_bfr_after (
		.din(new_net_16716),
		.dout(new_net_16717)
	);

	bfr new_net_16718_bfr_after (
		.din(new_net_16717),
		.dout(new_net_16718)
	);

	bfr new_net_16719_bfr_after (
		.din(new_net_16718),
		.dout(new_net_16719)
	);

	bfr new_net_16720_bfr_after (
		.din(new_net_16719),
		.dout(new_net_16720)
	);

	bfr new_net_16721_bfr_after (
		.din(new_net_16720),
		.dout(new_net_16721)
	);

	bfr new_net_16722_bfr_after (
		.din(new_net_16721),
		.dout(new_net_16722)
	);

	bfr new_net_16723_bfr_after (
		.din(new_net_16722),
		.dout(new_net_16723)
	);

	bfr new_net_16724_bfr_after (
		.din(new_net_16723),
		.dout(new_net_16724)
	);

	bfr new_net_16725_bfr_after (
		.din(new_net_16724),
		.dout(new_net_16725)
	);

	bfr new_net_16726_bfr_after (
		.din(new_net_16725),
		.dout(new_net_16726)
	);

	bfr new_net_16727_bfr_after (
		.din(new_net_16726),
		.dout(new_net_16727)
	);

	bfr new_net_16728_bfr_after (
		.din(new_net_16727),
		.dout(new_net_16728)
	);

	bfr new_net_16729_bfr_after (
		.din(new_net_16728),
		.dout(new_net_16729)
	);

	bfr new_net_16730_bfr_after (
		.din(new_net_16729),
		.dout(new_net_16730)
	);

	bfr new_net_16731_bfr_after (
		.din(new_net_16730),
		.dout(new_net_16731)
	);

	bfr new_net_16732_bfr_after (
		.din(new_net_16731),
		.dout(new_net_16732)
	);

	bfr new_net_16733_bfr_after (
		.din(new_net_16732),
		.dout(new_net_16733)
	);

	bfr new_net_16734_bfr_after (
		.din(new_net_16733),
		.dout(new_net_16734)
	);

	bfr new_net_16735_bfr_after (
		.din(new_net_16734),
		.dout(new_net_16735)
	);

	bfr new_net_16736_bfr_after (
		.din(new_net_16735),
		.dout(new_net_16736)
	);

	bfr new_net_16737_bfr_after (
		.din(new_net_16736),
		.dout(new_net_16737)
	);

	bfr new_net_16738_bfr_after (
		.din(new_net_16737),
		.dout(new_net_16738)
	);

	bfr new_net_16739_bfr_after (
		.din(new_net_16738),
		.dout(new_net_16739)
	);

	bfr new_net_16740_bfr_after (
		.din(new_net_16739),
		.dout(new_net_16740)
	);

	bfr new_net_16741_bfr_after (
		.din(new_net_16740),
		.dout(new_net_16741)
	);

	bfr new_net_16742_bfr_after (
		.din(new_net_16741),
		.dout(new_net_16742)
	);

	bfr new_net_16743_bfr_after (
		.din(new_net_16742),
		.dout(new_net_16743)
	);

	bfr new_net_16744_bfr_after (
		.din(new_net_16743),
		.dout(new_net_16744)
	);

	bfr new_net_16745_bfr_after (
		.din(new_net_16744),
		.dout(new_net_16745)
	);

	bfr new_net_16746_bfr_after (
		.din(new_net_16745),
		.dout(new_net_16746)
	);

	bfr new_net_16747_bfr_after (
		.din(new_net_16746),
		.dout(new_net_16747)
	);

	bfr new_net_16748_bfr_after (
		.din(new_net_16747),
		.dout(new_net_16748)
	);

	bfr new_net_16749_bfr_after (
		.din(new_net_16748),
		.dout(new_net_16749)
	);

	bfr new_net_16750_bfr_after (
		.din(new_net_16749),
		.dout(new_net_16750)
	);

	bfr new_net_16751_bfr_after (
		.din(new_net_16750),
		.dout(new_net_16751)
	);

	bfr new_net_16752_bfr_after (
		.din(new_net_16751),
		.dout(new_net_16752)
	);

	bfr new_net_16753_bfr_after (
		.din(new_net_16752),
		.dout(new_net_16753)
	);

	bfr new_net_16754_bfr_after (
		.din(new_net_16753),
		.dout(new_net_16754)
	);

	bfr new_net_16755_bfr_after (
		.din(new_net_16754),
		.dout(new_net_16755)
	);

	bfr new_net_16756_bfr_after (
		.din(new_net_16755),
		.dout(new_net_16756)
	);

	spl2 _1361__v_fanout (
		.a(new_net_16756),
		.b(new_net_3059),
		.c(new_net_3060)
	);

	bfr new_net_16757_bfr_after (
		.din(_0216_),
		.dout(new_net_16757)
	);

	bfr new_net_16758_bfr_after (
		.din(new_net_16757),
		.dout(new_net_16758)
	);

	bfr new_net_16759_bfr_after (
		.din(new_net_16758),
		.dout(new_net_16759)
	);

	bfr new_net_16760_bfr_after (
		.din(new_net_16759),
		.dout(new_net_16760)
	);

	bfr new_net_16761_bfr_after (
		.din(new_net_16760),
		.dout(new_net_16761)
	);

	bfr new_net_16762_bfr_after (
		.din(new_net_16761),
		.dout(new_net_16762)
	);

	bfr new_net_16763_bfr_after (
		.din(new_net_16762),
		.dout(new_net_16763)
	);

	bfr new_net_16764_bfr_after (
		.din(new_net_16763),
		.dout(new_net_16764)
	);

	bfr new_net_16765_bfr_after (
		.din(new_net_16764),
		.dout(new_net_16765)
	);

	bfr new_net_16766_bfr_after (
		.din(new_net_16765),
		.dout(new_net_16766)
	);

	bfr new_net_16767_bfr_after (
		.din(new_net_16766),
		.dout(new_net_16767)
	);

	bfr new_net_16768_bfr_after (
		.din(new_net_16767),
		.dout(new_net_16768)
	);

	bfr new_net_16769_bfr_after (
		.din(new_net_16768),
		.dout(new_net_16769)
	);

	bfr new_net_16770_bfr_after (
		.din(new_net_16769),
		.dout(new_net_16770)
	);

	bfr new_net_16771_bfr_after (
		.din(new_net_16770),
		.dout(new_net_16771)
	);

	bfr new_net_16772_bfr_after (
		.din(new_net_16771),
		.dout(new_net_16772)
	);

	bfr new_net_16773_bfr_after (
		.din(new_net_16772),
		.dout(new_net_16773)
	);

	bfr new_net_16774_bfr_after (
		.din(new_net_16773),
		.dout(new_net_16774)
	);

	bfr new_net_16775_bfr_after (
		.din(new_net_16774),
		.dout(new_net_16775)
	);

	bfr new_net_16776_bfr_after (
		.din(new_net_16775),
		.dout(new_net_16776)
	);

	bfr new_net_16777_bfr_after (
		.din(new_net_16776),
		.dout(new_net_16777)
	);

	bfr new_net_16778_bfr_after (
		.din(new_net_16777),
		.dout(new_net_16778)
	);

	bfr new_net_16779_bfr_after (
		.din(new_net_16778),
		.dout(new_net_16779)
	);

	bfr new_net_16780_bfr_after (
		.din(new_net_16779),
		.dout(new_net_16780)
	);

	bfr new_net_16781_bfr_after (
		.din(new_net_16780),
		.dout(new_net_16781)
	);

	bfr new_net_16782_bfr_after (
		.din(new_net_16781),
		.dout(new_net_16782)
	);

	bfr new_net_16783_bfr_after (
		.din(new_net_16782),
		.dout(new_net_16783)
	);

	bfr new_net_16784_bfr_after (
		.din(new_net_16783),
		.dout(new_net_16784)
	);

	bfr new_net_16785_bfr_after (
		.din(new_net_16784),
		.dout(new_net_16785)
	);

	bfr new_net_16786_bfr_after (
		.din(new_net_16785),
		.dout(new_net_16786)
	);

	bfr new_net_16787_bfr_after (
		.din(new_net_16786),
		.dout(new_net_16787)
	);

	bfr new_net_16788_bfr_after (
		.din(new_net_16787),
		.dout(new_net_16788)
	);

	bfr new_net_16789_bfr_after (
		.din(new_net_16788),
		.dout(new_net_16789)
	);

	bfr new_net_16790_bfr_after (
		.din(new_net_16789),
		.dout(new_net_16790)
	);

	bfr new_net_16791_bfr_after (
		.din(new_net_16790),
		.dout(new_net_16791)
	);

	bfr new_net_16792_bfr_after (
		.din(new_net_16791),
		.dout(new_net_16792)
	);

	bfr new_net_16793_bfr_after (
		.din(new_net_16792),
		.dout(new_net_16793)
	);

	bfr new_net_16794_bfr_after (
		.din(new_net_16793),
		.dout(new_net_16794)
	);

	bfr new_net_16795_bfr_after (
		.din(new_net_16794),
		.dout(new_net_16795)
	);

	bfr new_net_16796_bfr_after (
		.din(new_net_16795),
		.dout(new_net_16796)
	);

	bfr new_net_16797_bfr_after (
		.din(new_net_16796),
		.dout(new_net_16797)
	);

	bfr new_net_16798_bfr_after (
		.din(new_net_16797),
		.dout(new_net_16798)
	);

	bfr new_net_16799_bfr_after (
		.din(new_net_16798),
		.dout(new_net_16799)
	);

	bfr new_net_16800_bfr_after (
		.din(new_net_16799),
		.dout(new_net_16800)
	);

	bfr new_net_16801_bfr_after (
		.din(new_net_16800),
		.dout(new_net_16801)
	);

	bfr new_net_16802_bfr_after (
		.din(new_net_16801),
		.dout(new_net_16802)
	);

	bfr new_net_16803_bfr_after (
		.din(new_net_16802),
		.dout(new_net_16803)
	);

	bfr new_net_16804_bfr_after (
		.din(new_net_16803),
		.dout(new_net_16804)
	);

	bfr new_net_16805_bfr_after (
		.din(new_net_16804),
		.dout(new_net_16805)
	);

	bfr new_net_16806_bfr_after (
		.din(new_net_16805),
		.dout(new_net_16806)
	);

	bfr new_net_16807_bfr_after (
		.din(new_net_16806),
		.dout(new_net_16807)
	);

	bfr new_net_16808_bfr_after (
		.din(new_net_16807),
		.dout(new_net_16808)
	);

	bfr new_net_16809_bfr_after (
		.din(new_net_16808),
		.dout(new_net_16809)
	);

	bfr new_net_16810_bfr_after (
		.din(new_net_16809),
		.dout(new_net_16810)
	);

	bfr new_net_16811_bfr_after (
		.din(new_net_16810),
		.dout(new_net_16811)
	);

	bfr new_net_16812_bfr_after (
		.din(new_net_16811),
		.dout(new_net_16812)
	);

	bfr new_net_16813_bfr_after (
		.din(new_net_16812),
		.dout(new_net_16813)
	);

	bfr new_net_16814_bfr_after (
		.din(new_net_16813),
		.dout(new_net_16814)
	);

	bfr new_net_16815_bfr_after (
		.din(new_net_16814),
		.dout(new_net_16815)
	);

	bfr new_net_16816_bfr_after (
		.din(new_net_16815),
		.dout(new_net_16816)
	);

	bfr new_net_16817_bfr_after (
		.din(new_net_16816),
		.dout(new_net_16817)
	);

	bfr new_net_16818_bfr_after (
		.din(new_net_16817),
		.dout(new_net_16818)
	);

	bfr new_net_16819_bfr_after (
		.din(new_net_16818),
		.dout(new_net_16819)
	);

	bfr new_net_16820_bfr_after (
		.din(new_net_16819),
		.dout(new_net_16820)
	);

	bfr new_net_16821_bfr_after (
		.din(new_net_16820),
		.dout(new_net_16821)
	);

	bfr new_net_16822_bfr_after (
		.din(new_net_16821),
		.dout(new_net_16822)
	);

	bfr new_net_16823_bfr_after (
		.din(new_net_16822),
		.dout(new_net_16823)
	);

	bfr new_net_16824_bfr_after (
		.din(new_net_16823),
		.dout(new_net_16824)
	);

	bfr new_net_16825_bfr_after (
		.din(new_net_16824),
		.dout(new_net_16825)
	);

	bfr new_net_16826_bfr_after (
		.din(new_net_16825),
		.dout(new_net_16826)
	);

	bfr new_net_16827_bfr_after (
		.din(new_net_16826),
		.dout(new_net_16827)
	);

	bfr new_net_16828_bfr_after (
		.din(new_net_16827),
		.dout(new_net_16828)
	);

	bfr new_net_16829_bfr_after (
		.din(new_net_16828),
		.dout(new_net_16829)
	);

	bfr new_net_16830_bfr_after (
		.din(new_net_16829),
		.dout(new_net_16830)
	);

	bfr new_net_16831_bfr_after (
		.din(new_net_16830),
		.dout(new_net_16831)
	);

	bfr new_net_16832_bfr_after (
		.din(new_net_16831),
		.dout(new_net_16832)
	);

	bfr new_net_16833_bfr_after (
		.din(new_net_16832),
		.dout(new_net_16833)
	);

	bfr new_net_16834_bfr_after (
		.din(new_net_16833),
		.dout(new_net_16834)
	);

	bfr new_net_16835_bfr_after (
		.din(new_net_16834),
		.dout(new_net_16835)
	);

	bfr new_net_16836_bfr_after (
		.din(new_net_16835),
		.dout(new_net_16836)
	);

	bfr new_net_16837_bfr_after (
		.din(new_net_16836),
		.dout(new_net_16837)
	);

	bfr new_net_16838_bfr_after (
		.din(new_net_16837),
		.dout(new_net_16838)
	);

	bfr new_net_16839_bfr_after (
		.din(new_net_16838),
		.dout(new_net_16839)
	);

	bfr new_net_16840_bfr_after (
		.din(new_net_16839),
		.dout(new_net_16840)
	);

	bfr new_net_16841_bfr_after (
		.din(new_net_16840),
		.dout(new_net_16841)
	);

	bfr new_net_16842_bfr_after (
		.din(new_net_16841),
		.dout(new_net_16842)
	);

	bfr new_net_16843_bfr_after (
		.din(new_net_16842),
		.dout(new_net_16843)
	);

	bfr new_net_16844_bfr_after (
		.din(new_net_16843),
		.dout(new_net_16844)
	);

	bfr new_net_16845_bfr_after (
		.din(new_net_16844),
		.dout(new_net_16845)
	);

	bfr new_net_16846_bfr_after (
		.din(new_net_16845),
		.dout(new_net_16846)
	);

	bfr new_net_16847_bfr_after (
		.din(new_net_16846),
		.dout(new_net_16847)
	);

	bfr new_net_16848_bfr_after (
		.din(new_net_16847),
		.dout(new_net_16848)
	);

	bfr new_net_16849_bfr_after (
		.din(new_net_16848),
		.dout(new_net_16849)
	);

	bfr new_net_16850_bfr_after (
		.din(new_net_16849),
		.dout(new_net_16850)
	);

	bfr new_net_16851_bfr_after (
		.din(new_net_16850),
		.dout(new_net_16851)
	);

	bfr new_net_16852_bfr_after (
		.din(new_net_16851),
		.dout(new_net_16852)
	);

	spl2 _0216__v_fanout (
		.a(new_net_16852),
		.b(new_net_2331),
		.c(new_net_2332)
	);

	bfr new_net_16853_bfr_after (
		.din(_1702_),
		.dout(new_net_16853)
	);

	bfr new_net_16854_bfr_after (
		.din(new_net_16853),
		.dout(new_net_16854)
	);

	bfr new_net_16855_bfr_after (
		.din(new_net_16854),
		.dout(new_net_16855)
	);

	bfr new_net_16856_bfr_after (
		.din(new_net_16855),
		.dout(new_net_16856)
	);

	bfr new_net_16857_bfr_after (
		.din(new_net_16856),
		.dout(new_net_16857)
	);

	bfr new_net_16858_bfr_after (
		.din(new_net_16857),
		.dout(new_net_16858)
	);

	bfr new_net_16859_bfr_after (
		.din(new_net_16858),
		.dout(new_net_16859)
	);

	bfr new_net_16860_bfr_after (
		.din(new_net_16859),
		.dout(new_net_16860)
	);

	bfr new_net_16861_bfr_after (
		.din(new_net_16860),
		.dout(new_net_16861)
	);

	bfr new_net_16862_bfr_after (
		.din(new_net_16861),
		.dout(new_net_16862)
	);

	bfr new_net_16863_bfr_after (
		.din(new_net_16862),
		.dout(new_net_16863)
	);

	bfr new_net_16864_bfr_after (
		.din(new_net_16863),
		.dout(new_net_16864)
	);

	bfr new_net_16865_bfr_after (
		.din(new_net_16864),
		.dout(new_net_16865)
	);

	bfr new_net_16866_bfr_after (
		.din(new_net_16865),
		.dout(new_net_16866)
	);

	bfr new_net_16867_bfr_after (
		.din(new_net_16866),
		.dout(new_net_16867)
	);

	bfr new_net_16868_bfr_after (
		.din(new_net_16867),
		.dout(new_net_16868)
	);

	bfr new_net_16869_bfr_after (
		.din(new_net_16868),
		.dout(new_net_16869)
	);

	bfr new_net_16870_bfr_after (
		.din(new_net_16869),
		.dout(new_net_16870)
	);

	bfr new_net_16871_bfr_after (
		.din(new_net_16870),
		.dout(new_net_16871)
	);

	bfr new_net_16872_bfr_after (
		.din(new_net_16871),
		.dout(new_net_16872)
	);

	bfr new_net_16873_bfr_after (
		.din(new_net_16872),
		.dout(new_net_16873)
	);

	bfr new_net_16874_bfr_after (
		.din(new_net_16873),
		.dout(new_net_16874)
	);

	bfr new_net_16875_bfr_after (
		.din(new_net_16874),
		.dout(new_net_16875)
	);

	bfr new_net_16876_bfr_after (
		.din(new_net_16875),
		.dout(new_net_16876)
	);

	spl2 _1702__v_fanout (
		.a(new_net_16876),
		.b(new_net_1880),
		.c(new_net_1881)
	);

	spl2 _1145__v_fanout (
		.a(_1145_),
		.b(new_net_1467),
		.c(new_net_1468)
	);

	bfr new_net_16877_bfr_after (
		.din(_1562_),
		.dout(new_net_16877)
	);

	bfr new_net_16878_bfr_after (
		.din(new_net_16877),
		.dout(new_net_16878)
	);

	bfr new_net_16879_bfr_after (
		.din(new_net_16878),
		.dout(new_net_16879)
	);

	bfr new_net_16880_bfr_after (
		.din(new_net_16879),
		.dout(new_net_16880)
	);

	bfr new_net_16881_bfr_after (
		.din(new_net_16880),
		.dout(new_net_16881)
	);

	bfr new_net_16882_bfr_after (
		.din(new_net_16881),
		.dout(new_net_16882)
	);

	bfr new_net_16883_bfr_after (
		.din(new_net_16882),
		.dout(new_net_16883)
	);

	bfr new_net_16884_bfr_after (
		.din(new_net_16883),
		.dout(new_net_16884)
	);

	bfr new_net_16885_bfr_after (
		.din(new_net_16884),
		.dout(new_net_16885)
	);

	bfr new_net_16886_bfr_after (
		.din(new_net_16885),
		.dout(new_net_16886)
	);

	bfr new_net_16887_bfr_after (
		.din(new_net_16886),
		.dout(new_net_16887)
	);

	bfr new_net_16888_bfr_after (
		.din(new_net_16887),
		.dout(new_net_16888)
	);

	bfr new_net_16889_bfr_after (
		.din(new_net_16888),
		.dout(new_net_16889)
	);

	bfr new_net_16890_bfr_after (
		.din(new_net_16889),
		.dout(new_net_16890)
	);

	bfr new_net_16891_bfr_after (
		.din(new_net_16890),
		.dout(new_net_16891)
	);

	bfr new_net_16892_bfr_after (
		.din(new_net_16891),
		.dout(new_net_16892)
	);

	bfr new_net_16893_bfr_after (
		.din(new_net_16892),
		.dout(new_net_16893)
	);

	bfr new_net_16894_bfr_after (
		.din(new_net_16893),
		.dout(new_net_16894)
	);

	bfr new_net_16895_bfr_after (
		.din(new_net_16894),
		.dout(new_net_16895)
	);

	bfr new_net_16896_bfr_after (
		.din(new_net_16895),
		.dout(new_net_16896)
	);

	bfr new_net_16897_bfr_after (
		.din(new_net_16896),
		.dout(new_net_16897)
	);

	bfr new_net_16898_bfr_after (
		.din(new_net_16897),
		.dout(new_net_16898)
	);

	bfr new_net_16899_bfr_after (
		.din(new_net_16898),
		.dout(new_net_16899)
	);

	bfr new_net_16900_bfr_after (
		.din(new_net_16899),
		.dout(new_net_16900)
	);

	bfr new_net_16901_bfr_after (
		.din(new_net_16900),
		.dout(new_net_16901)
	);

	bfr new_net_16902_bfr_after (
		.din(new_net_16901),
		.dout(new_net_16902)
	);

	bfr new_net_16903_bfr_after (
		.din(new_net_16902),
		.dout(new_net_16903)
	);

	bfr new_net_16904_bfr_after (
		.din(new_net_16903),
		.dout(new_net_16904)
	);

	bfr new_net_16905_bfr_after (
		.din(new_net_16904),
		.dout(new_net_16905)
	);

	bfr new_net_16906_bfr_after (
		.din(new_net_16905),
		.dout(new_net_16906)
	);

	bfr new_net_16907_bfr_after (
		.din(new_net_16906),
		.dout(new_net_16907)
	);

	bfr new_net_16908_bfr_after (
		.din(new_net_16907),
		.dout(new_net_16908)
	);

	bfr new_net_16909_bfr_after (
		.din(new_net_16908),
		.dout(new_net_16909)
	);

	bfr new_net_16910_bfr_after (
		.din(new_net_16909),
		.dout(new_net_16910)
	);

	bfr new_net_16911_bfr_after (
		.din(new_net_16910),
		.dout(new_net_16911)
	);

	bfr new_net_16912_bfr_after (
		.din(new_net_16911),
		.dout(new_net_16912)
	);

	bfr new_net_16913_bfr_after (
		.din(new_net_16912),
		.dout(new_net_16913)
	);

	bfr new_net_16914_bfr_after (
		.din(new_net_16913),
		.dout(new_net_16914)
	);

	bfr new_net_16915_bfr_after (
		.din(new_net_16914),
		.dout(new_net_16915)
	);

	bfr new_net_16916_bfr_after (
		.din(new_net_16915),
		.dout(new_net_16916)
	);

	bfr new_net_16917_bfr_after (
		.din(new_net_16916),
		.dout(new_net_16917)
	);

	bfr new_net_16918_bfr_after (
		.din(new_net_16917),
		.dout(new_net_16918)
	);

	bfr new_net_16919_bfr_after (
		.din(new_net_16918),
		.dout(new_net_16919)
	);

	bfr new_net_16920_bfr_after (
		.din(new_net_16919),
		.dout(new_net_16920)
	);

	bfr new_net_16921_bfr_after (
		.din(new_net_16920),
		.dout(new_net_16921)
	);

	bfr new_net_16922_bfr_after (
		.din(new_net_16921),
		.dout(new_net_16922)
	);

	bfr new_net_16923_bfr_after (
		.din(new_net_16922),
		.dout(new_net_16923)
	);

	bfr new_net_16924_bfr_after (
		.din(new_net_16923),
		.dout(new_net_16924)
	);

	bfr new_net_16925_bfr_after (
		.din(new_net_16924),
		.dout(new_net_16925)
	);

	bfr new_net_16926_bfr_after (
		.din(new_net_16925),
		.dout(new_net_16926)
	);

	bfr new_net_16927_bfr_after (
		.din(new_net_16926),
		.dout(new_net_16927)
	);

	bfr new_net_16928_bfr_after (
		.din(new_net_16927),
		.dout(new_net_16928)
	);

	bfr new_net_16929_bfr_after (
		.din(new_net_16928),
		.dout(new_net_16929)
	);

	bfr new_net_16930_bfr_after (
		.din(new_net_16929),
		.dout(new_net_16930)
	);

	bfr new_net_16931_bfr_after (
		.din(new_net_16930),
		.dout(new_net_16931)
	);

	bfr new_net_16932_bfr_after (
		.din(new_net_16931),
		.dout(new_net_16932)
	);

	bfr new_net_16933_bfr_after (
		.din(new_net_16932),
		.dout(new_net_16933)
	);

	bfr new_net_16934_bfr_after (
		.din(new_net_16933),
		.dout(new_net_16934)
	);

	bfr new_net_16935_bfr_after (
		.din(new_net_16934),
		.dout(new_net_16935)
	);

	bfr new_net_16936_bfr_after (
		.din(new_net_16935),
		.dout(new_net_16936)
	);

	bfr new_net_16937_bfr_after (
		.din(new_net_16936),
		.dout(new_net_16937)
	);

	bfr new_net_16938_bfr_after (
		.din(new_net_16937),
		.dout(new_net_16938)
	);

	bfr new_net_16939_bfr_after (
		.din(new_net_16938),
		.dout(new_net_16939)
	);

	bfr new_net_16940_bfr_after (
		.din(new_net_16939),
		.dout(new_net_16940)
	);

	bfr new_net_16941_bfr_after (
		.din(new_net_16940),
		.dout(new_net_16941)
	);

	bfr new_net_16942_bfr_after (
		.din(new_net_16941),
		.dout(new_net_16942)
	);

	bfr new_net_16943_bfr_after (
		.din(new_net_16942),
		.dout(new_net_16943)
	);

	bfr new_net_16944_bfr_after (
		.din(new_net_16943),
		.dout(new_net_16944)
	);

	bfr new_net_16945_bfr_after (
		.din(new_net_16944),
		.dout(new_net_16945)
	);

	bfr new_net_16946_bfr_after (
		.din(new_net_16945),
		.dout(new_net_16946)
	);

	bfr new_net_16947_bfr_after (
		.din(new_net_16946),
		.dout(new_net_16947)
	);

	bfr new_net_16948_bfr_after (
		.din(new_net_16947),
		.dout(new_net_16948)
	);

	bfr new_net_16949_bfr_after (
		.din(new_net_16948),
		.dout(new_net_16949)
	);

	bfr new_net_16950_bfr_after (
		.din(new_net_16949),
		.dout(new_net_16950)
	);

	bfr new_net_16951_bfr_after (
		.din(new_net_16950),
		.dout(new_net_16951)
	);

	bfr new_net_16952_bfr_after (
		.din(new_net_16951),
		.dout(new_net_16952)
	);

	bfr new_net_16953_bfr_after (
		.din(new_net_16952),
		.dout(new_net_16953)
	);

	bfr new_net_16954_bfr_after (
		.din(new_net_16953),
		.dout(new_net_16954)
	);

	bfr new_net_16955_bfr_after (
		.din(new_net_16954),
		.dout(new_net_16955)
	);

	bfr new_net_16956_bfr_after (
		.din(new_net_16955),
		.dout(new_net_16956)
	);

	bfr new_net_16957_bfr_after (
		.din(new_net_16956),
		.dout(new_net_16957)
	);

	bfr new_net_16958_bfr_after (
		.din(new_net_16957),
		.dout(new_net_16958)
	);

	bfr new_net_16959_bfr_after (
		.din(new_net_16958),
		.dout(new_net_16959)
	);

	bfr new_net_16960_bfr_after (
		.din(new_net_16959),
		.dout(new_net_16960)
	);

	bfr new_net_16961_bfr_after (
		.din(new_net_16960),
		.dout(new_net_16961)
	);

	bfr new_net_16962_bfr_after (
		.din(new_net_16961),
		.dout(new_net_16962)
	);

	bfr new_net_16963_bfr_after (
		.din(new_net_16962),
		.dout(new_net_16963)
	);

	bfr new_net_16964_bfr_after (
		.din(new_net_16963),
		.dout(new_net_16964)
	);

	bfr new_net_16965_bfr_after (
		.din(new_net_16964),
		.dout(new_net_16965)
	);

	bfr new_net_16966_bfr_after (
		.din(new_net_16965),
		.dout(new_net_16966)
	);

	bfr new_net_16967_bfr_after (
		.din(new_net_16966),
		.dout(new_net_16967)
	);

	bfr new_net_16968_bfr_after (
		.din(new_net_16967),
		.dout(new_net_16968)
	);

	bfr new_net_16969_bfr_after (
		.din(new_net_16968),
		.dout(new_net_16969)
	);

	bfr new_net_16970_bfr_after (
		.din(new_net_16969),
		.dout(new_net_16970)
	);

	bfr new_net_16971_bfr_after (
		.din(new_net_16970),
		.dout(new_net_16971)
	);

	bfr new_net_16972_bfr_after (
		.din(new_net_16971),
		.dout(new_net_16972)
	);

	spl2 _1562__v_fanout (
		.a(new_net_16972),
		.b(new_net_3001),
		.c(new_net_3002)
	);

	bfr new_net_16973_bfr_after (
		.din(_1693_),
		.dout(new_net_16973)
	);

	bfr new_net_16974_bfr_after (
		.din(new_net_16973),
		.dout(new_net_16974)
	);

	bfr new_net_16975_bfr_after (
		.din(new_net_16974),
		.dout(new_net_16975)
	);

	bfr new_net_16976_bfr_after (
		.din(new_net_16975),
		.dout(new_net_16976)
	);

	bfr new_net_16977_bfr_after (
		.din(new_net_16976),
		.dout(new_net_16977)
	);

	bfr new_net_16978_bfr_after (
		.din(new_net_16977),
		.dout(new_net_16978)
	);

	bfr new_net_16979_bfr_after (
		.din(new_net_16978),
		.dout(new_net_16979)
	);

	bfr new_net_16980_bfr_after (
		.din(new_net_16979),
		.dout(new_net_16980)
	);

	bfr new_net_16981_bfr_after (
		.din(new_net_16980),
		.dout(new_net_16981)
	);

	bfr new_net_16982_bfr_after (
		.din(new_net_16981),
		.dout(new_net_16982)
	);

	bfr new_net_16983_bfr_after (
		.din(new_net_16982),
		.dout(new_net_16983)
	);

	bfr new_net_16984_bfr_after (
		.din(new_net_16983),
		.dout(new_net_16984)
	);

	bfr new_net_16985_bfr_after (
		.din(new_net_16984),
		.dout(new_net_16985)
	);

	bfr new_net_16986_bfr_after (
		.din(new_net_16985),
		.dout(new_net_16986)
	);

	bfr new_net_16987_bfr_after (
		.din(new_net_16986),
		.dout(new_net_16987)
	);

	bfr new_net_16988_bfr_after (
		.din(new_net_16987),
		.dout(new_net_16988)
	);

	bfr new_net_16989_bfr_after (
		.din(new_net_16988),
		.dout(new_net_16989)
	);

	bfr new_net_16990_bfr_after (
		.din(new_net_16989),
		.dout(new_net_16990)
	);

	bfr new_net_16991_bfr_after (
		.din(new_net_16990),
		.dout(new_net_16991)
	);

	bfr new_net_16992_bfr_after (
		.din(new_net_16991),
		.dout(new_net_16992)
	);

	bfr new_net_16993_bfr_after (
		.din(new_net_16992),
		.dout(new_net_16993)
	);

	bfr new_net_16994_bfr_after (
		.din(new_net_16993),
		.dout(new_net_16994)
	);

	bfr new_net_16995_bfr_after (
		.din(new_net_16994),
		.dout(new_net_16995)
	);

	bfr new_net_16996_bfr_after (
		.din(new_net_16995),
		.dout(new_net_16996)
	);

	bfr new_net_16997_bfr_after (
		.din(new_net_16996),
		.dout(new_net_16997)
	);

	bfr new_net_16998_bfr_after (
		.din(new_net_16997),
		.dout(new_net_16998)
	);

	bfr new_net_16999_bfr_after (
		.din(new_net_16998),
		.dout(new_net_16999)
	);

	bfr new_net_17000_bfr_after (
		.din(new_net_16999),
		.dout(new_net_17000)
	);

	bfr new_net_17001_bfr_after (
		.din(new_net_17000),
		.dout(new_net_17001)
	);

	bfr new_net_17002_bfr_after (
		.din(new_net_17001),
		.dout(new_net_17002)
	);

	bfr new_net_17003_bfr_after (
		.din(new_net_17002),
		.dout(new_net_17003)
	);

	bfr new_net_17004_bfr_after (
		.din(new_net_17003),
		.dout(new_net_17004)
	);

	bfr new_net_17005_bfr_after (
		.din(new_net_17004),
		.dout(new_net_17005)
	);

	bfr new_net_17006_bfr_after (
		.din(new_net_17005),
		.dout(new_net_17006)
	);

	bfr new_net_17007_bfr_after (
		.din(new_net_17006),
		.dout(new_net_17007)
	);

	bfr new_net_17008_bfr_after (
		.din(new_net_17007),
		.dout(new_net_17008)
	);

	bfr new_net_17009_bfr_after (
		.din(new_net_17008),
		.dout(new_net_17009)
	);

	bfr new_net_17010_bfr_after (
		.din(new_net_17009),
		.dout(new_net_17010)
	);

	bfr new_net_17011_bfr_after (
		.din(new_net_17010),
		.dout(new_net_17011)
	);

	bfr new_net_17012_bfr_after (
		.din(new_net_17011),
		.dout(new_net_17012)
	);

	bfr new_net_17013_bfr_after (
		.din(new_net_17012),
		.dout(new_net_17013)
	);

	bfr new_net_17014_bfr_after (
		.din(new_net_17013),
		.dout(new_net_17014)
	);

	bfr new_net_17015_bfr_after (
		.din(new_net_17014),
		.dout(new_net_17015)
	);

	bfr new_net_17016_bfr_after (
		.din(new_net_17015),
		.dout(new_net_17016)
	);

	bfr new_net_17017_bfr_after (
		.din(new_net_17016),
		.dout(new_net_17017)
	);

	bfr new_net_17018_bfr_after (
		.din(new_net_17017),
		.dout(new_net_17018)
	);

	bfr new_net_17019_bfr_after (
		.din(new_net_17018),
		.dout(new_net_17019)
	);

	bfr new_net_17020_bfr_after (
		.din(new_net_17019),
		.dout(new_net_17020)
	);

	bfr new_net_17021_bfr_after (
		.din(new_net_17020),
		.dout(new_net_17021)
	);

	bfr new_net_17022_bfr_after (
		.din(new_net_17021),
		.dout(new_net_17022)
	);

	bfr new_net_17023_bfr_after (
		.din(new_net_17022),
		.dout(new_net_17023)
	);

	bfr new_net_17024_bfr_after (
		.din(new_net_17023),
		.dout(new_net_17024)
	);

	bfr new_net_17025_bfr_after (
		.din(new_net_17024),
		.dout(new_net_17025)
	);

	bfr new_net_17026_bfr_after (
		.din(new_net_17025),
		.dout(new_net_17026)
	);

	bfr new_net_17027_bfr_after (
		.din(new_net_17026),
		.dout(new_net_17027)
	);

	bfr new_net_17028_bfr_after (
		.din(new_net_17027),
		.dout(new_net_17028)
	);

	spl2 _1693__v_fanout (
		.a(new_net_17028),
		.b(new_net_1573),
		.c(new_net_1574)
	);

	bfr new_net_17029_bfr_after (
		.din(_1678_),
		.dout(new_net_17029)
	);

	bfr new_net_17030_bfr_after (
		.din(new_net_17029),
		.dout(new_net_17030)
	);

	bfr new_net_17031_bfr_after (
		.din(new_net_17030),
		.dout(new_net_17031)
	);

	bfr new_net_17032_bfr_after (
		.din(new_net_17031),
		.dout(new_net_17032)
	);

	bfr new_net_17033_bfr_after (
		.din(new_net_17032),
		.dout(new_net_17033)
	);

	bfr new_net_17034_bfr_after (
		.din(new_net_17033),
		.dout(new_net_17034)
	);

	bfr new_net_17035_bfr_after (
		.din(new_net_17034),
		.dout(new_net_17035)
	);

	bfr new_net_17036_bfr_after (
		.din(new_net_17035),
		.dout(new_net_17036)
	);

	bfr new_net_17037_bfr_after (
		.din(new_net_17036),
		.dout(new_net_17037)
	);

	bfr new_net_17038_bfr_after (
		.din(new_net_17037),
		.dout(new_net_17038)
	);

	bfr new_net_17039_bfr_after (
		.din(new_net_17038),
		.dout(new_net_17039)
	);

	bfr new_net_17040_bfr_after (
		.din(new_net_17039),
		.dout(new_net_17040)
	);

	bfr new_net_17041_bfr_after (
		.din(new_net_17040),
		.dout(new_net_17041)
	);

	bfr new_net_17042_bfr_after (
		.din(new_net_17041),
		.dout(new_net_17042)
	);

	bfr new_net_17043_bfr_after (
		.din(new_net_17042),
		.dout(new_net_17043)
	);

	bfr new_net_17044_bfr_after (
		.din(new_net_17043),
		.dout(new_net_17044)
	);

	bfr new_net_17045_bfr_after (
		.din(new_net_17044),
		.dout(new_net_17045)
	);

	bfr new_net_17046_bfr_after (
		.din(new_net_17045),
		.dout(new_net_17046)
	);

	bfr new_net_17047_bfr_after (
		.din(new_net_17046),
		.dout(new_net_17047)
	);

	bfr new_net_17048_bfr_after (
		.din(new_net_17047),
		.dout(new_net_17048)
	);

	bfr new_net_17049_bfr_after (
		.din(new_net_17048),
		.dout(new_net_17049)
	);

	bfr new_net_17050_bfr_after (
		.din(new_net_17049),
		.dout(new_net_17050)
	);

	bfr new_net_17051_bfr_after (
		.din(new_net_17050),
		.dout(new_net_17051)
	);

	bfr new_net_17052_bfr_after (
		.din(new_net_17051),
		.dout(new_net_17052)
	);

	bfr new_net_17053_bfr_after (
		.din(new_net_17052),
		.dout(new_net_17053)
	);

	bfr new_net_17054_bfr_after (
		.din(new_net_17053),
		.dout(new_net_17054)
	);

	bfr new_net_17055_bfr_after (
		.din(new_net_17054),
		.dout(new_net_17055)
	);

	bfr new_net_17056_bfr_after (
		.din(new_net_17055),
		.dout(new_net_17056)
	);

	bfr new_net_17057_bfr_after (
		.din(new_net_17056),
		.dout(new_net_17057)
	);

	bfr new_net_17058_bfr_after (
		.din(new_net_17057),
		.dout(new_net_17058)
	);

	bfr new_net_17059_bfr_after (
		.din(new_net_17058),
		.dout(new_net_17059)
	);

	bfr new_net_17060_bfr_after (
		.din(new_net_17059),
		.dout(new_net_17060)
	);

	bfr new_net_17061_bfr_after (
		.din(new_net_17060),
		.dout(new_net_17061)
	);

	bfr new_net_17062_bfr_after (
		.din(new_net_17061),
		.dout(new_net_17062)
	);

	bfr new_net_17063_bfr_after (
		.din(new_net_17062),
		.dout(new_net_17063)
	);

	bfr new_net_17064_bfr_after (
		.din(new_net_17063),
		.dout(new_net_17064)
	);

	bfr new_net_17065_bfr_after (
		.din(new_net_17064),
		.dout(new_net_17065)
	);

	bfr new_net_17066_bfr_after (
		.din(new_net_17065),
		.dout(new_net_17066)
	);

	bfr new_net_17067_bfr_after (
		.din(new_net_17066),
		.dout(new_net_17067)
	);

	bfr new_net_17068_bfr_after (
		.din(new_net_17067),
		.dout(new_net_17068)
	);

	bfr new_net_17069_bfr_after (
		.din(new_net_17068),
		.dout(new_net_17069)
	);

	bfr new_net_17070_bfr_after (
		.din(new_net_17069),
		.dout(new_net_17070)
	);

	bfr new_net_17071_bfr_after (
		.din(new_net_17070),
		.dout(new_net_17071)
	);

	bfr new_net_17072_bfr_after (
		.din(new_net_17071),
		.dout(new_net_17072)
	);

	bfr new_net_17073_bfr_after (
		.din(new_net_17072),
		.dout(new_net_17073)
	);

	bfr new_net_17074_bfr_after (
		.din(new_net_17073),
		.dout(new_net_17074)
	);

	bfr new_net_17075_bfr_after (
		.din(new_net_17074),
		.dout(new_net_17075)
	);

	bfr new_net_17076_bfr_after (
		.din(new_net_17075),
		.dout(new_net_17076)
	);

	bfr new_net_17077_bfr_after (
		.din(new_net_17076),
		.dout(new_net_17077)
	);

	bfr new_net_17078_bfr_after (
		.din(new_net_17077),
		.dout(new_net_17078)
	);

	bfr new_net_17079_bfr_after (
		.din(new_net_17078),
		.dout(new_net_17079)
	);

	bfr new_net_17080_bfr_after (
		.din(new_net_17079),
		.dout(new_net_17080)
	);

	bfr new_net_17081_bfr_after (
		.din(new_net_17080),
		.dout(new_net_17081)
	);

	bfr new_net_17082_bfr_after (
		.din(new_net_17081),
		.dout(new_net_17082)
	);

	bfr new_net_17083_bfr_after (
		.din(new_net_17082),
		.dout(new_net_17083)
	);

	bfr new_net_17084_bfr_after (
		.din(new_net_17083),
		.dout(new_net_17084)
	);

	bfr new_net_17085_bfr_after (
		.din(new_net_17084),
		.dout(new_net_17085)
	);

	bfr new_net_17086_bfr_after (
		.din(new_net_17085),
		.dout(new_net_17086)
	);

	bfr new_net_17087_bfr_after (
		.din(new_net_17086),
		.dout(new_net_17087)
	);

	bfr new_net_17088_bfr_after (
		.din(new_net_17087),
		.dout(new_net_17088)
	);

	bfr new_net_17089_bfr_after (
		.din(new_net_17088),
		.dout(new_net_17089)
	);

	bfr new_net_17090_bfr_after (
		.din(new_net_17089),
		.dout(new_net_17090)
	);

	bfr new_net_17091_bfr_after (
		.din(new_net_17090),
		.dout(new_net_17091)
	);

	bfr new_net_17092_bfr_after (
		.din(new_net_17091),
		.dout(new_net_17092)
	);

	bfr new_net_17093_bfr_after (
		.din(new_net_17092),
		.dout(new_net_17093)
	);

	bfr new_net_17094_bfr_after (
		.din(new_net_17093),
		.dout(new_net_17094)
	);

	bfr new_net_17095_bfr_after (
		.din(new_net_17094),
		.dout(new_net_17095)
	);

	bfr new_net_17096_bfr_after (
		.din(new_net_17095),
		.dout(new_net_17096)
	);

	bfr new_net_17097_bfr_after (
		.din(new_net_17096),
		.dout(new_net_17097)
	);

	bfr new_net_17098_bfr_after (
		.din(new_net_17097),
		.dout(new_net_17098)
	);

	bfr new_net_17099_bfr_after (
		.din(new_net_17098),
		.dout(new_net_17099)
	);

	bfr new_net_17100_bfr_after (
		.din(new_net_17099),
		.dout(new_net_17100)
	);

	bfr new_net_17101_bfr_after (
		.din(new_net_17100),
		.dout(new_net_17101)
	);

	bfr new_net_17102_bfr_after (
		.din(new_net_17101),
		.dout(new_net_17102)
	);

	bfr new_net_17103_bfr_after (
		.din(new_net_17102),
		.dout(new_net_17103)
	);

	bfr new_net_17104_bfr_after (
		.din(new_net_17103),
		.dout(new_net_17104)
	);

	bfr new_net_17105_bfr_after (
		.din(new_net_17104),
		.dout(new_net_17105)
	);

	bfr new_net_17106_bfr_after (
		.din(new_net_17105),
		.dout(new_net_17106)
	);

	bfr new_net_17107_bfr_after (
		.din(new_net_17106),
		.dout(new_net_17107)
	);

	bfr new_net_17108_bfr_after (
		.din(new_net_17107),
		.dout(new_net_17108)
	);

	bfr new_net_17109_bfr_after (
		.din(new_net_17108),
		.dout(new_net_17109)
	);

	bfr new_net_17110_bfr_after (
		.din(new_net_17109),
		.dout(new_net_17110)
	);

	bfr new_net_17111_bfr_after (
		.din(new_net_17110),
		.dout(new_net_17111)
	);

	bfr new_net_17112_bfr_after (
		.din(new_net_17111),
		.dout(new_net_17112)
	);

	bfr new_net_17113_bfr_after (
		.din(new_net_17112),
		.dout(new_net_17113)
	);

	bfr new_net_17114_bfr_after (
		.din(new_net_17113),
		.dout(new_net_17114)
	);

	bfr new_net_17115_bfr_after (
		.din(new_net_17114),
		.dout(new_net_17115)
	);

	bfr new_net_17116_bfr_after (
		.din(new_net_17115),
		.dout(new_net_17116)
	);

	bfr new_net_17117_bfr_after (
		.din(new_net_17116),
		.dout(new_net_17117)
	);

	bfr new_net_17118_bfr_after (
		.din(new_net_17117),
		.dout(new_net_17118)
	);

	bfr new_net_17119_bfr_after (
		.din(new_net_17118),
		.dout(new_net_17119)
	);

	bfr new_net_17120_bfr_after (
		.din(new_net_17119),
		.dout(new_net_17120)
	);

	bfr new_net_17121_bfr_after (
		.din(new_net_17120),
		.dout(new_net_17121)
	);

	bfr new_net_17122_bfr_after (
		.din(new_net_17121),
		.dout(new_net_17122)
	);

	bfr new_net_17123_bfr_after (
		.din(new_net_17122),
		.dout(new_net_17123)
	);

	bfr new_net_17124_bfr_after (
		.din(new_net_17123),
		.dout(new_net_17124)
	);

	bfr new_net_17125_bfr_after (
		.din(new_net_17124),
		.dout(new_net_17125)
	);

	bfr new_net_17126_bfr_after (
		.din(new_net_17125),
		.dout(new_net_17126)
	);

	bfr new_net_17127_bfr_after (
		.din(new_net_17126),
		.dout(new_net_17127)
	);

	bfr new_net_17128_bfr_after (
		.din(new_net_17127),
		.dout(new_net_17128)
	);

	bfr new_net_17129_bfr_after (
		.din(new_net_17128),
		.dout(new_net_17129)
	);

	bfr new_net_17130_bfr_after (
		.din(new_net_17129),
		.dout(new_net_17130)
	);

	bfr new_net_17131_bfr_after (
		.din(new_net_17130),
		.dout(new_net_17131)
	);

	bfr new_net_17132_bfr_after (
		.din(new_net_17131),
		.dout(new_net_17132)
	);

	bfr new_net_17133_bfr_after (
		.din(new_net_17132),
		.dout(new_net_17133)
	);

	bfr new_net_17134_bfr_after (
		.din(new_net_17133),
		.dout(new_net_17134)
	);

	bfr new_net_17135_bfr_after (
		.din(new_net_17134),
		.dout(new_net_17135)
	);

	bfr new_net_17136_bfr_after (
		.din(new_net_17135),
		.dout(new_net_17136)
	);

	bfr new_net_17137_bfr_after (
		.din(new_net_17136),
		.dout(new_net_17137)
	);

	bfr new_net_17138_bfr_after (
		.din(new_net_17137),
		.dout(new_net_17138)
	);

	bfr new_net_17139_bfr_after (
		.din(new_net_17138),
		.dout(new_net_17139)
	);

	bfr new_net_17140_bfr_after (
		.din(new_net_17139),
		.dout(new_net_17140)
	);

	spl2 _1678__v_fanout (
		.a(new_net_17140),
		.b(new_net_992),
		.c(new_net_993)
	);

	bfr new_net_17141_bfr_after (
		.din(_0988_),
		.dout(new_net_17141)
	);

	bfr new_net_17142_bfr_after (
		.din(new_net_17141),
		.dout(new_net_17142)
	);

	bfr new_net_17143_bfr_after (
		.din(new_net_17142),
		.dout(new_net_17143)
	);

	bfr new_net_17144_bfr_after (
		.din(new_net_17143),
		.dout(new_net_17144)
	);

	bfr new_net_17145_bfr_after (
		.din(new_net_17144),
		.dout(new_net_17145)
	);

	bfr new_net_17146_bfr_after (
		.din(new_net_17145),
		.dout(new_net_17146)
	);

	bfr new_net_17147_bfr_after (
		.din(new_net_17146),
		.dout(new_net_17147)
	);

	bfr new_net_17148_bfr_after (
		.din(new_net_17147),
		.dout(new_net_17148)
	);

	bfr new_net_17149_bfr_after (
		.din(new_net_17148),
		.dout(new_net_17149)
	);

	bfr new_net_17150_bfr_after (
		.din(new_net_17149),
		.dout(new_net_17150)
	);

	bfr new_net_17151_bfr_after (
		.din(new_net_17150),
		.dout(new_net_17151)
	);

	bfr new_net_17152_bfr_after (
		.din(new_net_17151),
		.dout(new_net_17152)
	);

	bfr new_net_17153_bfr_after (
		.din(new_net_17152),
		.dout(new_net_17153)
	);

	bfr new_net_17154_bfr_after (
		.din(new_net_17153),
		.dout(new_net_17154)
	);

	bfr new_net_17155_bfr_after (
		.din(new_net_17154),
		.dout(new_net_17155)
	);

	bfr new_net_17156_bfr_after (
		.din(new_net_17155),
		.dout(new_net_17156)
	);

	bfr new_net_17157_bfr_after (
		.din(new_net_17156),
		.dout(new_net_17157)
	);

	bfr new_net_17158_bfr_after (
		.din(new_net_17157),
		.dout(new_net_17158)
	);

	bfr new_net_17159_bfr_after (
		.din(new_net_17158),
		.dout(new_net_17159)
	);

	bfr new_net_17160_bfr_after (
		.din(new_net_17159),
		.dout(new_net_17160)
	);

	bfr new_net_17161_bfr_after (
		.din(new_net_17160),
		.dout(new_net_17161)
	);

	bfr new_net_17162_bfr_after (
		.din(new_net_17161),
		.dout(new_net_17162)
	);

	bfr new_net_17163_bfr_after (
		.din(new_net_17162),
		.dout(new_net_17163)
	);

	bfr new_net_17164_bfr_after (
		.din(new_net_17163),
		.dout(new_net_17164)
	);

	bfr new_net_17165_bfr_after (
		.din(new_net_17164),
		.dout(new_net_17165)
	);

	bfr new_net_17166_bfr_after (
		.din(new_net_17165),
		.dout(new_net_17166)
	);

	bfr new_net_17167_bfr_after (
		.din(new_net_17166),
		.dout(new_net_17167)
	);

	bfr new_net_17168_bfr_after (
		.din(new_net_17167),
		.dout(new_net_17168)
	);

	bfr new_net_17169_bfr_after (
		.din(new_net_17168),
		.dout(new_net_17169)
	);

	bfr new_net_17170_bfr_after (
		.din(new_net_17169),
		.dout(new_net_17170)
	);

	bfr new_net_17171_bfr_after (
		.din(new_net_17170),
		.dout(new_net_17171)
	);

	bfr new_net_17172_bfr_after (
		.din(new_net_17171),
		.dout(new_net_17172)
	);

	bfr new_net_17173_bfr_after (
		.din(new_net_17172),
		.dout(new_net_17173)
	);

	bfr new_net_17174_bfr_after (
		.din(new_net_17173),
		.dout(new_net_17174)
	);

	bfr new_net_17175_bfr_after (
		.din(new_net_17174),
		.dout(new_net_17175)
	);

	bfr new_net_17176_bfr_after (
		.din(new_net_17175),
		.dout(new_net_17176)
	);

	bfr new_net_17177_bfr_after (
		.din(new_net_17176),
		.dout(new_net_17177)
	);

	bfr new_net_17178_bfr_after (
		.din(new_net_17177),
		.dout(new_net_17178)
	);

	bfr new_net_17179_bfr_after (
		.din(new_net_17178),
		.dout(new_net_17179)
	);

	bfr new_net_17180_bfr_after (
		.din(new_net_17179),
		.dout(new_net_17180)
	);

	bfr new_net_17181_bfr_after (
		.din(new_net_17180),
		.dout(new_net_17181)
	);

	bfr new_net_17182_bfr_after (
		.din(new_net_17181),
		.dout(new_net_17182)
	);

	bfr new_net_17183_bfr_after (
		.din(new_net_17182),
		.dout(new_net_17183)
	);

	bfr new_net_17184_bfr_after (
		.din(new_net_17183),
		.dout(new_net_17184)
	);

	bfr new_net_17185_bfr_after (
		.din(new_net_17184),
		.dout(new_net_17185)
	);

	bfr new_net_17186_bfr_after (
		.din(new_net_17185),
		.dout(new_net_17186)
	);

	bfr new_net_17187_bfr_after (
		.din(new_net_17186),
		.dout(new_net_17187)
	);

	bfr new_net_17188_bfr_after (
		.din(new_net_17187),
		.dout(new_net_17188)
	);

	bfr new_net_17189_bfr_after (
		.din(new_net_17188),
		.dout(new_net_17189)
	);

	bfr new_net_17190_bfr_after (
		.din(new_net_17189),
		.dout(new_net_17190)
	);

	bfr new_net_17191_bfr_after (
		.din(new_net_17190),
		.dout(new_net_17191)
	);

	bfr new_net_17192_bfr_after (
		.din(new_net_17191),
		.dout(new_net_17192)
	);

	bfr new_net_17193_bfr_after (
		.din(new_net_17192),
		.dout(new_net_17193)
	);

	bfr new_net_17194_bfr_after (
		.din(new_net_17193),
		.dout(new_net_17194)
	);

	bfr new_net_17195_bfr_after (
		.din(new_net_17194),
		.dout(new_net_17195)
	);

	bfr new_net_17196_bfr_after (
		.din(new_net_17195),
		.dout(new_net_17196)
	);

	bfr new_net_17197_bfr_after (
		.din(new_net_17196),
		.dout(new_net_17197)
	);

	bfr new_net_17198_bfr_after (
		.din(new_net_17197),
		.dout(new_net_17198)
	);

	bfr new_net_17199_bfr_after (
		.din(new_net_17198),
		.dout(new_net_17199)
	);

	bfr new_net_17200_bfr_after (
		.din(new_net_17199),
		.dout(new_net_17200)
	);

	bfr new_net_17201_bfr_after (
		.din(new_net_17200),
		.dout(new_net_17201)
	);

	bfr new_net_17202_bfr_after (
		.din(new_net_17201),
		.dout(new_net_17202)
	);

	bfr new_net_17203_bfr_after (
		.din(new_net_17202),
		.dout(new_net_17203)
	);

	bfr new_net_17204_bfr_after (
		.din(new_net_17203),
		.dout(new_net_17204)
	);

	bfr new_net_17205_bfr_after (
		.din(new_net_17204),
		.dout(new_net_17205)
	);

	bfr new_net_17206_bfr_after (
		.din(new_net_17205),
		.dout(new_net_17206)
	);

	bfr new_net_17207_bfr_after (
		.din(new_net_17206),
		.dout(new_net_17207)
	);

	bfr new_net_17208_bfr_after (
		.din(new_net_17207),
		.dout(new_net_17208)
	);

	bfr new_net_17209_bfr_after (
		.din(new_net_17208),
		.dout(new_net_17209)
	);

	bfr new_net_17210_bfr_after (
		.din(new_net_17209),
		.dout(new_net_17210)
	);

	bfr new_net_17211_bfr_after (
		.din(new_net_17210),
		.dout(new_net_17211)
	);

	bfr new_net_17212_bfr_after (
		.din(new_net_17211),
		.dout(new_net_17212)
	);

	bfr new_net_17213_bfr_after (
		.din(new_net_17212),
		.dout(new_net_17213)
	);

	bfr new_net_17214_bfr_after (
		.din(new_net_17213),
		.dout(new_net_17214)
	);

	bfr new_net_17215_bfr_after (
		.din(new_net_17214),
		.dout(new_net_17215)
	);

	bfr new_net_17216_bfr_after (
		.din(new_net_17215),
		.dout(new_net_17216)
	);

	bfr new_net_17217_bfr_after (
		.din(new_net_17216),
		.dout(new_net_17217)
	);

	bfr new_net_17218_bfr_after (
		.din(new_net_17217),
		.dout(new_net_17218)
	);

	bfr new_net_17219_bfr_after (
		.din(new_net_17218),
		.dout(new_net_17219)
	);

	bfr new_net_17220_bfr_after (
		.din(new_net_17219),
		.dout(new_net_17220)
	);

	bfr new_net_17221_bfr_after (
		.din(new_net_17220),
		.dout(new_net_17221)
	);

	bfr new_net_17222_bfr_after (
		.din(new_net_17221),
		.dout(new_net_17222)
	);

	bfr new_net_17223_bfr_after (
		.din(new_net_17222),
		.dout(new_net_17223)
	);

	bfr new_net_17224_bfr_after (
		.din(new_net_17223),
		.dout(new_net_17224)
	);

	bfr new_net_17225_bfr_after (
		.din(new_net_17224),
		.dout(new_net_17225)
	);

	bfr new_net_17226_bfr_after (
		.din(new_net_17225),
		.dout(new_net_17226)
	);

	bfr new_net_17227_bfr_after (
		.din(new_net_17226),
		.dout(new_net_17227)
	);

	bfr new_net_17228_bfr_after (
		.din(new_net_17227),
		.dout(new_net_17228)
	);

	bfr new_net_17229_bfr_after (
		.din(new_net_17228),
		.dout(new_net_17229)
	);

	bfr new_net_17230_bfr_after (
		.din(new_net_17229),
		.dout(new_net_17230)
	);

	bfr new_net_17231_bfr_after (
		.din(new_net_17230),
		.dout(new_net_17231)
	);

	bfr new_net_17232_bfr_after (
		.din(new_net_17231),
		.dout(new_net_17232)
	);

	bfr new_net_17233_bfr_after (
		.din(new_net_17232),
		.dout(new_net_17233)
	);

	bfr new_net_17234_bfr_after (
		.din(new_net_17233),
		.dout(new_net_17234)
	);

	bfr new_net_17235_bfr_after (
		.din(new_net_17234),
		.dout(new_net_17235)
	);

	bfr new_net_17236_bfr_after (
		.din(new_net_17235),
		.dout(new_net_17236)
	);

	bfr new_net_17237_bfr_after (
		.din(new_net_17236),
		.dout(new_net_17237)
	);

	bfr new_net_17238_bfr_after (
		.din(new_net_17237),
		.dout(new_net_17238)
	);

	bfr new_net_17239_bfr_after (
		.din(new_net_17238),
		.dout(new_net_17239)
	);

	bfr new_net_17240_bfr_after (
		.din(new_net_17239),
		.dout(new_net_17240)
	);

	bfr new_net_17241_bfr_after (
		.din(new_net_17240),
		.dout(new_net_17241)
	);

	bfr new_net_17242_bfr_after (
		.din(new_net_17241),
		.dout(new_net_17242)
	);

	spl2 _0988__v_fanout (
		.a(new_net_17242),
		.b(new_net_1998),
		.c(new_net_1999)
	);

	bfr new_net_17243_bfr_after (
		.din(_1828_),
		.dout(new_net_17243)
	);

	bfr new_net_17244_bfr_after (
		.din(new_net_17243),
		.dout(new_net_17244)
	);

	bfr new_net_17245_bfr_after (
		.din(new_net_17244),
		.dout(new_net_17245)
	);

	bfr new_net_17246_bfr_after (
		.din(new_net_17245),
		.dout(new_net_17246)
	);

	bfr new_net_17247_bfr_after (
		.din(new_net_17246),
		.dout(new_net_17247)
	);

	bfr new_net_17248_bfr_after (
		.din(new_net_17247),
		.dout(new_net_17248)
	);

	bfr new_net_17249_bfr_after (
		.din(new_net_17248),
		.dout(new_net_17249)
	);

	bfr new_net_17250_bfr_after (
		.din(new_net_17249),
		.dout(new_net_17250)
	);

	bfr new_net_17251_bfr_after (
		.din(new_net_17250),
		.dout(new_net_17251)
	);

	bfr new_net_17252_bfr_after (
		.din(new_net_17251),
		.dout(new_net_17252)
	);

	bfr new_net_17253_bfr_after (
		.din(new_net_17252),
		.dout(new_net_17253)
	);

	bfr new_net_17254_bfr_after (
		.din(new_net_17253),
		.dout(new_net_17254)
	);

	bfr new_net_17255_bfr_after (
		.din(new_net_17254),
		.dout(new_net_17255)
	);

	bfr new_net_17256_bfr_after (
		.din(new_net_17255),
		.dout(new_net_17256)
	);

	spl2 _1828__v_fanout (
		.a(new_net_17256),
		.b(new_net_1868),
		.c(new_net_1869)
	);

	bfr new_net_17257_bfr_after (
		.din(_0776_),
		.dout(new_net_17257)
	);

	bfr new_net_17258_bfr_after (
		.din(new_net_17257),
		.dout(new_net_17258)
	);

	bfr new_net_17259_bfr_after (
		.din(new_net_17258),
		.dout(new_net_17259)
	);

	bfr new_net_17260_bfr_after (
		.din(new_net_17259),
		.dout(new_net_17260)
	);

	bfr new_net_17261_bfr_after (
		.din(new_net_17260),
		.dout(new_net_17261)
	);

	bfr new_net_17262_bfr_after (
		.din(new_net_17261),
		.dout(new_net_17262)
	);

	bfr new_net_17263_bfr_after (
		.din(new_net_17262),
		.dout(new_net_17263)
	);

	bfr new_net_17264_bfr_after (
		.din(new_net_17263),
		.dout(new_net_17264)
	);

	bfr new_net_17265_bfr_after (
		.din(new_net_17264),
		.dout(new_net_17265)
	);

	bfr new_net_17266_bfr_after (
		.din(new_net_17265),
		.dout(new_net_17266)
	);

	bfr new_net_17267_bfr_after (
		.din(new_net_17266),
		.dout(new_net_17267)
	);

	bfr new_net_17268_bfr_after (
		.din(new_net_17267),
		.dout(new_net_17268)
	);

	bfr new_net_17269_bfr_after (
		.din(new_net_17268),
		.dout(new_net_17269)
	);

	bfr new_net_17270_bfr_after (
		.din(new_net_17269),
		.dout(new_net_17270)
	);

	bfr new_net_17271_bfr_after (
		.din(new_net_17270),
		.dout(new_net_17271)
	);

	bfr new_net_17272_bfr_after (
		.din(new_net_17271),
		.dout(new_net_17272)
	);

	bfr new_net_17273_bfr_after (
		.din(new_net_17272),
		.dout(new_net_17273)
	);

	bfr new_net_17274_bfr_after (
		.din(new_net_17273),
		.dout(new_net_17274)
	);

	bfr new_net_17275_bfr_after (
		.din(new_net_17274),
		.dout(new_net_17275)
	);

	bfr new_net_17276_bfr_after (
		.din(new_net_17275),
		.dout(new_net_17276)
	);

	bfr new_net_17277_bfr_after (
		.din(new_net_17276),
		.dout(new_net_17277)
	);

	bfr new_net_17278_bfr_after (
		.din(new_net_17277),
		.dout(new_net_17278)
	);

	bfr new_net_17279_bfr_after (
		.din(new_net_17278),
		.dout(new_net_17279)
	);

	bfr new_net_17280_bfr_after (
		.din(new_net_17279),
		.dout(new_net_17280)
	);

	bfr new_net_17281_bfr_after (
		.din(new_net_17280),
		.dout(new_net_17281)
	);

	bfr new_net_17282_bfr_after (
		.din(new_net_17281),
		.dout(new_net_17282)
	);

	bfr new_net_17283_bfr_after (
		.din(new_net_17282),
		.dout(new_net_17283)
	);

	bfr new_net_17284_bfr_after (
		.din(new_net_17283),
		.dout(new_net_17284)
	);

	bfr new_net_17285_bfr_after (
		.din(new_net_17284),
		.dout(new_net_17285)
	);

	bfr new_net_17286_bfr_after (
		.din(new_net_17285),
		.dout(new_net_17286)
	);

	bfr new_net_17287_bfr_after (
		.din(new_net_17286),
		.dout(new_net_17287)
	);

	bfr new_net_17288_bfr_after (
		.din(new_net_17287),
		.dout(new_net_17288)
	);

	bfr new_net_17289_bfr_after (
		.din(new_net_17288),
		.dout(new_net_17289)
	);

	bfr new_net_17290_bfr_after (
		.din(new_net_17289),
		.dout(new_net_17290)
	);

	bfr new_net_17291_bfr_after (
		.din(new_net_17290),
		.dout(new_net_17291)
	);

	bfr new_net_17292_bfr_after (
		.din(new_net_17291),
		.dout(new_net_17292)
	);

	bfr new_net_17293_bfr_after (
		.din(new_net_17292),
		.dout(new_net_17293)
	);

	bfr new_net_17294_bfr_after (
		.din(new_net_17293),
		.dout(new_net_17294)
	);

	bfr new_net_17295_bfr_after (
		.din(new_net_17294),
		.dout(new_net_17295)
	);

	bfr new_net_17296_bfr_after (
		.din(new_net_17295),
		.dout(new_net_17296)
	);

	bfr new_net_17297_bfr_after (
		.din(new_net_17296),
		.dout(new_net_17297)
	);

	bfr new_net_17298_bfr_after (
		.din(new_net_17297),
		.dout(new_net_17298)
	);

	bfr new_net_17299_bfr_after (
		.din(new_net_17298),
		.dout(new_net_17299)
	);

	bfr new_net_17300_bfr_after (
		.din(new_net_17299),
		.dout(new_net_17300)
	);

	bfr new_net_17301_bfr_after (
		.din(new_net_17300),
		.dout(new_net_17301)
	);

	bfr new_net_17302_bfr_after (
		.din(new_net_17301),
		.dout(new_net_17302)
	);

	bfr new_net_17303_bfr_after (
		.din(new_net_17302),
		.dout(new_net_17303)
	);

	bfr new_net_17304_bfr_after (
		.din(new_net_17303),
		.dout(new_net_17304)
	);

	bfr new_net_17305_bfr_after (
		.din(new_net_17304),
		.dout(new_net_17305)
	);

	bfr new_net_17306_bfr_after (
		.din(new_net_17305),
		.dout(new_net_17306)
	);

	bfr new_net_17307_bfr_after (
		.din(new_net_17306),
		.dout(new_net_17307)
	);

	bfr new_net_17308_bfr_after (
		.din(new_net_17307),
		.dout(new_net_17308)
	);

	bfr new_net_17309_bfr_after (
		.din(new_net_17308),
		.dout(new_net_17309)
	);

	bfr new_net_17310_bfr_after (
		.din(new_net_17309),
		.dout(new_net_17310)
	);

	bfr new_net_17311_bfr_after (
		.din(new_net_17310),
		.dout(new_net_17311)
	);

	bfr new_net_17312_bfr_after (
		.din(new_net_17311),
		.dout(new_net_17312)
	);

	bfr new_net_17313_bfr_after (
		.din(new_net_17312),
		.dout(new_net_17313)
	);

	bfr new_net_17314_bfr_after (
		.din(new_net_17313),
		.dout(new_net_17314)
	);

	bfr new_net_17315_bfr_after (
		.din(new_net_17314),
		.dout(new_net_17315)
	);

	bfr new_net_17316_bfr_after (
		.din(new_net_17315),
		.dout(new_net_17316)
	);

	bfr new_net_17317_bfr_after (
		.din(new_net_17316),
		.dout(new_net_17317)
	);

	bfr new_net_17318_bfr_after (
		.din(new_net_17317),
		.dout(new_net_17318)
	);

	bfr new_net_17319_bfr_after (
		.din(new_net_17318),
		.dout(new_net_17319)
	);

	bfr new_net_17320_bfr_after (
		.din(new_net_17319),
		.dout(new_net_17320)
	);

	bfr new_net_17321_bfr_after (
		.din(new_net_17320),
		.dout(new_net_17321)
	);

	bfr new_net_17322_bfr_after (
		.din(new_net_17321),
		.dout(new_net_17322)
	);

	bfr new_net_17323_bfr_after (
		.din(new_net_17322),
		.dout(new_net_17323)
	);

	bfr new_net_17324_bfr_after (
		.din(new_net_17323),
		.dout(new_net_17324)
	);

	bfr new_net_17325_bfr_after (
		.din(new_net_17324),
		.dout(new_net_17325)
	);

	bfr new_net_17326_bfr_after (
		.din(new_net_17325),
		.dout(new_net_17326)
	);

	bfr new_net_17327_bfr_after (
		.din(new_net_17326),
		.dout(new_net_17327)
	);

	bfr new_net_17328_bfr_after (
		.din(new_net_17327),
		.dout(new_net_17328)
	);

	bfr new_net_17329_bfr_after (
		.din(new_net_17328),
		.dout(new_net_17329)
	);

	bfr new_net_17330_bfr_after (
		.din(new_net_17329),
		.dout(new_net_17330)
	);

	bfr new_net_17331_bfr_after (
		.din(new_net_17330),
		.dout(new_net_17331)
	);

	bfr new_net_17332_bfr_after (
		.din(new_net_17331),
		.dout(new_net_17332)
	);

	bfr new_net_17333_bfr_after (
		.din(new_net_17332),
		.dout(new_net_17333)
	);

	bfr new_net_17334_bfr_after (
		.din(new_net_17333),
		.dout(new_net_17334)
	);

	spl2 _0776__v_fanout (
		.a(new_net_17334),
		.b(new_net_1888),
		.c(new_net_1889)
	);

	bfr new_net_17335_bfr_after (
		.din(_1371_),
		.dout(new_net_17335)
	);

	bfr new_net_17336_bfr_after (
		.din(new_net_17335),
		.dout(new_net_17336)
	);

	bfr new_net_17337_bfr_after (
		.din(new_net_17336),
		.dout(new_net_17337)
	);

	bfr new_net_17338_bfr_after (
		.din(new_net_17337),
		.dout(new_net_17338)
	);

	bfr new_net_17339_bfr_after (
		.din(new_net_17338),
		.dout(new_net_17339)
	);

	bfr new_net_17340_bfr_after (
		.din(new_net_17339),
		.dout(new_net_17340)
	);

	bfr new_net_17341_bfr_after (
		.din(new_net_17340),
		.dout(new_net_17341)
	);

	bfr new_net_17342_bfr_after (
		.din(new_net_17341),
		.dout(new_net_17342)
	);

	bfr new_net_17343_bfr_after (
		.din(new_net_17342),
		.dout(new_net_17343)
	);

	bfr new_net_17344_bfr_after (
		.din(new_net_17343),
		.dout(new_net_17344)
	);

	bfr new_net_17345_bfr_after (
		.din(new_net_17344),
		.dout(new_net_17345)
	);

	bfr new_net_17346_bfr_after (
		.din(new_net_17345),
		.dout(new_net_17346)
	);

	bfr new_net_17347_bfr_after (
		.din(new_net_17346),
		.dout(new_net_17347)
	);

	bfr new_net_17348_bfr_after (
		.din(new_net_17347),
		.dout(new_net_17348)
	);

	bfr new_net_17349_bfr_after (
		.din(new_net_17348),
		.dout(new_net_17349)
	);

	bfr new_net_17350_bfr_after (
		.din(new_net_17349),
		.dout(new_net_17350)
	);

	bfr new_net_17351_bfr_after (
		.din(new_net_17350),
		.dout(new_net_17351)
	);

	bfr new_net_17352_bfr_after (
		.din(new_net_17351),
		.dout(new_net_17352)
	);

	bfr new_net_17353_bfr_after (
		.din(new_net_17352),
		.dout(new_net_17353)
	);

	bfr new_net_17354_bfr_after (
		.din(new_net_17353),
		.dout(new_net_17354)
	);

	bfr new_net_17355_bfr_after (
		.din(new_net_17354),
		.dout(new_net_17355)
	);

	bfr new_net_17356_bfr_after (
		.din(new_net_17355),
		.dout(new_net_17356)
	);

	bfr new_net_17357_bfr_after (
		.din(new_net_17356),
		.dout(new_net_17357)
	);

	bfr new_net_17358_bfr_after (
		.din(new_net_17357),
		.dout(new_net_17358)
	);

	bfr new_net_17359_bfr_after (
		.din(new_net_17358),
		.dout(new_net_17359)
	);

	bfr new_net_17360_bfr_after (
		.din(new_net_17359),
		.dout(new_net_17360)
	);

	bfr new_net_17361_bfr_after (
		.din(new_net_17360),
		.dout(new_net_17361)
	);

	bfr new_net_17362_bfr_after (
		.din(new_net_17361),
		.dout(new_net_17362)
	);

	bfr new_net_17363_bfr_after (
		.din(new_net_17362),
		.dout(new_net_17363)
	);

	bfr new_net_17364_bfr_after (
		.din(new_net_17363),
		.dout(new_net_17364)
	);

	bfr new_net_17365_bfr_after (
		.din(new_net_17364),
		.dout(new_net_17365)
	);

	bfr new_net_17366_bfr_after (
		.din(new_net_17365),
		.dout(new_net_17366)
	);

	bfr new_net_17367_bfr_after (
		.din(new_net_17366),
		.dout(new_net_17367)
	);

	bfr new_net_17368_bfr_after (
		.din(new_net_17367),
		.dout(new_net_17368)
	);

	bfr new_net_17369_bfr_after (
		.din(new_net_17368),
		.dout(new_net_17369)
	);

	bfr new_net_17370_bfr_after (
		.din(new_net_17369),
		.dout(new_net_17370)
	);

	bfr new_net_17371_bfr_after (
		.din(new_net_17370),
		.dout(new_net_17371)
	);

	bfr new_net_17372_bfr_after (
		.din(new_net_17371),
		.dout(new_net_17372)
	);

	bfr new_net_17373_bfr_after (
		.din(new_net_17372),
		.dout(new_net_17373)
	);

	bfr new_net_17374_bfr_after (
		.din(new_net_17373),
		.dout(new_net_17374)
	);

	bfr new_net_17375_bfr_after (
		.din(new_net_17374),
		.dout(new_net_17375)
	);

	bfr new_net_17376_bfr_after (
		.din(new_net_17375),
		.dout(new_net_17376)
	);

	bfr new_net_17377_bfr_after (
		.din(new_net_17376),
		.dout(new_net_17377)
	);

	bfr new_net_17378_bfr_after (
		.din(new_net_17377),
		.dout(new_net_17378)
	);

	bfr new_net_17379_bfr_after (
		.din(new_net_17378),
		.dout(new_net_17379)
	);

	bfr new_net_17380_bfr_after (
		.din(new_net_17379),
		.dout(new_net_17380)
	);

	bfr new_net_17381_bfr_after (
		.din(new_net_17380),
		.dout(new_net_17381)
	);

	bfr new_net_17382_bfr_after (
		.din(new_net_17381),
		.dout(new_net_17382)
	);

	spl2 _1371__v_fanout (
		.a(new_net_17382),
		.b(new_net_2076),
		.c(new_net_2077)
	);

	bfr new_net_17383_bfr_after (
		.din(_1452_),
		.dout(new_net_17383)
	);

	bfr new_net_17384_bfr_after (
		.din(new_net_17383),
		.dout(new_net_17384)
	);

	bfr new_net_17385_bfr_after (
		.din(new_net_17384),
		.dout(new_net_17385)
	);

	bfr new_net_17386_bfr_after (
		.din(new_net_17385),
		.dout(new_net_17386)
	);

	bfr new_net_17387_bfr_after (
		.din(new_net_17386),
		.dout(new_net_17387)
	);

	bfr new_net_17388_bfr_after (
		.din(new_net_17387),
		.dout(new_net_17388)
	);

	bfr new_net_17389_bfr_after (
		.din(new_net_17388),
		.dout(new_net_17389)
	);

	bfr new_net_17390_bfr_after (
		.din(new_net_17389),
		.dout(new_net_17390)
	);

	bfr new_net_17391_bfr_after (
		.din(new_net_17390),
		.dout(new_net_17391)
	);

	bfr new_net_17392_bfr_after (
		.din(new_net_17391),
		.dout(new_net_17392)
	);

	bfr new_net_17393_bfr_after (
		.din(new_net_17392),
		.dout(new_net_17393)
	);

	bfr new_net_17394_bfr_after (
		.din(new_net_17393),
		.dout(new_net_17394)
	);

	bfr new_net_17395_bfr_after (
		.din(new_net_17394),
		.dout(new_net_17395)
	);

	bfr new_net_17396_bfr_after (
		.din(new_net_17395),
		.dout(new_net_17396)
	);

	bfr new_net_17397_bfr_after (
		.din(new_net_17396),
		.dout(new_net_17397)
	);

	bfr new_net_17398_bfr_after (
		.din(new_net_17397),
		.dout(new_net_17398)
	);

	bfr new_net_17399_bfr_after (
		.din(new_net_17398),
		.dout(new_net_17399)
	);

	bfr new_net_17400_bfr_after (
		.din(new_net_17399),
		.dout(new_net_17400)
	);

	bfr new_net_17401_bfr_after (
		.din(new_net_17400),
		.dout(new_net_17401)
	);

	bfr new_net_17402_bfr_after (
		.din(new_net_17401),
		.dout(new_net_17402)
	);

	bfr new_net_17403_bfr_after (
		.din(new_net_17402),
		.dout(new_net_17403)
	);

	bfr new_net_17404_bfr_after (
		.din(new_net_17403),
		.dout(new_net_17404)
	);

	bfr new_net_17405_bfr_after (
		.din(new_net_17404),
		.dout(new_net_17405)
	);

	bfr new_net_17406_bfr_after (
		.din(new_net_17405),
		.dout(new_net_17406)
	);

	bfr new_net_17407_bfr_after (
		.din(new_net_17406),
		.dout(new_net_17407)
	);

	bfr new_net_17408_bfr_after (
		.din(new_net_17407),
		.dout(new_net_17408)
	);

	bfr new_net_17409_bfr_after (
		.din(new_net_17408),
		.dout(new_net_17409)
	);

	bfr new_net_17410_bfr_after (
		.din(new_net_17409),
		.dout(new_net_17410)
	);

	bfr new_net_17411_bfr_after (
		.din(new_net_17410),
		.dout(new_net_17411)
	);

	bfr new_net_17412_bfr_after (
		.din(new_net_17411),
		.dout(new_net_17412)
	);

	bfr new_net_17413_bfr_after (
		.din(new_net_17412),
		.dout(new_net_17413)
	);

	bfr new_net_17414_bfr_after (
		.din(new_net_17413),
		.dout(new_net_17414)
	);

	bfr new_net_17415_bfr_after (
		.din(new_net_17414),
		.dout(new_net_17415)
	);

	bfr new_net_17416_bfr_after (
		.din(new_net_17415),
		.dout(new_net_17416)
	);

	bfr new_net_17417_bfr_after (
		.din(new_net_17416),
		.dout(new_net_17417)
	);

	bfr new_net_17418_bfr_after (
		.din(new_net_17417),
		.dout(new_net_17418)
	);

	bfr new_net_17419_bfr_after (
		.din(new_net_17418),
		.dout(new_net_17419)
	);

	bfr new_net_17420_bfr_after (
		.din(new_net_17419),
		.dout(new_net_17420)
	);

	bfr new_net_17421_bfr_after (
		.din(new_net_17420),
		.dout(new_net_17421)
	);

	bfr new_net_17422_bfr_after (
		.din(new_net_17421),
		.dout(new_net_17422)
	);

	bfr new_net_17423_bfr_after (
		.din(new_net_17422),
		.dout(new_net_17423)
	);

	bfr new_net_17424_bfr_after (
		.din(new_net_17423),
		.dout(new_net_17424)
	);

	bfr new_net_17425_bfr_after (
		.din(new_net_17424),
		.dout(new_net_17425)
	);

	bfr new_net_17426_bfr_after (
		.din(new_net_17425),
		.dout(new_net_17426)
	);

	bfr new_net_17427_bfr_after (
		.din(new_net_17426),
		.dout(new_net_17427)
	);

	bfr new_net_17428_bfr_after (
		.din(new_net_17427),
		.dout(new_net_17428)
	);

	bfr new_net_17429_bfr_after (
		.din(new_net_17428),
		.dout(new_net_17429)
	);

	bfr new_net_17430_bfr_after (
		.din(new_net_17429),
		.dout(new_net_17430)
	);

	bfr new_net_17431_bfr_after (
		.din(new_net_17430),
		.dout(new_net_17431)
	);

	bfr new_net_17432_bfr_after (
		.din(new_net_17431),
		.dout(new_net_17432)
	);

	bfr new_net_17433_bfr_after (
		.din(new_net_17432),
		.dout(new_net_17433)
	);

	bfr new_net_17434_bfr_after (
		.din(new_net_17433),
		.dout(new_net_17434)
	);

	bfr new_net_17435_bfr_after (
		.din(new_net_17434),
		.dout(new_net_17435)
	);

	bfr new_net_17436_bfr_after (
		.din(new_net_17435),
		.dout(new_net_17436)
	);

	bfr new_net_17437_bfr_after (
		.din(new_net_17436),
		.dout(new_net_17437)
	);

	bfr new_net_17438_bfr_after (
		.din(new_net_17437),
		.dout(new_net_17438)
	);

	bfr new_net_17439_bfr_after (
		.din(new_net_17438),
		.dout(new_net_17439)
	);

	bfr new_net_17440_bfr_after (
		.din(new_net_17439),
		.dout(new_net_17440)
	);

	bfr new_net_17441_bfr_after (
		.din(new_net_17440),
		.dout(new_net_17441)
	);

	bfr new_net_17442_bfr_after (
		.din(new_net_17441),
		.dout(new_net_17442)
	);

	bfr new_net_17443_bfr_after (
		.din(new_net_17442),
		.dout(new_net_17443)
	);

	bfr new_net_17444_bfr_after (
		.din(new_net_17443),
		.dout(new_net_17444)
	);

	bfr new_net_17445_bfr_after (
		.din(new_net_17444),
		.dout(new_net_17445)
	);

	bfr new_net_17446_bfr_after (
		.din(new_net_17445),
		.dout(new_net_17446)
	);

	bfr new_net_17447_bfr_after (
		.din(new_net_17446),
		.dout(new_net_17447)
	);

	bfr new_net_17448_bfr_after (
		.din(new_net_17447),
		.dout(new_net_17448)
	);

	bfr new_net_17449_bfr_after (
		.din(new_net_17448),
		.dout(new_net_17449)
	);

	bfr new_net_17450_bfr_after (
		.din(new_net_17449),
		.dout(new_net_17450)
	);

	bfr new_net_17451_bfr_after (
		.din(new_net_17450),
		.dout(new_net_17451)
	);

	bfr new_net_17452_bfr_after (
		.din(new_net_17451),
		.dout(new_net_17452)
	);

	bfr new_net_17453_bfr_after (
		.din(new_net_17452),
		.dout(new_net_17453)
	);

	bfr new_net_17454_bfr_after (
		.din(new_net_17453),
		.dout(new_net_17454)
	);

	bfr new_net_17455_bfr_after (
		.din(new_net_17454),
		.dout(new_net_17455)
	);

	bfr new_net_17456_bfr_after (
		.din(new_net_17455),
		.dout(new_net_17456)
	);

	bfr new_net_17457_bfr_after (
		.din(new_net_17456),
		.dout(new_net_17457)
	);

	bfr new_net_17458_bfr_after (
		.din(new_net_17457),
		.dout(new_net_17458)
	);

	bfr new_net_17459_bfr_after (
		.din(new_net_17458),
		.dout(new_net_17459)
	);

	bfr new_net_17460_bfr_after (
		.din(new_net_17459),
		.dout(new_net_17460)
	);

	bfr new_net_17461_bfr_after (
		.din(new_net_17460),
		.dout(new_net_17461)
	);

	bfr new_net_17462_bfr_after (
		.din(new_net_17461),
		.dout(new_net_17462)
	);

	bfr new_net_17463_bfr_after (
		.din(new_net_17462),
		.dout(new_net_17463)
	);

	bfr new_net_17464_bfr_after (
		.din(new_net_17463),
		.dout(new_net_17464)
	);

	bfr new_net_17465_bfr_after (
		.din(new_net_17464),
		.dout(new_net_17465)
	);

	bfr new_net_17466_bfr_after (
		.din(new_net_17465),
		.dout(new_net_17466)
	);

	bfr new_net_17467_bfr_after (
		.din(new_net_17466),
		.dout(new_net_17467)
	);

	bfr new_net_17468_bfr_after (
		.din(new_net_17467),
		.dout(new_net_17468)
	);

	bfr new_net_17469_bfr_after (
		.din(new_net_17468),
		.dout(new_net_17469)
	);

	bfr new_net_17470_bfr_after (
		.din(new_net_17469),
		.dout(new_net_17470)
	);

	bfr new_net_17471_bfr_after (
		.din(new_net_17470),
		.dout(new_net_17471)
	);

	bfr new_net_17472_bfr_after (
		.din(new_net_17471),
		.dout(new_net_17472)
	);

	bfr new_net_17473_bfr_after (
		.din(new_net_17472),
		.dout(new_net_17473)
	);

	bfr new_net_17474_bfr_after (
		.din(new_net_17473),
		.dout(new_net_17474)
	);

	bfr new_net_17475_bfr_after (
		.din(new_net_17474),
		.dout(new_net_17475)
	);

	bfr new_net_17476_bfr_after (
		.din(new_net_17475),
		.dout(new_net_17476)
	);

	bfr new_net_17477_bfr_after (
		.din(new_net_17476),
		.dout(new_net_17477)
	);

	bfr new_net_17478_bfr_after (
		.din(new_net_17477),
		.dout(new_net_17478)
	);

	spl2 _1452__v_fanout (
		.a(new_net_17478),
		.b(new_net_1493),
		.c(new_net_1494)
	);

	bfr new_net_17479_bfr_after (
		.din(_0329_),
		.dout(new_net_17479)
	);

	bfr new_net_17480_bfr_after (
		.din(new_net_17479),
		.dout(new_net_17480)
	);

	bfr new_net_17481_bfr_after (
		.din(new_net_17480),
		.dout(new_net_17481)
	);

	bfr new_net_17482_bfr_after (
		.din(new_net_17481),
		.dout(new_net_17482)
	);

	bfr new_net_17483_bfr_after (
		.din(new_net_17482),
		.dout(new_net_17483)
	);

	bfr new_net_17484_bfr_after (
		.din(new_net_17483),
		.dout(new_net_17484)
	);

	bfr new_net_17485_bfr_after (
		.din(new_net_17484),
		.dout(new_net_17485)
	);

	bfr new_net_17486_bfr_after (
		.din(new_net_17485),
		.dout(new_net_17486)
	);

	bfr new_net_17487_bfr_after (
		.din(new_net_17486),
		.dout(new_net_17487)
	);

	bfr new_net_17488_bfr_after (
		.din(new_net_17487),
		.dout(new_net_17488)
	);

	bfr new_net_17489_bfr_after (
		.din(new_net_17488),
		.dout(new_net_17489)
	);

	bfr new_net_17490_bfr_after (
		.din(new_net_17489),
		.dout(new_net_17490)
	);

	bfr new_net_17491_bfr_after (
		.din(new_net_17490),
		.dout(new_net_17491)
	);

	bfr new_net_17492_bfr_after (
		.din(new_net_17491),
		.dout(new_net_17492)
	);

	bfr new_net_17493_bfr_after (
		.din(new_net_17492),
		.dout(new_net_17493)
	);

	bfr new_net_17494_bfr_after (
		.din(new_net_17493),
		.dout(new_net_17494)
	);

	bfr new_net_17495_bfr_after (
		.din(new_net_17494),
		.dout(new_net_17495)
	);

	bfr new_net_17496_bfr_after (
		.din(new_net_17495),
		.dout(new_net_17496)
	);

	bfr new_net_17497_bfr_after (
		.din(new_net_17496),
		.dout(new_net_17497)
	);

	bfr new_net_17498_bfr_after (
		.din(new_net_17497),
		.dout(new_net_17498)
	);

	bfr new_net_17499_bfr_after (
		.din(new_net_17498),
		.dout(new_net_17499)
	);

	bfr new_net_17500_bfr_after (
		.din(new_net_17499),
		.dout(new_net_17500)
	);

	bfr new_net_17501_bfr_after (
		.din(new_net_17500),
		.dout(new_net_17501)
	);

	bfr new_net_17502_bfr_after (
		.din(new_net_17501),
		.dout(new_net_17502)
	);

	bfr new_net_17503_bfr_after (
		.din(new_net_17502),
		.dout(new_net_17503)
	);

	bfr new_net_17504_bfr_after (
		.din(new_net_17503),
		.dout(new_net_17504)
	);

	bfr new_net_17505_bfr_after (
		.din(new_net_17504),
		.dout(new_net_17505)
	);

	bfr new_net_17506_bfr_after (
		.din(new_net_17505),
		.dout(new_net_17506)
	);

	bfr new_net_17507_bfr_after (
		.din(new_net_17506),
		.dout(new_net_17507)
	);

	bfr new_net_17508_bfr_after (
		.din(new_net_17507),
		.dout(new_net_17508)
	);

	bfr new_net_17509_bfr_after (
		.din(new_net_17508),
		.dout(new_net_17509)
	);

	bfr new_net_17510_bfr_after (
		.din(new_net_17509),
		.dout(new_net_17510)
	);

	bfr new_net_17511_bfr_after (
		.din(new_net_17510),
		.dout(new_net_17511)
	);

	bfr new_net_17512_bfr_after (
		.din(new_net_17511),
		.dout(new_net_17512)
	);

	bfr new_net_17513_bfr_after (
		.din(new_net_17512),
		.dout(new_net_17513)
	);

	bfr new_net_17514_bfr_after (
		.din(new_net_17513),
		.dout(new_net_17514)
	);

	bfr new_net_17515_bfr_after (
		.din(new_net_17514),
		.dout(new_net_17515)
	);

	bfr new_net_17516_bfr_after (
		.din(new_net_17515),
		.dout(new_net_17516)
	);

	bfr new_net_17517_bfr_after (
		.din(new_net_17516),
		.dout(new_net_17517)
	);

	bfr new_net_17518_bfr_after (
		.din(new_net_17517),
		.dout(new_net_17518)
	);

	bfr new_net_17519_bfr_after (
		.din(new_net_17518),
		.dout(new_net_17519)
	);

	bfr new_net_17520_bfr_after (
		.din(new_net_17519),
		.dout(new_net_17520)
	);

	bfr new_net_17521_bfr_after (
		.din(new_net_17520),
		.dout(new_net_17521)
	);

	bfr new_net_17522_bfr_after (
		.din(new_net_17521),
		.dout(new_net_17522)
	);

	bfr new_net_17523_bfr_after (
		.din(new_net_17522),
		.dout(new_net_17523)
	);

	bfr new_net_17524_bfr_after (
		.din(new_net_17523),
		.dout(new_net_17524)
	);

	bfr new_net_17525_bfr_after (
		.din(new_net_17524),
		.dout(new_net_17525)
	);

	bfr new_net_17526_bfr_after (
		.din(new_net_17525),
		.dout(new_net_17526)
	);

	bfr new_net_17527_bfr_after (
		.din(new_net_17526),
		.dout(new_net_17527)
	);

	bfr new_net_17528_bfr_after (
		.din(new_net_17527),
		.dout(new_net_17528)
	);

	bfr new_net_17529_bfr_after (
		.din(new_net_17528),
		.dout(new_net_17529)
	);

	bfr new_net_17530_bfr_after (
		.din(new_net_17529),
		.dout(new_net_17530)
	);

	bfr new_net_17531_bfr_after (
		.din(new_net_17530),
		.dout(new_net_17531)
	);

	bfr new_net_17532_bfr_after (
		.din(new_net_17531),
		.dout(new_net_17532)
	);

	bfr new_net_17533_bfr_after (
		.din(new_net_17532),
		.dout(new_net_17533)
	);

	bfr new_net_17534_bfr_after (
		.din(new_net_17533),
		.dout(new_net_17534)
	);

	bfr new_net_17535_bfr_after (
		.din(new_net_17534),
		.dout(new_net_17535)
	);

	bfr new_net_17536_bfr_after (
		.din(new_net_17535),
		.dout(new_net_17536)
	);

	bfr new_net_17537_bfr_after (
		.din(new_net_17536),
		.dout(new_net_17537)
	);

	bfr new_net_17538_bfr_after (
		.din(new_net_17537),
		.dout(new_net_17538)
	);

	bfr new_net_17539_bfr_after (
		.din(new_net_17538),
		.dout(new_net_17539)
	);

	bfr new_net_17540_bfr_after (
		.din(new_net_17539),
		.dout(new_net_17540)
	);

	bfr new_net_17541_bfr_after (
		.din(new_net_17540),
		.dout(new_net_17541)
	);

	bfr new_net_17542_bfr_after (
		.din(new_net_17541),
		.dout(new_net_17542)
	);

	bfr new_net_17543_bfr_after (
		.din(new_net_17542),
		.dout(new_net_17543)
	);

	bfr new_net_17544_bfr_after (
		.din(new_net_17543),
		.dout(new_net_17544)
	);

	bfr new_net_17545_bfr_after (
		.din(new_net_17544),
		.dout(new_net_17545)
	);

	bfr new_net_17546_bfr_after (
		.din(new_net_17545),
		.dout(new_net_17546)
	);

	bfr new_net_17547_bfr_after (
		.din(new_net_17546),
		.dout(new_net_17547)
	);

	bfr new_net_17548_bfr_after (
		.din(new_net_17547),
		.dout(new_net_17548)
	);

	bfr new_net_17549_bfr_after (
		.din(new_net_17548),
		.dout(new_net_17549)
	);

	bfr new_net_17550_bfr_after (
		.din(new_net_17549),
		.dout(new_net_17550)
	);

	bfr new_net_17551_bfr_after (
		.din(new_net_17550),
		.dout(new_net_17551)
	);

	bfr new_net_17552_bfr_after (
		.din(new_net_17551),
		.dout(new_net_17552)
	);

	bfr new_net_17553_bfr_after (
		.din(new_net_17552),
		.dout(new_net_17553)
	);

	bfr new_net_17554_bfr_after (
		.din(new_net_17553),
		.dout(new_net_17554)
	);

	bfr new_net_17555_bfr_after (
		.din(new_net_17554),
		.dout(new_net_17555)
	);

	bfr new_net_17556_bfr_after (
		.din(new_net_17555),
		.dout(new_net_17556)
	);

	bfr new_net_17557_bfr_after (
		.din(new_net_17556),
		.dout(new_net_17557)
	);

	bfr new_net_17558_bfr_after (
		.din(new_net_17557),
		.dout(new_net_17558)
	);

	bfr new_net_17559_bfr_after (
		.din(new_net_17558),
		.dout(new_net_17559)
	);

	bfr new_net_17560_bfr_after (
		.din(new_net_17559),
		.dout(new_net_17560)
	);

	bfr new_net_17561_bfr_after (
		.din(new_net_17560),
		.dout(new_net_17561)
	);

	bfr new_net_17562_bfr_after (
		.din(new_net_17561),
		.dout(new_net_17562)
	);

	bfr new_net_17563_bfr_after (
		.din(new_net_17562),
		.dout(new_net_17563)
	);

	bfr new_net_17564_bfr_after (
		.din(new_net_17563),
		.dout(new_net_17564)
	);

	bfr new_net_17565_bfr_after (
		.din(new_net_17564),
		.dout(new_net_17565)
	);

	bfr new_net_17566_bfr_after (
		.din(new_net_17565),
		.dout(new_net_17566)
	);

	bfr new_net_17567_bfr_after (
		.din(new_net_17566),
		.dout(new_net_17567)
	);

	bfr new_net_17568_bfr_after (
		.din(new_net_17567),
		.dout(new_net_17568)
	);

	bfr new_net_17569_bfr_after (
		.din(new_net_17568),
		.dout(new_net_17569)
	);

	bfr new_net_17570_bfr_after (
		.din(new_net_17569),
		.dout(new_net_17570)
	);

	bfr new_net_17571_bfr_after (
		.din(new_net_17570),
		.dout(new_net_17571)
	);

	bfr new_net_17572_bfr_after (
		.din(new_net_17571),
		.dout(new_net_17572)
	);

	bfr new_net_17573_bfr_after (
		.din(new_net_17572),
		.dout(new_net_17573)
	);

	bfr new_net_17574_bfr_after (
		.din(new_net_17573),
		.dout(new_net_17574)
	);

	bfr new_net_17575_bfr_after (
		.din(new_net_17574),
		.dout(new_net_17575)
	);

	bfr new_net_17576_bfr_after (
		.din(new_net_17575),
		.dout(new_net_17576)
	);

	bfr new_net_17577_bfr_after (
		.din(new_net_17576),
		.dout(new_net_17577)
	);

	bfr new_net_17578_bfr_after (
		.din(new_net_17577),
		.dout(new_net_17578)
	);

	bfr new_net_17579_bfr_after (
		.din(new_net_17578),
		.dout(new_net_17579)
	);

	bfr new_net_17580_bfr_after (
		.din(new_net_17579),
		.dout(new_net_17580)
	);

	bfr new_net_17581_bfr_after (
		.din(new_net_17580),
		.dout(new_net_17581)
	);

	bfr new_net_17582_bfr_after (
		.din(new_net_17581),
		.dout(new_net_17582)
	);

	spl2 _0329__v_fanout (
		.a(new_net_17582),
		.b(new_net_2327),
		.c(new_net_2328)
	);

	bfr new_net_17583_bfr_after (
		.din(_1706_),
		.dout(new_net_17583)
	);

	bfr new_net_17584_bfr_after (
		.din(new_net_17583),
		.dout(new_net_17584)
	);

	bfr new_net_17585_bfr_after (
		.din(new_net_17584),
		.dout(new_net_17585)
	);

	bfr new_net_17586_bfr_after (
		.din(new_net_17585),
		.dout(new_net_17586)
	);

	bfr new_net_17587_bfr_after (
		.din(new_net_17586),
		.dout(new_net_17587)
	);

	bfr new_net_17588_bfr_after (
		.din(new_net_17587),
		.dout(new_net_17588)
	);

	spl2 _1706__v_fanout (
		.a(new_net_17588),
		.b(new_net_2022),
		.c(new_net_2023)
	);

	bfr new_net_17589_bfr_after (
		.din(_0711_),
		.dout(new_net_17589)
	);

	bfr new_net_17590_bfr_after (
		.din(new_net_17589),
		.dout(new_net_17590)
	);

	bfr new_net_17591_bfr_after (
		.din(new_net_17590),
		.dout(new_net_17591)
	);

	bfr new_net_17592_bfr_after (
		.din(new_net_17591),
		.dout(new_net_17592)
	);

	bfr new_net_17593_bfr_after (
		.din(new_net_17592),
		.dout(new_net_17593)
	);

	bfr new_net_17594_bfr_after (
		.din(new_net_17593),
		.dout(new_net_17594)
	);

	bfr new_net_17595_bfr_after (
		.din(new_net_17594),
		.dout(new_net_17595)
	);

	bfr new_net_17596_bfr_after (
		.din(new_net_17595),
		.dout(new_net_17596)
	);

	bfr new_net_17597_bfr_after (
		.din(new_net_17596),
		.dout(new_net_17597)
	);

	bfr new_net_17598_bfr_after (
		.din(new_net_17597),
		.dout(new_net_17598)
	);

	bfr new_net_17599_bfr_after (
		.din(new_net_17598),
		.dout(new_net_17599)
	);

	bfr new_net_17600_bfr_after (
		.din(new_net_17599),
		.dout(new_net_17600)
	);

	bfr new_net_17601_bfr_after (
		.din(new_net_17600),
		.dout(new_net_17601)
	);

	bfr new_net_17602_bfr_after (
		.din(new_net_17601),
		.dout(new_net_17602)
	);

	bfr new_net_17603_bfr_after (
		.din(new_net_17602),
		.dout(new_net_17603)
	);

	bfr new_net_17604_bfr_after (
		.din(new_net_17603),
		.dout(new_net_17604)
	);

	bfr new_net_17605_bfr_after (
		.din(new_net_17604),
		.dout(new_net_17605)
	);

	bfr new_net_17606_bfr_after (
		.din(new_net_17605),
		.dout(new_net_17606)
	);

	bfr new_net_17607_bfr_after (
		.din(new_net_17606),
		.dout(new_net_17607)
	);

	bfr new_net_17608_bfr_after (
		.din(new_net_17607),
		.dout(new_net_17608)
	);

	bfr new_net_17609_bfr_after (
		.din(new_net_17608),
		.dout(new_net_17609)
	);

	bfr new_net_17610_bfr_after (
		.din(new_net_17609),
		.dout(new_net_17610)
	);

	bfr new_net_17611_bfr_after (
		.din(new_net_17610),
		.dout(new_net_17611)
	);

	bfr new_net_17612_bfr_after (
		.din(new_net_17611),
		.dout(new_net_17612)
	);

	bfr new_net_17613_bfr_after (
		.din(new_net_17612),
		.dout(new_net_17613)
	);

	bfr new_net_17614_bfr_after (
		.din(new_net_17613),
		.dout(new_net_17614)
	);

	bfr new_net_17615_bfr_after (
		.din(new_net_17614),
		.dout(new_net_17615)
	);

	bfr new_net_17616_bfr_after (
		.din(new_net_17615),
		.dout(new_net_17616)
	);

	bfr new_net_17617_bfr_after (
		.din(new_net_17616),
		.dout(new_net_17617)
	);

	bfr new_net_17618_bfr_after (
		.din(new_net_17617),
		.dout(new_net_17618)
	);

	bfr new_net_17619_bfr_after (
		.din(new_net_17618),
		.dout(new_net_17619)
	);

	bfr new_net_17620_bfr_after (
		.din(new_net_17619),
		.dout(new_net_17620)
	);

	bfr new_net_17621_bfr_after (
		.din(new_net_17620),
		.dout(new_net_17621)
	);

	bfr new_net_17622_bfr_after (
		.din(new_net_17621),
		.dout(new_net_17622)
	);

	bfr new_net_17623_bfr_after (
		.din(new_net_17622),
		.dout(new_net_17623)
	);

	bfr new_net_17624_bfr_after (
		.din(new_net_17623),
		.dout(new_net_17624)
	);

	bfr new_net_17625_bfr_after (
		.din(new_net_17624),
		.dout(new_net_17625)
	);

	bfr new_net_17626_bfr_after (
		.din(new_net_17625),
		.dout(new_net_17626)
	);

	bfr new_net_17627_bfr_after (
		.din(new_net_17626),
		.dout(new_net_17627)
	);

	bfr new_net_17628_bfr_after (
		.din(new_net_17627),
		.dout(new_net_17628)
	);

	bfr new_net_17629_bfr_after (
		.din(new_net_17628),
		.dout(new_net_17629)
	);

	bfr new_net_17630_bfr_after (
		.din(new_net_17629),
		.dout(new_net_17630)
	);

	bfr new_net_17631_bfr_after (
		.din(new_net_17630),
		.dout(new_net_17631)
	);

	bfr new_net_17632_bfr_after (
		.din(new_net_17631),
		.dout(new_net_17632)
	);

	bfr new_net_17633_bfr_after (
		.din(new_net_17632),
		.dout(new_net_17633)
	);

	bfr new_net_17634_bfr_after (
		.din(new_net_17633),
		.dout(new_net_17634)
	);

	bfr new_net_17635_bfr_after (
		.din(new_net_17634),
		.dout(new_net_17635)
	);

	bfr new_net_17636_bfr_after (
		.din(new_net_17635),
		.dout(new_net_17636)
	);

	bfr new_net_17637_bfr_after (
		.din(new_net_17636),
		.dout(new_net_17637)
	);

	bfr new_net_17638_bfr_after (
		.din(new_net_17637),
		.dout(new_net_17638)
	);

	bfr new_net_17639_bfr_after (
		.din(new_net_17638),
		.dout(new_net_17639)
	);

	bfr new_net_17640_bfr_after (
		.din(new_net_17639),
		.dout(new_net_17640)
	);

	bfr new_net_17641_bfr_after (
		.din(new_net_17640),
		.dout(new_net_17641)
	);

	bfr new_net_17642_bfr_after (
		.din(new_net_17641),
		.dout(new_net_17642)
	);

	spl2 _0711__v_fanout (
		.a(new_net_17642),
		.b(new_net_974),
		.c(new_net_975)
	);

	bfr new_net_17643_bfr_after (
		.din(_0829_),
		.dout(new_net_17643)
	);

	bfr new_net_17644_bfr_after (
		.din(new_net_17643),
		.dout(new_net_17644)
	);

	bfr new_net_17645_bfr_after (
		.din(new_net_17644),
		.dout(new_net_17645)
	);

	bfr new_net_17646_bfr_after (
		.din(new_net_17645),
		.dout(new_net_17646)
	);

	bfr new_net_17647_bfr_after (
		.din(new_net_17646),
		.dout(new_net_17647)
	);

	bfr new_net_17648_bfr_after (
		.din(new_net_17647),
		.dout(new_net_17648)
	);

	bfr new_net_17649_bfr_after (
		.din(new_net_17648),
		.dout(new_net_17649)
	);

	bfr new_net_17650_bfr_after (
		.din(new_net_17649),
		.dout(new_net_17650)
	);

	bfr new_net_17651_bfr_after (
		.din(new_net_17650),
		.dout(new_net_17651)
	);

	bfr new_net_17652_bfr_after (
		.din(new_net_17651),
		.dout(new_net_17652)
	);

	bfr new_net_17653_bfr_after (
		.din(new_net_17652),
		.dout(new_net_17653)
	);

	bfr new_net_17654_bfr_after (
		.din(new_net_17653),
		.dout(new_net_17654)
	);

	bfr new_net_17655_bfr_after (
		.din(new_net_17654),
		.dout(new_net_17655)
	);

	bfr new_net_17656_bfr_after (
		.din(new_net_17655),
		.dout(new_net_17656)
	);

	bfr new_net_17657_bfr_after (
		.din(new_net_17656),
		.dout(new_net_17657)
	);

	bfr new_net_17658_bfr_after (
		.din(new_net_17657),
		.dout(new_net_17658)
	);

	bfr new_net_17659_bfr_after (
		.din(new_net_17658),
		.dout(new_net_17659)
	);

	bfr new_net_17660_bfr_after (
		.din(new_net_17659),
		.dout(new_net_17660)
	);

	bfr new_net_17661_bfr_after (
		.din(new_net_17660),
		.dout(new_net_17661)
	);

	bfr new_net_17662_bfr_after (
		.din(new_net_17661),
		.dout(new_net_17662)
	);

	bfr new_net_17663_bfr_after (
		.din(new_net_17662),
		.dout(new_net_17663)
	);

	bfr new_net_17664_bfr_after (
		.din(new_net_17663),
		.dout(new_net_17664)
	);

	bfr new_net_17665_bfr_after (
		.din(new_net_17664),
		.dout(new_net_17665)
	);

	bfr new_net_17666_bfr_after (
		.din(new_net_17665),
		.dout(new_net_17666)
	);

	bfr new_net_17667_bfr_after (
		.din(new_net_17666),
		.dout(new_net_17667)
	);

	bfr new_net_17668_bfr_after (
		.din(new_net_17667),
		.dout(new_net_17668)
	);

	bfr new_net_17669_bfr_after (
		.din(new_net_17668),
		.dout(new_net_17669)
	);

	bfr new_net_17670_bfr_after (
		.din(new_net_17669),
		.dout(new_net_17670)
	);

	bfr new_net_17671_bfr_after (
		.din(new_net_17670),
		.dout(new_net_17671)
	);

	bfr new_net_17672_bfr_after (
		.din(new_net_17671),
		.dout(new_net_17672)
	);

	bfr new_net_17673_bfr_after (
		.din(new_net_17672),
		.dout(new_net_17673)
	);

	bfr new_net_17674_bfr_after (
		.din(new_net_17673),
		.dout(new_net_17674)
	);

	bfr new_net_17675_bfr_after (
		.din(new_net_17674),
		.dout(new_net_17675)
	);

	bfr new_net_17676_bfr_after (
		.din(new_net_17675),
		.dout(new_net_17676)
	);

	bfr new_net_17677_bfr_after (
		.din(new_net_17676),
		.dout(new_net_17677)
	);

	bfr new_net_17678_bfr_after (
		.din(new_net_17677),
		.dout(new_net_17678)
	);

	bfr new_net_17679_bfr_after (
		.din(new_net_17678),
		.dout(new_net_17679)
	);

	bfr new_net_17680_bfr_after (
		.din(new_net_17679),
		.dout(new_net_17680)
	);

	bfr new_net_17681_bfr_after (
		.din(new_net_17680),
		.dout(new_net_17681)
	);

	bfr new_net_17682_bfr_after (
		.din(new_net_17681),
		.dout(new_net_17682)
	);

	bfr new_net_17683_bfr_after (
		.din(new_net_17682),
		.dout(new_net_17683)
	);

	bfr new_net_17684_bfr_after (
		.din(new_net_17683),
		.dout(new_net_17684)
	);

	bfr new_net_17685_bfr_after (
		.din(new_net_17684),
		.dout(new_net_17685)
	);

	bfr new_net_17686_bfr_after (
		.din(new_net_17685),
		.dout(new_net_17686)
	);

	bfr new_net_17687_bfr_after (
		.din(new_net_17686),
		.dout(new_net_17687)
	);

	bfr new_net_17688_bfr_after (
		.din(new_net_17687),
		.dout(new_net_17688)
	);

	bfr new_net_17689_bfr_after (
		.din(new_net_17688),
		.dout(new_net_17689)
	);

	bfr new_net_17690_bfr_after (
		.din(new_net_17689),
		.dout(new_net_17690)
	);

	bfr new_net_17691_bfr_after (
		.din(new_net_17690),
		.dout(new_net_17691)
	);

	bfr new_net_17692_bfr_after (
		.din(new_net_17691),
		.dout(new_net_17692)
	);

	bfr new_net_17693_bfr_after (
		.din(new_net_17692),
		.dout(new_net_17693)
	);

	bfr new_net_17694_bfr_after (
		.din(new_net_17693),
		.dout(new_net_17694)
	);

	bfr new_net_17695_bfr_after (
		.din(new_net_17694),
		.dout(new_net_17695)
	);

	bfr new_net_17696_bfr_after (
		.din(new_net_17695),
		.dout(new_net_17696)
	);

	bfr new_net_17697_bfr_after (
		.din(new_net_17696),
		.dout(new_net_17697)
	);

	bfr new_net_17698_bfr_after (
		.din(new_net_17697),
		.dout(new_net_17698)
	);

	bfr new_net_17699_bfr_after (
		.din(new_net_17698),
		.dout(new_net_17699)
	);

	bfr new_net_17700_bfr_after (
		.din(new_net_17699),
		.dout(new_net_17700)
	);

	bfr new_net_17701_bfr_after (
		.din(new_net_17700),
		.dout(new_net_17701)
	);

	bfr new_net_17702_bfr_after (
		.din(new_net_17701),
		.dout(new_net_17702)
	);

	bfr new_net_17703_bfr_after (
		.din(new_net_17702),
		.dout(new_net_17703)
	);

	bfr new_net_17704_bfr_after (
		.din(new_net_17703),
		.dout(new_net_17704)
	);

	bfr new_net_17705_bfr_after (
		.din(new_net_17704),
		.dout(new_net_17705)
	);

	bfr new_net_17706_bfr_after (
		.din(new_net_17705),
		.dout(new_net_17706)
	);

	bfr new_net_17707_bfr_after (
		.din(new_net_17706),
		.dout(new_net_17707)
	);

	bfr new_net_17708_bfr_after (
		.din(new_net_17707),
		.dout(new_net_17708)
	);

	bfr new_net_17709_bfr_after (
		.din(new_net_17708),
		.dout(new_net_17709)
	);

	bfr new_net_17710_bfr_after (
		.din(new_net_17709),
		.dout(new_net_17710)
	);

	bfr new_net_17711_bfr_after (
		.din(new_net_17710),
		.dout(new_net_17711)
	);

	bfr new_net_17712_bfr_after (
		.din(new_net_17711),
		.dout(new_net_17712)
	);

	bfr new_net_17713_bfr_after (
		.din(new_net_17712),
		.dout(new_net_17713)
	);

	bfr new_net_17714_bfr_after (
		.din(new_net_17713),
		.dout(new_net_17714)
	);

	bfr new_net_17715_bfr_after (
		.din(new_net_17714),
		.dout(new_net_17715)
	);

	bfr new_net_17716_bfr_after (
		.din(new_net_17715),
		.dout(new_net_17716)
	);

	bfr new_net_17717_bfr_after (
		.din(new_net_17716),
		.dout(new_net_17717)
	);

	bfr new_net_17718_bfr_after (
		.din(new_net_17717),
		.dout(new_net_17718)
	);

	bfr new_net_17719_bfr_after (
		.din(new_net_17718),
		.dout(new_net_17719)
	);

	bfr new_net_17720_bfr_after (
		.din(new_net_17719),
		.dout(new_net_17720)
	);

	bfr new_net_17721_bfr_after (
		.din(new_net_17720),
		.dout(new_net_17721)
	);

	bfr new_net_17722_bfr_after (
		.din(new_net_17721),
		.dout(new_net_17722)
	);

	bfr new_net_17723_bfr_after (
		.din(new_net_17722),
		.dout(new_net_17723)
	);

	bfr new_net_17724_bfr_after (
		.din(new_net_17723),
		.dout(new_net_17724)
	);

	bfr new_net_17725_bfr_after (
		.din(new_net_17724),
		.dout(new_net_17725)
	);

	bfr new_net_17726_bfr_after (
		.din(new_net_17725),
		.dout(new_net_17726)
	);

	bfr new_net_17727_bfr_after (
		.din(new_net_17726),
		.dout(new_net_17727)
	);

	bfr new_net_17728_bfr_after (
		.din(new_net_17727),
		.dout(new_net_17728)
	);

	bfr new_net_17729_bfr_after (
		.din(new_net_17728),
		.dout(new_net_17729)
	);

	bfr new_net_17730_bfr_after (
		.din(new_net_17729),
		.dout(new_net_17730)
	);

	bfr new_net_17731_bfr_after (
		.din(new_net_17730),
		.dout(new_net_17731)
	);

	bfr new_net_17732_bfr_after (
		.din(new_net_17731),
		.dout(new_net_17732)
	);

	bfr new_net_17733_bfr_after (
		.din(new_net_17732),
		.dout(new_net_17733)
	);

	bfr new_net_17734_bfr_after (
		.din(new_net_17733),
		.dout(new_net_17734)
	);

	bfr new_net_17735_bfr_after (
		.din(new_net_17734),
		.dout(new_net_17735)
	);

	bfr new_net_17736_bfr_after (
		.din(new_net_17735),
		.dout(new_net_17736)
	);

	bfr new_net_17737_bfr_after (
		.din(new_net_17736),
		.dout(new_net_17737)
	);

	bfr new_net_17738_bfr_after (
		.din(new_net_17737),
		.dout(new_net_17738)
	);

	bfr new_net_17739_bfr_after (
		.din(new_net_17738),
		.dout(new_net_17739)
	);

	bfr new_net_17740_bfr_after (
		.din(new_net_17739),
		.dout(new_net_17740)
	);

	bfr new_net_17741_bfr_after (
		.din(new_net_17740),
		.dout(new_net_17741)
	);

	bfr new_net_17742_bfr_after (
		.din(new_net_17741),
		.dout(new_net_17742)
	);

	bfr new_net_17743_bfr_after (
		.din(new_net_17742),
		.dout(new_net_17743)
	);

	bfr new_net_17744_bfr_after (
		.din(new_net_17743),
		.dout(new_net_17744)
	);

	bfr new_net_17745_bfr_after (
		.din(new_net_17744),
		.dout(new_net_17745)
	);

	bfr new_net_17746_bfr_after (
		.din(new_net_17745),
		.dout(new_net_17746)
	);

	bfr new_net_17747_bfr_after (
		.din(new_net_17746),
		.dout(new_net_17747)
	);

	bfr new_net_17748_bfr_after (
		.din(new_net_17747),
		.dout(new_net_17748)
	);

	bfr new_net_17749_bfr_after (
		.din(new_net_17748),
		.dout(new_net_17749)
	);

	bfr new_net_17750_bfr_after (
		.din(new_net_17749),
		.dout(new_net_17750)
	);

	bfr new_net_17751_bfr_after (
		.din(new_net_17750),
		.dout(new_net_17751)
	);

	bfr new_net_17752_bfr_after (
		.din(new_net_17751),
		.dout(new_net_17752)
	);

	bfr new_net_17753_bfr_after (
		.din(new_net_17752),
		.dout(new_net_17753)
	);

	bfr new_net_17754_bfr_after (
		.din(new_net_17753),
		.dout(new_net_17754)
	);

	spl2 _0829__v_fanout (
		.a(new_net_17754),
		.b(new_net_2232),
		.c(new_net_2233)
	);

	bfr new_net_17755_bfr_after (
		.din(_0931_),
		.dout(new_net_17755)
	);

	bfr new_net_17756_bfr_after (
		.din(new_net_17755),
		.dout(new_net_17756)
	);

	bfr new_net_17757_bfr_after (
		.din(new_net_17756),
		.dout(new_net_17757)
	);

	bfr new_net_17758_bfr_after (
		.din(new_net_17757),
		.dout(new_net_17758)
	);

	bfr new_net_17759_bfr_after (
		.din(new_net_17758),
		.dout(new_net_17759)
	);

	bfr new_net_17760_bfr_after (
		.din(new_net_17759),
		.dout(new_net_17760)
	);

	bfr new_net_17761_bfr_after (
		.din(new_net_17760),
		.dout(new_net_17761)
	);

	bfr new_net_17762_bfr_after (
		.din(new_net_17761),
		.dout(new_net_17762)
	);

	bfr new_net_17763_bfr_after (
		.din(new_net_17762),
		.dout(new_net_17763)
	);

	bfr new_net_17764_bfr_after (
		.din(new_net_17763),
		.dout(new_net_17764)
	);

	bfr new_net_17765_bfr_after (
		.din(new_net_17764),
		.dout(new_net_17765)
	);

	bfr new_net_17766_bfr_after (
		.din(new_net_17765),
		.dout(new_net_17766)
	);

	bfr new_net_17767_bfr_after (
		.din(new_net_17766),
		.dout(new_net_17767)
	);

	bfr new_net_17768_bfr_after (
		.din(new_net_17767),
		.dout(new_net_17768)
	);

	bfr new_net_17769_bfr_after (
		.din(new_net_17768),
		.dout(new_net_17769)
	);

	bfr new_net_17770_bfr_after (
		.din(new_net_17769),
		.dout(new_net_17770)
	);

	bfr new_net_17771_bfr_after (
		.din(new_net_17770),
		.dout(new_net_17771)
	);

	bfr new_net_17772_bfr_after (
		.din(new_net_17771),
		.dout(new_net_17772)
	);

	bfr new_net_17773_bfr_after (
		.din(new_net_17772),
		.dout(new_net_17773)
	);

	bfr new_net_17774_bfr_after (
		.din(new_net_17773),
		.dout(new_net_17774)
	);

	bfr new_net_17775_bfr_after (
		.din(new_net_17774),
		.dout(new_net_17775)
	);

	bfr new_net_17776_bfr_after (
		.din(new_net_17775),
		.dout(new_net_17776)
	);

	bfr new_net_17777_bfr_after (
		.din(new_net_17776),
		.dout(new_net_17777)
	);

	bfr new_net_17778_bfr_after (
		.din(new_net_17777),
		.dout(new_net_17778)
	);

	bfr new_net_17779_bfr_after (
		.din(new_net_17778),
		.dout(new_net_17779)
	);

	bfr new_net_17780_bfr_after (
		.din(new_net_17779),
		.dout(new_net_17780)
	);

	bfr new_net_17781_bfr_after (
		.din(new_net_17780),
		.dout(new_net_17781)
	);

	bfr new_net_17782_bfr_after (
		.din(new_net_17781),
		.dout(new_net_17782)
	);

	bfr new_net_17783_bfr_after (
		.din(new_net_17782),
		.dout(new_net_17783)
	);

	bfr new_net_17784_bfr_after (
		.din(new_net_17783),
		.dout(new_net_17784)
	);

	bfr new_net_17785_bfr_after (
		.din(new_net_17784),
		.dout(new_net_17785)
	);

	bfr new_net_17786_bfr_after (
		.din(new_net_17785),
		.dout(new_net_17786)
	);

	bfr new_net_17787_bfr_after (
		.din(new_net_17786),
		.dout(new_net_17787)
	);

	bfr new_net_17788_bfr_after (
		.din(new_net_17787),
		.dout(new_net_17788)
	);

	bfr new_net_17789_bfr_after (
		.din(new_net_17788),
		.dout(new_net_17789)
	);

	bfr new_net_17790_bfr_after (
		.din(new_net_17789),
		.dout(new_net_17790)
	);

	bfr new_net_17791_bfr_after (
		.din(new_net_17790),
		.dout(new_net_17791)
	);

	bfr new_net_17792_bfr_after (
		.din(new_net_17791),
		.dout(new_net_17792)
	);

	bfr new_net_17793_bfr_after (
		.din(new_net_17792),
		.dout(new_net_17793)
	);

	bfr new_net_17794_bfr_after (
		.din(new_net_17793),
		.dout(new_net_17794)
	);

	bfr new_net_17795_bfr_after (
		.din(new_net_17794),
		.dout(new_net_17795)
	);

	bfr new_net_17796_bfr_after (
		.din(new_net_17795),
		.dout(new_net_17796)
	);

	bfr new_net_17797_bfr_after (
		.din(new_net_17796),
		.dout(new_net_17797)
	);

	bfr new_net_17798_bfr_after (
		.din(new_net_17797),
		.dout(new_net_17798)
	);

	bfr new_net_17799_bfr_after (
		.din(new_net_17798),
		.dout(new_net_17799)
	);

	bfr new_net_17800_bfr_after (
		.din(new_net_17799),
		.dout(new_net_17800)
	);

	bfr new_net_17801_bfr_after (
		.din(new_net_17800),
		.dout(new_net_17801)
	);

	bfr new_net_17802_bfr_after (
		.din(new_net_17801),
		.dout(new_net_17802)
	);

	bfr new_net_17803_bfr_after (
		.din(new_net_17802),
		.dout(new_net_17803)
	);

	bfr new_net_17804_bfr_after (
		.din(new_net_17803),
		.dout(new_net_17804)
	);

	bfr new_net_17805_bfr_after (
		.din(new_net_17804),
		.dout(new_net_17805)
	);

	bfr new_net_17806_bfr_after (
		.din(new_net_17805),
		.dout(new_net_17806)
	);

	bfr new_net_17807_bfr_after (
		.din(new_net_17806),
		.dout(new_net_17807)
	);

	bfr new_net_17808_bfr_after (
		.din(new_net_17807),
		.dout(new_net_17808)
	);

	bfr new_net_17809_bfr_after (
		.din(new_net_17808),
		.dout(new_net_17809)
	);

	bfr new_net_17810_bfr_after (
		.din(new_net_17809),
		.dout(new_net_17810)
	);

	bfr new_net_17811_bfr_after (
		.din(new_net_17810),
		.dout(new_net_17811)
	);

	bfr new_net_17812_bfr_after (
		.din(new_net_17811),
		.dout(new_net_17812)
	);

	bfr new_net_17813_bfr_after (
		.din(new_net_17812),
		.dout(new_net_17813)
	);

	bfr new_net_17814_bfr_after (
		.din(new_net_17813),
		.dout(new_net_17814)
	);

	bfr new_net_17815_bfr_after (
		.din(new_net_17814),
		.dout(new_net_17815)
	);

	bfr new_net_17816_bfr_after (
		.din(new_net_17815),
		.dout(new_net_17816)
	);

	bfr new_net_17817_bfr_after (
		.din(new_net_17816),
		.dout(new_net_17817)
	);

	bfr new_net_17818_bfr_after (
		.din(new_net_17817),
		.dout(new_net_17818)
	);

	bfr new_net_17819_bfr_after (
		.din(new_net_17818),
		.dout(new_net_17819)
	);

	bfr new_net_17820_bfr_after (
		.din(new_net_17819),
		.dout(new_net_17820)
	);

	bfr new_net_17821_bfr_after (
		.din(new_net_17820),
		.dout(new_net_17821)
	);

	bfr new_net_17822_bfr_after (
		.din(new_net_17821),
		.dout(new_net_17822)
	);

	bfr new_net_17823_bfr_after (
		.din(new_net_17822),
		.dout(new_net_17823)
	);

	bfr new_net_17824_bfr_after (
		.din(new_net_17823),
		.dout(new_net_17824)
	);

	bfr new_net_17825_bfr_after (
		.din(new_net_17824),
		.dout(new_net_17825)
	);

	bfr new_net_17826_bfr_after (
		.din(new_net_17825),
		.dout(new_net_17826)
	);

	bfr new_net_17827_bfr_after (
		.din(new_net_17826),
		.dout(new_net_17827)
	);

	bfr new_net_17828_bfr_after (
		.din(new_net_17827),
		.dout(new_net_17828)
	);

	bfr new_net_17829_bfr_after (
		.din(new_net_17828),
		.dout(new_net_17829)
	);

	bfr new_net_17830_bfr_after (
		.din(new_net_17829),
		.dout(new_net_17830)
	);

	bfr new_net_17831_bfr_after (
		.din(new_net_17830),
		.dout(new_net_17831)
	);

	bfr new_net_17832_bfr_after (
		.din(new_net_17831),
		.dout(new_net_17832)
	);

	bfr new_net_17833_bfr_after (
		.din(new_net_17832),
		.dout(new_net_17833)
	);

	bfr new_net_17834_bfr_after (
		.din(new_net_17833),
		.dout(new_net_17834)
	);

	bfr new_net_17835_bfr_after (
		.din(new_net_17834),
		.dout(new_net_17835)
	);

	bfr new_net_17836_bfr_after (
		.din(new_net_17835),
		.dout(new_net_17836)
	);

	bfr new_net_17837_bfr_after (
		.din(new_net_17836),
		.dout(new_net_17837)
	);

	bfr new_net_17838_bfr_after (
		.din(new_net_17837),
		.dout(new_net_17838)
	);

	bfr new_net_17839_bfr_after (
		.din(new_net_17838),
		.dout(new_net_17839)
	);

	bfr new_net_17840_bfr_after (
		.din(new_net_17839),
		.dout(new_net_17840)
	);

	spl2 _0931__v_fanout (
		.a(new_net_17840),
		.b(new_net_1507),
		.c(new_net_1508)
	);

	bfr new_net_17841_bfr_after (
		.din(_0079_),
		.dout(new_net_17841)
	);

	bfr new_net_17842_bfr_after (
		.din(new_net_17841),
		.dout(new_net_17842)
	);

	bfr new_net_17843_bfr_after (
		.din(new_net_17842),
		.dout(new_net_17843)
	);

	bfr new_net_17844_bfr_after (
		.din(new_net_17843),
		.dout(new_net_17844)
	);

	bfr new_net_17845_bfr_after (
		.din(new_net_17844),
		.dout(new_net_17845)
	);

	bfr new_net_17846_bfr_after (
		.din(new_net_17845),
		.dout(new_net_17846)
	);

	bfr new_net_17847_bfr_after (
		.din(new_net_17846),
		.dout(new_net_17847)
	);

	bfr new_net_17848_bfr_after (
		.din(new_net_17847),
		.dout(new_net_17848)
	);

	bfr new_net_17849_bfr_after (
		.din(new_net_17848),
		.dout(new_net_17849)
	);

	bfr new_net_17850_bfr_after (
		.din(new_net_17849),
		.dout(new_net_17850)
	);

	bfr new_net_17851_bfr_after (
		.din(new_net_17850),
		.dout(new_net_17851)
	);

	bfr new_net_17852_bfr_after (
		.din(new_net_17851),
		.dout(new_net_17852)
	);

	bfr new_net_17853_bfr_after (
		.din(new_net_17852),
		.dout(new_net_17853)
	);

	bfr new_net_17854_bfr_after (
		.din(new_net_17853),
		.dout(new_net_17854)
	);

	bfr new_net_17855_bfr_after (
		.din(new_net_17854),
		.dout(new_net_17855)
	);

	bfr new_net_17856_bfr_after (
		.din(new_net_17855),
		.dout(new_net_17856)
	);

	bfr new_net_17857_bfr_after (
		.din(new_net_17856),
		.dout(new_net_17857)
	);

	bfr new_net_17858_bfr_after (
		.din(new_net_17857),
		.dout(new_net_17858)
	);

	bfr new_net_17859_bfr_after (
		.din(new_net_17858),
		.dout(new_net_17859)
	);

	bfr new_net_17860_bfr_after (
		.din(new_net_17859),
		.dout(new_net_17860)
	);

	bfr new_net_17861_bfr_after (
		.din(new_net_17860),
		.dout(new_net_17861)
	);

	bfr new_net_17862_bfr_after (
		.din(new_net_17861),
		.dout(new_net_17862)
	);

	bfr new_net_17863_bfr_after (
		.din(new_net_17862),
		.dout(new_net_17863)
	);

	bfr new_net_17864_bfr_after (
		.din(new_net_17863),
		.dout(new_net_17864)
	);

	bfr new_net_17865_bfr_after (
		.din(new_net_17864),
		.dout(new_net_17865)
	);

	bfr new_net_17866_bfr_after (
		.din(new_net_17865),
		.dout(new_net_17866)
	);

	bfr new_net_17867_bfr_after (
		.din(new_net_17866),
		.dout(new_net_17867)
	);

	bfr new_net_17868_bfr_after (
		.din(new_net_17867),
		.dout(new_net_17868)
	);

	bfr new_net_17869_bfr_after (
		.din(new_net_17868),
		.dout(new_net_17869)
	);

	bfr new_net_17870_bfr_after (
		.din(new_net_17869),
		.dout(new_net_17870)
	);

	bfr new_net_17871_bfr_after (
		.din(new_net_17870),
		.dout(new_net_17871)
	);

	bfr new_net_17872_bfr_after (
		.din(new_net_17871),
		.dout(new_net_17872)
	);

	bfr new_net_17873_bfr_after (
		.din(new_net_17872),
		.dout(new_net_17873)
	);

	bfr new_net_17874_bfr_after (
		.din(new_net_17873),
		.dout(new_net_17874)
	);

	bfr new_net_17875_bfr_after (
		.din(new_net_17874),
		.dout(new_net_17875)
	);

	bfr new_net_17876_bfr_after (
		.din(new_net_17875),
		.dout(new_net_17876)
	);

	bfr new_net_17877_bfr_after (
		.din(new_net_17876),
		.dout(new_net_17877)
	);

	bfr new_net_17878_bfr_after (
		.din(new_net_17877),
		.dout(new_net_17878)
	);

	bfr new_net_17879_bfr_after (
		.din(new_net_17878),
		.dout(new_net_17879)
	);

	bfr new_net_17880_bfr_after (
		.din(new_net_17879),
		.dout(new_net_17880)
	);

	bfr new_net_17881_bfr_after (
		.din(new_net_17880),
		.dout(new_net_17881)
	);

	bfr new_net_17882_bfr_after (
		.din(new_net_17881),
		.dout(new_net_17882)
	);

	bfr new_net_17883_bfr_after (
		.din(new_net_17882),
		.dout(new_net_17883)
	);

	bfr new_net_17884_bfr_after (
		.din(new_net_17883),
		.dout(new_net_17884)
	);

	bfr new_net_17885_bfr_after (
		.din(new_net_17884),
		.dout(new_net_17885)
	);

	bfr new_net_17886_bfr_after (
		.din(new_net_17885),
		.dout(new_net_17886)
	);

	bfr new_net_17887_bfr_after (
		.din(new_net_17886),
		.dout(new_net_17887)
	);

	bfr new_net_17888_bfr_after (
		.din(new_net_17887),
		.dout(new_net_17888)
	);

	bfr new_net_17889_bfr_after (
		.din(new_net_17888),
		.dout(new_net_17889)
	);

	bfr new_net_17890_bfr_after (
		.din(new_net_17889),
		.dout(new_net_17890)
	);

	bfr new_net_17891_bfr_after (
		.din(new_net_17890),
		.dout(new_net_17891)
	);

	bfr new_net_17892_bfr_after (
		.din(new_net_17891),
		.dout(new_net_17892)
	);

	bfr new_net_17893_bfr_after (
		.din(new_net_17892),
		.dout(new_net_17893)
	);

	bfr new_net_17894_bfr_after (
		.din(new_net_17893),
		.dout(new_net_17894)
	);

	bfr new_net_17895_bfr_after (
		.din(new_net_17894),
		.dout(new_net_17895)
	);

	bfr new_net_17896_bfr_after (
		.din(new_net_17895),
		.dout(new_net_17896)
	);

	bfr new_net_17897_bfr_after (
		.din(new_net_17896),
		.dout(new_net_17897)
	);

	bfr new_net_17898_bfr_after (
		.din(new_net_17897),
		.dout(new_net_17898)
	);

	bfr new_net_17899_bfr_after (
		.din(new_net_17898),
		.dout(new_net_17899)
	);

	bfr new_net_17900_bfr_after (
		.din(new_net_17899),
		.dout(new_net_17900)
	);

	bfr new_net_17901_bfr_after (
		.din(new_net_17900),
		.dout(new_net_17901)
	);

	bfr new_net_17902_bfr_after (
		.din(new_net_17901),
		.dout(new_net_17902)
	);

	bfr new_net_17903_bfr_after (
		.din(new_net_17902),
		.dout(new_net_17903)
	);

	bfr new_net_17904_bfr_after (
		.din(new_net_17903),
		.dout(new_net_17904)
	);

	bfr new_net_17905_bfr_after (
		.din(new_net_17904),
		.dout(new_net_17905)
	);

	bfr new_net_17906_bfr_after (
		.din(new_net_17905),
		.dout(new_net_17906)
	);

	bfr new_net_17907_bfr_after (
		.din(new_net_17906),
		.dout(new_net_17907)
	);

	bfr new_net_17908_bfr_after (
		.din(new_net_17907),
		.dout(new_net_17908)
	);

	bfr new_net_17909_bfr_after (
		.din(new_net_17908),
		.dout(new_net_17909)
	);

	bfr new_net_17910_bfr_after (
		.din(new_net_17909),
		.dout(new_net_17910)
	);

	bfr new_net_17911_bfr_after (
		.din(new_net_17910),
		.dout(new_net_17911)
	);

	bfr new_net_17912_bfr_after (
		.din(new_net_17911),
		.dout(new_net_17912)
	);

	bfr new_net_17913_bfr_after (
		.din(new_net_17912),
		.dout(new_net_17913)
	);

	bfr new_net_17914_bfr_after (
		.din(new_net_17913),
		.dout(new_net_17914)
	);

	bfr new_net_17915_bfr_after (
		.din(new_net_17914),
		.dout(new_net_17915)
	);

	bfr new_net_17916_bfr_after (
		.din(new_net_17915),
		.dout(new_net_17916)
	);

	bfr new_net_17917_bfr_after (
		.din(new_net_17916),
		.dout(new_net_17917)
	);

	bfr new_net_17918_bfr_after (
		.din(new_net_17917),
		.dout(new_net_17918)
	);

	bfr new_net_17919_bfr_after (
		.din(new_net_17918),
		.dout(new_net_17919)
	);

	bfr new_net_17920_bfr_after (
		.din(new_net_17919),
		.dout(new_net_17920)
	);

	bfr new_net_17921_bfr_after (
		.din(new_net_17920),
		.dout(new_net_17921)
	);

	bfr new_net_17922_bfr_after (
		.din(new_net_17921),
		.dout(new_net_17922)
	);

	bfr new_net_17923_bfr_after (
		.din(new_net_17922),
		.dout(new_net_17923)
	);

	bfr new_net_17924_bfr_after (
		.din(new_net_17923),
		.dout(new_net_17924)
	);

	bfr new_net_17925_bfr_after (
		.din(new_net_17924),
		.dout(new_net_17925)
	);

	bfr new_net_17926_bfr_after (
		.din(new_net_17925),
		.dout(new_net_17926)
	);

	bfr new_net_17927_bfr_after (
		.din(new_net_17926),
		.dout(new_net_17927)
	);

	bfr new_net_17928_bfr_after (
		.din(new_net_17927),
		.dout(new_net_17928)
	);

	bfr new_net_17929_bfr_after (
		.din(new_net_17928),
		.dout(new_net_17929)
	);

	bfr new_net_17930_bfr_after (
		.din(new_net_17929),
		.dout(new_net_17930)
	);

	bfr new_net_17931_bfr_after (
		.din(new_net_17930),
		.dout(new_net_17931)
	);

	bfr new_net_17932_bfr_after (
		.din(new_net_17931),
		.dout(new_net_17932)
	);

	bfr new_net_17933_bfr_after (
		.din(new_net_17932),
		.dout(new_net_17933)
	);

	bfr new_net_17934_bfr_after (
		.din(new_net_17933),
		.dout(new_net_17934)
	);

	bfr new_net_17935_bfr_after (
		.din(new_net_17934),
		.dout(new_net_17935)
	);

	bfr new_net_17936_bfr_after (
		.din(new_net_17935),
		.dout(new_net_17936)
	);

	bfr new_net_17937_bfr_after (
		.din(new_net_17936),
		.dout(new_net_17937)
	);

	bfr new_net_17938_bfr_after (
		.din(new_net_17937),
		.dout(new_net_17938)
	);

	bfr new_net_17939_bfr_after (
		.din(new_net_17938),
		.dout(new_net_17939)
	);

	bfr new_net_17940_bfr_after (
		.din(new_net_17939),
		.dout(new_net_17940)
	);

	bfr new_net_17941_bfr_after (
		.din(new_net_17940),
		.dout(new_net_17941)
	);

	bfr new_net_17942_bfr_after (
		.din(new_net_17941),
		.dout(new_net_17942)
	);

	bfr new_net_17943_bfr_after (
		.din(new_net_17942),
		.dout(new_net_17943)
	);

	bfr new_net_17944_bfr_after (
		.din(new_net_17943),
		.dout(new_net_17944)
	);

	bfr new_net_17945_bfr_after (
		.din(new_net_17944),
		.dout(new_net_17945)
	);

	bfr new_net_17946_bfr_after (
		.din(new_net_17945),
		.dout(new_net_17946)
	);

	bfr new_net_17947_bfr_after (
		.din(new_net_17946),
		.dout(new_net_17947)
	);

	bfr new_net_17948_bfr_after (
		.din(new_net_17947),
		.dout(new_net_17948)
	);

	bfr new_net_17949_bfr_after (
		.din(new_net_17948),
		.dout(new_net_17949)
	);

	bfr new_net_17950_bfr_after (
		.din(new_net_17949),
		.dout(new_net_17950)
	);

	bfr new_net_17951_bfr_after (
		.din(new_net_17950),
		.dout(new_net_17951)
	);

	bfr new_net_17952_bfr_after (
		.din(new_net_17951),
		.dout(new_net_17952)
	);

	spl2 _0079__v_fanout (
		.a(new_net_17952),
		.b(new_net_2460),
		.c(new_net_2461)
	);

	bfr new_net_17953_bfr_after (
		.din(_0833_),
		.dout(new_net_17953)
	);

	bfr new_net_17954_bfr_after (
		.din(new_net_17953),
		.dout(new_net_17954)
	);

	bfr new_net_17955_bfr_after (
		.din(new_net_17954),
		.dout(new_net_17955)
	);

	bfr new_net_17956_bfr_after (
		.din(new_net_17955),
		.dout(new_net_17956)
	);

	bfr new_net_17957_bfr_after (
		.din(new_net_17956),
		.dout(new_net_17957)
	);

	bfr new_net_17958_bfr_after (
		.din(new_net_17957),
		.dout(new_net_17958)
	);

	bfr new_net_17959_bfr_after (
		.din(new_net_17958),
		.dout(new_net_17959)
	);

	bfr new_net_17960_bfr_after (
		.din(new_net_17959),
		.dout(new_net_17960)
	);

	bfr new_net_17961_bfr_after (
		.din(new_net_17960),
		.dout(new_net_17961)
	);

	bfr new_net_17962_bfr_after (
		.din(new_net_17961),
		.dout(new_net_17962)
	);

	bfr new_net_17963_bfr_after (
		.din(new_net_17962),
		.dout(new_net_17963)
	);

	bfr new_net_17964_bfr_after (
		.din(new_net_17963),
		.dout(new_net_17964)
	);

	bfr new_net_17965_bfr_after (
		.din(new_net_17964),
		.dout(new_net_17965)
	);

	bfr new_net_17966_bfr_after (
		.din(new_net_17965),
		.dout(new_net_17966)
	);

	bfr new_net_17967_bfr_after (
		.din(new_net_17966),
		.dout(new_net_17967)
	);

	bfr new_net_17968_bfr_after (
		.din(new_net_17967),
		.dout(new_net_17968)
	);

	bfr new_net_17969_bfr_after (
		.din(new_net_17968),
		.dout(new_net_17969)
	);

	bfr new_net_17970_bfr_after (
		.din(new_net_17969),
		.dout(new_net_17970)
	);

	bfr new_net_17971_bfr_after (
		.din(new_net_17970),
		.dout(new_net_17971)
	);

	bfr new_net_17972_bfr_after (
		.din(new_net_17971),
		.dout(new_net_17972)
	);

	bfr new_net_17973_bfr_after (
		.din(new_net_17972),
		.dout(new_net_17973)
	);

	bfr new_net_17974_bfr_after (
		.din(new_net_17973),
		.dout(new_net_17974)
	);

	bfr new_net_17975_bfr_after (
		.din(new_net_17974),
		.dout(new_net_17975)
	);

	bfr new_net_17976_bfr_after (
		.din(new_net_17975),
		.dout(new_net_17976)
	);

	bfr new_net_17977_bfr_after (
		.din(new_net_17976),
		.dout(new_net_17977)
	);

	bfr new_net_17978_bfr_after (
		.din(new_net_17977),
		.dout(new_net_17978)
	);

	bfr new_net_17979_bfr_after (
		.din(new_net_17978),
		.dout(new_net_17979)
	);

	bfr new_net_17980_bfr_after (
		.din(new_net_17979),
		.dout(new_net_17980)
	);

	bfr new_net_17981_bfr_after (
		.din(new_net_17980),
		.dout(new_net_17981)
	);

	bfr new_net_17982_bfr_after (
		.din(new_net_17981),
		.dout(new_net_17982)
	);

	bfr new_net_17983_bfr_after (
		.din(new_net_17982),
		.dout(new_net_17983)
	);

	bfr new_net_17984_bfr_after (
		.din(new_net_17983),
		.dout(new_net_17984)
	);

	bfr new_net_17985_bfr_after (
		.din(new_net_17984),
		.dout(new_net_17985)
	);

	bfr new_net_17986_bfr_after (
		.din(new_net_17985),
		.dout(new_net_17986)
	);

	bfr new_net_17987_bfr_after (
		.din(new_net_17986),
		.dout(new_net_17987)
	);

	bfr new_net_17988_bfr_after (
		.din(new_net_17987),
		.dout(new_net_17988)
	);

	bfr new_net_17989_bfr_after (
		.din(new_net_17988),
		.dout(new_net_17989)
	);

	bfr new_net_17990_bfr_after (
		.din(new_net_17989),
		.dout(new_net_17990)
	);

	bfr new_net_17991_bfr_after (
		.din(new_net_17990),
		.dout(new_net_17991)
	);

	bfr new_net_17992_bfr_after (
		.din(new_net_17991),
		.dout(new_net_17992)
	);

	bfr new_net_17993_bfr_after (
		.din(new_net_17992),
		.dout(new_net_17993)
	);

	bfr new_net_17994_bfr_after (
		.din(new_net_17993),
		.dout(new_net_17994)
	);

	bfr new_net_17995_bfr_after (
		.din(new_net_17994),
		.dout(new_net_17995)
	);

	bfr new_net_17996_bfr_after (
		.din(new_net_17995),
		.dout(new_net_17996)
	);

	bfr new_net_17997_bfr_after (
		.din(new_net_17996),
		.dout(new_net_17997)
	);

	bfr new_net_17998_bfr_after (
		.din(new_net_17997),
		.dout(new_net_17998)
	);

	bfr new_net_17999_bfr_after (
		.din(new_net_17998),
		.dout(new_net_17999)
	);

	bfr new_net_18000_bfr_after (
		.din(new_net_17999),
		.dout(new_net_18000)
	);

	bfr new_net_18001_bfr_after (
		.din(new_net_18000),
		.dout(new_net_18001)
	);

	bfr new_net_18002_bfr_after (
		.din(new_net_18001),
		.dout(new_net_18002)
	);

	bfr new_net_18003_bfr_after (
		.din(new_net_18002),
		.dout(new_net_18003)
	);

	bfr new_net_18004_bfr_after (
		.din(new_net_18003),
		.dout(new_net_18004)
	);

	bfr new_net_18005_bfr_after (
		.din(new_net_18004),
		.dout(new_net_18005)
	);

	bfr new_net_18006_bfr_after (
		.din(new_net_18005),
		.dout(new_net_18006)
	);

	bfr new_net_18007_bfr_after (
		.din(new_net_18006),
		.dout(new_net_18007)
	);

	bfr new_net_18008_bfr_after (
		.din(new_net_18007),
		.dout(new_net_18008)
	);

	bfr new_net_18009_bfr_after (
		.din(new_net_18008),
		.dout(new_net_18009)
	);

	bfr new_net_18010_bfr_after (
		.din(new_net_18009),
		.dout(new_net_18010)
	);

	bfr new_net_18011_bfr_after (
		.din(new_net_18010),
		.dout(new_net_18011)
	);

	bfr new_net_18012_bfr_after (
		.din(new_net_18011),
		.dout(new_net_18012)
	);

	bfr new_net_18013_bfr_after (
		.din(new_net_18012),
		.dout(new_net_18013)
	);

	bfr new_net_18014_bfr_after (
		.din(new_net_18013),
		.dout(new_net_18014)
	);

	bfr new_net_18015_bfr_after (
		.din(new_net_18014),
		.dout(new_net_18015)
	);

	bfr new_net_18016_bfr_after (
		.din(new_net_18015),
		.dout(new_net_18016)
	);

	bfr new_net_18017_bfr_after (
		.din(new_net_18016),
		.dout(new_net_18017)
	);

	bfr new_net_18018_bfr_after (
		.din(new_net_18017),
		.dout(new_net_18018)
	);

	bfr new_net_18019_bfr_after (
		.din(new_net_18018),
		.dout(new_net_18019)
	);

	bfr new_net_18020_bfr_after (
		.din(new_net_18019),
		.dout(new_net_18020)
	);

	bfr new_net_18021_bfr_after (
		.din(new_net_18020),
		.dout(new_net_18021)
	);

	bfr new_net_18022_bfr_after (
		.din(new_net_18021),
		.dout(new_net_18022)
	);

	bfr new_net_18023_bfr_after (
		.din(new_net_18022),
		.dout(new_net_18023)
	);

	bfr new_net_18024_bfr_after (
		.din(new_net_18023),
		.dout(new_net_18024)
	);

	bfr new_net_18025_bfr_after (
		.din(new_net_18024),
		.dout(new_net_18025)
	);

	bfr new_net_18026_bfr_after (
		.din(new_net_18025),
		.dout(new_net_18026)
	);

	bfr new_net_18027_bfr_after (
		.din(new_net_18026),
		.dout(new_net_18027)
	);

	bfr new_net_18028_bfr_after (
		.din(new_net_18027),
		.dout(new_net_18028)
	);

	bfr new_net_18029_bfr_after (
		.din(new_net_18028),
		.dout(new_net_18029)
	);

	bfr new_net_18030_bfr_after (
		.din(new_net_18029),
		.dout(new_net_18030)
	);

	bfr new_net_18031_bfr_after (
		.din(new_net_18030),
		.dout(new_net_18031)
	);

	bfr new_net_18032_bfr_after (
		.din(new_net_18031),
		.dout(new_net_18032)
	);

	bfr new_net_18033_bfr_after (
		.din(new_net_18032),
		.dout(new_net_18033)
	);

	bfr new_net_18034_bfr_after (
		.din(new_net_18033),
		.dout(new_net_18034)
	);

	bfr new_net_18035_bfr_after (
		.din(new_net_18034),
		.dout(new_net_18035)
	);

	bfr new_net_18036_bfr_after (
		.din(new_net_18035),
		.dout(new_net_18036)
	);

	bfr new_net_18037_bfr_after (
		.din(new_net_18036),
		.dout(new_net_18037)
	);

	bfr new_net_18038_bfr_after (
		.din(new_net_18037),
		.dout(new_net_18038)
	);

	bfr new_net_18039_bfr_after (
		.din(new_net_18038),
		.dout(new_net_18039)
	);

	bfr new_net_18040_bfr_after (
		.din(new_net_18039),
		.dout(new_net_18040)
	);

	bfr new_net_18041_bfr_after (
		.din(new_net_18040),
		.dout(new_net_18041)
	);

	bfr new_net_18042_bfr_after (
		.din(new_net_18041),
		.dout(new_net_18042)
	);

	bfr new_net_18043_bfr_after (
		.din(new_net_18042),
		.dout(new_net_18043)
	);

	bfr new_net_18044_bfr_after (
		.din(new_net_18043),
		.dout(new_net_18044)
	);

	bfr new_net_18045_bfr_after (
		.din(new_net_18044),
		.dout(new_net_18045)
	);

	bfr new_net_18046_bfr_after (
		.din(new_net_18045),
		.dout(new_net_18046)
	);

	bfr new_net_18047_bfr_after (
		.din(new_net_18046),
		.dout(new_net_18047)
	);

	bfr new_net_18048_bfr_after (
		.din(new_net_18047),
		.dout(new_net_18048)
	);

	spl2 _0833__v_fanout (
		.a(new_net_18048),
		.b(new_net_2392),
		.c(new_net_2393)
	);

	bfr new_net_18049_bfr_after (
		.din(_0223_),
		.dout(new_net_18049)
	);

	bfr new_net_18050_bfr_after (
		.din(new_net_18049),
		.dout(new_net_18050)
	);

	bfr new_net_18051_bfr_after (
		.din(new_net_18050),
		.dout(new_net_18051)
	);

	bfr new_net_18052_bfr_after (
		.din(new_net_18051),
		.dout(new_net_18052)
	);

	bfr new_net_18053_bfr_after (
		.din(new_net_18052),
		.dout(new_net_18053)
	);

	bfr new_net_18054_bfr_after (
		.din(new_net_18053),
		.dout(new_net_18054)
	);

	bfr new_net_18055_bfr_after (
		.din(new_net_18054),
		.dout(new_net_18055)
	);

	bfr new_net_18056_bfr_after (
		.din(new_net_18055),
		.dout(new_net_18056)
	);

	bfr new_net_18057_bfr_after (
		.din(new_net_18056),
		.dout(new_net_18057)
	);

	bfr new_net_18058_bfr_after (
		.din(new_net_18057),
		.dout(new_net_18058)
	);

	bfr new_net_18059_bfr_after (
		.din(new_net_18058),
		.dout(new_net_18059)
	);

	bfr new_net_18060_bfr_after (
		.din(new_net_18059),
		.dout(new_net_18060)
	);

	bfr new_net_18061_bfr_after (
		.din(new_net_18060),
		.dout(new_net_18061)
	);

	bfr new_net_18062_bfr_after (
		.din(new_net_18061),
		.dout(new_net_18062)
	);

	bfr new_net_18063_bfr_after (
		.din(new_net_18062),
		.dout(new_net_18063)
	);

	bfr new_net_18064_bfr_after (
		.din(new_net_18063),
		.dout(new_net_18064)
	);

	bfr new_net_18065_bfr_after (
		.din(new_net_18064),
		.dout(new_net_18065)
	);

	bfr new_net_18066_bfr_after (
		.din(new_net_18065),
		.dout(new_net_18066)
	);

	bfr new_net_18067_bfr_after (
		.din(new_net_18066),
		.dout(new_net_18067)
	);

	bfr new_net_18068_bfr_after (
		.din(new_net_18067),
		.dout(new_net_18068)
	);

	bfr new_net_18069_bfr_after (
		.din(new_net_18068),
		.dout(new_net_18069)
	);

	bfr new_net_18070_bfr_after (
		.din(new_net_18069),
		.dout(new_net_18070)
	);

	bfr new_net_18071_bfr_after (
		.din(new_net_18070),
		.dout(new_net_18071)
	);

	bfr new_net_18072_bfr_after (
		.din(new_net_18071),
		.dout(new_net_18072)
	);

	bfr new_net_18073_bfr_after (
		.din(new_net_18072),
		.dout(new_net_18073)
	);

	bfr new_net_18074_bfr_after (
		.din(new_net_18073),
		.dout(new_net_18074)
	);

	bfr new_net_18075_bfr_after (
		.din(new_net_18074),
		.dout(new_net_18075)
	);

	bfr new_net_18076_bfr_after (
		.din(new_net_18075),
		.dout(new_net_18076)
	);

	bfr new_net_18077_bfr_after (
		.din(new_net_18076),
		.dout(new_net_18077)
	);

	bfr new_net_18078_bfr_after (
		.din(new_net_18077),
		.dout(new_net_18078)
	);

	bfr new_net_18079_bfr_after (
		.din(new_net_18078),
		.dout(new_net_18079)
	);

	bfr new_net_18080_bfr_after (
		.din(new_net_18079),
		.dout(new_net_18080)
	);

	bfr new_net_18081_bfr_after (
		.din(new_net_18080),
		.dout(new_net_18081)
	);

	bfr new_net_18082_bfr_after (
		.din(new_net_18081),
		.dout(new_net_18082)
	);

	bfr new_net_18083_bfr_after (
		.din(new_net_18082),
		.dout(new_net_18083)
	);

	bfr new_net_18084_bfr_after (
		.din(new_net_18083),
		.dout(new_net_18084)
	);

	bfr new_net_18085_bfr_after (
		.din(new_net_18084),
		.dout(new_net_18085)
	);

	bfr new_net_18086_bfr_after (
		.din(new_net_18085),
		.dout(new_net_18086)
	);

	bfr new_net_18087_bfr_after (
		.din(new_net_18086),
		.dout(new_net_18087)
	);

	bfr new_net_18088_bfr_after (
		.din(new_net_18087),
		.dout(new_net_18088)
	);

	bfr new_net_18089_bfr_after (
		.din(new_net_18088),
		.dout(new_net_18089)
	);

	bfr new_net_18090_bfr_after (
		.din(new_net_18089),
		.dout(new_net_18090)
	);

	bfr new_net_18091_bfr_after (
		.din(new_net_18090),
		.dout(new_net_18091)
	);

	bfr new_net_18092_bfr_after (
		.din(new_net_18091),
		.dout(new_net_18092)
	);

	bfr new_net_18093_bfr_after (
		.din(new_net_18092),
		.dout(new_net_18093)
	);

	bfr new_net_18094_bfr_after (
		.din(new_net_18093),
		.dout(new_net_18094)
	);

	bfr new_net_18095_bfr_after (
		.din(new_net_18094),
		.dout(new_net_18095)
	);

	bfr new_net_18096_bfr_after (
		.din(new_net_18095),
		.dout(new_net_18096)
	);

	bfr new_net_18097_bfr_after (
		.din(new_net_18096),
		.dout(new_net_18097)
	);

	bfr new_net_18098_bfr_after (
		.din(new_net_18097),
		.dout(new_net_18098)
	);

	bfr new_net_18099_bfr_after (
		.din(new_net_18098),
		.dout(new_net_18099)
	);

	bfr new_net_18100_bfr_after (
		.din(new_net_18099),
		.dout(new_net_18100)
	);

	bfr new_net_18101_bfr_after (
		.din(new_net_18100),
		.dout(new_net_18101)
	);

	bfr new_net_18102_bfr_after (
		.din(new_net_18101),
		.dout(new_net_18102)
	);

	bfr new_net_18103_bfr_after (
		.din(new_net_18102),
		.dout(new_net_18103)
	);

	bfr new_net_18104_bfr_after (
		.din(new_net_18103),
		.dout(new_net_18104)
	);

	bfr new_net_18105_bfr_after (
		.din(new_net_18104),
		.dout(new_net_18105)
	);

	bfr new_net_18106_bfr_after (
		.din(new_net_18105),
		.dout(new_net_18106)
	);

	bfr new_net_18107_bfr_after (
		.din(new_net_18106),
		.dout(new_net_18107)
	);

	bfr new_net_18108_bfr_after (
		.din(new_net_18107),
		.dout(new_net_18108)
	);

	bfr new_net_18109_bfr_after (
		.din(new_net_18108),
		.dout(new_net_18109)
	);

	bfr new_net_18110_bfr_after (
		.din(new_net_18109),
		.dout(new_net_18110)
	);

	bfr new_net_18111_bfr_after (
		.din(new_net_18110),
		.dout(new_net_18111)
	);

	bfr new_net_18112_bfr_after (
		.din(new_net_18111),
		.dout(new_net_18112)
	);

	bfr new_net_18113_bfr_after (
		.din(new_net_18112),
		.dout(new_net_18113)
	);

	bfr new_net_18114_bfr_after (
		.din(new_net_18113),
		.dout(new_net_18114)
	);

	bfr new_net_18115_bfr_after (
		.din(new_net_18114),
		.dout(new_net_18115)
	);

	bfr new_net_18116_bfr_after (
		.din(new_net_18115),
		.dout(new_net_18116)
	);

	bfr new_net_18117_bfr_after (
		.din(new_net_18116),
		.dout(new_net_18117)
	);

	bfr new_net_18118_bfr_after (
		.din(new_net_18117),
		.dout(new_net_18118)
	);

	bfr new_net_18119_bfr_after (
		.din(new_net_18118),
		.dout(new_net_18119)
	);

	bfr new_net_18120_bfr_after (
		.din(new_net_18119),
		.dout(new_net_18120)
	);

	spl2 _0223__v_fanout (
		.a(new_net_18120),
		.b(new_net_480),
		.c(new_net_481)
	);

	bfr new_net_18121_bfr_after (
		.din(_1022_),
		.dout(new_net_18121)
	);

	bfr new_net_18122_bfr_after (
		.din(new_net_18121),
		.dout(new_net_18122)
	);

	bfr new_net_18123_bfr_after (
		.din(new_net_18122),
		.dout(new_net_18123)
	);

	bfr new_net_18124_bfr_after (
		.din(new_net_18123),
		.dout(new_net_18124)
	);

	bfr new_net_18125_bfr_after (
		.din(new_net_18124),
		.dout(new_net_18125)
	);

	bfr new_net_18126_bfr_after (
		.din(new_net_18125),
		.dout(new_net_18126)
	);

	bfr new_net_18127_bfr_after (
		.din(new_net_18126),
		.dout(new_net_18127)
	);

	bfr new_net_18128_bfr_after (
		.din(new_net_18127),
		.dout(new_net_18128)
	);

	bfr new_net_18129_bfr_after (
		.din(new_net_18128),
		.dout(new_net_18129)
	);

	bfr new_net_18130_bfr_after (
		.din(new_net_18129),
		.dout(new_net_18130)
	);

	bfr new_net_18131_bfr_after (
		.din(new_net_18130),
		.dout(new_net_18131)
	);

	bfr new_net_18132_bfr_after (
		.din(new_net_18131),
		.dout(new_net_18132)
	);

	bfr new_net_18133_bfr_after (
		.din(new_net_18132),
		.dout(new_net_18133)
	);

	bfr new_net_18134_bfr_after (
		.din(new_net_18133),
		.dout(new_net_18134)
	);

	bfr new_net_18135_bfr_after (
		.din(new_net_18134),
		.dout(new_net_18135)
	);

	bfr new_net_18136_bfr_after (
		.din(new_net_18135),
		.dout(new_net_18136)
	);

	bfr new_net_18137_bfr_after (
		.din(new_net_18136),
		.dout(new_net_18137)
	);

	bfr new_net_18138_bfr_after (
		.din(new_net_18137),
		.dout(new_net_18138)
	);

	bfr new_net_18139_bfr_after (
		.din(new_net_18138),
		.dout(new_net_18139)
	);

	bfr new_net_18140_bfr_after (
		.din(new_net_18139),
		.dout(new_net_18140)
	);

	bfr new_net_18141_bfr_after (
		.din(new_net_18140),
		.dout(new_net_18141)
	);

	bfr new_net_18142_bfr_after (
		.din(new_net_18141),
		.dout(new_net_18142)
	);

	bfr new_net_18143_bfr_after (
		.din(new_net_18142),
		.dout(new_net_18143)
	);

	bfr new_net_18144_bfr_after (
		.din(new_net_18143),
		.dout(new_net_18144)
	);

	bfr new_net_18145_bfr_after (
		.din(new_net_18144),
		.dout(new_net_18145)
	);

	bfr new_net_18146_bfr_after (
		.din(new_net_18145),
		.dout(new_net_18146)
	);

	bfr new_net_18147_bfr_after (
		.din(new_net_18146),
		.dout(new_net_18147)
	);

	bfr new_net_18148_bfr_after (
		.din(new_net_18147),
		.dout(new_net_18148)
	);

	bfr new_net_18149_bfr_after (
		.din(new_net_18148),
		.dout(new_net_18149)
	);

	bfr new_net_18150_bfr_after (
		.din(new_net_18149),
		.dout(new_net_18150)
	);

	bfr new_net_18151_bfr_after (
		.din(new_net_18150),
		.dout(new_net_18151)
	);

	bfr new_net_18152_bfr_after (
		.din(new_net_18151),
		.dout(new_net_18152)
	);

	bfr new_net_18153_bfr_after (
		.din(new_net_18152),
		.dout(new_net_18153)
	);

	bfr new_net_18154_bfr_after (
		.din(new_net_18153),
		.dout(new_net_18154)
	);

	bfr new_net_18155_bfr_after (
		.din(new_net_18154),
		.dout(new_net_18155)
	);

	bfr new_net_18156_bfr_after (
		.din(new_net_18155),
		.dout(new_net_18156)
	);

	bfr new_net_18157_bfr_after (
		.din(new_net_18156),
		.dout(new_net_18157)
	);

	bfr new_net_18158_bfr_after (
		.din(new_net_18157),
		.dout(new_net_18158)
	);

	bfr new_net_18159_bfr_after (
		.din(new_net_18158),
		.dout(new_net_18159)
	);

	bfr new_net_18160_bfr_after (
		.din(new_net_18159),
		.dout(new_net_18160)
	);

	spl2 _1022__v_fanout (
		.a(new_net_18160),
		.b(new_net_998),
		.c(new_net_999)
	);

	bfr new_net_18161_bfr_after (
		.din(_0093_),
		.dout(new_net_18161)
	);

	bfr new_net_18162_bfr_after (
		.din(new_net_18161),
		.dout(new_net_18162)
	);

	bfr new_net_18163_bfr_after (
		.din(new_net_18162),
		.dout(new_net_18163)
	);

	bfr new_net_18164_bfr_after (
		.din(new_net_18163),
		.dout(new_net_18164)
	);

	bfr new_net_18165_bfr_after (
		.din(new_net_18164),
		.dout(new_net_18165)
	);

	bfr new_net_18166_bfr_after (
		.din(new_net_18165),
		.dout(new_net_18166)
	);

	bfr new_net_18167_bfr_after (
		.din(new_net_18166),
		.dout(new_net_18167)
	);

	bfr new_net_18168_bfr_after (
		.din(new_net_18167),
		.dout(new_net_18168)
	);

	bfr new_net_18169_bfr_after (
		.din(new_net_18168),
		.dout(new_net_18169)
	);

	bfr new_net_18170_bfr_after (
		.din(new_net_18169),
		.dout(new_net_18170)
	);

	bfr new_net_18171_bfr_after (
		.din(new_net_18170),
		.dout(new_net_18171)
	);

	bfr new_net_18172_bfr_after (
		.din(new_net_18171),
		.dout(new_net_18172)
	);

	bfr new_net_18173_bfr_after (
		.din(new_net_18172),
		.dout(new_net_18173)
	);

	bfr new_net_18174_bfr_after (
		.din(new_net_18173),
		.dout(new_net_18174)
	);

	bfr new_net_18175_bfr_after (
		.din(new_net_18174),
		.dout(new_net_18175)
	);

	bfr new_net_18176_bfr_after (
		.din(new_net_18175),
		.dout(new_net_18176)
	);

	bfr new_net_18177_bfr_after (
		.din(new_net_18176),
		.dout(new_net_18177)
	);

	bfr new_net_18178_bfr_after (
		.din(new_net_18177),
		.dout(new_net_18178)
	);

	bfr new_net_18179_bfr_after (
		.din(new_net_18178),
		.dout(new_net_18179)
	);

	bfr new_net_18180_bfr_after (
		.din(new_net_18179),
		.dout(new_net_18180)
	);

	bfr new_net_18181_bfr_after (
		.din(new_net_18180),
		.dout(new_net_18181)
	);

	bfr new_net_18182_bfr_after (
		.din(new_net_18181),
		.dout(new_net_18182)
	);

	bfr new_net_18183_bfr_after (
		.din(new_net_18182),
		.dout(new_net_18183)
	);

	bfr new_net_18184_bfr_after (
		.din(new_net_18183),
		.dout(new_net_18184)
	);

	bfr new_net_18185_bfr_after (
		.din(new_net_18184),
		.dout(new_net_18185)
	);

	bfr new_net_18186_bfr_after (
		.din(new_net_18185),
		.dout(new_net_18186)
	);

	bfr new_net_18187_bfr_after (
		.din(new_net_18186),
		.dout(new_net_18187)
	);

	bfr new_net_18188_bfr_after (
		.din(new_net_18187),
		.dout(new_net_18188)
	);

	bfr new_net_18189_bfr_after (
		.din(new_net_18188),
		.dout(new_net_18189)
	);

	bfr new_net_18190_bfr_after (
		.din(new_net_18189),
		.dout(new_net_18190)
	);

	bfr new_net_18191_bfr_after (
		.din(new_net_18190),
		.dout(new_net_18191)
	);

	bfr new_net_18192_bfr_after (
		.din(new_net_18191),
		.dout(new_net_18192)
	);

	bfr new_net_18193_bfr_after (
		.din(new_net_18192),
		.dout(new_net_18193)
	);

	bfr new_net_18194_bfr_after (
		.din(new_net_18193),
		.dout(new_net_18194)
	);

	bfr new_net_18195_bfr_after (
		.din(new_net_18194),
		.dout(new_net_18195)
	);

	bfr new_net_18196_bfr_after (
		.din(new_net_18195),
		.dout(new_net_18196)
	);

	bfr new_net_18197_bfr_after (
		.din(new_net_18196),
		.dout(new_net_18197)
	);

	bfr new_net_18198_bfr_after (
		.din(new_net_18197),
		.dout(new_net_18198)
	);

	bfr new_net_18199_bfr_after (
		.din(new_net_18198),
		.dout(new_net_18199)
	);

	bfr new_net_18200_bfr_after (
		.din(new_net_18199),
		.dout(new_net_18200)
	);

	bfr new_net_18201_bfr_after (
		.din(new_net_18200),
		.dout(new_net_18201)
	);

	bfr new_net_18202_bfr_after (
		.din(new_net_18201),
		.dout(new_net_18202)
	);

	bfr new_net_18203_bfr_after (
		.din(new_net_18202),
		.dout(new_net_18203)
	);

	bfr new_net_18204_bfr_after (
		.din(new_net_18203),
		.dout(new_net_18204)
	);

	bfr new_net_18205_bfr_after (
		.din(new_net_18204),
		.dout(new_net_18205)
	);

	bfr new_net_18206_bfr_after (
		.din(new_net_18205),
		.dout(new_net_18206)
	);

	bfr new_net_18207_bfr_after (
		.din(new_net_18206),
		.dout(new_net_18207)
	);

	bfr new_net_18208_bfr_after (
		.din(new_net_18207),
		.dout(new_net_18208)
	);

	bfr new_net_18209_bfr_after (
		.din(new_net_18208),
		.dout(new_net_18209)
	);

	bfr new_net_18210_bfr_after (
		.din(new_net_18209),
		.dout(new_net_18210)
	);

	bfr new_net_18211_bfr_after (
		.din(new_net_18210),
		.dout(new_net_18211)
	);

	bfr new_net_18212_bfr_after (
		.din(new_net_18211),
		.dout(new_net_18212)
	);

	bfr new_net_18213_bfr_after (
		.din(new_net_18212),
		.dout(new_net_18213)
	);

	bfr new_net_18214_bfr_after (
		.din(new_net_18213),
		.dout(new_net_18214)
	);

	bfr new_net_18215_bfr_after (
		.din(new_net_18214),
		.dout(new_net_18215)
	);

	bfr new_net_18216_bfr_after (
		.din(new_net_18215),
		.dout(new_net_18216)
	);

	bfr new_net_18217_bfr_after (
		.din(new_net_18216),
		.dout(new_net_18217)
	);

	bfr new_net_18218_bfr_after (
		.din(new_net_18217),
		.dout(new_net_18218)
	);

	bfr new_net_18219_bfr_after (
		.din(new_net_18218),
		.dout(new_net_18219)
	);

	bfr new_net_18220_bfr_after (
		.din(new_net_18219),
		.dout(new_net_18220)
	);

	bfr new_net_18221_bfr_after (
		.din(new_net_18220),
		.dout(new_net_18221)
	);

	bfr new_net_18222_bfr_after (
		.din(new_net_18221),
		.dout(new_net_18222)
	);

	bfr new_net_18223_bfr_after (
		.din(new_net_18222),
		.dout(new_net_18223)
	);

	bfr new_net_18224_bfr_after (
		.din(new_net_18223),
		.dout(new_net_18224)
	);

	bfr new_net_18225_bfr_after (
		.din(new_net_18224),
		.dout(new_net_18225)
	);

	bfr new_net_18226_bfr_after (
		.din(new_net_18225),
		.dout(new_net_18226)
	);

	bfr new_net_18227_bfr_after (
		.din(new_net_18226),
		.dout(new_net_18227)
	);

	bfr new_net_18228_bfr_after (
		.din(new_net_18227),
		.dout(new_net_18228)
	);

	bfr new_net_18229_bfr_after (
		.din(new_net_18228),
		.dout(new_net_18229)
	);

	bfr new_net_18230_bfr_after (
		.din(new_net_18229),
		.dout(new_net_18230)
	);

	bfr new_net_18231_bfr_after (
		.din(new_net_18230),
		.dout(new_net_18231)
	);

	bfr new_net_18232_bfr_after (
		.din(new_net_18231),
		.dout(new_net_18232)
	);

	bfr new_net_18233_bfr_after (
		.din(new_net_18232),
		.dout(new_net_18233)
	);

	bfr new_net_18234_bfr_after (
		.din(new_net_18233),
		.dout(new_net_18234)
	);

	bfr new_net_18235_bfr_after (
		.din(new_net_18234),
		.dout(new_net_18235)
	);

	bfr new_net_18236_bfr_after (
		.din(new_net_18235),
		.dout(new_net_18236)
	);

	bfr new_net_18237_bfr_after (
		.din(new_net_18236),
		.dout(new_net_18237)
	);

	bfr new_net_18238_bfr_after (
		.din(new_net_18237),
		.dout(new_net_18238)
	);

	bfr new_net_18239_bfr_after (
		.din(new_net_18238),
		.dout(new_net_18239)
	);

	bfr new_net_18240_bfr_after (
		.din(new_net_18239),
		.dout(new_net_18240)
	);

	spl2 _0093__v_fanout (
		.a(new_net_18240),
		.b(new_net_3045),
		.c(new_net_3046)
	);

	bfr new_net_18241_bfr_after (
		.din(_1003_),
		.dout(new_net_18241)
	);

	bfr new_net_18242_bfr_after (
		.din(new_net_18241),
		.dout(new_net_18242)
	);

	bfr new_net_18243_bfr_after (
		.din(new_net_18242),
		.dout(new_net_18243)
	);

	bfr new_net_18244_bfr_after (
		.din(new_net_18243),
		.dout(new_net_18244)
	);

	bfr new_net_18245_bfr_after (
		.din(new_net_18244),
		.dout(new_net_18245)
	);

	bfr new_net_18246_bfr_after (
		.din(new_net_18245),
		.dout(new_net_18246)
	);

	bfr new_net_18247_bfr_after (
		.din(new_net_18246),
		.dout(new_net_18247)
	);

	bfr new_net_18248_bfr_after (
		.din(new_net_18247),
		.dout(new_net_18248)
	);

	bfr new_net_18249_bfr_after (
		.din(new_net_18248),
		.dout(new_net_18249)
	);

	bfr new_net_18250_bfr_after (
		.din(new_net_18249),
		.dout(new_net_18250)
	);

	bfr new_net_18251_bfr_after (
		.din(new_net_18250),
		.dout(new_net_18251)
	);

	bfr new_net_18252_bfr_after (
		.din(new_net_18251),
		.dout(new_net_18252)
	);

	bfr new_net_18253_bfr_after (
		.din(new_net_18252),
		.dout(new_net_18253)
	);

	bfr new_net_18254_bfr_after (
		.din(new_net_18253),
		.dout(new_net_18254)
	);

	bfr new_net_18255_bfr_after (
		.din(new_net_18254),
		.dout(new_net_18255)
	);

	bfr new_net_18256_bfr_after (
		.din(new_net_18255),
		.dout(new_net_18256)
	);

	bfr new_net_18257_bfr_after (
		.din(new_net_18256),
		.dout(new_net_18257)
	);

	bfr new_net_18258_bfr_after (
		.din(new_net_18257),
		.dout(new_net_18258)
	);

	bfr new_net_18259_bfr_after (
		.din(new_net_18258),
		.dout(new_net_18259)
	);

	bfr new_net_18260_bfr_after (
		.din(new_net_18259),
		.dout(new_net_18260)
	);

	bfr new_net_18261_bfr_after (
		.din(new_net_18260),
		.dout(new_net_18261)
	);

	bfr new_net_18262_bfr_after (
		.din(new_net_18261),
		.dout(new_net_18262)
	);

	bfr new_net_18263_bfr_after (
		.din(new_net_18262),
		.dout(new_net_18263)
	);

	bfr new_net_18264_bfr_after (
		.din(new_net_18263),
		.dout(new_net_18264)
	);

	bfr new_net_18265_bfr_after (
		.din(new_net_18264),
		.dout(new_net_18265)
	);

	bfr new_net_18266_bfr_after (
		.din(new_net_18265),
		.dout(new_net_18266)
	);

	bfr new_net_18267_bfr_after (
		.din(new_net_18266),
		.dout(new_net_18267)
	);

	bfr new_net_18268_bfr_after (
		.din(new_net_18267),
		.dout(new_net_18268)
	);

	bfr new_net_18269_bfr_after (
		.din(new_net_18268),
		.dout(new_net_18269)
	);

	bfr new_net_18270_bfr_after (
		.din(new_net_18269),
		.dout(new_net_18270)
	);

	bfr new_net_18271_bfr_after (
		.din(new_net_18270),
		.dout(new_net_18271)
	);

	bfr new_net_18272_bfr_after (
		.din(new_net_18271),
		.dout(new_net_18272)
	);

	bfr new_net_18273_bfr_after (
		.din(new_net_18272),
		.dout(new_net_18273)
	);

	bfr new_net_18274_bfr_after (
		.din(new_net_18273),
		.dout(new_net_18274)
	);

	bfr new_net_18275_bfr_after (
		.din(new_net_18274),
		.dout(new_net_18275)
	);

	bfr new_net_18276_bfr_after (
		.din(new_net_18275),
		.dout(new_net_18276)
	);

	bfr new_net_18277_bfr_after (
		.din(new_net_18276),
		.dout(new_net_18277)
	);

	bfr new_net_18278_bfr_after (
		.din(new_net_18277),
		.dout(new_net_18278)
	);

	bfr new_net_18279_bfr_after (
		.din(new_net_18278),
		.dout(new_net_18279)
	);

	bfr new_net_18280_bfr_after (
		.din(new_net_18279),
		.dout(new_net_18280)
	);

	bfr new_net_18281_bfr_after (
		.din(new_net_18280),
		.dout(new_net_18281)
	);

	bfr new_net_18282_bfr_after (
		.din(new_net_18281),
		.dout(new_net_18282)
	);

	bfr new_net_18283_bfr_after (
		.din(new_net_18282),
		.dout(new_net_18283)
	);

	bfr new_net_18284_bfr_after (
		.din(new_net_18283),
		.dout(new_net_18284)
	);

	bfr new_net_18285_bfr_after (
		.din(new_net_18284),
		.dout(new_net_18285)
	);

	bfr new_net_18286_bfr_after (
		.din(new_net_18285),
		.dout(new_net_18286)
	);

	bfr new_net_18287_bfr_after (
		.din(new_net_18286),
		.dout(new_net_18287)
	);

	bfr new_net_18288_bfr_after (
		.din(new_net_18287),
		.dout(new_net_18288)
	);

	bfr new_net_18289_bfr_after (
		.din(new_net_18288),
		.dout(new_net_18289)
	);

	bfr new_net_18290_bfr_after (
		.din(new_net_18289),
		.dout(new_net_18290)
	);

	bfr new_net_18291_bfr_after (
		.din(new_net_18290),
		.dout(new_net_18291)
	);

	bfr new_net_18292_bfr_after (
		.din(new_net_18291),
		.dout(new_net_18292)
	);

	bfr new_net_18293_bfr_after (
		.din(new_net_18292),
		.dout(new_net_18293)
	);

	bfr new_net_18294_bfr_after (
		.din(new_net_18293),
		.dout(new_net_18294)
	);

	bfr new_net_18295_bfr_after (
		.din(new_net_18294),
		.dout(new_net_18295)
	);

	bfr new_net_18296_bfr_after (
		.din(new_net_18295),
		.dout(new_net_18296)
	);

	bfr new_net_18297_bfr_after (
		.din(new_net_18296),
		.dout(new_net_18297)
	);

	bfr new_net_18298_bfr_after (
		.din(new_net_18297),
		.dout(new_net_18298)
	);

	bfr new_net_18299_bfr_after (
		.din(new_net_18298),
		.dout(new_net_18299)
	);

	bfr new_net_18300_bfr_after (
		.din(new_net_18299),
		.dout(new_net_18300)
	);

	bfr new_net_18301_bfr_after (
		.din(new_net_18300),
		.dout(new_net_18301)
	);

	bfr new_net_18302_bfr_after (
		.din(new_net_18301),
		.dout(new_net_18302)
	);

	bfr new_net_18303_bfr_after (
		.din(new_net_18302),
		.dout(new_net_18303)
	);

	bfr new_net_18304_bfr_after (
		.din(new_net_18303),
		.dout(new_net_18304)
	);

	bfr new_net_18305_bfr_after (
		.din(new_net_18304),
		.dout(new_net_18305)
	);

	bfr new_net_18306_bfr_after (
		.din(new_net_18305),
		.dout(new_net_18306)
	);

	bfr new_net_18307_bfr_after (
		.din(new_net_18306),
		.dout(new_net_18307)
	);

	bfr new_net_18308_bfr_after (
		.din(new_net_18307),
		.dout(new_net_18308)
	);

	bfr new_net_18309_bfr_after (
		.din(new_net_18308),
		.dout(new_net_18309)
	);

	bfr new_net_18310_bfr_after (
		.din(new_net_18309),
		.dout(new_net_18310)
	);

	bfr new_net_18311_bfr_after (
		.din(new_net_18310),
		.dout(new_net_18311)
	);

	bfr new_net_18312_bfr_after (
		.din(new_net_18311),
		.dout(new_net_18312)
	);

	bfr new_net_18313_bfr_after (
		.din(new_net_18312),
		.dout(new_net_18313)
	);

	bfr new_net_18314_bfr_after (
		.din(new_net_18313),
		.dout(new_net_18314)
	);

	bfr new_net_18315_bfr_after (
		.din(new_net_18314),
		.dout(new_net_18315)
	);

	bfr new_net_18316_bfr_after (
		.din(new_net_18315),
		.dout(new_net_18316)
	);

	bfr new_net_18317_bfr_after (
		.din(new_net_18316),
		.dout(new_net_18317)
	);

	bfr new_net_18318_bfr_after (
		.din(new_net_18317),
		.dout(new_net_18318)
	);

	bfr new_net_18319_bfr_after (
		.din(new_net_18318),
		.dout(new_net_18319)
	);

	bfr new_net_18320_bfr_after (
		.din(new_net_18319),
		.dout(new_net_18320)
	);

	bfr new_net_18321_bfr_after (
		.din(new_net_18320),
		.dout(new_net_18321)
	);

	bfr new_net_18322_bfr_after (
		.din(new_net_18321),
		.dout(new_net_18322)
	);

	bfr new_net_18323_bfr_after (
		.din(new_net_18322),
		.dout(new_net_18323)
	);

	bfr new_net_18324_bfr_after (
		.din(new_net_18323),
		.dout(new_net_18324)
	);

	bfr new_net_18325_bfr_after (
		.din(new_net_18324),
		.dout(new_net_18325)
	);

	bfr new_net_18326_bfr_after (
		.din(new_net_18325),
		.dout(new_net_18326)
	);

	bfr new_net_18327_bfr_after (
		.din(new_net_18326),
		.dout(new_net_18327)
	);

	bfr new_net_18328_bfr_after (
		.din(new_net_18327),
		.dout(new_net_18328)
	);

	bfr new_net_18329_bfr_after (
		.din(new_net_18328),
		.dout(new_net_18329)
	);

	bfr new_net_18330_bfr_after (
		.din(new_net_18329),
		.dout(new_net_18330)
	);

	bfr new_net_18331_bfr_after (
		.din(new_net_18330),
		.dout(new_net_18331)
	);

	bfr new_net_18332_bfr_after (
		.din(new_net_18331),
		.dout(new_net_18332)
	);

	bfr new_net_18333_bfr_after (
		.din(new_net_18332),
		.dout(new_net_18333)
	);

	bfr new_net_18334_bfr_after (
		.din(new_net_18333),
		.dout(new_net_18334)
	);

	bfr new_net_18335_bfr_after (
		.din(new_net_18334),
		.dout(new_net_18335)
	);

	bfr new_net_18336_bfr_after (
		.din(new_net_18335),
		.dout(new_net_18336)
	);

	bfr new_net_18337_bfr_after (
		.din(new_net_18336),
		.dout(new_net_18337)
	);

	bfr new_net_18338_bfr_after (
		.din(new_net_18337),
		.dout(new_net_18338)
	);

	bfr new_net_18339_bfr_after (
		.din(new_net_18338),
		.dout(new_net_18339)
	);

	bfr new_net_18340_bfr_after (
		.din(new_net_18339),
		.dout(new_net_18340)
	);

	bfr new_net_18341_bfr_after (
		.din(new_net_18340),
		.dout(new_net_18341)
	);

	bfr new_net_18342_bfr_after (
		.din(new_net_18341),
		.dout(new_net_18342)
	);

	bfr new_net_18343_bfr_after (
		.din(new_net_18342),
		.dout(new_net_18343)
	);

	bfr new_net_18344_bfr_after (
		.din(new_net_18343),
		.dout(new_net_18344)
	);

	bfr new_net_18345_bfr_after (
		.din(new_net_18344),
		.dout(new_net_18345)
	);

	bfr new_net_18346_bfr_after (
		.din(new_net_18345),
		.dout(new_net_18346)
	);

	bfr new_net_18347_bfr_after (
		.din(new_net_18346),
		.dout(new_net_18347)
	);

	bfr new_net_18348_bfr_after (
		.din(new_net_18347),
		.dout(new_net_18348)
	);

	bfr new_net_18349_bfr_after (
		.din(new_net_18348),
		.dout(new_net_18349)
	);

	bfr new_net_18350_bfr_after (
		.din(new_net_18349),
		.dout(new_net_18350)
	);

	spl2 _1003__v_fanout (
		.a(new_net_18350),
		.b(new_net_1664),
		.c(new_net_1665)
	);

	bfr new_net_18351_bfr_after (
		.din(_1078_),
		.dout(new_net_18351)
	);

	bfr new_net_18352_bfr_after (
		.din(new_net_18351),
		.dout(new_net_18352)
	);

	bfr new_net_18353_bfr_after (
		.din(new_net_18352),
		.dout(new_net_18353)
	);

	bfr new_net_18354_bfr_after (
		.din(new_net_18353),
		.dout(new_net_18354)
	);

	bfr new_net_18355_bfr_after (
		.din(new_net_18354),
		.dout(new_net_18355)
	);

	bfr new_net_18356_bfr_after (
		.din(new_net_18355),
		.dout(new_net_18356)
	);

	bfr new_net_18357_bfr_after (
		.din(new_net_18356),
		.dout(new_net_18357)
	);

	bfr new_net_18358_bfr_after (
		.din(new_net_18357),
		.dout(new_net_18358)
	);

	bfr new_net_18359_bfr_after (
		.din(new_net_18358),
		.dout(new_net_18359)
	);

	bfr new_net_18360_bfr_after (
		.din(new_net_18359),
		.dout(new_net_18360)
	);

	bfr new_net_18361_bfr_after (
		.din(new_net_18360),
		.dout(new_net_18361)
	);

	bfr new_net_18362_bfr_after (
		.din(new_net_18361),
		.dout(new_net_18362)
	);

	bfr new_net_18363_bfr_after (
		.din(new_net_18362),
		.dout(new_net_18363)
	);

	bfr new_net_18364_bfr_after (
		.din(new_net_18363),
		.dout(new_net_18364)
	);

	bfr new_net_18365_bfr_after (
		.din(new_net_18364),
		.dout(new_net_18365)
	);

	bfr new_net_18366_bfr_after (
		.din(new_net_18365),
		.dout(new_net_18366)
	);

	bfr new_net_18367_bfr_after (
		.din(new_net_18366),
		.dout(new_net_18367)
	);

	bfr new_net_18368_bfr_after (
		.din(new_net_18367),
		.dout(new_net_18368)
	);

	bfr new_net_18369_bfr_after (
		.din(new_net_18368),
		.dout(new_net_18369)
	);

	bfr new_net_18370_bfr_after (
		.din(new_net_18369),
		.dout(new_net_18370)
	);

	bfr new_net_18371_bfr_after (
		.din(new_net_18370),
		.dout(new_net_18371)
	);

	bfr new_net_18372_bfr_after (
		.din(new_net_18371),
		.dout(new_net_18372)
	);

	bfr new_net_18373_bfr_after (
		.din(new_net_18372),
		.dout(new_net_18373)
	);

	bfr new_net_18374_bfr_after (
		.din(new_net_18373),
		.dout(new_net_18374)
	);

	bfr new_net_18375_bfr_after (
		.din(new_net_18374),
		.dout(new_net_18375)
	);

	spl2 _1078__v_fanout (
		.a(new_net_18375),
		.b(new_net_1261),
		.c(new_net_1262)
	);

	bfr new_net_18376_bfr_after (
		.din(_1136_),
		.dout(new_net_18376)
	);

	bfr new_net_18377_bfr_after (
		.din(new_net_18376),
		.dout(new_net_18377)
	);

	bfr new_net_18378_bfr_after (
		.din(new_net_18377),
		.dout(new_net_18378)
	);

	bfr new_net_18379_bfr_after (
		.din(new_net_18378),
		.dout(new_net_18379)
	);

	bfr new_net_18380_bfr_after (
		.din(new_net_18379),
		.dout(new_net_18380)
	);

	bfr new_net_18381_bfr_after (
		.din(new_net_18380),
		.dout(new_net_18381)
	);

	bfr new_net_18382_bfr_after (
		.din(new_net_18381),
		.dout(new_net_18382)
	);

	bfr new_net_18383_bfr_after (
		.din(new_net_18382),
		.dout(new_net_18383)
	);

	bfr new_net_18384_bfr_after (
		.din(new_net_18383),
		.dout(new_net_18384)
	);

	bfr new_net_18385_bfr_after (
		.din(new_net_18384),
		.dout(new_net_18385)
	);

	bfr new_net_18386_bfr_after (
		.din(new_net_18385),
		.dout(new_net_18386)
	);

	bfr new_net_18387_bfr_after (
		.din(new_net_18386),
		.dout(new_net_18387)
	);

	bfr new_net_18388_bfr_after (
		.din(new_net_18387),
		.dout(new_net_18388)
	);

	bfr new_net_18389_bfr_after (
		.din(new_net_18388),
		.dout(new_net_18389)
	);

	bfr new_net_18390_bfr_after (
		.din(new_net_18389),
		.dout(new_net_18390)
	);

	bfr new_net_18391_bfr_after (
		.din(new_net_18390),
		.dout(new_net_18391)
	);

	bfr new_net_18392_bfr_after (
		.din(new_net_18391),
		.dout(new_net_18392)
	);

	bfr new_net_18393_bfr_after (
		.din(new_net_18392),
		.dout(new_net_18393)
	);

	bfr new_net_18394_bfr_after (
		.din(new_net_18393),
		.dout(new_net_18394)
	);

	bfr new_net_18395_bfr_after (
		.din(new_net_18394),
		.dout(new_net_18395)
	);

	bfr new_net_18396_bfr_after (
		.din(new_net_18395),
		.dout(new_net_18396)
	);

	bfr new_net_18397_bfr_after (
		.din(new_net_18396),
		.dout(new_net_18397)
	);

	bfr new_net_18398_bfr_after (
		.din(new_net_18397),
		.dout(new_net_18398)
	);

	bfr new_net_18399_bfr_after (
		.din(new_net_18398),
		.dout(new_net_18399)
	);

	bfr new_net_18400_bfr_after (
		.din(new_net_18399),
		.dout(new_net_18400)
	);

	bfr new_net_18401_bfr_after (
		.din(new_net_18400),
		.dout(new_net_18401)
	);

	bfr new_net_18402_bfr_after (
		.din(new_net_18401),
		.dout(new_net_18402)
	);

	bfr new_net_18403_bfr_after (
		.din(new_net_18402),
		.dout(new_net_18403)
	);

	bfr new_net_18404_bfr_after (
		.din(new_net_18403),
		.dout(new_net_18404)
	);

	bfr new_net_18405_bfr_after (
		.din(new_net_18404),
		.dout(new_net_18405)
	);

	bfr new_net_18406_bfr_after (
		.din(new_net_18405),
		.dout(new_net_18406)
	);

	bfr new_net_18407_bfr_after (
		.din(new_net_18406),
		.dout(new_net_18407)
	);

	bfr new_net_18408_bfr_after (
		.din(new_net_18407),
		.dout(new_net_18408)
	);

	spl2 _1136__v_fanout (
		.a(new_net_18408),
		.b(new_net_1110),
		.c(new_net_1111)
	);

	bfr new_net_18409_bfr_after (
		.din(_1211_),
		.dout(new_net_18409)
	);

	bfr new_net_18410_bfr_after (
		.din(new_net_18409),
		.dout(new_net_18410)
	);

	bfr new_net_18411_bfr_after (
		.din(new_net_18410),
		.dout(new_net_18411)
	);

	bfr new_net_18412_bfr_after (
		.din(new_net_18411),
		.dout(new_net_18412)
	);

	bfr new_net_18413_bfr_after (
		.din(new_net_18412),
		.dout(new_net_18413)
	);

	bfr new_net_18414_bfr_after (
		.din(new_net_18413),
		.dout(new_net_18414)
	);

	bfr new_net_18415_bfr_after (
		.din(new_net_18414),
		.dout(new_net_18415)
	);

	bfr new_net_18416_bfr_after (
		.din(new_net_18415),
		.dout(new_net_18416)
	);

	bfr new_net_18417_bfr_after (
		.din(new_net_18416),
		.dout(new_net_18417)
	);

	bfr new_net_18418_bfr_after (
		.din(new_net_18417),
		.dout(new_net_18418)
	);

	bfr new_net_18419_bfr_after (
		.din(new_net_18418),
		.dout(new_net_18419)
	);

	bfr new_net_18420_bfr_after (
		.din(new_net_18419),
		.dout(new_net_18420)
	);

	bfr new_net_18421_bfr_after (
		.din(new_net_18420),
		.dout(new_net_18421)
	);

	bfr new_net_18422_bfr_after (
		.din(new_net_18421),
		.dout(new_net_18422)
	);

	bfr new_net_18423_bfr_after (
		.din(new_net_18422),
		.dout(new_net_18423)
	);

	bfr new_net_18424_bfr_after (
		.din(new_net_18423),
		.dout(new_net_18424)
	);

	bfr new_net_18425_bfr_after (
		.din(new_net_18424),
		.dout(new_net_18425)
	);

	bfr new_net_18426_bfr_after (
		.din(new_net_18425),
		.dout(new_net_18426)
	);

	bfr new_net_18427_bfr_after (
		.din(new_net_18426),
		.dout(new_net_18427)
	);

	bfr new_net_18428_bfr_after (
		.din(new_net_18427),
		.dout(new_net_18428)
	);

	bfr new_net_18429_bfr_after (
		.din(new_net_18428),
		.dout(new_net_18429)
	);

	bfr new_net_18430_bfr_after (
		.din(new_net_18429),
		.dout(new_net_18430)
	);

	bfr new_net_18431_bfr_after (
		.din(new_net_18430),
		.dout(new_net_18431)
	);

	bfr new_net_18432_bfr_after (
		.din(new_net_18431),
		.dout(new_net_18432)
	);

	bfr new_net_18433_bfr_after (
		.din(new_net_18432),
		.dout(new_net_18433)
	);

	bfr new_net_18434_bfr_after (
		.din(new_net_18433),
		.dout(new_net_18434)
	);

	bfr new_net_18435_bfr_after (
		.din(new_net_18434),
		.dout(new_net_18435)
	);

	bfr new_net_18436_bfr_after (
		.din(new_net_18435),
		.dout(new_net_18436)
	);

	bfr new_net_18437_bfr_after (
		.din(new_net_18436),
		.dout(new_net_18437)
	);

	bfr new_net_18438_bfr_after (
		.din(new_net_18437),
		.dout(new_net_18438)
	);

	bfr new_net_18439_bfr_after (
		.din(new_net_18438),
		.dout(new_net_18439)
	);

	bfr new_net_18440_bfr_after (
		.din(new_net_18439),
		.dout(new_net_18440)
	);

	bfr new_net_18441_bfr_after (
		.din(new_net_18440),
		.dout(new_net_18441)
	);

	bfr new_net_18442_bfr_after (
		.din(new_net_18441),
		.dout(new_net_18442)
	);

	bfr new_net_18443_bfr_after (
		.din(new_net_18442),
		.dout(new_net_18443)
	);

	bfr new_net_18444_bfr_after (
		.din(new_net_18443),
		.dout(new_net_18444)
	);

	bfr new_net_18445_bfr_after (
		.din(new_net_18444),
		.dout(new_net_18445)
	);

	bfr new_net_18446_bfr_after (
		.din(new_net_18445),
		.dout(new_net_18446)
	);

	bfr new_net_18447_bfr_after (
		.din(new_net_18446),
		.dout(new_net_18447)
	);

	bfr new_net_18448_bfr_after (
		.din(new_net_18447),
		.dout(new_net_18448)
	);

	bfr new_net_18449_bfr_after (
		.din(new_net_18448),
		.dout(new_net_18449)
	);

	spl2 _1211__v_fanout (
		.a(new_net_18449),
		.b(new_net_1212),
		.c(new_net_1213)
	);

	bfr new_net_18450_bfr_after (
		.din(_1687_),
		.dout(new_net_18450)
	);

	bfr new_net_18451_bfr_after (
		.din(new_net_18450),
		.dout(new_net_18451)
	);

	bfr new_net_18452_bfr_after (
		.din(new_net_18451),
		.dout(new_net_18452)
	);

	bfr new_net_18453_bfr_after (
		.din(new_net_18452),
		.dout(new_net_18453)
	);

	bfr new_net_18454_bfr_after (
		.din(new_net_18453),
		.dout(new_net_18454)
	);

	bfr new_net_18455_bfr_after (
		.din(new_net_18454),
		.dout(new_net_18455)
	);

	bfr new_net_18456_bfr_after (
		.din(new_net_18455),
		.dout(new_net_18456)
	);

	bfr new_net_18457_bfr_after (
		.din(new_net_18456),
		.dout(new_net_18457)
	);

	bfr new_net_18458_bfr_after (
		.din(new_net_18457),
		.dout(new_net_18458)
	);

	bfr new_net_18459_bfr_after (
		.din(new_net_18458),
		.dout(new_net_18459)
	);

	bfr new_net_18460_bfr_after (
		.din(new_net_18459),
		.dout(new_net_18460)
	);

	bfr new_net_18461_bfr_after (
		.din(new_net_18460),
		.dout(new_net_18461)
	);

	bfr new_net_18462_bfr_after (
		.din(new_net_18461),
		.dout(new_net_18462)
	);

	bfr new_net_18463_bfr_after (
		.din(new_net_18462),
		.dout(new_net_18463)
	);

	bfr new_net_18464_bfr_after (
		.din(new_net_18463),
		.dout(new_net_18464)
	);

	bfr new_net_18465_bfr_after (
		.din(new_net_18464),
		.dout(new_net_18465)
	);

	bfr new_net_18466_bfr_after (
		.din(new_net_18465),
		.dout(new_net_18466)
	);

	bfr new_net_18467_bfr_after (
		.din(new_net_18466),
		.dout(new_net_18467)
	);

	bfr new_net_18468_bfr_after (
		.din(new_net_18467),
		.dout(new_net_18468)
	);

	bfr new_net_18469_bfr_after (
		.din(new_net_18468),
		.dout(new_net_18469)
	);

	bfr new_net_18470_bfr_after (
		.din(new_net_18469),
		.dout(new_net_18470)
	);

	bfr new_net_18471_bfr_after (
		.din(new_net_18470),
		.dout(new_net_18471)
	);

	bfr new_net_18472_bfr_after (
		.din(new_net_18471),
		.dout(new_net_18472)
	);

	bfr new_net_18473_bfr_after (
		.din(new_net_18472),
		.dout(new_net_18473)
	);

	bfr new_net_18474_bfr_after (
		.din(new_net_18473),
		.dout(new_net_18474)
	);

	bfr new_net_18475_bfr_after (
		.din(new_net_18474),
		.dout(new_net_18475)
	);

	bfr new_net_18476_bfr_after (
		.din(new_net_18475),
		.dout(new_net_18476)
	);

	bfr new_net_18477_bfr_after (
		.din(new_net_18476),
		.dout(new_net_18477)
	);

	bfr new_net_18478_bfr_after (
		.din(new_net_18477),
		.dout(new_net_18478)
	);

	bfr new_net_18479_bfr_after (
		.din(new_net_18478),
		.dout(new_net_18479)
	);

	bfr new_net_18480_bfr_after (
		.din(new_net_18479),
		.dout(new_net_18480)
	);

	bfr new_net_18481_bfr_after (
		.din(new_net_18480),
		.dout(new_net_18481)
	);

	bfr new_net_18482_bfr_after (
		.din(new_net_18481),
		.dout(new_net_18482)
	);

	bfr new_net_18483_bfr_after (
		.din(new_net_18482),
		.dout(new_net_18483)
	);

	bfr new_net_18484_bfr_after (
		.din(new_net_18483),
		.dout(new_net_18484)
	);

	bfr new_net_18485_bfr_after (
		.din(new_net_18484),
		.dout(new_net_18485)
	);

	bfr new_net_18486_bfr_after (
		.din(new_net_18485),
		.dout(new_net_18486)
	);

	bfr new_net_18487_bfr_after (
		.din(new_net_18486),
		.dout(new_net_18487)
	);

	bfr new_net_18488_bfr_after (
		.din(new_net_18487),
		.dout(new_net_18488)
	);

	bfr new_net_18489_bfr_after (
		.din(new_net_18488),
		.dout(new_net_18489)
	);

	bfr new_net_18490_bfr_after (
		.din(new_net_18489),
		.dout(new_net_18490)
	);

	bfr new_net_18491_bfr_after (
		.din(new_net_18490),
		.dout(new_net_18491)
	);

	bfr new_net_18492_bfr_after (
		.din(new_net_18491),
		.dout(new_net_18492)
	);

	bfr new_net_18493_bfr_after (
		.din(new_net_18492),
		.dout(new_net_18493)
	);

	bfr new_net_18494_bfr_after (
		.din(new_net_18493),
		.dout(new_net_18494)
	);

	bfr new_net_18495_bfr_after (
		.din(new_net_18494),
		.dout(new_net_18495)
	);

	bfr new_net_18496_bfr_after (
		.din(new_net_18495),
		.dout(new_net_18496)
	);

	bfr new_net_18497_bfr_after (
		.din(new_net_18496),
		.dout(new_net_18497)
	);

	bfr new_net_18498_bfr_after (
		.din(new_net_18497),
		.dout(new_net_18498)
	);

	bfr new_net_18499_bfr_after (
		.din(new_net_18498),
		.dout(new_net_18499)
	);

	bfr new_net_18500_bfr_after (
		.din(new_net_18499),
		.dout(new_net_18500)
	);

	bfr new_net_18501_bfr_after (
		.din(new_net_18500),
		.dout(new_net_18501)
	);

	bfr new_net_18502_bfr_after (
		.din(new_net_18501),
		.dout(new_net_18502)
	);

	bfr new_net_18503_bfr_after (
		.din(new_net_18502),
		.dout(new_net_18503)
	);

	bfr new_net_18504_bfr_after (
		.din(new_net_18503),
		.dout(new_net_18504)
	);

	bfr new_net_18505_bfr_after (
		.din(new_net_18504),
		.dout(new_net_18505)
	);

	bfr new_net_18506_bfr_after (
		.din(new_net_18505),
		.dout(new_net_18506)
	);

	bfr new_net_18507_bfr_after (
		.din(new_net_18506),
		.dout(new_net_18507)
	);

	bfr new_net_18508_bfr_after (
		.din(new_net_18507),
		.dout(new_net_18508)
	);

	bfr new_net_18509_bfr_after (
		.din(new_net_18508),
		.dout(new_net_18509)
	);

	bfr new_net_18510_bfr_after (
		.din(new_net_18509),
		.dout(new_net_18510)
	);

	bfr new_net_18511_bfr_after (
		.din(new_net_18510),
		.dout(new_net_18511)
	);

	bfr new_net_18512_bfr_after (
		.din(new_net_18511),
		.dout(new_net_18512)
	);

	bfr new_net_18513_bfr_after (
		.din(new_net_18512),
		.dout(new_net_18513)
	);

	bfr new_net_18514_bfr_after (
		.din(new_net_18513),
		.dout(new_net_18514)
	);

	bfr new_net_18515_bfr_after (
		.din(new_net_18514),
		.dout(new_net_18515)
	);

	bfr new_net_18516_bfr_after (
		.din(new_net_18515),
		.dout(new_net_18516)
	);

	bfr new_net_18517_bfr_after (
		.din(new_net_18516),
		.dout(new_net_18517)
	);

	bfr new_net_18518_bfr_after (
		.din(new_net_18517),
		.dout(new_net_18518)
	);

	bfr new_net_18519_bfr_after (
		.din(new_net_18518),
		.dout(new_net_18519)
	);

	bfr new_net_18520_bfr_after (
		.din(new_net_18519),
		.dout(new_net_18520)
	);

	bfr new_net_18521_bfr_after (
		.din(new_net_18520),
		.dout(new_net_18521)
	);

	bfr new_net_18522_bfr_after (
		.din(new_net_18521),
		.dout(new_net_18522)
	);

	bfr new_net_18523_bfr_after (
		.din(new_net_18522),
		.dout(new_net_18523)
	);

	bfr new_net_18524_bfr_after (
		.din(new_net_18523),
		.dout(new_net_18524)
	);

	bfr new_net_18525_bfr_after (
		.din(new_net_18524),
		.dout(new_net_18525)
	);

	bfr new_net_18526_bfr_after (
		.din(new_net_18525),
		.dout(new_net_18526)
	);

	bfr new_net_18527_bfr_after (
		.din(new_net_18526),
		.dout(new_net_18527)
	);

	bfr new_net_18528_bfr_after (
		.din(new_net_18527),
		.dout(new_net_18528)
	);

	bfr new_net_18529_bfr_after (
		.din(new_net_18528),
		.dout(new_net_18529)
	);

	bfr new_net_18530_bfr_after (
		.din(new_net_18529),
		.dout(new_net_18530)
	);

	spl2 _1687__v_fanout (
		.a(new_net_18530),
		.b(new_net_190),
		.c(new_net_191)
	);

	bfr new_net_18531_bfr_after (
		.din(_0214_),
		.dout(new_net_18531)
	);

	bfr new_net_18532_bfr_after (
		.din(new_net_18531),
		.dout(new_net_18532)
	);

	bfr new_net_18533_bfr_after (
		.din(new_net_18532),
		.dout(new_net_18533)
	);

	bfr new_net_18534_bfr_after (
		.din(new_net_18533),
		.dout(new_net_18534)
	);

	bfr new_net_18535_bfr_after (
		.din(new_net_18534),
		.dout(new_net_18535)
	);

	bfr new_net_18536_bfr_after (
		.din(new_net_18535),
		.dout(new_net_18536)
	);

	bfr new_net_18537_bfr_after (
		.din(new_net_18536),
		.dout(new_net_18537)
	);

	bfr new_net_18538_bfr_after (
		.din(new_net_18537),
		.dout(new_net_18538)
	);

	bfr new_net_18539_bfr_after (
		.din(new_net_18538),
		.dout(new_net_18539)
	);

	bfr new_net_18540_bfr_after (
		.din(new_net_18539),
		.dout(new_net_18540)
	);

	bfr new_net_18541_bfr_after (
		.din(new_net_18540),
		.dout(new_net_18541)
	);

	bfr new_net_18542_bfr_after (
		.din(new_net_18541),
		.dout(new_net_18542)
	);

	bfr new_net_18543_bfr_after (
		.din(new_net_18542),
		.dout(new_net_18543)
	);

	bfr new_net_18544_bfr_after (
		.din(new_net_18543),
		.dout(new_net_18544)
	);

	bfr new_net_18545_bfr_after (
		.din(new_net_18544),
		.dout(new_net_18545)
	);

	bfr new_net_18546_bfr_after (
		.din(new_net_18545),
		.dout(new_net_18546)
	);

	bfr new_net_18547_bfr_after (
		.din(new_net_18546),
		.dout(new_net_18547)
	);

	bfr new_net_18548_bfr_after (
		.din(new_net_18547),
		.dout(new_net_18548)
	);

	bfr new_net_18549_bfr_after (
		.din(new_net_18548),
		.dout(new_net_18549)
	);

	bfr new_net_18550_bfr_after (
		.din(new_net_18549),
		.dout(new_net_18550)
	);

	bfr new_net_18551_bfr_after (
		.din(new_net_18550),
		.dout(new_net_18551)
	);

	bfr new_net_18552_bfr_after (
		.din(new_net_18551),
		.dout(new_net_18552)
	);

	bfr new_net_18553_bfr_after (
		.din(new_net_18552),
		.dout(new_net_18553)
	);

	bfr new_net_18554_bfr_after (
		.din(new_net_18553),
		.dout(new_net_18554)
	);

	bfr new_net_18555_bfr_after (
		.din(new_net_18554),
		.dout(new_net_18555)
	);

	bfr new_net_18556_bfr_after (
		.din(new_net_18555),
		.dout(new_net_18556)
	);

	bfr new_net_18557_bfr_after (
		.din(new_net_18556),
		.dout(new_net_18557)
	);

	bfr new_net_18558_bfr_after (
		.din(new_net_18557),
		.dout(new_net_18558)
	);

	bfr new_net_18559_bfr_after (
		.din(new_net_18558),
		.dout(new_net_18559)
	);

	bfr new_net_18560_bfr_after (
		.din(new_net_18559),
		.dout(new_net_18560)
	);

	bfr new_net_18561_bfr_after (
		.din(new_net_18560),
		.dout(new_net_18561)
	);

	bfr new_net_18562_bfr_after (
		.din(new_net_18561),
		.dout(new_net_18562)
	);

	bfr new_net_18563_bfr_after (
		.din(new_net_18562),
		.dout(new_net_18563)
	);

	bfr new_net_18564_bfr_after (
		.din(new_net_18563),
		.dout(new_net_18564)
	);

	bfr new_net_18565_bfr_after (
		.din(new_net_18564),
		.dout(new_net_18565)
	);

	bfr new_net_18566_bfr_after (
		.din(new_net_18565),
		.dout(new_net_18566)
	);

	bfr new_net_18567_bfr_after (
		.din(new_net_18566),
		.dout(new_net_18567)
	);

	bfr new_net_18568_bfr_after (
		.din(new_net_18567),
		.dout(new_net_18568)
	);

	bfr new_net_18569_bfr_after (
		.din(new_net_18568),
		.dout(new_net_18569)
	);

	bfr new_net_18570_bfr_after (
		.din(new_net_18569),
		.dout(new_net_18570)
	);

	bfr new_net_18571_bfr_after (
		.din(new_net_18570),
		.dout(new_net_18571)
	);

	bfr new_net_18572_bfr_after (
		.din(new_net_18571),
		.dout(new_net_18572)
	);

	bfr new_net_18573_bfr_after (
		.din(new_net_18572),
		.dout(new_net_18573)
	);

	bfr new_net_18574_bfr_after (
		.din(new_net_18573),
		.dout(new_net_18574)
	);

	bfr new_net_18575_bfr_after (
		.din(new_net_18574),
		.dout(new_net_18575)
	);

	bfr new_net_18576_bfr_after (
		.din(new_net_18575),
		.dout(new_net_18576)
	);

	bfr new_net_18577_bfr_after (
		.din(new_net_18576),
		.dout(new_net_18577)
	);

	bfr new_net_18578_bfr_after (
		.din(new_net_18577),
		.dout(new_net_18578)
	);

	bfr new_net_18579_bfr_after (
		.din(new_net_18578),
		.dout(new_net_18579)
	);

	bfr new_net_18580_bfr_after (
		.din(new_net_18579),
		.dout(new_net_18580)
	);

	bfr new_net_18581_bfr_after (
		.din(new_net_18580),
		.dout(new_net_18581)
	);

	bfr new_net_18582_bfr_after (
		.din(new_net_18581),
		.dout(new_net_18582)
	);

	bfr new_net_18583_bfr_after (
		.din(new_net_18582),
		.dout(new_net_18583)
	);

	bfr new_net_18584_bfr_after (
		.din(new_net_18583),
		.dout(new_net_18584)
	);

	bfr new_net_18585_bfr_after (
		.din(new_net_18584),
		.dout(new_net_18585)
	);

	bfr new_net_18586_bfr_after (
		.din(new_net_18585),
		.dout(new_net_18586)
	);

	bfr new_net_18587_bfr_after (
		.din(new_net_18586),
		.dout(new_net_18587)
	);

	bfr new_net_18588_bfr_after (
		.din(new_net_18587),
		.dout(new_net_18588)
	);

	bfr new_net_18589_bfr_after (
		.din(new_net_18588),
		.dout(new_net_18589)
	);

	bfr new_net_18590_bfr_after (
		.din(new_net_18589),
		.dout(new_net_18590)
	);

	bfr new_net_18591_bfr_after (
		.din(new_net_18590),
		.dout(new_net_18591)
	);

	bfr new_net_18592_bfr_after (
		.din(new_net_18591),
		.dout(new_net_18592)
	);

	bfr new_net_18593_bfr_after (
		.din(new_net_18592),
		.dout(new_net_18593)
	);

	bfr new_net_18594_bfr_after (
		.din(new_net_18593),
		.dout(new_net_18594)
	);

	bfr new_net_18595_bfr_after (
		.din(new_net_18594),
		.dout(new_net_18595)
	);

	bfr new_net_18596_bfr_after (
		.din(new_net_18595),
		.dout(new_net_18596)
	);

	bfr new_net_18597_bfr_after (
		.din(new_net_18596),
		.dout(new_net_18597)
	);

	bfr new_net_18598_bfr_after (
		.din(new_net_18597),
		.dout(new_net_18598)
	);

	bfr new_net_18599_bfr_after (
		.din(new_net_18598),
		.dout(new_net_18599)
	);

	bfr new_net_18600_bfr_after (
		.din(new_net_18599),
		.dout(new_net_18600)
	);

	bfr new_net_18601_bfr_after (
		.din(new_net_18600),
		.dout(new_net_18601)
	);

	bfr new_net_18602_bfr_after (
		.din(new_net_18601),
		.dout(new_net_18602)
	);

	bfr new_net_18603_bfr_after (
		.din(new_net_18602),
		.dout(new_net_18603)
	);

	bfr new_net_18604_bfr_after (
		.din(new_net_18603),
		.dout(new_net_18604)
	);

	bfr new_net_18605_bfr_after (
		.din(new_net_18604),
		.dout(new_net_18605)
	);

	bfr new_net_18606_bfr_after (
		.din(new_net_18605),
		.dout(new_net_18606)
	);

	bfr new_net_18607_bfr_after (
		.din(new_net_18606),
		.dout(new_net_18607)
	);

	bfr new_net_18608_bfr_after (
		.din(new_net_18607),
		.dout(new_net_18608)
	);

	bfr new_net_18609_bfr_after (
		.din(new_net_18608),
		.dout(new_net_18609)
	);

	bfr new_net_18610_bfr_after (
		.din(new_net_18609),
		.dout(new_net_18610)
	);

	bfr new_net_18611_bfr_after (
		.din(new_net_18610),
		.dout(new_net_18611)
	);

	bfr new_net_18612_bfr_after (
		.din(new_net_18611),
		.dout(new_net_18612)
	);

	bfr new_net_18613_bfr_after (
		.din(new_net_18612),
		.dout(new_net_18613)
	);

	bfr new_net_18614_bfr_after (
		.din(new_net_18613),
		.dout(new_net_18614)
	);

	bfr new_net_18615_bfr_after (
		.din(new_net_18614),
		.dout(new_net_18615)
	);

	bfr new_net_18616_bfr_after (
		.din(new_net_18615),
		.dout(new_net_18616)
	);

	bfr new_net_18617_bfr_after (
		.din(new_net_18616),
		.dout(new_net_18617)
	);

	bfr new_net_18618_bfr_after (
		.din(new_net_18617),
		.dout(new_net_18618)
	);

	bfr new_net_18619_bfr_after (
		.din(new_net_18618),
		.dout(new_net_18619)
	);

	bfr new_net_18620_bfr_after (
		.din(new_net_18619),
		.dout(new_net_18620)
	);

	bfr new_net_18621_bfr_after (
		.din(new_net_18620),
		.dout(new_net_18621)
	);

	bfr new_net_18622_bfr_after (
		.din(new_net_18621),
		.dout(new_net_18622)
	);

	bfr new_net_18623_bfr_after (
		.din(new_net_18622),
		.dout(new_net_18623)
	);

	bfr new_net_18624_bfr_after (
		.din(new_net_18623),
		.dout(new_net_18624)
	);

	bfr new_net_18625_bfr_after (
		.din(new_net_18624),
		.dout(new_net_18625)
	);

	bfr new_net_18626_bfr_after (
		.din(new_net_18625),
		.dout(new_net_18626)
	);

	bfr new_net_18627_bfr_after (
		.din(new_net_18626),
		.dout(new_net_18627)
	);

	bfr new_net_18628_bfr_after (
		.din(new_net_18627),
		.dout(new_net_18628)
	);

	bfr new_net_18629_bfr_after (
		.din(new_net_18628),
		.dout(new_net_18629)
	);

	bfr new_net_18630_bfr_after (
		.din(new_net_18629),
		.dout(new_net_18630)
	);

	bfr new_net_18631_bfr_after (
		.din(new_net_18630),
		.dout(new_net_18631)
	);

	bfr new_net_18632_bfr_after (
		.din(new_net_18631),
		.dout(new_net_18632)
	);

	bfr new_net_18633_bfr_after (
		.din(new_net_18632),
		.dout(new_net_18633)
	);

	bfr new_net_18634_bfr_after (
		.din(new_net_18633),
		.dout(new_net_18634)
	);

	bfr new_net_18635_bfr_after (
		.din(new_net_18634),
		.dout(new_net_18635)
	);

	spl2 _0214__v_fanout (
		.a(new_net_18635),
		.b(new_net_2815),
		.c(new_net_2816)
	);

	bfr new_net_18636_bfr_after (
		.din(_1569_),
		.dout(new_net_18636)
	);

	bfr new_net_18637_bfr_after (
		.din(new_net_18636),
		.dout(new_net_18637)
	);

	bfr new_net_18638_bfr_after (
		.din(new_net_18637),
		.dout(new_net_18638)
	);

	bfr new_net_18639_bfr_after (
		.din(new_net_18638),
		.dout(new_net_18639)
	);

	bfr new_net_18640_bfr_after (
		.din(new_net_18639),
		.dout(new_net_18640)
	);

	bfr new_net_18641_bfr_after (
		.din(new_net_18640),
		.dout(new_net_18641)
	);

	bfr new_net_18642_bfr_after (
		.din(new_net_18641),
		.dout(new_net_18642)
	);

	bfr new_net_18643_bfr_after (
		.din(new_net_18642),
		.dout(new_net_18643)
	);

	bfr new_net_18644_bfr_after (
		.din(new_net_18643),
		.dout(new_net_18644)
	);

	bfr new_net_18645_bfr_after (
		.din(new_net_18644),
		.dout(new_net_18645)
	);

	bfr new_net_18646_bfr_after (
		.din(new_net_18645),
		.dout(new_net_18646)
	);

	bfr new_net_18647_bfr_after (
		.din(new_net_18646),
		.dout(new_net_18647)
	);

	bfr new_net_18648_bfr_after (
		.din(new_net_18647),
		.dout(new_net_18648)
	);

	bfr new_net_18649_bfr_after (
		.din(new_net_18648),
		.dout(new_net_18649)
	);

	bfr new_net_18650_bfr_after (
		.din(new_net_18649),
		.dout(new_net_18650)
	);

	bfr new_net_18651_bfr_after (
		.din(new_net_18650),
		.dout(new_net_18651)
	);

	bfr new_net_18652_bfr_after (
		.din(new_net_18651),
		.dout(new_net_18652)
	);

	bfr new_net_18653_bfr_after (
		.din(new_net_18652),
		.dout(new_net_18653)
	);

	bfr new_net_18654_bfr_after (
		.din(new_net_18653),
		.dout(new_net_18654)
	);

	bfr new_net_18655_bfr_after (
		.din(new_net_18654),
		.dout(new_net_18655)
	);

	bfr new_net_18656_bfr_after (
		.din(new_net_18655),
		.dout(new_net_18656)
	);

	bfr new_net_18657_bfr_after (
		.din(new_net_18656),
		.dout(new_net_18657)
	);

	bfr new_net_18658_bfr_after (
		.din(new_net_18657),
		.dout(new_net_18658)
	);

	bfr new_net_18659_bfr_after (
		.din(new_net_18658),
		.dout(new_net_18659)
	);

	bfr new_net_18660_bfr_after (
		.din(new_net_18659),
		.dout(new_net_18660)
	);

	bfr new_net_18661_bfr_after (
		.din(new_net_18660),
		.dout(new_net_18661)
	);

	bfr new_net_18662_bfr_after (
		.din(new_net_18661),
		.dout(new_net_18662)
	);

	bfr new_net_18663_bfr_after (
		.din(new_net_18662),
		.dout(new_net_18663)
	);

	bfr new_net_18664_bfr_after (
		.din(new_net_18663),
		.dout(new_net_18664)
	);

	bfr new_net_18665_bfr_after (
		.din(new_net_18664),
		.dout(new_net_18665)
	);

	bfr new_net_18666_bfr_after (
		.din(new_net_18665),
		.dout(new_net_18666)
	);

	bfr new_net_18667_bfr_after (
		.din(new_net_18666),
		.dout(new_net_18667)
	);

	bfr new_net_18668_bfr_after (
		.din(new_net_18667),
		.dout(new_net_18668)
	);

	bfr new_net_18669_bfr_after (
		.din(new_net_18668),
		.dout(new_net_18669)
	);

	bfr new_net_18670_bfr_after (
		.din(new_net_18669),
		.dout(new_net_18670)
	);

	bfr new_net_18671_bfr_after (
		.din(new_net_18670),
		.dout(new_net_18671)
	);

	bfr new_net_18672_bfr_after (
		.din(new_net_18671),
		.dout(new_net_18672)
	);

	bfr new_net_18673_bfr_after (
		.din(new_net_18672),
		.dout(new_net_18673)
	);

	bfr new_net_18674_bfr_after (
		.din(new_net_18673),
		.dout(new_net_18674)
	);

	bfr new_net_18675_bfr_after (
		.din(new_net_18674),
		.dout(new_net_18675)
	);

	bfr new_net_18676_bfr_after (
		.din(new_net_18675),
		.dout(new_net_18676)
	);

	bfr new_net_18677_bfr_after (
		.din(new_net_18676),
		.dout(new_net_18677)
	);

	bfr new_net_18678_bfr_after (
		.din(new_net_18677),
		.dout(new_net_18678)
	);

	bfr new_net_18679_bfr_after (
		.din(new_net_18678),
		.dout(new_net_18679)
	);

	bfr new_net_18680_bfr_after (
		.din(new_net_18679),
		.dout(new_net_18680)
	);

	bfr new_net_18681_bfr_after (
		.din(new_net_18680),
		.dout(new_net_18681)
	);

	bfr new_net_18682_bfr_after (
		.din(new_net_18681),
		.dout(new_net_18682)
	);

	bfr new_net_18683_bfr_after (
		.din(new_net_18682),
		.dout(new_net_18683)
	);

	bfr new_net_18684_bfr_after (
		.din(new_net_18683),
		.dout(new_net_18684)
	);

	bfr new_net_18685_bfr_after (
		.din(new_net_18684),
		.dout(new_net_18685)
	);

	bfr new_net_18686_bfr_after (
		.din(new_net_18685),
		.dout(new_net_18686)
	);

	bfr new_net_18687_bfr_after (
		.din(new_net_18686),
		.dout(new_net_18687)
	);

	bfr new_net_18688_bfr_after (
		.din(new_net_18687),
		.dout(new_net_18688)
	);

	bfr new_net_18689_bfr_after (
		.din(new_net_18688),
		.dout(new_net_18689)
	);

	bfr new_net_18690_bfr_after (
		.din(new_net_18689),
		.dout(new_net_18690)
	);

	bfr new_net_18691_bfr_after (
		.din(new_net_18690),
		.dout(new_net_18691)
	);

	bfr new_net_18692_bfr_after (
		.din(new_net_18691),
		.dout(new_net_18692)
	);

	bfr new_net_18693_bfr_after (
		.din(new_net_18692),
		.dout(new_net_18693)
	);

	bfr new_net_18694_bfr_after (
		.din(new_net_18693),
		.dout(new_net_18694)
	);

	bfr new_net_18695_bfr_after (
		.din(new_net_18694),
		.dout(new_net_18695)
	);

	bfr new_net_18696_bfr_after (
		.din(new_net_18695),
		.dout(new_net_18696)
	);

	bfr new_net_18697_bfr_after (
		.din(new_net_18696),
		.dout(new_net_18697)
	);

	bfr new_net_18698_bfr_after (
		.din(new_net_18697),
		.dout(new_net_18698)
	);

	bfr new_net_18699_bfr_after (
		.din(new_net_18698),
		.dout(new_net_18699)
	);

	bfr new_net_18700_bfr_after (
		.din(new_net_18699),
		.dout(new_net_18700)
	);

	bfr new_net_18701_bfr_after (
		.din(new_net_18700),
		.dout(new_net_18701)
	);

	bfr new_net_18702_bfr_after (
		.din(new_net_18701),
		.dout(new_net_18702)
	);

	bfr new_net_18703_bfr_after (
		.din(new_net_18702),
		.dout(new_net_18703)
	);

	bfr new_net_18704_bfr_after (
		.din(new_net_18703),
		.dout(new_net_18704)
	);

	bfr new_net_18705_bfr_after (
		.din(new_net_18704),
		.dout(new_net_18705)
	);

	bfr new_net_18706_bfr_after (
		.din(new_net_18705),
		.dout(new_net_18706)
	);

	bfr new_net_18707_bfr_after (
		.din(new_net_18706),
		.dout(new_net_18707)
	);

	bfr new_net_18708_bfr_after (
		.din(new_net_18707),
		.dout(new_net_18708)
	);

	spl2 _1569__v_fanout (
		.a(new_net_18708),
		.b(new_net_1648),
		.c(new_net_1649)
	);

	bfr new_net_18709_bfr_after (
		.din(_1461_),
		.dout(new_net_18709)
	);

	bfr new_net_18710_bfr_after (
		.din(new_net_18709),
		.dout(new_net_18710)
	);

	bfr new_net_18711_bfr_after (
		.din(new_net_18710),
		.dout(new_net_18711)
	);

	bfr new_net_18712_bfr_after (
		.din(new_net_18711),
		.dout(new_net_18712)
	);

	bfr new_net_18713_bfr_after (
		.din(new_net_18712),
		.dout(new_net_18713)
	);

	bfr new_net_18714_bfr_after (
		.din(new_net_18713),
		.dout(new_net_18714)
	);

	bfr new_net_18715_bfr_after (
		.din(new_net_18714),
		.dout(new_net_18715)
	);

	bfr new_net_18716_bfr_after (
		.din(new_net_18715),
		.dout(new_net_18716)
	);

	bfr new_net_18717_bfr_after (
		.din(new_net_18716),
		.dout(new_net_18717)
	);

	bfr new_net_18718_bfr_after (
		.din(new_net_18717),
		.dout(new_net_18718)
	);

	bfr new_net_18719_bfr_after (
		.din(new_net_18718),
		.dout(new_net_18719)
	);

	bfr new_net_18720_bfr_after (
		.din(new_net_18719),
		.dout(new_net_18720)
	);

	bfr new_net_18721_bfr_after (
		.din(new_net_18720),
		.dout(new_net_18721)
	);

	bfr new_net_18722_bfr_after (
		.din(new_net_18721),
		.dout(new_net_18722)
	);

	bfr new_net_18723_bfr_after (
		.din(new_net_18722),
		.dout(new_net_18723)
	);

	bfr new_net_18724_bfr_after (
		.din(new_net_18723),
		.dout(new_net_18724)
	);

	bfr new_net_18725_bfr_after (
		.din(new_net_18724),
		.dout(new_net_18725)
	);

	bfr new_net_18726_bfr_after (
		.din(new_net_18725),
		.dout(new_net_18726)
	);

	bfr new_net_18727_bfr_after (
		.din(new_net_18726),
		.dout(new_net_18727)
	);

	bfr new_net_18728_bfr_after (
		.din(new_net_18727),
		.dout(new_net_18728)
	);

	bfr new_net_18729_bfr_after (
		.din(new_net_18728),
		.dout(new_net_18729)
	);

	bfr new_net_18730_bfr_after (
		.din(new_net_18729),
		.dout(new_net_18730)
	);

	bfr new_net_18731_bfr_after (
		.din(new_net_18730),
		.dout(new_net_18731)
	);

	bfr new_net_18732_bfr_after (
		.din(new_net_18731),
		.dout(new_net_18732)
	);

	bfr new_net_18733_bfr_after (
		.din(new_net_18732),
		.dout(new_net_18733)
	);

	bfr new_net_18734_bfr_after (
		.din(new_net_18733),
		.dout(new_net_18734)
	);

	bfr new_net_18735_bfr_after (
		.din(new_net_18734),
		.dout(new_net_18735)
	);

	bfr new_net_18736_bfr_after (
		.din(new_net_18735),
		.dout(new_net_18736)
	);

	bfr new_net_18737_bfr_after (
		.din(new_net_18736),
		.dout(new_net_18737)
	);

	bfr new_net_18738_bfr_after (
		.din(new_net_18737),
		.dout(new_net_18738)
	);

	bfr new_net_18739_bfr_after (
		.din(new_net_18738),
		.dout(new_net_18739)
	);

	bfr new_net_18740_bfr_after (
		.din(new_net_18739),
		.dout(new_net_18740)
	);

	bfr new_net_18741_bfr_after (
		.din(new_net_18740),
		.dout(new_net_18741)
	);

	bfr new_net_18742_bfr_after (
		.din(new_net_18741),
		.dout(new_net_18742)
	);

	bfr new_net_18743_bfr_after (
		.din(new_net_18742),
		.dout(new_net_18743)
	);

	bfr new_net_18744_bfr_after (
		.din(new_net_18743),
		.dout(new_net_18744)
	);

	bfr new_net_18745_bfr_after (
		.din(new_net_18744),
		.dout(new_net_18745)
	);

	bfr new_net_18746_bfr_after (
		.din(new_net_18745),
		.dout(new_net_18746)
	);

	bfr new_net_18747_bfr_after (
		.din(new_net_18746),
		.dout(new_net_18747)
	);

	bfr new_net_18748_bfr_after (
		.din(new_net_18747),
		.dout(new_net_18748)
	);

	bfr new_net_18749_bfr_after (
		.din(new_net_18748),
		.dout(new_net_18749)
	);

	bfr new_net_18750_bfr_after (
		.din(new_net_18749),
		.dout(new_net_18750)
	);

	bfr new_net_18751_bfr_after (
		.din(new_net_18750),
		.dout(new_net_18751)
	);

	bfr new_net_18752_bfr_after (
		.din(new_net_18751),
		.dout(new_net_18752)
	);

	bfr new_net_18753_bfr_after (
		.din(new_net_18752),
		.dout(new_net_18753)
	);

	bfr new_net_18754_bfr_after (
		.din(new_net_18753),
		.dout(new_net_18754)
	);

	bfr new_net_18755_bfr_after (
		.din(new_net_18754),
		.dout(new_net_18755)
	);

	bfr new_net_18756_bfr_after (
		.din(new_net_18755),
		.dout(new_net_18756)
	);

	bfr new_net_18757_bfr_after (
		.din(new_net_18756),
		.dout(new_net_18757)
	);

	bfr new_net_18758_bfr_after (
		.din(new_net_18757),
		.dout(new_net_18758)
	);

	bfr new_net_18759_bfr_after (
		.din(new_net_18758),
		.dout(new_net_18759)
	);

	bfr new_net_18760_bfr_after (
		.din(new_net_18759),
		.dout(new_net_18760)
	);

	bfr new_net_18761_bfr_after (
		.din(new_net_18760),
		.dout(new_net_18761)
	);

	bfr new_net_18762_bfr_after (
		.din(new_net_18761),
		.dout(new_net_18762)
	);

	bfr new_net_18763_bfr_after (
		.din(new_net_18762),
		.dout(new_net_18763)
	);

	bfr new_net_18764_bfr_after (
		.din(new_net_18763),
		.dout(new_net_18764)
	);

	bfr new_net_18765_bfr_after (
		.din(new_net_18764),
		.dout(new_net_18765)
	);

	bfr new_net_18766_bfr_after (
		.din(new_net_18765),
		.dout(new_net_18766)
	);

	bfr new_net_18767_bfr_after (
		.din(new_net_18766),
		.dout(new_net_18767)
	);

	bfr new_net_18768_bfr_after (
		.din(new_net_18767),
		.dout(new_net_18768)
	);

	bfr new_net_18769_bfr_after (
		.din(new_net_18768),
		.dout(new_net_18769)
	);

	bfr new_net_18770_bfr_after (
		.din(new_net_18769),
		.dout(new_net_18770)
	);

	bfr new_net_18771_bfr_after (
		.din(new_net_18770),
		.dout(new_net_18771)
	);

	bfr new_net_18772_bfr_after (
		.din(new_net_18771),
		.dout(new_net_18772)
	);

	bfr new_net_18773_bfr_after (
		.din(new_net_18772),
		.dout(new_net_18773)
	);

	spl2 _1461__v_fanout (
		.a(new_net_18773),
		.b(new_net_769),
		.c(new_net_770)
	);

	bfr new_net_18774_bfr_after (
		.din(_0066_),
		.dout(new_net_18774)
	);

	spl2 _0066__v_fanout (
		.a(new_net_18774),
		.b(new_net_1632),
		.c(new_net_1633)
	);

	bfr new_net_18775_bfr_after (
		.din(_0044_),
		.dout(new_net_18775)
	);

	spl2 _0044__v_fanout (
		.a(new_net_18775),
		.b(new_net_888),
		.c(new_net_889)
	);

	bfr new_net_18776_bfr_after (
		.din(_1809_),
		.dout(new_net_18776)
	);

	bfr new_net_18777_bfr_after (
		.din(new_net_18776),
		.dout(new_net_18777)
	);

	bfr new_net_18778_bfr_after (
		.din(new_net_18777),
		.dout(new_net_18778)
	);

	bfr new_net_18779_bfr_after (
		.din(new_net_18778),
		.dout(new_net_18779)
	);

	bfr new_net_18780_bfr_after (
		.din(new_net_18779),
		.dout(new_net_18780)
	);

	bfr new_net_18781_bfr_after (
		.din(new_net_18780),
		.dout(new_net_18781)
	);

	bfr new_net_18782_bfr_after (
		.din(new_net_18781),
		.dout(new_net_18782)
	);

	bfr new_net_18783_bfr_after (
		.din(new_net_18782),
		.dout(new_net_18783)
	);

	bfr new_net_18784_bfr_after (
		.din(new_net_18783),
		.dout(new_net_18784)
	);

	bfr new_net_18785_bfr_after (
		.din(new_net_18784),
		.dout(new_net_18785)
	);

	bfr new_net_18786_bfr_after (
		.din(new_net_18785),
		.dout(new_net_18786)
	);

	bfr new_net_18787_bfr_after (
		.din(new_net_18786),
		.dout(new_net_18787)
	);

	bfr new_net_18788_bfr_after (
		.din(new_net_18787),
		.dout(new_net_18788)
	);

	bfr new_net_18789_bfr_after (
		.din(new_net_18788),
		.dout(new_net_18789)
	);

	bfr new_net_18790_bfr_after (
		.din(new_net_18789),
		.dout(new_net_18790)
	);

	bfr new_net_18791_bfr_after (
		.din(new_net_18790),
		.dout(new_net_18791)
	);

	bfr new_net_18792_bfr_after (
		.din(new_net_18791),
		.dout(new_net_18792)
	);

	bfr new_net_18793_bfr_after (
		.din(new_net_18792),
		.dout(new_net_18793)
	);

	bfr new_net_18794_bfr_after (
		.din(new_net_18793),
		.dout(new_net_18794)
	);

	bfr new_net_18795_bfr_after (
		.din(new_net_18794),
		.dout(new_net_18795)
	);

	bfr new_net_18796_bfr_after (
		.din(new_net_18795),
		.dout(new_net_18796)
	);

	bfr new_net_18797_bfr_after (
		.din(new_net_18796),
		.dout(new_net_18797)
	);

	bfr new_net_18798_bfr_after (
		.din(new_net_18797),
		.dout(new_net_18798)
	);

	bfr new_net_18799_bfr_after (
		.din(new_net_18798),
		.dout(new_net_18799)
	);

	bfr new_net_18800_bfr_after (
		.din(new_net_18799),
		.dout(new_net_18800)
	);

	bfr new_net_18801_bfr_after (
		.din(new_net_18800),
		.dout(new_net_18801)
	);

	bfr new_net_18802_bfr_after (
		.din(new_net_18801),
		.dout(new_net_18802)
	);

	bfr new_net_18803_bfr_after (
		.din(new_net_18802),
		.dout(new_net_18803)
	);

	bfr new_net_18804_bfr_after (
		.din(new_net_18803),
		.dout(new_net_18804)
	);

	bfr new_net_18805_bfr_after (
		.din(new_net_18804),
		.dout(new_net_18805)
	);

	bfr new_net_18806_bfr_after (
		.din(new_net_18805),
		.dout(new_net_18806)
	);

	bfr new_net_18807_bfr_after (
		.din(new_net_18806),
		.dout(new_net_18807)
	);

	bfr new_net_18808_bfr_after (
		.din(new_net_18807),
		.dout(new_net_18808)
	);

	bfr new_net_18809_bfr_after (
		.din(new_net_18808),
		.dout(new_net_18809)
	);

	bfr new_net_18810_bfr_after (
		.din(new_net_18809),
		.dout(new_net_18810)
	);

	bfr new_net_18811_bfr_after (
		.din(new_net_18810),
		.dout(new_net_18811)
	);

	bfr new_net_18812_bfr_after (
		.din(new_net_18811),
		.dout(new_net_18812)
	);

	bfr new_net_18813_bfr_after (
		.din(new_net_18812),
		.dout(new_net_18813)
	);

	bfr new_net_18814_bfr_after (
		.din(new_net_18813),
		.dout(new_net_18814)
	);

	bfr new_net_18815_bfr_after (
		.din(new_net_18814),
		.dout(new_net_18815)
	);

	bfr new_net_18816_bfr_after (
		.din(new_net_18815),
		.dout(new_net_18816)
	);

	bfr new_net_18817_bfr_after (
		.din(new_net_18816),
		.dout(new_net_18817)
	);

	bfr new_net_18818_bfr_after (
		.din(new_net_18817),
		.dout(new_net_18818)
	);

	bfr new_net_18819_bfr_after (
		.din(new_net_18818),
		.dout(new_net_18819)
	);

	bfr new_net_18820_bfr_after (
		.din(new_net_18819),
		.dout(new_net_18820)
	);

	bfr new_net_18821_bfr_after (
		.din(new_net_18820),
		.dout(new_net_18821)
	);

	bfr new_net_18822_bfr_after (
		.din(new_net_18821),
		.dout(new_net_18822)
	);

	bfr new_net_18823_bfr_after (
		.din(new_net_18822),
		.dout(new_net_18823)
	);

	bfr new_net_18824_bfr_after (
		.din(new_net_18823),
		.dout(new_net_18824)
	);

	bfr new_net_18825_bfr_after (
		.din(new_net_18824),
		.dout(new_net_18825)
	);

	bfr new_net_18826_bfr_after (
		.din(new_net_18825),
		.dout(new_net_18826)
	);

	bfr new_net_18827_bfr_after (
		.din(new_net_18826),
		.dout(new_net_18827)
	);

	bfr new_net_18828_bfr_after (
		.din(new_net_18827),
		.dout(new_net_18828)
	);

	bfr new_net_18829_bfr_after (
		.din(new_net_18828),
		.dout(new_net_18829)
	);

	bfr new_net_18830_bfr_after (
		.din(new_net_18829),
		.dout(new_net_18830)
	);

	bfr new_net_18831_bfr_after (
		.din(new_net_18830),
		.dout(new_net_18831)
	);

	bfr new_net_18832_bfr_after (
		.din(new_net_18831),
		.dout(new_net_18832)
	);

	bfr new_net_18833_bfr_after (
		.din(new_net_18832),
		.dout(new_net_18833)
	);

	bfr new_net_18834_bfr_after (
		.din(new_net_18833),
		.dout(new_net_18834)
	);

	bfr new_net_18835_bfr_after (
		.din(new_net_18834),
		.dout(new_net_18835)
	);

	bfr new_net_18836_bfr_after (
		.din(new_net_18835),
		.dout(new_net_18836)
	);

	bfr new_net_18837_bfr_after (
		.din(new_net_18836),
		.dout(new_net_18837)
	);

	bfr new_net_18838_bfr_after (
		.din(new_net_18837),
		.dout(new_net_18838)
	);

	bfr new_net_18839_bfr_after (
		.din(new_net_18838),
		.dout(new_net_18839)
	);

	bfr new_net_18840_bfr_after (
		.din(new_net_18839),
		.dout(new_net_18840)
	);

	bfr new_net_18841_bfr_after (
		.din(new_net_18840),
		.dout(new_net_18841)
	);

	bfr new_net_18842_bfr_after (
		.din(new_net_18841),
		.dout(new_net_18842)
	);

	bfr new_net_18843_bfr_after (
		.din(new_net_18842),
		.dout(new_net_18843)
	);

	bfr new_net_18844_bfr_after (
		.din(new_net_18843),
		.dout(new_net_18844)
	);

	bfr new_net_18845_bfr_after (
		.din(new_net_18844),
		.dout(new_net_18845)
	);

	bfr new_net_18846_bfr_after (
		.din(new_net_18845),
		.dout(new_net_18846)
	);

	bfr new_net_18847_bfr_after (
		.din(new_net_18846),
		.dout(new_net_18847)
	);

	bfr new_net_18848_bfr_after (
		.din(new_net_18847),
		.dout(new_net_18848)
	);

	bfr new_net_18849_bfr_after (
		.din(new_net_18848),
		.dout(new_net_18849)
	);

	bfr new_net_18850_bfr_after (
		.din(new_net_18849),
		.dout(new_net_18850)
	);

	bfr new_net_18851_bfr_after (
		.din(new_net_18850),
		.dout(new_net_18851)
	);

	bfr new_net_18852_bfr_after (
		.din(new_net_18851),
		.dout(new_net_18852)
	);

	bfr new_net_18853_bfr_after (
		.din(new_net_18852),
		.dout(new_net_18853)
	);

	bfr new_net_18854_bfr_after (
		.din(new_net_18853),
		.dout(new_net_18854)
	);

	bfr new_net_18855_bfr_after (
		.din(new_net_18854),
		.dout(new_net_18855)
	);

	bfr new_net_18856_bfr_after (
		.din(new_net_18855),
		.dout(new_net_18856)
	);

	bfr new_net_18857_bfr_after (
		.din(new_net_18856),
		.dout(new_net_18857)
	);

	bfr new_net_18858_bfr_after (
		.din(new_net_18857),
		.dout(new_net_18858)
	);

	bfr new_net_18859_bfr_after (
		.din(new_net_18858),
		.dout(new_net_18859)
	);

	bfr new_net_18860_bfr_after (
		.din(new_net_18859),
		.dout(new_net_18860)
	);

	bfr new_net_18861_bfr_after (
		.din(new_net_18860),
		.dout(new_net_18861)
	);

	bfr new_net_18862_bfr_after (
		.din(new_net_18861),
		.dout(new_net_18862)
	);

	bfr new_net_18863_bfr_after (
		.din(new_net_18862),
		.dout(new_net_18863)
	);

	bfr new_net_18864_bfr_after (
		.din(new_net_18863),
		.dout(new_net_18864)
	);

	spl2 _1809__v_fanout (
		.a(new_net_18864),
		.b(new_net_1154),
		.c(new_net_1155)
	);

	bfr new_net_18865_bfr_after (
		.din(_1028_),
		.dout(new_net_18865)
	);

	bfr new_net_18866_bfr_after (
		.din(new_net_18865),
		.dout(new_net_18866)
	);

	bfr new_net_18867_bfr_after (
		.din(new_net_18866),
		.dout(new_net_18867)
	);

	bfr new_net_18868_bfr_after (
		.din(new_net_18867),
		.dout(new_net_18868)
	);

	bfr new_net_18869_bfr_after (
		.din(new_net_18868),
		.dout(new_net_18869)
	);

	bfr new_net_18870_bfr_after (
		.din(new_net_18869),
		.dout(new_net_18870)
	);

	bfr new_net_18871_bfr_after (
		.din(new_net_18870),
		.dout(new_net_18871)
	);

	bfr new_net_18872_bfr_after (
		.din(new_net_18871),
		.dout(new_net_18872)
	);

	bfr new_net_18873_bfr_after (
		.din(new_net_18872),
		.dout(new_net_18873)
	);

	bfr new_net_18874_bfr_after (
		.din(new_net_18873),
		.dout(new_net_18874)
	);

	bfr new_net_18875_bfr_after (
		.din(new_net_18874),
		.dout(new_net_18875)
	);

	bfr new_net_18876_bfr_after (
		.din(new_net_18875),
		.dout(new_net_18876)
	);

	bfr new_net_18877_bfr_after (
		.din(new_net_18876),
		.dout(new_net_18877)
	);

	bfr new_net_18878_bfr_after (
		.din(new_net_18877),
		.dout(new_net_18878)
	);

	bfr new_net_18879_bfr_after (
		.din(new_net_18878),
		.dout(new_net_18879)
	);

	bfr new_net_18880_bfr_after (
		.din(new_net_18879),
		.dout(new_net_18880)
	);

	bfr new_net_18881_bfr_after (
		.din(new_net_18880),
		.dout(new_net_18881)
	);

	spl2 _1028__v_fanout (
		.a(new_net_18881),
		.b(new_net_2096),
		.c(new_net_2097)
	);

	bfr new_net_18882_bfr_after (
		.din(_0326_),
		.dout(new_net_18882)
	);

	bfr new_net_18883_bfr_after (
		.din(new_net_18882),
		.dout(new_net_18883)
	);

	bfr new_net_18884_bfr_after (
		.din(new_net_18883),
		.dout(new_net_18884)
	);

	bfr new_net_18885_bfr_after (
		.din(new_net_18884),
		.dout(new_net_18885)
	);

	bfr new_net_18886_bfr_after (
		.din(new_net_18885),
		.dout(new_net_18886)
	);

	bfr new_net_18887_bfr_after (
		.din(new_net_18886),
		.dout(new_net_18887)
	);

	bfr new_net_18888_bfr_after (
		.din(new_net_18887),
		.dout(new_net_18888)
	);

	bfr new_net_18889_bfr_after (
		.din(new_net_18888),
		.dout(new_net_18889)
	);

	bfr new_net_18890_bfr_after (
		.din(new_net_18889),
		.dout(new_net_18890)
	);

	bfr new_net_18891_bfr_after (
		.din(new_net_18890),
		.dout(new_net_18891)
	);

	bfr new_net_18892_bfr_after (
		.din(new_net_18891),
		.dout(new_net_18892)
	);

	bfr new_net_18893_bfr_after (
		.din(new_net_18892),
		.dout(new_net_18893)
	);

	bfr new_net_18894_bfr_after (
		.din(new_net_18893),
		.dout(new_net_18894)
	);

	bfr new_net_18895_bfr_after (
		.din(new_net_18894),
		.dout(new_net_18895)
	);

	bfr new_net_18896_bfr_after (
		.din(new_net_18895),
		.dout(new_net_18896)
	);

	bfr new_net_18897_bfr_after (
		.din(new_net_18896),
		.dout(new_net_18897)
	);

	bfr new_net_18898_bfr_after (
		.din(new_net_18897),
		.dout(new_net_18898)
	);

	bfr new_net_18899_bfr_after (
		.din(new_net_18898),
		.dout(new_net_18899)
	);

	bfr new_net_18900_bfr_after (
		.din(new_net_18899),
		.dout(new_net_18900)
	);

	bfr new_net_18901_bfr_after (
		.din(new_net_18900),
		.dout(new_net_18901)
	);

	bfr new_net_18902_bfr_after (
		.din(new_net_18901),
		.dout(new_net_18902)
	);

	bfr new_net_18903_bfr_after (
		.din(new_net_18902),
		.dout(new_net_18903)
	);

	bfr new_net_18904_bfr_after (
		.din(new_net_18903),
		.dout(new_net_18904)
	);

	bfr new_net_18905_bfr_after (
		.din(new_net_18904),
		.dout(new_net_18905)
	);

	bfr new_net_18906_bfr_after (
		.din(new_net_18905),
		.dout(new_net_18906)
	);

	bfr new_net_18907_bfr_after (
		.din(new_net_18906),
		.dout(new_net_18907)
	);

	bfr new_net_18908_bfr_after (
		.din(new_net_18907),
		.dout(new_net_18908)
	);

	bfr new_net_18909_bfr_after (
		.din(new_net_18908),
		.dout(new_net_18909)
	);

	bfr new_net_18910_bfr_after (
		.din(new_net_18909),
		.dout(new_net_18910)
	);

	bfr new_net_18911_bfr_after (
		.din(new_net_18910),
		.dout(new_net_18911)
	);

	bfr new_net_18912_bfr_after (
		.din(new_net_18911),
		.dout(new_net_18912)
	);

	bfr new_net_18913_bfr_after (
		.din(new_net_18912),
		.dout(new_net_18913)
	);

	bfr new_net_18914_bfr_after (
		.din(new_net_18913),
		.dout(new_net_18914)
	);

	bfr new_net_18915_bfr_after (
		.din(new_net_18914),
		.dout(new_net_18915)
	);

	bfr new_net_18916_bfr_after (
		.din(new_net_18915),
		.dout(new_net_18916)
	);

	bfr new_net_18917_bfr_after (
		.din(new_net_18916),
		.dout(new_net_18917)
	);

	bfr new_net_18918_bfr_after (
		.din(new_net_18917),
		.dout(new_net_18918)
	);

	bfr new_net_18919_bfr_after (
		.din(new_net_18918),
		.dout(new_net_18919)
	);

	bfr new_net_18920_bfr_after (
		.din(new_net_18919),
		.dout(new_net_18920)
	);

	bfr new_net_18921_bfr_after (
		.din(new_net_18920),
		.dout(new_net_18921)
	);

	bfr new_net_18922_bfr_after (
		.din(new_net_18921),
		.dout(new_net_18922)
	);

	bfr new_net_18923_bfr_after (
		.din(new_net_18922),
		.dout(new_net_18923)
	);

	bfr new_net_18924_bfr_after (
		.din(new_net_18923),
		.dout(new_net_18924)
	);

	bfr new_net_18925_bfr_after (
		.din(new_net_18924),
		.dout(new_net_18925)
	);

	bfr new_net_18926_bfr_after (
		.din(new_net_18925),
		.dout(new_net_18926)
	);

	bfr new_net_18927_bfr_after (
		.din(new_net_18926),
		.dout(new_net_18927)
	);

	bfr new_net_18928_bfr_after (
		.din(new_net_18927),
		.dout(new_net_18928)
	);

	bfr new_net_18929_bfr_after (
		.din(new_net_18928),
		.dout(new_net_18929)
	);

	bfr new_net_18930_bfr_after (
		.din(new_net_18929),
		.dout(new_net_18930)
	);

	bfr new_net_18931_bfr_after (
		.din(new_net_18930),
		.dout(new_net_18931)
	);

	bfr new_net_18932_bfr_after (
		.din(new_net_18931),
		.dout(new_net_18932)
	);

	bfr new_net_18933_bfr_after (
		.din(new_net_18932),
		.dout(new_net_18933)
	);

	bfr new_net_18934_bfr_after (
		.din(new_net_18933),
		.dout(new_net_18934)
	);

	bfr new_net_18935_bfr_after (
		.din(new_net_18934),
		.dout(new_net_18935)
	);

	bfr new_net_18936_bfr_after (
		.din(new_net_18935),
		.dout(new_net_18936)
	);

	bfr new_net_18937_bfr_after (
		.din(new_net_18936),
		.dout(new_net_18937)
	);

	bfr new_net_18938_bfr_after (
		.din(new_net_18937),
		.dout(new_net_18938)
	);

	bfr new_net_18939_bfr_after (
		.din(new_net_18938),
		.dout(new_net_18939)
	);

	bfr new_net_18940_bfr_after (
		.din(new_net_18939),
		.dout(new_net_18940)
	);

	bfr new_net_18941_bfr_after (
		.din(new_net_18940),
		.dout(new_net_18941)
	);

	bfr new_net_18942_bfr_after (
		.din(new_net_18941),
		.dout(new_net_18942)
	);

	bfr new_net_18943_bfr_after (
		.din(new_net_18942),
		.dout(new_net_18943)
	);

	bfr new_net_18944_bfr_after (
		.din(new_net_18943),
		.dout(new_net_18944)
	);

	bfr new_net_18945_bfr_after (
		.din(new_net_18944),
		.dout(new_net_18945)
	);

	bfr new_net_18946_bfr_after (
		.din(new_net_18945),
		.dout(new_net_18946)
	);

	bfr new_net_18947_bfr_after (
		.din(new_net_18946),
		.dout(new_net_18947)
	);

	bfr new_net_18948_bfr_after (
		.din(new_net_18947),
		.dout(new_net_18948)
	);

	bfr new_net_18949_bfr_after (
		.din(new_net_18948),
		.dout(new_net_18949)
	);

	bfr new_net_18950_bfr_after (
		.din(new_net_18949),
		.dout(new_net_18950)
	);

	bfr new_net_18951_bfr_after (
		.din(new_net_18950),
		.dout(new_net_18951)
	);

	bfr new_net_18952_bfr_after (
		.din(new_net_18951),
		.dout(new_net_18952)
	);

	bfr new_net_18953_bfr_after (
		.din(new_net_18952),
		.dout(new_net_18953)
	);

	bfr new_net_18954_bfr_after (
		.din(new_net_18953),
		.dout(new_net_18954)
	);

	bfr new_net_18955_bfr_after (
		.din(new_net_18954),
		.dout(new_net_18955)
	);

	bfr new_net_18956_bfr_after (
		.din(new_net_18955),
		.dout(new_net_18956)
	);

	bfr new_net_18957_bfr_after (
		.din(new_net_18956),
		.dout(new_net_18957)
	);

	bfr new_net_18958_bfr_after (
		.din(new_net_18957),
		.dout(new_net_18958)
	);

	bfr new_net_18959_bfr_after (
		.din(new_net_18958),
		.dout(new_net_18959)
	);

	bfr new_net_18960_bfr_after (
		.din(new_net_18959),
		.dout(new_net_18960)
	);

	bfr new_net_18961_bfr_after (
		.din(new_net_18960),
		.dout(new_net_18961)
	);

	bfr new_net_18962_bfr_after (
		.din(new_net_18961),
		.dout(new_net_18962)
	);

	bfr new_net_18963_bfr_after (
		.din(new_net_18962),
		.dout(new_net_18963)
	);

	bfr new_net_18964_bfr_after (
		.din(new_net_18963),
		.dout(new_net_18964)
	);

	bfr new_net_18965_bfr_after (
		.din(new_net_18964),
		.dout(new_net_18965)
	);

	bfr new_net_18966_bfr_after (
		.din(new_net_18965),
		.dout(new_net_18966)
	);

	bfr new_net_18967_bfr_after (
		.din(new_net_18966),
		.dout(new_net_18967)
	);

	bfr new_net_18968_bfr_after (
		.din(new_net_18967),
		.dout(new_net_18968)
	);

	bfr new_net_18969_bfr_after (
		.din(new_net_18968),
		.dout(new_net_18969)
	);

	bfr new_net_18970_bfr_after (
		.din(new_net_18969),
		.dout(new_net_18970)
	);

	bfr new_net_18971_bfr_after (
		.din(new_net_18970),
		.dout(new_net_18971)
	);

	bfr new_net_18972_bfr_after (
		.din(new_net_18971),
		.dout(new_net_18972)
	);

	bfr new_net_18973_bfr_after (
		.din(new_net_18972),
		.dout(new_net_18973)
	);

	bfr new_net_18974_bfr_after (
		.din(new_net_18973),
		.dout(new_net_18974)
	);

	bfr new_net_18975_bfr_after (
		.din(new_net_18974),
		.dout(new_net_18975)
	);

	bfr new_net_18976_bfr_after (
		.din(new_net_18975),
		.dout(new_net_18976)
	);

	bfr new_net_18977_bfr_after (
		.din(new_net_18976),
		.dout(new_net_18977)
	);

	bfr new_net_18978_bfr_after (
		.din(new_net_18977),
		.dout(new_net_18978)
	);

	bfr new_net_18979_bfr_after (
		.din(new_net_18978),
		.dout(new_net_18979)
	);

	bfr new_net_18980_bfr_after (
		.din(new_net_18979),
		.dout(new_net_18980)
	);

	bfr new_net_18981_bfr_after (
		.din(new_net_18980),
		.dout(new_net_18981)
	);

	bfr new_net_18982_bfr_after (
		.din(new_net_18981),
		.dout(new_net_18982)
	);

	bfr new_net_18983_bfr_after (
		.din(new_net_18982),
		.dout(new_net_18983)
	);

	bfr new_net_18984_bfr_after (
		.din(new_net_18983),
		.dout(new_net_18984)
	);

	bfr new_net_18985_bfr_after (
		.din(new_net_18984),
		.dout(new_net_18985)
	);

	bfr new_net_18986_bfr_after (
		.din(new_net_18985),
		.dout(new_net_18986)
	);

	bfr new_net_18987_bfr_after (
		.din(new_net_18986),
		.dout(new_net_18987)
	);

	bfr new_net_18988_bfr_after (
		.din(new_net_18987),
		.dout(new_net_18988)
	);

	bfr new_net_18989_bfr_after (
		.din(new_net_18988),
		.dout(new_net_18989)
	);

	bfr new_net_18990_bfr_after (
		.din(new_net_18989),
		.dout(new_net_18990)
	);

	bfr new_net_18991_bfr_after (
		.din(new_net_18990),
		.dout(new_net_18991)
	);

	bfr new_net_18992_bfr_after (
		.din(new_net_18991),
		.dout(new_net_18992)
	);

	bfr new_net_18993_bfr_after (
		.din(new_net_18992),
		.dout(new_net_18993)
	);

	bfr new_net_18994_bfr_after (
		.din(new_net_18993),
		.dout(new_net_18994)
	);

	spl2 _0326__v_fanout (
		.a(new_net_18994),
		.b(new_net_711),
		.c(new_net_712)
	);

	bfr new_net_18995_bfr_after (
		.din(_1369_),
		.dout(new_net_18995)
	);

	bfr new_net_18996_bfr_after (
		.din(new_net_18995),
		.dout(new_net_18996)
	);

	bfr new_net_18997_bfr_after (
		.din(new_net_18996),
		.dout(new_net_18997)
	);

	bfr new_net_18998_bfr_after (
		.din(new_net_18997),
		.dout(new_net_18998)
	);

	bfr new_net_18999_bfr_after (
		.din(new_net_18998),
		.dout(new_net_18999)
	);

	bfr new_net_19000_bfr_after (
		.din(new_net_18999),
		.dout(new_net_19000)
	);

	bfr new_net_19001_bfr_after (
		.din(new_net_19000),
		.dout(new_net_19001)
	);

	bfr new_net_19002_bfr_after (
		.din(new_net_19001),
		.dout(new_net_19002)
	);

	bfr new_net_19003_bfr_after (
		.din(new_net_19002),
		.dout(new_net_19003)
	);

	bfr new_net_19004_bfr_after (
		.din(new_net_19003),
		.dout(new_net_19004)
	);

	bfr new_net_19005_bfr_after (
		.din(new_net_19004),
		.dout(new_net_19005)
	);

	bfr new_net_19006_bfr_after (
		.din(new_net_19005),
		.dout(new_net_19006)
	);

	bfr new_net_19007_bfr_after (
		.din(new_net_19006),
		.dout(new_net_19007)
	);

	bfr new_net_19008_bfr_after (
		.din(new_net_19007),
		.dout(new_net_19008)
	);

	bfr new_net_19009_bfr_after (
		.din(new_net_19008),
		.dout(new_net_19009)
	);

	bfr new_net_19010_bfr_after (
		.din(new_net_19009),
		.dout(new_net_19010)
	);

	bfr new_net_19011_bfr_after (
		.din(new_net_19010),
		.dout(new_net_19011)
	);

	bfr new_net_19012_bfr_after (
		.din(new_net_19011),
		.dout(new_net_19012)
	);

	bfr new_net_19013_bfr_after (
		.din(new_net_19012),
		.dout(new_net_19013)
	);

	bfr new_net_19014_bfr_after (
		.din(new_net_19013),
		.dout(new_net_19014)
	);

	bfr new_net_19015_bfr_after (
		.din(new_net_19014),
		.dout(new_net_19015)
	);

	bfr new_net_19016_bfr_after (
		.din(new_net_19015),
		.dout(new_net_19016)
	);

	bfr new_net_19017_bfr_after (
		.din(new_net_19016),
		.dout(new_net_19017)
	);

	bfr new_net_19018_bfr_after (
		.din(new_net_19017),
		.dout(new_net_19018)
	);

	bfr new_net_19019_bfr_after (
		.din(new_net_19018),
		.dout(new_net_19019)
	);

	bfr new_net_19020_bfr_after (
		.din(new_net_19019),
		.dout(new_net_19020)
	);

	bfr new_net_19021_bfr_after (
		.din(new_net_19020),
		.dout(new_net_19021)
	);

	bfr new_net_19022_bfr_after (
		.din(new_net_19021),
		.dout(new_net_19022)
	);

	bfr new_net_19023_bfr_after (
		.din(new_net_19022),
		.dout(new_net_19023)
	);

	bfr new_net_19024_bfr_after (
		.din(new_net_19023),
		.dout(new_net_19024)
	);

	bfr new_net_19025_bfr_after (
		.din(new_net_19024),
		.dout(new_net_19025)
	);

	bfr new_net_19026_bfr_after (
		.din(new_net_19025),
		.dout(new_net_19026)
	);

	bfr new_net_19027_bfr_after (
		.din(new_net_19026),
		.dout(new_net_19027)
	);

	bfr new_net_19028_bfr_after (
		.din(new_net_19027),
		.dout(new_net_19028)
	);

	bfr new_net_19029_bfr_after (
		.din(new_net_19028),
		.dout(new_net_19029)
	);

	bfr new_net_19030_bfr_after (
		.din(new_net_19029),
		.dout(new_net_19030)
	);

	bfr new_net_19031_bfr_after (
		.din(new_net_19030),
		.dout(new_net_19031)
	);

	bfr new_net_19032_bfr_after (
		.din(new_net_19031),
		.dout(new_net_19032)
	);

	bfr new_net_19033_bfr_after (
		.din(new_net_19032),
		.dout(new_net_19033)
	);

	bfr new_net_19034_bfr_after (
		.din(new_net_19033),
		.dout(new_net_19034)
	);

	bfr new_net_19035_bfr_after (
		.din(new_net_19034),
		.dout(new_net_19035)
	);

	bfr new_net_19036_bfr_after (
		.din(new_net_19035),
		.dout(new_net_19036)
	);

	bfr new_net_19037_bfr_after (
		.din(new_net_19036),
		.dout(new_net_19037)
	);

	bfr new_net_19038_bfr_after (
		.din(new_net_19037),
		.dout(new_net_19038)
	);

	bfr new_net_19039_bfr_after (
		.din(new_net_19038),
		.dout(new_net_19039)
	);

	bfr new_net_19040_bfr_after (
		.din(new_net_19039),
		.dout(new_net_19040)
	);

	bfr new_net_19041_bfr_after (
		.din(new_net_19040),
		.dout(new_net_19041)
	);

	bfr new_net_19042_bfr_after (
		.din(new_net_19041),
		.dout(new_net_19042)
	);

	bfr new_net_19043_bfr_after (
		.din(new_net_19042),
		.dout(new_net_19043)
	);

	bfr new_net_19044_bfr_after (
		.din(new_net_19043),
		.dout(new_net_19044)
	);

	bfr new_net_19045_bfr_after (
		.din(new_net_19044),
		.dout(new_net_19045)
	);

	bfr new_net_19046_bfr_after (
		.din(new_net_19045),
		.dout(new_net_19046)
	);

	bfr new_net_19047_bfr_after (
		.din(new_net_19046),
		.dout(new_net_19047)
	);

	bfr new_net_19048_bfr_after (
		.din(new_net_19047),
		.dout(new_net_19048)
	);

	bfr new_net_19049_bfr_after (
		.din(new_net_19048),
		.dout(new_net_19049)
	);

	bfr new_net_19050_bfr_after (
		.din(new_net_19049),
		.dout(new_net_19050)
	);

	bfr new_net_19051_bfr_after (
		.din(new_net_19050),
		.dout(new_net_19051)
	);

	spl2 _1369__v_fanout (
		.a(new_net_19051),
		.b(new_net_1304),
		.c(new_net_1305)
	);

	bfr new_net_19052_bfr_after (
		.din(_0089_),
		.dout(new_net_19052)
	);

	bfr new_net_19053_bfr_after (
		.din(new_net_19052),
		.dout(new_net_19053)
	);

	bfr new_net_19054_bfr_after (
		.din(new_net_19053),
		.dout(new_net_19054)
	);

	bfr new_net_19055_bfr_after (
		.din(new_net_19054),
		.dout(new_net_19055)
	);

	bfr new_net_19056_bfr_after (
		.din(new_net_19055),
		.dout(new_net_19056)
	);

	bfr new_net_19057_bfr_after (
		.din(new_net_19056),
		.dout(new_net_19057)
	);

	bfr new_net_19058_bfr_after (
		.din(new_net_19057),
		.dout(new_net_19058)
	);

	bfr new_net_19059_bfr_after (
		.din(new_net_19058),
		.dout(new_net_19059)
	);

	bfr new_net_19060_bfr_after (
		.din(new_net_19059),
		.dout(new_net_19060)
	);

	bfr new_net_19061_bfr_after (
		.din(new_net_19060),
		.dout(new_net_19061)
	);

	bfr new_net_19062_bfr_after (
		.din(new_net_19061),
		.dout(new_net_19062)
	);

	bfr new_net_19063_bfr_after (
		.din(new_net_19062),
		.dout(new_net_19063)
	);

	bfr new_net_19064_bfr_after (
		.din(new_net_19063),
		.dout(new_net_19064)
	);

	bfr new_net_19065_bfr_after (
		.din(new_net_19064),
		.dout(new_net_19065)
	);

	bfr new_net_19066_bfr_after (
		.din(new_net_19065),
		.dout(new_net_19066)
	);

	bfr new_net_19067_bfr_after (
		.din(new_net_19066),
		.dout(new_net_19067)
	);

	bfr new_net_19068_bfr_after (
		.din(new_net_19067),
		.dout(new_net_19068)
	);

	bfr new_net_19069_bfr_after (
		.din(new_net_19068),
		.dout(new_net_19069)
	);

	bfr new_net_19070_bfr_after (
		.din(new_net_19069),
		.dout(new_net_19070)
	);

	bfr new_net_19071_bfr_after (
		.din(new_net_19070),
		.dout(new_net_19071)
	);

	bfr new_net_19072_bfr_after (
		.din(new_net_19071),
		.dout(new_net_19072)
	);

	bfr new_net_19073_bfr_after (
		.din(new_net_19072),
		.dout(new_net_19073)
	);

	bfr new_net_19074_bfr_after (
		.din(new_net_19073),
		.dout(new_net_19074)
	);

	bfr new_net_19075_bfr_after (
		.din(new_net_19074),
		.dout(new_net_19075)
	);

	bfr new_net_19076_bfr_after (
		.din(new_net_19075),
		.dout(new_net_19076)
	);

	bfr new_net_19077_bfr_after (
		.din(new_net_19076),
		.dout(new_net_19077)
	);

	bfr new_net_19078_bfr_after (
		.din(new_net_19077),
		.dout(new_net_19078)
	);

	bfr new_net_19079_bfr_after (
		.din(new_net_19078),
		.dout(new_net_19079)
	);

	bfr new_net_19080_bfr_after (
		.din(new_net_19079),
		.dout(new_net_19080)
	);

	bfr new_net_19081_bfr_after (
		.din(new_net_19080),
		.dout(new_net_19081)
	);

	bfr new_net_19082_bfr_after (
		.din(new_net_19081),
		.dout(new_net_19082)
	);

	bfr new_net_19083_bfr_after (
		.din(new_net_19082),
		.dout(new_net_19083)
	);

	bfr new_net_19084_bfr_after (
		.din(new_net_19083),
		.dout(new_net_19084)
	);

	bfr new_net_19085_bfr_after (
		.din(new_net_19084),
		.dout(new_net_19085)
	);

	bfr new_net_19086_bfr_after (
		.din(new_net_19085),
		.dout(new_net_19086)
	);

	bfr new_net_19087_bfr_after (
		.din(new_net_19086),
		.dout(new_net_19087)
	);

	bfr new_net_19088_bfr_after (
		.din(new_net_19087),
		.dout(new_net_19088)
	);

	bfr new_net_19089_bfr_after (
		.din(new_net_19088),
		.dout(new_net_19089)
	);

	bfr new_net_19090_bfr_after (
		.din(new_net_19089),
		.dout(new_net_19090)
	);

	bfr new_net_19091_bfr_after (
		.din(new_net_19090),
		.dout(new_net_19091)
	);

	bfr new_net_19092_bfr_after (
		.din(new_net_19091),
		.dout(new_net_19092)
	);

	bfr new_net_19093_bfr_after (
		.din(new_net_19092),
		.dout(new_net_19093)
	);

	bfr new_net_19094_bfr_after (
		.din(new_net_19093),
		.dout(new_net_19094)
	);

	bfr new_net_19095_bfr_after (
		.din(new_net_19094),
		.dout(new_net_19095)
	);

	bfr new_net_19096_bfr_after (
		.din(new_net_19095),
		.dout(new_net_19096)
	);

	bfr new_net_19097_bfr_after (
		.din(new_net_19096),
		.dout(new_net_19097)
	);

	bfr new_net_19098_bfr_after (
		.din(new_net_19097),
		.dout(new_net_19098)
	);

	bfr new_net_19099_bfr_after (
		.din(new_net_19098),
		.dout(new_net_19099)
	);

	bfr new_net_19100_bfr_after (
		.din(new_net_19099),
		.dout(new_net_19100)
	);

	bfr new_net_19101_bfr_after (
		.din(new_net_19100),
		.dout(new_net_19101)
	);

	bfr new_net_19102_bfr_after (
		.din(new_net_19101),
		.dout(new_net_19102)
	);

	bfr new_net_19103_bfr_after (
		.din(new_net_19102),
		.dout(new_net_19103)
	);

	bfr new_net_19104_bfr_after (
		.din(new_net_19103),
		.dout(new_net_19104)
	);

	bfr new_net_19105_bfr_after (
		.din(new_net_19104),
		.dout(new_net_19105)
	);

	bfr new_net_19106_bfr_after (
		.din(new_net_19105),
		.dout(new_net_19106)
	);

	bfr new_net_19107_bfr_after (
		.din(new_net_19106),
		.dout(new_net_19107)
	);

	bfr new_net_19108_bfr_after (
		.din(new_net_19107),
		.dout(new_net_19108)
	);

	bfr new_net_19109_bfr_after (
		.din(new_net_19108),
		.dout(new_net_19109)
	);

	bfr new_net_19110_bfr_after (
		.din(new_net_19109),
		.dout(new_net_19110)
	);

	bfr new_net_19111_bfr_after (
		.din(new_net_19110),
		.dout(new_net_19111)
	);

	bfr new_net_19112_bfr_after (
		.din(new_net_19111),
		.dout(new_net_19112)
	);

	bfr new_net_19113_bfr_after (
		.din(new_net_19112),
		.dout(new_net_19113)
	);

	bfr new_net_19114_bfr_after (
		.din(new_net_19113),
		.dout(new_net_19114)
	);

	bfr new_net_19115_bfr_after (
		.din(new_net_19114),
		.dout(new_net_19115)
	);

	bfr new_net_19116_bfr_after (
		.din(new_net_19115),
		.dout(new_net_19116)
	);

	bfr new_net_19117_bfr_after (
		.din(new_net_19116),
		.dout(new_net_19117)
	);

	bfr new_net_19118_bfr_after (
		.din(new_net_19117),
		.dout(new_net_19118)
	);

	bfr new_net_19119_bfr_after (
		.din(new_net_19118),
		.dout(new_net_19119)
	);

	bfr new_net_19120_bfr_after (
		.din(new_net_19119),
		.dout(new_net_19120)
	);

	bfr new_net_19121_bfr_after (
		.din(new_net_19120),
		.dout(new_net_19121)
	);

	bfr new_net_19122_bfr_after (
		.din(new_net_19121),
		.dout(new_net_19122)
	);

	bfr new_net_19123_bfr_after (
		.din(new_net_19122),
		.dout(new_net_19123)
	);

	bfr new_net_19124_bfr_after (
		.din(new_net_19123),
		.dout(new_net_19124)
	);

	bfr new_net_19125_bfr_after (
		.din(new_net_19124),
		.dout(new_net_19125)
	);

	bfr new_net_19126_bfr_after (
		.din(new_net_19125),
		.dout(new_net_19126)
	);

	bfr new_net_19127_bfr_after (
		.din(new_net_19126),
		.dout(new_net_19127)
	);

	bfr new_net_19128_bfr_after (
		.din(new_net_19127),
		.dout(new_net_19128)
	);

	bfr new_net_19129_bfr_after (
		.din(new_net_19128),
		.dout(new_net_19129)
	);

	bfr new_net_19130_bfr_after (
		.din(new_net_19129),
		.dout(new_net_19130)
	);

	bfr new_net_19131_bfr_after (
		.din(new_net_19130),
		.dout(new_net_19131)
	);

	bfr new_net_19132_bfr_after (
		.din(new_net_19131),
		.dout(new_net_19132)
	);

	bfr new_net_19133_bfr_after (
		.din(new_net_19132),
		.dout(new_net_19133)
	);

	bfr new_net_19134_bfr_after (
		.din(new_net_19133),
		.dout(new_net_19134)
	);

	bfr new_net_19135_bfr_after (
		.din(new_net_19134),
		.dout(new_net_19135)
	);

	bfr new_net_19136_bfr_after (
		.din(new_net_19135),
		.dout(new_net_19136)
	);

	bfr new_net_19137_bfr_after (
		.din(new_net_19136),
		.dout(new_net_19137)
	);

	bfr new_net_19138_bfr_after (
		.din(new_net_19137),
		.dout(new_net_19138)
	);

	bfr new_net_19139_bfr_after (
		.din(new_net_19138),
		.dout(new_net_19139)
	);

	bfr new_net_19140_bfr_after (
		.din(new_net_19139),
		.dout(new_net_19140)
	);

	bfr new_net_19141_bfr_after (
		.din(new_net_19140),
		.dout(new_net_19141)
	);

	bfr new_net_19142_bfr_after (
		.din(new_net_19141),
		.dout(new_net_19142)
	);

	bfr new_net_19143_bfr_after (
		.din(new_net_19142),
		.dout(new_net_19143)
	);

	bfr new_net_19144_bfr_after (
		.din(new_net_19143),
		.dout(new_net_19144)
	);

	bfr new_net_19145_bfr_after (
		.din(new_net_19144),
		.dout(new_net_19145)
	);

	bfr new_net_19146_bfr_after (
		.din(new_net_19145),
		.dout(new_net_19146)
	);

	bfr new_net_19147_bfr_after (
		.din(new_net_19146),
		.dout(new_net_19147)
	);

	bfr new_net_19148_bfr_after (
		.din(new_net_19147),
		.dout(new_net_19148)
	);

	spl2 _0089__v_fanout (
		.a(new_net_19148),
		.b(new_net_2857),
		.c(new_net_2858)
	);

	bfr new_net_19149_bfr_after (
		.din(_1143_),
		.dout(new_net_19149)
	);

	spl2 _1143__v_fanout (
		.a(new_net_19149),
		.b(new_net_1368),
		.c(new_net_1369)
	);

	bfr new_net_19150_bfr_after (
		.din(_1286_),
		.dout(new_net_19150)
	);

	bfr new_net_19151_bfr_after (
		.din(new_net_19150),
		.dout(new_net_19151)
	);

	bfr new_net_19152_bfr_after (
		.din(new_net_19151),
		.dout(new_net_19152)
	);

	bfr new_net_19153_bfr_after (
		.din(new_net_19152),
		.dout(new_net_19153)
	);

	bfr new_net_19154_bfr_after (
		.din(new_net_19153),
		.dout(new_net_19154)
	);

	bfr new_net_19155_bfr_after (
		.din(new_net_19154),
		.dout(new_net_19155)
	);

	bfr new_net_19156_bfr_after (
		.din(new_net_19155),
		.dout(new_net_19156)
	);

	bfr new_net_19157_bfr_after (
		.din(new_net_19156),
		.dout(new_net_19157)
	);

	bfr new_net_19158_bfr_after (
		.din(new_net_19157),
		.dout(new_net_19158)
	);

	bfr new_net_19159_bfr_after (
		.din(new_net_19158),
		.dout(new_net_19159)
	);

	bfr new_net_19160_bfr_after (
		.din(new_net_19159),
		.dout(new_net_19160)
	);

	bfr new_net_19161_bfr_after (
		.din(new_net_19160),
		.dout(new_net_19161)
	);

	bfr new_net_19162_bfr_after (
		.din(new_net_19161),
		.dout(new_net_19162)
	);

	bfr new_net_19163_bfr_after (
		.din(new_net_19162),
		.dout(new_net_19163)
	);

	bfr new_net_19164_bfr_after (
		.din(new_net_19163),
		.dout(new_net_19164)
	);

	bfr new_net_19165_bfr_after (
		.din(new_net_19164),
		.dout(new_net_19165)
	);

	bfr new_net_19166_bfr_after (
		.din(new_net_19165),
		.dout(new_net_19166)
	);

	bfr new_net_19167_bfr_after (
		.din(new_net_19166),
		.dout(new_net_19167)
	);

	bfr new_net_19168_bfr_after (
		.din(new_net_19167),
		.dout(new_net_19168)
	);

	bfr new_net_19169_bfr_after (
		.din(new_net_19168),
		.dout(new_net_19169)
	);

	bfr new_net_19170_bfr_after (
		.din(new_net_19169),
		.dout(new_net_19170)
	);

	bfr new_net_19171_bfr_after (
		.din(new_net_19170),
		.dout(new_net_19171)
	);

	bfr new_net_19172_bfr_after (
		.din(new_net_19171),
		.dout(new_net_19172)
	);

	bfr new_net_19173_bfr_after (
		.din(new_net_19172),
		.dout(new_net_19173)
	);

	bfr new_net_19174_bfr_after (
		.din(new_net_19173),
		.dout(new_net_19174)
	);

	bfr new_net_19175_bfr_after (
		.din(new_net_19174),
		.dout(new_net_19175)
	);

	bfr new_net_19176_bfr_after (
		.din(new_net_19175),
		.dout(new_net_19176)
	);

	bfr new_net_19177_bfr_after (
		.din(new_net_19176),
		.dout(new_net_19177)
	);

	bfr new_net_19178_bfr_after (
		.din(new_net_19177),
		.dout(new_net_19178)
	);

	bfr new_net_19179_bfr_after (
		.din(new_net_19178),
		.dout(new_net_19179)
	);

	bfr new_net_19180_bfr_after (
		.din(new_net_19179),
		.dout(new_net_19180)
	);

	bfr new_net_19181_bfr_after (
		.din(new_net_19180),
		.dout(new_net_19181)
	);

	bfr new_net_19182_bfr_after (
		.din(new_net_19181),
		.dout(new_net_19182)
	);

	bfr new_net_19183_bfr_after (
		.din(new_net_19182),
		.dout(new_net_19183)
	);

	bfr new_net_19184_bfr_after (
		.din(new_net_19183),
		.dout(new_net_19184)
	);

	bfr new_net_19185_bfr_after (
		.din(new_net_19184),
		.dout(new_net_19185)
	);

	bfr new_net_19186_bfr_after (
		.din(new_net_19185),
		.dout(new_net_19186)
	);

	bfr new_net_19187_bfr_after (
		.din(new_net_19186),
		.dout(new_net_19187)
	);

	bfr new_net_19188_bfr_after (
		.din(new_net_19187),
		.dout(new_net_19188)
	);

	bfr new_net_19189_bfr_after (
		.din(new_net_19188),
		.dout(new_net_19189)
	);

	bfr new_net_19190_bfr_after (
		.din(new_net_19189),
		.dout(new_net_19190)
	);

	bfr new_net_19191_bfr_after (
		.din(new_net_19190),
		.dout(new_net_19191)
	);

	bfr new_net_19192_bfr_after (
		.din(new_net_19191),
		.dout(new_net_19192)
	);

	bfr new_net_19193_bfr_after (
		.din(new_net_19192),
		.dout(new_net_19193)
	);

	bfr new_net_19194_bfr_after (
		.din(new_net_19193),
		.dout(new_net_19194)
	);

	bfr new_net_19195_bfr_after (
		.din(new_net_19194),
		.dout(new_net_19195)
	);

	bfr new_net_19196_bfr_after (
		.din(new_net_19195),
		.dout(new_net_19196)
	);

	bfr new_net_19197_bfr_after (
		.din(new_net_19196),
		.dout(new_net_19197)
	);

	bfr new_net_19198_bfr_after (
		.din(new_net_19197),
		.dout(new_net_19198)
	);

	spl2 _1286__v_fanout (
		.a(new_net_19198),
		.b(new_net_1580),
		.c(new_net_1581)
	);

	bfr new_net_19199_bfr_after (
		.din(_0731_),
		.dout(new_net_19199)
	);

	bfr new_net_19200_bfr_after (
		.din(new_net_19199),
		.dout(new_net_19200)
	);

	bfr new_net_19201_bfr_after (
		.din(new_net_19200),
		.dout(new_net_19201)
	);

	bfr new_net_19202_bfr_after (
		.din(new_net_19201),
		.dout(new_net_19202)
	);

	bfr new_net_19203_bfr_after (
		.din(new_net_19202),
		.dout(new_net_19203)
	);

	bfr new_net_19204_bfr_after (
		.din(new_net_19203),
		.dout(new_net_19204)
	);

	bfr new_net_19205_bfr_after (
		.din(new_net_19204),
		.dout(new_net_19205)
	);

	bfr new_net_19206_bfr_after (
		.din(new_net_19205),
		.dout(new_net_19206)
	);

	bfr new_net_19207_bfr_after (
		.din(new_net_19206),
		.dout(new_net_19207)
	);

	spl2 _0731__v_fanout (
		.a(new_net_19207),
		.b(new_net_126),
		.c(new_net_127)
	);

	spl4L new_net_3434_v_fanout (
		.a(new_net_3434),
		.b(new_net_263),
		.c(new_net_271),
		.d(new_net_269),
		.e(new_net_261)
	);

	spl4L new_net_3428_v_fanout (
		.a(new_net_3428),
		.b(new_net_2047),
		.c(new_net_2056),
		.d(new_net_2046),
		.e(new_net_2057)
	);

	spl4L new_net_3396_v_fanout (
		.a(new_net_3396),
		.b(new_net_2490),
		.c(new_net_2491),
		.d(new_net_2500),
		.e(new_net_2496)
	);

	bfr new_net_19208_bfr_before (
		.din(new_net_19208),
		.dout(new_net_2870)
	);

	bfr new_net_19209_bfr_before (
		.din(new_net_19209),
		.dout(new_net_19208)
	);

	bfr new_net_19210_bfr_before (
		.din(new_net_19210),
		.dout(new_net_19209)
	);

	bfr new_net_19211_bfr_before (
		.din(new_net_19211),
		.dout(new_net_19210)
	);

	bfr new_net_19212_bfr_before (
		.din(new_net_19212),
		.dout(new_net_19211)
	);

	spl4L new_net_3355_v_fanout (
		.a(new_net_3355),
		.b(new_net_19212),
		.c(new_net_2867),
		.d(new_net_2862),
		.e(new_net_2875)
	);

	spl4L new_net_3381_v_fanout (
		.a(new_net_3381),
		.b(new_net_740),
		.c(new_net_748),
		.d(new_net_752),
		.e(new_net_745)
	);

	spl4L new_net_3328_v_fanout (
		.a(new_net_3328),
		.b(new_net_927),
		.c(new_net_916),
		.d(new_net_930),
		.e(new_net_924)
	);

	spl3L new_net_3318_v_fanout (
		.a(new_net_3318),
		.b(new_net_426),
		.c(new_net_441),
		.d(new_net_431)
	);

	spl4L new_net_3385_v_fanout (
		.a(new_net_3385),
		.b(new_net_3245),
		.c(new_net_3246),
		.d(new_net_3235),
		.e(new_net_3234)
	);

	spl4L new_net_3362_v_fanout (
		.a(new_net_3362),
		.b(new_net_3077),
		.c(new_net_3087),
		.d(new_net_3092),
		.e(new_net_3089)
	);

	spl4L new_net_3371_v_fanout (
		.a(new_net_3371),
		.b(new_net_541),
		.c(new_net_540),
		.d(new_net_529),
		.e(new_net_533)
	);

	spl3L new_net_3308_v_fanout (
		.a(new_net_3308),
		.b(new_net_3022),
		.c(new_net_3011),
		.d(new_net_3024)
	);

	spl4L new_net_3416_v_fanout (
		.a(new_net_3416),
		.b(new_net_1129),
		.c(new_net_1118),
		.d(new_net_1124),
		.e(new_net_1116)
	);

	spl3L new_net_3410_v_fanout (
		.a(new_net_3410),
		.b(new_net_1807),
		.c(new_net_1810),
		.d(new_net_1808)
	);

	spl2 new_net_3407_v_fanout (
		.a(new_net_3407),
		.b(new_net_1798),
		.c(new_net_1800)
	);

	spl4L new_net_3367_v_fanout (
		.a(new_net_3367),
		.b(new_net_2410),
		.c(new_net_2403),
		.d(new_net_2405),
		.e(new_net_2398)
	);

	spl4L new_net_3338_v_fanout (
		.a(new_net_3338),
		.b(new_net_395),
		.c(new_net_392),
		.d(new_net_398),
		.e(new_net_396)
	);

	spl3L new_net_3365_v_fanout (
		.a(new_net_3365),
		.b(new_net_2397),
		.c(new_net_2399),
		.d(new_net_2396)
	);

	spl4L new_net_3421_v_fanout (
		.a(new_net_3421),
		.b(new_net_42),
		.c(new_net_44),
		.d(new_net_39),
		.e(new_net_43)
	);

	spl4L new_net_3366_v_fanout (
		.a(new_net_3366),
		.b(new_net_2400),
		.c(new_net_2402),
		.d(new_net_2404),
		.e(new_net_2409)
	);

	spl4L new_net_3324_v_fanout (
		.a(new_net_3324),
		.b(new_net_2339),
		.c(new_net_2344),
		.d(new_net_2340),
		.e(new_net_2341)
	);

	spl3L new_net_3398_v_fanout (
		.a(new_net_3398),
		.b(new_net_2498),
		.c(new_net_2497),
		.d(new_net_2499)
	);

	spl3L new_net_3313_v_fanout (
		.a(new_net_3313),
		.b(new_net_2913),
		.c(new_net_2922),
		.d(new_net_2919)
	);

	spl3L new_net_3360_v_fanout (
		.a(new_net_3360),
		.b(new_net_3078),
		.c(new_net_3086),
		.d(new_net_3084)
	);

	spl4L new_net_3414_v_fanout (
		.a(new_net_3414),
		.b(new_net_1117),
		.c(new_net_1121),
		.d(new_net_1120),
		.e(new_net_1119)
	);

	spl4L new_net_3370_v_fanout (
		.a(new_net_3370),
		.b(new_net_539),
		.c(new_net_535),
		.d(new_net_530),
		.e(new_net_532)
	);

	spl4L new_net_3375_v_fanout (
		.a(new_net_3375),
		.b(new_net_1473),
		.c(new_net_1480),
		.d(new_net_1475),
		.e(new_net_1470)
	);

	spl2 new_net_3419_v_fanout (
		.a(new_net_3419),
		.b(new_net_49),
		.c(new_net_50)
	);

	spl4L new_net_3376_v_fanout (
		.a(new_net_3376),
		.b(new_net_1479),
		.c(new_net_1472),
		.d(new_net_1471),
		.e(new_net_1474)
	);

	spl4L new_net_3422_v_fanout (
		.a(new_net_3422),
		.b(new_net_37),
		.c(new_net_48),
		.d(new_net_38),
		.e(new_net_46)
	);

	spl3L new_net_3303_v_fanout (
		.a(new_net_3303),
		.b(new_net_1249),
		.c(new_net_1245),
		.d(new_net_1260)
	);

	bfr new_net_19213_bfr_before (
		.din(new_net_19213),
		.dout(new_net_2697)
	);

	bfr new_net_19214_bfr_before (
		.din(new_net_19214),
		.dout(new_net_19213)
	);

	spl2 new_net_3288_v_fanout (
		.a(new_net_3288),
		.b(new_net_19214),
		.c(new_net_2712)
	);

	spl4L new_net_3432_v_fanout (
		.a(new_net_3432),
		.b(new_net_258),
		.c(new_net_265),
		.d(new_net_260),
		.e(new_net_259)
	);

	spl3L new_net_3431_v_fanout (
		.a(new_net_3431),
		.b(new_net_272),
		.c(new_net_264),
		.d(new_net_262)
	);

	spl4L new_net_3333_v_fanout (
		.a(new_net_3333),
		.b(new_net_3178),
		.c(new_net_3177),
		.d(new_net_3182),
		.e(new_net_3180)
	);

	spl3L new_net_3425_v_fanout (
		.a(new_net_3425),
		.b(new_net_2052),
		.c(new_net_2050),
		.d(new_net_2054)
	);

	spl3L new_net_3323_v_fanout (
		.a(new_net_3323),
		.b(new_net_2346),
		.c(new_net_2351),
		.d(new_net_2354)
	);

	spl4L new_net_3344_v_fanout (
		.a(new_net_3344),
		.b(new_net_1550),
		.c(new_net_1557),
		.d(new_net_1546),
		.e(new_net_1548)
	);

	spl4L new_net_3415_v_fanout (
		.a(new_net_3415),
		.b(new_net_1125),
		.c(new_net_1126),
		.d(new_net_1123),
		.e(new_net_1127)
	);

	spl4L new_net_3408_v_fanout (
		.a(new_net_3408),
		.b(new_net_1796),
		.c(new_net_1801),
		.d(new_net_1802),
		.e(new_net_1806)
	);

	spl4L new_net_3427_v_fanout (
		.a(new_net_3427),
		.b(new_net_2049),
		.c(new_net_2051),
		.d(new_net_2055),
		.e(new_net_2044)
	);

	spl2 new_net_3349_v_fanout (
		.a(new_net_3349),
		.b(new_net_1442),
		.c(new_net_1453)
	);

	spl2 new_net_3343_v_fanout (
		.a(new_net_3343),
		.b(new_net_1552),
		.c(new_net_1559)
	);

	spl4L new_net_3426_v_fanout (
		.a(new_net_3426),
		.b(new_net_2042),
		.c(new_net_2048),
		.d(new_net_2045),
		.e(new_net_2043)
	);

	spl4L new_net_3392_v_fanout (
		.a(new_net_3392),
		.b(new_net_209),
		.c(new_net_215),
		.d(new_net_200),
		.e(new_net_214)
	);

	spl4L new_net_3403_v_fanout (
		.a(new_net_3403),
		.b(new_net_2554),
		.c(new_net_2562),
		.d(new_net_2547),
		.e(new_net_2561)
	);

	spl2 new_net_3401_v_fanout (
		.a(new_net_3401),
		.b(new_net_2557),
		.c(new_net_2560)
	);

	spl4L new_net_3386_v_fanout (
		.a(new_net_3386),
		.b(new_net_3244),
		.c(new_net_3232),
		.d(new_net_3241),
		.e(new_net_3242)
	);

	spl4L new_net_3356_v_fanout (
		.a(new_net_3356),
		.b(new_net_2861),
		.c(new_net_2873),
		.d(new_net_2863),
		.e(new_net_2872)
	);

	spl4L new_net_3402_v_fanout (
		.a(new_net_3402),
		.b(new_net_2558),
		.c(new_net_2552),
		.d(new_net_2556),
		.e(new_net_2559)
	);

	spl4L new_net_3433_v_fanout (
		.a(new_net_3433),
		.b(new_net_268),
		.c(new_net_257),
		.d(new_net_270),
		.e(new_net_267)
	);

	spl4L new_net_3380_v_fanout (
		.a(new_net_3380),
		.b(new_net_747),
		.c(new_net_751),
		.d(new_net_737),
		.e(new_net_749)
	);

	spl4L new_net_3361_v_fanout (
		.a(new_net_3361),
		.b(new_net_3085),
		.c(new_net_3080),
		.d(new_net_3079),
		.e(new_net_3090)
	);

	spl3L new_net_3390_v_fanout (
		.a(new_net_3390),
		.b(new_net_203),
		.c(new_net_205),
		.d(new_net_202)
	);

	spl4L new_net_3345_v_fanout (
		.a(new_net_3345),
		.b(new_net_1554),
		.c(new_net_1556),
		.d(new_net_1551),
		.e(new_net_1545)
	);

	spl3L new_net_3293_v_fanout (
		.a(new_net_3293),
		.b(new_net_2605),
		.c(new_net_2611),
		.d(new_net_2617)
	);

	spl4L new_net_3382_v_fanout (
		.a(new_net_3382),
		.b(new_net_739),
		.c(new_net_738),
		.d(new_net_741),
		.e(new_net_746)
	);

	spl2 new_net_3413_v_fanout (
		.a(new_net_3413),
		.b(new_net_1128),
		.c(new_net_1131)
	);

	spl3L new_net_3298_v_fanout (
		.a(new_net_3298),
		.b(new_net_161),
		.c(new_net_154),
		.d(new_net_146)
	);

	spl3L new_net_3350_v_fanout (
		.a(new_net_3350),
		.b(new_net_1449),
		.c(new_net_1448),
		.d(new_net_1444)
	);

	spl2 new_net_3395_v_fanout (
		.a(new_net_3395),
		.b(new_net_2502),
		.c(new_net_2494)
	);

	spl3L new_net_3404_v_fanout (
		.a(new_net_3404),
		.b(new_net_2551),
		.c(new_net_2549),
		.d(new_net_2555)
	);

	spl4L new_net_3397_v_fanout (
		.a(new_net_3397),
		.b(new_net_2503),
		.c(new_net_2493),
		.d(new_net_2504),
		.e(new_net_2505)
	);

	spl4L new_net_3409_v_fanout (
		.a(new_net_3409),
		.b(new_net_1799),
		.c(new_net_1805),
		.d(new_net_1803),
		.e(new_net_1797)
	);

	spl4L new_net_3357_v_fanout (
		.a(new_net_3357),
		.b(new_net_2877),
		.c(new_net_2876),
		.d(new_net_2868),
		.e(new_net_2874)
	);

	spl4L new_net_3420_v_fanout (
		.a(new_net_3420),
		.b(new_net_36),
		.c(new_net_45),
		.d(new_net_51),
		.e(new_net_47)
	);

	spl4L new_net_3387_v_fanout (
		.a(new_net_3387),
		.b(new_net_3238),
		.c(new_net_3239),
		.d(new_net_3243),
		.e(new_net_3240)
	);

	spl4L new_net_3391_v_fanout (
		.a(new_net_3391),
		.b(new_net_211),
		.c(new_net_201),
		.d(new_net_212),
		.e(new_net_204)
	);

	spl4L new_net_3377_v_fanout (
		.a(new_net_3377),
		.b(new_net_1483),
		.c(new_net_1481),
		.d(new_net_1484),
		.e(new_net_1469)
	);

	spl4L new_net_3285_v_fanout (
		.a(new_net_3285),
		.b(new_net_2831),
		.c(new_net_2835),
		.d(new_net_2838),
		.e(new_net_2841)
	);

	spl3L new_net_3337_v_fanout (
		.a(new_net_3337),
		.b(new_net_3192),
		.c(new_net_3191),
		.d(new_net_3185)
	);

	bfr new_net_19215_bfr_before (
		.din(new_net_19215),
		.dout(new_net_2550)
	);

	bfr new_net_19216_bfr_before (
		.din(new_net_19216),
		.dout(new_net_2548)
	);

	spl4L new_net_3406_v_fanout (
		.a(new_net_3406),
		.b(new_net_19215),
		.c(new_net_3404),
		.d(new_net_3403),
		.e(new_net_19216)
	);

	spl3L new_net_3332_v_fanout (
		.a(new_net_3332),
		.b(new_net_918),
		.c(new_net_919),
		.d(new_net_921)
	);

	spl4L new_net_3317_v_fanout (
		.a(new_net_3317),
		.b(new_net_2916),
		.c(new_net_2918),
		.d(new_net_2920),
		.e(new_net_2917)
	);

	bfr new_net_19217_bfr_before (
		.din(new_net_19217),
		.dout(new_net_2701)
	);

	bfr new_net_19218_bfr_before (
		.din(new_net_19218),
		.dout(new_net_2698)
	);

	bfr new_net_19219_bfr_before (
		.din(new_net_19219),
		.dout(new_net_2702)
	);

	spl4L new_net_3291_v_fanout (
		.a(new_net_3291),
		.b(new_net_3288),
		.c(new_net_19219),
		.d(new_net_19218),
		.e(new_net_19217)
	);

	spl2 new_net_3435_v_fanout (
		.a(new_net_3435),
		.b(new_net_3433),
		.c(new_net_3431)
	);

	bfr new_net_19220_bfr_before (
		.din(new_net_19220),
		.dout(new_net_1547)
	);

	bfr new_net_19221_bfr_before (
		.din(new_net_19221),
		.dout(new_net_1555)
	);

	spl4L new_net_3347_v_fanout (
		.a(new_net_3347),
		.b(new_net_3345),
		.c(new_net_3343),
		.d(new_net_19221),
		.e(new_net_19220)
	);

	spl4L new_net_3305_v_fanout (
		.a(new_net_3305),
		.b(new_net_1256),
		.c(new_net_1246),
		.d(new_net_1254),
		.e(new_net_1257)
	);

	bfr new_net_19222_bfr_before (
		.din(new_net_19222),
		.dout(new_net_40)
	);

	spl2 new_net_3423_v_fanout (
		.a(new_net_3423),
		.b(new_net_19222),
		.c(new_net_3419)
	);

	spl4L new_net_3424_v_fanout (
		.a(new_net_3424),
		.b(new_net_3421),
		.c(new_net_41),
		.d(new_net_3420),
		.e(new_net_3422)
	);

	bfr new_net_19223_bfr_before (
		.din(new_net_19223),
		.dout(new_net_1122)
	);

	spl4L new_net_3418_v_fanout (
		.a(new_net_3418),
		.b(new_net_19223),
		.c(new_net_3416),
		.d(new_net_3413),
		.e(new_net_3415)
	);

	spl4L new_net_3340_v_fanout (
		.a(new_net_3340),
		.b(new_net_393),
		.c(new_net_394),
		.d(new_net_402),
		.e(new_net_404)
	);

	bfr new_net_19224_bfr_before (
		.din(new_net_19224),
		.dout(new_net_3026)
	);

	bfr new_net_19225_bfr_before (
		.din(new_net_19225),
		.dout(new_net_3014)
	);

	bfr new_net_19226_bfr_before (
		.din(new_net_19226),
		.dout(new_net_3017)
	);

	spl4L new_net_3312_v_fanout (
		.a(new_net_3312),
		.b(new_net_19224),
		.c(new_net_19226),
		.d(new_net_3308),
		.e(new_net_19225)
	);

	spl4L new_net_3310_v_fanout (
		.a(new_net_3310),
		.b(new_net_3021),
		.c(new_net_3015),
		.d(new_net_3020),
		.e(new_net_3023)
	);

	bfr new_net_19227_bfr_before (
		.din(new_net_19227),
		.dout(new_net_2553)
	);

	spl3L new_net_3405_v_fanout (
		.a(new_net_3405),
		.b(new_net_3402),
		.c(new_net_3401),
		.d(new_net_19227)
	);

	spl4L new_net_3287_v_fanout (
		.a(new_net_3287),
		.b(new_net_2843),
		.c(new_net_2830),
		.d(new_net_2834),
		.e(new_net_2837)
	);

	spl4L new_net_3315_v_fanout (
		.a(new_net_3315),
		.b(new_net_2909),
		.c(new_net_2912),
		.d(new_net_2907),
		.e(new_net_2915)
	);

	bfr new_net_19228_bfr_before (
		.din(new_net_19228),
		.dout(new_net_2053)
	);

	spl3L new_net_3430_v_fanout (
		.a(new_net_3430),
		.b(new_net_3428),
		.c(new_net_3426),
		.d(new_net_19228)
	);

	bfr new_net_19229_bfr_before (
		.din(new_net_19229),
		.dout(new_net_1476)
	);

	bfr new_net_19230_bfr_before (
		.din(new_net_19230),
		.dout(new_net_1478)
	);

	spl4L new_net_3379_v_fanout (
		.a(new_net_3379),
		.b(new_net_19229),
		.c(new_net_3377),
		.d(new_net_3375),
		.e(new_net_19230)
	);

	spl4L new_net_3277_v_fanout (
		.a(new_net_3277),
		.b(new_net_379),
		.c(new_net_386),
		.d(new_net_387),
		.e(new_net_388)
	);

	bfr new_net_19231_bfr_before (
		.din(new_net_19231),
		.dout(new_net_2492)
	);

	bfr new_net_19232_bfr_before (
		.din(new_net_19232),
		.dout(new_net_2501)
	);

	bfr new_net_19233_bfr_before (
		.din(new_net_19233),
		.dout(new_net_2495)
	);

	spl4L new_net_3400_v_fanout (
		.a(new_net_3400),
		.b(new_net_3398),
		.c(new_net_19233),
		.d(new_net_19232),
		.e(new_net_19231)
	);

	bfr new_net_19234_bfr_before (
		.din(new_net_19234),
		.dout(new_net_2910)
	);

	bfr new_net_19235_bfr_before (
		.din(new_net_19235),
		.dout(new_net_2914)
	);

	bfr new_net_19236_bfr_before (
		.din(new_net_19236),
		.dout(new_net_2911)
	);

	spl4L new_net_3316_v_fanout (
		.a(new_net_3316),
		.b(new_net_19234),
		.c(new_net_2908),
		.d(new_net_19236),
		.e(new_net_19235)
	);

	spl4L new_net_3437_v_fanout (
		.a(new_net_3437),
		.b(new_net_1420),
		.c(new_net_1415),
		.d(new_net_1413),
		.e(new_net_1409)
	);

	bfr new_net_19237_bfr_before (
		.din(new_net_19237),
		.dout(new_net_2608)
	);

	bfr new_net_19238_bfr_before (
		.din(new_net_19238),
		.dout(new_net_2616)
	);

	spl4L new_net_3297_v_fanout (
		.a(new_net_3297),
		.b(new_net_2615),
		.c(new_net_19238),
		.d(new_net_3293),
		.e(new_net_19237)
	);

	bfr new_net_19239_bfr_before (
		.din(new_net_19239),
		.dout(new_net_1251)
	);

	spl2 new_net_3304_v_fanout (
		.a(new_net_3304),
		.b(new_net_1259),
		.c(new_net_19239)
	);

	bfr new_net_19240_bfr_before (
		.din(new_net_19240),
		.dout(new_net_434)
	);

	bfr new_net_19241_bfr_before (
		.din(new_net_19241),
		.dout(new_net_437)
	);

	bfr new_net_19242_bfr_before (
		.din(new_net_19242),
		.dout(new_net_435)
	);

	spl4L new_net_3320_v_fanout (
		.a(new_net_3320),
		.b(new_net_19240),
		.c(new_net_19242),
		.d(new_net_436),
		.e(new_net_19241)
	);

	spl4L new_net_3307_v_fanout (
		.a(new_net_3307),
		.b(new_net_1247),
		.c(new_net_1258),
		.d(new_net_1255),
		.e(new_net_1248)
	);

	bfr new_net_19243_bfr_before (
		.din(new_net_19243),
		.dout(new_net_2350)
	);

	bfr new_net_19244_bfr_before (
		.din(new_net_19244),
		.dout(new_net_2345)
	);

	bfr new_net_19245_bfr_before (
		.din(new_net_19245),
		.dout(new_net_2349)
	);

	spl4L new_net_3326_v_fanout (
		.a(new_net_3326),
		.b(new_net_19243),
		.c(new_net_3324),
		.d(new_net_19245),
		.e(new_net_19244)
	);

	bfr new_net_19246_bfr_before (
		.din(new_net_19246),
		.dout(new_net_527)
	);

	spl2 new_net_3372_v_fanout (
		.a(new_net_3372),
		.b(new_net_19246),
		.c(new_net_531)
	);

	spl2 new_net_3429_v_fanout (
		.a(new_net_3429),
		.b(new_net_3425),
		.c(new_net_3427)
	);

	spl3L new_net_3399_v_fanout (
		.a(new_net_3399),
		.b(new_net_3395),
		.c(new_net_3397),
		.d(new_net_3396)
	);

	spl2 new_net_3339_v_fanout (
		.a(new_net_3339),
		.b(new_net_400),
		.c(new_net_406)
	);

	spl4L new_net_3292_v_fanout (
		.a(new_net_3292),
		.b(new_net_2699),
		.c(new_net_2703),
		.d(new_net_2706),
		.e(new_net_2704)
	);

	bfr new_net_19247_bfr_before (
		.din(new_net_19247),
		.dout(new_net_156)
	);

	spl2 new_net_3299_v_fanout (
		.a(new_net_3299),
		.b(new_net_19247),
		.c(new_net_157)
	);

	bfr new_net_19248_bfr_before (
		.din(new_net_19248),
		.dout(new_net_2864)
	);

	bfr new_net_19249_bfr_before (
		.din(new_net_19249),
		.dout(new_net_2865)
	);

	bfr new_net_19250_bfr_before (
		.din(new_net_19250),
		.dout(new_net_2871)
	);

	spl4L new_net_3358_v_fanout (
		.a(new_net_3358),
		.b(new_net_19248),
		.c(new_net_19250),
		.d(new_net_3356),
		.e(new_net_19249)
	);

	spl4L new_net_3439_v_fanout (
		.a(new_net_3439),
		.b(new_net_1410),
		.c(new_net_1418),
		.d(new_net_1416),
		.e(new_net_1419)
	);

	spl4L new_net_3331_v_fanout (
		.a(new_net_3331),
		.b(new_net_920),
		.c(new_net_928),
		.d(new_net_922),
		.e(new_net_923)
	);

	bfr new_net_19251_bfr_before (
		.din(new_net_19251),
		.dout(new_net_3233)
	);

	bfr new_net_19252_bfr_before (
		.din(new_net_19252),
		.dout(new_net_3247)
	);

	spl4L new_net_3389_v_fanout (
		.a(new_net_3389),
		.b(new_net_19251),
		.c(new_net_3387),
		.d(new_net_3385),
		.e(new_net_19252)
	);

	spl4L new_net_3364_v_fanout (
		.a(new_net_3364),
		.b(new_net_3082),
		.c(new_net_3083),
		.d(new_net_3088),
		.e(new_net_3081)
	);

	bfr new_net_19253_bfr_before (
		.din(new_net_19253),
		.dout(new_net_403)
	);

	spl3L new_net_3342_v_fanout (
		.a(new_net_3342),
		.b(new_net_19253),
		.c(new_net_405),
		.d(new_net_3338)
	);

	spl4L new_net_3438_v_fanout (
		.a(new_net_3438),
		.b(new_net_1406),
		.c(new_net_1417),
		.d(new_net_1407),
		.e(new_net_1408)
	);

	spl3L new_net_3383_v_fanout (
		.a(new_net_3383),
		.b(new_net_3381),
		.c(new_net_3380),
		.d(new_net_3382)
	);

	spl4L new_net_3286_v_fanout (
		.a(new_net_3286),
		.b(new_net_2842),
		.c(new_net_2836),
		.d(new_net_2832),
		.e(new_net_2839)
	);

	bfr new_net_19254_bfr_before (
		.din(new_net_19254),
		.dout(new_net_152)
	);

	bfr new_net_19255_bfr_before (
		.din(new_net_19255),
		.dout(new_net_160)
	);

	bfr new_net_19256_bfr_before (
		.din(new_net_19256),
		.dout(new_net_159)
	);

	spl4L new_net_3301_v_fanout (
		.a(new_net_3301),
		.b(new_net_19254),
		.c(new_net_19256),
		.d(new_net_3298),
		.e(new_net_19255)
	);

	spl4L new_net_3311_v_fanout (
		.a(new_net_3311),
		.b(new_net_3013),
		.c(new_net_3012),
		.d(new_net_3025),
		.e(new_net_3016)
	);

	spl4L new_net_3330_v_fanout (
		.a(new_net_3330),
		.b(new_net_925),
		.c(new_net_931),
		.d(new_net_929),
		.e(new_net_926)
	);

	spl2 new_net_3319_v_fanout (
		.a(new_net_3319),
		.b(new_net_432),
		.c(new_net_433)
	);

	spl4L new_net_3295_v_fanout (
		.a(new_net_3295),
		.b(new_net_2612),
		.c(new_net_2609),
		.d(new_net_2614),
		.e(new_net_2613)
	);

	spl2 new_net_3351_v_fanout (
		.a(new_net_3351),
		.b(new_net_1441),
		.c(new_net_1454)
	);

	spl4L new_net_3368_v_fanout (
		.a(new_net_3368),
		.b(new_net_2406),
		.c(new_net_2411),
		.d(new_net_2407),
		.e(new_net_2401)
	);

	bfr new_net_19257_bfr_before (
		.din(new_net_19257),
		.dout(new_net_1452)
	);

	bfr new_net_19258_bfr_before (
		.din(new_net_19258),
		.dout(new_net_1447)
	);

	spl4L new_net_3352_v_fanout (
		.a(new_net_3352),
		.b(new_net_1450),
		.c(new_net_3350),
		.d(new_net_19258),
		.e(new_net_19257)
	);

	bfr new_net_19259_bfr_before (
		.din(new_net_19259),
		.dout(new_net_1455)
	);

	bfr new_net_19260_bfr_before (
		.din(new_net_19260),
		.dout(new_net_1456)
	);

	spl3L new_net_3354_v_fanout (
		.a(new_net_3354),
		.b(new_net_19259),
		.c(new_net_19260),
		.d(new_net_3349)
	);

	bfr new_net_19261_bfr_before (
		.din(new_net_19261),
		.dout(new_net_206)
	);

	bfr new_net_19262_bfr_before (
		.din(new_net_19262),
		.dout(new_net_208)
	);

	bfr new_net_19263_bfr_before (
		.din(new_net_19263),
		.dout(new_net_213)
	);

	spl4L new_net_3394_v_fanout (
		.a(new_net_3394),
		.b(new_net_19261),
		.c(new_net_3391),
		.d(new_net_19263),
		.e(new_net_19262)
	);

	bfr new_net_19264_bfr_before (
		.din(new_net_19264),
		.dout(new_net_1130)
	);

	spl2 new_net_3417_v_fanout (
		.a(new_net_3417),
		.b(new_net_19264),
		.c(new_net_3414)
	);

	spl4L new_net_3278_v_fanout (
		.a(new_net_3278),
		.b(new_net_381),
		.c(new_net_382),
		.d(new_net_389),
		.e(new_net_378)
	);

	bfr new_net_19265_bfr_before (
		.din(new_net_19265),
		.dout(new_net_1809)
	);

	spl4L new_net_3412_v_fanout (
		.a(new_net_3412),
		.b(new_net_3410),
		.c(new_net_3408),
		.d(new_net_3409),
		.e(new_net_19265)
	);

	spl2 new_net_3334_v_fanout (
		.a(new_net_3334),
		.b(new_net_3188),
		.c(new_net_3190)
	);

	spl4L new_net_3289_v_fanout (
		.a(new_net_3289),
		.b(new_net_2700),
		.c(new_net_2713),
		.d(new_net_2710),
		.e(new_net_2705)
	);

	spl4L new_net_3300_v_fanout (
		.a(new_net_3300),
		.b(new_net_149),
		.c(new_net_151),
		.d(new_net_147),
		.e(new_net_155)
	);

	spl2 new_net_3294_v_fanout (
		.a(new_net_3294),
		.b(new_net_2610),
		.c(new_net_2619)
	);

	spl4L new_net_3327_v_fanout (
		.a(new_net_3327),
		.b(new_net_2343),
		.c(new_net_2353),
		.d(new_net_2352),
		.e(new_net_2342)
	);

	bfr new_net_19266_bfr_before (
		.din(new_net_19266),
		.dout(new_net_3181)
	);

	bfr new_net_19267_bfr_before (
		.din(new_net_19267),
		.dout(new_net_3189)
	);

	bfr new_net_19268_bfr_before (
		.din(new_net_19268),
		.dout(new_net_3183)
	);

	spl4L new_net_3335_v_fanout (
		.a(new_net_3335),
		.b(new_net_19266),
		.c(new_net_19268),
		.d(new_net_3333),
		.e(new_net_19267)
	);

	bfr new_net_19269_bfr_before (
		.din(new_net_19269),
		.dout(new_net_2347)
	);

	bfr new_net_19270_bfr_before (
		.din(new_net_19270),
		.dout(new_net_2348)
	);

	spl3L new_net_3325_v_fanout (
		.a(new_net_3325),
		.b(new_net_19269),
		.c(new_net_3323),
		.d(new_net_19270)
	);

	bfr new_net_19271_bfr_before (
		.din(new_net_19271),
		.dout(new_net_1482)
	);

	bfr new_net_19272_bfr_before (
		.din(new_net_19272),
		.dout(new_net_1477)
	);

	spl3L new_net_3378_v_fanout (
		.a(new_net_3378),
		.b(new_net_19271),
		.c(new_net_3376),
		.d(new_net_19272)
	);

	bfr new_net_19273_bfr_before (
		.din(new_net_19273),
		.dout(new_net_3091)
	);

	spl4L new_net_3363_v_fanout (
		.a(new_net_3363),
		.b(new_net_19273),
		.c(new_net_3361),
		.d(new_net_3362),
		.e(new_net_3360)
	);

	spl2 new_net_3329_v_fanout (
		.a(new_net_3329),
		.b(new_net_917),
		.c(new_net_3328)
	);

	spl4L new_net_3296_v_fanout (
		.a(new_net_3296),
		.b(new_net_2618),
		.c(new_net_2620),
		.d(new_net_2607),
		.e(new_net_2606)
	);

	spl4L new_net_3384_v_fanout (
		.a(new_net_3384),
		.b(new_net_742),
		.c(new_net_750),
		.d(new_net_744),
		.e(new_net_743)
	);

	bfr new_net_19274_bfr_before (
		.din(new_net_19274),
		.dout(new_net_1553)
	);

	spl2 new_net_3346_v_fanout (
		.a(new_net_3346),
		.b(new_net_19274),
		.c(new_net_3344)
	);

	spl4L new_net_3283_v_fanout (
		.a(new_net_3283),
		.b(new_net_3108),
		.c(new_net_3093),
		.d(new_net_3101),
		.e(new_net_3102)
	);

	bfr new_net_19275_bfr_before (
		.din(new_net_19275),
		.dout(new_net_430)
	);

	bfr new_net_19276_bfr_before (
		.din(new_net_19276),
		.dout(new_net_427)
	);

	bfr new_net_19277_bfr_before (
		.din(new_net_19277),
		.dout(new_net_429)
	);

	spl4L new_net_3322_v_fanout (
		.a(new_net_3322),
		.b(new_net_3318),
		.c(new_net_19277),
		.d(new_net_19276),
		.e(new_net_19275)
	);

	bfr new_net_19278_bfr_before (
		.din(new_net_19278),
		.dout(new_net_526)
	);

	bfr new_net_19279_bfr_before (
		.din(new_net_19279),
		.dout(new_net_534)
	);

	spl4L new_net_3374_v_fanout (
		.a(new_net_3374),
		.b(new_net_19278),
		.c(new_net_19279),
		.d(new_net_3370),
		.e(new_net_3371)
	);

	spl4L new_net_3280_v_fanout (
		.a(new_net_3280),
		.b(new_net_3094),
		.c(new_net_3107),
		.d(new_net_3099),
		.e(new_net_3098)
	);

	bfr new_net_19280_bfr_before (
		.din(new_net_19280),
		.dout(new_net_2921)
	);

	spl2 new_net_3314_v_fanout (
		.a(new_net_3314),
		.b(new_net_3313),
		.c(new_net_19280)
	);

	spl4L new_net_3279_v_fanout (
		.a(new_net_3279),
		.b(new_net_385),
		.c(new_net_391),
		.d(new_net_377),
		.e(new_net_376)
	);

	bfr new_net_19281_bfr_before (
		.din(new_net_19281),
		.dout(new_net_380)
	);

	bfr new_net_19282_bfr_before (
		.din(new_net_19282),
		.dout(new_net_383)
	);

	bfr new_net_19283_bfr_before (
		.din(new_net_19283),
		.dout(new_net_390)
	);

	spl4L new_net_3276_v_fanout (
		.a(new_net_3276),
		.b(new_net_19281),
		.c(new_net_19283),
		.d(new_net_384),
		.e(new_net_19282)
	);

	spl4L new_net_3373_v_fanout (
		.a(new_net_3373),
		.b(new_net_528),
		.c(new_net_538),
		.d(new_net_536),
		.e(new_net_537)
	);

	spl4L new_net_3321_v_fanout (
		.a(new_net_3321),
		.b(new_net_439),
		.c(new_net_438),
		.d(new_net_428),
		.e(new_net_440)
	);

	bfr new_net_19284_bfr_before (
		.din(new_net_19284),
		.dout(new_net_3237)
	);

	bfr new_net_19285_bfr_before (
		.din(new_net_19285),
		.dout(new_net_3236)
	);

	spl3L new_net_3388_v_fanout (
		.a(new_net_3388),
		.b(new_net_19284),
		.c(new_net_3386),
		.d(new_net_19285)
	);

	bfr new_net_19286_bfr_before (
		.din(new_net_19286),
		.dout(new_net_3106)
	);

	bfr new_net_19287_bfr_before (
		.din(new_net_19287),
		.dout(new_net_3104)
	);

	bfr new_net_19288_bfr_before (
		.din(new_net_19288),
		.dout(new_net_3103)
	);

	spl4L new_net_3282_v_fanout (
		.a(new_net_3282),
		.b(new_net_3097),
		.c(new_net_19288),
		.d(new_net_19287),
		.e(new_net_19286)
	);

	bfr new_net_19289_bfr_before (
		.din(new_net_19289),
		.dout(new_net_2829)
	);

	bfr new_net_19290_bfr_before (
		.din(new_net_19290),
		.dout(new_net_2833)
	);

	bfr new_net_19291_bfr_before (
		.din(new_net_19291),
		.dout(new_net_2840)
	);

	spl4L new_net_3284_v_fanout (
		.a(new_net_3284),
		.b(new_net_19289),
		.c(new_net_2844),
		.d(new_net_19291),
		.e(new_net_19290)
	);

	spl3L new_net_3348_v_fanout (
		.a(new_net_3348),
		.b(new_net_1549),
		.c(new_net_1560),
		.d(new_net_1558)
	);

	bfr new_net_19292_bfr_before (
		.din(new_net_19292),
		.dout(new_net_2408)
	);

	spl4L new_net_3369_v_fanout (
		.a(new_net_3369),
		.b(new_net_19292),
		.c(new_net_3366),
		.d(new_net_3367),
		.e(new_net_3365)
	);

	spl4L new_net_3302_v_fanout (
		.a(new_net_3302),
		.b(new_net_158),
		.c(new_net_153),
		.d(new_net_150),
		.e(new_net_148)
	);

	spl3L new_net_3436_v_fanout (
		.a(new_net_3436),
		.b(new_net_3432),
		.c(new_net_266),
		.d(new_net_3434)
	);

	bfr new_net_19293_bfr_before (
		.din(new_net_19293),
		.dout(new_net_1250)
	);

	bfr new_net_19294_bfr_before (
		.din(new_net_19294),
		.dout(new_net_1252)
	);

	bfr new_net_19295_bfr_before (
		.din(new_net_19295),
		.dout(new_net_1253)
	);

	spl4L new_net_3306_v_fanout (
		.a(new_net_3306),
		.b(new_net_19293),
		.c(new_net_19295),
		.d(new_net_3303),
		.e(new_net_19294)
	);

	bfr new_net_19296_bfr_before (
		.din(new_net_19296),
		.dout(new_net_3019)
	);

	spl2 new_net_3309_v_fanout (
		.a(new_net_3309),
		.b(new_net_3018),
		.c(new_net_19296)
	);

	spl4L new_net_3353_v_fanout (
		.a(new_net_3353),
		.b(new_net_1446),
		.c(new_net_1451),
		.d(new_net_1445),
		.e(new_net_1443)
	);

	bfr new_net_19297_bfr_before (
		.din(new_net_19297),
		.dout(new_net_1811)
	);

	spl3L new_net_3411_v_fanout (
		.a(new_net_3411),
		.b(new_net_3407),
		.c(new_net_19297),
		.d(new_net_1804)
	);

	spl4L new_net_3341_v_fanout (
		.a(new_net_3341),
		.b(new_net_399),
		.c(new_net_407),
		.d(new_net_401),
		.e(new_net_397)
	);

	bfr new_net_19298_bfr_before (
		.din(new_net_19298),
		.dout(new_net_2866)
	);

	bfr new_net_19299_bfr_before (
		.din(new_net_19299),
		.dout(new_net_2869)
	);

	spl4L new_net_3359_v_fanout (
		.a(new_net_3359),
		.b(new_net_19298),
		.c(new_net_19299),
		.d(new_net_3357),
		.e(new_net_3355)
	);

	bfr new_net_19300_bfr_before (
		.din(new_net_19300),
		.dout(new_net_207)
	);

	spl4L new_net_3393_v_fanout (
		.a(new_net_3393),
		.b(new_net_3390),
		.c(new_net_19300),
		.d(new_net_3392),
		.e(new_net_210)
	);

	bfr new_net_19301_bfr_before (
		.din(new_net_19301),
		.dout(new_net_3179)
	);

	bfr new_net_19302_bfr_before (
		.din(new_net_19302),
		.dout(new_net_3187)
	);

	bfr new_net_19303_bfr_before (
		.din(new_net_19303),
		.dout(new_net_3186)
	);

	spl4L new_net_3336_v_fanout (
		.a(new_net_3336),
		.b(new_net_19301),
		.c(new_net_3184),
		.d(new_net_19303),
		.e(new_net_19302)
	);

	spl4L new_net_3290_v_fanout (
		.a(new_net_3290),
		.b(new_net_2707),
		.c(new_net_2708),
		.d(new_net_2709),
		.e(new_net_2711)
	);

	spl4L new_net_3440_v_fanout (
		.a(new_net_3440),
		.b(new_net_1405),
		.c(new_net_1411),
		.d(new_net_1414),
		.e(new_net_1412)
	);

	bfr new_net_19304_bfr_before (
		.din(new_net_19304),
		.dout(new_net_3105)
	);

	bfr new_net_19305_bfr_before (
		.din(new_net_19305),
		.dout(new_net_3095)
	);

	spl4L new_net_3281_v_fanout (
		.a(new_net_3281),
		.b(new_net_3096),
		.c(new_net_3100),
		.d(new_net_19305),
		.e(new_net_19304)
	);

	bfr new_net_19306_bfr_before (
		.din(new_net_19306),
		.dout(new_net_3279)
	);

	bfr new_net_19307_bfr_before (
		.din(new_net_19307),
		.dout(new_net_3278)
	);

	bfr new_net_19308_bfr_before (
		.din(new_net_19308),
		.dout(new_net_3277)
	);

	spl4L N154_v_fanout (
		.a(N154),
		.b(new_net_19306),
		.c(new_net_3276),
		.d(new_net_19308),
		.e(new_net_19307)
	);

	bfr new_net_19309_bfr_before (
		.din(new_net_19309),
		.dout(new_net_3283)
	);

	bfr new_net_19310_bfr_before (
		.din(new_net_19310),
		.dout(new_net_3280)
	);

	spl4L N290_v_fanout (
		.a(N290),
		.b(new_net_19309),
		.c(new_net_19310),
		.d(new_net_3282),
		.e(new_net_3281)
	);

	bfr new_net_19311_bfr_before (
		.din(new_net_19311),
		.dout(new_net_3287)
	);

	bfr new_net_19312_bfr_before (
		.din(new_net_19312),
		.dout(new_net_3286)
	);

	bfr new_net_19313_bfr_before (
		.din(new_net_19313),
		.dout(new_net_3285)
	);

	spl4L N1_v_fanout (
		.a(N1),
		.b(new_net_19311),
		.c(new_net_19313),
		.d(new_net_19312),
		.e(new_net_3284)
	);

	bfr new_net_19314_bfr_before (
		.din(new_net_19314),
		.dout(new_net_3290)
	);

	bfr new_net_19315_bfr_before (
		.din(new_net_19315),
		.dout(new_net_3292)
	);

	bfr new_net_19316_bfr_before (
		.din(new_net_19316),
		.dout(new_net_3289)
	);

	spl4L N222_v_fanout (
		.a(N222),
		.b(new_net_19314),
		.c(new_net_19316),
		.d(new_net_3291),
		.e(new_net_19315)
	);

	bfr new_net_19317_bfr_before (
		.din(new_net_19317),
		.dout(new_net_3295)
	);

	bfr new_net_19318_bfr_before (
		.din(new_net_19318),
		.dout(new_net_3296)
	);

	bfr new_net_19319_bfr_before (
		.din(new_net_19319),
		.dout(new_net_3294)
	);

	spl4L N443_v_fanout (
		.a(N443),
		.b(new_net_3297),
		.c(new_net_19319),
		.d(new_net_19318),
		.e(new_net_19317)
	);

	bfr new_net_19320_bfr_before (
		.din(new_net_19320),
		.dout(new_net_3300)
	);

	bfr new_net_19321_bfr_before (
		.din(new_net_19321),
		.dout(new_net_3302)
	);

	spl4L N494_v_fanout (
		.a(N494),
		.b(new_net_3301),
		.c(new_net_3299),
		.d(new_net_19321),
		.e(new_net_19320)
	);

	bfr new_net_19322_bfr_before (
		.din(new_net_19322),
		.dout(new_net_3305)
	);

	bfr new_net_19323_bfr_before (
		.din(new_net_19323),
		.dout(new_net_3307)
	);

	spl4L N358_v_fanout (
		.a(N358),
		.b(new_net_19322),
		.c(new_net_3304),
		.d(new_net_3306),
		.e(new_net_19323)
	);

	bfr new_net_19324_bfr_before (
		.din(new_net_19324),
		.dout(new_net_3311)
	);

	bfr new_net_19325_bfr_before (
		.din(new_net_19325),
		.dout(new_net_3310)
	);

	spl4L N460_v_fanout (
		.a(N460),
		.b(new_net_19324),
		.c(new_net_19325),
		.d(new_net_3312),
		.e(new_net_3309)
	);

	bfr new_net_19326_bfr_before (
		.din(new_net_19326),
		.dout(new_net_3317)
	);

	bfr new_net_19327_bfr_before (
		.din(new_net_19327),
		.dout(new_net_3315)
	);

	spl4L N273_v_fanout (
		.a(N273),
		.b(new_net_3316),
		.c(new_net_19327),
		.d(new_net_19326),
		.e(new_net_3314)
	);

	bfr new_net_19328_bfr_before (
		.din(new_net_19328),
		.dout(new_net_3321)
	);

	bfr new_net_19329_bfr_before (
		.din(new_net_19329),
		.dout(new_net_3319)
	);

	spl4L N477_v_fanout (
		.a(N477),
		.b(new_net_19328),
		.c(new_net_3320),
		.d(new_net_19329),
		.e(new_net_3322)
	);

	bfr new_net_19330_bfr_before (
		.din(new_net_19330),
		.dout(new_net_3327)
	);

	spl3L N120_v_fanout (
		.a(N120),
		.b(new_net_19330),
		.c(new_net_3325),
		.d(new_net_3326)
	);

	bfr new_net_19331_bfr_before (
		.din(new_net_19331),
		.dout(new_net_3331)
	);

	bfr new_net_19332_bfr_before (
		.din(new_net_19332),
		.dout(new_net_3330)
	);

	bfr new_net_19333_bfr_before (
		.din(new_net_19333),
		.dout(new_net_3332)
	);

	spl4L N528_v_fanout (
		.a(N528),
		.b(new_net_19331),
		.c(new_net_19333),
		.d(new_net_3329),
		.e(new_net_19332)
	);

	bfr new_net_19334_bfr_before (
		.din(new_net_19334),
		.dout(new_net_3337)
	);

	bfr new_net_19335_bfr_before (
		.din(new_net_19335),
		.dout(new_net_3334)
	);

	spl4L N341_v_fanout (
		.a(N341),
		.b(new_net_19334),
		.c(new_net_19335),
		.d(new_net_3335),
		.e(new_net_3336)
	);

	bfr new_net_19336_bfr_before (
		.din(new_net_19336),
		.dout(new_net_3341)
	);

	bfr new_net_19337_bfr_before (
		.din(new_net_19337),
		.dout(new_net_3339)
	);

	bfr new_net_19338_bfr_before (
		.din(new_net_19338),
		.dout(new_net_3340)
	);

	spl4L N324_v_fanout (
		.a(N324),
		.b(new_net_3342),
		.c(new_net_19338),
		.d(new_net_19337),
		.e(new_net_19336)
	);

	bfr new_net_19339_bfr_before (
		.din(new_net_19339),
		.dout(new_net_3348)
	);

	spl3L N205_v_fanout (
		.a(N205),
		.b(new_net_19339),
		.c(new_net_3346),
		.d(new_net_3347)
	);

	bfr new_net_19340_bfr_before (
		.din(new_net_19340),
		.dout(new_net_3351)
	);

	bfr new_net_19341_bfr_before (
		.din(new_net_19341),
		.dout(new_net_3353)
	);

	spl4L N375_v_fanout (
		.a(N375),
		.b(new_net_3354),
		.c(new_net_19341),
		.d(new_net_19340),
		.e(new_net_3352)
	);

	spl2 N256_v_fanout (
		.a(N256),
		.b(new_net_3359),
		.c(new_net_3358)
	);

	bfr new_net_19342_bfr_before (
		.din(new_net_19342),
		.dout(new_net_3364)
	);

	spl2 N103_v_fanout (
		.a(N103),
		.b(new_net_19342),
		.c(new_net_3363)
	);

	bfr new_net_19343_bfr_before (
		.din(new_net_19343),
		.dout(new_net_3368)
	);

	spl2 N137_v_fanout (
		.a(N137),
		.b(new_net_3369),
		.c(new_net_19343)
	);

	bfr new_net_19344_bfr_before (
		.din(new_net_19344),
		.dout(new_net_3373)
	);

	spl3L N511_v_fanout (
		.a(N511),
		.b(new_net_3372),
		.c(new_net_19344),
		.d(new_net_3374)
	);

	spl2 N86_v_fanout (
		.a(N86),
		.b(new_net_3378),
		.c(new_net_3379)
	);

	bfr new_net_19345_bfr_before (
		.din(new_net_19345),
		.dout(new_net_3384)
	);

	spl2 N52_v_fanout (
		.a(N52),
		.b(new_net_3383),
		.c(new_net_19345)
	);

	spl2 N35_v_fanout (
		.a(N35),
		.b(new_net_3388),
		.c(new_net_3389)
	);

	spl2 N409_v_fanout (
		.a(N409),
		.b(new_net_3393),
		.c(new_net_3394)
	);

	spl2 N171_v_fanout (
		.a(N171),
		.b(new_net_3400),
		.c(new_net_3399)
	);

	spl2 N18_v_fanout (
		.a(N18),
		.b(new_net_3405),
		.c(new_net_3406)
	);

	spl2 N392_v_fanout (
		.a(N392),
		.b(new_net_3411),
		.c(new_net_3412)
	);

	spl2 N188_v_fanout (
		.a(N188),
		.b(new_net_3418),
		.c(new_net_3417)
	);

	spl2 N307_v_fanout (
		.a(N307),
		.b(new_net_3423),
		.c(new_net_3424)
	);

	spl2 N239_v_fanout (
		.a(N239),
		.b(new_net_3430),
		.c(new_net_3429)
	);

	spl2 N426_v_fanout (
		.a(N426),
		.b(new_net_3436),
		.c(new_net_3435)
	);

	spl4L N69_v_fanout (
		.a(N69),
		.b(new_net_3440),
		.c(new_net_3438),
		.d(new_net_3437),
		.e(new_net_3439)
	);

	bfr new_net_3470_bfr_after (
		.din(_0448_),
		.dout(new_net_3470)
	);

	bfr new_net_3580_bfr_after (
		.din(_1394_),
		.dout(new_net_3580)
	);

	bfr new_net_3724_bfr_after (
		.din(_0174_),
		.dout(new_net_3724)
	);

	bfr new_net_3808_bfr_after (
		.din(_0554_),
		.dout(new_net_3808)
	);

	bfr new_net_3874_bfr_after (
		.din(_0825_),
		.dout(new_net_3874)
	);

	bfr new_net_3469_bfr_after (
		.din(_0416_),
		.dout(new_net_3469)
	);

	bfr new_net_3480_bfr_after (
		.din(_0904_),
		.dout(new_net_3480)
	);

	bfr new_net_3534_bfr_after (
		.din(_1200_),
		.dout(new_net_3534)
	);

	bfr new_net_3656_bfr_after (
		.din(_1726_),
		.dout(new_net_3656)
	);

	bfr new_net_3756_bfr_after (
		.din(_0310_),
		.dout(new_net_3756)
	);

	bfr new_net_3799_bfr_after (
		.din(_0502_),
		.dout(new_net_3799)
	);

	bfr new_net_3483_bfr_after (
		.din(_1000_),
		.dout(new_net_3483)
	);

	bfr new_net_3765_bfr_after (
		.din(_0366_),
		.dout(new_net_3765)
	);

	bfr new_net_3866_bfr_after (
		.din(_0799_),
		.dout(new_net_3866)
	);

	bfr new_net_19346_bfr_after (
		.din(new_net_3954),
		.dout(new_net_19346)
	);

	bfr new_net_19347_bfr_after (
		.din(new_net_19346),
		.dout(new_net_19347)
	);

	bfr new_net_19348_bfr_after (
		.din(new_net_19347),
		.dout(new_net_19348)
	);

	bfr new_net_19349_bfr_after (
		.din(new_net_19348),
		.dout(new_net_19349)
	);

	bfr new_net_19350_bfr_after (
		.din(new_net_19349),
		.dout(new_net_19350)
	);

	bfr new_net_19351_bfr_after (
		.din(new_net_19350),
		.dout(new_net_19351)
	);

	bfr new_net_19352_bfr_after (
		.din(new_net_19351),
		.dout(new_net_19352)
	);

	bfr new_net_19353_bfr_after (
		.din(new_net_19352),
		.dout(new_net_19353)
	);

	bfr new_net_19354_bfr_after (
		.din(new_net_19353),
		.dout(new_net_19354)
	);

	bfr new_net_19355_bfr_after (
		.din(new_net_19354),
		.dout(new_net_19355)
	);

	bfr new_net_19356_bfr_after (
		.din(new_net_19355),
		.dout(new_net_19356)
	);

	bfr new_net_19357_bfr_after (
		.din(new_net_19356),
		.dout(new_net_19357)
	);

	bfr new_net_19358_bfr_after (
		.din(new_net_19357),
		.dout(new_net_19358)
	);

	bfr new_net_19359_bfr_after (
		.din(new_net_19358),
		.dout(new_net_19359)
	);

	bfr new_net_19360_bfr_after (
		.din(new_net_19359),
		.dout(new_net_19360)
	);

	bfr new_net_19361_bfr_after (
		.din(new_net_19360),
		.dout(new_net_19361)
	);

	bfr new_net_19362_bfr_after (
		.din(new_net_19361),
		.dout(new_net_19362)
	);

	bfr new_net_19363_bfr_after (
		.din(new_net_19362),
		.dout(new_net_19363)
	);

	bfr new_net_19364_bfr_after (
		.din(new_net_19363),
		.dout(new_net_19364)
	);

	bfr new_net_19365_bfr_after (
		.din(new_net_19364),
		.dout(new_net_19365)
	);

	bfr new_net_19366_bfr_after (
		.din(new_net_19365),
		.dout(new_net_19366)
	);

	bfr new_net_19367_bfr_after (
		.din(new_net_19366),
		.dout(new_net_19367)
	);

	bfr new_net_19368_bfr_after (
		.din(new_net_19367),
		.dout(new_net_19368)
	);

	bfr new_net_19369_bfr_after (
		.din(new_net_19368),
		.dout(new_net_19369)
	);

	bfr new_net_19370_bfr_after (
		.din(new_net_19369),
		.dout(new_net_19370)
	);

	bfr new_net_19371_bfr_after (
		.din(new_net_19370),
		.dout(new_net_19371)
	);

	bfr new_net_19372_bfr_after (
		.din(new_net_19371),
		.dout(new_net_19372)
	);

	bfr new_net_19373_bfr_after (
		.din(new_net_19372),
		.dout(new_net_19373)
	);

	bfr new_net_19374_bfr_after (
		.din(new_net_19373),
		.dout(new_net_19374)
	);

	bfr new_net_19375_bfr_after (
		.din(new_net_19374),
		.dout(new_net_19375)
	);

	bfr new_net_19376_bfr_after (
		.din(new_net_19375),
		.dout(new_net_19376)
	);

	bfr new_net_19377_bfr_after (
		.din(new_net_19376),
		.dout(new_net_19377)
	);

	bfr new_net_19378_bfr_after (
		.din(new_net_19377),
		.dout(new_net_19378)
	);

	bfr new_net_19379_bfr_after (
		.din(new_net_19378),
		.dout(new_net_19379)
	);

	bfr new_net_19380_bfr_after (
		.din(new_net_19379),
		.dout(new_net_19380)
	);

	bfr new_net_19381_bfr_after (
		.din(new_net_19380),
		.dout(new_net_19381)
	);

	bfr new_net_19382_bfr_after (
		.din(new_net_19381),
		.dout(new_net_19382)
	);

	bfr new_net_19383_bfr_after (
		.din(new_net_19382),
		.dout(new_net_19383)
	);

	bfr new_net_19384_bfr_after (
		.din(new_net_19383),
		.dout(new_net_19384)
	);

	bfr new_net_19385_bfr_after (
		.din(new_net_19384),
		.dout(new_net_19385)
	);

	bfr new_net_19386_bfr_after (
		.din(new_net_19385),
		.dout(new_net_19386)
	);

	bfr new_net_19387_bfr_after (
		.din(new_net_19386),
		.dout(new_net_19387)
	);

	bfr new_net_19388_bfr_after (
		.din(new_net_19387),
		.dout(new_net_19388)
	);

	bfr new_net_19389_bfr_after (
		.din(new_net_19388),
		.dout(new_net_19389)
	);

	bfr new_net_19390_bfr_after (
		.din(new_net_19389),
		.dout(new_net_19390)
	);

	bfr new_net_19391_bfr_after (
		.din(new_net_19390),
		.dout(new_net_19391)
	);

	bfr new_net_19392_bfr_after (
		.din(new_net_19391),
		.dout(new_net_19392)
	);

	bfr new_net_19393_bfr_after (
		.din(new_net_19392),
		.dout(new_net_19393)
	);

	bfr new_net_19394_bfr_after (
		.din(new_net_19393),
		.dout(new_net_19394)
	);

	bfr new_net_19395_bfr_after (
		.din(new_net_19394),
		.dout(new_net_19395)
	);

	bfr new_net_19396_bfr_after (
		.din(new_net_19395),
		.dout(new_net_19396)
	);

	bfr new_net_19397_bfr_after (
		.din(new_net_19396),
		.dout(new_net_19397)
	);

	bfr new_net_19398_bfr_after (
		.din(new_net_19397),
		.dout(new_net_19398)
	);

	bfr new_net_19399_bfr_after (
		.din(new_net_19398),
		.dout(new_net_19399)
	);

	bfr new_net_19400_bfr_after (
		.din(new_net_19399),
		.dout(new_net_19400)
	);

	bfr new_net_19401_bfr_after (
		.din(new_net_19400),
		.dout(new_net_19401)
	);

	bfr new_net_19402_bfr_after (
		.din(new_net_19401),
		.dout(new_net_19402)
	);

	bfr new_net_19403_bfr_after (
		.din(new_net_19402),
		.dout(new_net_19403)
	);

	bfr new_net_19404_bfr_after (
		.din(new_net_19403),
		.dout(new_net_19404)
	);

	bfr new_net_19405_bfr_after (
		.din(new_net_19404),
		.dout(new_net_19405)
	);

	bfr new_net_19406_bfr_after (
		.din(new_net_19405),
		.dout(new_net_19406)
	);

	bfr new_net_19407_bfr_after (
		.din(new_net_19406),
		.dout(new_net_19407)
	);

	bfr new_net_19408_bfr_after (
		.din(new_net_19407),
		.dout(new_net_19408)
	);

	bfr new_net_19409_bfr_after (
		.din(new_net_19408),
		.dout(new_net_19409)
	);

	bfr new_net_19410_bfr_after (
		.din(new_net_19409),
		.dout(new_net_19410)
	);

	bfr new_net_19411_bfr_after (
		.din(new_net_19410),
		.dout(new_net_19411)
	);

	bfr new_net_19412_bfr_after (
		.din(new_net_19411),
		.dout(new_net_19412)
	);

	bfr new_net_19413_bfr_after (
		.din(new_net_19412),
		.dout(new_net_19413)
	);

	bfr new_net_19414_bfr_after (
		.din(new_net_19413),
		.dout(new_net_19414)
	);

	bfr new_net_19415_bfr_after (
		.din(new_net_19414),
		.dout(new_net_19415)
	);

	bfr new_net_19416_bfr_after (
		.din(new_net_19415),
		.dout(new_net_19416)
	);

	bfr new_net_19417_bfr_after (
		.din(new_net_19416),
		.dout(new_net_19417)
	);

	bfr new_net_19418_bfr_after (
		.din(new_net_19417),
		.dout(new_net_19418)
	);

	bfr new_net_19419_bfr_after (
		.din(new_net_19418),
		.dout(new_net_19419)
	);

	bfr new_net_19420_bfr_after (
		.din(new_net_19419),
		.dout(new_net_19420)
	);

	bfr new_net_19421_bfr_after (
		.din(new_net_19420),
		.dout(new_net_19421)
	);

	bfr new_net_19422_bfr_after (
		.din(new_net_19421),
		.dout(new_net_19422)
	);

	bfr new_net_19423_bfr_after (
		.din(new_net_19422),
		.dout(new_net_19423)
	);

	bfr new_net_19424_bfr_after (
		.din(new_net_19423),
		.dout(new_net_19424)
	);

	bfr new_net_19425_bfr_after (
		.din(new_net_19424),
		.dout(new_net_19425)
	);

	bfr new_net_19426_bfr_after (
		.din(new_net_19425),
		.dout(new_net_19426)
	);

	bfr new_net_19427_bfr_after (
		.din(new_net_19426),
		.dout(new_net_19427)
	);

	bfr new_net_19428_bfr_after (
		.din(new_net_19427),
		.dout(new_net_19428)
	);

	bfr new_net_19429_bfr_after (
		.din(new_net_19428),
		.dout(new_net_19429)
	);

	bfr new_net_19430_bfr_after (
		.din(new_net_19429),
		.dout(new_net_19430)
	);

	bfr new_net_19431_bfr_after (
		.din(new_net_19430),
		.dout(new_net_19431)
	);

	bfr new_net_19432_bfr_after (
		.din(new_net_19431),
		.dout(new_net_19432)
	);

	bfr new_net_19433_bfr_after (
		.din(new_net_19432),
		.dout(new_net_19433)
	);

	bfr new_net_19434_bfr_after (
		.din(new_net_19433),
		.dout(new_net_19434)
	);

	bfr new_net_19435_bfr_after (
		.din(new_net_19434),
		.dout(new_net_19435)
	);

	bfr new_net_19436_bfr_after (
		.din(new_net_19435),
		.dout(new_net_19436)
	);

	bfr new_net_19437_bfr_after (
		.din(new_net_19436),
		.dout(new_net_19437)
	);

	bfr new_net_19438_bfr_after (
		.din(new_net_19437),
		.dout(new_net_19438)
	);

	bfr new_net_19439_bfr_after (
		.din(new_net_19438),
		.dout(new_net_19439)
	);

	bfr new_net_19440_bfr_after (
		.din(new_net_19439),
		.dout(new_net_19440)
	);

	bfr new_net_19441_bfr_after (
		.din(new_net_19440),
		.dout(new_net_19441)
	);

	bfr new_net_19442_bfr_after (
		.din(new_net_19441),
		.dout(new_net_19442)
	);

	bfr new_net_19443_bfr_after (
		.din(new_net_19442),
		.dout(new_net_19443)
	);

	bfr new_net_19444_bfr_after (
		.din(new_net_19443),
		.dout(new_net_19444)
	);

	bfr new_net_19445_bfr_after (
		.din(new_net_19444),
		.dout(new_net_19445)
	);

	bfr new_net_19446_bfr_after (
		.din(new_net_19445),
		.dout(new_net_19446)
	);

	bfr new_net_19447_bfr_after (
		.din(new_net_19446),
		.dout(new_net_19447)
	);

	bfr new_net_19448_bfr_after (
		.din(new_net_19447),
		.dout(new_net_19448)
	);

	bfr new_net_19449_bfr_after (
		.din(new_net_19448),
		.dout(new_net_19449)
	);

	bfr new_net_19450_bfr_after (
		.din(new_net_19449),
		.dout(new_net_19450)
	);

	bfr new_net_19451_bfr_after (
		.din(new_net_19450),
		.dout(new_net_19451)
	);

	bfr new_net_19452_bfr_after (
		.din(new_net_19451),
		.dout(new_net_19452)
	);

	bfr new_net_19453_bfr_after (
		.din(new_net_19452),
		.dout(new_net_19453)
	);

	bfr new_net_19454_bfr_after (
		.din(new_net_19453),
		.dout(new_net_19454)
	);

	bfr new_net_19455_bfr_after (
		.din(new_net_19454),
		.dout(new_net_19455)
	);

	bfr new_net_19456_bfr_after (
		.din(new_net_19455),
		.dout(new_net_19456)
	);

	bfr new_net_19457_bfr_after (
		.din(new_net_19456),
		.dout(new_net_19457)
	);

	bfr new_net_19458_bfr_after (
		.din(new_net_19457),
		.dout(new_net_19458)
	);

	bfr new_net_19459_bfr_after (
		.din(new_net_19458),
		.dout(new_net_19459)
	);

	bfr new_net_19460_bfr_after (
		.din(new_net_19459),
		.dout(new_net_19460)
	);

	bfr new_net_19461_bfr_after (
		.din(new_net_19460),
		.dout(new_net_19461)
	);

	bfr new_net_19462_bfr_after (
		.din(new_net_19461),
		.dout(new_net_19462)
	);

	bfr new_net_19463_bfr_after (
		.din(new_net_19462),
		.dout(new_net_19463)
	);

	bfr new_net_19464_bfr_after (
		.din(new_net_19463),
		.dout(new_net_19464)
	);

	bfr new_net_19465_bfr_after (
		.din(new_net_19464),
		.dout(new_net_19465)
	);

	bfr new_net_19466_bfr_after (
		.din(new_net_19465),
		.dout(new_net_19466)
	);

	bfr new_net_19467_bfr_after (
		.din(new_net_19466),
		.dout(new_net_19467)
	);

	bfr new_net_19468_bfr_after (
		.din(new_net_19467),
		.dout(new_net_19468)
	);

	bfr new_net_19469_bfr_after (
		.din(new_net_19468),
		.dout(new_net_19469)
	);

	bfr new_net_19470_bfr_after (
		.din(new_net_19469),
		.dout(new_net_19470)
	);

	bfr new_net_19471_bfr_after (
		.din(new_net_19470),
		.dout(new_net_19471)
	);

	bfr new_net_19472_bfr_after (
		.din(new_net_19471),
		.dout(new_net_19472)
	);

	bfr new_net_19473_bfr_after (
		.din(new_net_19472),
		.dout(new_net_19473)
	);

	bfr new_net_19474_bfr_after (
		.din(new_net_19473),
		.dout(new_net_19474)
	);

	bfr new_net_19475_bfr_after (
		.din(new_net_19474),
		.dout(new_net_19475)
	);

	bfr new_net_19476_bfr_after (
		.din(new_net_19475),
		.dout(new_net_19476)
	);

	bfr new_net_19477_bfr_after (
		.din(new_net_19476),
		.dout(new_net_19477)
	);

	bfr new_net_19478_bfr_after (
		.din(new_net_19477),
		.dout(new_net_19478)
	);

	bfr new_net_19479_bfr_after (
		.din(new_net_19478),
		.dout(new_net_19479)
	);

	bfr new_net_19480_bfr_after (
		.din(new_net_19479),
		.dout(new_net_19480)
	);

	bfr new_net_19481_bfr_after (
		.din(new_net_19480),
		.dout(new_net_19481)
	);

	bfr new_net_19482_bfr_after (
		.din(new_net_19481),
		.dout(new_net_19482)
	);

	bfr new_net_19483_bfr_after (
		.din(new_net_19482),
		.dout(new_net_19483)
	);

	bfr new_net_19484_bfr_after (
		.din(new_net_19483),
		.dout(new_net_19484)
	);

	bfr N2877_bfr_after (
		.din(new_net_19484),
		.dout(N2877)
	);

	bfr new_net_3458_bfr_after (
		.din(_1708_),
		.dout(new_net_3458)
	);

	bfr new_net_3497_bfr_after (
		.din(_1068_),
		.dout(new_net_3497)
	);

	bfr new_net_3784_bfr_after (
		.din(_0429_),
		.dout(new_net_3784)
	);

	bfr new_net_3830_bfr_after (
		.din(_0647_),
		.dout(new_net_3830)
	);

	bfr new_net_3868_bfr_after (
		.din(_0805_),
		.dout(new_net_3868)
	);

	bfr new_net_19485_bfr_after (
		.din(new_net_3942),
		.dout(new_net_19485)
	);

	bfr new_net_19486_bfr_after (
		.din(new_net_19485),
		.dout(new_net_19486)
	);

	bfr new_net_19487_bfr_after (
		.din(new_net_19486),
		.dout(new_net_19487)
	);

	bfr new_net_19488_bfr_after (
		.din(new_net_19487),
		.dout(new_net_19488)
	);

	bfr new_net_19489_bfr_after (
		.din(new_net_19488),
		.dout(new_net_19489)
	);

	bfr new_net_19490_bfr_after (
		.din(new_net_19489),
		.dout(new_net_19490)
	);

	bfr new_net_19491_bfr_after (
		.din(new_net_19490),
		.dout(new_net_19491)
	);

	bfr new_net_19492_bfr_after (
		.din(new_net_19491),
		.dout(new_net_19492)
	);

	bfr new_net_19493_bfr_after (
		.din(new_net_19492),
		.dout(new_net_19493)
	);

	bfr new_net_19494_bfr_after (
		.din(new_net_19493),
		.dout(new_net_19494)
	);

	bfr new_net_19495_bfr_after (
		.din(new_net_19494),
		.dout(new_net_19495)
	);

	bfr new_net_19496_bfr_after (
		.din(new_net_19495),
		.dout(new_net_19496)
	);

	bfr new_net_19497_bfr_after (
		.din(new_net_19496),
		.dout(new_net_19497)
	);

	bfr new_net_19498_bfr_after (
		.din(new_net_19497),
		.dout(new_net_19498)
	);

	bfr new_net_19499_bfr_after (
		.din(new_net_19498),
		.dout(new_net_19499)
	);

	bfr new_net_19500_bfr_after (
		.din(new_net_19499),
		.dout(new_net_19500)
	);

	bfr new_net_19501_bfr_after (
		.din(new_net_19500),
		.dout(new_net_19501)
	);

	bfr new_net_19502_bfr_after (
		.din(new_net_19501),
		.dout(new_net_19502)
	);

	bfr new_net_19503_bfr_after (
		.din(new_net_19502),
		.dout(new_net_19503)
	);

	bfr new_net_19504_bfr_after (
		.din(new_net_19503),
		.dout(new_net_19504)
	);

	bfr new_net_19505_bfr_after (
		.din(new_net_19504),
		.dout(new_net_19505)
	);

	bfr new_net_19506_bfr_after (
		.din(new_net_19505),
		.dout(new_net_19506)
	);

	bfr new_net_19507_bfr_after (
		.din(new_net_19506),
		.dout(new_net_19507)
	);

	bfr new_net_19508_bfr_after (
		.din(new_net_19507),
		.dout(new_net_19508)
	);

	bfr new_net_19509_bfr_after (
		.din(new_net_19508),
		.dout(new_net_19509)
	);

	bfr new_net_19510_bfr_after (
		.din(new_net_19509),
		.dout(new_net_19510)
	);

	bfr new_net_19511_bfr_after (
		.din(new_net_19510),
		.dout(new_net_19511)
	);

	bfr new_net_19512_bfr_after (
		.din(new_net_19511),
		.dout(new_net_19512)
	);

	bfr new_net_19513_bfr_after (
		.din(new_net_19512),
		.dout(new_net_19513)
	);

	bfr new_net_19514_bfr_after (
		.din(new_net_19513),
		.dout(new_net_19514)
	);

	bfr new_net_19515_bfr_after (
		.din(new_net_19514),
		.dout(new_net_19515)
	);

	bfr new_net_19516_bfr_after (
		.din(new_net_19515),
		.dout(new_net_19516)
	);

	bfr new_net_19517_bfr_after (
		.din(new_net_19516),
		.dout(new_net_19517)
	);

	bfr new_net_19518_bfr_after (
		.din(new_net_19517),
		.dout(new_net_19518)
	);

	bfr new_net_19519_bfr_after (
		.din(new_net_19518),
		.dout(new_net_19519)
	);

	bfr new_net_19520_bfr_after (
		.din(new_net_19519),
		.dout(new_net_19520)
	);

	bfr new_net_19521_bfr_after (
		.din(new_net_19520),
		.dout(new_net_19521)
	);

	bfr new_net_19522_bfr_after (
		.din(new_net_19521),
		.dout(new_net_19522)
	);

	bfr new_net_19523_bfr_after (
		.din(new_net_19522),
		.dout(new_net_19523)
	);

	bfr new_net_19524_bfr_after (
		.din(new_net_19523),
		.dout(new_net_19524)
	);

	bfr new_net_19525_bfr_after (
		.din(new_net_19524),
		.dout(new_net_19525)
	);

	bfr new_net_19526_bfr_after (
		.din(new_net_19525),
		.dout(new_net_19526)
	);

	bfr new_net_19527_bfr_after (
		.din(new_net_19526),
		.dout(new_net_19527)
	);

	bfr new_net_19528_bfr_after (
		.din(new_net_19527),
		.dout(new_net_19528)
	);

	bfr new_net_19529_bfr_after (
		.din(new_net_19528),
		.dout(new_net_19529)
	);

	bfr new_net_19530_bfr_after (
		.din(new_net_19529),
		.dout(new_net_19530)
	);

	bfr new_net_19531_bfr_after (
		.din(new_net_19530),
		.dout(new_net_19531)
	);

	bfr new_net_19532_bfr_after (
		.din(new_net_19531),
		.dout(new_net_19532)
	);

	bfr new_net_19533_bfr_after (
		.din(new_net_19532),
		.dout(new_net_19533)
	);

	bfr new_net_19534_bfr_after (
		.din(new_net_19533),
		.dout(new_net_19534)
	);

	bfr new_net_19535_bfr_after (
		.din(new_net_19534),
		.dout(new_net_19535)
	);

	bfr new_net_19536_bfr_after (
		.din(new_net_19535),
		.dout(new_net_19536)
	);

	bfr new_net_19537_bfr_after (
		.din(new_net_19536),
		.dout(new_net_19537)
	);

	bfr new_net_19538_bfr_after (
		.din(new_net_19537),
		.dout(new_net_19538)
	);

	bfr new_net_19539_bfr_after (
		.din(new_net_19538),
		.dout(new_net_19539)
	);

	bfr new_net_19540_bfr_after (
		.din(new_net_19539),
		.dout(new_net_19540)
	);

	bfr new_net_19541_bfr_after (
		.din(new_net_19540),
		.dout(new_net_19541)
	);

	bfr new_net_19542_bfr_after (
		.din(new_net_19541),
		.dout(new_net_19542)
	);

	bfr new_net_19543_bfr_after (
		.din(new_net_19542),
		.dout(new_net_19543)
	);

	bfr new_net_19544_bfr_after (
		.din(new_net_19543),
		.dout(new_net_19544)
	);

	bfr new_net_19545_bfr_after (
		.din(new_net_19544),
		.dout(new_net_19545)
	);

	bfr new_net_19546_bfr_after (
		.din(new_net_19545),
		.dout(new_net_19546)
	);

	bfr new_net_19547_bfr_after (
		.din(new_net_19546),
		.dout(new_net_19547)
	);

	bfr new_net_19548_bfr_after (
		.din(new_net_19547),
		.dout(new_net_19548)
	);

	bfr new_net_19549_bfr_after (
		.din(new_net_19548),
		.dout(new_net_19549)
	);

	bfr new_net_19550_bfr_after (
		.din(new_net_19549),
		.dout(new_net_19550)
	);

	bfr new_net_19551_bfr_after (
		.din(new_net_19550),
		.dout(new_net_19551)
	);

	bfr N5971_bfr_after (
		.din(new_net_19551),
		.dout(N5971)
	);

	bfr new_net_3596_bfr_after (
		.din(_1442_),
		.dout(new_net_3596)
	);

	bfr new_net_3636_bfr_after (
		.din(_1627_),
		.dout(new_net_3636)
	);

	bfr new_net_3673_bfr_after (
		.din(_1782_),
		.dout(new_net_3673)
	);

	bfr new_net_3771_bfr_after (
		.din(_0386_),
		.dout(new_net_3771)
	);

	bfr new_net_3821_bfr_after (
		.din(_0597_),
		.dout(new_net_3821)
	);

	bfr new_net_3825_bfr_after (
		.din(_0610_),
		.dout(new_net_3825)
	);

	bfr new_net_3811_bfr_after (
		.din(_0564_),
		.dout(new_net_3811)
	);

	bfr new_net_3847_bfr_after (
		.din(_0721_),
		.dout(new_net_3847)
	);

	bfr new_net_3875_bfr_after (
		.din(_0842_),
		.dout(new_net_3875)
	);

	bfr new_net_3455_bfr_after (
		.din(_1524_),
		.dout(new_net_3455)
	);

	bfr new_net_3460_bfr_after (
		.din(_1774_),
		.dout(new_net_3460)
	);

	bfr new_net_3516_bfr_after (
		.din(_1158_),
		.dout(new_net_3516)
	);

	bfr new_net_3595_bfr_after (
		.din(_1439_),
		.dout(new_net_3595)
	);

	bfr new_net_3679_bfr_after (
		.din(_1802_),
		.dout(new_net_3679)
	);

	bfr new_net_3720_bfr_after (
		.din(_0161_),
		.dout(new_net_3720)
	);

	bfr new_net_3774_bfr_after (
		.din(_0396_),
		.dout(new_net_3774)
	);

	bfr new_net_19552_bfr_after (
		.din(new_net_3962),
		.dout(new_net_19552)
	);

	bfr new_net_19553_bfr_after (
		.din(new_net_19552),
		.dout(new_net_19553)
	);

	bfr new_net_19554_bfr_after (
		.din(new_net_19553),
		.dout(new_net_19554)
	);

	bfr new_net_19555_bfr_after (
		.din(new_net_19554),
		.dout(new_net_19555)
	);

	bfr new_net_19556_bfr_after (
		.din(new_net_19555),
		.dout(new_net_19556)
	);

	bfr new_net_19557_bfr_after (
		.din(new_net_19556),
		.dout(new_net_19557)
	);

	bfr new_net_19558_bfr_after (
		.din(new_net_19557),
		.dout(new_net_19558)
	);

	bfr new_net_19559_bfr_after (
		.din(new_net_19558),
		.dout(new_net_19559)
	);

	bfr new_net_19560_bfr_after (
		.din(new_net_19559),
		.dout(new_net_19560)
	);

	bfr new_net_19561_bfr_after (
		.din(new_net_19560),
		.dout(new_net_19561)
	);

	bfr new_net_19562_bfr_after (
		.din(new_net_19561),
		.dout(new_net_19562)
	);

	bfr new_net_19563_bfr_after (
		.din(new_net_19562),
		.dout(new_net_19563)
	);

	bfr new_net_19564_bfr_after (
		.din(new_net_19563),
		.dout(new_net_19564)
	);

	bfr new_net_19565_bfr_after (
		.din(new_net_19564),
		.dout(new_net_19565)
	);

	bfr new_net_19566_bfr_after (
		.din(new_net_19565),
		.dout(new_net_19566)
	);

	bfr new_net_19567_bfr_after (
		.din(new_net_19566),
		.dout(new_net_19567)
	);

	bfr new_net_19568_bfr_after (
		.din(new_net_19567),
		.dout(new_net_19568)
	);

	bfr new_net_19569_bfr_after (
		.din(new_net_19568),
		.dout(new_net_19569)
	);

	bfr new_net_19570_bfr_after (
		.din(new_net_19569),
		.dout(new_net_19570)
	);

	bfr new_net_19571_bfr_after (
		.din(new_net_19570),
		.dout(new_net_19571)
	);

	bfr new_net_19572_bfr_after (
		.din(new_net_19571),
		.dout(new_net_19572)
	);

	bfr new_net_19573_bfr_after (
		.din(new_net_19572),
		.dout(new_net_19573)
	);

	bfr new_net_19574_bfr_after (
		.din(new_net_19573),
		.dout(new_net_19574)
	);

	bfr new_net_19575_bfr_after (
		.din(new_net_19574),
		.dout(new_net_19575)
	);

	bfr new_net_19576_bfr_after (
		.din(new_net_19575),
		.dout(new_net_19576)
	);

	bfr new_net_19577_bfr_after (
		.din(new_net_19576),
		.dout(new_net_19577)
	);

	bfr new_net_19578_bfr_after (
		.din(new_net_19577),
		.dout(new_net_19578)
	);

	bfr new_net_19579_bfr_after (
		.din(new_net_19578),
		.dout(new_net_19579)
	);

	bfr new_net_19580_bfr_after (
		.din(new_net_19579),
		.dout(new_net_19580)
	);

	bfr new_net_19581_bfr_after (
		.din(new_net_19580),
		.dout(new_net_19581)
	);

	bfr new_net_19582_bfr_after (
		.din(new_net_19581),
		.dout(new_net_19582)
	);

	bfr new_net_19583_bfr_after (
		.din(new_net_19582),
		.dout(new_net_19583)
	);

	bfr new_net_19584_bfr_after (
		.din(new_net_19583),
		.dout(new_net_19584)
	);

	bfr new_net_19585_bfr_after (
		.din(new_net_19584),
		.dout(new_net_19585)
	);

	bfr new_net_19586_bfr_after (
		.din(new_net_19585),
		.dout(new_net_19586)
	);

	bfr new_net_19587_bfr_after (
		.din(new_net_19586),
		.dout(new_net_19587)
	);

	bfr new_net_19588_bfr_after (
		.din(new_net_19587),
		.dout(new_net_19588)
	);

	bfr new_net_19589_bfr_after (
		.din(new_net_19588),
		.dout(new_net_19589)
	);

	bfr new_net_19590_bfr_after (
		.din(new_net_19589),
		.dout(new_net_19590)
	);

	bfr new_net_19591_bfr_after (
		.din(new_net_19590),
		.dout(new_net_19591)
	);

	bfr new_net_19592_bfr_after (
		.din(new_net_19591),
		.dout(new_net_19592)
	);

	bfr new_net_19593_bfr_after (
		.din(new_net_19592),
		.dout(new_net_19593)
	);

	bfr new_net_19594_bfr_after (
		.din(new_net_19593),
		.dout(new_net_19594)
	);

	bfr new_net_19595_bfr_after (
		.din(new_net_19594),
		.dout(new_net_19595)
	);

	bfr new_net_19596_bfr_after (
		.din(new_net_19595),
		.dout(new_net_19596)
	);

	bfr new_net_19597_bfr_after (
		.din(new_net_19596),
		.dout(new_net_19597)
	);

	bfr new_net_19598_bfr_after (
		.din(new_net_19597),
		.dout(new_net_19598)
	);

	bfr new_net_19599_bfr_after (
		.din(new_net_19598),
		.dout(new_net_19599)
	);

	bfr new_net_19600_bfr_after (
		.din(new_net_19599),
		.dout(new_net_19600)
	);

	bfr new_net_19601_bfr_after (
		.din(new_net_19600),
		.dout(new_net_19601)
	);

	bfr new_net_19602_bfr_after (
		.din(new_net_19601),
		.dout(new_net_19602)
	);

	bfr new_net_19603_bfr_after (
		.din(new_net_19602),
		.dout(new_net_19603)
	);

	bfr new_net_19604_bfr_after (
		.din(new_net_19603),
		.dout(new_net_19604)
	);

	bfr new_net_19605_bfr_after (
		.din(new_net_19604),
		.dout(new_net_19605)
	);

	bfr new_net_19606_bfr_after (
		.din(new_net_19605),
		.dout(new_net_19606)
	);

	bfr new_net_19607_bfr_after (
		.din(new_net_19606),
		.dout(new_net_19607)
	);

	bfr new_net_19608_bfr_after (
		.din(new_net_19607),
		.dout(new_net_19608)
	);

	bfr new_net_19609_bfr_after (
		.din(new_net_19608),
		.dout(new_net_19609)
	);

	bfr new_net_19610_bfr_after (
		.din(new_net_19609),
		.dout(new_net_19610)
	);

	bfr new_net_19611_bfr_after (
		.din(new_net_19610),
		.dout(new_net_19611)
	);

	bfr new_net_19612_bfr_after (
		.din(new_net_19611),
		.dout(new_net_19612)
	);

	bfr new_net_19613_bfr_after (
		.din(new_net_19612),
		.dout(new_net_19613)
	);

	bfr new_net_19614_bfr_after (
		.din(new_net_19613),
		.dout(new_net_19614)
	);

	bfr new_net_19615_bfr_after (
		.din(new_net_19614),
		.dout(new_net_19615)
	);

	bfr new_net_19616_bfr_after (
		.din(new_net_19615),
		.dout(new_net_19616)
	);

	bfr new_net_19617_bfr_after (
		.din(new_net_19616),
		.dout(new_net_19617)
	);

	bfr new_net_19618_bfr_after (
		.din(new_net_19617),
		.dout(new_net_19618)
	);

	bfr new_net_19619_bfr_after (
		.din(new_net_19618),
		.dout(new_net_19619)
	);

	bfr new_net_19620_bfr_after (
		.din(new_net_19619),
		.dout(new_net_19620)
	);

	bfr new_net_19621_bfr_after (
		.din(new_net_19620),
		.dout(new_net_19621)
	);

	bfr new_net_19622_bfr_after (
		.din(new_net_19621),
		.dout(new_net_19622)
	);

	bfr new_net_19623_bfr_after (
		.din(new_net_19622),
		.dout(new_net_19623)
	);

	bfr new_net_19624_bfr_after (
		.din(new_net_19623),
		.dout(new_net_19624)
	);

	bfr new_net_19625_bfr_after (
		.din(new_net_19624),
		.dout(new_net_19625)
	);

	bfr new_net_19626_bfr_after (
		.din(new_net_19625),
		.dout(new_net_19626)
	);

	bfr N5672_bfr_after (
		.din(new_net_19626),
		.dout(N5672)
	);

	bfr new_net_3461_bfr_after (
		.din(_1806_),
		.dout(new_net_3461)
	);

	bfr new_net_3502_bfr_after (
		.din(_1098_),
		.dout(new_net_3502)
	);

	bfr new_net_3545_bfr_after (
		.din(_1247_),
		.dout(new_net_3545)
	);

	bfr new_net_3820_bfr_after (
		.din(_0594_),
		.dout(new_net_3820)
	);

	bfr new_net_3842_bfr_after (
		.din(_0686_),
		.dout(new_net_3842)
	);

	bfr new_net_3878_bfr_after (
		.din(_0852_),
		.dout(new_net_3878)
	);

	bfr new_net_3880_bfr_after (
		.din(_0858_),
		.dout(new_net_3880)
	);

	bfr new_net_3585_bfr_after (
		.din(_1409_),
		.dout(new_net_3585)
	);

	bfr new_net_3652_bfr_after (
		.din(_1710_),
		.dout(new_net_3652)
	);

	bfr new_net_3798_bfr_after (
		.din(_0499_),
		.dout(new_net_3798)
	);

	bfr new_net_3815_bfr_after (
		.din(_0577_),
		.dout(new_net_3815)
	);

	bfr new_net_3831_bfr_after (
		.din(_0650_),
		.dout(new_net_3831)
	);

	bfr new_net_3716_bfr_after (
		.din(_0148_),
		.dout(new_net_3716)
	);

	bfr new_net_3796_bfr_after (
		.din(_0493_),
		.dout(new_net_3796)
	);

	bfr new_net_3917_bfr_after (
		.din(_1012_),
		.dout(new_net_3917)
	);

	bfr new_net_3684_bfr_after (
		.din(_0009_),
		.dout(new_net_3684)
	);

	bfr new_net_3729_bfr_after (
		.din(_0191_),
		.dout(new_net_3729)
	);

	bfr new_net_3761_bfr_after (
		.din(_0353_),
		.dout(new_net_3761)
	);

	bfr new_net_3510_bfr_after (
		.din(_1122_),
		.dout(new_net_3510)
	);

	bfr new_net_3536_bfr_after (
		.din(_1202_),
		.dout(new_net_3536)
	);

	bfr new_net_3547_bfr_after (
		.din(_1253_),
		.dout(new_net_3547)
	);

	bfr new_net_3600_bfr_after (
		.din(_1481_),
		.dout(new_net_3600)
	);

	bfr new_net_3624_bfr_after (
		.din(_1559_),
		.dout(new_net_3624)
	);

	bfr new_net_3665_bfr_after (
		.din(_1756_),
		.dout(new_net_3665)
	);

	bfr new_net_3791_bfr_after (
		.din(_0476_),
		.dout(new_net_3791)
	);

	bfr new_net_19627_bfr_after (
		.din(new_net_3964),
		.dout(new_net_19627)
	);

	bfr new_net_19628_bfr_after (
		.din(new_net_19627),
		.dout(new_net_19628)
	);

	bfr new_net_19629_bfr_after (
		.din(new_net_19628),
		.dout(new_net_19629)
	);

	bfr new_net_19630_bfr_after (
		.din(new_net_19629),
		.dout(new_net_19630)
	);

	bfr new_net_19631_bfr_after (
		.din(new_net_19630),
		.dout(new_net_19631)
	);

	bfr new_net_19632_bfr_after (
		.din(new_net_19631),
		.dout(new_net_19632)
	);

	bfr new_net_19633_bfr_after (
		.din(new_net_19632),
		.dout(new_net_19633)
	);

	bfr new_net_19634_bfr_after (
		.din(new_net_19633),
		.dout(new_net_19634)
	);

	bfr new_net_19635_bfr_after (
		.din(new_net_19634),
		.dout(new_net_19635)
	);

	bfr new_net_19636_bfr_after (
		.din(new_net_19635),
		.dout(new_net_19636)
	);

	bfr new_net_19637_bfr_after (
		.din(new_net_19636),
		.dout(new_net_19637)
	);

	bfr new_net_19638_bfr_after (
		.din(new_net_19637),
		.dout(new_net_19638)
	);

	bfr new_net_19639_bfr_after (
		.din(new_net_19638),
		.dout(new_net_19639)
	);

	bfr new_net_19640_bfr_after (
		.din(new_net_19639),
		.dout(new_net_19640)
	);

	bfr new_net_19641_bfr_after (
		.din(new_net_19640),
		.dout(new_net_19641)
	);

	bfr new_net_19642_bfr_after (
		.din(new_net_19641),
		.dout(new_net_19642)
	);

	bfr new_net_19643_bfr_after (
		.din(new_net_19642),
		.dout(new_net_19643)
	);

	bfr new_net_19644_bfr_after (
		.din(new_net_19643),
		.dout(new_net_19644)
	);

	bfr new_net_19645_bfr_after (
		.din(new_net_19644),
		.dout(new_net_19645)
	);

	bfr N6240_bfr_after (
		.din(new_net_19645),
		.dout(N6240)
	);

	bfr new_net_3501_bfr_after (
		.din(_1095_),
		.dout(new_net_3501)
	);

	bfr new_net_3546_bfr_after (
		.din(_1250_),
		.dout(new_net_3546)
	);

	bfr new_net_3576_bfr_after (
		.din(_1360_),
		.dout(new_net_3576)
	);

	bfr new_net_3594_bfr_after (
		.din(_1436_),
		.dout(new_net_3594)
	);

	bfr new_net_3620_bfr_after (
		.din(_1546_),
		.dout(new_net_3620)
	);

	bfr new_net_3680_bfr_after (
		.din(_1834_),
		.dout(new_net_3680)
	);

	bfr new_net_3715_bfr_after (
		.din(_0145_),
		.dout(new_net_3715)
	);

	bfr new_net_3608_bfr_after (
		.din(_1507_),
		.dout(new_net_3608)
	);

	bfr new_net_3669_bfr_after (
		.din(_1769_),
		.dout(new_net_3669)
	);

	bfr new_net_3688_bfr_after (
		.din(_0023_),
		.dout(new_net_3688)
	);

	bfr new_net_3780_bfr_after (
		.din(_0415_),
		.dout(new_net_3780)
	);

	bfr new_net_3913_bfr_after (
		.din(_0998_),
		.dout(new_net_3913)
	);

	bfr new_net_3856_bfr_after (
		.din(_0750_),
		.dout(new_net_3856)
	);

	bfr new_net_3707_bfr_after (
		.din(_0118_),
		.dout(new_net_3707)
	);

	bfr new_net_3742_bfr_after (
		.din(_0264_),
		.dout(new_net_3742)
	);

	bfr new_net_3507_bfr_after (
		.din(_1113_),
		.dout(new_net_3507)
	);

	bfr new_net_3525_bfr_after (
		.din(_1185_),
		.dout(new_net_3525)
	);

	bfr new_net_3686_bfr_after (
		.din(_0016_),
		.dout(new_net_3686)
	);

	bfr new_net_3848_bfr_after (
		.din(_0724_),
		.dout(new_net_3848)
	);

	bfr new_net_3862_bfr_after (
		.din(_0786_),
		.dout(new_net_3862)
	);

	bfr new_net_3494_bfr_after (
		.din(_1058_),
		.dout(new_net_3494)
	);

	bfr new_net_3561_bfr_after (
		.din(_1315_),
		.dout(new_net_3561)
	);

	bfr new_net_3775_bfr_after (
		.din(_0399_),
		.dout(new_net_3775)
	);

	bfr new_net_3824_bfr_after (
		.din(_0607_),
		.dout(new_net_3824)
	);

	bfr new_net_3841_bfr_after (
		.din(_0683_),
		.dout(new_net_3841)
	);

	bfr new_net_3900_bfr_after (
		.din(_0944_),
		.dout(new_net_3900)
	);

	bfr new_net_3687_bfr_after (
		.din(_0019_),
		.dout(new_net_3687)
	);

	bfr new_net_3698_bfr_after (
		.din(_0056_),
		.dout(new_net_3698)
	);

	bfr new_net_3542_bfr_after (
		.din(_1238_),
		.dout(new_net_3542)
	);

	bfr new_net_3678_bfr_after (
		.din(_1799_),
		.dout(new_net_3678)
	);

	bfr new_net_3804_bfr_after (
		.din(_0519_),
		.dout(new_net_3804)
	);

	bfr new_net_3823_bfr_after (
		.din(_0604_),
		.dout(new_net_3823)
	);

	bfr new_net_3894_bfr_after (
		.din(_0916_),
		.dout(new_net_3894)
	);

	bfr new_net_3809_bfr_after (
		.din(_0558_),
		.dout(new_net_3809)
	);

	bfr new_net_3500_bfr_after (
		.din(_1092_),
		.dout(new_net_3500)
	);

	bfr new_net_3515_bfr_after (
		.din(_1155_),
		.dout(new_net_3515)
	);

	bfr new_net_3526_bfr_after (
		.din(_1188_),
		.dout(new_net_3526)
	);

	bfr new_net_3567_bfr_after (
		.din(_1333_),
		.dout(new_net_3567)
	);

	bfr new_net_3601_bfr_after (
		.din(_1484_),
		.dout(new_net_3601)
	);

	bfr new_net_3604_bfr_after (
		.din(_1494_),
		.dout(new_net_3604)
	);

	bfr new_net_3851_bfr_after (
		.din(_0734_),
		.dout(new_net_3851)
	);

	bfr new_net_3869_bfr_after (
		.din(_0809_),
		.dout(new_net_3869)
	);

	bfr new_net_3476_bfr_after (
		.din(_0774_),
		.dout(new_net_3476)
	);

	bfr new_net_3581_bfr_after (
		.din(_1397_),
		.dout(new_net_3581)
	);

	bfr new_net_3668_bfr_after (
		.din(_1766_),
		.dout(new_net_3668)
	);

	bfr new_net_3712_bfr_after (
		.din(_0135_),
		.dout(new_net_3712)
	);

	bfr new_net_3779_bfr_after (
		.din(_0412_),
		.dout(new_net_3779)
	);

	bfr new_net_3907_bfr_after (
		.din(_0974_),
		.dout(new_net_3907)
	);

	bfr new_net_3589_bfr_after (
		.din(_1421_),
		.dout(new_net_3589)
	);

	bfr new_net_3635_bfr_after (
		.din(_1624_),
		.dout(new_net_3635)
	);

	bfr new_net_3766_bfr_after (
		.din(_0369_),
		.dout(new_net_3766)
	);

	bfr new_net_3795_bfr_after (
		.din(_0489_),
		.dout(new_net_3795)
	);

	bfr new_net_3839_bfr_after (
		.din(_0676_),
		.dout(new_net_3839)
	);

	bfr new_net_3897_bfr_after (
		.din(_0934_),
		.dout(new_net_3897)
	);

	bfr new_net_3459_bfr_after (
		.din(_1741_),
		.dout(new_net_3459)
	);

	bfr new_net_3487_bfr_after (
		.din(_1037_),
		.dout(new_net_3487)
	);

	bfr new_net_3645_bfr_after (
		.din(_1657_),
		.dout(new_net_3645)
	);

	bfr new_net_3481_bfr_after (
		.din(_0936_),
		.dout(new_net_3481)
	);

	bfr new_net_3514_bfr_after (
		.din(_1152_),
		.dout(new_net_3514)
	);

	bfr new_net_3517_bfr_after (
		.din(_1161_),
		.dout(new_net_3517)
	);

	bfr new_net_3609_bfr_after (
		.din(_1510_),
		.dout(new_net_3609)
	);

	bfr new_net_3794_bfr_after (
		.din(_0486_),
		.dout(new_net_3794)
	);

	bfr new_net_3496_bfr_after (
		.din(_1064_),
		.dout(new_net_3496)
	);

	bfr new_net_3518_bfr_after (
		.din(_1164_),
		.dout(new_net_3518)
	);

	bfr new_net_3558_bfr_after (
		.din(_1306_),
		.dout(new_net_3558)
	);

	bfr new_net_3579_bfr_after (
		.din(_1391_),
		.dout(new_net_3579)
	);

	bfr new_net_3593_bfr_after (
		.din(_1433_),
		.dout(new_net_3593)
	);

	bfr new_net_3638_bfr_after (
		.din(_1634_),
		.dout(new_net_3638)
	);

	bfr new_net_3471_bfr_after (
		.din(_0481_),
		.dout(new_net_3471)
	);

	bfr new_net_3531_bfr_after (
		.din(_1197_),
		.dout(new_net_3531)
	);

	bfr new_net_3694_bfr_after (
		.din(_0042_),
		.dout(new_net_3694)
	);

	bfr new_net_3705_bfr_after (
		.din(_0080_),
		.dout(new_net_3705)
	);

	bfr new_net_3740_bfr_after (
		.din(_0257_),
		.dout(new_net_3740)
	);

	bfr new_net_3770_bfr_after (
		.din(_0382_),
		.dout(new_net_3770)
	);

	bfr new_net_3782_bfr_after (
		.din(_0422_),
		.dout(new_net_3782)
	);

	bfr new_net_3909_bfr_after (
		.din(_0981_),
		.dout(new_net_3909)
	);

	bfr new_net_3623_bfr_after (
		.din(_1555_),
		.dout(new_net_3623)
	);

	bfr new_net_3666_bfr_after (
		.din(_1759_),
		.dout(new_net_3666)
	);

	bfr new_net_3681_bfr_after (
		.din(_1837_),
		.dout(new_net_3681)
	);

	bfr new_net_3696_bfr_after (
		.din(_0049_),
		.dout(new_net_3696)
	);

	bfr new_net_3758_bfr_after (
		.din(_0316_),
		.dout(new_net_3758)
	);

	bfr new_net_3805_bfr_after (
		.din(_0522_),
		.dout(new_net_3805)
	);

	bfr new_net_19646_bfr_after (
		.din(new_net_3938),
		.dout(new_net_19646)
	);

	bfr new_net_19647_bfr_after (
		.din(new_net_19646),
		.dout(new_net_19647)
	);

	bfr new_net_19648_bfr_after (
		.din(new_net_19647),
		.dout(new_net_19648)
	);

	bfr N6280_bfr_after (
		.din(new_net_19648),
		.dout(N6280)
	);

	bfr new_net_3602_bfr_after (
		.din(_1487_),
		.dout(new_net_3602)
	);

	bfr new_net_3753_bfr_after (
		.din(_0300_),
		.dout(new_net_3753)
	);

	bfr new_net_3910_bfr_after (
		.din(_0984_),
		.dout(new_net_3910)
	);

	bfr new_net_3554_bfr_after (
		.din(_1274_),
		.dout(new_net_3554)
	);

	bfr new_net_3621_bfr_after (
		.din(_1549_),
		.dout(new_net_3621)
	);

	bfr new_net_3661_bfr_after (
		.din(_1743_),
		.dout(new_net_3661)
	);

	bfr new_net_3760_bfr_after (
		.din(_0323_),
		.dout(new_net_3760)
	);

	bfr new_net_3833_bfr_after (
		.din(_0657_),
		.dout(new_net_3833)
	);

	bfr new_net_19649_bfr_after (
		.din(new_net_3960),
		.dout(new_net_19649)
	);

	bfr new_net_19650_bfr_after (
		.din(new_net_19649),
		.dout(new_net_19650)
	);

	bfr new_net_19651_bfr_after (
		.din(new_net_19650),
		.dout(new_net_19651)
	);

	bfr new_net_19652_bfr_after (
		.din(new_net_19651),
		.dout(new_net_19652)
	);

	bfr new_net_19653_bfr_after (
		.din(new_net_19652),
		.dout(new_net_19653)
	);

	bfr new_net_19654_bfr_after (
		.din(new_net_19653),
		.dout(new_net_19654)
	);

	bfr new_net_19655_bfr_after (
		.din(new_net_19654),
		.dout(new_net_19655)
	);

	bfr new_net_19656_bfr_after (
		.din(new_net_19655),
		.dout(new_net_19656)
	);

	bfr new_net_19657_bfr_after (
		.din(new_net_19656),
		.dout(new_net_19657)
	);

	bfr new_net_19658_bfr_after (
		.din(new_net_19657),
		.dout(new_net_19658)
	);

	bfr new_net_19659_bfr_after (
		.din(new_net_19658),
		.dout(new_net_19659)
	);

	bfr new_net_19660_bfr_after (
		.din(new_net_19659),
		.dout(new_net_19660)
	);

	bfr new_net_19661_bfr_after (
		.din(new_net_19660),
		.dout(new_net_19661)
	);

	bfr new_net_19662_bfr_after (
		.din(new_net_19661),
		.dout(new_net_19662)
	);

	bfr new_net_19663_bfr_after (
		.din(new_net_19662),
		.dout(new_net_19663)
	);

	bfr new_net_19664_bfr_after (
		.din(new_net_19663),
		.dout(new_net_19664)
	);

	bfr new_net_19665_bfr_after (
		.din(new_net_19664),
		.dout(new_net_19665)
	);

	bfr new_net_19666_bfr_after (
		.din(new_net_19665),
		.dout(new_net_19666)
	);

	bfr new_net_19667_bfr_after (
		.din(new_net_19666),
		.dout(new_net_19667)
	);

	bfr new_net_19668_bfr_after (
		.din(new_net_19667),
		.dout(new_net_19668)
	);

	bfr new_net_19669_bfr_after (
		.din(new_net_19668),
		.dout(new_net_19669)
	);

	bfr new_net_19670_bfr_after (
		.din(new_net_19669),
		.dout(new_net_19670)
	);

	bfr new_net_19671_bfr_after (
		.din(new_net_19670),
		.dout(new_net_19671)
	);

	bfr new_net_19672_bfr_after (
		.din(new_net_19671),
		.dout(new_net_19672)
	);

	bfr new_net_19673_bfr_after (
		.din(new_net_19672),
		.dout(new_net_19673)
	);

	bfr new_net_19674_bfr_after (
		.din(new_net_19673),
		.dout(new_net_19674)
	);

	bfr new_net_19675_bfr_after (
		.din(new_net_19674),
		.dout(new_net_19675)
	);

	bfr new_net_19676_bfr_after (
		.din(new_net_19675),
		.dout(new_net_19676)
	);

	bfr new_net_19677_bfr_after (
		.din(new_net_19676),
		.dout(new_net_19677)
	);

	bfr new_net_19678_bfr_after (
		.din(new_net_19677),
		.dout(new_net_19678)
	);

	bfr new_net_19679_bfr_after (
		.din(new_net_19678),
		.dout(new_net_19679)
	);

	bfr new_net_19680_bfr_after (
		.din(new_net_19679),
		.dout(new_net_19680)
	);

	bfr new_net_19681_bfr_after (
		.din(new_net_19680),
		.dout(new_net_19681)
	);

	bfr new_net_19682_bfr_after (
		.din(new_net_19681),
		.dout(new_net_19682)
	);

	bfr new_net_19683_bfr_after (
		.din(new_net_19682),
		.dout(new_net_19683)
	);

	bfr new_net_19684_bfr_after (
		.din(new_net_19683),
		.dout(new_net_19684)
	);

	bfr new_net_19685_bfr_after (
		.din(new_net_19684),
		.dout(new_net_19685)
	);

	bfr new_net_19686_bfr_after (
		.din(new_net_19685),
		.dout(new_net_19686)
	);

	bfr new_net_19687_bfr_after (
		.din(new_net_19686),
		.dout(new_net_19687)
	);

	bfr new_net_19688_bfr_after (
		.din(new_net_19687),
		.dout(new_net_19688)
	);

	bfr new_net_19689_bfr_after (
		.din(new_net_19688),
		.dout(new_net_19689)
	);

	bfr new_net_19690_bfr_after (
		.din(new_net_19689),
		.dout(new_net_19690)
	);

	bfr new_net_19691_bfr_after (
		.din(new_net_19690),
		.dout(new_net_19691)
	);

	bfr new_net_19692_bfr_after (
		.din(new_net_19691),
		.dout(new_net_19692)
	);

	bfr new_net_19693_bfr_after (
		.din(new_net_19692),
		.dout(new_net_19693)
	);

	bfr new_net_19694_bfr_after (
		.din(new_net_19693),
		.dout(new_net_19694)
	);

	bfr new_net_19695_bfr_after (
		.din(new_net_19694),
		.dout(new_net_19695)
	);

	bfr N6170_bfr_after (
		.din(new_net_19695),
		.dout(N6170)
	);

	bfr new_net_3482_bfr_after (
		.din(_0968_),
		.dout(new_net_3482)
	);

	bfr new_net_3570_bfr_after (
		.din(_1342_),
		.dout(new_net_3570)
	);

	bfr new_net_3612_bfr_after (
		.din(_1520_),
		.dout(new_net_3612)
	);

	bfr new_net_3649_bfr_after (
		.din(_1670_),
		.dout(new_net_3649)
	);

	bfr new_net_3739_bfr_after (
		.din(_0254_),
		.dout(new_net_3739)
	);

	bfr new_net_3683_bfr_after (
		.din(_0006_),
		.dout(new_net_3683)
	);

	bfr new_net_3714_bfr_after (
		.din(_0141_),
		.dout(new_net_3714)
	);

	bfr new_net_3793_bfr_after (
		.din(_0483_),
		.dout(new_net_3793)
	);

	bfr new_net_3871_bfr_after (
		.din(_0815_),
		.dout(new_net_3871)
	);

	bfr new_net_19696_bfr_after (
		.din(new_net_3950),
		.dout(new_net_19696)
	);

	bfr new_net_19697_bfr_after (
		.din(new_net_19696),
		.dout(new_net_19697)
	);

	bfr new_net_19698_bfr_after (
		.din(new_net_19697),
		.dout(new_net_19698)
	);

	bfr new_net_19699_bfr_after (
		.din(new_net_19698),
		.dout(new_net_19699)
	);

	bfr new_net_19700_bfr_after (
		.din(new_net_19699),
		.dout(new_net_19700)
	);

	bfr new_net_19701_bfr_after (
		.din(new_net_19700),
		.dout(new_net_19701)
	);

	bfr new_net_19702_bfr_after (
		.din(new_net_19701),
		.dout(new_net_19702)
	);

	bfr new_net_19703_bfr_after (
		.din(new_net_19702),
		.dout(new_net_19703)
	);

	bfr new_net_19704_bfr_after (
		.din(new_net_19703),
		.dout(new_net_19704)
	);

	bfr new_net_19705_bfr_after (
		.din(new_net_19704),
		.dout(new_net_19705)
	);

	bfr new_net_19706_bfr_after (
		.din(new_net_19705),
		.dout(new_net_19706)
	);

	bfr new_net_19707_bfr_after (
		.din(new_net_19706),
		.dout(new_net_19707)
	);

	bfr new_net_19708_bfr_after (
		.din(new_net_19707),
		.dout(new_net_19708)
	);

	bfr new_net_19709_bfr_after (
		.din(new_net_19708),
		.dout(new_net_19709)
	);

	bfr new_net_19710_bfr_after (
		.din(new_net_19709),
		.dout(new_net_19710)
	);

	bfr new_net_19711_bfr_after (
		.din(new_net_19710),
		.dout(new_net_19711)
	);

	bfr new_net_19712_bfr_after (
		.din(new_net_19711),
		.dout(new_net_19712)
	);

	bfr new_net_19713_bfr_after (
		.din(new_net_19712),
		.dout(new_net_19713)
	);

	bfr new_net_19714_bfr_after (
		.din(new_net_19713),
		.dout(new_net_19714)
	);

	bfr new_net_19715_bfr_after (
		.din(new_net_19714),
		.dout(new_net_19715)
	);

	bfr new_net_19716_bfr_after (
		.din(new_net_19715),
		.dout(new_net_19716)
	);

	bfr new_net_19717_bfr_after (
		.din(new_net_19716),
		.dout(new_net_19717)
	);

	bfr new_net_19718_bfr_after (
		.din(new_net_19717),
		.dout(new_net_19718)
	);

	bfr new_net_19719_bfr_after (
		.din(new_net_19718),
		.dout(new_net_19719)
	);

	bfr new_net_19720_bfr_after (
		.din(new_net_19719),
		.dout(new_net_19720)
	);

	bfr new_net_19721_bfr_after (
		.din(new_net_19720),
		.dout(new_net_19721)
	);

	bfr new_net_19722_bfr_after (
		.din(new_net_19721),
		.dout(new_net_19722)
	);

	bfr new_net_19723_bfr_after (
		.din(new_net_19722),
		.dout(new_net_19723)
	);

	bfr new_net_19724_bfr_after (
		.din(new_net_19723),
		.dout(new_net_19724)
	);

	bfr new_net_19725_bfr_after (
		.din(new_net_19724),
		.dout(new_net_19725)
	);

	bfr new_net_19726_bfr_after (
		.din(new_net_19725),
		.dout(new_net_19726)
	);

	bfr new_net_19727_bfr_after (
		.din(new_net_19726),
		.dout(new_net_19727)
	);

	bfr new_net_19728_bfr_after (
		.din(new_net_19727),
		.dout(new_net_19728)
	);

	bfr new_net_19729_bfr_after (
		.din(new_net_19728),
		.dout(new_net_19729)
	);

	bfr new_net_19730_bfr_after (
		.din(new_net_19729),
		.dout(new_net_19730)
	);

	bfr new_net_19731_bfr_after (
		.din(new_net_19730),
		.dout(new_net_19731)
	);

	bfr new_net_19732_bfr_after (
		.din(new_net_19731),
		.dout(new_net_19732)
	);

	bfr new_net_19733_bfr_after (
		.din(new_net_19732),
		.dout(new_net_19733)
	);

	bfr new_net_19734_bfr_after (
		.din(new_net_19733),
		.dout(new_net_19734)
	);

	bfr new_net_19735_bfr_after (
		.din(new_net_19734),
		.dout(new_net_19735)
	);

	bfr new_net_19736_bfr_after (
		.din(new_net_19735),
		.dout(new_net_19736)
	);

	bfr new_net_19737_bfr_after (
		.din(new_net_19736),
		.dout(new_net_19737)
	);

	bfr new_net_19738_bfr_after (
		.din(new_net_19737),
		.dout(new_net_19738)
	);

	bfr new_net_19739_bfr_after (
		.din(new_net_19738),
		.dout(new_net_19739)
	);

	bfr new_net_19740_bfr_after (
		.din(new_net_19739),
		.dout(new_net_19740)
	);

	bfr new_net_19741_bfr_after (
		.din(new_net_19740),
		.dout(new_net_19741)
	);

	bfr new_net_19742_bfr_after (
		.din(new_net_19741),
		.dout(new_net_19742)
	);

	bfr new_net_19743_bfr_after (
		.din(new_net_19742),
		.dout(new_net_19743)
	);

	bfr new_net_19744_bfr_after (
		.din(new_net_19743),
		.dout(new_net_19744)
	);

	bfr new_net_19745_bfr_after (
		.din(new_net_19744),
		.dout(new_net_19745)
	);

	bfr new_net_19746_bfr_after (
		.din(new_net_19745),
		.dout(new_net_19746)
	);

	bfr new_net_19747_bfr_after (
		.din(new_net_19746),
		.dout(new_net_19747)
	);

	bfr new_net_19748_bfr_after (
		.din(new_net_19747),
		.dout(new_net_19748)
	);

	bfr new_net_19749_bfr_after (
		.din(new_net_19748),
		.dout(new_net_19749)
	);

	bfr new_net_19750_bfr_after (
		.din(new_net_19749),
		.dout(new_net_19750)
	);

	bfr new_net_19751_bfr_after (
		.din(new_net_19750),
		.dout(new_net_19751)
	);

	bfr new_net_19752_bfr_after (
		.din(new_net_19751),
		.dout(new_net_19752)
	);

	bfr new_net_19753_bfr_after (
		.din(new_net_19752),
		.dout(new_net_19753)
	);

	bfr new_net_19754_bfr_after (
		.din(new_net_19753),
		.dout(new_net_19754)
	);

	bfr new_net_19755_bfr_after (
		.din(new_net_19754),
		.dout(new_net_19755)
	);

	bfr new_net_19756_bfr_after (
		.din(new_net_19755),
		.dout(new_net_19756)
	);

	bfr new_net_19757_bfr_after (
		.din(new_net_19756),
		.dout(new_net_19757)
	);

	bfr new_net_19758_bfr_after (
		.din(new_net_19757),
		.dout(new_net_19758)
	);

	bfr new_net_19759_bfr_after (
		.din(new_net_19758),
		.dout(new_net_19759)
	);

	bfr new_net_19760_bfr_after (
		.din(new_net_19759),
		.dout(new_net_19760)
	);

	bfr new_net_19761_bfr_after (
		.din(new_net_19760),
		.dout(new_net_19761)
	);

	bfr new_net_19762_bfr_after (
		.din(new_net_19761),
		.dout(new_net_19762)
	);

	bfr new_net_19763_bfr_after (
		.din(new_net_19762),
		.dout(new_net_19763)
	);

	bfr new_net_19764_bfr_after (
		.din(new_net_19763),
		.dout(new_net_19764)
	);

	bfr new_net_19765_bfr_after (
		.din(new_net_19764),
		.dout(new_net_19765)
	);

	bfr new_net_19766_bfr_after (
		.din(new_net_19765),
		.dout(new_net_19766)
	);

	bfr new_net_19767_bfr_after (
		.din(new_net_19766),
		.dout(new_net_19767)
	);

	bfr new_net_19768_bfr_after (
		.din(new_net_19767),
		.dout(new_net_19768)
	);

	bfr new_net_19769_bfr_after (
		.din(new_net_19768),
		.dout(new_net_19769)
	);

	bfr new_net_19770_bfr_after (
		.din(new_net_19769),
		.dout(new_net_19770)
	);

	bfr new_net_19771_bfr_after (
		.din(new_net_19770),
		.dout(new_net_19771)
	);

	bfr new_net_19772_bfr_after (
		.din(new_net_19771),
		.dout(new_net_19772)
	);

	bfr new_net_19773_bfr_after (
		.din(new_net_19772),
		.dout(new_net_19773)
	);

	bfr new_net_19774_bfr_after (
		.din(new_net_19773),
		.dout(new_net_19774)
	);

	bfr new_net_19775_bfr_after (
		.din(new_net_19774),
		.dout(new_net_19775)
	);

	bfr new_net_19776_bfr_after (
		.din(new_net_19775),
		.dout(new_net_19776)
	);

	bfr new_net_19777_bfr_after (
		.din(new_net_19776),
		.dout(new_net_19777)
	);

	bfr new_net_19778_bfr_after (
		.din(new_net_19777),
		.dout(new_net_19778)
	);

	bfr new_net_19779_bfr_after (
		.din(new_net_19778),
		.dout(new_net_19779)
	);

	bfr new_net_19780_bfr_after (
		.din(new_net_19779),
		.dout(new_net_19780)
	);

	bfr new_net_19781_bfr_after (
		.din(new_net_19780),
		.dout(new_net_19781)
	);

	bfr new_net_19782_bfr_after (
		.din(new_net_19781),
		.dout(new_net_19782)
	);

	bfr new_net_19783_bfr_after (
		.din(new_net_19782),
		.dout(new_net_19783)
	);

	bfr new_net_19784_bfr_after (
		.din(new_net_19783),
		.dout(new_net_19784)
	);

	bfr new_net_19785_bfr_after (
		.din(new_net_19784),
		.dout(new_net_19785)
	);

	bfr new_net_19786_bfr_after (
		.din(new_net_19785),
		.dout(new_net_19786)
	);

	bfr new_net_19787_bfr_after (
		.din(new_net_19786),
		.dout(new_net_19787)
	);

	bfr new_net_19788_bfr_after (
		.din(new_net_19787),
		.dout(new_net_19788)
	);

	bfr new_net_19789_bfr_after (
		.din(new_net_19788),
		.dout(new_net_19789)
	);

	bfr new_net_19790_bfr_after (
		.din(new_net_19789),
		.dout(new_net_19790)
	);

	bfr new_net_19791_bfr_after (
		.din(new_net_19790),
		.dout(new_net_19791)
	);

	bfr new_net_19792_bfr_after (
		.din(new_net_19791),
		.dout(new_net_19792)
	);

	bfr new_net_19793_bfr_after (
		.din(new_net_19792),
		.dout(new_net_19793)
	);

	bfr new_net_19794_bfr_after (
		.din(new_net_19793),
		.dout(new_net_19794)
	);

	bfr new_net_19795_bfr_after (
		.din(new_net_19794),
		.dout(new_net_19795)
	);

	bfr new_net_19796_bfr_after (
		.din(new_net_19795),
		.dout(new_net_19796)
	);

	bfr new_net_19797_bfr_after (
		.din(new_net_19796),
		.dout(new_net_19797)
	);

	bfr new_net_19798_bfr_after (
		.din(new_net_19797),
		.dout(new_net_19798)
	);

	bfr new_net_19799_bfr_after (
		.din(new_net_19798),
		.dout(new_net_19799)
	);

	bfr new_net_19800_bfr_after (
		.din(new_net_19799),
		.dout(new_net_19800)
	);

	bfr new_net_19801_bfr_after (
		.din(new_net_19800),
		.dout(new_net_19801)
	);

	bfr new_net_19802_bfr_after (
		.din(new_net_19801),
		.dout(new_net_19802)
	);

	bfr new_net_19803_bfr_after (
		.din(new_net_19802),
		.dout(new_net_19803)
	);

	bfr new_net_19804_bfr_after (
		.din(new_net_19803),
		.dout(new_net_19804)
	);

	bfr new_net_19805_bfr_after (
		.din(new_net_19804),
		.dout(new_net_19805)
	);

	bfr new_net_19806_bfr_after (
		.din(new_net_19805),
		.dout(new_net_19806)
	);

	bfr new_net_19807_bfr_after (
		.din(new_net_19806),
		.dout(new_net_19807)
	);

	bfr new_net_19808_bfr_after (
		.din(new_net_19807),
		.dout(new_net_19808)
	);

	bfr new_net_19809_bfr_after (
		.din(new_net_19808),
		.dout(new_net_19809)
	);

	bfr new_net_19810_bfr_after (
		.din(new_net_19809),
		.dout(new_net_19810)
	);

	bfr new_net_19811_bfr_after (
		.din(new_net_19810),
		.dout(new_net_19811)
	);

	bfr new_net_19812_bfr_after (
		.din(new_net_19811),
		.dout(new_net_19812)
	);

	bfr new_net_19813_bfr_after (
		.din(new_net_19812),
		.dout(new_net_19813)
	);

	bfr new_net_19814_bfr_after (
		.din(new_net_19813),
		.dout(new_net_19814)
	);

	bfr new_net_19815_bfr_after (
		.din(new_net_19814),
		.dout(new_net_19815)
	);

	bfr new_net_19816_bfr_after (
		.din(new_net_19815),
		.dout(new_net_19816)
	);

	bfr new_net_19817_bfr_after (
		.din(new_net_19816),
		.dout(new_net_19817)
	);

	bfr new_net_19818_bfr_after (
		.din(new_net_19817),
		.dout(new_net_19818)
	);

	bfr new_net_19819_bfr_after (
		.din(new_net_19818),
		.dout(new_net_19819)
	);

	bfr new_net_19820_bfr_after (
		.din(new_net_19819),
		.dout(new_net_19820)
	);

	bfr new_net_19821_bfr_after (
		.din(new_net_19820),
		.dout(new_net_19821)
	);

	bfr new_net_19822_bfr_after (
		.din(new_net_19821),
		.dout(new_net_19822)
	);

	bfr new_net_19823_bfr_after (
		.din(new_net_19822),
		.dout(new_net_19823)
	);

	bfr new_net_19824_bfr_after (
		.din(new_net_19823),
		.dout(new_net_19824)
	);

	bfr new_net_19825_bfr_after (
		.din(new_net_19824),
		.dout(new_net_19825)
	);

	bfr new_net_19826_bfr_after (
		.din(new_net_19825),
		.dout(new_net_19826)
	);

	bfr N3211_bfr_after (
		.din(new_net_19826),
		.dout(N3211)
	);

	bfr new_net_3505_bfr_after (
		.din(_1107_),
		.dout(new_net_3505)
	);

	bfr new_net_3540_bfr_after (
		.din(_1232_),
		.dout(new_net_3540)
	);

	bfr new_net_3571_bfr_after (
		.din(_1345_),
		.dout(new_net_3571)
	);

	bfr new_net_3592_bfr_after (
		.din(_1430_),
		.dout(new_net_3592)
	);

	bfr new_net_3618_bfr_after (
		.din(_1540_),
		.dout(new_net_3618)
	);

	bfr new_net_3651_bfr_after (
		.din(_1677_),
		.dout(new_net_3651)
	);

	bfr new_net_3703_bfr_after (
		.din(_0072_),
		.dout(new_net_3703)
	);

	bfr new_net_3750_bfr_after (
		.din(_0290_),
		.dout(new_net_3750)
	);

	bfr new_net_3888_bfr_after (
		.din(_0896_),
		.dout(new_net_3888)
	);

	bfr new_net_3472_bfr_after (
		.din(_0514_),
		.dout(new_net_3472)
	);

	bfr new_net_3598_bfr_after (
		.din(_1448_),
		.dout(new_net_3598)
	);

	bfr new_net_3607_bfr_after (
		.din(_1504_),
		.dout(new_net_3607)
	);

	bfr new_net_3682_bfr_after (
		.din(_0003_),
		.dout(new_net_3682)
	);

	bfr new_net_3843_bfr_after (
		.din(_0690_),
		.dout(new_net_3843)
	);

	bfr new_net_19827_bfr_after (
		.din(new_net_3970),
		.dout(new_net_19827)
	);

	bfr new_net_19828_bfr_after (
		.din(new_net_19827),
		.dout(new_net_19828)
	);

	bfr new_net_19829_bfr_after (
		.din(new_net_19828),
		.dout(new_net_19829)
	);

	bfr new_net_19830_bfr_after (
		.din(new_net_19829),
		.dout(new_net_19830)
	);

	bfr new_net_19831_bfr_after (
		.din(new_net_19830),
		.dout(new_net_19831)
	);

	bfr new_net_19832_bfr_after (
		.din(new_net_19831),
		.dout(new_net_19832)
	);

	bfr new_net_19833_bfr_after (
		.din(new_net_19832),
		.dout(new_net_19833)
	);

	bfr new_net_19834_bfr_after (
		.din(new_net_19833),
		.dout(new_net_19834)
	);

	bfr new_net_19835_bfr_after (
		.din(new_net_19834),
		.dout(new_net_19835)
	);

	bfr new_net_19836_bfr_after (
		.din(new_net_19835),
		.dout(new_net_19836)
	);

	bfr new_net_19837_bfr_after (
		.din(new_net_19836),
		.dout(new_net_19837)
	);

	bfr new_net_19838_bfr_after (
		.din(new_net_19837),
		.dout(new_net_19838)
	);

	bfr new_net_19839_bfr_after (
		.din(new_net_19838),
		.dout(new_net_19839)
	);

	bfr new_net_19840_bfr_after (
		.din(new_net_19839),
		.dout(new_net_19840)
	);

	bfr new_net_19841_bfr_after (
		.din(new_net_19840),
		.dout(new_net_19841)
	);

	bfr new_net_19842_bfr_after (
		.din(new_net_19841),
		.dout(new_net_19842)
	);

	bfr new_net_19843_bfr_after (
		.din(new_net_19842),
		.dout(new_net_19843)
	);

	bfr new_net_19844_bfr_after (
		.din(new_net_19843),
		.dout(new_net_19844)
	);

	bfr new_net_19845_bfr_after (
		.din(new_net_19844),
		.dout(new_net_19845)
	);

	bfr new_net_19846_bfr_after (
		.din(new_net_19845),
		.dout(new_net_19846)
	);

	bfr new_net_19847_bfr_after (
		.din(new_net_19846),
		.dout(new_net_19847)
	);

	bfr new_net_19848_bfr_after (
		.din(new_net_19847),
		.dout(new_net_19848)
	);

	bfr new_net_19849_bfr_after (
		.din(new_net_19848),
		.dout(new_net_19849)
	);

	bfr new_net_19850_bfr_after (
		.din(new_net_19849),
		.dout(new_net_19850)
	);

	bfr new_net_19851_bfr_after (
		.din(new_net_19850),
		.dout(new_net_19851)
	);

	bfr new_net_19852_bfr_after (
		.din(new_net_19851),
		.dout(new_net_19852)
	);

	bfr new_net_19853_bfr_after (
		.din(new_net_19852),
		.dout(new_net_19853)
	);

	bfr new_net_19854_bfr_after (
		.din(new_net_19853),
		.dout(new_net_19854)
	);

	bfr new_net_19855_bfr_after (
		.din(new_net_19854),
		.dout(new_net_19855)
	);

	bfr new_net_19856_bfr_after (
		.din(new_net_19855),
		.dout(new_net_19856)
	);

	bfr new_net_19857_bfr_after (
		.din(new_net_19856),
		.dout(new_net_19857)
	);

	bfr new_net_19858_bfr_after (
		.din(new_net_19857),
		.dout(new_net_19858)
	);

	bfr new_net_19859_bfr_after (
		.din(new_net_19858),
		.dout(new_net_19859)
	);

	bfr new_net_19860_bfr_after (
		.din(new_net_19859),
		.dout(new_net_19860)
	);

	bfr new_net_19861_bfr_after (
		.din(new_net_19860),
		.dout(new_net_19861)
	);

	bfr new_net_19862_bfr_after (
		.din(new_net_19861),
		.dout(new_net_19862)
	);

	bfr new_net_19863_bfr_after (
		.din(new_net_19862),
		.dout(new_net_19863)
	);

	bfr new_net_19864_bfr_after (
		.din(new_net_19863),
		.dout(new_net_19864)
	);

	bfr new_net_19865_bfr_after (
		.din(new_net_19864),
		.dout(new_net_19865)
	);

	bfr N6190_bfr_after (
		.din(new_net_19865),
		.dout(N6190)
	);

	bfr new_net_3504_bfr_after (
		.din(_1104_),
		.dout(new_net_3504)
	);

	bfr new_net_3722_bfr_after (
		.din(_0168_),
		.dout(new_net_3722)
	);

	bfr new_net_3741_bfr_after (
		.din(_0260_),
		.dout(new_net_3741)
	);

	bfr new_net_3769_bfr_after (
		.din(_0379_),
		.dout(new_net_3769)
	);

	bfr new_net_3816_bfr_after (
		.din(_0581_),
		.dout(new_net_3816)
	);

	bfr new_net_3879_bfr_after (
		.din(_0855_),
		.dout(new_net_3879)
	);

	bfr new_net_19866_bfr_after (
		.din(new_net_3958),
		.dout(new_net_19866)
	);

	bfr new_net_19867_bfr_after (
		.din(new_net_19866),
		.dout(new_net_19867)
	);

	bfr new_net_19868_bfr_after (
		.din(new_net_19867),
		.dout(new_net_19868)
	);

	bfr new_net_19869_bfr_after (
		.din(new_net_19868),
		.dout(new_net_19869)
	);

	bfr new_net_19870_bfr_after (
		.din(new_net_19869),
		.dout(new_net_19870)
	);

	bfr new_net_19871_bfr_after (
		.din(new_net_19870),
		.dout(new_net_19871)
	);

	bfr new_net_19872_bfr_after (
		.din(new_net_19871),
		.dout(new_net_19872)
	);

	bfr new_net_19873_bfr_after (
		.din(new_net_19872),
		.dout(new_net_19873)
	);

	bfr new_net_19874_bfr_after (
		.din(new_net_19873),
		.dout(new_net_19874)
	);

	bfr new_net_19875_bfr_after (
		.din(new_net_19874),
		.dout(new_net_19875)
	);

	bfr new_net_19876_bfr_after (
		.din(new_net_19875),
		.dout(new_net_19876)
	);

	bfr new_net_19877_bfr_after (
		.din(new_net_19876),
		.dout(new_net_19877)
	);

	bfr new_net_19878_bfr_after (
		.din(new_net_19877),
		.dout(new_net_19878)
	);

	bfr new_net_19879_bfr_after (
		.din(new_net_19878),
		.dout(new_net_19879)
	);

	bfr new_net_19880_bfr_after (
		.din(new_net_19879),
		.dout(new_net_19880)
	);

	bfr new_net_19881_bfr_after (
		.din(new_net_19880),
		.dout(new_net_19881)
	);

	bfr new_net_19882_bfr_after (
		.din(new_net_19881),
		.dout(new_net_19882)
	);

	bfr new_net_19883_bfr_after (
		.din(new_net_19882),
		.dout(new_net_19883)
	);

	bfr new_net_19884_bfr_after (
		.din(new_net_19883),
		.dout(new_net_19884)
	);

	bfr new_net_19885_bfr_after (
		.din(new_net_19884),
		.dout(new_net_19885)
	);

	bfr new_net_19886_bfr_after (
		.din(new_net_19885),
		.dout(new_net_19886)
	);

	bfr new_net_19887_bfr_after (
		.din(new_net_19886),
		.dout(new_net_19887)
	);

	bfr new_net_19888_bfr_after (
		.din(new_net_19887),
		.dout(new_net_19888)
	);

	bfr new_net_19889_bfr_after (
		.din(new_net_19888),
		.dout(new_net_19889)
	);

	bfr new_net_19890_bfr_after (
		.din(new_net_19889),
		.dout(new_net_19890)
	);

	bfr new_net_19891_bfr_after (
		.din(new_net_19890),
		.dout(new_net_19891)
	);

	bfr new_net_19892_bfr_after (
		.din(new_net_19891),
		.dout(new_net_19892)
	);

	bfr new_net_19893_bfr_after (
		.din(new_net_19892),
		.dout(new_net_19893)
	);

	bfr new_net_19894_bfr_after (
		.din(new_net_19893),
		.dout(new_net_19894)
	);

	bfr new_net_19895_bfr_after (
		.din(new_net_19894),
		.dout(new_net_19895)
	);

	bfr new_net_19896_bfr_after (
		.din(new_net_19895),
		.dout(new_net_19896)
	);

	bfr new_net_19897_bfr_after (
		.din(new_net_19896),
		.dout(new_net_19897)
	);

	bfr new_net_19898_bfr_after (
		.din(new_net_19897),
		.dout(new_net_19898)
	);

	bfr new_net_19899_bfr_after (
		.din(new_net_19898),
		.dout(new_net_19899)
	);

	bfr new_net_19900_bfr_after (
		.din(new_net_19899),
		.dout(new_net_19900)
	);

	bfr new_net_19901_bfr_after (
		.din(new_net_19900),
		.dout(new_net_19901)
	);

	bfr new_net_19902_bfr_after (
		.din(new_net_19901),
		.dout(new_net_19902)
	);

	bfr new_net_19903_bfr_after (
		.din(new_net_19902),
		.dout(new_net_19903)
	);

	bfr new_net_19904_bfr_after (
		.din(new_net_19903),
		.dout(new_net_19904)
	);

	bfr new_net_19905_bfr_after (
		.din(new_net_19904),
		.dout(new_net_19905)
	);

	bfr new_net_19906_bfr_after (
		.din(new_net_19905),
		.dout(new_net_19906)
	);

	bfr new_net_19907_bfr_after (
		.din(new_net_19906),
		.dout(new_net_19907)
	);

	bfr new_net_19908_bfr_after (
		.din(new_net_19907),
		.dout(new_net_19908)
	);

	bfr new_net_19909_bfr_after (
		.din(new_net_19908),
		.dout(new_net_19909)
	);

	bfr new_net_19910_bfr_after (
		.din(new_net_19909),
		.dout(new_net_19910)
	);

	bfr new_net_19911_bfr_after (
		.din(new_net_19910),
		.dout(new_net_19911)
	);

	bfr new_net_19912_bfr_after (
		.din(new_net_19911),
		.dout(new_net_19912)
	);

	bfr new_net_19913_bfr_after (
		.din(new_net_19912),
		.dout(new_net_19913)
	);

	bfr new_net_19914_bfr_after (
		.din(new_net_19913),
		.dout(new_net_19914)
	);

	bfr new_net_19915_bfr_after (
		.din(new_net_19914),
		.dout(new_net_19915)
	);

	bfr new_net_19916_bfr_after (
		.din(new_net_19915),
		.dout(new_net_19916)
	);

	bfr new_net_19917_bfr_after (
		.din(new_net_19916),
		.dout(new_net_19917)
	);

	bfr new_net_19918_bfr_after (
		.din(new_net_19917),
		.dout(new_net_19918)
	);

	bfr new_net_19919_bfr_after (
		.din(new_net_19918),
		.dout(new_net_19919)
	);

	bfr new_net_19920_bfr_after (
		.din(new_net_19919),
		.dout(new_net_19920)
	);

	bfr new_net_19921_bfr_after (
		.din(new_net_19920),
		.dout(new_net_19921)
	);

	bfr new_net_19922_bfr_after (
		.din(new_net_19921),
		.dout(new_net_19922)
	);

	bfr new_net_19923_bfr_after (
		.din(new_net_19922),
		.dout(new_net_19923)
	);

	bfr new_net_19924_bfr_after (
		.din(new_net_19923),
		.dout(new_net_19924)
	);

	bfr new_net_19925_bfr_after (
		.din(new_net_19924),
		.dout(new_net_19925)
	);

	bfr new_net_19926_bfr_after (
		.din(new_net_19925),
		.dout(new_net_19926)
	);

	bfr new_net_19927_bfr_after (
		.din(new_net_19926),
		.dout(new_net_19927)
	);

	bfr new_net_19928_bfr_after (
		.din(new_net_19927),
		.dout(new_net_19928)
	);

	bfr new_net_19929_bfr_after (
		.din(new_net_19928),
		.dout(new_net_19929)
	);

	bfr new_net_19930_bfr_after (
		.din(new_net_19929),
		.dout(new_net_19930)
	);

	bfr new_net_19931_bfr_after (
		.din(new_net_19930),
		.dout(new_net_19931)
	);

	bfr new_net_19932_bfr_after (
		.din(new_net_19931),
		.dout(new_net_19932)
	);

	bfr new_net_19933_bfr_after (
		.din(new_net_19932),
		.dout(new_net_19933)
	);

	bfr new_net_19934_bfr_after (
		.din(new_net_19933),
		.dout(new_net_19934)
	);

	bfr new_net_19935_bfr_after (
		.din(new_net_19934),
		.dout(new_net_19935)
	);

	bfr new_net_19936_bfr_after (
		.din(new_net_19935),
		.dout(new_net_19936)
	);

	bfr new_net_19937_bfr_after (
		.din(new_net_19936),
		.dout(new_net_19937)
	);

	bfr new_net_19938_bfr_after (
		.din(new_net_19937),
		.dout(new_net_19938)
	);

	bfr new_net_19939_bfr_after (
		.din(new_net_19938),
		.dout(new_net_19939)
	);

	bfr new_net_19940_bfr_after (
		.din(new_net_19939),
		.dout(new_net_19940)
	);

	bfr new_net_19941_bfr_after (
		.din(new_net_19940),
		.dout(new_net_19941)
	);

	bfr new_net_19942_bfr_after (
		.din(new_net_19941),
		.dout(new_net_19942)
	);

	bfr new_net_19943_bfr_after (
		.din(new_net_19942),
		.dout(new_net_19943)
	);

	bfr new_net_19944_bfr_after (
		.din(new_net_19943),
		.dout(new_net_19944)
	);

	bfr new_net_19945_bfr_after (
		.din(new_net_19944),
		.dout(new_net_19945)
	);

	bfr new_net_19946_bfr_after (
		.din(new_net_19945),
		.dout(new_net_19946)
	);

	bfr new_net_19947_bfr_after (
		.din(new_net_19946),
		.dout(new_net_19947)
	);

	bfr new_net_19948_bfr_after (
		.din(new_net_19947),
		.dout(new_net_19948)
	);

	bfr new_net_19949_bfr_after (
		.din(new_net_19948),
		.dout(new_net_19949)
	);

	bfr new_net_19950_bfr_after (
		.din(new_net_19949),
		.dout(new_net_19950)
	);

	bfr new_net_19951_bfr_after (
		.din(new_net_19950),
		.dout(new_net_19951)
	);

	bfr new_net_19952_bfr_after (
		.din(new_net_19951),
		.dout(new_net_19952)
	);

	bfr new_net_19953_bfr_after (
		.din(new_net_19952),
		.dout(new_net_19953)
	);

	bfr new_net_19954_bfr_after (
		.din(new_net_19953),
		.dout(new_net_19954)
	);

	bfr new_net_19955_bfr_after (
		.din(new_net_19954),
		.dout(new_net_19955)
	);

	bfr new_net_19956_bfr_after (
		.din(new_net_19955),
		.dout(new_net_19956)
	);

	bfr new_net_19957_bfr_after (
		.din(new_net_19956),
		.dout(new_net_19957)
	);

	bfr new_net_19958_bfr_after (
		.din(new_net_19957),
		.dout(new_net_19958)
	);

	bfr new_net_19959_bfr_after (
		.din(new_net_19958),
		.dout(new_net_19959)
	);

	bfr new_net_19960_bfr_after (
		.din(new_net_19959),
		.dout(new_net_19960)
	);

	bfr new_net_19961_bfr_after (
		.din(new_net_19960),
		.dout(new_net_19961)
	);

	bfr new_net_19962_bfr_after (
		.din(new_net_19961),
		.dout(new_net_19962)
	);

	bfr new_net_19963_bfr_after (
		.din(new_net_19962),
		.dout(new_net_19963)
	);

	bfr new_net_19964_bfr_after (
		.din(new_net_19963),
		.dout(new_net_19964)
	);

	bfr new_net_19965_bfr_after (
		.din(new_net_19964),
		.dout(new_net_19965)
	);

	bfr new_net_19966_bfr_after (
		.din(new_net_19965),
		.dout(new_net_19966)
	);

	bfr new_net_19967_bfr_after (
		.din(new_net_19966),
		.dout(new_net_19967)
	);

	bfr new_net_19968_bfr_after (
		.din(new_net_19967),
		.dout(new_net_19968)
	);

	bfr new_net_19969_bfr_after (
		.din(new_net_19968),
		.dout(new_net_19969)
	);

	bfr new_net_19970_bfr_after (
		.din(new_net_19969),
		.dout(new_net_19970)
	);

	bfr new_net_19971_bfr_after (
		.din(new_net_19970),
		.dout(new_net_19971)
	);

	bfr new_net_19972_bfr_after (
		.din(new_net_19971),
		.dout(new_net_19972)
	);

	bfr new_net_19973_bfr_after (
		.din(new_net_19972),
		.dout(new_net_19973)
	);

	bfr new_net_19974_bfr_after (
		.din(new_net_19973),
		.dout(new_net_19974)
	);

	bfr new_net_19975_bfr_after (
		.din(new_net_19974),
		.dout(new_net_19975)
	);

	bfr new_net_19976_bfr_after (
		.din(new_net_19975),
		.dout(new_net_19976)
	);

	bfr new_net_19977_bfr_after (
		.din(new_net_19976),
		.dout(new_net_19977)
	);

	bfr new_net_19978_bfr_after (
		.din(new_net_19977),
		.dout(new_net_19978)
	);

	bfr new_net_19979_bfr_after (
		.din(new_net_19978),
		.dout(new_net_19979)
	);

	bfr new_net_19980_bfr_after (
		.din(new_net_19979),
		.dout(new_net_19980)
	);

	bfr new_net_19981_bfr_after (
		.din(new_net_19980),
		.dout(new_net_19981)
	);

	bfr new_net_19982_bfr_after (
		.din(new_net_19981),
		.dout(new_net_19982)
	);

	bfr new_net_19983_bfr_after (
		.din(new_net_19982),
		.dout(new_net_19983)
	);

	bfr new_net_19984_bfr_after (
		.din(new_net_19983),
		.dout(new_net_19984)
	);

	bfr new_net_19985_bfr_after (
		.din(new_net_19984),
		.dout(new_net_19985)
	);

	bfr new_net_19986_bfr_after (
		.din(new_net_19985),
		.dout(new_net_19986)
	);

	bfr new_net_19987_bfr_after (
		.din(new_net_19986),
		.dout(new_net_19987)
	);

	bfr new_net_19988_bfr_after (
		.din(new_net_19987),
		.dout(new_net_19988)
	);

	bfr new_net_19989_bfr_after (
		.din(new_net_19988),
		.dout(new_net_19989)
	);

	bfr new_net_19990_bfr_after (
		.din(new_net_19989),
		.dout(new_net_19990)
	);

	bfr new_net_19991_bfr_after (
		.din(new_net_19990),
		.dout(new_net_19991)
	);

	bfr new_net_19992_bfr_after (
		.din(new_net_19991),
		.dout(new_net_19992)
	);

	bfr new_net_19993_bfr_after (
		.din(new_net_19992),
		.dout(new_net_19993)
	);

	bfr new_net_19994_bfr_after (
		.din(new_net_19993),
		.dout(new_net_19994)
	);

	bfr new_net_19995_bfr_after (
		.din(new_net_19994),
		.dout(new_net_19995)
	);

	bfr new_net_19996_bfr_after (
		.din(new_net_19995),
		.dout(new_net_19996)
	);

	bfr new_net_19997_bfr_after (
		.din(new_net_19996),
		.dout(new_net_19997)
	);

	bfr new_net_19998_bfr_after (
		.din(new_net_19997),
		.dout(new_net_19998)
	);

	bfr new_net_19999_bfr_after (
		.din(new_net_19998),
		.dout(new_net_19999)
	);

	bfr new_net_20000_bfr_after (
		.din(new_net_19999),
		.dout(new_net_20000)
	);

	bfr new_net_20001_bfr_after (
		.din(new_net_20000),
		.dout(new_net_20001)
	);

	bfr new_net_20002_bfr_after (
		.din(new_net_20001),
		.dout(new_net_20002)
	);

	bfr new_net_20003_bfr_after (
		.din(new_net_20002),
		.dout(new_net_20003)
	);

	bfr new_net_20004_bfr_after (
		.din(new_net_20003),
		.dout(new_net_20004)
	);

	bfr new_net_20005_bfr_after (
		.din(new_net_20004),
		.dout(new_net_20005)
	);

	bfr new_net_20006_bfr_after (
		.din(new_net_20005),
		.dout(new_net_20006)
	);

	bfr new_net_20007_bfr_after (
		.din(new_net_20006),
		.dout(new_net_20007)
	);

	bfr new_net_20008_bfr_after (
		.din(new_net_20007),
		.dout(new_net_20008)
	);

	bfr new_net_20009_bfr_after (
		.din(new_net_20008),
		.dout(new_net_20009)
	);

	bfr new_net_20010_bfr_after (
		.din(new_net_20009),
		.dout(new_net_20010)
	);

	bfr new_net_20011_bfr_after (
		.din(new_net_20010),
		.dout(new_net_20011)
	);

	bfr new_net_20012_bfr_after (
		.din(new_net_20011),
		.dout(new_net_20012)
	);

	bfr new_net_20013_bfr_after (
		.din(new_net_20012),
		.dout(new_net_20013)
	);

	bfr new_net_20014_bfr_after (
		.din(new_net_20013),
		.dout(new_net_20014)
	);

	bfr new_net_20015_bfr_after (
		.din(new_net_20014),
		.dout(new_net_20015)
	);

	bfr new_net_20016_bfr_after (
		.din(new_net_20015),
		.dout(new_net_20016)
	);

	bfr new_net_20017_bfr_after (
		.din(new_net_20016),
		.dout(new_net_20017)
	);

	bfr new_net_20018_bfr_after (
		.din(new_net_20017),
		.dout(new_net_20018)
	);

	bfr new_net_20019_bfr_after (
		.din(new_net_20018),
		.dout(new_net_20019)
	);

	bfr new_net_20020_bfr_after (
		.din(new_net_20019),
		.dout(new_net_20020)
	);

	bfr new_net_20021_bfr_after (
		.din(new_net_20020),
		.dout(new_net_20021)
	);

	bfr new_net_20022_bfr_after (
		.din(new_net_20021),
		.dout(new_net_20022)
	);

	bfr new_net_20023_bfr_after (
		.din(new_net_20022),
		.dout(new_net_20023)
	);

	bfr new_net_20024_bfr_after (
		.din(new_net_20023),
		.dout(new_net_20024)
	);

	bfr new_net_20025_bfr_after (
		.din(new_net_20024),
		.dout(new_net_20025)
	);

	bfr new_net_20026_bfr_after (
		.din(new_net_20025),
		.dout(new_net_20026)
	);

	bfr new_net_20027_bfr_after (
		.din(new_net_20026),
		.dout(new_net_20027)
	);

	bfr new_net_20028_bfr_after (
		.din(new_net_20027),
		.dout(new_net_20028)
	);

	bfr new_net_20029_bfr_after (
		.din(new_net_20028),
		.dout(new_net_20029)
	);

	bfr new_net_20030_bfr_after (
		.din(new_net_20029),
		.dout(new_net_20030)
	);

	bfr new_net_20031_bfr_after (
		.din(new_net_20030),
		.dout(new_net_20031)
	);

	bfr new_net_20032_bfr_after (
		.din(new_net_20031),
		.dout(new_net_20032)
	);

	bfr new_net_20033_bfr_after (
		.din(new_net_20032),
		.dout(new_net_20033)
	);

	bfr new_net_20034_bfr_after (
		.din(new_net_20033),
		.dout(new_net_20034)
	);

	bfr new_net_20035_bfr_after (
		.din(new_net_20034),
		.dout(new_net_20035)
	);

	bfr new_net_20036_bfr_after (
		.din(new_net_20035),
		.dout(new_net_20036)
	);

	bfr N1581_bfr_after (
		.din(new_net_20036),
		.dout(N1581)
	);

	bfr new_net_3692_bfr_after (
		.din(_0036_),
		.dout(new_net_3692)
	);

	bfr new_net_3754_bfr_after (
		.din(_0303_),
		.dout(new_net_3754)
	);

	bfr new_net_3491_bfr_after (
		.din(_1049_),
		.dout(new_net_3491)
	);

	bfr new_net_3555_bfr_after (
		.din(_1277_),
		.dout(new_net_3555)
	);

	bfr new_net_3840_bfr_after (
		.din(_0680_),
		.dout(new_net_3840)
	);

	bfr new_net_3911_bfr_after (
		.din(_0992_),
		.dout(new_net_3911)
	);

	bfr new_net_3549_bfr_after (
		.din(_1259_),
		.dout(new_net_3549)
	);

	bfr new_net_3719_bfr_after (
		.din(_0158_),
		.dout(new_net_3719)
	);

	bfr new_net_3778_bfr_after (
		.din(_0409_),
		.dout(new_net_3778)
	);

	bfr new_net_3837_bfr_after (
		.din(_0670_),
		.dout(new_net_3837)
	);

	bfr new_net_3853_bfr_after (
		.din(_0740_),
		.dout(new_net_3853)
	);

	bfr new_net_3902_bfr_after (
		.din(_0951_),
		.dout(new_net_3902)
	);

	bfr new_net_3744_bfr_after (
		.din(_0270_),
		.dout(new_net_3744)
	);

	bfr new_net_3568_bfr_after (
		.din(_1336_),
		.dout(new_net_3568)
	);

	bfr new_net_3676_bfr_after (
		.din(_1792_),
		.dout(new_net_3676)
	);

	bfr new_net_3699_bfr_after (
		.din(_0059_),
		.dout(new_net_3699)
	);

	bfr new_net_3797_bfr_after (
		.din(_0496_),
		.dout(new_net_3797)
	);

	bfr new_net_3520_bfr_after (
		.din(_1170_),
		.dout(new_net_3520)
	);

	bfr new_net_3614_bfr_after (
		.din(_1527_),
		.dout(new_net_3614)
	);

	bfr new_net_3667_bfr_after (
		.din(_1762_),
		.dout(new_net_3667)
	);

	bfr new_net_3749_bfr_after (
		.din(_0287_),
		.dout(new_net_3749)
	);

	bfr new_net_20037_bfr_after (
		.din(new_net_3922),
		.dout(new_net_20037)
	);

	bfr new_net_20038_bfr_after (
		.din(new_net_20037),
		.dout(new_net_20038)
	);

	bfr new_net_20039_bfr_after (
		.din(new_net_20038),
		.dout(new_net_20039)
	);

	bfr new_net_20040_bfr_after (
		.din(new_net_20039),
		.dout(new_net_20040)
	);

	bfr new_net_20041_bfr_after (
		.din(new_net_20040),
		.dout(new_net_20041)
	);

	bfr new_net_20042_bfr_after (
		.din(new_net_20041),
		.dout(new_net_20042)
	);

	bfr new_net_20043_bfr_after (
		.din(new_net_20042),
		.dout(new_net_20043)
	);

	bfr new_net_20044_bfr_after (
		.din(new_net_20043),
		.dout(new_net_20044)
	);

	bfr new_net_20045_bfr_after (
		.din(new_net_20044),
		.dout(new_net_20045)
	);

	bfr new_net_20046_bfr_after (
		.din(new_net_20045),
		.dout(new_net_20046)
	);

	bfr new_net_20047_bfr_after (
		.din(new_net_20046),
		.dout(new_net_20047)
	);

	bfr new_net_20048_bfr_after (
		.din(new_net_20047),
		.dout(new_net_20048)
	);

	bfr new_net_20049_bfr_after (
		.din(new_net_20048),
		.dout(new_net_20049)
	);

	bfr new_net_20050_bfr_after (
		.din(new_net_20049),
		.dout(new_net_20050)
	);

	bfr new_net_20051_bfr_after (
		.din(new_net_20050),
		.dout(new_net_20051)
	);

	bfr new_net_20052_bfr_after (
		.din(new_net_20051),
		.dout(new_net_20052)
	);

	bfr new_net_20053_bfr_after (
		.din(new_net_20052),
		.dout(new_net_20053)
	);

	bfr new_net_20054_bfr_after (
		.din(new_net_20053),
		.dout(new_net_20054)
	);

	bfr new_net_20055_bfr_after (
		.din(new_net_20054),
		.dout(new_net_20055)
	);

	bfr new_net_20056_bfr_after (
		.din(new_net_20055),
		.dout(new_net_20056)
	);

	bfr new_net_20057_bfr_after (
		.din(new_net_20056),
		.dout(new_net_20057)
	);

	bfr new_net_20058_bfr_after (
		.din(new_net_20057),
		.dout(new_net_20058)
	);

	bfr new_net_20059_bfr_after (
		.din(new_net_20058),
		.dout(new_net_20059)
	);

	bfr new_net_20060_bfr_after (
		.din(new_net_20059),
		.dout(new_net_20060)
	);

	bfr new_net_20061_bfr_after (
		.din(new_net_20060),
		.dout(new_net_20061)
	);

	bfr new_net_20062_bfr_after (
		.din(new_net_20061),
		.dout(new_net_20062)
	);

	bfr new_net_20063_bfr_after (
		.din(new_net_20062),
		.dout(new_net_20063)
	);

	bfr new_net_20064_bfr_after (
		.din(new_net_20063),
		.dout(new_net_20064)
	);

	bfr new_net_20065_bfr_after (
		.din(new_net_20064),
		.dout(new_net_20065)
	);

	bfr new_net_20066_bfr_after (
		.din(new_net_20065),
		.dout(new_net_20066)
	);

	bfr new_net_20067_bfr_after (
		.din(new_net_20066),
		.dout(new_net_20067)
	);

	bfr new_net_20068_bfr_after (
		.din(new_net_20067),
		.dout(new_net_20068)
	);

	bfr new_net_20069_bfr_after (
		.din(new_net_20068),
		.dout(new_net_20069)
	);

	bfr new_net_20070_bfr_after (
		.din(new_net_20069),
		.dout(new_net_20070)
	);

	bfr new_net_20071_bfr_after (
		.din(new_net_20070),
		.dout(new_net_20071)
	);

	bfr new_net_20072_bfr_after (
		.din(new_net_20071),
		.dout(new_net_20072)
	);

	bfr new_net_20073_bfr_after (
		.din(new_net_20072),
		.dout(new_net_20073)
	);

	bfr new_net_20074_bfr_after (
		.din(new_net_20073),
		.dout(new_net_20074)
	);

	bfr new_net_20075_bfr_after (
		.din(new_net_20074),
		.dout(new_net_20075)
	);

	bfr new_net_20076_bfr_after (
		.din(new_net_20075),
		.dout(new_net_20076)
	);

	bfr new_net_20077_bfr_after (
		.din(new_net_20076),
		.dout(new_net_20077)
	);

	bfr new_net_20078_bfr_after (
		.din(new_net_20077),
		.dout(new_net_20078)
	);

	bfr new_net_20079_bfr_after (
		.din(new_net_20078),
		.dout(new_net_20079)
	);

	bfr new_net_20080_bfr_after (
		.din(new_net_20079),
		.dout(new_net_20080)
	);

	bfr new_net_20081_bfr_after (
		.din(new_net_20080),
		.dout(new_net_20081)
	);

	bfr new_net_20082_bfr_after (
		.din(new_net_20081),
		.dout(new_net_20082)
	);

	bfr new_net_20083_bfr_after (
		.din(new_net_20082),
		.dout(new_net_20083)
	);

	bfr new_net_20084_bfr_after (
		.din(new_net_20083),
		.dout(new_net_20084)
	);

	bfr new_net_20085_bfr_after (
		.din(new_net_20084),
		.dout(new_net_20085)
	);

	bfr new_net_20086_bfr_after (
		.din(new_net_20085),
		.dout(new_net_20086)
	);

	bfr new_net_20087_bfr_after (
		.din(new_net_20086),
		.dout(new_net_20087)
	);

	bfr new_net_20088_bfr_after (
		.din(new_net_20087),
		.dout(new_net_20088)
	);

	bfr new_net_20089_bfr_after (
		.din(new_net_20088),
		.dout(new_net_20089)
	);

	bfr new_net_20090_bfr_after (
		.din(new_net_20089),
		.dout(new_net_20090)
	);

	bfr new_net_20091_bfr_after (
		.din(new_net_20090),
		.dout(new_net_20091)
	);

	bfr new_net_20092_bfr_after (
		.din(new_net_20091),
		.dout(new_net_20092)
	);

	bfr new_net_20093_bfr_after (
		.din(new_net_20092),
		.dout(new_net_20093)
	);

	bfr new_net_20094_bfr_after (
		.din(new_net_20093),
		.dout(new_net_20094)
	);

	bfr new_net_20095_bfr_after (
		.din(new_net_20094),
		.dout(new_net_20095)
	);

	bfr new_net_20096_bfr_after (
		.din(new_net_20095),
		.dout(new_net_20096)
	);

	bfr new_net_20097_bfr_after (
		.din(new_net_20096),
		.dout(new_net_20097)
	);

	bfr new_net_20098_bfr_after (
		.din(new_net_20097),
		.dout(new_net_20098)
	);

	bfr new_net_20099_bfr_after (
		.din(new_net_20098),
		.dout(new_net_20099)
	);

	bfr new_net_20100_bfr_after (
		.din(new_net_20099),
		.dout(new_net_20100)
	);

	bfr new_net_20101_bfr_after (
		.din(new_net_20100),
		.dout(new_net_20101)
	);

	bfr new_net_20102_bfr_after (
		.din(new_net_20101),
		.dout(new_net_20102)
	);

	bfr new_net_20103_bfr_after (
		.din(new_net_20102),
		.dout(new_net_20103)
	);

	bfr new_net_20104_bfr_after (
		.din(new_net_20103),
		.dout(new_net_20104)
	);

	bfr new_net_20105_bfr_after (
		.din(new_net_20104),
		.dout(new_net_20105)
	);

	bfr new_net_20106_bfr_after (
		.din(new_net_20105),
		.dout(new_net_20106)
	);

	bfr new_net_20107_bfr_after (
		.din(new_net_20106),
		.dout(new_net_20107)
	);

	bfr new_net_20108_bfr_after (
		.din(new_net_20107),
		.dout(new_net_20108)
	);

	bfr new_net_20109_bfr_after (
		.din(new_net_20108),
		.dout(new_net_20109)
	);

	bfr new_net_20110_bfr_after (
		.din(new_net_20109),
		.dout(new_net_20110)
	);

	bfr new_net_20111_bfr_after (
		.din(new_net_20110),
		.dout(new_net_20111)
	);

	bfr new_net_20112_bfr_after (
		.din(new_net_20111),
		.dout(new_net_20112)
	);

	bfr new_net_20113_bfr_after (
		.din(new_net_20112),
		.dout(new_net_20113)
	);

	bfr new_net_20114_bfr_after (
		.din(new_net_20113),
		.dout(new_net_20114)
	);

	bfr new_net_20115_bfr_after (
		.din(new_net_20114),
		.dout(new_net_20115)
	);

	bfr new_net_20116_bfr_after (
		.din(new_net_20115),
		.dout(new_net_20116)
	);

	bfr new_net_20117_bfr_after (
		.din(new_net_20116),
		.dout(new_net_20117)
	);

	bfr new_net_20118_bfr_after (
		.din(new_net_20117),
		.dout(new_net_20118)
	);

	bfr new_net_20119_bfr_after (
		.din(new_net_20118),
		.dout(new_net_20119)
	);

	bfr new_net_20120_bfr_after (
		.din(new_net_20119),
		.dout(new_net_20120)
	);

	bfr new_net_20121_bfr_after (
		.din(new_net_20120),
		.dout(new_net_20121)
	);

	bfr new_net_20122_bfr_after (
		.din(new_net_20121),
		.dout(new_net_20122)
	);

	bfr new_net_20123_bfr_after (
		.din(new_net_20122),
		.dout(new_net_20123)
	);

	bfr new_net_20124_bfr_after (
		.din(new_net_20123),
		.dout(new_net_20124)
	);

	bfr new_net_20125_bfr_after (
		.din(new_net_20124),
		.dout(new_net_20125)
	);

	bfr new_net_20126_bfr_after (
		.din(new_net_20125),
		.dout(new_net_20126)
	);

	bfr new_net_20127_bfr_after (
		.din(new_net_20126),
		.dout(new_net_20127)
	);

	bfr new_net_20128_bfr_after (
		.din(new_net_20127),
		.dout(new_net_20128)
	);

	bfr new_net_20129_bfr_after (
		.din(new_net_20128),
		.dout(new_net_20129)
	);

	bfr new_net_20130_bfr_after (
		.din(new_net_20129),
		.dout(new_net_20130)
	);

	bfr new_net_20131_bfr_after (
		.din(new_net_20130),
		.dout(new_net_20131)
	);

	bfr new_net_20132_bfr_after (
		.din(new_net_20131),
		.dout(new_net_20132)
	);

	bfr new_net_20133_bfr_after (
		.din(new_net_20132),
		.dout(new_net_20133)
	);

	bfr new_net_20134_bfr_after (
		.din(new_net_20133),
		.dout(new_net_20134)
	);

	bfr new_net_20135_bfr_after (
		.din(new_net_20134),
		.dout(new_net_20135)
	);

	bfr N4591_bfr_after (
		.din(new_net_20135),
		.dout(N4591)
	);

	bfr new_net_3553_bfr_after (
		.din(_1271_),
		.dout(new_net_3553)
	);

	bfr new_net_3646_bfr_after (
		.din(_1660_),
		.dout(new_net_3646)
	);

	bfr new_net_3835_bfr_after (
		.din(_0663_),
		.dout(new_net_3835)
	);

	bfr new_net_3891_bfr_after (
		.din(_0906_),
		.dout(new_net_3891)
	);

	bfr new_net_3915_bfr_after (
		.din(_1007_),
		.dout(new_net_3915)
	);

	bfr new_net_3457_bfr_after (
		.din(_1676_),
		.dout(new_net_3457)
	);

	bfr new_net_3466_bfr_after (
		.din(_0209_),
		.dout(new_net_3466)
	);

	bfr new_net_3735_bfr_after (
		.din(_0240_),
		.dout(new_net_3735)
	);

	bfr new_net_3747_bfr_after (
		.din(_0280_),
		.dout(new_net_3747)
	);

	bfr new_net_3772_bfr_after (
		.din(_0389_),
		.dout(new_net_3772)
	);

	bfr new_net_3781_bfr_after (
		.din(_0419_),
		.dout(new_net_3781)
	);

	bfr new_net_3822_bfr_after (
		.din(_0600_),
		.dout(new_net_3822)
	);

	bfr new_net_3914_bfr_after (
		.din(_1002_),
		.dout(new_net_3914)
	);

	bfr new_net_3478_bfr_after (
		.din(_0839_),
		.dout(new_net_3478)
	);

	bfr new_net_3615_bfr_after (
		.din(_1530_),
		.dout(new_net_3615)
	);

	bfr new_net_3818_bfr_after (
		.din(_0587_),
		.dout(new_net_3818)
	);

	bfr new_net_3860_bfr_after (
		.din(_0763_),
		.dout(new_net_3860)
	);

	bfr new_net_3544_bfr_after (
		.din(_1244_),
		.dout(new_net_3544)
	);

	bfr new_net_3586_bfr_after (
		.din(_1412_),
		.dout(new_net_3586)
	);

	bfr new_net_3641_bfr_after (
		.din(_1644_),
		.dout(new_net_3641)
	);

	bfr new_net_3777_bfr_after (
		.din(_0406_),
		.dout(new_net_3777)
	);

	bfr new_net_3806_bfr_after (
		.din(_0526_),
		.dout(new_net_3806)
	);

	bfr new_net_3873_bfr_after (
		.din(_0822_),
		.dout(new_net_3873)
	);

	bfr new_net_3611_bfr_after (
		.din(_1517_),
		.dout(new_net_3611)
	);

	bfr new_net_3826_bfr_after (
		.din(_0614_),
		.dout(new_net_3826)
	);

	bfr new_net_3895_bfr_after (
		.din(_0919_),
		.dout(new_net_3895)
	);

	bfr new_net_3557_bfr_after (
		.din(_1303_),
		.dout(new_net_3557)
	);

	bfr new_net_3577_bfr_after (
		.din(_1385_),
		.dout(new_net_3577)
	);

	bfr new_net_3632_bfr_after (
		.din(_1614_),
		.dout(new_net_3632)
	);

	bfr new_net_3643_bfr_after (
		.din(_1650_),
		.dout(new_net_3643)
	);

	bfr new_net_3670_bfr_after (
		.din(_1772_),
		.dout(new_net_3670)
	);

	bfr new_net_3858_bfr_after (
		.din(_0757_),
		.dout(new_net_3858)
	);

	bfr new_net_20136_bfr_after (
		.din(new_net_3930),
		.dout(new_net_20136)
	);

	bfr new_net_20137_bfr_after (
		.din(new_net_20136),
		.dout(new_net_20137)
	);

	bfr new_net_20138_bfr_after (
		.din(new_net_20137),
		.dout(new_net_20138)
	);

	bfr new_net_20139_bfr_after (
		.din(new_net_20138),
		.dout(new_net_20139)
	);

	bfr new_net_20140_bfr_after (
		.din(new_net_20139),
		.dout(new_net_20140)
	);

	bfr new_net_20141_bfr_after (
		.din(new_net_20140),
		.dout(new_net_20141)
	);

	bfr new_net_20142_bfr_after (
		.din(new_net_20141),
		.dout(new_net_20142)
	);

	bfr new_net_20143_bfr_after (
		.din(new_net_20142),
		.dout(new_net_20143)
	);

	bfr new_net_20144_bfr_after (
		.din(new_net_20143),
		.dout(new_net_20144)
	);

	bfr new_net_20145_bfr_after (
		.din(new_net_20144),
		.dout(new_net_20145)
	);

	bfr new_net_20146_bfr_after (
		.din(new_net_20145),
		.dout(new_net_20146)
	);

	bfr new_net_20147_bfr_after (
		.din(new_net_20146),
		.dout(new_net_20147)
	);

	bfr new_net_20148_bfr_after (
		.din(new_net_20147),
		.dout(new_net_20148)
	);

	bfr new_net_20149_bfr_after (
		.din(new_net_20148),
		.dout(new_net_20149)
	);

	bfr new_net_20150_bfr_after (
		.din(new_net_20149),
		.dout(new_net_20150)
	);

	bfr new_net_20151_bfr_after (
		.din(new_net_20150),
		.dout(new_net_20151)
	);

	bfr new_net_20152_bfr_after (
		.din(new_net_20151),
		.dout(new_net_20152)
	);

	bfr new_net_20153_bfr_after (
		.din(new_net_20152),
		.dout(new_net_20153)
	);

	bfr new_net_20154_bfr_after (
		.din(new_net_20153),
		.dout(new_net_20154)
	);

	bfr new_net_20155_bfr_after (
		.din(new_net_20154),
		.dout(new_net_20155)
	);

	bfr new_net_20156_bfr_after (
		.din(new_net_20155),
		.dout(new_net_20156)
	);

	bfr new_net_20157_bfr_after (
		.din(new_net_20156),
		.dout(new_net_20157)
	);

	bfr new_net_20158_bfr_after (
		.din(new_net_20157),
		.dout(new_net_20158)
	);

	bfr new_net_20159_bfr_after (
		.din(new_net_20158),
		.dout(new_net_20159)
	);

	bfr new_net_20160_bfr_after (
		.din(new_net_20159),
		.dout(new_net_20160)
	);

	bfr new_net_20161_bfr_after (
		.din(new_net_20160),
		.dout(new_net_20161)
	);

	bfr new_net_20162_bfr_after (
		.din(new_net_20161),
		.dout(new_net_20162)
	);

	bfr new_net_20163_bfr_after (
		.din(new_net_20162),
		.dout(new_net_20163)
	);

	bfr new_net_20164_bfr_after (
		.din(new_net_20163),
		.dout(new_net_20164)
	);

	bfr new_net_20165_bfr_after (
		.din(new_net_20164),
		.dout(new_net_20165)
	);

	bfr new_net_20166_bfr_after (
		.din(new_net_20165),
		.dout(new_net_20166)
	);

	bfr new_net_20167_bfr_after (
		.din(new_net_20166),
		.dout(new_net_20167)
	);

	bfr new_net_20168_bfr_after (
		.din(new_net_20167),
		.dout(new_net_20168)
	);

	bfr new_net_20169_bfr_after (
		.din(new_net_20168),
		.dout(new_net_20169)
	);

	bfr new_net_20170_bfr_after (
		.din(new_net_20169),
		.dout(new_net_20170)
	);

	bfr new_net_20171_bfr_after (
		.din(new_net_20170),
		.dout(new_net_20171)
	);

	bfr new_net_20172_bfr_after (
		.din(new_net_20171),
		.dout(new_net_20172)
	);

	bfr new_net_20173_bfr_after (
		.din(new_net_20172),
		.dout(new_net_20173)
	);

	bfr new_net_20174_bfr_after (
		.din(new_net_20173),
		.dout(new_net_20174)
	);

	bfr new_net_20175_bfr_after (
		.din(new_net_20174),
		.dout(new_net_20175)
	);

	bfr new_net_20176_bfr_after (
		.din(new_net_20175),
		.dout(new_net_20176)
	);

	bfr new_net_20177_bfr_after (
		.din(new_net_20176),
		.dout(new_net_20177)
	);

	bfr new_net_20178_bfr_after (
		.din(new_net_20177),
		.dout(new_net_20178)
	);

	bfr new_net_20179_bfr_after (
		.din(new_net_20178),
		.dout(new_net_20179)
	);

	bfr new_net_20180_bfr_after (
		.din(new_net_20179),
		.dout(new_net_20180)
	);

	bfr new_net_20181_bfr_after (
		.din(new_net_20180),
		.dout(new_net_20181)
	);

	bfr new_net_20182_bfr_after (
		.din(new_net_20181),
		.dout(new_net_20182)
	);

	bfr new_net_20183_bfr_after (
		.din(new_net_20182),
		.dout(new_net_20183)
	);

	bfr new_net_20184_bfr_after (
		.din(new_net_20183),
		.dout(new_net_20184)
	);

	bfr new_net_20185_bfr_after (
		.din(new_net_20184),
		.dout(new_net_20185)
	);

	bfr new_net_20186_bfr_after (
		.din(new_net_20185),
		.dout(new_net_20186)
	);

	bfr new_net_20187_bfr_after (
		.din(new_net_20186),
		.dout(new_net_20187)
	);

	bfr new_net_20188_bfr_after (
		.din(new_net_20187),
		.dout(new_net_20188)
	);

	bfr new_net_20189_bfr_after (
		.din(new_net_20188),
		.dout(new_net_20189)
	);

	bfr new_net_20190_bfr_after (
		.din(new_net_20189),
		.dout(new_net_20190)
	);

	bfr new_net_20191_bfr_after (
		.din(new_net_20190),
		.dout(new_net_20191)
	);

	bfr new_net_20192_bfr_after (
		.din(new_net_20191),
		.dout(new_net_20192)
	);

	bfr new_net_20193_bfr_after (
		.din(new_net_20192),
		.dout(new_net_20193)
	);

	bfr new_net_20194_bfr_after (
		.din(new_net_20193),
		.dout(new_net_20194)
	);

	bfr new_net_20195_bfr_after (
		.din(new_net_20194),
		.dout(new_net_20195)
	);

	bfr new_net_20196_bfr_after (
		.din(new_net_20195),
		.dout(new_net_20196)
	);

	bfr new_net_20197_bfr_after (
		.din(new_net_20196),
		.dout(new_net_20197)
	);

	bfr new_net_20198_bfr_after (
		.din(new_net_20197),
		.dout(new_net_20198)
	);

	bfr new_net_20199_bfr_after (
		.din(new_net_20198),
		.dout(new_net_20199)
	);

	bfr new_net_20200_bfr_after (
		.din(new_net_20199),
		.dout(new_net_20200)
	);

	bfr new_net_20201_bfr_after (
		.din(new_net_20200),
		.dout(new_net_20201)
	);

	bfr new_net_20202_bfr_after (
		.din(new_net_20201),
		.dout(new_net_20202)
	);

	bfr new_net_20203_bfr_after (
		.din(new_net_20202),
		.dout(new_net_20203)
	);

	bfr new_net_20204_bfr_after (
		.din(new_net_20203),
		.dout(new_net_20204)
	);

	bfr new_net_20205_bfr_after (
		.din(new_net_20204),
		.dout(new_net_20205)
	);

	bfr new_net_20206_bfr_after (
		.din(new_net_20205),
		.dout(new_net_20206)
	);

	bfr new_net_20207_bfr_after (
		.din(new_net_20206),
		.dout(new_net_20207)
	);

	bfr new_net_20208_bfr_after (
		.din(new_net_20207),
		.dout(new_net_20208)
	);

	bfr new_net_20209_bfr_after (
		.din(new_net_20208),
		.dout(new_net_20209)
	);

	bfr new_net_20210_bfr_after (
		.din(new_net_20209),
		.dout(new_net_20210)
	);

	bfr new_net_20211_bfr_after (
		.din(new_net_20210),
		.dout(new_net_20211)
	);

	bfr new_net_20212_bfr_after (
		.din(new_net_20211),
		.dout(new_net_20212)
	);

	bfr new_net_20213_bfr_after (
		.din(new_net_20212),
		.dout(new_net_20213)
	);

	bfr new_net_20214_bfr_after (
		.din(new_net_20213),
		.dout(new_net_20214)
	);

	bfr new_net_20215_bfr_after (
		.din(new_net_20214),
		.dout(new_net_20215)
	);

	bfr new_net_20216_bfr_after (
		.din(new_net_20215),
		.dout(new_net_20216)
	);

	bfr new_net_20217_bfr_after (
		.din(new_net_20216),
		.dout(new_net_20217)
	);

	bfr new_net_20218_bfr_after (
		.din(new_net_20217),
		.dout(new_net_20218)
	);

	bfr new_net_20219_bfr_after (
		.din(new_net_20218),
		.dout(new_net_20219)
	);

	bfr new_net_20220_bfr_after (
		.din(new_net_20219),
		.dout(new_net_20220)
	);

	bfr new_net_20221_bfr_after (
		.din(new_net_20220),
		.dout(new_net_20221)
	);

	bfr new_net_20222_bfr_after (
		.din(new_net_20221),
		.dout(new_net_20222)
	);

	bfr new_net_20223_bfr_after (
		.din(new_net_20222),
		.dout(new_net_20223)
	);

	bfr new_net_20224_bfr_after (
		.din(new_net_20223),
		.dout(new_net_20224)
	);

	bfr new_net_20225_bfr_after (
		.din(new_net_20224),
		.dout(new_net_20225)
	);

	bfr new_net_20226_bfr_after (
		.din(new_net_20225),
		.dout(new_net_20226)
	);

	bfr new_net_20227_bfr_after (
		.din(new_net_20226),
		.dout(new_net_20227)
	);

	bfr new_net_20228_bfr_after (
		.din(new_net_20227),
		.dout(new_net_20228)
	);

	bfr new_net_20229_bfr_after (
		.din(new_net_20228),
		.dout(new_net_20229)
	);

	bfr new_net_20230_bfr_after (
		.din(new_net_20229),
		.dout(new_net_20230)
	);

	bfr new_net_20231_bfr_after (
		.din(new_net_20230),
		.dout(new_net_20231)
	);

	bfr new_net_20232_bfr_after (
		.din(new_net_20231),
		.dout(new_net_20232)
	);

	bfr new_net_20233_bfr_after (
		.din(new_net_20232),
		.dout(new_net_20233)
	);

	bfr new_net_20234_bfr_after (
		.din(new_net_20233),
		.dout(new_net_20234)
	);

	bfr new_net_20235_bfr_after (
		.din(new_net_20234),
		.dout(new_net_20235)
	);

	bfr new_net_20236_bfr_after (
		.din(new_net_20235),
		.dout(new_net_20236)
	);

	bfr new_net_20237_bfr_after (
		.din(new_net_20236),
		.dout(new_net_20237)
	);

	bfr new_net_20238_bfr_after (
		.din(new_net_20237),
		.dout(new_net_20238)
	);

	bfr new_net_20239_bfr_after (
		.din(new_net_20238),
		.dout(new_net_20239)
	);

	bfr new_net_20240_bfr_after (
		.din(new_net_20239),
		.dout(new_net_20240)
	);

	bfr new_net_20241_bfr_after (
		.din(new_net_20240),
		.dout(new_net_20241)
	);

	bfr new_net_20242_bfr_after (
		.din(new_net_20241),
		.dout(new_net_20242)
	);

	bfr new_net_20243_bfr_after (
		.din(new_net_20242),
		.dout(new_net_20243)
	);

	bfr new_net_20244_bfr_after (
		.din(new_net_20243),
		.dout(new_net_20244)
	);

	bfr new_net_20245_bfr_after (
		.din(new_net_20244),
		.dout(new_net_20245)
	);

	bfr new_net_20246_bfr_after (
		.din(new_net_20245),
		.dout(new_net_20246)
	);

	bfr new_net_20247_bfr_after (
		.din(new_net_20246),
		.dout(new_net_20247)
	);

	bfr new_net_20248_bfr_after (
		.din(new_net_20247),
		.dout(new_net_20248)
	);

	bfr new_net_20249_bfr_after (
		.din(new_net_20248),
		.dout(new_net_20249)
	);

	bfr new_net_20250_bfr_after (
		.din(new_net_20249),
		.dout(new_net_20250)
	);

	bfr new_net_20251_bfr_after (
		.din(new_net_20250),
		.dout(new_net_20251)
	);

	bfr new_net_20252_bfr_after (
		.din(new_net_20251),
		.dout(new_net_20252)
	);

	bfr new_net_20253_bfr_after (
		.din(new_net_20252),
		.dout(new_net_20253)
	);

	bfr new_net_20254_bfr_after (
		.din(new_net_20253),
		.dout(new_net_20254)
	);

	bfr new_net_20255_bfr_after (
		.din(new_net_20254),
		.dout(new_net_20255)
	);

	bfr new_net_20256_bfr_after (
		.din(new_net_20255),
		.dout(new_net_20256)
	);

	bfr new_net_20257_bfr_after (
		.din(new_net_20256),
		.dout(new_net_20257)
	);

	bfr new_net_20258_bfr_after (
		.din(new_net_20257),
		.dout(new_net_20258)
	);

	bfr new_net_20259_bfr_after (
		.din(new_net_20258),
		.dout(new_net_20259)
	);

	bfr new_net_20260_bfr_after (
		.din(new_net_20259),
		.dout(new_net_20260)
	);

	bfr new_net_20261_bfr_after (
		.din(new_net_20260),
		.dout(new_net_20261)
	);

	bfr new_net_20262_bfr_after (
		.din(new_net_20261),
		.dout(new_net_20262)
	);

	bfr new_net_20263_bfr_after (
		.din(new_net_20262),
		.dout(new_net_20263)
	);

	bfr new_net_20264_bfr_after (
		.din(new_net_20263),
		.dout(new_net_20264)
	);

	bfr new_net_20265_bfr_after (
		.din(new_net_20264),
		.dout(new_net_20265)
	);

	bfr new_net_20266_bfr_after (
		.din(new_net_20265),
		.dout(new_net_20266)
	);

	bfr new_net_20267_bfr_after (
		.din(new_net_20266),
		.dout(new_net_20267)
	);

	bfr new_net_20268_bfr_after (
		.din(new_net_20267),
		.dout(new_net_20268)
	);

	bfr new_net_20269_bfr_after (
		.din(new_net_20268),
		.dout(new_net_20269)
	);

	bfr new_net_20270_bfr_after (
		.din(new_net_20269),
		.dout(new_net_20270)
	);

	bfr new_net_20271_bfr_after (
		.din(new_net_20270),
		.dout(new_net_20271)
	);

	bfr new_net_20272_bfr_after (
		.din(new_net_20271),
		.dout(new_net_20272)
	);

	bfr new_net_20273_bfr_after (
		.din(new_net_20272),
		.dout(new_net_20273)
	);

	bfr new_net_20274_bfr_after (
		.din(new_net_20273),
		.dout(new_net_20274)
	);

	bfr new_net_20275_bfr_after (
		.din(new_net_20274),
		.dout(new_net_20275)
	);

	bfr new_net_20276_bfr_after (
		.din(new_net_20275),
		.dout(new_net_20276)
	);

	bfr new_net_20277_bfr_after (
		.din(new_net_20276),
		.dout(new_net_20277)
	);

	bfr new_net_20278_bfr_after (
		.din(new_net_20277),
		.dout(new_net_20278)
	);

	bfr new_net_20279_bfr_after (
		.din(new_net_20278),
		.dout(new_net_20279)
	);

	bfr new_net_20280_bfr_after (
		.din(new_net_20279),
		.dout(new_net_20280)
	);

	bfr new_net_20281_bfr_after (
		.din(new_net_20280),
		.dout(new_net_20281)
	);

	bfr new_net_20282_bfr_after (
		.din(new_net_20281),
		.dout(new_net_20282)
	);

	bfr new_net_20283_bfr_after (
		.din(new_net_20282),
		.dout(new_net_20283)
	);

	bfr new_net_20284_bfr_after (
		.din(new_net_20283),
		.dout(new_net_20284)
	);

	bfr new_net_20285_bfr_after (
		.din(new_net_20284),
		.dout(new_net_20285)
	);

	bfr new_net_20286_bfr_after (
		.din(new_net_20285),
		.dout(new_net_20286)
	);

	bfr new_net_20287_bfr_after (
		.din(new_net_20286),
		.dout(new_net_20287)
	);

	bfr new_net_20288_bfr_after (
		.din(new_net_20287),
		.dout(new_net_20288)
	);

	bfr new_net_20289_bfr_after (
		.din(new_net_20288),
		.dout(new_net_20289)
	);

	bfr new_net_20290_bfr_after (
		.din(new_net_20289),
		.dout(new_net_20290)
	);

	bfr new_net_20291_bfr_after (
		.din(new_net_20290),
		.dout(new_net_20291)
	);

	bfr new_net_20292_bfr_after (
		.din(new_net_20291),
		.dout(new_net_20292)
	);

	bfr new_net_20293_bfr_after (
		.din(new_net_20292),
		.dout(new_net_20293)
	);

	bfr new_net_20294_bfr_after (
		.din(new_net_20293),
		.dout(new_net_20294)
	);

	bfr new_net_20295_bfr_after (
		.din(new_net_20294),
		.dout(new_net_20295)
	);

	bfr new_net_20296_bfr_after (
		.din(new_net_20295),
		.dout(new_net_20296)
	);

	bfr new_net_20297_bfr_after (
		.din(new_net_20296),
		.dout(new_net_20297)
	);

	bfr new_net_20298_bfr_after (
		.din(new_net_20297),
		.dout(new_net_20298)
	);

	bfr N1901_bfr_after (
		.din(new_net_20298),
		.dout(N1901)
	);

	bfr new_net_3700_bfr_after (
		.din(_0062_),
		.dout(new_net_3700)
	);

	bfr new_net_3733_bfr_after (
		.din(_0204_),
		.dout(new_net_3733)
	);

	bfr new_net_3872_bfr_after (
		.din(_0819_),
		.dout(new_net_3872)
	);

	bfr new_net_3899_bfr_after (
		.din(_0941_),
		.dout(new_net_3899)
	);

	bfr new_net_3473_bfr_after (
		.din(_0546_),
		.dout(new_net_3473)
	);

	bfr new_net_3565_bfr_after (
		.din(_1327_),
		.dout(new_net_3565)
	);

	bfr new_net_3575_bfr_after (
		.din(_1357_),
		.dout(new_net_3575)
	);

	bfr new_net_3695_bfr_after (
		.din(_0046_),
		.dout(new_net_3695)
	);

	bfr new_net_3829_bfr_after (
		.din(_0643_),
		.dout(new_net_3829)
	);

	bfr new_net_3905_bfr_after (
		.din(_0967_),
		.dout(new_net_3905)
	);

	bfr new_net_20299_bfr_after (
		.din(new_net_3940),
		.dout(new_net_20299)
	);

	bfr new_net_20300_bfr_after (
		.din(new_net_20299),
		.dout(new_net_20300)
	);

	bfr new_net_20301_bfr_after (
		.din(new_net_20300),
		.dout(new_net_20301)
	);

	bfr new_net_20302_bfr_after (
		.din(new_net_20301),
		.dout(new_net_20302)
	);

	bfr new_net_20303_bfr_after (
		.din(new_net_20302),
		.dout(new_net_20303)
	);

	bfr new_net_20304_bfr_after (
		.din(new_net_20303),
		.dout(new_net_20304)
	);

	bfr new_net_20305_bfr_after (
		.din(new_net_20304),
		.dout(new_net_20305)
	);

	bfr new_net_20306_bfr_after (
		.din(new_net_20305),
		.dout(new_net_20306)
	);

	bfr new_net_20307_bfr_after (
		.din(new_net_20306),
		.dout(new_net_20307)
	);

	bfr new_net_20308_bfr_after (
		.din(new_net_20307),
		.dout(new_net_20308)
	);

	bfr new_net_20309_bfr_after (
		.din(new_net_20308),
		.dout(new_net_20309)
	);

	bfr new_net_20310_bfr_after (
		.din(new_net_20309),
		.dout(new_net_20310)
	);

	bfr new_net_20311_bfr_after (
		.din(new_net_20310),
		.dout(new_net_20311)
	);

	bfr new_net_20312_bfr_after (
		.din(new_net_20311),
		.dout(new_net_20312)
	);

	bfr new_net_20313_bfr_after (
		.din(new_net_20312),
		.dout(new_net_20313)
	);

	bfr new_net_20314_bfr_after (
		.din(new_net_20313),
		.dout(new_net_20314)
	);

	bfr new_net_20315_bfr_after (
		.din(new_net_20314),
		.dout(new_net_20315)
	);

	bfr new_net_20316_bfr_after (
		.din(new_net_20315),
		.dout(new_net_20316)
	);

	bfr new_net_20317_bfr_after (
		.din(new_net_20316),
		.dout(new_net_20317)
	);

	bfr new_net_20318_bfr_after (
		.din(new_net_20317),
		.dout(new_net_20318)
	);

	bfr new_net_20319_bfr_after (
		.din(new_net_20318),
		.dout(new_net_20319)
	);

	bfr new_net_20320_bfr_after (
		.din(new_net_20319),
		.dout(new_net_20320)
	);

	bfr new_net_20321_bfr_after (
		.din(new_net_20320),
		.dout(new_net_20321)
	);

	bfr new_net_20322_bfr_after (
		.din(new_net_20321),
		.dout(new_net_20322)
	);

	bfr new_net_20323_bfr_after (
		.din(new_net_20322),
		.dout(new_net_20323)
	);

	bfr new_net_20324_bfr_after (
		.din(new_net_20323),
		.dout(new_net_20324)
	);

	bfr new_net_20325_bfr_after (
		.din(new_net_20324),
		.dout(new_net_20325)
	);

	bfr new_net_20326_bfr_after (
		.din(new_net_20325),
		.dout(new_net_20326)
	);

	bfr new_net_20327_bfr_after (
		.din(new_net_20326),
		.dout(new_net_20327)
	);

	bfr new_net_20328_bfr_after (
		.din(new_net_20327),
		.dout(new_net_20328)
	);

	bfr new_net_20329_bfr_after (
		.din(new_net_20328),
		.dout(new_net_20329)
	);

	bfr new_net_20330_bfr_after (
		.din(new_net_20329),
		.dout(new_net_20330)
	);

	bfr new_net_20331_bfr_after (
		.din(new_net_20330),
		.dout(new_net_20331)
	);

	bfr new_net_20332_bfr_after (
		.din(new_net_20331),
		.dout(new_net_20332)
	);

	bfr new_net_20333_bfr_after (
		.din(new_net_20332),
		.dout(new_net_20333)
	);

	bfr new_net_20334_bfr_after (
		.din(new_net_20333),
		.dout(new_net_20334)
	);

	bfr new_net_20335_bfr_after (
		.din(new_net_20334),
		.dout(new_net_20335)
	);

	bfr new_net_20336_bfr_after (
		.din(new_net_20335),
		.dout(new_net_20336)
	);

	bfr new_net_20337_bfr_after (
		.din(new_net_20336),
		.dout(new_net_20337)
	);

	bfr new_net_20338_bfr_after (
		.din(new_net_20337),
		.dout(new_net_20338)
	);

	bfr new_net_20339_bfr_after (
		.din(new_net_20338),
		.dout(new_net_20339)
	);

	bfr new_net_20340_bfr_after (
		.din(new_net_20339),
		.dout(new_net_20340)
	);

	bfr new_net_20341_bfr_after (
		.din(new_net_20340),
		.dout(new_net_20341)
	);

	bfr new_net_20342_bfr_after (
		.din(new_net_20341),
		.dout(new_net_20342)
	);

	bfr new_net_20343_bfr_after (
		.din(new_net_20342),
		.dout(new_net_20343)
	);

	bfr new_net_20344_bfr_after (
		.din(new_net_20343),
		.dout(new_net_20344)
	);

	bfr new_net_20345_bfr_after (
		.din(new_net_20344),
		.dout(new_net_20345)
	);

	bfr new_net_20346_bfr_after (
		.din(new_net_20345),
		.dout(new_net_20346)
	);

	bfr new_net_20347_bfr_after (
		.din(new_net_20346),
		.dout(new_net_20347)
	);

	bfr new_net_20348_bfr_after (
		.din(new_net_20347),
		.dout(new_net_20348)
	);

	bfr new_net_20349_bfr_after (
		.din(new_net_20348),
		.dout(new_net_20349)
	);

	bfr new_net_20350_bfr_after (
		.din(new_net_20349),
		.dout(new_net_20350)
	);

	bfr new_net_20351_bfr_after (
		.din(new_net_20350),
		.dout(new_net_20351)
	);

	bfr new_net_20352_bfr_after (
		.din(new_net_20351),
		.dout(new_net_20352)
	);

	bfr new_net_20353_bfr_after (
		.din(new_net_20352),
		.dout(new_net_20353)
	);

	bfr N6150_bfr_after (
		.din(new_net_20353),
		.dout(N6150)
	);

	bfr new_net_20354_bfr_after (
		.din(new_net_3972),
		.dout(new_net_20354)
	);

	bfr new_net_20355_bfr_after (
		.din(new_net_20354),
		.dout(new_net_20355)
	);

	bfr new_net_20356_bfr_after (
		.din(new_net_20355),
		.dout(new_net_20356)
	);

	bfr new_net_20357_bfr_after (
		.din(new_net_20356),
		.dout(new_net_20357)
	);

	bfr new_net_20358_bfr_after (
		.din(new_net_20357),
		.dout(new_net_20358)
	);

	bfr new_net_20359_bfr_after (
		.din(new_net_20358),
		.dout(new_net_20359)
	);

	bfr new_net_20360_bfr_after (
		.din(new_net_20359),
		.dout(new_net_20360)
	);

	bfr N6270_bfr_after (
		.din(new_net_20360),
		.dout(N6270)
	);

	bfr new_net_3484_bfr_after (
		.din(_1014_),
		.dout(new_net_3484)
	);

	bfr new_net_3587_bfr_after (
		.din(_1415_),
		.dout(new_net_3587)
	);

	bfr new_net_3658_bfr_after (
		.din(_1733_),
		.dout(new_net_3658)
	);

	bfr new_net_3854_bfr_after (
		.din(_0744_),
		.dout(new_net_3854)
	);

	bfr new_net_3870_bfr_after (
		.din(_0812_),
		.dout(new_net_3870)
	);

	bfr new_net_3906_bfr_after (
		.din(_0971_),
		.dout(new_net_3906)
	);

	bfr new_net_3503_bfr_after (
		.din(_1101_),
		.dout(new_net_3503)
	);

	bfr new_net_3569_bfr_after (
		.din(_1339_),
		.dout(new_net_3569)
	);

	bfr new_net_3654_bfr_after (
		.din(_1720_),
		.dout(new_net_3654)
	);

	bfr new_net_3702_bfr_after (
		.din(_0069_),
		.dout(new_net_3702)
	);

	bfr new_net_3762_bfr_after (
		.din(_0356_),
		.dout(new_net_3762)
	);

	bfr new_net_3773_bfr_after (
		.din(_0392_),
		.dout(new_net_3773)
	);

	bfr new_net_3783_bfr_after (
		.din(_0425_),
		.dout(new_net_3783)
	);

	bfr new_net_20361_bfr_after (
		.din(new_net_3966),
		.dout(new_net_20361)
	);

	bfr new_net_20362_bfr_after (
		.din(new_net_20361),
		.dout(new_net_20362)
	);

	bfr new_net_20363_bfr_after (
		.din(new_net_20362),
		.dout(new_net_20363)
	);

	bfr new_net_20364_bfr_after (
		.din(new_net_20363),
		.dout(new_net_20364)
	);

	bfr new_net_20365_bfr_after (
		.din(new_net_20364),
		.dout(new_net_20365)
	);

	bfr new_net_20366_bfr_after (
		.din(new_net_20365),
		.dout(new_net_20366)
	);

	bfr new_net_20367_bfr_after (
		.din(new_net_20366),
		.dout(new_net_20367)
	);

	bfr new_net_20368_bfr_after (
		.din(new_net_20367),
		.dout(new_net_20368)
	);

	bfr new_net_20369_bfr_after (
		.din(new_net_20368),
		.dout(new_net_20369)
	);

	bfr new_net_20370_bfr_after (
		.din(new_net_20369),
		.dout(new_net_20370)
	);

	bfr new_net_20371_bfr_after (
		.din(new_net_20370),
		.dout(new_net_20371)
	);

	bfr new_net_20372_bfr_after (
		.din(new_net_20371),
		.dout(new_net_20372)
	);

	bfr new_net_20373_bfr_after (
		.din(new_net_20372),
		.dout(new_net_20373)
	);

	bfr new_net_20374_bfr_after (
		.din(new_net_20373),
		.dout(new_net_20374)
	);

	bfr new_net_20375_bfr_after (
		.din(new_net_20374),
		.dout(new_net_20375)
	);

	bfr new_net_20376_bfr_after (
		.din(new_net_20375),
		.dout(new_net_20376)
	);

	bfr new_net_20377_bfr_after (
		.din(new_net_20376),
		.dout(new_net_20377)
	);

	bfr new_net_20378_bfr_after (
		.din(new_net_20377),
		.dout(new_net_20378)
	);

	bfr new_net_20379_bfr_after (
		.din(new_net_20378),
		.dout(new_net_20379)
	);

	bfr new_net_20380_bfr_after (
		.din(new_net_20379),
		.dout(new_net_20380)
	);

	bfr new_net_20381_bfr_after (
		.din(new_net_20380),
		.dout(new_net_20381)
	);

	bfr new_net_20382_bfr_after (
		.din(new_net_20381),
		.dout(new_net_20382)
	);

	bfr new_net_20383_bfr_after (
		.din(new_net_20382),
		.dout(new_net_20383)
	);

	bfr new_net_20384_bfr_after (
		.din(new_net_20383),
		.dout(new_net_20384)
	);

	bfr new_net_20385_bfr_after (
		.din(new_net_20384),
		.dout(new_net_20385)
	);

	bfr new_net_20386_bfr_after (
		.din(new_net_20385),
		.dout(new_net_20386)
	);

	bfr new_net_20387_bfr_after (
		.din(new_net_20386),
		.dout(new_net_20387)
	);

	bfr new_net_20388_bfr_after (
		.din(new_net_20387),
		.dout(new_net_20388)
	);

	bfr new_net_20389_bfr_after (
		.din(new_net_20388),
		.dout(new_net_20389)
	);

	bfr new_net_20390_bfr_after (
		.din(new_net_20389),
		.dout(new_net_20390)
	);

	bfr new_net_20391_bfr_after (
		.din(new_net_20390),
		.dout(new_net_20391)
	);

	bfr new_net_20392_bfr_after (
		.din(new_net_20391),
		.dout(new_net_20392)
	);

	bfr new_net_20393_bfr_after (
		.din(new_net_20392),
		.dout(new_net_20393)
	);

	bfr new_net_20394_bfr_after (
		.din(new_net_20393),
		.dout(new_net_20394)
	);

	bfr new_net_20395_bfr_after (
		.din(new_net_20394),
		.dout(new_net_20395)
	);

	bfr N6200_bfr_after (
		.din(new_net_20395),
		.dout(N6200)
	);

	bfr new_net_3465_bfr_after (
		.din(_0176_),
		.dout(new_net_3465)
	);

	bfr new_net_3644_bfr_after (
		.din(_1653_),
		.dout(new_net_3644)
	);

	bfr new_net_3759_bfr_after (
		.din(_0320_),
		.dout(new_net_3759)
	);

	bfr new_net_3803_bfr_after (
		.din(_0516_),
		.dout(new_net_3803)
	);

	bfr new_net_3867_bfr_after (
		.din(_0802_),
		.dout(new_net_3867)
	);

	bfr new_net_3882_bfr_after (
		.din(_0865_),
		.dout(new_net_3882)
	);

	bfr new_net_3610_bfr_after (
		.din(_1514_),
		.dout(new_net_3610)
	);

	bfr new_net_3671_bfr_after (
		.din(_1776_),
		.dout(new_net_3671)
	);

	bfr new_net_3685_bfr_after (
		.din(_0013_),
		.dout(new_net_3685)
	);

	bfr new_net_3737_bfr_after (
		.din(_0247_),
		.dout(new_net_3737)
	);

	bfr new_net_3844_bfr_after (
		.din(_0693_),
		.dout(new_net_3844)
	);

	bfr new_net_3864_bfr_after (
		.din(_0792_),
		.dout(new_net_3864)
	);

	bfr new_net_3896_bfr_after (
		.din(_0922_),
		.dout(new_net_3896)
	);

	bfr new_net_20396_bfr_after (
		.din(new_net_3936),
		.dout(new_net_20396)
	);

	bfr new_net_20397_bfr_after (
		.din(new_net_20396),
		.dout(new_net_20397)
	);

	bfr new_net_20398_bfr_after (
		.din(new_net_20397),
		.dout(new_net_20398)
	);

	bfr new_net_20399_bfr_after (
		.din(new_net_20398),
		.dout(new_net_20399)
	);

	bfr new_net_20400_bfr_after (
		.din(new_net_20399),
		.dout(new_net_20400)
	);

	bfr new_net_20401_bfr_after (
		.din(new_net_20400),
		.dout(new_net_20401)
	);

	bfr new_net_20402_bfr_after (
		.din(new_net_20401),
		.dout(new_net_20402)
	);

	bfr new_net_20403_bfr_after (
		.din(new_net_20402),
		.dout(new_net_20403)
	);

	bfr new_net_20404_bfr_after (
		.din(new_net_20403),
		.dout(new_net_20404)
	);

	bfr new_net_20405_bfr_after (
		.din(new_net_20404),
		.dout(new_net_20405)
	);

	bfr new_net_20406_bfr_after (
		.din(new_net_20405),
		.dout(new_net_20406)
	);

	bfr new_net_20407_bfr_after (
		.din(new_net_20406),
		.dout(new_net_20407)
	);

	bfr new_net_20408_bfr_after (
		.din(new_net_20407),
		.dout(new_net_20408)
	);

	bfr new_net_20409_bfr_after (
		.din(new_net_20408),
		.dout(new_net_20409)
	);

	bfr new_net_20410_bfr_after (
		.din(new_net_20409),
		.dout(new_net_20410)
	);

	bfr new_net_20411_bfr_after (
		.din(new_net_20410),
		.dout(new_net_20411)
	);

	bfr new_net_20412_bfr_after (
		.din(new_net_20411),
		.dout(new_net_20412)
	);

	bfr new_net_20413_bfr_after (
		.din(new_net_20412),
		.dout(new_net_20413)
	);

	bfr new_net_20414_bfr_after (
		.din(new_net_20413),
		.dout(new_net_20414)
	);

	bfr new_net_20415_bfr_after (
		.din(new_net_20414),
		.dout(new_net_20415)
	);

	bfr new_net_20416_bfr_after (
		.din(new_net_20415),
		.dout(new_net_20416)
	);

	bfr new_net_20417_bfr_after (
		.din(new_net_20416),
		.dout(new_net_20417)
	);

	bfr new_net_20418_bfr_after (
		.din(new_net_20417),
		.dout(new_net_20418)
	);

	bfr new_net_20419_bfr_after (
		.din(new_net_20418),
		.dout(new_net_20419)
	);

	bfr new_net_20420_bfr_after (
		.din(new_net_20419),
		.dout(new_net_20420)
	);

	bfr new_net_20421_bfr_after (
		.din(new_net_20420),
		.dout(new_net_20421)
	);

	bfr new_net_20422_bfr_after (
		.din(new_net_20421),
		.dout(new_net_20422)
	);

	bfr new_net_20423_bfr_after (
		.din(new_net_20422),
		.dout(new_net_20423)
	);

	bfr new_net_20424_bfr_after (
		.din(new_net_20423),
		.dout(new_net_20424)
	);

	bfr new_net_20425_bfr_after (
		.din(new_net_20424),
		.dout(new_net_20425)
	);

	bfr new_net_20426_bfr_after (
		.din(new_net_20425),
		.dout(new_net_20426)
	);

	bfr new_net_20427_bfr_after (
		.din(new_net_20426),
		.dout(new_net_20427)
	);

	bfr new_net_20428_bfr_after (
		.din(new_net_20427),
		.dout(new_net_20428)
	);

	bfr new_net_20429_bfr_after (
		.din(new_net_20428),
		.dout(new_net_20429)
	);

	bfr new_net_20430_bfr_after (
		.din(new_net_20429),
		.dout(new_net_20430)
	);

	bfr new_net_20431_bfr_after (
		.din(new_net_20430),
		.dout(new_net_20431)
	);

	bfr new_net_20432_bfr_after (
		.din(new_net_20431),
		.dout(new_net_20432)
	);

	bfr new_net_20433_bfr_after (
		.din(new_net_20432),
		.dout(new_net_20433)
	);

	bfr new_net_20434_bfr_after (
		.din(new_net_20433),
		.dout(new_net_20434)
	);

	bfr new_net_20435_bfr_after (
		.din(new_net_20434),
		.dout(new_net_20435)
	);

	bfr new_net_20436_bfr_after (
		.din(new_net_20435),
		.dout(new_net_20436)
	);

	bfr new_net_20437_bfr_after (
		.din(new_net_20436),
		.dout(new_net_20437)
	);

	bfr new_net_20438_bfr_after (
		.din(new_net_20437),
		.dout(new_net_20438)
	);

	bfr new_net_20439_bfr_after (
		.din(new_net_20438),
		.dout(new_net_20439)
	);

	bfr new_net_20440_bfr_after (
		.din(new_net_20439),
		.dout(new_net_20440)
	);

	bfr new_net_20441_bfr_after (
		.din(new_net_20440),
		.dout(new_net_20441)
	);

	bfr new_net_20442_bfr_after (
		.din(new_net_20441),
		.dout(new_net_20442)
	);

	bfr new_net_20443_bfr_after (
		.din(new_net_20442),
		.dout(new_net_20443)
	);

	bfr new_net_20444_bfr_after (
		.din(new_net_20443),
		.dout(new_net_20444)
	);

	bfr new_net_20445_bfr_after (
		.din(new_net_20444),
		.dout(new_net_20445)
	);

	bfr new_net_20446_bfr_after (
		.din(new_net_20445),
		.dout(new_net_20446)
	);

	bfr N6160_bfr_after (
		.din(new_net_20446),
		.dout(N6160)
	);

	bfr new_net_3511_bfr_after (
		.din(_1126_),
		.dout(new_net_3511)
	);

	bfr new_net_3532_bfr_after (
		.din(_1198_),
		.dout(new_net_3532)
	);

	bfr new_net_3550_bfr_after (
		.din(_1262_),
		.dout(new_net_3550)
	);

	bfr new_net_3559_bfr_after (
		.din(_1309_),
		.dout(new_net_3559)
	);

	bfr new_net_3573_bfr_after (
		.din(_1351_),
		.dout(new_net_3573)
	);

	bfr new_net_3626_bfr_after (
		.din(_1594_),
		.dout(new_net_3626)
	);

	bfr new_net_3832_bfr_after (
		.din(_0653_),
		.dout(new_net_3832)
	);

	bfr new_net_3530_bfr_after (
		.din(_1196_),
		.dout(new_net_3530)
	);

	bfr new_net_3495_bfr_after (
		.din(_1061_),
		.dout(new_net_3495)
	);

	bfr new_net_3583_bfr_after (
		.din(_1403_),
		.dout(new_net_3583)
	);

	bfr new_net_3792_bfr_after (
		.din(_0479_),
		.dout(new_net_3792)
	);

	bfr new_net_3845_bfr_after (
		.din(_0714_),
		.dout(new_net_3845)
	);

	bfr new_net_3883_bfr_after (
		.din(_0868_),
		.dout(new_net_3883)
	);

	bfr new_net_3599_bfr_after (
		.din(_1451_),
		.dout(new_net_3599)
	);

	bfr new_net_3617_bfr_after (
		.din(_1537_),
		.dout(new_net_3617)
	);

	bfr new_net_3659_bfr_after (
		.din(_1736_),
		.dout(new_net_3659)
	);

	bfr new_net_3672_bfr_after (
		.din(_1779_),
		.dout(new_net_3672)
	);

	bfr new_net_3711_bfr_after (
		.din(_0131_),
		.dout(new_net_3711)
	);

	bfr new_net_3889_bfr_after (
		.din(_0899_),
		.dout(new_net_3889)
	);

	bfr new_net_3730_bfr_after (
		.din(_0194_),
		.dout(new_net_3730)
	);

	bfr new_net_3468_bfr_after (
		.din(_0383_),
		.dout(new_net_3468)
	);

	bfr new_net_3560_bfr_after (
		.din(_1312_),
		.dout(new_net_3560)
	);

	bfr new_net_3582_bfr_after (
		.din(_1400_),
		.dout(new_net_3582)
	);

	bfr new_net_3675_bfr_after (
		.din(_1789_),
		.dout(new_net_3675)
	);

	bfr new_net_3887_bfr_after (
		.din(_0892_),
		.dout(new_net_3887)
	);

	bfr new_net_3748_bfr_after (
		.din(_0283_),
		.dout(new_net_3748)
	);

	bfr new_net_3528_bfr_after (
		.din(_1194_),
		.dout(new_net_3528)
	);

	bfr new_net_3474_bfr_after (
		.din(_0579_),
		.dout(new_net_3474)
	);

	bfr new_net_3479_bfr_after (
		.din(_0872_),
		.dout(new_net_3479)
	);

	bfr new_net_3639_bfr_after (
		.din(_1637_),
		.dout(new_net_3639)
	);

	bfr new_net_3655_bfr_after (
		.din(_1723_),
		.dout(new_net_3655)
	);

	bfr new_net_3736_bfr_after (
		.din(_0244_),
		.dout(new_net_3736)
	);

	bfr new_net_3768_bfr_after (
		.din(_0376_),
		.dout(new_net_3768)
	);

	bfr new_net_3807_bfr_after (
		.din(_0551_),
		.dout(new_net_3807)
	);

	bfr new_net_3817_bfr_after (
		.din(_0584_),
		.dout(new_net_3817)
	);

	bfr new_net_3548_bfr_after (
		.din(_1256_),
		.dout(new_net_3548)
	);

	bfr new_net_3662_bfr_after (
		.din(_1746_),
		.dout(new_net_3662)
	);

	bfr new_net_20447_bfr_after (
		.din(new_net_3952),
		.dout(new_net_20447)
	);

	bfr new_net_20448_bfr_after (
		.din(new_net_20447),
		.dout(new_net_20448)
	);

	bfr new_net_20449_bfr_after (
		.din(new_net_20448),
		.dout(new_net_20449)
	);

	bfr new_net_20450_bfr_after (
		.din(new_net_20449),
		.dout(new_net_20450)
	);

	bfr new_net_20451_bfr_after (
		.din(new_net_20450),
		.dout(new_net_20451)
	);

	bfr new_net_20452_bfr_after (
		.din(new_net_20451),
		.dout(new_net_20452)
	);

	bfr new_net_20453_bfr_after (
		.din(new_net_20452),
		.dout(new_net_20453)
	);

	bfr new_net_20454_bfr_after (
		.din(new_net_20453),
		.dout(new_net_20454)
	);

	bfr new_net_20455_bfr_after (
		.din(new_net_20454),
		.dout(new_net_20455)
	);

	bfr new_net_20456_bfr_after (
		.din(new_net_20455),
		.dout(new_net_20456)
	);

	bfr new_net_20457_bfr_after (
		.din(new_net_20456),
		.dout(new_net_20457)
	);

	bfr new_net_20458_bfr_after (
		.din(new_net_20457),
		.dout(new_net_20458)
	);

	bfr new_net_20459_bfr_after (
		.din(new_net_20458),
		.dout(new_net_20459)
	);

	bfr new_net_20460_bfr_after (
		.din(new_net_20459),
		.dout(new_net_20460)
	);

	bfr new_net_20461_bfr_after (
		.din(new_net_20460),
		.dout(new_net_20461)
	);

	bfr new_net_20462_bfr_after (
		.din(new_net_20461),
		.dout(new_net_20462)
	);

	bfr new_net_20463_bfr_after (
		.din(new_net_20462),
		.dout(new_net_20463)
	);

	bfr new_net_20464_bfr_after (
		.din(new_net_20463),
		.dout(new_net_20464)
	);

	bfr new_net_20465_bfr_after (
		.din(new_net_20464),
		.dout(new_net_20465)
	);

	bfr new_net_20466_bfr_after (
		.din(new_net_20465),
		.dout(new_net_20466)
	);

	bfr new_net_20467_bfr_after (
		.din(new_net_20466),
		.dout(new_net_20467)
	);

	bfr new_net_20468_bfr_after (
		.din(new_net_20467),
		.dout(new_net_20468)
	);

	bfr new_net_20469_bfr_after (
		.din(new_net_20468),
		.dout(new_net_20469)
	);

	bfr new_net_20470_bfr_after (
		.din(new_net_20469),
		.dout(new_net_20470)
	);

	bfr new_net_20471_bfr_after (
		.din(new_net_20470),
		.dout(new_net_20471)
	);

	bfr new_net_20472_bfr_after (
		.din(new_net_20471),
		.dout(new_net_20472)
	);

	bfr new_net_20473_bfr_after (
		.din(new_net_20472),
		.dout(new_net_20473)
	);

	bfr new_net_20474_bfr_after (
		.din(new_net_20473),
		.dout(new_net_20474)
	);

	bfr new_net_20475_bfr_after (
		.din(new_net_20474),
		.dout(new_net_20475)
	);

	bfr new_net_20476_bfr_after (
		.din(new_net_20475),
		.dout(new_net_20476)
	);

	bfr new_net_20477_bfr_after (
		.din(new_net_20476),
		.dout(new_net_20477)
	);

	bfr new_net_20478_bfr_after (
		.din(new_net_20477),
		.dout(new_net_20478)
	);

	bfr new_net_20479_bfr_after (
		.din(new_net_20478),
		.dout(new_net_20479)
	);

	bfr new_net_20480_bfr_after (
		.din(new_net_20479),
		.dout(new_net_20480)
	);

	bfr new_net_20481_bfr_after (
		.din(new_net_20480),
		.dout(new_net_20481)
	);

	bfr new_net_20482_bfr_after (
		.din(new_net_20481),
		.dout(new_net_20482)
	);

	bfr new_net_20483_bfr_after (
		.din(new_net_20482),
		.dout(new_net_20483)
	);

	bfr new_net_20484_bfr_after (
		.din(new_net_20483),
		.dout(new_net_20484)
	);

	bfr new_net_20485_bfr_after (
		.din(new_net_20484),
		.dout(new_net_20485)
	);

	bfr new_net_20486_bfr_after (
		.din(new_net_20485),
		.dout(new_net_20486)
	);

	bfr new_net_20487_bfr_after (
		.din(new_net_20486),
		.dout(new_net_20487)
	);

	bfr new_net_20488_bfr_after (
		.din(new_net_20487),
		.dout(new_net_20488)
	);

	bfr new_net_20489_bfr_after (
		.din(new_net_20488),
		.dout(new_net_20489)
	);

	bfr new_net_20490_bfr_after (
		.din(new_net_20489),
		.dout(new_net_20490)
	);

	bfr new_net_20491_bfr_after (
		.din(new_net_20490),
		.dout(new_net_20491)
	);

	bfr new_net_20492_bfr_after (
		.din(new_net_20491),
		.dout(new_net_20492)
	);

	bfr new_net_20493_bfr_after (
		.din(new_net_20492),
		.dout(new_net_20493)
	);

	bfr new_net_20494_bfr_after (
		.din(new_net_20493),
		.dout(new_net_20494)
	);

	bfr new_net_20495_bfr_after (
		.din(new_net_20494),
		.dout(new_net_20495)
	);

	bfr new_net_20496_bfr_after (
		.din(new_net_20495),
		.dout(new_net_20496)
	);

	bfr new_net_20497_bfr_after (
		.din(new_net_20496),
		.dout(new_net_20497)
	);

	bfr new_net_20498_bfr_after (
		.din(new_net_20497),
		.dout(new_net_20498)
	);

	bfr new_net_20499_bfr_after (
		.din(new_net_20498),
		.dout(new_net_20499)
	);

	bfr new_net_20500_bfr_after (
		.din(new_net_20499),
		.dout(new_net_20500)
	);

	bfr new_net_20501_bfr_after (
		.din(new_net_20500),
		.dout(new_net_20501)
	);

	bfr new_net_20502_bfr_after (
		.din(new_net_20501),
		.dout(new_net_20502)
	);

	bfr new_net_20503_bfr_after (
		.din(new_net_20502),
		.dout(new_net_20503)
	);

	bfr new_net_20504_bfr_after (
		.din(new_net_20503),
		.dout(new_net_20504)
	);

	bfr new_net_20505_bfr_after (
		.din(new_net_20504),
		.dout(new_net_20505)
	);

	bfr new_net_20506_bfr_after (
		.din(new_net_20505),
		.dout(new_net_20506)
	);

	bfr new_net_20507_bfr_after (
		.din(new_net_20506),
		.dout(new_net_20507)
	);

	bfr new_net_20508_bfr_after (
		.din(new_net_20507),
		.dout(new_net_20508)
	);

	bfr new_net_20509_bfr_after (
		.din(new_net_20508),
		.dout(new_net_20509)
	);

	bfr new_net_20510_bfr_after (
		.din(new_net_20509),
		.dout(new_net_20510)
	);

	bfr new_net_20511_bfr_after (
		.din(new_net_20510),
		.dout(new_net_20511)
	);

	bfr new_net_20512_bfr_after (
		.din(new_net_20511),
		.dout(new_net_20512)
	);

	bfr new_net_20513_bfr_after (
		.din(new_net_20512),
		.dout(new_net_20513)
	);

	bfr new_net_20514_bfr_after (
		.din(new_net_20513),
		.dout(new_net_20514)
	);

	bfr new_net_20515_bfr_after (
		.din(new_net_20514),
		.dout(new_net_20515)
	);

	bfr new_net_20516_bfr_after (
		.din(new_net_20515),
		.dout(new_net_20516)
	);

	bfr new_net_20517_bfr_after (
		.din(new_net_20516),
		.dout(new_net_20517)
	);

	bfr new_net_20518_bfr_after (
		.din(new_net_20517),
		.dout(new_net_20518)
	);

	bfr new_net_20519_bfr_after (
		.din(new_net_20518),
		.dout(new_net_20519)
	);

	bfr new_net_20520_bfr_after (
		.din(new_net_20519),
		.dout(new_net_20520)
	);

	bfr new_net_20521_bfr_after (
		.din(new_net_20520),
		.dout(new_net_20521)
	);

	bfr new_net_20522_bfr_after (
		.din(new_net_20521),
		.dout(new_net_20522)
	);

	bfr new_net_20523_bfr_after (
		.din(new_net_20522),
		.dout(new_net_20523)
	);

	bfr new_net_20524_bfr_after (
		.din(new_net_20523),
		.dout(new_net_20524)
	);

	bfr new_net_20525_bfr_after (
		.din(new_net_20524),
		.dout(new_net_20525)
	);

	bfr new_net_20526_bfr_after (
		.din(new_net_20525),
		.dout(new_net_20526)
	);

	bfr new_net_20527_bfr_after (
		.din(new_net_20526),
		.dout(new_net_20527)
	);

	bfr new_net_20528_bfr_after (
		.din(new_net_20527),
		.dout(new_net_20528)
	);

	bfr new_net_20529_bfr_after (
		.din(new_net_20528),
		.dout(new_net_20529)
	);

	bfr N5308_bfr_after (
		.din(new_net_20529),
		.dout(N5308)
	);

	bfr new_net_3477_bfr_after (
		.din(_0807_),
		.dout(new_net_3477)
	);

	bfr new_net_3493_bfr_after (
		.din(_1055_),
		.dout(new_net_3493)
	);

	bfr new_net_3538_bfr_after (
		.din(_1226_),
		.dout(new_net_3538)
	);

	bfr new_net_3838_bfr_after (
		.din(_0673_),
		.dout(new_net_3838)
	);

	bfr new_net_3908_bfr_after (
		.din(_0977_),
		.dout(new_net_3908)
	);

	bfr new_net_3738_bfr_after (
		.din(_0250_),
		.dout(new_net_3738)
	);

	bfr new_net_3631_bfr_after (
		.din(_1611_),
		.dout(new_net_3631)
	);

	bfr new_net_3509_bfr_after (
		.din(_1119_),
		.dout(new_net_3509)
	);

	bfr new_net_3552_bfr_after (
		.din(_1268_),
		.dout(new_net_3552)
	);

	bfr new_net_3563_bfr_after (
		.din(_1321_),
		.dout(new_net_3563)
	);

	bfr new_net_3590_bfr_after (
		.din(_1424_),
		.dout(new_net_3590)
	);

	bfr new_net_3660_bfr_after (
		.din(_1739_),
		.dout(new_net_3660)
	);

	bfr new_net_3708_bfr_after (
		.din(_0122_),
		.dout(new_net_3708)
	);

	bfr new_net_3814_bfr_after (
		.din(_0574_),
		.dout(new_net_3814)
	);

	bfr new_net_3463_bfr_after (
		.din(_0110_),
		.dout(new_net_3463)
	);

	bfr new_net_3490_bfr_after (
		.din(_1046_),
		.dout(new_net_3490)
	);

	bfr new_net_3512_bfr_after (
		.din(_1146_),
		.dout(new_net_3512)
	);

	bfr new_net_3713_bfr_after (
		.din(_0138_),
		.dout(new_net_3713)
	);

	bfr new_net_3802_bfr_after (
		.din(_0512_),
		.dout(new_net_3802)
	);

	bfr new_net_3819_bfr_after (
		.din(_0591_),
		.dout(new_net_3819)
	);

	bfr new_net_3691_bfr_after (
		.din(_0032_),
		.dout(new_net_3691)
	);

	bfr new_net_3524_bfr_after (
		.din(_1182_),
		.dout(new_net_3524)
	);

	bfr new_net_3535_bfr_after (
		.din(_1201_),
		.dout(new_net_3535)
	);

	bfr new_net_3562_bfr_after (
		.din(_1318_),
		.dout(new_net_3562)
	);

	bfr new_net_3597_bfr_after (
		.din(_1445_),
		.dout(new_net_3597)
	);

	bfr new_net_3627_bfr_after (
		.din(_1597_),
		.dout(new_net_3627)
	);

	bfr new_net_3846_bfr_after (
		.din(_0717_),
		.dout(new_net_3846)
	);

	bfr new_net_3865_bfr_after (
		.din(_0795_),
		.dout(new_net_3865)
	);

	bfr new_net_3886_bfr_after (
		.din(_0878_),
		.dout(new_net_3886)
	);

	bfr new_net_3893_bfr_after (
		.din(_0912_),
		.dout(new_net_3893)
	);

	bfr new_net_3521_bfr_after (
		.din(_1173_),
		.dout(new_net_3521)
	);

	bfr new_net_3556_bfr_after (
		.din(_1300_),
		.dout(new_net_3556)
	);

	bfr new_net_3653_bfr_after (
		.din(_1716_),
		.dout(new_net_3653)
	);

	bfr new_net_3801_bfr_after (
		.din(_0509_),
		.dout(new_net_3801)
	);

	bfr new_net_20530_bfr_after (
		.din(new_net_3926),
		.dout(new_net_20530)
	);

	bfr new_net_20531_bfr_after (
		.din(new_net_20530),
		.dout(new_net_20531)
	);

	bfr new_net_20532_bfr_after (
		.din(new_net_20531),
		.dout(new_net_20532)
	);

	bfr new_net_20533_bfr_after (
		.din(new_net_20532),
		.dout(new_net_20533)
	);

	bfr new_net_20534_bfr_after (
		.din(new_net_20533),
		.dout(new_net_20534)
	);

	bfr new_net_20535_bfr_after (
		.din(new_net_20534),
		.dout(new_net_20535)
	);

	bfr new_net_20536_bfr_after (
		.din(new_net_20535),
		.dout(new_net_20536)
	);

	bfr new_net_20537_bfr_after (
		.din(new_net_20536),
		.dout(new_net_20537)
	);

	bfr new_net_20538_bfr_after (
		.din(new_net_20537),
		.dout(new_net_20538)
	);

	bfr new_net_20539_bfr_after (
		.din(new_net_20538),
		.dout(new_net_20539)
	);

	bfr new_net_20540_bfr_after (
		.din(new_net_20539),
		.dout(new_net_20540)
	);

	bfr new_net_20541_bfr_after (
		.din(new_net_20540),
		.dout(new_net_20541)
	);

	bfr new_net_20542_bfr_after (
		.din(new_net_20541),
		.dout(new_net_20542)
	);

	bfr new_net_20543_bfr_after (
		.din(new_net_20542),
		.dout(new_net_20543)
	);

	bfr new_net_20544_bfr_after (
		.din(new_net_20543),
		.dout(new_net_20544)
	);

	bfr new_net_20545_bfr_after (
		.din(new_net_20544),
		.dout(new_net_20545)
	);

	bfr new_net_20546_bfr_after (
		.din(new_net_20545),
		.dout(new_net_20546)
	);

	bfr new_net_20547_bfr_after (
		.din(new_net_20546),
		.dout(new_net_20547)
	);

	bfr new_net_20548_bfr_after (
		.din(new_net_20547),
		.dout(new_net_20548)
	);

	bfr new_net_20549_bfr_after (
		.din(new_net_20548),
		.dout(new_net_20549)
	);

	bfr new_net_20550_bfr_after (
		.din(new_net_20549),
		.dout(new_net_20550)
	);

	bfr new_net_20551_bfr_after (
		.din(new_net_20550),
		.dout(new_net_20551)
	);

	bfr new_net_20552_bfr_after (
		.din(new_net_20551),
		.dout(new_net_20552)
	);

	bfr new_net_20553_bfr_after (
		.din(new_net_20552),
		.dout(new_net_20553)
	);

	bfr new_net_20554_bfr_after (
		.din(new_net_20553),
		.dout(new_net_20554)
	);

	bfr new_net_20555_bfr_after (
		.din(new_net_20554),
		.dout(new_net_20555)
	);

	bfr new_net_20556_bfr_after (
		.din(new_net_20555),
		.dout(new_net_20556)
	);

	bfr new_net_20557_bfr_after (
		.din(new_net_20556),
		.dout(new_net_20557)
	);

	bfr new_net_20558_bfr_after (
		.din(new_net_20557),
		.dout(new_net_20558)
	);

	bfr new_net_20559_bfr_after (
		.din(new_net_20558),
		.dout(new_net_20559)
	);

	bfr new_net_20560_bfr_after (
		.din(new_net_20559),
		.dout(new_net_20560)
	);

	bfr new_net_20561_bfr_after (
		.din(new_net_20560),
		.dout(new_net_20561)
	);

	bfr new_net_20562_bfr_after (
		.din(new_net_20561),
		.dout(new_net_20562)
	);

	bfr new_net_20563_bfr_after (
		.din(new_net_20562),
		.dout(new_net_20563)
	);

	bfr new_net_20564_bfr_after (
		.din(new_net_20563),
		.dout(new_net_20564)
	);

	bfr new_net_20565_bfr_after (
		.din(new_net_20564),
		.dout(new_net_20565)
	);

	bfr new_net_20566_bfr_after (
		.din(new_net_20565),
		.dout(new_net_20566)
	);

	bfr new_net_20567_bfr_after (
		.din(new_net_20566),
		.dout(new_net_20567)
	);

	bfr new_net_20568_bfr_after (
		.din(new_net_20567),
		.dout(new_net_20568)
	);

	bfr new_net_20569_bfr_after (
		.din(new_net_20568),
		.dout(new_net_20569)
	);

	bfr new_net_20570_bfr_after (
		.din(new_net_20569),
		.dout(new_net_20570)
	);

	bfr new_net_20571_bfr_after (
		.din(new_net_20570),
		.dout(new_net_20571)
	);

	bfr new_net_20572_bfr_after (
		.din(new_net_20571),
		.dout(new_net_20572)
	);

	bfr new_net_20573_bfr_after (
		.din(new_net_20572),
		.dout(new_net_20573)
	);

	bfr new_net_20574_bfr_after (
		.din(new_net_20573),
		.dout(new_net_20574)
	);

	bfr new_net_20575_bfr_after (
		.din(new_net_20574),
		.dout(new_net_20575)
	);

	bfr new_net_20576_bfr_after (
		.din(new_net_20575),
		.dout(new_net_20576)
	);

	bfr new_net_20577_bfr_after (
		.din(new_net_20576),
		.dout(new_net_20577)
	);

	bfr new_net_20578_bfr_after (
		.din(new_net_20577),
		.dout(new_net_20578)
	);

	bfr new_net_20579_bfr_after (
		.din(new_net_20578),
		.dout(new_net_20579)
	);

	bfr new_net_20580_bfr_after (
		.din(new_net_20579),
		.dout(new_net_20580)
	);

	bfr new_net_20581_bfr_after (
		.din(new_net_20580),
		.dout(new_net_20581)
	);

	bfr new_net_20582_bfr_after (
		.din(new_net_20581),
		.dout(new_net_20582)
	);

	bfr new_net_20583_bfr_after (
		.din(new_net_20582),
		.dout(new_net_20583)
	);

	bfr new_net_20584_bfr_after (
		.din(new_net_20583),
		.dout(new_net_20584)
	);

	bfr new_net_20585_bfr_after (
		.din(new_net_20584),
		.dout(new_net_20585)
	);

	bfr new_net_20586_bfr_after (
		.din(new_net_20585),
		.dout(new_net_20586)
	);

	bfr new_net_20587_bfr_after (
		.din(new_net_20586),
		.dout(new_net_20587)
	);

	bfr new_net_20588_bfr_after (
		.din(new_net_20587),
		.dout(new_net_20588)
	);

	bfr new_net_20589_bfr_after (
		.din(new_net_20588),
		.dout(new_net_20589)
	);

	bfr new_net_20590_bfr_after (
		.din(new_net_20589),
		.dout(new_net_20590)
	);

	bfr new_net_20591_bfr_after (
		.din(new_net_20590),
		.dout(new_net_20591)
	);

	bfr new_net_20592_bfr_after (
		.din(new_net_20591),
		.dout(new_net_20592)
	);

	bfr new_net_20593_bfr_after (
		.din(new_net_20592),
		.dout(new_net_20593)
	);

	bfr new_net_20594_bfr_after (
		.din(new_net_20593),
		.dout(new_net_20594)
	);

	bfr new_net_20595_bfr_after (
		.din(new_net_20594),
		.dout(new_net_20595)
	);

	bfr new_net_20596_bfr_after (
		.din(new_net_20595),
		.dout(new_net_20596)
	);

	bfr new_net_20597_bfr_after (
		.din(new_net_20596),
		.dout(new_net_20597)
	);

	bfr new_net_20598_bfr_after (
		.din(new_net_20597),
		.dout(new_net_20598)
	);

	bfr new_net_20599_bfr_after (
		.din(new_net_20598),
		.dout(new_net_20599)
	);

	bfr new_net_20600_bfr_after (
		.din(new_net_20599),
		.dout(new_net_20600)
	);

	bfr new_net_20601_bfr_after (
		.din(new_net_20600),
		.dout(new_net_20601)
	);

	bfr new_net_20602_bfr_after (
		.din(new_net_20601),
		.dout(new_net_20602)
	);

	bfr new_net_20603_bfr_after (
		.din(new_net_20602),
		.dout(new_net_20603)
	);

	bfr new_net_20604_bfr_after (
		.din(new_net_20603),
		.dout(new_net_20604)
	);

	bfr new_net_20605_bfr_after (
		.din(new_net_20604),
		.dout(new_net_20605)
	);

	bfr new_net_20606_bfr_after (
		.din(new_net_20605),
		.dout(new_net_20606)
	);

	bfr new_net_20607_bfr_after (
		.din(new_net_20606),
		.dout(new_net_20607)
	);

	bfr new_net_20608_bfr_after (
		.din(new_net_20607),
		.dout(new_net_20608)
	);

	bfr new_net_20609_bfr_after (
		.din(new_net_20608),
		.dout(new_net_20609)
	);

	bfr new_net_20610_bfr_after (
		.din(new_net_20609),
		.dout(new_net_20610)
	);

	bfr new_net_20611_bfr_after (
		.din(new_net_20610),
		.dout(new_net_20611)
	);

	bfr new_net_20612_bfr_after (
		.din(new_net_20611),
		.dout(new_net_20612)
	);

	bfr new_net_20613_bfr_after (
		.din(new_net_20612),
		.dout(new_net_20613)
	);

	bfr new_net_20614_bfr_after (
		.din(new_net_20613),
		.dout(new_net_20614)
	);

	bfr new_net_20615_bfr_after (
		.din(new_net_20614),
		.dout(new_net_20615)
	);

	bfr new_net_20616_bfr_after (
		.din(new_net_20615),
		.dout(new_net_20616)
	);

	bfr new_net_20617_bfr_after (
		.din(new_net_20616),
		.dout(new_net_20617)
	);

	bfr new_net_20618_bfr_after (
		.din(new_net_20617),
		.dout(new_net_20618)
	);

	bfr new_net_20619_bfr_after (
		.din(new_net_20618),
		.dout(new_net_20619)
	);

	bfr new_net_20620_bfr_after (
		.din(new_net_20619),
		.dout(new_net_20620)
	);

	bfr N4946_bfr_after (
		.din(new_net_20620),
		.dout(N4946)
	);

	bfr new_net_20621_bfr_after (
		.din(new_net_3968),
		.dout(new_net_20621)
	);

	bfr new_net_20622_bfr_after (
		.din(new_net_20621),
		.dout(new_net_20622)
	);

	bfr new_net_20623_bfr_after (
		.din(new_net_20622),
		.dout(new_net_20623)
	);

	bfr new_net_20624_bfr_after (
		.din(new_net_20623),
		.dout(new_net_20624)
	);

	bfr new_net_20625_bfr_after (
		.din(new_net_20624),
		.dout(new_net_20625)
	);

	bfr new_net_20626_bfr_after (
		.din(new_net_20625),
		.dout(new_net_20626)
	);

	bfr new_net_20627_bfr_after (
		.din(new_net_20626),
		.dout(new_net_20627)
	);

	bfr new_net_20628_bfr_after (
		.din(new_net_20627),
		.dout(new_net_20628)
	);

	bfr new_net_20629_bfr_after (
		.din(new_net_20628),
		.dout(new_net_20629)
	);

	bfr new_net_20630_bfr_after (
		.din(new_net_20629),
		.dout(new_net_20630)
	);

	bfr new_net_20631_bfr_after (
		.din(new_net_20630),
		.dout(new_net_20631)
	);

	bfr new_net_20632_bfr_after (
		.din(new_net_20631),
		.dout(new_net_20632)
	);

	bfr new_net_20633_bfr_after (
		.din(new_net_20632),
		.dout(new_net_20633)
	);

	bfr new_net_20634_bfr_after (
		.din(new_net_20633),
		.dout(new_net_20634)
	);

	bfr new_net_20635_bfr_after (
		.din(new_net_20634),
		.dout(new_net_20635)
	);

	bfr new_net_20636_bfr_after (
		.din(new_net_20635),
		.dout(new_net_20636)
	);

	bfr new_net_20637_bfr_after (
		.din(new_net_20636),
		.dout(new_net_20637)
	);

	bfr new_net_20638_bfr_after (
		.din(new_net_20637),
		.dout(new_net_20638)
	);

	bfr new_net_20639_bfr_after (
		.din(new_net_20638),
		.dout(new_net_20639)
	);

	bfr new_net_20640_bfr_after (
		.din(new_net_20639),
		.dout(new_net_20640)
	);

	bfr new_net_20641_bfr_after (
		.din(new_net_20640),
		.dout(new_net_20641)
	);

	bfr new_net_20642_bfr_after (
		.din(new_net_20641),
		.dout(new_net_20642)
	);

	bfr new_net_20643_bfr_after (
		.din(new_net_20642),
		.dout(new_net_20643)
	);

	bfr new_net_20644_bfr_after (
		.din(new_net_20643),
		.dout(new_net_20644)
	);

	bfr new_net_20645_bfr_after (
		.din(new_net_20644),
		.dout(new_net_20645)
	);

	bfr new_net_20646_bfr_after (
		.din(new_net_20645),
		.dout(new_net_20646)
	);

	bfr new_net_20647_bfr_after (
		.din(new_net_20646),
		.dout(new_net_20647)
	);

	bfr new_net_20648_bfr_after (
		.din(new_net_20647),
		.dout(new_net_20648)
	);

	bfr new_net_20649_bfr_after (
		.din(new_net_20648),
		.dout(new_net_20649)
	);

	bfr new_net_20650_bfr_after (
		.din(new_net_20649),
		.dout(new_net_20650)
	);

	bfr new_net_20651_bfr_after (
		.din(new_net_20650),
		.dout(new_net_20651)
	);

	bfr new_net_20652_bfr_after (
		.din(new_net_20651),
		.dout(new_net_20652)
	);

	bfr new_net_20653_bfr_after (
		.din(new_net_20652),
		.dout(new_net_20653)
	);

	bfr new_net_20654_bfr_after (
		.din(new_net_20653),
		.dout(new_net_20654)
	);

	bfr new_net_20655_bfr_after (
		.din(new_net_20654),
		.dout(new_net_20655)
	);

	bfr new_net_20656_bfr_after (
		.din(new_net_20655),
		.dout(new_net_20656)
	);

	bfr new_net_20657_bfr_after (
		.din(new_net_20656),
		.dout(new_net_20657)
	);

	bfr new_net_20658_bfr_after (
		.din(new_net_20657),
		.dout(new_net_20658)
	);

	bfr new_net_20659_bfr_after (
		.din(new_net_20658),
		.dout(new_net_20659)
	);

	bfr new_net_20660_bfr_after (
		.din(new_net_20659),
		.dout(new_net_20660)
	);

	bfr new_net_20661_bfr_after (
		.din(new_net_20660),
		.dout(new_net_20661)
	);

	bfr new_net_20662_bfr_after (
		.din(new_net_20661),
		.dout(new_net_20662)
	);

	bfr new_net_20663_bfr_after (
		.din(new_net_20662),
		.dout(new_net_20663)
	);

	bfr new_net_20664_bfr_after (
		.din(new_net_20663),
		.dout(new_net_20664)
	);

	bfr new_net_20665_bfr_after (
		.din(new_net_20664),
		.dout(new_net_20665)
	);

	bfr new_net_20666_bfr_after (
		.din(new_net_20665),
		.dout(new_net_20666)
	);

	bfr new_net_20667_bfr_after (
		.din(new_net_20666),
		.dout(new_net_20667)
	);

	bfr new_net_20668_bfr_after (
		.din(new_net_20667),
		.dout(new_net_20668)
	);

	bfr new_net_20669_bfr_after (
		.din(new_net_20668),
		.dout(new_net_20669)
	);

	bfr new_net_20670_bfr_after (
		.din(new_net_20669),
		.dout(new_net_20670)
	);

	bfr new_net_20671_bfr_after (
		.din(new_net_20670),
		.dout(new_net_20671)
	);

	bfr new_net_20672_bfr_after (
		.din(new_net_20671),
		.dout(new_net_20672)
	);

	bfr new_net_20673_bfr_after (
		.din(new_net_20672),
		.dout(new_net_20673)
	);

	bfr new_net_20674_bfr_after (
		.din(new_net_20673),
		.dout(new_net_20674)
	);

	bfr new_net_20675_bfr_after (
		.din(new_net_20674),
		.dout(new_net_20675)
	);

	bfr new_net_20676_bfr_after (
		.din(new_net_20675),
		.dout(new_net_20676)
	);

	bfr new_net_20677_bfr_after (
		.din(new_net_20676),
		.dout(new_net_20677)
	);

	bfr new_net_20678_bfr_after (
		.din(new_net_20677),
		.dout(new_net_20678)
	);

	bfr new_net_20679_bfr_after (
		.din(new_net_20678),
		.dout(new_net_20679)
	);

	bfr new_net_20680_bfr_after (
		.din(new_net_20679),
		.dout(new_net_20680)
	);

	bfr new_net_20681_bfr_after (
		.din(new_net_20680),
		.dout(new_net_20681)
	);

	bfr new_net_20682_bfr_after (
		.din(new_net_20681),
		.dout(new_net_20682)
	);

	bfr new_net_20683_bfr_after (
		.din(new_net_20682),
		.dout(new_net_20683)
	);

	bfr new_net_20684_bfr_after (
		.din(new_net_20683),
		.dout(new_net_20684)
	);

	bfr new_net_20685_bfr_after (
		.din(new_net_20684),
		.dout(new_net_20685)
	);

	bfr new_net_20686_bfr_after (
		.din(new_net_20685),
		.dout(new_net_20686)
	);

	bfr new_net_20687_bfr_after (
		.din(new_net_20686),
		.dout(new_net_20687)
	);

	bfr new_net_20688_bfr_after (
		.din(new_net_20687),
		.dout(new_net_20688)
	);

	bfr new_net_20689_bfr_after (
		.din(new_net_20688),
		.dout(new_net_20689)
	);

	bfr new_net_20690_bfr_after (
		.din(new_net_20689),
		.dout(new_net_20690)
	);

	bfr new_net_20691_bfr_after (
		.din(new_net_20690),
		.dout(new_net_20691)
	);

	bfr new_net_20692_bfr_after (
		.din(new_net_20691),
		.dout(new_net_20692)
	);

	bfr new_net_20693_bfr_after (
		.din(new_net_20692),
		.dout(new_net_20693)
	);

	bfr new_net_20694_bfr_after (
		.din(new_net_20693),
		.dout(new_net_20694)
	);

	bfr new_net_20695_bfr_after (
		.din(new_net_20694),
		.dout(new_net_20695)
	);

	bfr new_net_20696_bfr_after (
		.din(new_net_20695),
		.dout(new_net_20696)
	);

	bfr new_net_20697_bfr_after (
		.din(new_net_20696),
		.dout(new_net_20697)
	);

	bfr new_net_20698_bfr_after (
		.din(new_net_20697),
		.dout(new_net_20698)
	);

	bfr new_net_20699_bfr_after (
		.din(new_net_20698),
		.dout(new_net_20699)
	);

	bfr new_net_20700_bfr_after (
		.din(new_net_20699),
		.dout(new_net_20700)
	);

	bfr new_net_20701_bfr_after (
		.din(new_net_20700),
		.dout(new_net_20701)
	);

	bfr new_net_20702_bfr_after (
		.din(new_net_20701),
		.dout(new_net_20702)
	);

	bfr new_net_20703_bfr_after (
		.din(new_net_20702),
		.dout(new_net_20703)
	);

	bfr new_net_20704_bfr_after (
		.din(new_net_20703),
		.dout(new_net_20704)
	);

	bfr new_net_20705_bfr_after (
		.din(new_net_20704),
		.dout(new_net_20705)
	);

	bfr new_net_20706_bfr_after (
		.din(new_net_20705),
		.dout(new_net_20706)
	);

	bfr new_net_20707_bfr_after (
		.din(new_net_20706),
		.dout(new_net_20707)
	);

	bfr new_net_20708_bfr_after (
		.din(new_net_20707),
		.dout(new_net_20708)
	);

	bfr new_net_20709_bfr_after (
		.din(new_net_20708),
		.dout(new_net_20709)
	);

	bfr new_net_20710_bfr_after (
		.din(new_net_20709),
		.dout(new_net_20710)
	);

	bfr new_net_20711_bfr_after (
		.din(new_net_20710),
		.dout(new_net_20711)
	);

	bfr new_net_20712_bfr_after (
		.din(new_net_20711),
		.dout(new_net_20712)
	);

	bfr new_net_20713_bfr_after (
		.din(new_net_20712),
		.dout(new_net_20713)
	);

	bfr new_net_20714_bfr_after (
		.din(new_net_20713),
		.dout(new_net_20714)
	);

	bfr new_net_20715_bfr_after (
		.din(new_net_20714),
		.dout(new_net_20715)
	);

	bfr new_net_20716_bfr_after (
		.din(new_net_20715),
		.dout(new_net_20716)
	);

	bfr new_net_20717_bfr_after (
		.din(new_net_20716),
		.dout(new_net_20717)
	);

	bfr new_net_20718_bfr_after (
		.din(new_net_20717),
		.dout(new_net_20718)
	);

	bfr new_net_20719_bfr_after (
		.din(new_net_20718),
		.dout(new_net_20719)
	);

	bfr new_net_20720_bfr_after (
		.din(new_net_20719),
		.dout(new_net_20720)
	);

	bfr new_net_20721_bfr_after (
		.din(new_net_20720),
		.dout(new_net_20721)
	);

	bfr new_net_20722_bfr_after (
		.din(new_net_20721),
		.dout(new_net_20722)
	);

	bfr new_net_20723_bfr_after (
		.din(new_net_20722),
		.dout(new_net_20723)
	);

	bfr new_net_20724_bfr_after (
		.din(new_net_20723),
		.dout(new_net_20724)
	);

	bfr new_net_20725_bfr_after (
		.din(new_net_20724),
		.dout(new_net_20725)
	);

	bfr new_net_20726_bfr_after (
		.din(new_net_20725),
		.dout(new_net_20726)
	);

	bfr new_net_20727_bfr_after (
		.din(new_net_20726),
		.dout(new_net_20727)
	);

	bfr new_net_20728_bfr_after (
		.din(new_net_20727),
		.dout(new_net_20728)
	);

	bfr new_net_20729_bfr_after (
		.din(new_net_20728),
		.dout(new_net_20729)
	);

	bfr new_net_20730_bfr_after (
		.din(new_net_20729),
		.dout(new_net_20730)
	);

	bfr new_net_20731_bfr_after (
		.din(new_net_20730),
		.dout(new_net_20731)
	);

	bfr new_net_20732_bfr_after (
		.din(new_net_20731),
		.dout(new_net_20732)
	);

	bfr new_net_20733_bfr_after (
		.din(new_net_20732),
		.dout(new_net_20733)
	);

	bfr new_net_20734_bfr_after (
		.din(new_net_20733),
		.dout(new_net_20734)
	);

	bfr new_net_20735_bfr_after (
		.din(new_net_20734),
		.dout(new_net_20735)
	);

	bfr new_net_20736_bfr_after (
		.din(new_net_20735),
		.dout(new_net_20736)
	);

	bfr new_net_20737_bfr_after (
		.din(new_net_20736),
		.dout(new_net_20737)
	);

	bfr new_net_20738_bfr_after (
		.din(new_net_20737),
		.dout(new_net_20738)
	);

	bfr new_net_20739_bfr_after (
		.din(new_net_20738),
		.dout(new_net_20739)
	);

	bfr new_net_20740_bfr_after (
		.din(new_net_20739),
		.dout(new_net_20740)
	);

	bfr new_net_20741_bfr_after (
		.din(new_net_20740),
		.dout(new_net_20741)
	);

	bfr new_net_20742_bfr_after (
		.din(new_net_20741),
		.dout(new_net_20742)
	);

	bfr new_net_20743_bfr_after (
		.din(new_net_20742),
		.dout(new_net_20743)
	);

	bfr new_net_20744_bfr_after (
		.din(new_net_20743),
		.dout(new_net_20744)
	);

	bfr new_net_20745_bfr_after (
		.din(new_net_20744),
		.dout(new_net_20745)
	);

	bfr new_net_20746_bfr_after (
		.din(new_net_20745),
		.dout(new_net_20746)
	);

	bfr new_net_20747_bfr_after (
		.din(new_net_20746),
		.dout(new_net_20747)
	);

	bfr new_net_20748_bfr_after (
		.din(new_net_20747),
		.dout(new_net_20748)
	);

	bfr new_net_20749_bfr_after (
		.din(new_net_20748),
		.dout(new_net_20749)
	);

	bfr new_net_20750_bfr_after (
		.din(new_net_20749),
		.dout(new_net_20750)
	);

	bfr new_net_20751_bfr_after (
		.din(new_net_20750),
		.dout(new_net_20751)
	);

	bfr new_net_20752_bfr_after (
		.din(new_net_20751),
		.dout(new_net_20752)
	);

	bfr new_net_20753_bfr_after (
		.din(new_net_20752),
		.dout(new_net_20753)
	);

	bfr new_net_20754_bfr_after (
		.din(new_net_20753),
		.dout(new_net_20754)
	);

	bfr new_net_20755_bfr_after (
		.din(new_net_20754),
		.dout(new_net_20755)
	);

	bfr new_net_20756_bfr_after (
		.din(new_net_20755),
		.dout(new_net_20756)
	);

	bfr new_net_20757_bfr_after (
		.din(new_net_20756),
		.dout(new_net_20757)
	);

	bfr new_net_20758_bfr_after (
		.din(new_net_20757),
		.dout(new_net_20758)
	);

	bfr new_net_20759_bfr_after (
		.din(new_net_20758),
		.dout(new_net_20759)
	);

	bfr new_net_20760_bfr_after (
		.din(new_net_20759),
		.dout(new_net_20760)
	);

	bfr new_net_20761_bfr_after (
		.din(new_net_20760),
		.dout(new_net_20761)
	);

	bfr new_net_20762_bfr_after (
		.din(new_net_20761),
		.dout(new_net_20762)
	);

	bfr new_net_20763_bfr_after (
		.din(new_net_20762),
		.dout(new_net_20763)
	);

	bfr new_net_20764_bfr_after (
		.din(new_net_20763),
		.dout(new_net_20764)
	);

	bfr new_net_20765_bfr_after (
		.din(new_net_20764),
		.dout(new_net_20765)
	);

	bfr new_net_20766_bfr_after (
		.din(new_net_20765),
		.dout(new_net_20766)
	);

	bfr new_net_20767_bfr_after (
		.din(new_net_20766),
		.dout(new_net_20767)
	);

	bfr new_net_20768_bfr_after (
		.din(new_net_20767),
		.dout(new_net_20768)
	);

	bfr new_net_20769_bfr_after (
		.din(new_net_20768),
		.dout(new_net_20769)
	);

	bfr new_net_20770_bfr_after (
		.din(new_net_20769),
		.dout(new_net_20770)
	);

	bfr new_net_20771_bfr_after (
		.din(new_net_20770),
		.dout(new_net_20771)
	);

	bfr new_net_20772_bfr_after (
		.din(new_net_20771),
		.dout(new_net_20772)
	);

	bfr new_net_20773_bfr_after (
		.din(new_net_20772),
		.dout(new_net_20773)
	);

	bfr new_net_20774_bfr_after (
		.din(new_net_20773),
		.dout(new_net_20774)
	);

	bfr new_net_20775_bfr_after (
		.din(new_net_20774),
		.dout(new_net_20775)
	);

	bfr N2223_bfr_after (
		.din(new_net_20775),
		.dout(N2223)
	);

	bfr new_net_3492_bfr_after (
		.din(_1052_),
		.dout(new_net_3492)
	);

	bfr new_net_3537_bfr_after (
		.din(_1223_),
		.dout(new_net_3537)
	);

	bfr new_net_3605_bfr_after (
		.din(_1497_),
		.dout(new_net_3605)
	);

	bfr new_net_3630_bfr_after (
		.din(_1607_),
		.dout(new_net_3630)
	);

	bfr new_net_3657_bfr_after (
		.din(_1729_),
		.dout(new_net_3657)
	);

	bfr new_net_3810_bfr_after (
		.din(_0561_),
		.dout(new_net_3810)
	);

	bfr new_net_20776_bfr_after (
		.din(new_net_3924),
		.dout(new_net_20776)
	);

	bfr new_net_20777_bfr_after (
		.din(new_net_20776),
		.dout(new_net_20777)
	);

	bfr new_net_20778_bfr_after (
		.din(new_net_20777),
		.dout(new_net_20778)
	);

	bfr new_net_20779_bfr_after (
		.din(new_net_20778),
		.dout(new_net_20779)
	);

	bfr new_net_20780_bfr_after (
		.din(new_net_20779),
		.dout(new_net_20780)
	);

	bfr new_net_20781_bfr_after (
		.din(new_net_20780),
		.dout(new_net_20781)
	);

	bfr new_net_20782_bfr_after (
		.din(new_net_20781),
		.dout(new_net_20782)
	);

	bfr new_net_20783_bfr_after (
		.din(new_net_20782),
		.dout(new_net_20783)
	);

	bfr new_net_20784_bfr_after (
		.din(new_net_20783),
		.dout(new_net_20784)
	);

	bfr new_net_20785_bfr_after (
		.din(new_net_20784),
		.dout(new_net_20785)
	);

	bfr new_net_20786_bfr_after (
		.din(new_net_20785),
		.dout(new_net_20786)
	);

	bfr new_net_20787_bfr_after (
		.din(new_net_20786),
		.dout(new_net_20787)
	);

	bfr new_net_20788_bfr_after (
		.din(new_net_20787),
		.dout(new_net_20788)
	);

	bfr new_net_20789_bfr_after (
		.din(new_net_20788),
		.dout(new_net_20789)
	);

	bfr new_net_20790_bfr_after (
		.din(new_net_20789),
		.dout(new_net_20790)
	);

	bfr N6250_bfr_after (
		.din(new_net_20790),
		.dout(N6250)
	);

	bfr new_net_3642_bfr_after (
		.din(_1647_),
		.dout(new_net_3642)
	);

	bfr new_net_3903_bfr_after (
		.din(_0954_),
		.dout(new_net_3903)
	);

	bfr new_net_3706_bfr_after (
		.din(_0115_),
		.dout(new_net_3706)
	);

	bfr new_net_3751_bfr_after (
		.din(_0293_),
		.dout(new_net_3751)
	);

	bfr new_net_3850_bfr_after (
		.din(_0730_),
		.dout(new_net_3850)
	);

	bfr new_net_3456_bfr_after (
		.din(_1588_),
		.dout(new_net_3456)
	);

	bfr new_net_3485_bfr_after (
		.din(_1018_),
		.dout(new_net_3485)
	);

	bfr new_net_3541_bfr_after (
		.din(_1235_),
		.dout(new_net_3541)
	);

	bfr new_net_3690_bfr_after (
		.din(_0029_),
		.dout(new_net_3690)
	);

	bfr new_net_20791_bfr_after (
		.din(new_net_3928),
		.dout(new_net_20791)
	);

	bfr new_net_20792_bfr_after (
		.din(new_net_20791),
		.dout(new_net_20792)
	);

	bfr new_net_20793_bfr_after (
		.din(new_net_20792),
		.dout(new_net_20793)
	);

	bfr new_net_20794_bfr_after (
		.din(new_net_20793),
		.dout(new_net_20794)
	);

	bfr new_net_20795_bfr_after (
		.din(new_net_20794),
		.dout(new_net_20795)
	);

	bfr new_net_20796_bfr_after (
		.din(new_net_20795),
		.dout(new_net_20796)
	);

	bfr new_net_20797_bfr_after (
		.din(new_net_20796),
		.dout(new_net_20797)
	);

	bfr new_net_20798_bfr_after (
		.din(new_net_20797),
		.dout(new_net_20798)
	);

	bfr new_net_20799_bfr_after (
		.din(new_net_20798),
		.dout(new_net_20799)
	);

	bfr new_net_20800_bfr_after (
		.din(new_net_20799),
		.dout(new_net_20800)
	);

	bfr new_net_20801_bfr_after (
		.din(new_net_20800),
		.dout(new_net_20801)
	);

	bfr new_net_20802_bfr_after (
		.din(new_net_20801),
		.dout(new_net_20802)
	);

	bfr new_net_20803_bfr_after (
		.din(new_net_20802),
		.dout(new_net_20803)
	);

	bfr new_net_20804_bfr_after (
		.din(new_net_20803),
		.dout(new_net_20804)
	);

	bfr new_net_20805_bfr_after (
		.din(new_net_20804),
		.dout(new_net_20805)
	);

	bfr new_net_20806_bfr_after (
		.din(new_net_20805),
		.dout(new_net_20806)
	);

	bfr new_net_20807_bfr_after (
		.din(new_net_20806),
		.dout(new_net_20807)
	);

	bfr new_net_20808_bfr_after (
		.din(new_net_20807),
		.dout(new_net_20808)
	);

	bfr new_net_20809_bfr_after (
		.din(new_net_20808),
		.dout(new_net_20809)
	);

	bfr new_net_20810_bfr_after (
		.din(new_net_20809),
		.dout(new_net_20810)
	);

	bfr new_net_20811_bfr_after (
		.din(new_net_20810),
		.dout(new_net_20811)
	);

	bfr new_net_20812_bfr_after (
		.din(new_net_20811),
		.dout(new_net_20812)
	);

	bfr new_net_20813_bfr_after (
		.din(new_net_20812),
		.dout(new_net_20813)
	);

	bfr new_net_20814_bfr_after (
		.din(new_net_20813),
		.dout(new_net_20814)
	);

	bfr new_net_20815_bfr_after (
		.din(new_net_20814),
		.dout(new_net_20815)
	);

	bfr new_net_20816_bfr_after (
		.din(new_net_20815),
		.dout(new_net_20816)
	);

	bfr new_net_20817_bfr_after (
		.din(new_net_20816),
		.dout(new_net_20817)
	);

	bfr new_net_20818_bfr_after (
		.din(new_net_20817),
		.dout(new_net_20818)
	);

	bfr new_net_20819_bfr_after (
		.din(new_net_20818),
		.dout(new_net_20819)
	);

	bfr new_net_20820_bfr_after (
		.din(new_net_20819),
		.dout(new_net_20820)
	);

	bfr new_net_20821_bfr_after (
		.din(new_net_20820),
		.dout(new_net_20821)
	);

	bfr new_net_20822_bfr_after (
		.din(new_net_20821),
		.dout(new_net_20822)
	);

	bfr new_net_20823_bfr_after (
		.din(new_net_20822),
		.dout(new_net_20823)
	);

	bfr new_net_20824_bfr_after (
		.din(new_net_20823),
		.dout(new_net_20824)
	);

	bfr new_net_20825_bfr_after (
		.din(new_net_20824),
		.dout(new_net_20825)
	);

	bfr new_net_20826_bfr_after (
		.din(new_net_20825),
		.dout(new_net_20826)
	);

	bfr new_net_20827_bfr_after (
		.din(new_net_20826),
		.dout(new_net_20827)
	);

	bfr new_net_20828_bfr_after (
		.din(new_net_20827),
		.dout(new_net_20828)
	);

	bfr new_net_20829_bfr_after (
		.din(new_net_20828),
		.dout(new_net_20829)
	);

	bfr new_net_20830_bfr_after (
		.din(new_net_20829),
		.dout(new_net_20830)
	);

	bfr new_net_20831_bfr_after (
		.din(new_net_20830),
		.dout(new_net_20831)
	);

	bfr new_net_20832_bfr_after (
		.din(new_net_20831),
		.dout(new_net_20832)
	);

	bfr new_net_20833_bfr_after (
		.din(new_net_20832),
		.dout(new_net_20833)
	);

	bfr new_net_20834_bfr_after (
		.din(new_net_20833),
		.dout(new_net_20834)
	);

	bfr new_net_20835_bfr_after (
		.din(new_net_20834),
		.dout(new_net_20835)
	);

	bfr new_net_20836_bfr_after (
		.din(new_net_20835),
		.dout(new_net_20836)
	);

	bfr new_net_20837_bfr_after (
		.din(new_net_20836),
		.dout(new_net_20837)
	);

	bfr new_net_20838_bfr_after (
		.din(new_net_20837),
		.dout(new_net_20838)
	);

	bfr new_net_20839_bfr_after (
		.din(new_net_20838),
		.dout(new_net_20839)
	);

	bfr new_net_20840_bfr_after (
		.din(new_net_20839),
		.dout(new_net_20840)
	);

	bfr new_net_20841_bfr_after (
		.din(new_net_20840),
		.dout(new_net_20841)
	);

	bfr new_net_20842_bfr_after (
		.din(new_net_20841),
		.dout(new_net_20842)
	);

	bfr new_net_20843_bfr_after (
		.din(new_net_20842),
		.dout(new_net_20843)
	);

	bfr new_net_20844_bfr_after (
		.din(new_net_20843),
		.dout(new_net_20844)
	);

	bfr new_net_20845_bfr_after (
		.din(new_net_20844),
		.dout(new_net_20845)
	);

	bfr new_net_20846_bfr_after (
		.din(new_net_20845),
		.dout(new_net_20846)
	);

	bfr new_net_20847_bfr_after (
		.din(new_net_20846),
		.dout(new_net_20847)
	);

	bfr new_net_20848_bfr_after (
		.din(new_net_20847),
		.dout(new_net_20848)
	);

	bfr new_net_20849_bfr_after (
		.din(new_net_20848),
		.dout(new_net_20849)
	);

	bfr new_net_20850_bfr_after (
		.din(new_net_20849),
		.dout(new_net_20850)
	);

	bfr new_net_20851_bfr_after (
		.din(new_net_20850),
		.dout(new_net_20851)
	);

	bfr new_net_20852_bfr_after (
		.din(new_net_20851),
		.dout(new_net_20852)
	);

	bfr new_net_20853_bfr_after (
		.din(new_net_20852),
		.dout(new_net_20853)
	);

	bfr new_net_20854_bfr_after (
		.din(new_net_20853),
		.dout(new_net_20854)
	);

	bfr new_net_20855_bfr_after (
		.din(new_net_20854),
		.dout(new_net_20855)
	);

	bfr new_net_20856_bfr_after (
		.din(new_net_20855),
		.dout(new_net_20856)
	);

	bfr new_net_20857_bfr_after (
		.din(new_net_20856),
		.dout(new_net_20857)
	);

	bfr new_net_20858_bfr_after (
		.din(new_net_20857),
		.dout(new_net_20858)
	);

	bfr new_net_20859_bfr_after (
		.din(new_net_20858),
		.dout(new_net_20859)
	);

	bfr new_net_20860_bfr_after (
		.din(new_net_20859),
		.dout(new_net_20860)
	);

	bfr new_net_20861_bfr_after (
		.din(new_net_20860),
		.dout(new_net_20861)
	);

	bfr new_net_20862_bfr_after (
		.din(new_net_20861),
		.dout(new_net_20862)
	);

	bfr new_net_20863_bfr_after (
		.din(new_net_20862),
		.dout(new_net_20863)
	);

	bfr new_net_20864_bfr_after (
		.din(new_net_20863),
		.dout(new_net_20864)
	);

	bfr new_net_20865_bfr_after (
		.din(new_net_20864),
		.dout(new_net_20865)
	);

	bfr new_net_20866_bfr_after (
		.din(new_net_20865),
		.dout(new_net_20866)
	);

	bfr new_net_20867_bfr_after (
		.din(new_net_20866),
		.dout(new_net_20867)
	);

	bfr new_net_20868_bfr_after (
		.din(new_net_20867),
		.dout(new_net_20868)
	);

	bfr new_net_20869_bfr_after (
		.din(new_net_20868),
		.dout(new_net_20869)
	);

	bfr new_net_20870_bfr_after (
		.din(new_net_20869),
		.dout(new_net_20870)
	);

	bfr new_net_20871_bfr_after (
		.din(new_net_20870),
		.dout(new_net_20871)
	);

	bfr new_net_20872_bfr_after (
		.din(new_net_20871),
		.dout(new_net_20872)
	);

	bfr new_net_20873_bfr_after (
		.din(new_net_20872),
		.dout(new_net_20873)
	);

	bfr new_net_20874_bfr_after (
		.din(new_net_20873),
		.dout(new_net_20874)
	);

	bfr new_net_20875_bfr_after (
		.din(new_net_20874),
		.dout(new_net_20875)
	);

	bfr new_net_20876_bfr_after (
		.din(new_net_20875),
		.dout(new_net_20876)
	);

	bfr new_net_20877_bfr_after (
		.din(new_net_20876),
		.dout(new_net_20877)
	);

	bfr new_net_20878_bfr_after (
		.din(new_net_20877),
		.dout(new_net_20878)
	);

	bfr new_net_20879_bfr_after (
		.din(new_net_20878),
		.dout(new_net_20879)
	);

	bfr new_net_20880_bfr_after (
		.din(new_net_20879),
		.dout(new_net_20880)
	);

	bfr new_net_20881_bfr_after (
		.din(new_net_20880),
		.dout(new_net_20881)
	);

	bfr new_net_20882_bfr_after (
		.din(new_net_20881),
		.dout(new_net_20882)
	);

	bfr new_net_20883_bfr_after (
		.din(new_net_20882),
		.dout(new_net_20883)
	);

	bfr new_net_20884_bfr_after (
		.din(new_net_20883),
		.dout(new_net_20884)
	);

	bfr new_net_20885_bfr_after (
		.din(new_net_20884),
		.dout(new_net_20885)
	);

	bfr new_net_20886_bfr_after (
		.din(new_net_20885),
		.dout(new_net_20886)
	);

	bfr new_net_20887_bfr_after (
		.din(new_net_20886),
		.dout(new_net_20887)
	);

	bfr new_net_20888_bfr_after (
		.din(new_net_20887),
		.dout(new_net_20888)
	);

	bfr new_net_20889_bfr_after (
		.din(new_net_20888),
		.dout(new_net_20889)
	);

	bfr new_net_20890_bfr_after (
		.din(new_net_20889),
		.dout(new_net_20890)
	);

	bfr new_net_20891_bfr_after (
		.din(new_net_20890),
		.dout(new_net_20891)
	);

	bfr new_net_20892_bfr_after (
		.din(new_net_20891),
		.dout(new_net_20892)
	);

	bfr new_net_20893_bfr_after (
		.din(new_net_20892),
		.dout(new_net_20893)
	);

	bfr new_net_20894_bfr_after (
		.din(new_net_20893),
		.dout(new_net_20894)
	);

	bfr new_net_20895_bfr_after (
		.din(new_net_20894),
		.dout(new_net_20895)
	);

	bfr new_net_20896_bfr_after (
		.din(new_net_20895),
		.dout(new_net_20896)
	);

	bfr new_net_20897_bfr_after (
		.din(new_net_20896),
		.dout(new_net_20897)
	);

	bfr new_net_20898_bfr_after (
		.din(new_net_20897),
		.dout(new_net_20898)
	);

	bfr new_net_20899_bfr_after (
		.din(new_net_20898),
		.dout(new_net_20899)
	);

	bfr new_net_20900_bfr_after (
		.din(new_net_20899),
		.dout(new_net_20900)
	);

	bfr new_net_20901_bfr_after (
		.din(new_net_20900),
		.dout(new_net_20901)
	);

	bfr new_net_20902_bfr_after (
		.din(new_net_20901),
		.dout(new_net_20902)
	);

	bfr new_net_20903_bfr_after (
		.din(new_net_20902),
		.dout(new_net_20903)
	);

	bfr new_net_20904_bfr_after (
		.din(new_net_20903),
		.dout(new_net_20904)
	);

	bfr new_net_20905_bfr_after (
		.din(new_net_20904),
		.dout(new_net_20905)
	);

	bfr N3895_bfr_after (
		.din(new_net_20905),
		.dout(N3895)
	);

	bfr new_net_3731_bfr_after (
		.din(_0197_),
		.dout(new_net_3731)
	);

	bfr new_net_3499_bfr_after (
		.din(_1089_),
		.dout(new_net_3499)
	);

	bfr new_net_3616_bfr_after (
		.din(_1533_),
		.dout(new_net_3616)
	);

	bfr new_net_3674_bfr_after (
		.din(_1786_),
		.dout(new_net_3674)
	);

	bfr new_net_3689_bfr_after (
		.din(_0026_),
		.dout(new_net_3689)
	);

	bfr new_net_3693_bfr_after (
		.din(_0039_),
		.dout(new_net_3693)
	);

	bfr new_net_3764_bfr_after (
		.din(_0363_),
		.dout(new_net_3764)
	);

	bfr new_net_3827_bfr_after (
		.din(_0637_),
		.dout(new_net_3827)
	);

	bfr new_net_3892_bfr_after (
		.din(_0909_),
		.dout(new_net_3892)
	);

	bfr new_net_3464_bfr_after (
		.din(_0143_),
		.dout(new_net_3464)
	);

	bfr new_net_3566_bfr_after (
		.din(_1330_),
		.dout(new_net_3566)
	);

	bfr new_net_3588_bfr_after (
		.din(_1418_),
		.dout(new_net_3588)
	);

	bfr new_net_3704_bfr_after (
		.din(_0075_),
		.dout(new_net_3704)
	);

	bfr new_net_3789_bfr_after (
		.din(_0469_),
		.dout(new_net_3789)
	);

	bfr new_net_3828_bfr_after (
		.din(_0640_),
		.dout(new_net_3828)
	);

	bfr new_net_3861_bfr_after (
		.din(_0782_),
		.dout(new_net_3861)
	);

	bfr new_net_3901_bfr_after (
		.din(_0948_),
		.dout(new_net_3901)
	);

	bfr new_net_20906_bfr_after (
		.din(new_net_3918),
		.dout(new_net_20906)
	);

	bfr new_net_20907_bfr_after (
		.din(new_net_20906),
		.dout(new_net_20907)
	);

	bfr new_net_20908_bfr_after (
		.din(new_net_20907),
		.dout(new_net_20908)
	);

	bfr new_net_20909_bfr_after (
		.din(new_net_20908),
		.dout(new_net_20909)
	);

	bfr new_net_20910_bfr_after (
		.din(new_net_20909),
		.dout(new_net_20910)
	);

	bfr new_net_20911_bfr_after (
		.din(new_net_20910),
		.dout(new_net_20911)
	);

	bfr new_net_20912_bfr_after (
		.din(new_net_20911),
		.dout(new_net_20912)
	);

	bfr new_net_20913_bfr_after (
		.din(new_net_20912),
		.dout(new_net_20913)
	);

	bfr new_net_20914_bfr_after (
		.din(new_net_20913),
		.dout(new_net_20914)
	);

	bfr new_net_20915_bfr_after (
		.din(new_net_20914),
		.dout(new_net_20915)
	);

	bfr new_net_20916_bfr_after (
		.din(new_net_20915),
		.dout(new_net_20916)
	);

	bfr new_net_20917_bfr_after (
		.din(new_net_20916),
		.dout(new_net_20917)
	);

	bfr new_net_20918_bfr_after (
		.din(new_net_20917),
		.dout(new_net_20918)
	);

	bfr new_net_20919_bfr_after (
		.din(new_net_20918),
		.dout(new_net_20919)
	);

	bfr new_net_20920_bfr_after (
		.din(new_net_20919),
		.dout(new_net_20920)
	);

	bfr new_net_20921_bfr_after (
		.din(new_net_20920),
		.dout(new_net_20921)
	);

	bfr new_net_20922_bfr_after (
		.din(new_net_20921),
		.dout(new_net_20922)
	);

	bfr new_net_20923_bfr_after (
		.din(new_net_20922),
		.dout(new_net_20923)
	);

	bfr new_net_20924_bfr_after (
		.din(new_net_20923),
		.dout(new_net_20924)
	);

	bfr new_net_20925_bfr_after (
		.din(new_net_20924),
		.dout(new_net_20925)
	);

	bfr new_net_20926_bfr_after (
		.din(new_net_20925),
		.dout(new_net_20926)
	);

	bfr new_net_20927_bfr_after (
		.din(new_net_20926),
		.dout(new_net_20927)
	);

	bfr new_net_20928_bfr_after (
		.din(new_net_20927),
		.dout(new_net_20928)
	);

	bfr new_net_20929_bfr_after (
		.din(new_net_20928),
		.dout(new_net_20929)
	);

	bfr new_net_20930_bfr_after (
		.din(new_net_20929),
		.dout(new_net_20930)
	);

	bfr new_net_20931_bfr_after (
		.din(new_net_20930),
		.dout(new_net_20931)
	);

	bfr new_net_20932_bfr_after (
		.din(new_net_20931),
		.dout(new_net_20932)
	);

	bfr N6220_bfr_after (
		.din(new_net_20932),
		.dout(N6220)
	);

	bfr new_net_3863_bfr_after (
		.din(_0789_),
		.dout(new_net_3863)
	);

	bfr new_net_3574_bfr_after (
		.din(_1354_),
		.dout(new_net_3574)
	);

	bfr new_net_3717_bfr_after (
		.din(_0151_),
		.dout(new_net_3717)
	);

	bfr new_net_3757_bfr_after (
		.din(_0313_),
		.dout(new_net_3757)
	);

	bfr new_net_3912_bfr_after (
		.din(_0995_),
		.dout(new_net_3912)
	);

	bfr new_net_3564_bfr_after (
		.din(_1324_),
		.dout(new_net_3564)
	);

	bfr new_net_3584_bfr_after (
		.din(_1406_),
		.dout(new_net_3584)
	);

	bfr new_net_3640_bfr_after (
		.din(_1640_),
		.dout(new_net_3640)
	);

	bfr new_net_3648_bfr_after (
		.din(_1667_),
		.dout(new_net_3648)
	);

	bfr new_net_3664_bfr_after (
		.din(_1753_),
		.dout(new_net_3664)
	);

	bfr new_net_3745_bfr_after (
		.din(_0273_),
		.dout(new_net_3745)
	);

	bfr new_net_3812_bfr_after (
		.din(_0567_),
		.dout(new_net_3812)
	);

	bfr new_net_3849_bfr_after (
		.din(_0727_),
		.dout(new_net_3849)
	);

	bfr new_net_3855_bfr_after (
		.din(_0747_),
		.dout(new_net_3855)
	);

	bfr new_net_3857_bfr_after (
		.din(_0754_),
		.dout(new_net_3857)
	);

	bfr new_net_3462_bfr_after (
		.din(_0077_),
		.dout(new_net_3462)
	);

	bfr new_net_3723_bfr_after (
		.din(_0171_),
		.dout(new_net_3723)
	);

	bfr new_net_3506_bfr_after (
		.din(_1110_),
		.dout(new_net_3506)
	);

	bfr new_net_3551_bfr_after (
		.din(_1265_),
		.dout(new_net_3551)
	);

	bfr new_net_3697_bfr_after (
		.din(_0052_),
		.dout(new_net_3697)
	);

	bfr new_net_20933_bfr_after (
		.din(new_net_3956),
		.dout(new_net_20933)
	);

	bfr new_net_20934_bfr_after (
		.din(new_net_20933),
		.dout(new_net_20934)
	);

	bfr new_net_20935_bfr_after (
		.din(new_net_20934),
		.dout(new_net_20935)
	);

	bfr new_net_20936_bfr_after (
		.din(new_net_20935),
		.dout(new_net_20936)
	);

	bfr new_net_20937_bfr_after (
		.din(new_net_20936),
		.dout(new_net_20937)
	);

	bfr new_net_20938_bfr_after (
		.din(new_net_20937),
		.dout(new_net_20938)
	);

	bfr new_net_20939_bfr_after (
		.din(new_net_20938),
		.dout(new_net_20939)
	);

	bfr new_net_20940_bfr_after (
		.din(new_net_20939),
		.dout(new_net_20940)
	);

	bfr new_net_20941_bfr_after (
		.din(new_net_20940),
		.dout(new_net_20941)
	);

	bfr new_net_20942_bfr_after (
		.din(new_net_20941),
		.dout(new_net_20942)
	);

	bfr new_net_20943_bfr_after (
		.din(new_net_20942),
		.dout(new_net_20943)
	);

	bfr new_net_20944_bfr_after (
		.din(new_net_20943),
		.dout(new_net_20944)
	);

	bfr new_net_20945_bfr_after (
		.din(new_net_20944),
		.dout(new_net_20945)
	);

	bfr new_net_20946_bfr_after (
		.din(new_net_20945),
		.dout(new_net_20946)
	);

	bfr new_net_20947_bfr_after (
		.din(new_net_20946),
		.dout(new_net_20947)
	);

	bfr new_net_20948_bfr_after (
		.din(new_net_20947),
		.dout(new_net_20948)
	);

	bfr new_net_20949_bfr_after (
		.din(new_net_20948),
		.dout(new_net_20949)
	);

	bfr new_net_20950_bfr_after (
		.din(new_net_20949),
		.dout(new_net_20950)
	);

	bfr new_net_20951_bfr_after (
		.din(new_net_20950),
		.dout(new_net_20951)
	);

	bfr new_net_20952_bfr_after (
		.din(new_net_20951),
		.dout(new_net_20952)
	);

	bfr new_net_20953_bfr_after (
		.din(new_net_20952),
		.dout(new_net_20953)
	);

	bfr new_net_20954_bfr_after (
		.din(new_net_20953),
		.dout(new_net_20954)
	);

	bfr new_net_20955_bfr_after (
		.din(new_net_20954),
		.dout(new_net_20955)
	);

	bfr new_net_20956_bfr_after (
		.din(new_net_20955),
		.dout(new_net_20956)
	);

	bfr new_net_20957_bfr_after (
		.din(new_net_20956),
		.dout(new_net_20957)
	);

	bfr new_net_20958_bfr_after (
		.din(new_net_20957),
		.dout(new_net_20958)
	);

	bfr new_net_20959_bfr_after (
		.din(new_net_20958),
		.dout(new_net_20959)
	);

	bfr new_net_20960_bfr_after (
		.din(new_net_20959),
		.dout(new_net_20960)
	);

	bfr new_net_20961_bfr_after (
		.din(new_net_20960),
		.dout(new_net_20961)
	);

	bfr new_net_20962_bfr_after (
		.din(new_net_20961),
		.dout(new_net_20962)
	);

	bfr new_net_20963_bfr_after (
		.din(new_net_20962),
		.dout(new_net_20963)
	);

	bfr new_net_20964_bfr_after (
		.din(new_net_20963),
		.dout(new_net_20964)
	);

	bfr new_net_20965_bfr_after (
		.din(new_net_20964),
		.dout(new_net_20965)
	);

	bfr new_net_20966_bfr_after (
		.din(new_net_20965),
		.dout(new_net_20966)
	);

	bfr new_net_20967_bfr_after (
		.din(new_net_20966),
		.dout(new_net_20967)
	);

	bfr new_net_20968_bfr_after (
		.din(new_net_20967),
		.dout(new_net_20968)
	);

	bfr new_net_20969_bfr_after (
		.din(new_net_20968),
		.dout(new_net_20969)
	);

	bfr new_net_20970_bfr_after (
		.din(new_net_20969),
		.dout(new_net_20970)
	);

	bfr new_net_20971_bfr_after (
		.din(new_net_20970),
		.dout(new_net_20971)
	);

	bfr new_net_20972_bfr_after (
		.din(new_net_20971),
		.dout(new_net_20972)
	);

	bfr new_net_20973_bfr_after (
		.din(new_net_20972),
		.dout(new_net_20973)
	);

	bfr new_net_20974_bfr_after (
		.din(new_net_20973),
		.dout(new_net_20974)
	);

	bfr new_net_20975_bfr_after (
		.din(new_net_20974),
		.dout(new_net_20975)
	);

	bfr new_net_20976_bfr_after (
		.din(new_net_20975),
		.dout(new_net_20976)
	);

	bfr new_net_20977_bfr_after (
		.din(new_net_20976),
		.dout(new_net_20977)
	);

	bfr new_net_20978_bfr_after (
		.din(new_net_20977),
		.dout(new_net_20978)
	);

	bfr new_net_20979_bfr_after (
		.din(new_net_20978),
		.dout(new_net_20979)
	);

	bfr new_net_20980_bfr_after (
		.din(new_net_20979),
		.dout(new_net_20980)
	);

	bfr new_net_20981_bfr_after (
		.din(new_net_20980),
		.dout(new_net_20981)
	);

	bfr new_net_20982_bfr_after (
		.din(new_net_20981),
		.dout(new_net_20982)
	);

	bfr new_net_20983_bfr_after (
		.din(new_net_20982),
		.dout(new_net_20983)
	);

	bfr new_net_20984_bfr_after (
		.din(new_net_20983),
		.dout(new_net_20984)
	);

	bfr new_net_20985_bfr_after (
		.din(new_net_20984),
		.dout(new_net_20985)
	);

	bfr new_net_20986_bfr_after (
		.din(new_net_20985),
		.dout(new_net_20986)
	);

	bfr new_net_20987_bfr_after (
		.din(new_net_20986),
		.dout(new_net_20987)
	);

	bfr new_net_20988_bfr_after (
		.din(new_net_20987),
		.dout(new_net_20988)
	);

	bfr new_net_20989_bfr_after (
		.din(new_net_20988),
		.dout(new_net_20989)
	);

	bfr new_net_20990_bfr_after (
		.din(new_net_20989),
		.dout(new_net_20990)
	);

	bfr new_net_20991_bfr_after (
		.din(new_net_20990),
		.dout(new_net_20991)
	);

	bfr new_net_20992_bfr_after (
		.din(new_net_20991),
		.dout(new_net_20992)
	);

	bfr new_net_20993_bfr_after (
		.din(new_net_20992),
		.dout(new_net_20993)
	);

	bfr new_net_20994_bfr_after (
		.din(new_net_20993),
		.dout(new_net_20994)
	);

	bfr new_net_20995_bfr_after (
		.din(new_net_20994),
		.dout(new_net_20995)
	);

	bfr new_net_20996_bfr_after (
		.din(new_net_20995),
		.dout(new_net_20996)
	);

	bfr new_net_20997_bfr_after (
		.din(new_net_20996),
		.dout(new_net_20997)
	);

	bfr new_net_20998_bfr_after (
		.din(new_net_20997),
		.dout(new_net_20998)
	);

	bfr new_net_20999_bfr_after (
		.din(new_net_20998),
		.dout(new_net_20999)
	);

	bfr new_net_21000_bfr_after (
		.din(new_net_20999),
		.dout(new_net_21000)
	);

	bfr new_net_21001_bfr_after (
		.din(new_net_21000),
		.dout(new_net_21001)
	);

	bfr new_net_21002_bfr_after (
		.din(new_net_21001),
		.dout(new_net_21002)
	);

	bfr new_net_21003_bfr_after (
		.din(new_net_21002),
		.dout(new_net_21003)
	);

	bfr new_net_21004_bfr_after (
		.din(new_net_21003),
		.dout(new_net_21004)
	);

	bfr new_net_21005_bfr_after (
		.din(new_net_21004),
		.dout(new_net_21005)
	);

	bfr new_net_21006_bfr_after (
		.din(new_net_21005),
		.dout(new_net_21006)
	);

	bfr new_net_21007_bfr_after (
		.din(new_net_21006),
		.dout(new_net_21007)
	);

	bfr new_net_21008_bfr_after (
		.din(new_net_21007),
		.dout(new_net_21008)
	);

	bfr new_net_21009_bfr_after (
		.din(new_net_21008),
		.dout(new_net_21009)
	);

	bfr new_net_21010_bfr_after (
		.din(new_net_21009),
		.dout(new_net_21010)
	);

	bfr new_net_21011_bfr_after (
		.din(new_net_21010),
		.dout(new_net_21011)
	);

	bfr new_net_21012_bfr_after (
		.din(new_net_21011),
		.dout(new_net_21012)
	);

	bfr new_net_21013_bfr_after (
		.din(new_net_21012),
		.dout(new_net_21013)
	);

	bfr new_net_21014_bfr_after (
		.din(new_net_21013),
		.dout(new_net_21014)
	);

	bfr new_net_21015_bfr_after (
		.din(new_net_21014),
		.dout(new_net_21015)
	);

	bfr new_net_21016_bfr_after (
		.din(new_net_21015),
		.dout(new_net_21016)
	);

	bfr new_net_21017_bfr_after (
		.din(new_net_21016),
		.dout(new_net_21017)
	);

	bfr new_net_21018_bfr_after (
		.din(new_net_21017),
		.dout(new_net_21018)
	);

	bfr new_net_21019_bfr_after (
		.din(new_net_21018),
		.dout(new_net_21019)
	);

	bfr new_net_21020_bfr_after (
		.din(new_net_21019),
		.dout(new_net_21020)
	);

	bfr new_net_21021_bfr_after (
		.din(new_net_21020),
		.dout(new_net_21021)
	);

	bfr new_net_21022_bfr_after (
		.din(new_net_21021),
		.dout(new_net_21022)
	);

	bfr new_net_21023_bfr_after (
		.din(new_net_21022),
		.dout(new_net_21023)
	);

	bfr new_net_21024_bfr_after (
		.din(new_net_21023),
		.dout(new_net_21024)
	);

	bfr new_net_21025_bfr_after (
		.din(new_net_21024),
		.dout(new_net_21025)
	);

	bfr new_net_21026_bfr_after (
		.din(new_net_21025),
		.dout(new_net_21026)
	);

	bfr new_net_21027_bfr_after (
		.din(new_net_21026),
		.dout(new_net_21027)
	);

	bfr new_net_21028_bfr_after (
		.din(new_net_21027),
		.dout(new_net_21028)
	);

	bfr new_net_21029_bfr_after (
		.din(new_net_21028),
		.dout(new_net_21029)
	);

	bfr new_net_21030_bfr_after (
		.din(new_net_21029),
		.dout(new_net_21030)
	);

	bfr new_net_21031_bfr_after (
		.din(new_net_21030),
		.dout(new_net_21031)
	);

	bfr new_net_21032_bfr_after (
		.din(new_net_21031),
		.dout(new_net_21032)
	);

	bfr new_net_21033_bfr_after (
		.din(new_net_21032),
		.dout(new_net_21033)
	);

	bfr new_net_21034_bfr_after (
		.din(new_net_21033),
		.dout(new_net_21034)
	);

	bfr new_net_21035_bfr_after (
		.din(new_net_21034),
		.dout(new_net_21035)
	);

	bfr new_net_21036_bfr_after (
		.din(new_net_21035),
		.dout(new_net_21036)
	);

	bfr new_net_21037_bfr_after (
		.din(new_net_21036),
		.dout(new_net_21037)
	);

	bfr new_net_21038_bfr_after (
		.din(new_net_21037),
		.dout(new_net_21038)
	);

	bfr new_net_21039_bfr_after (
		.din(new_net_21038),
		.dout(new_net_21039)
	);

	bfr N4241_bfr_after (
		.din(new_net_21039),
		.dout(N4241)
	);

	bfr new_net_3776_bfr_after (
		.din(_0402_),
		.dout(new_net_3776)
	);

	bfr new_net_21040_bfr_after (
		.din(new_net_3974),
		.dout(new_net_21040)
	);

	bfr new_net_21041_bfr_after (
		.din(new_net_21040),
		.dout(new_net_21041)
	);

	bfr new_net_21042_bfr_after (
		.din(new_net_21041),
		.dout(new_net_21042)
	);

	bfr new_net_21043_bfr_after (
		.din(new_net_21042),
		.dout(new_net_21043)
	);

	bfr new_net_21044_bfr_after (
		.din(new_net_21043),
		.dout(new_net_21044)
	);

	bfr new_net_21045_bfr_after (
		.din(new_net_21044),
		.dout(new_net_21045)
	);

	bfr new_net_21046_bfr_after (
		.din(new_net_21045),
		.dout(new_net_21046)
	);

	bfr new_net_21047_bfr_after (
		.din(new_net_21046),
		.dout(new_net_21047)
	);

	bfr new_net_21048_bfr_after (
		.din(new_net_21047),
		.dout(new_net_21048)
	);

	bfr new_net_21049_bfr_after (
		.din(new_net_21048),
		.dout(new_net_21049)
	);

	bfr new_net_21050_bfr_after (
		.din(new_net_21049),
		.dout(new_net_21050)
	);

	bfr new_net_21051_bfr_after (
		.din(new_net_21050),
		.dout(new_net_21051)
	);

	bfr new_net_21052_bfr_after (
		.din(new_net_21051),
		.dout(new_net_21052)
	);

	bfr new_net_21053_bfr_after (
		.din(new_net_21052),
		.dout(new_net_21053)
	);

	bfr new_net_21054_bfr_after (
		.din(new_net_21053),
		.dout(new_net_21054)
	);

	bfr new_net_21055_bfr_after (
		.din(new_net_21054),
		.dout(new_net_21055)
	);

	bfr new_net_21056_bfr_after (
		.din(new_net_21055),
		.dout(new_net_21056)
	);

	bfr new_net_21057_bfr_after (
		.din(new_net_21056),
		.dout(new_net_21057)
	);

	bfr new_net_21058_bfr_after (
		.din(new_net_21057),
		.dout(new_net_21058)
	);

	bfr new_net_21059_bfr_after (
		.din(new_net_21058),
		.dout(new_net_21059)
	);

	bfr new_net_21060_bfr_after (
		.din(new_net_21059),
		.dout(new_net_21060)
	);

	bfr new_net_21061_bfr_after (
		.din(new_net_21060),
		.dout(new_net_21061)
	);

	bfr new_net_21062_bfr_after (
		.din(new_net_21061),
		.dout(new_net_21062)
	);

	bfr new_net_21063_bfr_after (
		.din(new_net_21062),
		.dout(new_net_21063)
	);

	bfr new_net_21064_bfr_after (
		.din(new_net_21063),
		.dout(new_net_21064)
	);

	bfr new_net_21065_bfr_after (
		.din(new_net_21064),
		.dout(new_net_21065)
	);

	bfr new_net_21066_bfr_after (
		.din(new_net_21065),
		.dout(new_net_21066)
	);

	bfr new_net_21067_bfr_after (
		.din(new_net_21066),
		.dout(new_net_21067)
	);

	bfr new_net_21068_bfr_after (
		.din(new_net_21067),
		.dout(new_net_21068)
	);

	bfr new_net_21069_bfr_after (
		.din(new_net_21068),
		.dout(new_net_21069)
	);

	bfr new_net_21070_bfr_after (
		.din(new_net_21069),
		.dout(new_net_21070)
	);

	bfr new_net_21071_bfr_after (
		.din(new_net_21070),
		.dout(new_net_21071)
	);

	bfr new_net_21072_bfr_after (
		.din(new_net_21071),
		.dout(new_net_21072)
	);

	bfr new_net_21073_bfr_after (
		.din(new_net_21072),
		.dout(new_net_21073)
	);

	bfr new_net_21074_bfr_after (
		.din(new_net_21073),
		.dout(new_net_21074)
	);

	bfr new_net_21075_bfr_after (
		.din(new_net_21074),
		.dout(new_net_21075)
	);

	bfr new_net_21076_bfr_after (
		.din(new_net_21075),
		.dout(new_net_21076)
	);

	bfr new_net_21077_bfr_after (
		.din(new_net_21076),
		.dout(new_net_21077)
	);

	bfr new_net_21078_bfr_after (
		.din(new_net_21077),
		.dout(new_net_21078)
	);

	bfr new_net_21079_bfr_after (
		.din(new_net_21078),
		.dout(new_net_21079)
	);

	bfr new_net_21080_bfr_after (
		.din(new_net_21079),
		.dout(new_net_21080)
	);

	bfr new_net_21081_bfr_after (
		.din(new_net_21080),
		.dout(new_net_21081)
	);

	bfr new_net_21082_bfr_after (
		.din(new_net_21081),
		.dout(new_net_21082)
	);

	bfr new_net_21083_bfr_after (
		.din(new_net_21082),
		.dout(new_net_21083)
	);

	bfr new_net_21084_bfr_after (
		.din(new_net_21083),
		.dout(new_net_21084)
	);

	bfr new_net_21085_bfr_after (
		.din(new_net_21084),
		.dout(new_net_21085)
	);

	bfr new_net_21086_bfr_after (
		.din(new_net_21085),
		.dout(new_net_21086)
	);

	bfr new_net_21087_bfr_after (
		.din(new_net_21086),
		.dout(new_net_21087)
	);

	bfr new_net_21088_bfr_after (
		.din(new_net_21087),
		.dout(new_net_21088)
	);

	bfr new_net_21089_bfr_after (
		.din(new_net_21088),
		.dout(new_net_21089)
	);

	bfr new_net_21090_bfr_after (
		.din(new_net_21089),
		.dout(new_net_21090)
	);

	bfr new_net_21091_bfr_after (
		.din(new_net_21090),
		.dout(new_net_21091)
	);

	bfr new_net_21092_bfr_after (
		.din(new_net_21091),
		.dout(new_net_21092)
	);

	bfr new_net_21093_bfr_after (
		.din(new_net_21092),
		.dout(new_net_21093)
	);

	bfr new_net_21094_bfr_after (
		.din(new_net_21093),
		.dout(new_net_21094)
	);

	bfr new_net_21095_bfr_after (
		.din(new_net_21094),
		.dout(new_net_21095)
	);

	bfr new_net_21096_bfr_after (
		.din(new_net_21095),
		.dout(new_net_21096)
	);

	bfr new_net_21097_bfr_after (
		.din(new_net_21096),
		.dout(new_net_21097)
	);

	bfr new_net_21098_bfr_after (
		.din(new_net_21097),
		.dout(new_net_21098)
	);

	bfr new_net_21099_bfr_after (
		.din(new_net_21098),
		.dout(new_net_21099)
	);

	bfr new_net_21100_bfr_after (
		.din(new_net_21099),
		.dout(new_net_21100)
	);

	bfr new_net_21101_bfr_after (
		.din(new_net_21100),
		.dout(new_net_21101)
	);

	bfr new_net_21102_bfr_after (
		.din(new_net_21101),
		.dout(new_net_21102)
	);

	bfr new_net_21103_bfr_after (
		.din(new_net_21102),
		.dout(new_net_21103)
	);

	bfr new_net_21104_bfr_after (
		.din(new_net_21103),
		.dout(new_net_21104)
	);

	bfr new_net_21105_bfr_after (
		.din(new_net_21104),
		.dout(new_net_21105)
	);

	bfr new_net_21106_bfr_after (
		.din(new_net_21105),
		.dout(new_net_21106)
	);

	bfr new_net_21107_bfr_after (
		.din(new_net_21106),
		.dout(new_net_21107)
	);

	bfr new_net_21108_bfr_after (
		.din(new_net_21107),
		.dout(new_net_21108)
	);

	bfr new_net_21109_bfr_after (
		.din(new_net_21108),
		.dout(new_net_21109)
	);

	bfr new_net_21110_bfr_after (
		.din(new_net_21109),
		.dout(new_net_21110)
	);

	bfr new_net_21111_bfr_after (
		.din(new_net_21110),
		.dout(new_net_21111)
	);

	bfr new_net_21112_bfr_after (
		.din(new_net_21111),
		.dout(new_net_21112)
	);

	bfr new_net_21113_bfr_after (
		.din(new_net_21112),
		.dout(new_net_21113)
	);

	bfr new_net_21114_bfr_after (
		.din(new_net_21113),
		.dout(new_net_21114)
	);

	bfr new_net_21115_bfr_after (
		.din(new_net_21114),
		.dout(new_net_21115)
	);

	bfr new_net_21116_bfr_after (
		.din(new_net_21115),
		.dout(new_net_21116)
	);

	bfr new_net_21117_bfr_after (
		.din(new_net_21116),
		.dout(new_net_21117)
	);

	bfr new_net_21118_bfr_after (
		.din(new_net_21117),
		.dout(new_net_21118)
	);

	bfr new_net_21119_bfr_after (
		.din(new_net_21118),
		.dout(new_net_21119)
	);

	bfr new_net_21120_bfr_after (
		.din(new_net_21119),
		.dout(new_net_21120)
	);

	bfr new_net_21121_bfr_after (
		.din(new_net_21120),
		.dout(new_net_21121)
	);

	bfr new_net_21122_bfr_after (
		.din(new_net_21121),
		.dout(new_net_21122)
	);

	bfr new_net_21123_bfr_after (
		.din(new_net_21122),
		.dout(new_net_21123)
	);

	bfr new_net_21124_bfr_after (
		.din(new_net_21123),
		.dout(new_net_21124)
	);

	bfr new_net_21125_bfr_after (
		.din(new_net_21124),
		.dout(new_net_21125)
	);

	bfr new_net_21126_bfr_after (
		.din(new_net_21125),
		.dout(new_net_21126)
	);

	bfr new_net_21127_bfr_after (
		.din(new_net_21126),
		.dout(new_net_21127)
	);

	bfr new_net_21128_bfr_after (
		.din(new_net_21127),
		.dout(new_net_21128)
	);

	bfr new_net_21129_bfr_after (
		.din(new_net_21128),
		.dout(new_net_21129)
	);

	bfr new_net_21130_bfr_after (
		.din(new_net_21129),
		.dout(new_net_21130)
	);

	bfr new_net_21131_bfr_after (
		.din(new_net_21130),
		.dout(new_net_21131)
	);

	bfr new_net_21132_bfr_after (
		.din(new_net_21131),
		.dout(new_net_21132)
	);

	bfr new_net_21133_bfr_after (
		.din(new_net_21132),
		.dout(new_net_21133)
	);

	bfr new_net_21134_bfr_after (
		.din(new_net_21133),
		.dout(new_net_21134)
	);

	bfr new_net_21135_bfr_after (
		.din(new_net_21134),
		.dout(new_net_21135)
	);

	bfr new_net_21136_bfr_after (
		.din(new_net_21135),
		.dout(new_net_21136)
	);

	bfr new_net_21137_bfr_after (
		.din(new_net_21136),
		.dout(new_net_21137)
	);

	bfr new_net_21138_bfr_after (
		.din(new_net_21137),
		.dout(new_net_21138)
	);

	bfr new_net_21139_bfr_after (
		.din(new_net_21138),
		.dout(new_net_21139)
	);

	bfr new_net_21140_bfr_after (
		.din(new_net_21139),
		.dout(new_net_21140)
	);

	bfr new_net_21141_bfr_after (
		.din(new_net_21140),
		.dout(new_net_21141)
	);

	bfr new_net_21142_bfr_after (
		.din(new_net_21141),
		.dout(new_net_21142)
	);

	bfr new_net_21143_bfr_after (
		.din(new_net_21142),
		.dout(new_net_21143)
	);

	bfr new_net_21144_bfr_after (
		.din(new_net_21143),
		.dout(new_net_21144)
	);

	bfr new_net_21145_bfr_after (
		.din(new_net_21144),
		.dout(new_net_21145)
	);

	bfr new_net_21146_bfr_after (
		.din(new_net_21145),
		.dout(new_net_21146)
	);

	bfr new_net_21147_bfr_after (
		.din(new_net_21146),
		.dout(new_net_21147)
	);

	bfr new_net_21148_bfr_after (
		.din(new_net_21147),
		.dout(new_net_21148)
	);

	bfr new_net_21149_bfr_after (
		.din(new_net_21148),
		.dout(new_net_21149)
	);

	bfr new_net_21150_bfr_after (
		.din(new_net_21149),
		.dout(new_net_21150)
	);

	bfr new_net_21151_bfr_after (
		.din(new_net_21150),
		.dout(new_net_21151)
	);

	bfr new_net_21152_bfr_after (
		.din(new_net_21151),
		.dout(new_net_21152)
	);

	bfr new_net_21153_bfr_after (
		.din(new_net_21152),
		.dout(new_net_21153)
	);

	bfr new_net_21154_bfr_after (
		.din(new_net_21153),
		.dout(new_net_21154)
	);

	bfr new_net_21155_bfr_after (
		.din(new_net_21154),
		.dout(new_net_21155)
	);

	bfr new_net_21156_bfr_after (
		.din(new_net_21155),
		.dout(new_net_21156)
	);

	bfr new_net_21157_bfr_after (
		.din(new_net_21156),
		.dout(new_net_21157)
	);

	bfr new_net_21158_bfr_after (
		.din(new_net_21157),
		.dout(new_net_21158)
	);

	bfr new_net_21159_bfr_after (
		.din(new_net_21158),
		.dout(new_net_21159)
	);

	bfr new_net_21160_bfr_after (
		.din(new_net_21159),
		.dout(new_net_21160)
	);

	bfr new_net_21161_bfr_after (
		.din(new_net_21160),
		.dout(new_net_21161)
	);

	bfr new_net_21162_bfr_after (
		.din(new_net_21161),
		.dout(new_net_21162)
	);

	bfr new_net_21163_bfr_after (
		.din(new_net_21162),
		.dout(new_net_21163)
	);

	bfr new_net_21164_bfr_after (
		.din(new_net_21163),
		.dout(new_net_21164)
	);

	bfr new_net_21165_bfr_after (
		.din(new_net_21164),
		.dout(new_net_21165)
	);

	bfr new_net_21166_bfr_after (
		.din(new_net_21165),
		.dout(new_net_21166)
	);

	bfr new_net_21167_bfr_after (
		.din(new_net_21166),
		.dout(new_net_21167)
	);

	bfr new_net_21168_bfr_after (
		.din(new_net_21167),
		.dout(new_net_21168)
	);

	bfr new_net_21169_bfr_after (
		.din(new_net_21168),
		.dout(new_net_21169)
	);

	bfr new_net_21170_bfr_after (
		.din(new_net_21169),
		.dout(new_net_21170)
	);

	bfr new_net_21171_bfr_after (
		.din(new_net_21170),
		.dout(new_net_21171)
	);

	bfr new_net_21172_bfr_after (
		.din(new_net_21171),
		.dout(new_net_21172)
	);

	bfr new_net_21173_bfr_after (
		.din(new_net_21172),
		.dout(new_net_21173)
	);

	bfr new_net_21174_bfr_after (
		.din(new_net_21173),
		.dout(new_net_21174)
	);

	bfr new_net_21175_bfr_after (
		.din(new_net_21174),
		.dout(new_net_21175)
	);

	bfr new_net_21176_bfr_after (
		.din(new_net_21175),
		.dout(new_net_21176)
	);

	bfr new_net_21177_bfr_after (
		.din(new_net_21176),
		.dout(new_net_21177)
	);

	bfr new_net_21178_bfr_after (
		.din(new_net_21177),
		.dout(new_net_21178)
	);

	bfr new_net_21179_bfr_after (
		.din(new_net_21178),
		.dout(new_net_21179)
	);

	bfr new_net_21180_bfr_after (
		.din(new_net_21179),
		.dout(new_net_21180)
	);

	bfr new_net_21181_bfr_after (
		.din(new_net_21180),
		.dout(new_net_21181)
	);

	bfr new_net_21182_bfr_after (
		.din(new_net_21181),
		.dout(new_net_21182)
	);

	bfr new_net_21183_bfr_after (
		.din(new_net_21182),
		.dout(new_net_21183)
	);

	bfr new_net_21184_bfr_after (
		.din(new_net_21183),
		.dout(new_net_21184)
	);

	bfr new_net_21185_bfr_after (
		.din(new_net_21184),
		.dout(new_net_21185)
	);

	bfr new_net_21186_bfr_after (
		.din(new_net_21185),
		.dout(new_net_21186)
	);

	bfr N2548_bfr_after (
		.din(new_net_21186),
		.dout(N2548)
	);

	bfr new_net_3513_bfr_after (
		.din(_1149_),
		.dout(new_net_3513)
	);

	bfr new_net_3523_bfr_after (
		.din(_1179_),
		.dout(new_net_3523)
	);

	bfr new_net_3743_bfr_after (
		.din(_0267_),
		.dout(new_net_3743)
	);

	bfr new_net_3785_bfr_after (
		.din(_0456_),
		.dout(new_net_3785)
	);

	bfr new_net_21187_bfr_after (
		.din(new_net_3948),
		.dout(new_net_21187)
	);

	bfr new_net_21188_bfr_after (
		.din(new_net_21187),
		.dout(new_net_21188)
	);

	bfr new_net_21189_bfr_after (
		.din(new_net_21188),
		.dout(new_net_21189)
	);

	bfr new_net_21190_bfr_after (
		.din(new_net_21189),
		.dout(new_net_21190)
	);

	bfr new_net_21191_bfr_after (
		.din(new_net_21190),
		.dout(new_net_21191)
	);

	bfr new_net_21192_bfr_after (
		.din(new_net_21191),
		.dout(new_net_21192)
	);

	bfr new_net_21193_bfr_after (
		.din(new_net_21192),
		.dout(new_net_21193)
	);

	bfr new_net_21194_bfr_after (
		.din(new_net_21193),
		.dout(new_net_21194)
	);

	bfr new_net_21195_bfr_after (
		.din(new_net_21194),
		.dout(new_net_21195)
	);

	bfr new_net_21196_bfr_after (
		.din(new_net_21195),
		.dout(new_net_21196)
	);

	bfr new_net_21197_bfr_after (
		.din(new_net_21196),
		.dout(new_net_21197)
	);

	bfr N6260_bfr_after (
		.din(new_net_21197),
		.dout(N6260)
	);

	bfr new_net_3508_bfr_after (
		.din(_1116_),
		.dout(new_net_3508)
	);

	bfr new_net_3629_bfr_after (
		.din(_1604_),
		.dout(new_net_3629)
	);

	bfr new_net_3734_bfr_after (
		.din(_0208_),
		.dout(new_net_3734)
	);

	bfr new_net_3813_bfr_after (
		.din(_0571_),
		.dout(new_net_3813)
	);

	bfr new_net_3859_bfr_after (
		.din(_0760_),
		.dout(new_net_3859)
	);

	bfr new_net_3489_bfr_after (
		.din(_1043_),
		.dout(new_net_3489)
	);

	bfr new_net_3519_bfr_after (
		.din(_1167_),
		.dout(new_net_3519)
	);

	bfr new_net_3622_bfr_after (
		.din(_1552_),
		.dout(new_net_3622)
	);

	bfr new_net_3725_bfr_after (
		.din(_0178_),
		.dout(new_net_3725)
	);

	bfr new_net_3788_bfr_after (
		.din(_0466_),
		.dout(new_net_3788)
	);

	bfr new_net_21198_bfr_after (
		.din(new_net_3946),
		.dout(new_net_21198)
	);

	bfr new_net_21199_bfr_after (
		.din(new_net_21198),
		.dout(new_net_21199)
	);

	bfr new_net_21200_bfr_after (
		.din(new_net_21199),
		.dout(new_net_21200)
	);

	bfr new_net_21201_bfr_after (
		.din(new_net_21200),
		.dout(new_net_21201)
	);

	bfr new_net_21202_bfr_after (
		.din(new_net_21201),
		.dout(new_net_21202)
	);

	bfr new_net_21203_bfr_after (
		.din(new_net_21202),
		.dout(new_net_21203)
	);

	bfr new_net_21204_bfr_after (
		.din(new_net_21203),
		.dout(new_net_21204)
	);

	bfr new_net_21205_bfr_after (
		.din(new_net_21204),
		.dout(new_net_21205)
	);

	bfr new_net_21206_bfr_after (
		.din(new_net_21205),
		.dout(new_net_21206)
	);

	bfr new_net_21207_bfr_after (
		.din(new_net_21206),
		.dout(new_net_21207)
	);

	bfr new_net_21208_bfr_after (
		.din(new_net_21207),
		.dout(new_net_21208)
	);

	bfr new_net_21209_bfr_after (
		.din(new_net_21208),
		.dout(new_net_21209)
	);

	bfr new_net_21210_bfr_after (
		.din(new_net_21209),
		.dout(new_net_21210)
	);

	bfr new_net_21211_bfr_after (
		.din(new_net_21210),
		.dout(new_net_21211)
	);

	bfr new_net_21212_bfr_after (
		.din(new_net_21211),
		.dout(new_net_21212)
	);

	bfr new_net_21213_bfr_after (
		.din(new_net_21212),
		.dout(new_net_21213)
	);

	bfr new_net_21214_bfr_after (
		.din(new_net_21213),
		.dout(new_net_21214)
	);

	bfr new_net_21215_bfr_after (
		.din(new_net_21214),
		.dout(new_net_21215)
	);

	bfr new_net_21216_bfr_after (
		.din(new_net_21215),
		.dout(new_net_21216)
	);

	bfr new_net_21217_bfr_after (
		.din(new_net_21216),
		.dout(new_net_21217)
	);

	bfr new_net_21218_bfr_after (
		.din(new_net_21217),
		.dout(new_net_21218)
	);

	bfr new_net_21219_bfr_after (
		.din(new_net_21218),
		.dout(new_net_21219)
	);

	bfr new_net_21220_bfr_after (
		.din(new_net_21219),
		.dout(new_net_21220)
	);

	bfr N6230_bfr_after (
		.din(new_net_21220),
		.dout(N6230)
	);

	bfr new_net_21221_bfr_after (
		.din(_1195_),
		.dout(new_net_21221)
	);

	bfr new_net_3529_bfr_after (
		.din(new_net_21221),
		.dout(new_net_3529)
	);

	bfr new_net_3637_bfr_after (
		.din(_1630_),
		.dout(new_net_3637)
	);

	bfr new_net_3726_bfr_after (
		.din(_0181_),
		.dout(new_net_3726)
	);

	bfr new_net_3755_bfr_after (
		.din(_0306_),
		.dout(new_net_3755)
	);

	bfr new_net_3533_bfr_after (
		.din(_1199_),
		.dout(new_net_3533)
	);

	bfr new_net_3628_bfr_after (
		.din(_1601_),
		.dout(new_net_3628)
	);

	bfr new_net_3677_bfr_after (
		.din(_1795_),
		.dout(new_net_3677)
	);

	bfr new_net_3800_bfr_after (
		.din(_0506_),
		.dout(new_net_3800)
	);

	bfr new_net_3475_bfr_after (
		.din(_0632_),
		.dout(new_net_3475)
	);

	bfr new_net_3543_bfr_after (
		.din(_1241_),
		.dout(new_net_3543)
	);

	bfr new_net_3710_bfr_after (
		.din(_0128_),
		.dout(new_net_3710)
	);

	bfr new_net_3721_bfr_after (
		.din(_0164_),
		.dout(new_net_3721)
	);

	bfr new_net_3898_bfr_after (
		.din(_0938_),
		.dout(new_net_3898)
	);

	bfr new_net_3663_bfr_after (
		.din(_1749_),
		.dout(new_net_3663)
	);

	bfr new_net_3619_bfr_after (
		.din(_1543_),
		.dout(new_net_3619)
	);

	bfr new_net_3732_bfr_after (
		.din(_0201_),
		.dout(new_net_3732)
	);

	bfr new_net_3767_bfr_after (
		.din(_0373_),
		.dout(new_net_3767)
	);

	bfr new_net_21222_bfr_after (
		.din(new_net_3944),
		.dout(new_net_21222)
	);

	bfr new_net_21223_bfr_after (
		.din(new_net_21222),
		.dout(new_net_21223)
	);

	bfr new_net_21224_bfr_after (
		.din(new_net_21223),
		.dout(new_net_21224)
	);

	bfr new_net_21225_bfr_after (
		.din(new_net_21224),
		.dout(new_net_21225)
	);

	bfr new_net_21226_bfr_after (
		.din(new_net_21225),
		.dout(new_net_21226)
	);

	bfr new_net_21227_bfr_after (
		.din(new_net_21226),
		.dout(new_net_21227)
	);

	bfr new_net_21228_bfr_after (
		.din(new_net_21227),
		.dout(new_net_21228)
	);

	bfr new_net_21229_bfr_after (
		.din(new_net_21228),
		.dout(new_net_21229)
	);

	bfr new_net_21230_bfr_after (
		.din(new_net_21229),
		.dout(new_net_21230)
	);

	bfr new_net_21231_bfr_after (
		.din(new_net_21230),
		.dout(new_net_21231)
	);

	bfr new_net_21232_bfr_after (
		.din(new_net_21231),
		.dout(new_net_21232)
	);

	bfr new_net_21233_bfr_after (
		.din(new_net_21232),
		.dout(new_net_21233)
	);

	bfr new_net_21234_bfr_after (
		.din(new_net_21233),
		.dout(new_net_21234)
	);

	bfr new_net_21235_bfr_after (
		.din(new_net_21234),
		.dout(new_net_21235)
	);

	bfr new_net_21236_bfr_after (
		.din(new_net_21235),
		.dout(new_net_21236)
	);

	bfr new_net_21237_bfr_after (
		.din(new_net_21236),
		.dout(new_net_21237)
	);

	bfr new_net_21238_bfr_after (
		.din(new_net_21237),
		.dout(new_net_21238)
	);

	bfr new_net_21239_bfr_after (
		.din(new_net_21238),
		.dout(new_net_21239)
	);

	bfr new_net_21240_bfr_after (
		.din(new_net_21239),
		.dout(new_net_21240)
	);

	bfr new_net_21241_bfr_after (
		.din(new_net_21240),
		.dout(new_net_21241)
	);

	bfr new_net_21242_bfr_after (
		.din(new_net_21241),
		.dout(new_net_21242)
	);

	bfr new_net_21243_bfr_after (
		.din(new_net_21242),
		.dout(new_net_21243)
	);

	bfr new_net_21244_bfr_after (
		.din(new_net_21243),
		.dout(new_net_21244)
	);

	bfr new_net_21245_bfr_after (
		.din(new_net_21244),
		.dout(new_net_21245)
	);

	bfr new_net_21246_bfr_after (
		.din(new_net_21245),
		.dout(new_net_21246)
	);

	bfr new_net_21247_bfr_after (
		.din(new_net_21246),
		.dout(new_net_21247)
	);

	bfr new_net_21248_bfr_after (
		.din(new_net_21247),
		.dout(new_net_21248)
	);

	bfr new_net_21249_bfr_after (
		.din(new_net_21248),
		.dout(new_net_21249)
	);

	bfr new_net_21250_bfr_after (
		.din(new_net_21249),
		.dout(new_net_21250)
	);

	bfr new_net_21251_bfr_after (
		.din(new_net_21250),
		.dout(new_net_21251)
	);

	bfr new_net_21252_bfr_after (
		.din(new_net_21251),
		.dout(new_net_21252)
	);

	bfr N6210_bfr_after (
		.din(new_net_21252),
		.dout(N6210)
	);

	bfr new_net_3488_bfr_after (
		.din(_1040_),
		.dout(new_net_3488)
	);

	bfr new_net_3527_bfr_after (
		.din(_1191_),
		.dout(new_net_3527)
	);

	bfr new_net_3539_bfr_after (
		.din(_1229_),
		.dout(new_net_3539)
	);

	bfr new_net_3625_bfr_after (
		.din(_1591_),
		.dout(new_net_3625)
	);

	bfr new_net_3728_bfr_after (
		.din(_0188_),
		.dout(new_net_3728)
	);

	bfr new_net_3790_bfr_after (
		.din(_0473_),
		.dout(new_net_3790)
	);

	bfr new_net_3836_bfr_after (
		.din(_0667_),
		.dout(new_net_3836)
	);

	bfr new_net_3916_bfr_after (
		.din(_1011_),
		.dout(new_net_3916)
	);

	bfr new_net_3727_bfr_after (
		.din(_0184_),
		.dout(new_net_3727)
	);

	bfr new_net_3522_bfr_after (
		.din(_1176_),
		.dout(new_net_3522)
	);

	bfr new_net_3606_bfr_after (
		.din(_1500_),
		.dout(new_net_3606)
	);

	bfr new_net_3650_bfr_after (
		.din(_1673_),
		.dout(new_net_3650)
	);

	bfr new_net_21253_bfr_after (
		.din(new_net_3934),
		.dout(new_net_21253)
	);

	bfr new_net_21254_bfr_after (
		.din(new_net_21253),
		.dout(new_net_21254)
	);

	bfr new_net_21255_bfr_after (
		.din(new_net_21254),
		.dout(new_net_21255)
	);

	bfr new_net_21256_bfr_after (
		.din(new_net_21255),
		.dout(new_net_21256)
	);

	bfr new_net_21257_bfr_after (
		.din(new_net_21256),
		.dout(new_net_21257)
	);

	bfr new_net_21258_bfr_after (
		.din(new_net_21257),
		.dout(new_net_21258)
	);

	bfr new_net_21259_bfr_after (
		.din(new_net_21258),
		.dout(new_net_21259)
	);

	bfr new_net_21260_bfr_after (
		.din(new_net_21259),
		.dout(new_net_21260)
	);

	bfr new_net_21261_bfr_after (
		.din(new_net_21260),
		.dout(new_net_21261)
	);

	bfr new_net_21262_bfr_after (
		.din(new_net_21261),
		.dout(new_net_21262)
	);

	bfr new_net_21263_bfr_after (
		.din(new_net_21262),
		.dout(new_net_21263)
	);

	bfr new_net_21264_bfr_after (
		.din(new_net_21263),
		.dout(new_net_21264)
	);

	bfr new_net_21265_bfr_after (
		.din(new_net_21264),
		.dout(new_net_21265)
	);

	bfr new_net_21266_bfr_after (
		.din(new_net_21265),
		.dout(new_net_21266)
	);

	bfr new_net_21267_bfr_after (
		.din(new_net_21266),
		.dout(new_net_21267)
	);

	bfr new_net_21268_bfr_after (
		.din(new_net_21267),
		.dout(new_net_21268)
	);

	bfr new_net_21269_bfr_after (
		.din(new_net_21268),
		.dout(new_net_21269)
	);

	bfr new_net_21270_bfr_after (
		.din(new_net_21269),
		.dout(new_net_21270)
	);

	bfr new_net_21271_bfr_after (
		.din(new_net_21270),
		.dout(new_net_21271)
	);

	bfr new_net_21272_bfr_after (
		.din(new_net_21271),
		.dout(new_net_21272)
	);

	bfr new_net_21273_bfr_after (
		.din(new_net_21272),
		.dout(new_net_21273)
	);

	bfr new_net_21274_bfr_after (
		.din(new_net_21273),
		.dout(new_net_21274)
	);

	bfr new_net_21275_bfr_after (
		.din(new_net_21274),
		.dout(new_net_21275)
	);

	bfr new_net_21276_bfr_after (
		.din(new_net_21275),
		.dout(new_net_21276)
	);

	bfr new_net_21277_bfr_after (
		.din(new_net_21276),
		.dout(new_net_21277)
	);

	bfr new_net_21278_bfr_after (
		.din(new_net_21277),
		.dout(new_net_21278)
	);

	bfr new_net_21279_bfr_after (
		.din(new_net_21278),
		.dout(new_net_21279)
	);

	bfr new_net_21280_bfr_after (
		.din(new_net_21279),
		.dout(new_net_21280)
	);

	bfr new_net_21281_bfr_after (
		.din(new_net_21280),
		.dout(new_net_21281)
	);

	bfr new_net_21282_bfr_after (
		.din(new_net_21281),
		.dout(new_net_21282)
	);

	bfr new_net_21283_bfr_after (
		.din(new_net_21282),
		.dout(new_net_21283)
	);

	bfr new_net_21284_bfr_after (
		.din(new_net_21283),
		.dout(new_net_21284)
	);

	bfr new_net_21285_bfr_after (
		.din(new_net_21284),
		.dout(new_net_21285)
	);

	bfr new_net_21286_bfr_after (
		.din(new_net_21285),
		.dout(new_net_21286)
	);

	bfr new_net_21287_bfr_after (
		.din(new_net_21286),
		.dout(new_net_21287)
	);

	bfr new_net_21288_bfr_after (
		.din(new_net_21287),
		.dout(new_net_21288)
	);

	bfr new_net_21289_bfr_after (
		.din(new_net_21288),
		.dout(new_net_21289)
	);

	bfr new_net_21290_bfr_after (
		.din(new_net_21289),
		.dout(new_net_21290)
	);

	bfr new_net_21291_bfr_after (
		.din(new_net_21290),
		.dout(new_net_21291)
	);

	bfr new_net_21292_bfr_after (
		.din(new_net_21291),
		.dout(new_net_21292)
	);

	bfr new_net_21293_bfr_after (
		.din(new_net_21292),
		.dout(new_net_21293)
	);

	bfr new_net_21294_bfr_after (
		.din(new_net_21293),
		.dout(new_net_21294)
	);

	bfr new_net_21295_bfr_after (
		.din(new_net_21294),
		.dout(new_net_21295)
	);

	bfr N6180_bfr_after (
		.din(new_net_21295),
		.dout(N6180)
	);

	bfr new_net_3613_bfr_after (
		.din(_1523_),
		.dout(new_net_3613)
	);

	bfr new_net_3752_bfr_after (
		.din(_0297_),
		.dout(new_net_3752)
	);

	bfr new_net_3786_bfr_after (
		.din(_0460_),
		.dout(new_net_3786)
	);

	bfr new_net_3709_bfr_after (
		.din(_0125_),
		.dout(new_net_3709)
	);

	bfr new_net_3467_bfr_after (
		.din(_0252_),
		.dout(new_net_3467)
	);

	bfr new_net_3572_bfr_after (
		.din(_1348_),
		.dout(new_net_3572)
	);

	bfr new_net_3591_bfr_after (
		.din(_1427_),
		.dout(new_net_3591)
	);

	bfr new_net_3634_bfr_after (
		.din(_1620_),
		.dout(new_net_3634)
	);

	bfr new_net_3834_bfr_after (
		.din(_0660_),
		.dout(new_net_3834)
	);

	bfr new_net_3904_bfr_after (
		.din(_0957_),
		.dout(new_net_3904)
	);

	bfr new_net_3718_bfr_after (
		.din(_0155_),
		.dout(new_net_3718)
	);

	bfr new_net_3603_bfr_after (
		.din(_1490_),
		.dout(new_net_3603)
	);

	bfr new_net_3647_bfr_after (
		.din(_1663_),
		.dout(new_net_3647)
	);

	bfr new_net_3890_bfr_after (
		.din(_0902_),
		.dout(new_net_3890)
	);

	bfr new_net_21296_bfr_after (
		.din(new_net_3920),
		.dout(new_net_21296)
	);

	bfr new_net_21297_bfr_after (
		.din(new_net_21296),
		.dout(new_net_21297)
	);

	bfr new_net_21298_bfr_after (
		.din(new_net_21297),
		.dout(new_net_21298)
	);

	bfr new_net_21299_bfr_after (
		.din(new_net_21298),
		.dout(new_net_21299)
	);

	bfr new_net_21300_bfr_after (
		.din(new_net_21299),
		.dout(new_net_21300)
	);

	bfr new_net_21301_bfr_after (
		.din(new_net_21300),
		.dout(new_net_21301)
	);

	bfr new_net_21302_bfr_after (
		.din(new_net_21301),
		.dout(new_net_21302)
	);

	bfr new_net_21303_bfr_after (
		.din(new_net_21302),
		.dout(new_net_21303)
	);

	bfr new_net_21304_bfr_after (
		.din(new_net_21303),
		.dout(new_net_21304)
	);

	bfr new_net_21305_bfr_after (
		.din(new_net_21304),
		.dout(new_net_21305)
	);

	bfr new_net_21306_bfr_after (
		.din(new_net_21305),
		.dout(new_net_21306)
	);

	bfr new_net_21307_bfr_after (
		.din(new_net_21306),
		.dout(new_net_21307)
	);

	bfr new_net_21308_bfr_after (
		.din(new_net_21307),
		.dout(new_net_21308)
	);

	bfr new_net_21309_bfr_after (
		.din(new_net_21308),
		.dout(new_net_21309)
	);

	bfr new_net_21310_bfr_after (
		.din(new_net_21309),
		.dout(new_net_21310)
	);

	bfr new_net_21311_bfr_after (
		.din(new_net_21310),
		.dout(new_net_21311)
	);

	bfr new_net_21312_bfr_after (
		.din(new_net_21311),
		.dout(new_net_21312)
	);

	bfr new_net_21313_bfr_after (
		.din(new_net_21312),
		.dout(new_net_21313)
	);

	bfr new_net_21314_bfr_after (
		.din(new_net_21313),
		.dout(new_net_21314)
	);

	bfr new_net_21315_bfr_after (
		.din(new_net_21314),
		.dout(new_net_21315)
	);

	bfr new_net_21316_bfr_after (
		.din(new_net_21315),
		.dout(new_net_21316)
	);

	bfr new_net_21317_bfr_after (
		.din(new_net_21316),
		.dout(new_net_21317)
	);

	bfr new_net_21318_bfr_after (
		.din(new_net_21317),
		.dout(new_net_21318)
	);

	bfr new_net_21319_bfr_after (
		.din(new_net_21318),
		.dout(new_net_21319)
	);

	bfr new_net_21320_bfr_after (
		.din(new_net_21319),
		.dout(new_net_21320)
	);

	bfr new_net_21321_bfr_after (
		.din(new_net_21320),
		.dout(new_net_21321)
	);

	bfr new_net_21322_bfr_after (
		.din(new_net_21321),
		.dout(new_net_21322)
	);

	bfr new_net_21323_bfr_after (
		.din(new_net_21322),
		.dout(new_net_21323)
	);

	bfr new_net_21324_bfr_after (
		.din(new_net_21323),
		.dout(new_net_21324)
	);

	bfr new_net_21325_bfr_after (
		.din(new_net_21324),
		.dout(new_net_21325)
	);

	bfr new_net_21326_bfr_after (
		.din(new_net_21325),
		.dout(new_net_21326)
	);

	bfr new_net_21327_bfr_after (
		.din(new_net_21326),
		.dout(new_net_21327)
	);

	bfr new_net_21328_bfr_after (
		.din(new_net_21327),
		.dout(new_net_21328)
	);

	bfr new_net_21329_bfr_after (
		.din(new_net_21328),
		.dout(new_net_21329)
	);

	bfr new_net_21330_bfr_after (
		.din(new_net_21329),
		.dout(new_net_21330)
	);

	bfr new_net_21331_bfr_after (
		.din(new_net_21330),
		.dout(new_net_21331)
	);

	bfr new_net_21332_bfr_after (
		.din(new_net_21331),
		.dout(new_net_21332)
	);

	bfr new_net_21333_bfr_after (
		.din(new_net_21332),
		.dout(new_net_21333)
	);

	bfr new_net_21334_bfr_after (
		.din(new_net_21333),
		.dout(new_net_21334)
	);

	bfr new_net_21335_bfr_after (
		.din(new_net_21334),
		.dout(new_net_21335)
	);

	bfr new_net_21336_bfr_after (
		.din(new_net_21335),
		.dout(new_net_21336)
	);

	bfr new_net_21337_bfr_after (
		.din(new_net_21336),
		.dout(new_net_21337)
	);

	bfr new_net_21338_bfr_after (
		.din(new_net_21337),
		.dout(new_net_21338)
	);

	bfr new_net_21339_bfr_after (
		.din(new_net_21338),
		.dout(new_net_21339)
	);

	bfr new_net_21340_bfr_after (
		.din(new_net_21339),
		.dout(new_net_21340)
	);

	bfr new_net_21341_bfr_after (
		.din(new_net_21340),
		.dout(new_net_21341)
	);

	bfr new_net_21342_bfr_after (
		.din(new_net_21341),
		.dout(new_net_21342)
	);

	bfr new_net_21343_bfr_after (
		.din(new_net_21342),
		.dout(new_net_21343)
	);

	bfr new_net_21344_bfr_after (
		.din(new_net_21343),
		.dout(new_net_21344)
	);

	bfr new_net_21345_bfr_after (
		.din(new_net_21344),
		.dout(new_net_21345)
	);

	bfr new_net_21346_bfr_after (
		.din(new_net_21345),
		.dout(new_net_21346)
	);

	bfr new_net_21347_bfr_after (
		.din(new_net_21346),
		.dout(new_net_21347)
	);

	bfr new_net_21348_bfr_after (
		.din(new_net_21347),
		.dout(new_net_21348)
	);

	bfr new_net_21349_bfr_after (
		.din(new_net_21348),
		.dout(new_net_21349)
	);

	bfr new_net_21350_bfr_after (
		.din(new_net_21349),
		.dout(new_net_21350)
	);

	bfr new_net_21351_bfr_after (
		.din(new_net_21350),
		.dout(new_net_21351)
	);

	bfr new_net_21352_bfr_after (
		.din(new_net_21351),
		.dout(new_net_21352)
	);

	bfr new_net_21353_bfr_after (
		.din(new_net_21352),
		.dout(new_net_21353)
	);

	bfr new_net_21354_bfr_after (
		.din(new_net_21353),
		.dout(new_net_21354)
	);

	bfr N6123_bfr_after (
		.din(new_net_21354),
		.dout(N6123)
	);

	bfr new_net_3763_bfr_after (
		.din(_0359_),
		.dout(new_net_3763)
	);

	bfr new_net_3884_bfr_after (
		.din(_0871_),
		.dout(new_net_3884)
	);

	bfr new_net_21355_bfr_after (
		.din(new_net_3932),
		.dout(new_net_21355)
	);

	bfr new_net_21356_bfr_after (
		.din(new_net_21355),
		.dout(new_net_21356)
	);

	bfr new_net_21357_bfr_after (
		.din(new_net_21356),
		.dout(new_net_21357)
	);

	bfr new_net_21358_bfr_after (
		.din(new_net_21357),
		.dout(new_net_21358)
	);

	bfr new_net_21359_bfr_after (
		.din(new_net_21358),
		.dout(new_net_21359)
	);

	bfr new_net_21360_bfr_after (
		.din(new_net_21359),
		.dout(new_net_21360)
	);

	bfr new_net_21361_bfr_after (
		.din(new_net_21360),
		.dout(new_net_21361)
	);

	bfr new_net_21362_bfr_after (
		.din(new_net_21361),
		.dout(new_net_21362)
	);

	bfr new_net_21363_bfr_after (
		.din(new_net_21362),
		.dout(new_net_21363)
	);

	bfr new_net_21364_bfr_after (
		.din(new_net_21363),
		.dout(new_net_21364)
	);

	bfr new_net_21365_bfr_after (
		.din(new_net_21364),
		.dout(new_net_21365)
	);

	bfr new_net_21366_bfr_after (
		.din(new_net_21365),
		.dout(new_net_21366)
	);

	bfr new_net_21367_bfr_after (
		.din(new_net_21366),
		.dout(new_net_21367)
	);

	bfr new_net_21368_bfr_after (
		.din(new_net_21367),
		.dout(new_net_21368)
	);

	bfr new_net_21369_bfr_after (
		.din(new_net_21368),
		.dout(new_net_21369)
	);

	bfr new_net_21370_bfr_after (
		.din(new_net_21369),
		.dout(new_net_21370)
	);

	bfr new_net_21371_bfr_after (
		.din(new_net_21370),
		.dout(new_net_21371)
	);

	bfr new_net_21372_bfr_after (
		.din(new_net_21371),
		.dout(new_net_21372)
	);

	bfr new_net_21373_bfr_after (
		.din(new_net_21372),
		.dout(new_net_21373)
	);

	bfr new_net_21374_bfr_after (
		.din(new_net_21373),
		.dout(new_net_21374)
	);

	bfr new_net_21375_bfr_after (
		.din(new_net_21374),
		.dout(new_net_21375)
	);

	bfr new_net_21376_bfr_after (
		.din(new_net_21375),
		.dout(new_net_21376)
	);

	bfr new_net_21377_bfr_after (
		.din(new_net_21376),
		.dout(new_net_21377)
	);

	bfr new_net_21378_bfr_after (
		.din(new_net_21377),
		.dout(new_net_21378)
	);

	bfr new_net_21379_bfr_after (
		.din(new_net_21378),
		.dout(new_net_21379)
	);

	bfr new_net_21380_bfr_after (
		.din(new_net_21379),
		.dout(new_net_21380)
	);

	bfr new_net_21381_bfr_after (
		.din(new_net_21380),
		.dout(new_net_21381)
	);

	bfr new_net_21382_bfr_after (
		.din(new_net_21381),
		.dout(new_net_21382)
	);

	bfr new_net_21383_bfr_after (
		.din(new_net_21382),
		.dout(new_net_21383)
	);

	bfr new_net_21384_bfr_after (
		.din(new_net_21383),
		.dout(new_net_21384)
	);

	bfr new_net_21385_bfr_after (
		.din(new_net_21384),
		.dout(new_net_21385)
	);

	bfr new_net_21386_bfr_after (
		.din(new_net_21385),
		.dout(new_net_21386)
	);

	bfr new_net_21387_bfr_after (
		.din(new_net_21386),
		.dout(new_net_21387)
	);

	bfr new_net_21388_bfr_after (
		.din(new_net_21387),
		.dout(new_net_21388)
	);

	bfr new_net_21389_bfr_after (
		.din(new_net_21388),
		.dout(new_net_21389)
	);

	bfr new_net_21390_bfr_after (
		.din(new_net_21389),
		.dout(new_net_21390)
	);

	bfr new_net_21391_bfr_after (
		.din(new_net_21390),
		.dout(new_net_21391)
	);

	bfr new_net_21392_bfr_after (
		.din(new_net_21391),
		.dout(new_net_21392)
	);

	bfr new_net_21393_bfr_after (
		.din(new_net_21392),
		.dout(new_net_21393)
	);

	bfr new_net_21394_bfr_after (
		.din(new_net_21393),
		.dout(new_net_21394)
	);

	bfr new_net_21395_bfr_after (
		.din(new_net_21394),
		.dout(new_net_21395)
	);

	bfr new_net_21396_bfr_after (
		.din(new_net_21395),
		.dout(new_net_21396)
	);

	bfr new_net_21397_bfr_after (
		.din(new_net_21396),
		.dout(new_net_21397)
	);

	bfr new_net_21398_bfr_after (
		.din(new_net_21397),
		.dout(new_net_21398)
	);

	bfr new_net_21399_bfr_after (
		.din(new_net_21398),
		.dout(new_net_21399)
	);

	bfr new_net_21400_bfr_after (
		.din(new_net_21399),
		.dout(new_net_21400)
	);

	bfr new_net_21401_bfr_after (
		.din(new_net_21400),
		.dout(new_net_21401)
	);

	bfr new_net_21402_bfr_after (
		.din(new_net_21401),
		.dout(new_net_21402)
	);

	bfr new_net_21403_bfr_after (
		.din(new_net_21402),
		.dout(new_net_21403)
	);

	bfr new_net_21404_bfr_after (
		.din(new_net_21403),
		.dout(new_net_21404)
	);

	bfr new_net_21405_bfr_after (
		.din(new_net_21404),
		.dout(new_net_21405)
	);

	bfr new_net_21406_bfr_after (
		.din(new_net_21405),
		.dout(new_net_21406)
	);

	bfr new_net_21407_bfr_after (
		.din(new_net_21406),
		.dout(new_net_21407)
	);

	bfr new_net_21408_bfr_after (
		.din(new_net_21407),
		.dout(new_net_21408)
	);

	bfr new_net_21409_bfr_after (
		.din(new_net_21408),
		.dout(new_net_21409)
	);

	bfr new_net_21410_bfr_after (
		.din(new_net_21409),
		.dout(new_net_21410)
	);

	bfr new_net_21411_bfr_after (
		.din(new_net_21410),
		.dout(new_net_21411)
	);

	bfr new_net_21412_bfr_after (
		.din(new_net_21411),
		.dout(new_net_21412)
	);

	bfr new_net_21413_bfr_after (
		.din(new_net_21412),
		.dout(new_net_21413)
	);

	bfr new_net_21414_bfr_after (
		.din(new_net_21413),
		.dout(new_net_21414)
	);

	bfr new_net_21415_bfr_after (
		.din(new_net_21414),
		.dout(new_net_21415)
	);

	bfr new_net_21416_bfr_after (
		.din(new_net_21415),
		.dout(new_net_21416)
	);

	bfr new_net_21417_bfr_after (
		.din(new_net_21416),
		.dout(new_net_21417)
	);

	bfr new_net_21418_bfr_after (
		.din(new_net_21417),
		.dout(new_net_21418)
	);

	bfr new_net_21419_bfr_after (
		.din(new_net_21418),
		.dout(new_net_21419)
	);

	bfr new_net_21420_bfr_after (
		.din(new_net_21419),
		.dout(new_net_21420)
	);

	bfr new_net_21421_bfr_after (
		.din(new_net_21420),
		.dout(new_net_21421)
	);

	bfr new_net_21422_bfr_after (
		.din(new_net_21421),
		.dout(new_net_21422)
	);

	bfr new_net_21423_bfr_after (
		.din(new_net_21422),
		.dout(new_net_21423)
	);

	bfr new_net_21424_bfr_after (
		.din(new_net_21423),
		.dout(new_net_21424)
	);

	bfr new_net_21425_bfr_after (
		.din(new_net_21424),
		.dout(new_net_21425)
	);

	bfr new_net_21426_bfr_after (
		.din(new_net_21425),
		.dout(new_net_21426)
	);

	bfr new_net_21427_bfr_after (
		.din(new_net_21426),
		.dout(new_net_21427)
	);

	bfr new_net_21428_bfr_after (
		.din(new_net_21427),
		.dout(new_net_21428)
	);

	bfr new_net_21429_bfr_after (
		.din(new_net_21428),
		.dout(new_net_21429)
	);

	bfr new_net_21430_bfr_after (
		.din(new_net_21429),
		.dout(new_net_21430)
	);

	bfr new_net_21431_bfr_after (
		.din(new_net_21430),
		.dout(new_net_21431)
	);

	bfr new_net_21432_bfr_after (
		.din(new_net_21431),
		.dout(new_net_21432)
	);

	bfr new_net_21433_bfr_after (
		.din(new_net_21432),
		.dout(new_net_21433)
	);

	bfr new_net_21434_bfr_after (
		.din(new_net_21433),
		.dout(new_net_21434)
	);

	bfr new_net_21435_bfr_after (
		.din(new_net_21434),
		.dout(new_net_21435)
	);

	bfr new_net_21436_bfr_after (
		.din(new_net_21435),
		.dout(new_net_21436)
	);

	bfr new_net_21437_bfr_after (
		.din(new_net_21436),
		.dout(new_net_21437)
	);

	bfr new_net_21438_bfr_after (
		.din(new_net_21437),
		.dout(new_net_21438)
	);

	bfr new_net_21439_bfr_after (
		.din(new_net_21438),
		.dout(new_net_21439)
	);

	bfr new_net_21440_bfr_after (
		.din(new_net_21439),
		.dout(new_net_21440)
	);

	bfr new_net_21441_bfr_after (
		.din(new_net_21440),
		.dout(new_net_21441)
	);

	bfr new_net_21442_bfr_after (
		.din(new_net_21441),
		.dout(new_net_21442)
	);

	bfr new_net_21443_bfr_after (
		.din(new_net_21442),
		.dout(new_net_21443)
	);

	bfr new_net_21444_bfr_after (
		.din(new_net_21443),
		.dout(new_net_21444)
	);

	bfr new_net_21445_bfr_after (
		.din(new_net_21444),
		.dout(new_net_21445)
	);

	bfr new_net_21446_bfr_after (
		.din(new_net_21445),
		.dout(new_net_21446)
	);

	bfr new_net_21447_bfr_after (
		.din(new_net_21446),
		.dout(new_net_21447)
	);

	bfr new_net_21448_bfr_after (
		.din(new_net_21447),
		.dout(new_net_21448)
	);

	bfr new_net_21449_bfr_after (
		.din(new_net_21448),
		.dout(new_net_21449)
	);

	bfr new_net_21450_bfr_after (
		.din(new_net_21449),
		.dout(new_net_21450)
	);

	bfr new_net_21451_bfr_after (
		.din(new_net_21450),
		.dout(new_net_21451)
	);

	bfr new_net_21452_bfr_after (
		.din(new_net_21451),
		.dout(new_net_21452)
	);

	bfr new_net_21453_bfr_after (
		.din(new_net_21452),
		.dout(new_net_21453)
	);

	bfr new_net_21454_bfr_after (
		.din(new_net_21453),
		.dout(new_net_21454)
	);

	bfr new_net_21455_bfr_after (
		.din(new_net_21454),
		.dout(new_net_21455)
	);

	bfr new_net_21456_bfr_after (
		.din(new_net_21455),
		.dout(new_net_21456)
	);

	bfr new_net_21457_bfr_after (
		.din(new_net_21456),
		.dout(new_net_21457)
	);

	bfr new_net_21458_bfr_after (
		.din(new_net_21457),
		.dout(new_net_21458)
	);

	bfr new_net_21459_bfr_after (
		.din(new_net_21458),
		.dout(new_net_21459)
	);

	bfr new_net_21460_bfr_after (
		.din(new_net_21459),
		.dout(new_net_21460)
	);

	bfr new_net_21461_bfr_after (
		.din(new_net_21460),
		.dout(new_net_21461)
	);

	bfr new_net_21462_bfr_after (
		.din(new_net_21461),
		.dout(new_net_21462)
	);

	bfr new_net_21463_bfr_after (
		.din(new_net_21462),
		.dout(new_net_21463)
	);

	bfr new_net_21464_bfr_after (
		.din(new_net_21463),
		.dout(new_net_21464)
	);

	bfr new_net_21465_bfr_after (
		.din(new_net_21464),
		.dout(new_net_21465)
	);

	bfr new_net_21466_bfr_after (
		.din(new_net_21465),
		.dout(new_net_21466)
	);

	bfr new_net_21467_bfr_after (
		.din(new_net_21466),
		.dout(new_net_21467)
	);

	bfr new_net_21468_bfr_after (
		.din(new_net_21467),
		.dout(new_net_21468)
	);

	bfr new_net_21469_bfr_after (
		.din(new_net_21468),
		.dout(new_net_21469)
	);

	bfr new_net_21470_bfr_after (
		.din(new_net_21469),
		.dout(new_net_21470)
	);

	bfr new_net_21471_bfr_after (
		.din(new_net_21470),
		.dout(new_net_21471)
	);

	bfr new_net_21472_bfr_after (
		.din(new_net_21471),
		.dout(new_net_21472)
	);

	bfr new_net_21473_bfr_after (
		.din(new_net_21472),
		.dout(new_net_21473)
	);

	bfr new_net_21474_bfr_after (
		.din(new_net_21473),
		.dout(new_net_21474)
	);

	bfr new_net_21475_bfr_after (
		.din(new_net_21474),
		.dout(new_net_21475)
	);

	bfr new_net_21476_bfr_after (
		.din(new_net_21475),
		.dout(new_net_21476)
	);

	bfr new_net_21477_bfr_after (
		.din(new_net_21476),
		.dout(new_net_21477)
	);

	bfr N3552_bfr_after (
		.din(new_net_21477),
		.dout(N3552)
	);

	bfr new_net_3578_bfr_after (
		.din(_1388_),
		.dout(new_net_3578)
	);

	bfr new_net_3633_bfr_after (
		.din(_1617_),
		.dout(new_net_3633)
	);

	bfr new_net_3701_bfr_after (
		.din(_0065_),
		.dout(new_net_3701)
	);

	bfr new_net_3852_bfr_after (
		.din(_0737_),
		.dout(new_net_3852)
	);

	bfr new_net_3876_bfr_after (
		.din(_0845_),
		.dout(new_net_3876)
	);

	bfr new_net_3885_bfr_after (
		.din(_0875_),
		.dout(new_net_3885)
	);

	bfr new_net_3746_bfr_after (
		.din(_0277_),
		.dout(new_net_3746)
	);

	bfr new_net_3486_bfr_after (
		.din(_1034_),
		.dout(new_net_3486)
	);

	bfr new_net_3498_bfr_after (
		.din(_1086_),
		.dout(new_net_3498)
	);

	bfr new_net_3787_bfr_after (
		.din(_0463_),
		.dout(new_net_3787)
	);

	bfr new_net_3877_bfr_after (
		.din(_0848_),
		.dout(new_net_3877)
	);

	bfr new_net_3881_bfr_after (
		.din(_0862_),
		.dout(new_net_3881)
	);

endmodule