module c7552(N1, N5, N9, N12, N15, N18, N23, N26, N29, N32, N35, N38, N41, N44, N47, N50, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N69, N70, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N94, N97, N100, N103, N106, N109, N110, N111, N112, N113, N114, N115, N118, N121, N124, N127, N130, N133, N134, N135, N138, N141, N144, N147, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N242, N245, N248, N251, N254, N257, N260, N263, N267, N271, N274, N277, N280, N283, N286, N289, N293, N296, N299, N303, N307, N310, N313, N316, N319, N322, N325, N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N358, N361, N364, N367, N382, N241_I, N387, N388, N478, N482, N484, N486, N489, N492, N501, N505, N507, N509, N511, N513, N515, N517, N519, N535, N537, N539, N541, N543, N545, N547, N549, N551, N553, N556, N559, N561, N563, N565, N567, N569, N571, N573, N582, N643, N707, N813, N881, N882, N883, N884, N885, N889, N945, N1110, N1111, N1112, N1113, N1114, N1489, N1490, N1781, N10025, N10101, N10102, N10103, N10104, N10109, N10110, N10111, N10112, N10350, N10351, N10352, N10353, N10574, N10575, N10576, N10628, N10632, N10641, N10704, N10706, N10711, N10712, N10713, N10714, N10715, N10716, N10717, N10718, N10729, N10759, N10760, N10761, N10762, N10763, N10827, N10837, N10838, N10839, N10840, N10868, N10869, N10870, N10871, N10905, N10906, N10907, N10908, N11333, N11334, N11340, N11342, N241_O);
	wire new_net_6599;
	wire new_net_10260;
	wire new_net_6689;
	wire new_net_7351;
	wire new_net_8888;
	wire new_net_6561;
	wire new_net_9090;
	wire new_net_7400;
	wire new_net_8712;
	wire new_net_9247;
	wire n_0009_;
	wire n_0219_;
	wire n_0723_;
	wire n_1227_;
	wire new_net_2999;
	wire new_net_1365;
	wire new_net_1629;
	wire new_net_6208;
	wire new_net_6776;
	wire new_net_8139;
	wire new_net_4318;
	wire new_net_8156;
	wire new_net_9134;
	wire new_net_9644;
	wire new_net_7252;
	wire new_net_9821;
	wire new_net_4412;
	wire new_net_7859;
	wire new_net_8769;
	wire new_net_6466;
	wire new_net_771;
	wire new_net_2937;
	wire new_net_5061;
	wire new_net_5291;
	wire new_net_6005;
	wire new_net_5093;
	wire new_net_7642;
	wire new_net_7666;
	wire new_net_7805;
	wire new_net_7994;
	wire new_net_5710;
	wire new_net_8289;
	wire new_net_9547;
	wire new_net_7801;
	wire new_net_7977;
	wire new_net_7970;
	wire new_net_9871;
	wire new_net_9195;
	wire new_net_4434;
	wire n_0010_;
	wire n_0220_;
	wire n_0724_;
	wire n_1228_;
	wire new_net_1742;
	wire new_net_3564;
	wire new_net_952;
	wire new_net_2871;
	wire new_net_3793;
	wire new_net_4125;
	wire new_net_5584;
	wire new_net_6411;
	wire new_net_7439;
	wire new_net_8784;
	wire new_net_5974;
	wire new_net_6752;
	wire new_net_10599;
	wire new_net_2417;
	wire new_net_86;
	wire new_net_1251;
	wire new_net_1398;
	wire new_net_1890;
	wire new_net_3885;
	wire new_net_3932;
	wire new_net_4392;
	wire new_net_4513;
	wire new_net_5099;
	wire new_net_9217;
	wire new_net_9424;
	wire new_net_10683;
	wire new_net_8693;
	wire new_net_7303;
	wire n_1042_;
	wire n_0011_;
	wire n_0221_;
	wire n_0725_;
	wire new_net_2146;
	wire n_1229_;
	wire new_net_3204;
	wire new_net_4301;
	wire new_net_6103;
	wire new_net_6977;
	wire new_net_7001;
	wire new_net_6940;
	wire new_net_10145;
	wire new_net_7521;
	wire new_net_4014;
	wire new_net_7519;
	wire new_net_5514;
	wire new_net_9608;
	wire new_net_10307;
	wire new_net_7031;
	wire new_net_9606;
	wire new_net_8643;
	wire new_net_772;
	wire new_net_1217;
	wire new_net_3630;
	wire new_net_3585;
	wire new_net_4070;
	wire new_net_4327;
	wire new_net_5081;
	wire new_net_5856;
	wire new_net_6712;
	wire new_net_6795;
	wire new_net_10053;
	wire new_net_6585;
	wire new_net_10210;
	wire new_net_7541;
	wire new_net_8833;
	wire n_0222_;
	wire n_0012_;
	wire n_0726_;
	wire n_1230_;
	wire new_net_1743;
	wire new_net_953;
	wire new_net_3794;
	wire new_net_4348;
	wire new_net_4867;
	wire new_net_9178;
	wire new_net_7887;
	wire new_net_8251;
	wire new_net_7391;
	wire new_net_8703;
	wire new_net_10467;
	wire new_net_2065;
	wire new_net_1252;
	wire new_net_1366;
	wire new_net_1399;
	wire new_net_1630;
	wire new_net_3000;
	wire new_net_6777;
	wire new_net_8140;
	wire new_net_8687;
	wire new_net_9057;
	wire new_net_10389;
	wire new_net_9920;
	wire new_net_6353;
	wire new_net_10440;
	wire new_net_4111;
	wire new_net_6452;
	wire new_net_8437;
	wire new_net_10519;
	wire n_0727_;
	wire n_0223_;
	wire n_0013_;
	wire new_net_2938;
	wire n_1231_;
	wire new_net_3205;
	wire new_net_5062;
	wire new_net_5292;
	wire new_net_6006;
	wire new_net_7643;
	wire new_net_8608;
	wire new_net_9142;
	wire new_net_8804;
	wire new_net_10328;
	wire new_net_3852;
	wire new_net_5741;
	wire new_net_5570;
	wire new_net_9118;
	wire new_net_773;
	wire new_net_1218;
	wire new_net_2872;
	wire new_net_3565;
	wire new_net_4126;
	wire new_net_4885;
	wire new_net_5857;
	wire new_net_6630;
	wire new_net_6961;
	wire new_net_7058;
	wire new_net_9164;
	wire new_net_4724;
	wire new_net_4390;
	wire new_net_10348;
	wire new_net_7149;
	wire new_net_9717;
	wire new_net_5215;
	wire n_0014_;
	wire n_0224_;
	wire n_0728_;
	wire new_net_7;
	wire new_net_1891;
	wire n_1232_;
	wire new_net_87;
	wire new_net_1744;
	wire new_net_3886;
	wire new_net_3933;
	wire new_net_10674;
	wire new_net_6540;
	wire new_net_10013;
	wire new_net_7664;
	wire new_net_5005;
	wire new_net_6149;
	wire new_net_1727;
	wire new_net_1367;
	wire new_net_1400;
	wire new_net_1631;
	wire new_net_2418;
	wire new_net_4470;
	wire new_net_6104;
	wire new_net_6978;
	wire new_net_7002;
	wire new_net_7121;
	wire new_net_7145;
	wire new_net_10254;
	wire new_net_6926;
	wire new_net_10421;
	wire new_net_6473;
	wire n_1223_;
	wire new_net_8629;
	wire new_net_3586;
	wire n_0015_;
	wire n_0225_;
	wire n_0729_;
	wire new_net_2958;
	wire n_1233_;
	wire new_net_3631;
	wire new_net_4328;
	wire new_net_5082;
	wire new_net_6713;
	wire new_net_9022;
	wire new_net_5559;
	wire new_net_9020;
	wire new_net_9290;
	wire new_net_9974;
	wire new_net_7701;
	wire new_net_954;
	wire new_net_1219;
	wire new_net_3795;
	wire new_net_4349;
	wire new_net_4868;
	wire new_net_8461;
	wire new_net_9074;
	wire new_net_10075;
	wire new_net_10660;
	wire new_net_5602;
	wire new_net_5819;
	wire new_net_9042;
	wire n_1043_;
	wire new_net_8493;
	wire new_net_9749;
	wire new_net_9474;
	wire n_0226_;
	wire n_0016_;
	wire n_0730_;
	wire new_net_1892;
	wire new_net_1253;
	wire n_1234_;
	wire new_net_88;
	wire new_net_3001;
	wire new_net_6778;
	wire new_net_8141;
	wire new_net_8013;
	wire new_net_4396;
	wire new_net_6232;
	wire new_net_8462;
	wire new_net_8067;
	wire new_net_3964;
	wire new_net_8423;
	wire new_net_8348;
	wire new_net_8981;
	wire new_net_3206;
	wire new_net_2939;
	wire new_net_2676;
	wire new_net_4471;
	wire new_net_5063;
	wire new_net_5293;
	wire new_net_5388;
	wire new_net_6007;
	wire new_net_6621;
	wire new_net_7644;
	wire new_net_8858;
	wire new_net_9771;
	wire new_net_6286;
	wire new_net_8322;
	wire new_net_6097;
	wire new_net_10168;
	wire new_net_8320;
	wire new_net_9179;
	wire new_net_9109;
	wire new_net_3183;
	wire new_net_3566;
	wire n_0731_;
	wire n_0227_;
	wire n_0017_;
	wire new_net_2873;
	wire new_net_774;
	wire n_1235_;
	wire new_net_4127;
	wire new_net_4886;
	wire new_net_7049;
	wire new_net_5328;
	wire new_net_4091;
	wire new_net_5326;
	wire new_net_4978;
	wire new_net_6437;
	wire new_net_6729;
	wire new_net_955;
	wire new_net_1745;
	wire new_net_3887;
	wire new_net_3934;
	wire new_net_4515;
	wire new_net_2978;
	wire new_net_5101;
	wire new_net_5117;
	wire new_net_6185;
	wire new_net_6526;
	wire new_net_8851;
	wire new_net_9949;
	wire n_0732_;
	wire n_0228_;
	wire n_0018_;
	wire new_net_1368;
	wire new_net_2021;
	wire new_net_1401;
	wire new_net_1632;
	wire new_net_1254;
	wire new_net_2149;
	wire n_1236_;
	wire new_net_6917;
	wire new_net_8241;
	wire new_net_6845;
	wire new_net_4257;
	wire new_net_10491;
	wire new_net_3587;
	wire new_net_2419;
	wire new_net_3632;
	wire new_net_4329;
	wire new_net_5083;
	wire new_net_6714;
	wire new_net_6797;
	wire new_net_7376;
	wire new_net_7498;
	wire new_net_8707;
	wire new_net_10187;
	wire new_net_6562;
	wire new_net_9521;
	wire new_net_6618;
	wire new_net_10238;
	wire n_1237_;
	wire n_0019_;
	wire n_0229_;
	wire n_0733_;
	wire new_net_3184;
	wire new_net_2026;
	wire new_net_775;
	wire new_net_1220;
	wire n_0840_;
	wire new_net_3428;
	wire new_net_7864;
	wire new_net_9411;
	wire new_net_7862;
	wire new_net_5115;
	wire new_net_8952;
	wire new_net_7368;
	wire new_net_8950;
	wire new_net_10575;
	wire new_net_8484;
	wire new_net_1746;
	wire new_net_3002;
	wire new_net_1893;
	wire new_net_6779;
	wire new_net_8122;
	wire new_net_8142;
	wire new_net_9854;
	wire new_net_8004;
	wire new_net_8539;
	wire new_net_6218;
	wire new_net_8173;
	wire new_net_9668;
	wire new_net_7276;
	wire n_1238_;
	wire new_net_90;
	wire n_0230_;
	wire n_0020_;
	wire n_0734_;
	wire new_net_1369;
	wire new_net_3438;
	wire new_net_2940;
	wire new_net_1402;
	wire new_net_1633;
	wire new_net_9762;
	wire new_net_6206;
	wire new_net_6412;
	wire new_net_8107;
	wire new_net_4599;
	wire new_net_10550;
	wire new_net_5734;
	wire new_net_10159;
	wire new_net_6870;
	wire new_net_2874;
	wire new_net_4128;
	wire new_net_4887;
	wire new_net_5859;
	wire new_net_6137;
	wire new_net_6632;
	wire new_net_6963;
	wire new_net_6288;
	wire new_net_8277;
	wire new_net_8301;
	wire new_net_8871;
	wire new_net_4374;
	wire new_net_7133;
	wire new_net_10062;
	wire new_net_6423;
	wire new_net_7126;
	wire new_net_7096;
	wire new_net_6421;
	wire new_net_4170;
	wire new_net_7779;
	wire new_net_5916;
	wire n_1239_;
	wire n_0021_;
	wire n_0231_;
	wire n_0735_;
	wire new_net_8;
	wire new_net_956;
	wire new_net_1221;
	wire new_net_3888;
	wire new_net_3935;
	wire new_net_4516;
	wire new_net_9364;
	wire new_net_9397;
	wire new_net_10515;
	wire new_net_8236;
	wire new_net_5144;
	wire new_net_7327;
	wire new_net_7697;
	wire new_net_1255;
	wire new_net_1894;
	wire new_net_6106;
	wire new_net_6980;
	wire new_net_7004;
	wire new_net_7123;
	wire new_net_7147;
	wire new_net_9261;
	wire new_net_4071;
	wire new_net_9715;
	wire new_net_6831;
	wire new_net_6180;
	wire new_net_8910;
	wire new_net_5640;
	wire new_net_7915;
	wire n_0736_;
	wire n_0022_;
	wire n_0232_;
	wire n_1240_;
	wire new_net_3588;
	wire new_net_1370;
	wire new_net_1403;
	wire new_net_3633;
	wire new_net_4330;
	wire new_net_6715;
	wire new_net_9269;
	wire new_net_8666;
	wire new_net_9267;
	wire new_net_9794;
	wire new_net_9083;
	wire new_net_9792;
	wire new_net_10072;
	wire new_net_5424;
	wire new_net_7563;
	wire new_net_776;
	wire new_net_3185;
	wire new_net_2420;
	wire new_net_3797;
	wire new_net_4351;
	wire new_net_4757;
	wire new_net_4870;
	wire new_net_5381;
	wire new_net_9076;
	wire new_net_9525;
	wire new_net_9407;
	wire new_net_10005;
	wire new_net_3824;
	wire new_net_7904;
	wire new_net_5267;
	wire new_net_9731;
	wire n_0737_;
	wire n_0023_;
	wire n_0233_;
	wire n_1241_;
	wire new_net_1747;
	wire new_net_3003;
	wire new_net_957;
	wire new_net_6780;
	wire new_net_7099;
	wire new_net_8143;
	wire new_net_4770;
	wire new_net_7290;
	wire new_net_7754;
	wire new_net_10287;
	wire new_net_8766;
	wire new_net_9944;
	wire new_net_10285;
	wire new_net_4541;
	wire new_net_6370;
	wire new_net_8579;
	wire new_net_2941;
	wire new_net_1256;
	wire new_net_91;
	wire new_net_3208;
	wire new_net_1634;
	wire new_net_4473;
	wire new_net_5065;
	wire new_net_5134;
	wire new_net_5295;
	wire new_net_6009;
	wire new_net_10033;
	wire new_net_10031;
	wire new_net_8098;
	wire new_net_8299;
	wire new_net_8931;
	wire new_net_9564;
	wire new_net_9557;
	wire new_net_8929;
	wire new_net_9446;
	wire new_net_7811;
	wire new_net_8463;
	wire new_net_10345;
	wire new_net_9888;
	wire new_net_2959;
	wire n_0738_;
	wire n_0234_;
	wire n_0024_;
	wire n_1242_;
	wire new_net_2074;
	wire new_net_2875;
	wire new_net_1404;
	wire new_net_4888;
	wire new_net_5860;
	wire new_net_6272;
	wire new_net_4957;
	wire new_net_5594;
	wire new_net_4955;
	wire new_net_7082;
	wire new_net_5989;
	wire new_net_777;
	wire new_net_1222;
	wire new_net_3439;
	wire new_net_3889;
	wire new_net_3936;
	wire new_net_4517;
	wire new_net_5103;
	wire new_net_6187;
	wire new_net_6563;
	wire new_net_6587;
	wire new_net_8368;
	wire new_net_9355;
	wire new_net_4502;
	wire new_net_5956;
	wire new_net_7221;
	wire new_net_6727;
	wire new_net_8973;
	wire n_0025_;
	wire n_0235_;
	wire n_1243_;
	wire new_net_1748;
	wire n_0739_;
	wire new_net_1895;
	wire new_net_5029;
	wire new_net_6107;
	wire new_net_6981;
	wire new_net_7005;
	wire new_net_6822;
	wire new_net_7480;
	wire new_net_4234;
	wire new_net_6950;
	wire new_net_9171;
	wire new_net_6497;
	wire new_net_5624;
	wire new_net_2589;
	wire new_net_92;
	wire new_net_2153;
	wire new_net_3589;
	wire new_net_1371;
	wire new_net_2071;
	wire new_net_1635;
	wire new_net_3634;
	wire new_net_4331;
	wire new_net_6716;
	wire new_net_8653;
	wire new_net_9803;
	wire new_net_10133;
	wire new_net_4456;
	wire new_net_5680;
	wire new_net_9505;
	wire new_net_9702;
	wire new_net_6600;
	wire n_0740_;
	wire n_0026_;
	wire n_0236_;
	wire new_net_2960;
	wire n_1244_;
	wire new_net_2645;
	wire new_net_3186;
	wire new_net_3567;
	wire new_net_3798;
	wire new_net_4352;
	wire new_net_7470;
	wire new_net_6690;
	wire new_net_7352;
	wire new_net_4514;
	wire new_net_5100;
	wire new_net_6085;
	wire new_net_4965;
	wire new_net_9091;
	wire new_net_7401;
	wire new_net_5843;
	wire new_net_9248;
	wire new_net_778;
	wire new_net_958;
	wire new_net_1223;
	wire new_net_2148;
	wire new_net_3004;
	wire new_net_2069;
	wire new_net_2421;
	wire new_net_5118;
	wire new_net_6781;
	wire new_net_8144;
	wire new_net_10477;
	wire new_net_8517;
	wire new_net_9135;
	wire new_net_8157;
	wire new_net_9645;
	wire new_net_10639;
	wire new_net_3928;
	wire new_net_8037;
	wire new_net_7253;
	wire new_net_5272;
	wire new_net_1896;
	wire n_0741_;
	wire n_0027_;
	wire n_0237_;
	wire new_net_1257;
	wire n_1245_;
	wire new_net_2942;
	wire new_net_3209;
	wire new_net_3988;
	wire new_net_4474;
	wire new_net_6467;
	wire new_net_8290;
	wire new_net_9548;
	wire new_net_9432;
	wire new_net_7802;
	wire new_net_7978;
	wire new_net_5130;
	wire new_net_93;
	wire new_net_1372;
	wire new_net_1405;
	wire new_net_1636;
	wire new_net_2876;
	wire new_net_5084;
	wire new_net_5861;
	wire new_net_6634;
	wire new_net_6965;
	wire new_net_5296;
	wire new_net_7971;
	wire new_net_5585;
	wire new_net_7442;
	wire new_net_5225;
	wire new_net_6753;
	wire n_0742_;
	wire n_0238_;
	wire n_0028_;
	wire n_1246_;
	wire new_net_3568;
	wire new_net_9;
	wire new_net_3440;
	wire new_net_3890;
	wire new_net_3937;
	wire new_net_4518;
	wire new_net_10600;
	wire new_net_9218;
	wire new_net_10684;
	wire new_net_5947;
	wire new_net_6211;
	wire new_net_8694;
	wire new_net_779;
	wire new_net_959;
	wire new_net_1224;
	wire new_net_1749;
	wire new_net_6108;
	wire new_net_6982;
	wire new_net_7006;
	wire new_net_6159;
	wire new_net_7101;
	wire new_net_7125;
	wire new_net_4895;
	wire new_net_4302;
	wire new_net_6941;
	wire new_net_7522;
	wire new_net_10310;
	wire new_net_5515;
	wire new_net_10308;
	wire n_0743_;
	wire n_0239_;
	wire n_0029_;
	wire new_net_1258;
	wire n_1247_;
	wire new_net_3590;
	wire new_net_2076;
	wire new_net_3635;
	wire new_net_4332;
	wire new_net_4875;
	wire new_net_7032;
	wire new_net_8644;
	wire new_net_9491;
	wire new_net_10054;
	wire new_net_6586;
	wire new_net_10448;
	wire new_net_3792;
	wire new_net_7542;
	wire new_net_3187;
	wire new_net_1406;
	wire new_net_1637;
	wire new_net_2147;
	wire new_net_2961;
	wire new_net_3799;
	wire new_net_4353;
	wire new_net_4872;
	wire new_net_5085;
	wire new_net_8124;
	wire new_net_8792;
	wire new_net_7888;
	wire new_net_10449;
	wire new_net_8252;
	wire new_net_7881;
	wire new_net_8812;
	wire new_net_5829;
	wire new_net_7392;
	wire new_net_10259;
	wire n_1226_;
	wire new_net_8704;
	wire n_0030_;
	wire n_0240_;
	wire n_0744_;
	wire n_1248_;
	wire new_net_2629;
	wire new_net_3005;
	wire new_net_2590;
	wire new_net_6782;
	wire new_net_8145;
	wire new_net_8503;
	wire new_net_10392;
	wire new_net_10390;
	wire new_net_9921;
	wire new_net_6354;
	wire new_net_6242;
	wire new_net_8199;
	wire new_net_10441;
	wire new_net_8197;
	wire new_net_8077;
	wire new_net_2086;
	wire new_net_2422;
	wire new_net_780;
	wire new_net_1750;
	wire new_net_2943;
	wire new_net_2646;
	wire new_net_4130;
	wire new_net_4475;
	wire new_net_5067;
	wire new_net_5136;
	wire new_net_6453;
	wire new_net_6962;
	wire new_net_8276;
	wire new_net_10520;
	wire new_net_8805;
	wire new_net_10329;
	wire new_net_3853;
	wire new_net_4616;
	wire new_net_5742;
	wire new_net_1373;
	wire new_net_2877;
	wire n_0031_;
	wire n_0241_;
	wire n_0745_;
	wire n_1249_;
	wire new_net_94;
	wire new_net_5571;
	wire new_net_5862;
	wire new_net_6635;
	wire new_net_7059;
	wire new_net_9165;
	wire new_net_7150;
	wire new_net_9718;
	wire new_net_2132;
	wire new_net_3569;
	wire new_net_3891;
	wire new_net_3938;
	wire new_net_4519;
	wire new_net_6189;
	wire new_net_6565;
	wire new_net_6589;
	wire new_net_9061;
	wire new_net_9144;
	wire new_net_10675;
	wire new_net_10014;
	wire new_net_7667;
	wire n_0287_;
	wire new_net_7665;
	wire new_net_8834;
	wire new_net_5006;
	wire new_net_960;
	wire new_net_2090;
	wire n_0242_;
	wire n_0032_;
	wire n_0746_;
	wire new_net_1225;
	wire n_1250_;
	wire new_net_6109;
	wire new_net_6150;
	wire new_net_6983;
	wire new_net_4890;
	wire new_net_10255;
	wire new_net_10422;
	wire new_net_6474;
	wire new_net_3999;
	wire new_net_3591;
	wire new_net_781;
	wire new_net_1259;
	wire new_net_1898;
	wire new_net_3636;
	wire new_net_4333;
	wire new_net_6718;
	wire new_net_6801;
	wire new_net_7380;
	wire new_net_7502;
	wire new_net_8630;
	wire new_net_9023;
	wire new_net_9293;
	wire new_net_9021;
	wire new_net_9291;
	wire new_net_5351;
	wire new_net_1374;
	wire new_net_2056;
	wire n_0243_;
	wire n_0033_;
	wire n_0747_;
	wire new_net_1407;
	wire new_net_1638;
	wire new_net_2962;
	wire n_1251_;
	wire new_net_95;
	wire new_net_5820;
	wire new_net_9043;
	wire new_net_6721;
	wire new_net_7383;
	wire new_net_2055;
	wire new_net_3006;
	wire new_net_6783;
	wire new_net_8146;
	wire new_net_9077;
	wire new_net_8494;
	wire new_net_9750;
	wire new_net_9475;
	wire new_net_9858;
	wire new_net_8014;
	wire new_net_7776;
	wire new_net_2647;
	wire new_net_961;
	wire new_net_3441;
	wire n_0748_;
	wire n_0244_;
	wire n_0034_;
	wire new_net_2944;
	wire new_net_2163;
	wire n_1252_;
	wire new_net_1751;
	wire new_net_6622;
	wire new_net_8982;
	wire new_net_10478;
	wire new_net_9772;
	wire new_net_8396;
	wire new_net_8323;
	wire new_net_6098;
	wire new_net_10169;
	wire new_net_8321;
	wire new_net_9180;
	wire new_net_2878;
	wire new_net_782;
	wire new_net_1260;
	wire new_net_1899;
	wire new_net_2423;
	wire new_net_5273;
	wire new_net_5863;
	wire new_net_6636;
	wire new_net_6967;
	wire new_net_8281;
	wire new_net_9110;
	wire new_net_4581;
	wire new_net_9698;
	wire new_net_7050;
	wire new_net_4979;
	wire new_net_6730;
	wire n_0035_;
	wire n_0245_;
	wire n_0749_;
	wire new_net_10;
	wire new_net_1375;
	wire new_net_1408;
	wire new_net_1639;
	wire new_net_3570;
	wire n_1253_;
	wire new_net_96;
	wire new_net_6008;
	wire new_net_7191;
	wire new_net_8224;
	wire new_net_8782;
	wire new_net_6527;
	wire new_net_6110;
	wire new_net_6984;
	wire new_net_7008;
	wire new_net_7103;
	wire new_net_7127;
	wire new_net_7151;
	wire new_net_9167;
	wire new_net_9528;
	wire new_net_9719;
	wire new_net_10118;
	wire new_net_10246;
	wire n_0427_;
	wire new_net_6918;
	wire new_net_6846;
	wire new_net_4258;
	wire new_net_10492;
	wire n_1254_;
	wire new_net_1752;
	wire new_net_3592;
	wire n_0246_;
	wire n_0036_;
	wire n_0750_;
	wire new_net_962;
	wire new_net_1227;
	wire new_net_3637;
	wire new_net_4334;
	wire new_net_8261;
	wire new_net_3189;
	wire new_net_1261;
	wire new_net_2150;
	wire new_net_2963;
	wire new_net_3801;
	wire new_net_4355;
	wire new_net_4874;
	wire new_net_4889;
	wire new_net_5087;
	wire new_net_5104;
	wire new_net_6055;
	wire new_net_10239;
	wire new_net_7865;
	wire new_net_9412;
	wire new_net_9384;
	wire new_net_5116;
	wire new_net_8953;
	wire new_net_7369;
	wire new_net_7626;
	wire new_net_8951;
	wire n_1255_;
	wire new_net_97;
	wire new_net_3007;
	wire n_0247_;
	wire n_0037_;
	wire n_0751_;
	wire new_net_2062;
	wire new_net_6784;
	wire new_net_8126;
	wire new_net_8147;
	wire new_net_8485;
	wire new_net_7713;
	wire new_net_8005;
	wire new_net_8540;
	wire new_net_9669;
	wire new_net_2630;
	wire new_net_2648;
	wire new_net_2945;
	wire new_net_4477;
	wire new_net_5069;
	wire new_net_5131;
	wire new_net_5138;
	wire new_net_5275;
	wire new_net_5299;
	wire new_net_6013;
	wire new_net_6385;
	wire new_net_7277;
	wire new_net_9483;
	wire new_net_10232;
	wire new_net_9763;
	wire new_net_8108;
	wire new_net_4600;
	wire new_net_10551;
	wire new_net_5735;
	wire new_net_6873;
	wire new_net_10160;
	wire n_1256_;
	wire new_net_2637;
	wire n_0038_;
	wire n_0248_;
	wire n_0752_;
	wire new_net_963;
	wire new_net_2879;
	wire new_net_783;
	wire new_net_1900;
	wire new_net_1228;
	wire new_net_6289;
	wire new_net_4375;
	wire new_net_8872;
	wire new_net_6424;
	wire new_net_7097;
	wire new_net_6422;
	wire new_net_9314;
	wire new_net_3571;
	wire new_net_1262;
	wire new_net_1376;
	wire new_net_3442;
	wire new_net_1409;
	wire new_net_1640;
	wire new_net_2424;
	wire new_net_3893;
	wire new_net_3940;
	wire new_net_4521;
	wire new_net_9365;
	wire new_net_4896;
	wire new_net_3774;
	wire new_net_5971;
	wire n_1257_;
	wire n_0753_;
	wire n_0039_;
	wire n_0249_;
	wire new_net_3210;
	wire new_net_5145;
	wire new_net_6111;
	wire new_net_6985;
	wire new_net_7009;
	wire new_net_7104;
	wire new_net_7698;
	wire new_net_6832;
	wire n_0574_;
	wire new_net_6181;
	wire new_net_4845;
	wire new_net_5191;
	wire new_net_8911;
	wire new_net_5700;
	wire new_net_1753;
	wire new_net_2631;
	wire new_net_3593;
	wire new_net_3638;
	wire new_net_4335;
	wire new_net_6720;
	wire new_net_6803;
	wire new_net_7382;
	wire new_net_7504;
	wire new_net_8713;
	wire new_net_9270;
	wire new_net_9268;
	wire new_net_9795;
	wire new_net_9084;
	wire new_net_10073;
	wire new_net_2964;
	wire n_1258_;
	wire new_net_3190;
	wire n_0754_;
	wire n_0250_;
	wire n_0040_;
	wire new_net_784;
	wire new_net_1901;
	wire new_net_3802;
	wire new_net_4356;
	wire new_net_7564;
	wire new_net_4758;
	wire new_net_5382;
	wire new_net_9128;
	wire new_net_9408;
	wire new_net_10006;
	wire new_net_3825;
	wire new_net_8287;
	wire new_net_98;
	wire new_net_2054;
	wire new_net_1377;
	wire new_net_1410;
	wire new_net_1641;
	wire new_net_3008;
	wire new_net_5268;
	wire new_net_5853;
	wire new_net_6785;
	wire new_net_8148;
	wire new_net_9732;
	wire n_0428_;
	wire new_net_3796;
	wire new_net_7992;
	wire new_net_4771;
	wire new_net_8527;
	wire new_net_9425;
	wire new_net_3945;
	wire new_net_7755;
	wire new_net_10288;
	wire new_net_8047;
	wire new_net_9945;
	wire new_net_10286;
	wire new_net_2946;
	wire n_1259_;
	wire n_0041_;
	wire n_0251_;
	wire n_0755_;
	wire new_net_2070;
	wire n_1048_;
	wire new_net_4478;
	wire new_net_4542;
	wire new_net_5070;
	wire new_net_8580;
	wire new_net_10034;
	wire new_net_6202;
	wire new_net_8099;
	wire new_net_8300;
	wire new_net_8932;
	wire new_net_9565;
	wire new_net_9558;
	wire new_net_10146;
	wire new_net_7812;
	wire new_net_8464;
	wire new_net_1754;
	wire new_net_964;
	wire new_net_1229;
	wire new_net_5120;
	wire new_net_5865;
	wire new_net_6638;
	wire new_net_6969;
	wire new_net_8283;
	wire new_net_8307;
	wire new_net_8331;
	wire new_net_9609;
	wire new_net_9889;
	wire new_net_5390;
	wire new_net_5595;
	wire new_net_6273;
	wire new_net_4956;
	wire new_net_7083;
	wire new_net_8394;
	wire new_net_9383;
	wire new_net_5487;
	wire new_net_10211;
	wire new_net_1263;
	wire n_1260_;
	wire n_0042_;
	wire n_0252_;
	wire n_0756_;
	wire new_net_3572;
	wire new_net_11;
	wire new_net_3443;
	wire new_net_785;
	wire new_net_3894;
	wire new_net_9356;
	wire new_net_10610;
	wire new_net_8369;
	wire new_net_6871;
	wire new_net_99;
	wire new_net_1411;
	wire new_net_2151;
	wire new_net_2425;
	wire new_net_6112;
	wire new_net_6986;
	wire new_net_7010;
	wire new_net_7105;
	wire new_net_7129;
	wire new_net_7153;
	wire new_net_8974;
	wire new_net_5030;
	wire new_net_8222;
	wire new_net_6823;
	wire new_net_7481;
	wire new_net_5627;
	wire new_net_7532;
	wire n_0757_;
	wire n_0043_;
	wire n_0253_;
	wire n_1261_;
	wire new_net_2632;
	wire new_net_3594;
	wire new_net_3639;
	wire new_net_4336;
	wire new_net_5121;
	wire new_net_6498;
	wire new_net_8654;
	wire new_net_10134;
	wire new_net_9506;
	wire new_net_9143;
	wire new_net_9703;
	wire new_net_10571;
	wire new_net_1902;
	wire new_net_2965;
	wire new_net_965;
	wire new_net_1230;
	wire new_net_1755;
	wire new_net_2649;
	wire new_net_3191;
	wire new_net_3803;
	wire new_net_4132;
	wire new_net_4357;
	wire new_net_6601;
	wire new_net_7920;
	wire new_net_9119;
	wire new_net_6691;
	wire new_net_7353;
	wire new_net_8259;
	wire new_net_8822;
	wire new_net_786;
	wire new_net_1264;
	wire n_0758_;
	wire n_0254_;
	wire n_0044_;
	wire n_1262_;
	wire new_net_3009;
	wire new_net_1378;
	wire new_net_1642;
	wire new_net_5844;
	wire new_net_7774;
	wire new_net_8714;
	wire new_net_9249;
	wire new_net_10214;
	wire n_0845_;
	wire new_net_8518;
	wire new_net_9136;
	wire new_net_8158;
	wire new_net_9646;
	wire new_net_10640;
	wire new_net_8038;
	wire new_net_1412;
	wire new_net_4479;
	wire new_net_5071;
	wire new_net_5140;
	wire new_net_5277;
	wire new_net_5301;
	wire new_net_6015;
	wire new_net_4414;
	wire new_net_7254;
	wire new_net_7652;
	wire new_net_7916;
	wire new_net_10648;
	wire new_net_8771;
	wire new_net_6468;
	wire new_net_8291;
	wire new_net_5712;
	wire new_net_9549;
	wire new_net_9433;
	wire new_net_7803;
	wire n_0759_;
	wire n_0255_;
	wire n_0045_;
	wire n_1263_;
	wire new_net_5106;
	wire new_net_5866;
	wire new_net_6639;
	wire new_net_6970;
	wire new_net_7979;
	wire new_net_8284;
	wire new_net_9875;
	wire new_net_7972;
	wire new_net_9873;
	wire new_net_8940;
	wire new_net_5297;
	wire new_net_5586;
	wire new_net_9455;
	wire new_net_5976;
	wire new_net_3444;
	wire new_net_1903;
	wire new_net_3573;
	wire new_net_3895;
	wire new_net_3942;
	wire new_net_4523;
	wire new_net_6193;
	wire new_net_6569;
	wire new_net_6593;
	wire new_net_6754;
	wire new_net_10601;
	wire new_net_9219;
	wire new_net_10685;
	wire new_net_9078;
	wire new_net_1643;
	wire new_net_787;
	wire n_0046_;
	wire n_0256_;
	wire n_0760_;
	wire new_net_1265;
	wire n_1264_;
	wire new_net_100;
	wire new_net_3211;
	wire new_net_1379;
	wire new_net_7305;
	wire new_net_7552;
	wire new_net_7983;
	wire new_net_6160;
	wire new_net_4303;
	wire new_net_6979;
	wire new_net_7347;
	wire new_net_6942;
	wire new_net_7523;
	wire new_net_10311;
	wire new_net_2426;
	wire new_net_2633;
	wire new_net_3595;
	wire new_net_3640;
	wire new_net_4337;
	wire new_net_5122;
	wire new_net_5516;
	wire new_net_6722;
	wire new_net_4634;
	wire new_net_6805;
	wire new_net_4876;
	wire new_net_6667;
	wire new_net_10309;
	wire new_net_7033;
	wire new_net_966;
	wire new_net_2083;
	wire new_net_1231;
	wire n_0761_;
	wire n_0047_;
	wire n_0257_;
	wire new_net_2966;
	wire n_1265_;
	wire new_net_1756;
	wire new_net_3192;
	wire new_net_7543;
	wire n_0910_;
	wire new_net_7889;
	wire new_net_7882;
	wire new_net_5247;
	wire new_net_8813;
	wire new_net_3010;
	wire new_net_3212;
	wire new_net_6787;
	wire new_net_8150;
	wire new_net_7393;
	wire new_net_9169;
	wire new_net_9315;
	wire new_net_9573;
	wire new_net_9862;
	wire new_net_3732;
	wire new_net_10393;
	wire new_net_10391;
	wire new_net_9922;
	wire new_net_6355;
	wire new_net_4115;
	wire new_net_6243;
	wire new_net_1380;
	wire new_net_1413;
	wire n_0762_;
	wire n_0258_;
	wire n_0048_;
	wire n_1266_;
	wire new_net_101;
	wire new_net_2650;
	wire new_net_4133;
	wire new_net_4480;
	wire new_net_6454;
	wire new_net_7702;
	wire new_net_10521;
	wire new_net_8806;
	wire new_net_10330;
	wire new_net_4617;
	wire new_net_2880;
	wire new_net_3854;
	wire new_net_5867;
	wire new_net_6113;
	wire new_net_5743;
	wire new_net_6640;
	wire new_net_6971;
	wire new_net_6897;
	wire new_net_8285;
	wire new_net_8309;
	wire new_net_5572;
	wire new_net_12;
	wire new_net_967;
	wire new_net_3445;
	wire new_net_1904;
	wire n_0763_;
	wire n_0259_;
	wire n_0049_;
	wire new_net_1232;
	wire n_1267_;
	wire new_net_1757;
	wire new_net_5217;
	wire new_net_6740;
	wire new_net_10676;
	wire new_net_7668;
	wire new_net_1644;
	wire new_net_788;
	wire new_net_1266;
	wire new_net_6114;
	wire new_net_6988;
	wire new_net_7012;
	wire new_net_7107;
	wire new_net_7131;
	wire new_net_7155;
	wire new_net_8835;
	wire new_net_5007;
	wire new_net_4891;
	wire new_net_10256;
	wire new_net_6928;
	wire new_net_6482;
	wire new_net_10423;
	wire new_net_6475;
	wire new_net_3596;
	wire new_net_1381;
	wire new_net_2072;
	wire new_net_1414;
	wire n_0764_;
	wire n_0260_;
	wire n_0050_;
	wire n_1268_;
	wire new_net_2634;
	wire new_net_3641;
	wire new_net_6653;
	wire new_net_8631;
	wire new_net_9024;
	wire new_net_9294;
	wire new_net_9292;
	wire new_net_5352;
	wire new_net_2139;
	wire new_net_2427;
	wire new_net_2967;
	wire new_net_3193;
	wire new_net_3805;
	wire new_net_4359;
	wire new_net_4892;
	wire new_net_5091;
	wire new_net_8129;
	wire new_net_9065;
	wire new_net_9976;
	wire new_net_10063;
	wire new_net_5864;
	wire new_net_7384;
	wire n_1050_;
	wire new_net_8495;
	wire new_net_9751;
	wire new_net_9476;
	wire new_net_9398;
	wire new_net_10261;
	wire new_net_8015;
	wire new_net_8550;
	wire new_net_8889;
	wire new_net_4398;
	wire new_net_6234;
	wire new_net_3968;
	wire new_net_8069;
	wire new_net_7775;
	wire new_net_8425;
	wire n_1311_;
	wire n_0513_;
	wire n_0807_;
	wire new_net_3423;
	wire n_0303_;
	wire n_1017_;
	wire new_net_3495;
	wire new_net_3128;
	wire new_net_1515;
	wire new_net_3869;
	wire new_net_6623;
	wire new_net_9773;
	wire new_net_8860;
	wire new_net_8324;
	wire new_net_6099;
	wire new_net_10170;
	wire new_net_9181;
	wire new_net_5281;
	wire new_net_9822;
	wire new_net_5274;
	wire new_net_1102;
	wire new_net_2916;
	wire new_net_3541;
	wire new_net_4493;
	wire new_net_5213;
	wire new_net_5315;
	wire new_net_5563;
	wire new_net_6029;
	wire new_net_7540;
	wire new_net_7562;
	wire new_net_7051;
	wire new_net_9699;
	wire new_net_4980;
	wire new_net_6439;
	wire new_net_6731;
	wire n_1312_;
	wire n_0514_;
	wire n_0808_;
	wire new_net_160;
	wire new_net_2164;
	wire n_0304_;
	wire n_1018_;
	wire new_net_1694;
	wire new_net_1922;
	wire new_net_838;
	wire new_net_7192;
	wire new_net_8787;
	wire new_net_9196;
	wire new_net_8785;
	wire new_net_3784;
	wire new_net_2354;
	wire new_net_2552;
	wire new_net_302;
	wire new_net_575;
	wire new_net_1019;
	wire new_net_1284;
	wire new_net_1431;
	wire new_net_1662;
	wire new_net_2739;
	wire new_net_1464;
	wire new_net_10247;
	wire new_net_6919;
	wire new_net_6847;
	wire new_net_8695;
	wire new_net_5651;
	wire new_net_10493;
	wire new_net_7921;
	wire new_net_1516;
	wire n_1313_;
	wire new_net_2833;
	wire new_net_690;
	wire n_0305_;
	wire n_0515_;
	wire n_0809_;
	wire n_1019_;
	wire new_net_2578;
	wire new_net_3730;
	wire new_net_9633;
	wire new_net_5338;
	wire new_net_6571;
	wire new_net_9805;
	wire new_net_6564;
	wire new_net_1775;
	wire new_net_607;
	wire new_net_1103;
	wire new_net_1316;
	wire new_net_2682;
	wire new_net_4810;
	wire new_net_5445;
	wire new_net_5639;
	wire new_net_6042;
	wire new_net_6676;
	wire new_net_7573;
	wire new_net_7866;
	wire new_net_9413;
	wire new_net_8954;
	wire new_net_7370;
	wire new_net_10088;
	wire new_net_8486;
	wire new_net_2980;
	wire new_net_3164;
	wire new_net_3294;
	wire n_1314_;
	wire new_net_119;
	wire new_net_422;
	wire new_net_3403;
	wire n_0516_;
	wire n_0810_;
	wire new_net_161;
	wire new_net_7714;
	wire new_net_2183;
	wire new_net_3806;
	wire new_net_7224;
	wire new_net_8541;
	wire new_net_9670;
	wire new_net_4789;
	wire new_net_4552;
	wire new_net_6386;
	wire new_net_2260;
	wire new_net_2386;
	wire new_net_576;
	wire new_net_1285;
	wire new_net_3496;
	wire new_net_3846;
	wire new_net_4082;
	wire new_net_4395;
	wire new_net_4903;
	wire new_net_4927;
	wire new_net_7278;
	wire new_net_9484;
	wire new_net_9764;
	wire new_net_8109;
	wire new_net_4601;
	wire new_net_10552;
	wire new_net_5736;
	wire new_net_9172;
	wire new_net_10161;
	wire new_net_6874;
	wire new_net_6872;
	wire new_net_2023;
	wire new_net_1517;
	wire n_1315_;
	wire n_0517_;
	wire n_0811_;
	wire new_net_691;
	wire n_1021_;
	wire n_0307_;
	wire new_net_3542;
	wire new_net_2917;
	wire new_net_4376;
	wire new_net_4703;
	wire new_net_6425;
	wire new_net_7128;
	wire new_net_7098;
	wire new_net_4172;
	wire new_net_1776;
	wire new_net_608;
	wire new_net_839;
	wire new_net_1317;
	wire new_net_1923;
	wire new_net_3863;
	wire new_net_4103;
	wire new_net_5236;
	wire new_net_5703;
	wire new_net_5727;
	wire new_net_5918;
	wire new_net_9366;
	wire new_net_7645;
	wire new_net_3775;
	wire new_net_4992;
	wire new_net_9092;
	wire new_net_2787;
	wire n_1316_;
	wire new_net_120;
	wire new_net_423;
	wire n_0518_;
	wire n_0812_;
	wire new_net_162;
	wire n_0308_;
	wire new_net_987;
	wire n_1022_;
	wire new_net_7329;
	wire new_net_7699;
	wire new_net_4073;
	wire new_net_6833;
	wire new_net_7491;
	wire new_net_6182;
	wire new_net_7003;
	wire new_net_8912;
	wire new_net_5701;
	wire new_net_5642;
	wire new_net_2493;
	wire new_net_2541;
	wire new_net_2834;
	wire new_net_2355;
	wire new_net_577;
	wire new_net_1466;
	wire new_net_3731;
	wire new_net_4790;
	wire new_net_6506;
	wire new_net_6530;
	wire new_net_7792;
	wire new_net_9271;
	wire new_net_9796;
	wire new_net_9085;
	wire new_net_5426;
	wire n_1317_;
	wire new_net_1104;
	wire n_0519_;
	wire n_0813_;
	wire n_0309_;
	wire n_1023_;
	wire new_net_4037;
	wire new_net_4759;
	wire new_net_4811;
	wire new_net_5383;
	wire new_net_9129;
	wire new_net_9409;
	wire new_net_10007;
	wire new_net_4835;
	wire new_net_9735;
	wire new_net_5269;
	wire new_net_3121;
	wire new_net_3295;
	wire new_net_2981;
	wire new_net_2087;
	wire new_net_3404;
	wire new_net_840;
	wire new_net_1696;
	wire new_net_1924;
	wire new_net_3307;
	wire new_net_3165;
	wire new_net_6395;
	wire new_net_8528;
	wire new_net_9426;
	wire new_net_7756;
	wire new_net_10289;
	wire new_net_8048;
	wire new_net_9946;
	wire new_net_4543;
	wire new_net_6372;
	wire new_net_8581;
	wire new_net_3497;
	wire new_net_1286;
	wire new_net_2810;
	wire n_1318_;
	wire new_net_121;
	wire new_net_424;
	wire n_0310_;
	wire n_0520_;
	wire n_0814_;
	wire new_net_163;
	wire new_net_10035;
	wire new_net_6203;
	wire new_net_8933;
	wire new_net_9566;
	wire new_net_9559;
	wire new_net_10147;
	wire new_net_7813;
	wire new_net_9963;
	wire new_net_698;
	wire new_net_1467;
	wire new_net_2261;
	wire new_net_1518;
	wire new_net_3543;
	wire new_net_692;
	wire new_net_2387;
	wire new_net_2918;
	wire new_net_4495;
	wire new_net_4670;
	wire new_net_5317;
	wire new_net_5391;
	wire new_net_6276;
	wire new_net_8352;
	wire n_0848_;
	wire new_net_6274;
	wire new_net_4959;
	wire new_net_5596;
	wire new_net_7084;
	wire new_net_8395;
	wire new_net_5488;
	wire new_net_609;
	wire n_1319_;
	wire new_net_1318;
	wire new_net_1777;
	wire n_1025_;
	wire n_0311_;
	wire n_0521_;
	wire n_0815_;
	wire new_net_1105;
	wire new_net_3864;
	wire new_net_6764;
	wire new_net_9357;
	wire new_net_10611;
	wire new_net_4504;
	wire new_net_5958;
	wire new_net_7315;
	wire new_net_2741;
	wire new_net_1697;
	wire new_net_2788;
	wire new_net_988;
	wire new_net_2008;
	wire new_net_2554;
	wire new_net_3818;
	wire new_net_4535;
	wire new_net_6290;
	wire new_net_7708;
	wire new_net_5031;
	wire new_net_8223;
	wire new_net_6824;
	wire new_net_7482;
	wire new_net_6952;
	wire new_net_5628;
	wire new_net_10442;
	wire new_net_6499;
	wire new_net_305;
	wire new_net_1022;
	wire new_net_1665;
	wire new_net_1287;
	wire new_net_2811;
	wire n_1320_;
	wire new_net_122;
	wire new_net_425;
	wire n_1026_;
	wire n_0312_;
	wire new_net_8655;
	wire new_net_10135;
	wire new_net_4458;
	wire new_net_5047;
	wire new_net_8242;
	wire new_net_9507;
	wire new_net_9704;
	wire new_net_10572;
	wire n_1052_;
	wire new_net_1519;
	wire new_net_693;
	wire new_net_1468;
	wire new_net_2356;
	wire new_net_4038;
	wire new_net_4812;
	wire new_net_5641;
	wire new_net_6044;
	wire new_net_6602;
	wire new_net_6678;
	wire new_net_9120;
	wire new_net_6692;
	wire new_net_7354;
	wire new_net_5102;
	wire new_net_6087;
	wire new_net_8260;
	wire new_net_2982;
	wire new_net_3296;
	wire new_net_1925;
	wire new_net_3122;
	wire n_0313_;
	wire n_0523_;
	wire n_1027_;
	wire n_1321_;
	wire new_net_1319;
	wire new_net_1778;
	wire new_net_3870;
	wire new_net_8715;
	wire new_net_9250;
	wire new_net_8519;
	wire new_net_8159;
	wire new_net_9654;
	wire new_net_9647;
	wire new_net_10641;
	wire new_net_8039;
	wire new_net_7257;
	wire new_net_7255;
	wire new_net_3498;
	wire new_net_2131;
	wire new_net_989;
	wire new_net_4084;
	wire new_net_4397;
	wire new_net_4905;
	wire new_net_4929;
	wire new_net_5470;
	wire new_net_5494;
	wire new_net_6233;
	wire new_net_8132;
	wire new_net_6469;
	wire new_net_8772;
	wire new_net_8292;
	wire new_net_5713;
	wire new_net_9550;
	wire new_net_9434;
	wire new_net_7804;
	wire new_net_9876;
	wire n_1028_;
	wire new_net_306;
	wire new_net_1023;
	wire new_net_1666;
	wire n_0314_;
	wire new_net_3544;
	wire n_0524_;
	wire n_0818_;
	wire n_1322_;
	wire new_net_123;
	wire new_net_7973;
	wire new_net_7980;
	wire new_net_9874;
	wire new_net_5298;
	wire new_net_5587;
	wire new_net_7444;
	wire new_net_6413;
	wire new_net_9456;
	wire new_net_2262;
	wire new_net_1106;
	wire new_net_2388;
	wire new_net_3865;
	wire new_net_4105;
	wire new_net_4991;
	wire new_net_5238;
	wire new_net_5705;
	wire new_net_5729;
	wire new_net_5883;
	wire new_net_6755;
	wire new_net_7037;
	wire new_net_9898;
	wire new_net_10602;
	wire new_net_9220;
	wire new_net_10686;
	wire new_net_9079;
	wire new_net_7306;
	wire new_net_2572;
	wire new_net_2742;
	wire new_net_1698;
	wire new_net_1926;
	wire n_0315_;
	wire new_net_842;
	wire new_net_2789;
	wire n_1029_;
	wire n_0525_;
	wire n_0819_;
	wire new_net_6161;
	wire new_net_6943;
	wire new_net_10379;
	wire new_net_7524;
	wire new_net_4017;
	wire new_net_7777;
	wire new_net_10312;
	wire new_net_1435;
	wire new_net_2495;
	wire new_net_2543;
	wire new_net_426;
	wire new_net_990;
	wire new_net_1288;
	wire new_net_2812;
	wire new_net_3733;
	wire new_net_4792;
	wire new_net_5517;
	wire new_net_7034;
	wire new_net_9493;
	wire new_net_5362;
	wire new_net_6588;
	wire new_net_10450;
	wire new_net_7544;
	wire new_net_1469;
	wire n_0316_;
	wire n_1030_;
	wire new_net_1520;
	wire n_1324_;
	wire new_net_124;
	wire new_net_2000;
	wire n_0526_;
	wire n_0820_;
	wire new_net_166;
	wire new_net_9986;
	wire new_net_6073;
	wire new_net_7597;
	wire new_net_7890;
	wire new_net_8254;
	wire new_net_5248;
	wire new_net_7883;
	wire new_net_8814;
	wire new_net_9056;
	wire new_net_6371;
	wire new_net_5831;
	wire new_net_7394;
	wire new_net_3309;
	wire new_net_3123;
	wire new_net_611;
	wire new_net_1107;
	wire new_net_1320;
	wire new_net_2983;
	wire new_net_3167;
	wire new_net_3297;
	wire new_net_3406;
	wire new_net_2357;
	wire new_net_8505;
	wire new_net_10394;
	wire new_net_9923;
	wire new_net_3315;
	wire new_net_2007;
	wire new_net_1699;
	wire new_net_1927;
	wire new_net_3499;
	wire n_0317_;
	wire n_0527_;
	wire n_0821_;
	wire n_1031_;
	wire new_net_2128;
	wire n_1325_;
	wire new_net_6455;
	wire new_net_7703;
	wire new_net_8079;
	wire new_net_10522;
	wire new_net_6964;
	wire new_net_8278;
	wire new_net_8807;
	wire new_net_10331;
	wire new_net_5746;
	wire new_net_8334;
	wire new_net_5744;
	wire new_net_1436;
	wire new_net_1667;
	wire new_net_2920;
	wire new_net_307;
	wire new_net_427;
	wire new_net_580;
	wire new_net_991;
	wire new_net_1024;
	wire new_net_1289;
	wire new_net_3545;
	wire new_net_6898;
	wire new_net_5573;
	wire new_net_8216;
	wire new_net_5467;
	wire new_net_7061;
	wire new_net_9447;
	wire new_net_6741;
	wire new_net_7152;
	wire new_net_9720;
	wire new_net_167;
	wire new_net_695;
	wire n_1032_;
	wire new_net_1470;
	wire n_0528_;
	wire n_0822_;
	wire n_0318_;
	wire new_net_1521;
	wire n_1326_;
	wire new_net_125;
	wire new_net_8350;
	wire new_net_10240;
	wire new_net_9385;
	wire new_net_10677;
	wire new_net_6341;
	wire new_net_7669;
	wire n_0294_;
	wire new_net_2790;
	wire new_net_2263;
	wire new_net_2743;
	wire new_net_2556;
	wire new_net_2082;
	wire new_net_612;
	wire new_net_843;
	wire new_net_2389;
	wire new_net_1321;
	wire new_net_1780;
	wire new_net_3619;
	wire new_net_6152;
	wire new_net_4657;
	wire new_net_10424;
	wire new_net_1858;
	wire new_net_6483;
	wire new_net_6476;
	wire new_net_4001;
	wire new_net_5132;
	wire n_1033_;
	wire new_net_1928;
	wire n_0529_;
	wire n_0823_;
	wire n_0319_;
	wire new_net_2133;
	wire new_net_2813;
	wire n_1327_;
	wire new_net_2004;
	wire new_net_3734;
	wire new_net_8632;
	wire new_net_9295;
	wire new_net_5353;
	wire new_net_10358;
	wire new_net_308;
	wire new_net_428;
	wire new_net_581;
	wire new_net_1025;
	wire new_net_1668;
	wire new_net_1975;
	wire new_net_4040;
	wire new_net_4775;
	wire new_net_4814;
	wire new_net_5643;
	wire new_net_9977;
	wire new_net_10064;
	wire new_net_6723;
	wire new_net_7385;
	wire n_1328_;
	wire new_net_126;
	wire new_net_3407;
	wire n_0530_;
	wire n_0824_;
	wire new_net_168;
	wire new_net_1108;
	wire new_net_3310;
	wire new_net_1471;
	wire new_net_3124;
	wire n_0775_;
	wire new_net_8496;
	wire new_net_9477;
	wire new_net_9399;
	wire new_net_8018;
	wire new_net_10262;
	wire new_net_8551;
	wire new_net_6235;
	wire new_net_1322;
	wire new_net_1781;
	wire new_net_2358;
	wire new_net_1700;
	wire new_net_3500;
	wire new_net_613;
	wire new_net_844;
	wire new_net_4086;
	wire new_net_4399;
	wire new_net_4907;
	wire new_net_8070;
	wire new_net_8984;
	wire new_net_10122;
	wire new_net_6624;
	wire new_net_9774;
	wire new_net_8325;
	wire new_net_9825;
	wire new_net_10171;
	wire new_net_9182;
	wire n_1329_;
	wire n_0531_;
	wire n_0825_;
	wire new_net_992;
	wire new_net_2167;
	wire new_net_1437;
	wire new_net_2921;
	wire n_1035_;
	wire n_0321_;
	wire new_net_1290;
	wire new_net_5282;
	wire new_net_5564;
	wire new_net_8130;
	wire new_net_9760;
	wire new_net_9700;
	wire new_net_1731;
	wire new_net_7052;
	wire new_net_6300;
	wire new_net_4981;
	wire new_net_6851;
	wire new_net_6732;
	wire new_net_1669;
	wire new_net_309;
	wire new_net_429;
	wire new_net_696;
	wire new_net_1522;
	wire new_net_3867;
	wire new_net_4993;
	wire new_net_5216;
	wire new_net_5240;
	wire new_net_5562;
	wire new_net_6010;
	wire new_net_9199;
	wire new_net_9197;
	wire new_net_6788;
	wire new_net_8786;
	wire new_net_6414;
	wire new_net_6786;
	wire new_net_3785;
	wire n_1330_;
	wire new_net_127;
	wire new_net_169;
	wire new_net_1109;
	wire new_net_2744;
	wire n_0532_;
	wire n_0826_;
	wire n_1036_;
	wire n_0441_;
	wire new_net_1472;
	wire new_net_9999;
	wire new_net_10248;
	wire new_net_7993;
	wire new_net_6920;
	wire new_net_6848;
	wire new_net_7013;
	wire new_net_4260;
	wire new_net_4596;
	wire new_net_2814;
	wire new_net_1323;
	wire new_net_2390;
	wire new_net_614;
	wire new_net_1701;
	wire new_net_1929;
	wire new_net_2497;
	wire new_net_2264;
	wire new_net_2545;
	wire new_net_4794;
	wire new_net_5652;
	wire new_net_7922;
	wire new_net_10494;
	wire new_net_9634;
	wire new_net_6572;
	wire new_net_9806;
	wire new_net_1291;
	wire n_1331_;
	wire new_net_2835;
	wire new_net_993;
	wire n_1037_;
	wire new_net_1026;
	wire new_net_1438;
	wire n_0827_;
	wire n_0533_;
	wire new_net_582;
	wire new_net_7867;
	wire new_net_9414;
	wire new_net_10233;
	wire new_net_7371;
	wire new_net_1523;
	wire new_net_2985;
	wire new_net_3169;
	wire new_net_3299;
	wire new_net_3408;
	wire new_net_3311;
	wire new_net_310;
	wire new_net_430;
	wire new_net_697;
	wire new_net_3125;
	wire new_net_8487;
	wire new_net_7715;
	wire new_net_4094;
	wire new_net_7225;
	wire new_net_8542;
	wire new_net_9671;
	wire new_net_4669;
	wire new_net_8057;
	wire new_net_845;
	wire n_1332_;
	wire new_net_128;
	wire new_net_1782;
	wire n_0534_;
	wire n_0828_;
	wire n_0324_;
	wire n_1038_;
	wire new_net_1110;
	wire new_net_3501;
	wire new_net_7279;
	wire new_net_9485;
	wire new_net_8112;
	wire new_net_9765;
	wire new_net_8110;
	wire new_net_3172;
	wire new_net_4602;
	wire new_net_5737;
	wire new_net_9173;
	wire new_net_6875;
	wire new_net_10162;
	wire new_net_3547;
	wire new_net_2359;
	wire new_net_3425;
	wire new_net_2922;
	wire new_net_1930;
	wire new_net_4499;
	wire new_net_5321;
	wire new_net_6213;
	wire new_net_7567;
	wire new_net_7696;
	wire new_net_7038;
	wire new_net_6291;
	wire new_net_5606;
	wire new_net_4377;
	wire new_net_6426;
	wire new_net_1292;
	wire n_1333_;
	wire n_0535_;
	wire n_0829_;
	wire n_0325_;
	wire n_1039_;
	wire new_net_1027;
	wire new_net_1670;
	wire new_net_583;
	wire new_net_3868;
	wire new_net_9367;
	wire new_net_4898;
	wire new_net_8849;
	wire new_net_7646;
	wire new_net_9166;
	wire new_net_9093;
	wire new_net_2792;
	wire new_net_2558;
	wire new_net_431;
	wire new_net_1473;
	wire new_net_2745;
	wire new_net_3822;
	wire new_net_4931;
	wire new_net_6294;
	wire new_net_7712;
	wire new_net_5147;
	wire new_net_7330;
	wire new_net_7700;
	wire new_net_6834;
	wire new_net_9137;
	wire n_0581_;
	wire new_net_10015;
	wire new_net_4847;
	wire new_net_8913;
	wire new_net_1702;
	wire new_net_615;
	wire new_net_846;
	wire new_net_2815;
	wire n_1334_;
	wire new_net_129;
	wire new_net_1324;
	wire new_net_1783;
	wire new_net_171;
	wire n_0326_;
	wire new_net_5536;
	wire new_net_9272;
	wire new_net_8898;
	wire new_net_2053;
	wire new_net_9797;
	wire new_net_8263;
	wire new_net_2265;
	wire new_net_2391;
	wire new_net_994;
	wire new_net_1439;
	wire new_net_1931;
	wire new_net_4042;
	wire new_net_4776;
	wire new_net_4816;
	wire new_net_5645;
	wire new_net_5427;
	wire new_net_6043;
	wire new_net_5384;
	wire new_net_9410;
	wire new_net_10008;
	wire new_net_6707;
	wire new_net_3827;
	wire new_net_3126;
	wire new_net_2576;
	wire new_net_1293;
	wire new_net_1524;
	wire new_net_2986;
	wire new_net_3170;
	wire new_net_3300;
	wire n_1335_;
	wire new_net_3409;
	wire n_0537_;
	wire new_net_5270;
	wire new_net_9734;
	wire new_net_5855;
	wire new_net_8529;
	wire new_net_9427;
	wire new_net_3947;
	wire new_net_7757;
	wire new_net_8983;
	wire new_net_10290;
	wire n_1062_;
	wire new_net_8049;
	wire new_net_9947;
	wire new_net_2585;
	wire new_net_3502;
	wire new_net_2836;
	wire new_net_3430;
	wire new_net_432;
	wire new_net_1111;
	wire new_net_1474;
	wire n_1055_;
	wire new_net_3738;
	wire new_net_4088;
	wire new_net_4544;
	wire new_net_6373;
	wire new_net_8582;
	wire new_net_10036;
	wire new_net_4588;
	wire new_net_2280;
	wire new_net_8302;
	wire new_net_8934;
	wire new_net_9567;
	wire new_net_9560;
	wire new_net_10148;
	wire new_net_2923;
	wire new_net_1703;
	wire new_net_616;
	wire new_net_2130;
	wire new_net_3548;
	wire n_1336_;
	wire new_net_130;
	wire new_net_1325;
	wire new_net_1784;
	wire n_0538_;
	wire new_net_1352;
	wire new_net_7814;
	wire new_net_9611;
	wire new_net_9891;
	wire new_net_6277;
	wire new_net_5392;
	wire new_net_4960;
	wire new_net_5597;
	wire new_net_6275;
	wire new_net_7454;
	wire new_net_8563;
	wire new_net_5491;
	wire new_net_10563;
	wire new_net_7085;
	wire new_net_3517;
	wire new_net_5489;
	wire new_net_1440;
	wire new_net_1932;
	wire new_net_2360;
	wire new_net_584;
	wire new_net_995;
	wire new_net_4108;
	wire new_net_4995;
	wire new_net_5218;
	wire new_net_5242;
	wire new_net_5685;
	wire new_net_5992;
	wire new_net_1384;
	wire new_net_7555;
	wire new_net_6765;
	wire new_net_9358;
	wire new_net_10612;
	wire new_net_440;
	wire n_0916_;
	wire new_net_3426;
	wire new_net_312;
	wire new_net_2746;
	wire new_net_2793;
	wire new_net_1525;
	wire n_1337_;
	wire n_0539_;
	wire n_0833_;
	wire new_net_699;
	wire n_0329_;
	wire new_net_5133;
	wire new_net_7316;
	wire new_net_3643;
	wire new_net_6825;
	wire new_net_7483;
	wire new_net_9532;
	wire new_net_6953;
	wire new_net_5629;
	wire new_net_2547;
	wire new_net_2816;
	wire new_net_847;
	wire new_net_1112;
	wire new_net_2499;
	wire new_net_3312;
	wire new_net_6500;
	wire new_net_6512;
	wire new_net_6536;
	wire new_net_6560;
	wire new_net_10443;
	wire new_net_2032;
	wire new_net_3261;
	wire new_net_8656;
	wire new_net_10136;
	wire new_net_9508;
	wire new_net_9145;
	wire new_net_9705;
	wire new_net_10573;
	wire n_1044_;
	wire new_net_1704;
	wire n_1338_;
	wire new_net_131;
	wire new_net_173;
	wire n_0540_;
	wire n_0834_;
	wire n_0330_;
	wire new_net_4043;
	wire new_net_4817;
	wire new_net_6603;
	wire new_net_9121;
	wire new_net_8865;
	wire new_net_6693;
	wire new_net_7355;
	wire new_net_4726;
	wire new_net_1672;
	wire new_net_3127;
	wire new_net_2266;
	wire new_net_2987;
	wire new_net_3171;
	wire new_net_3301;
	wire new_net_3410;
	wire new_net_585;
	wire new_net_1294;
	wire new_net_1441;
	wire new_net_7404;
	wire new_net_8718;
	wire new_net_8716;
	wire new_net_9251;
	wire new_net_3871;
	wire new_net_10404;
	wire new_net_8520;
	wire new_net_8160;
	wire new_net_9655;
	wire n_0582_;
	wire new_net_4322;
	wire new_net_9648;
	wire n_1045_;
	wire new_net_1475;
	wire new_net_3503;
	wire n_0331_;
	wire n_1339_;
	wire new_net_433;
	wire new_net_2837;
	wire new_net_700;
	wire n_0541_;
	wire n_0835_;
	wire new_net_3711;
	wire new_net_6254;
	wire new_net_4416;
	wire new_net_7256;
	wire new_net_7918;
	wire new_net_8836;
	wire new_net_10650;
	wire new_net_4932;
	wire new_net_8773;
	wire new_net_8293;
	wire new_net_4982;
	wire new_net_6852;
	wire new_net_9435;
	wire new_net_2924;
	wire new_net_3549;
	wire new_net_1785;
	wire new_net_617;
	wire new_net_1982;
	wire new_net_1113;
	wire new_net_1326;
	wire new_net_4501;
	wire new_net_4674;
	wire new_net_4778;
	wire new_net_9877;
	wire new_net_7981;
	wire new_net_5588;
	wire new_net_996;
	wire new_net_0;
	wire n_1340_;
	wire new_net_132;
	wire new_net_2005;
	wire n_1046_;
	wire n_0332_;
	wire n_0713_;
	wire n_0542_;
	wire n_0836_;
	wire new_net_5978;
	wire new_net_6756;
	wire new_net_10603;
	wire new_net_2740;
	wire new_net_9899;
	wire new_net_2738;
	wire new_net_9221;
	wire new_net_10687;
	wire n_1063_;
	wire new_net_2560;
	wire new_net_1673;
	wire new_net_2747;
	wire new_net_2794;
	wire new_net_1526;
	wire new_net_313;
	wire new_net_1295;
	wire new_net_1442;
	wire new_net_2361;
	wire new_net_3427;
	wire n_1056_;
	wire new_net_7307;
	wire new_net_7554;
	wire new_net_6162;
	wire new_net_6944;
	wire new_net_7525;
	wire new_net_1476;
	wire n_0333_;
	wire new_net_2817;
	wire n_1341_;
	wire new_net_434;
	wire n_1047_;
	wire n_0543_;
	wire n_0837_;
	wire new_net_701;
	wire new_net_6513;
	wire new_net_10313;
	wire new_net_5518;
	wire new_net_6669;
	wire new_net_7035;
	wire new_net_8861;
	wire n_0297_;
	wire new_net_1705;
	wire new_net_1786;
	wire new_net_1327;
	wire new_net_618;
	wire new_net_4044;
	wire new_net_4818;
	wire new_net_5363;
	wire new_net_5647;
	wire new_net_6050;
	wire new_net_6684;
	wire new_net_4742;
	wire new_net_9987;
	wire new_net_9624;
	wire new_net_7598;
	wire new_net_3062;
	wire new_net_5330;
	wire new_net_7891;
	wire new_net_8255;
	wire new_net_5249;
	wire new_net_1934;
	wire n_0838_;
	wire new_net_133;
	wire n_0544_;
	wire new_net_997;
	wire new_net_3313;
	wire new_net_586;
	wire n_1342_;
	wire n_0334_;
	wire new_net_1030;
	wire new_net_7395;
	wire new_net_8506;
	wire new_net_10395;
	wire new_net_9924;
	wire new_net_3504;
	wire new_net_2393;
	wire new_net_2267;
	wire new_net_314;
	wire new_net_1527;
	wire new_net_4117;
	wire new_net_4403;
	wire new_net_4676;
	wire new_net_4911;
	wire new_net_5452;
	wire new_net_6183;
	wire new_net_7056;
	wire new_net_7906;
	wire new_net_8080;
	wire new_net_7704;
	wire n_0158_;
	wire new_net_10523;
	wire new_net_8279;
	wire new_net_2175;
	wire new_net_10332;
	wire new_net_1114;
	wire new_net_2009;
	wire n_0335_;
	wire new_net_849;
	wire new_net_3550;
	wire n_0545_;
	wire n_0839_;
	wire n_1049_;
	wire n_1343_;
	wire new_net_3856;
	wire new_net_5745;
	wire new_net_6899;
	wire new_net_5574;
	wire new_net_5468;
	wire new_net_7062;
	wire new_net_10086;
	wire new_net_1706;
	wire new_net_619;
	wire new_net_1328;
	wire new_net_4110;
	wire new_net_4997;
	wire new_net_2367;
	wire new_net_5220;
	wire new_net_5244;
	wire new_net_5687;
	wire new_net_5711;
	wire new_net_5219;
	wire new_net_6742;
	wire new_net_9721;
	wire new_net_8056;
	wire new_net_8351;
	wire new_net_10241;
	wire new_net_9386;
	wire new_net_10678;
	wire new_net_2786;
	wire new_net_7670;
	wire new_net_8955;
	wire n_1344_;
	wire new_net_134;
	wire new_net_176;
	wire new_net_998;
	wire new_net_1031;
	wire new_net_1443;
	wire new_net_1674;
	wire new_net_2748;
	wire new_net_587;
	wire n_0336_;
	wire new_net_5011;
	wire new_net_7545;
	wire new_net_7628;
	wire new_net_10103;
	wire new_net_3574;
	wire new_net_10427;
	wire new_net_6930;
	wire new_net_6484;
	wire new_net_10425;
	wire new_net_2362;
	wire new_net_2501;
	wire new_net_2549;
	wire new_net_315;
	wire new_net_435;
	wire new_net_702;
	wire new_net_1477;
	wire new_net_1528;
	wire new_net_2818;
	wire new_net_6477;
	wire new_net_6655;
	wire new_net_7565;
	wire new_net_5560;
	wire new_net_9809;
	wire new_net_9296;
	wire n_1345_;
	wire new_net_1787;
	wire n_0547_;
	wire n_0841_;
	wire new_net_1115;
	wire new_net_2570;
	wire new_net_1;
	wire n_0337_;
	wire new_net_850;
	wire n_1051_;
	wire n_0714_;
	wire new_net_10359;
	wire new_net_9978;
	wire new_net_6677;
	wire new_net_1958;
	wire new_net_1985;
	wire new_net_3412;
	wire new_net_1981;
	wire new_net_3303;
	wire new_net_3314;
	wire new_net_2925;
	wire new_net_3129;
	wire n_1064_;
	wire new_net_1935;
	wire new_net_2989;
	wire new_net_9235;
	wire n_1057_;
	wire new_net_8497;
	wire new_net_8019;
	wire new_net_10263;
	wire new_net_7856;
	wire new_net_8017;
	wire new_net_7235;
	wire new_net_8552;
	wire new_net_8891;
	wire n_1346_;
	wire new_net_135;
	wire n_0548_;
	wire n_0842_;
	wire new_net_177;
	wire new_net_999;
	wire new_net_1444;
	wire new_net_1675;
	wire new_net_588;
	wire new_net_3505;
	wire new_net_3970;
	wire new_net_4393;
	wire new_net_3132;
	wire new_net_7778;
	wire new_net_8071;
	wire new_net_8353;
	wire new_net_8465;
	wire new_net_8987;
	wire new_net_1708;
	wire new_net_3130;
	wire new_net_8985;
	wire new_net_10123;
	wire new_net_9775;
	wire new_net_1529;
	wire new_net_2394;
	wire new_net_2268;
	wire new_net_316;
	wire new_net_436;
	wire new_net_703;
	wire new_net_1478;
	wire new_net_4503;
	wire new_net_4780;
	wire new_net_5325;
	wire new_net_6885;
	wire new_net_9183;
	wire new_net_9826;
	wire new_net_10172;
	wire new_net_9824;
	wire new_net_1385;
	wire new_net_8131;
	wire new_net_5276;
	wire new_net_2392;
	wire new_net_5565;
	wire new_net_5459;
	wire new_net_7053;
	wire new_net_8370;
	wire new_net_6301;
	wire n_0918_;
	wire new_net_1860;
	wire n_0003_;
	wire n_1347_;
	wire new_net_1788;
	wire new_net_1329;
	wire new_net_1707;
	wire n_0339_;
	wire new_net_620;
	wire n_0549_;
	wire n_0843_;
	wire n_1053_;
	wire new_net_6733;
	wire new_net_9086;
	wire new_net_9328;
	wire new_net_9200;
	wire new_net_6011;
	wire new_net_2984;
	wire new_net_2039;
	wire new_net_9198;
	wire new_net_2006;
	wire new_net_3429;
	wire new_net_2562;
	wire new_net_2078;
	wire new_net_1936;
	wire new_net_1032;
	wire new_net_2796;
	wire new_net_2749;
	wire new_net_3739;
	wire new_net_3826;
	wire n_1302_;
	wire new_net_4262;
	wire new_net_6921;
	wire new_net_791;
	wire new_net_8450;
	wire new_net_6849;
	wire new_net_9845;
	wire n_0004_;
	wire new_net_2819;
	wire n_1348_;
	wire new_net_136;
	wire new_net_178;
	wire n_1054_;
	wire new_net_2025;
	wire n_0550_;
	wire n_0844_;
	wire n_0340_;
	wire new_net_10497;
	wire new_net_5653;
	wire new_net_10495;
	wire new_net_7923;
	wire new_net_9635;
	wire new_net_154;
	wire new_net_8676;
	wire new_net_5681;
	wire new_net_6573;
	wire new_net_9807;
	wire new_net_2038;
	wire new_net_2363;
	wire new_net_437;
	wire new_net_704;
	wire new_net_1116;
	wire new_net_4046;
	wire new_net_4796;
	wire new_net_4820;
	wire new_net_5649;
	wire new_net_6052;
	wire new_net_6566;
	wire new_net_2684;
	wire new_net_3433;
	wire new_net_7575;
	wire new_net_10479;
	wire new_net_9415;
	wire new_net_3348;
	wire n_0341_;
	wire new_net_621;
	wire n_0005_;
	wire new_net_2990;
	wire new_net_3174;
	wire new_net_3304;
	wire n_1349_;
	wire new_net_1330;
	wire new_net_1789;
	wire new_net_3413;
	wire new_net_8488;
	wire new_net_7718;
	wire new_net_7716;
	wire new_net_3808;
	wire new_net_8543;
	wire new_net_6222;
	wire new_net_1445;
	wire new_net_1676;
	wire new_net_3506;
	wire new_net_589;
	wire new_net_1000;
	wire new_net_1033;
	wire new_net_1298;
	wire new_net_4405;
	wire new_net_4913;
	wire new_net_4934;
	wire new_net_9672;
	wire new_net_4791;
	wire new_net_4554;
	wire new_net_7280;
	wire new_net_9766;
	wire new_net_8113;
	wire new_net_8111;
	wire new_net_3173;
	wire new_net_1005;
	wire new_net_4603;
	wire n_0342_;
	wire new_net_2574;
	wire n_0006_;
	wire new_net_1530;
	wire n_1350_;
	wire new_net_137;
	wire new_net_2010;
	wire n_0552_;
	wire n_0846_;
	wire new_net_179;
	wire new_net_6876;
	wire new_net_9174;
	wire new_net_10163;
	wire n_0445_;
	wire new_net_5778;
	wire new_net_7039;
	wire new_net_6292;
	wire new_net_4707;
	wire new_net_4378;
	wire new_net_2269;
	wire new_net_1117;
	wire new_net_2395;
	wire new_net_2568;
	wire new_net_438;
	wire new_net_705;
	wire new_net_852;
	wire new_net_4112;
	wire new_net_4179;
	wire new_net_5222;
	wire new_net_7130;
	wire new_net_915;
	wire new_net_4347;
	wire new_net_5920;
	wire new_net_9368;
	wire new_net_7647;
	wire new_net_1937;
	wire n_0343_;
	wire new_net_2797;
	wire n_0007_;
	wire n_1351_;
	wire new_net_2014;
	wire new_net_1790;
	wire new_net_2750;
	wire n_0553_;
	wire n_0847_;
	wire new_net_4994;
	wire new_net_9094;
	wire new_net_7331;
	wire new_net_4075;
	wire new_net_6835;
	wire new_net_7493;
	wire new_net_10016;
	wire n_0306_;
	wire new_net_2503;
	wire new_net_2820;
	wire new_net_2838;
	wire new_net_1677;
	wire new_net_2;
	wire new_net_590;
	wire n_0299_;
	wire new_net_1001;
	wire new_net_1299;
	wire new_net_1446;
	wire new_net_8914;
	wire new_net_5644;
	wire new_net_9273;
	wire n_0919_;
	wire new_net_5331;
	wire new_net_9798;
	wire new_net_1480;
	wire n_0344_;
	wire n_0008_;
	wire new_net_1531;
	wire n_1352_;
	wire new_net_138;
	wire new_net_180;
	wire n_1058_;
	wire new_net_318;
	wire n_0554_;
	wire new_net_10583;
	wire new_net_5428;
	wire new_net_8226;
	wire new_net_7566;
	wire new_net_5385;
	wire new_net_10009;
	wire new_net_1709;
	wire new_net_3131;
	wire new_net_3553;
	wire new_net_853;
	wire new_net_3316;
	wire new_net_2991;
	wire new_net_3305;
	wire new_net_2364;
	wire new_net_3175;
	wire new_net_2186;
	wire new_net_7534;
	wire new_net_9457;
	wire new_net_9737;
	wire new_net_4773;
	wire new_net_8530;
	wire new_net_3666;
	wire new_net_3948;
	wire new_net_7758;
	wire new_net_9080;
	wire new_net_10291;
	wire new_net_9948;
	wire new_net_4545;
	wire new_net_6374;
	wire new_net_8583;
	wire new_net_9752;
	wire new_net_10037;
	wire new_net_8303;
	wire new_net_8935;
	wire new_net_9568;
	wire new_net_9561;
	wire new_net_10149;
	wire new_net_7817;
	wire new_net_8554;
	wire new_net_7815;
	wire new_net_8466;
	wire new_net_9965;
	wire n_0093_;
	wire n_0597_;
	wire n_1101_;
	wire new_net_3359;
	wire new_net_3383;
	wire new_net_1134;
	wire new_net_1167;
	wire new_net_4418;
	wire new_net_8163;
	wire new_net_8187;
	wire new_net_9892;
	wire new_net_6278;
	wire new_net_4961;
	wire new_net_5598;
	wire new_net_9733;
	wire new_net_5492;
	wire new_net_7086;
	wire new_net_4131;
	wire new_net_10451;
	wire new_net_336;
	wire new_net_456;
	wire new_net_1051;
	wire new_net_2651;
	wire new_net_1807;
	wire new_net_4635;
	wire new_net_4704;
	wire new_net_5154;
	wire new_net_5279;
	wire new_net_6766;
	wire new_net_9359;
	wire new_net_10613;
	wire new_net_8371;
	wire new_net_5960;
	wire new_net_8815;
	wire n_1102_;
	wire n_0094_;
	wire n_0598_;
	wire new_net_673;
	wire new_net_1547;
	wire new_net_5758;
	wire new_net_5035;
	wire new_net_5782;
	wire new_net_7067;
	wire new_net_7233;
	wire new_net_7317;
	wire new_net_5033;
	wire new_net_8788;
	wire new_net_6826;
	wire new_net_4238;
	wire new_net_9533;
	wire new_net_6954;
	wire new_net_5630;
	wire new_net_10444;
	wire new_net_38;
	wire new_net_722;
	wire new_net_2717;
	wire new_net_3079;
	wire new_net_2459;
	wire new_net_2228;
	wire new_net_2763;
	wire new_net_2291;
	wire new_net_2564;
	wire new_net_3753;
	wire new_net_6501;
	wire new_net_9509;
	wire new_net_9146;
	wire new_net_9706;
	wire new_net_10574;
	wire n_0095_;
	wire n_1103_;
	wire n_0599_;
	wire new_net_1168;
	wire new_net_3274;
	wire new_net_3098;
	wire new_net_1996;
	wire new_net_1135;
	wire new_net_5926;
	wire new_net_6604;
	wire new_net_6694;
	wire new_net_7356;
	wire new_net_7349;
	wire new_net_8719;
	wire new_net_337;
	wire new_net_457;
	wire new_net_1052;
	wire new_net_1955;
	wire new_net_4060;
	wire new_net_5175;
	wire new_net_6066;
	wire new_net_6700;
	wire new_net_7398;
	wire new_net_7405;
	wire new_net_9252;
	wire new_net_3872;
	wire new_net_10405;
	wire new_net_8521;
	wire new_net_8161;
	wire new_net_9656;
	wire new_net_9890;
	wire new_net_8397;
	wire new_net_9649;
	wire new_net_8041;
	wire new_net_7259;
	wire new_net_3712;
	wire new_net_6255;
	wire n_0096_;
	wire n_1104_;
	wire n_0600_;
	wire new_net_2028;
	wire new_net_2900;
	wire new_net_674;
	wire new_net_1548;
	wire new_net_3776;
	wire new_net_4254;
	wire new_net_4417;
	wire new_net_8837;
	wire new_net_4933;
	wire new_net_8774;
	wire new_net_8294;
	wire new_net_4983;
	wire new_net_6853;
	wire new_net_9436;
	wire new_net_39;
	wire new_net_3360;
	wire new_net_2121;
	wire new_net_3384;
	wire new_net_2323;
	wire new_net_4419;
	wire new_net_8164;
	wire new_net_4785;
	wire new_net_6909;
	wire new_net_7982;
	wire new_net_9878;
	wire new_net_5300;
	wire new_net_5589;
	wire new_net_7446;
	wire new_net_9026;
	wire new_net_5979;
	wire n_0097_;
	wire n_0601_;
	wire n_1105_;
	wire new_net_4636;
	wire new_net_4681;
	wire new_net_4705;
	wire new_net_5155;
	wire new_net_5280;
	wire new_net_6757;
	wire new_net_8043;
	wire new_net_10649;
	wire new_net_10604;
	wire new_net_9222;
	wire new_net_10018;
	wire new_net_10688;
	wire new_net_458;
	wire new_net_1956;
	wire new_net_3140;
	wire new_net_5759;
	wire new_net_5783;
	wire new_net_7068;
	wire new_net_7234;
	wire new_net_7258;
	wire new_net_7308;
	wire new_net_8504;
	wire new_net_9400;
	wire new_net_5682;
	wire new_net_6945;
	wire new_net_8262;
	wire new_net_7526;
	wire new_net_10314;
	wire n_0098_;
	wire n_0602_;
	wire n_1106_;
	wire new_net_2718;
	wire new_net_3080;
	wire new_net_2764;
	wire new_net_675;
	wire new_net_3754;
	wire new_net_4015;
	wire new_net_5339;
	wire new_net_5519;
	wire new_net_7036;
	wire new_net_9495;
	wire new_net_9586;
	wire new_net_40;
	wire new_net_1136;
	wire new_net_1169;
	wire new_net_2229;
	wire new_net_2460;
	wire new_net_3099;
	wire new_net_3551;
	wire new_net_2292;
	wire new_net_5798;
	wire new_net_5927;
	wire new_net_6590;
	wire new_net_9988;
	wire new_net_9625;
	wire new_net_6075;
	wire new_net_7599;
	wire new_net_7892;
	wire new_net_7885;
	wire new_net_9058;
	wire new_net_1809;
	wire n_1107_;
	wire n_0099_;
	wire n_0603_;
	wire new_net_338;
	wire new_net_1053;
	wire new_net_3518;
	wire new_net_4061;
	wire new_net_5176;
	wire new_net_6067;
	wire new_net_4760;
	wire new_net_8507;
	wire new_net_10396;
	wire new_net_7047;
	wire new_net_7742;
	wire new_net_9925;
	wire new_net_6358;
	wire new_net_8562;
	wire new_net_6246;
	wire new_net_7907;
	wire new_net_459;
	wire new_net_1549;
	wire new_net_2652;
	wire new_net_2901;
	wire new_net_3283;
	wire new_net_3141;
	wire new_net_3777;
	wire new_net_4255;
	wire new_net_4559;
	wire new_net_4619;
	wire new_net_6184;
	wire new_net_6457;
	wire new_net_8081;
	wire new_net_7705;
	wire new_net_10524;
	wire new_net_6966;
	wire new_net_8280;
	wire new_net_10333;
	wire new_net_5748;
	wire n_0100_;
	wire n_1108_;
	wire n_0604_;
	wire new_net_724;
	wire new_net_3361;
	wire new_net_871;
	wire new_net_3385;
	wire new_net_4420;
	wire new_net_5799;
	wire new_net_6900;
	wire new_net_10659;
	wire new_net_5575;
	wire new_net_5469;
	wire new_net_7063;
	wire new_net_10087;
	wire new_net_7156;
	wire new_net_8596;
	wire new_net_9449;
	wire new_net_2324;
	wire new_net_1137;
	wire new_net_1170;
	wire new_net_3519;
	wire new_net_4637;
	wire new_net_4682;
	wire new_net_4706;
	wire new_net_4203;
	wire new_net_5156;
	wire new_net_5195;
	wire new_net_7154;
	wire new_net_9722;
	wire new_net_10242;
	wire new_net_9387;
	wire new_net_10679;
	wire new_net_7671;
	wire new_net_8956;
	wire n_0605_;
	wire n_0101_;
	wire n_1109_;
	wire new_net_1810;
	wire new_net_3275;
	wire new_net_339;
	wire new_net_1054;
	wire new_net_1957;
	wire new_net_5760;
	wire new_net_5784;
	wire new_net_7546;
	wire new_net_6154;
	wire new_net_8127;
	wire new_net_10426;
	wire new_net_6485;
	wire new_net_6478;
	wire new_net_676;
	wire new_net_1550;
	wire new_net_2566;
	wire new_net_2719;
	wire new_net_3081;
	wire new_net_3755;
	wire new_net_4016;
	wire new_net_4231;
	wire new_net_5340;
	wire new_net_5364;
	wire new_net_5663;
	wire new_net_6656;
	wire new_net_9610;
	wire new_net_9486;
	wire new_net_9297;
	wire new_net_5355;
	wire n_0606_;
	wire n_0102_;
	wire n_1110_;
	wire new_net_3100;
	wire new_net_41;
	wire new_net_872;
	wire new_net_5928;
	wire new_net_7110;
	wire new_net_7134;
	wire new_net_7193;
	wire new_net_9316;
	wire new_net_9979;
	wire new_net_9044;
	wire new_net_9236;
	wire new_net_2293;
	wire new_net_1138;
	wire new_net_2230;
	wire new_net_2461;
	wire new_net_4062;
	wire new_net_4693;
	wire new_net_5177;
	wire new_net_5621;
	wire new_net_6068;
	wire new_net_6702;
	wire new_net_7847;
	wire new_net_8020;
	wire new_net_7236;
	wire new_net_8553;
	wire new_net_8892;
	wire new_net_4401;
	wire new_net_6237;
	wire new_net_2137;
	wire n_1111_;
	wire n_0103_;
	wire n_0607_;
	wire new_net_460;
	wire new_net_2109;
	wire new_net_2489;
	wire new_net_2588;
	wire new_net_2902;
	wire new_net_3284;
	wire new_net_3971;
	wire new_net_8072;
	wire new_net_8354;
	wire new_net_8988;
	wire new_net_8986;
	wire new_net_6626;
	wire new_net_9776;
	wire new_net_8327;
	wire new_net_3386;
	wire new_net_677;
	wire new_net_725;
	wire new_net_3362;
	wire new_net_4421;
	wire new_net_5800;
	wire new_net_6886;
	wire new_net_7841;
	wire new_net_8166;
	wire new_net_5284;
	wire new_net_9184;
	wire new_net_5566;
	wire new_net_5460;
	wire new_net_7054;
	wire new_net_10257;
	wire new_net_6302;
	wire new_net_9087;
	wire new_net_9329;
	wire new_net_6442;
	wire n_1112_;
	wire n_0104_;
	wire new_net_2653;
	wire new_net_13;
	wire new_net_1171;
	wire new_net_42;
	wire new_net_2765;
	wire n_0608_;
	wire new_net_3520;
	wire new_net_4638;
	wire new_net_6734;
	wire new_net_4786;
	wire new_net_9201;
	wire new_net_6012;
	wire new_net_340;
	wire new_net_1139;
	wire new_net_1811;
	wire new_net_2325;
	wire n_0718_;
	wire new_net_4694;
	wire new_net_5761;
	wire new_net_5785;
	wire new_net_6329;
	wire new_net_6796;
	wire new_net_6922;
	wire new_net_8451;
	wire new_net_6850;
	wire new_net_9428;
	wire new_net_7015;
	wire new_net_1959;
	wire n_0609_;
	wire n_0105_;
	wire n_1113_;
	wire new_net_1551;
	wire new_net_461;
	wire new_net_2720;
	wire new_net_3082;
	wire new_net_1056;
	wire new_net_2085;
	wire new_net_5654;
	wire new_net_7926;
	wire new_net_7924;
	wire new_net_8361;
	wire new_net_10496;
	wire new_net_8677;
	wire new_net_5341;
	wire new_net_6574;
	wire new_net_9808;
	wire new_net_6567;
	wire new_net_8531;
	wire new_net_678;
	wire new_net_726;
	wire new_net_873;
	wire new_net_2143;
	wire new_net_3101;
	wire new_net_5929;
	wire new_net_7111;
	wire new_net_7135;
	wire new_net_7194;
	wire new_net_7443;
	wire new_net_4798;
	wire new_net_10480;
	wire new_net_7576;
	wire new_net_7869;
	wire new_net_9416;
	wire new_net_5119;
	wire new_net_7373;
	wire n_0610_;
	wire n_0106_;
	wire n_1114_;
	wire new_net_14;
	wire new_net_1172;
	wire new_net_3479;
	wire new_net_43;
	wire new_net_4063;
	wire new_net_5178;
	wire new_net_5622;
	wire new_net_8489;
	wire new_net_7719;
	wire new_net_8372;
	wire new_net_7717;
	wire new_net_5095;
	wire new_net_7227;
	wire new_net_8544;
	wire new_net_3143;
	wire new_net_341;
	wire new_net_2124;
	wire new_net_2294;
	wire new_net_1812;
	wire new_net_2623;
	wire new_net_2903;
	wire new_net_2462;
	wire new_net_3285;
	wire new_net_2231;
	wire new_net_9673;
	wire new_net_8114;
	wire new_net_9767;
	wire new_net_4604;
	wire new_net_2766;
	wire new_net_1960;
	wire new_net_3363;
	wire n_1115_;
	wire n_0611_;
	wire n_0107_;
	wire new_net_3387;
	wire new_net_1552;
	wire new_net_2111;
	wire new_net_4422;
	wire new_net_6877;
	wire new_net_7416;
	wire new_net_7040;
	wire new_net_8873;
	wire new_net_6293;
	wire new_net_10137;
	wire new_net_5608;
	wire new_net_4379;
	wire new_net_7138;
	wire new_net_3521;
	wire new_net_874;
	wire new_net_2654;
	wire new_net_4180;
	wire new_net_4639;
	wire new_net_4708;
	wire new_net_5283;
	wire new_net_8046;
	wire new_net_8068;
	wire new_net_9203;
	wire new_net_4902;
	wire new_net_9369;
	wire new_net_4900;
	wire new_net_7648;
	wire new_net_9168;
	wire new_net_44;
	wire n_1116_;
	wire n_0108_;
	wire n_0612_;
	wire new_net_1140;
	wire new_net_1173;
	wire new_net_4727;
	wire new_net_5762;
	wire new_net_5786;
	wire new_net_7071;
	wire new_net_5149;
	wire new_net_7332;
	wire new_net_8219;
	wire new_net_7496;
	wire new_net_6836;
	wire new_net_7494;
	wire new_net_10017;
	wire new_net_4849;
	wire new_net_1057;
	wire new_net_2326;
	wire new_net_1813;
	wire new_net_3083;
	wire new_net_3757;
	wire new_net_4018;
	wire new_net_5342;
	wire new_net_5366;
	wire new_net_6151;
	wire new_net_6575;
	wire new_net_8915;
	wire new_net_10651;
	wire new_net_5538;
	wire new_net_9907;
	wire new_net_4584;
	wire new_net_9274;
	wire new_net_6359;
	wire new_net_10074;
	wire new_net_5332;
	wire new_net_9799;
	wire new_net_3102;
	wire n_0613_;
	wire n_1117_;
	wire n_0109_;
	wire new_net_679;
	wire new_net_1553;
	wire new_net_5930;
	wire new_net_7112;
	wire new_net_7136;
	wire new_net_7195;
	wire new_net_6045;
	wire new_net_8227;
	wire new_net_4437;
	wire new_net_8225;
	wire new_net_6709;
	wire new_net_875;
	wire new_net_4064;
	wire new_net_4683;
	wire new_net_6070;
	wire new_net_6704;
	wire new_net_7402;
	wire new_net_7535;
	wire new_net_9458;
	wire new_net_9738;
	wire new_net_9900;
	wire new_net_3800;
	wire new_net_5086;
	wire new_net_4774;
	wire new_net_6214;
	wire new_net_3949;
	wire new_net_7759;
	wire new_net_9081;
	wire new_net_10292;
	wire new_net_3286;
	wire new_net_2904;
	wire new_net_342;
	wire n_0614_;
	wire n_1118_;
	wire n_0110_;
	wire new_net_3144;
	wire new_net_1141;
	wire new_net_1174;
	wire new_net_3780;
	wire new_net_4142;
	wire new_net_8051;
	wire new_net_8586;
	wire new_net_8584;
	wire new_net_9753;
	wire new_net_10038;
	wire new_net_9570;
	wire new_net_4590;
	wire new_net_8304;
	wire new_net_8936;
	wire new_net_9569;
	wire new_net_9562;
	wire new_net_10150;
	wire new_net_7818;
	wire new_net_2463;
	wire new_net_3480;
	wire new_net_15;
	wire new_net_463;
	wire new_net_1058;
	wire new_net_2232;
	wire new_net_3364;
	wire new_net_2295;
	wire new_net_1814;
	wire new_net_3388;
	wire new_net_7816;
	wire new_net_9966;
	wire new_net_9893;
	wire new_net_6279;
	wire new_net_5394;
	wire new_net_5599;
	wire new_net_7456;
	wire new_net_5493;
	wire new_net_7087;
	wire n_1119_;
	wire n_0615_;
	wire n_0111_;
	wire new_net_3522;
	wire new_net_2166;
	wire new_net_680;
	wire new_net_1554;
	wire new_net_2110;
	wire new_net_4640;
	wire new_net_4709;
	wire new_net_7179;
	wire new_net_10452;
	wire new_net_6767;
	wire new_net_6400;
	wire new_net_9360;
	wire new_net_10614;
	wire new_net_8816;
	wire new_net_45;
	wire new_net_2161;
	wire new_net_5763;
	wire new_net_5787;
	wire new_net_7072;
	wire new_net_7238;
	wire new_net_7262;
	wire new_net_8508;
	wire new_net_8555;
	wire new_net_5135;
	wire new_net_7318;
	wire new_net_5036;
	wire new_net_3645;
	wire new_net_8789;
	wire new_net_6827;
	wire new_net_4837;
	wire new_net_4239;
	wire new_net_6955;
	wire new_net_1175;
	wire new_net_3084;
	wire n_1120_;
	wire n_0616_;
	wire n_0112_;
	wire new_net_343;
	wire new_net_2767;
	wire new_net_3758;
	wire new_net_4019;
	wire new_net_5343;
	wire new_net_5631;
	wire new_net_10140;
	wire new_net_8727;
	wire new_net_10249;
	wire new_net_9510;
	wire new_net_9147;
	wire new_net_9707;
	wire new_net_3103;
	wire new_net_2327;
	wire new_net_5931;
	wire new_net_7113;
	wire new_net_7137;
	wire new_net_7196;
	wire new_net_7445;
	wire new_net_6607;
	wire new_net_9003;
	wire new_net_9471;
	wire new_net_6605;
	wire new_net_6695;
	wire new_net_7357;
	wire new_net_7609;
	wire n_1121_;
	wire n_0113_;
	wire n_0617_;
	wire new_net_876;
	wire new_net_681;
	wire new_net_4065;
	wire new_net_6071;
	wire new_net_6705;
	wire new_net_7403;
	wire new_net_8468;
	wire new_net_8720;
	wire new_net_9253;
	wire new_net_10406;
	wire new_net_8522;
	wire new_net_8162;
	wire new_net_9657;
	wire new_net_4324;
	wire new_net_8398;
	wire new_net_9650;
	wire new_net_2905;
	wire new_net_46;
	wire new_net_1142;
	wire new_net_3287;
	wire new_net_3145;
	wire new_net_2138;
	wire new_net_3781;
	wire new_net_4235;
	wire new_net_4259;
	wire new_net_4563;
	wire new_net_6256;
	wire new_net_7260;
	wire new_net_8838;
	wire new_net_8775;
	wire new_net_622;
	wire new_net_4201;
	wire new_net_8295;
	wire new_net_10428;
	wire new_net_4984;
	wire new_net_6854;
	wire new_net_9437;
	wire n_0114_;
	wire n_1122_;
	wire n_0618_;
	wire new_net_3481;
	wire new_net_1059;
	wire new_net_3365;
	wire new_net_3389;
	wire new_net_464;
	wire new_net_1815;
	wire new_net_4424;
	wire new_net_9879;
	wire new_net_6910;
	wire new_net_7237;
	wire new_net_5590;
	wire new_net_9027;
	wire new_net_2296;
	wire new_net_16;
	wire new_net_729;
	wire new_net_1555;
	wire new_net_2464;
	wire new_net_2233;
	wire new_net_3523;
	wire new_net_4641;
	wire new_net_4710;
	wire new_net_5158;
	wire new_net_5980;
	wire new_net_6758;
	wire new_net_7409;
	wire new_net_10605;
	wire new_net_5446;
	wire new_net_8244;
	wire new_net_10689;
	wire n_0115_;
	wire n_0619_;
	wire n_1123_;
	wire new_net_877;
	wire new_net_2136;
	wire new_net_4728;
	wire new_net_5764;
	wire new_net_5788;
	wire new_net_7073;
	wire new_net_7239;
	wire new_net_7681;
	wire new_net_6164;
	wire new_net_9401;
	wire new_net_5683;
	wire new_net_6946;
	wire new_net_344;
	wire new_net_1143;
	wire new_net_1176;
	wire new_net_3085;
	wire new_net_2768;
	wire new_net_3759;
	wire new_net_4020;
	wire new_net_5344;
	wire new_net_5368;
	wire new_net_6153;
	wire new_net_7527;
	wire new_net_10315;
	wire new_net_5520;
	wire new_net_7950;
	wire new_net_10429;
	wire new_net_10124;
	wire new_net_9496;
	wire new_net_9587;
	wire new_net_465;
	wire new_net_1816;
	wire n_0116_;
	wire n_1124_;
	wire n_0620_;
	wire new_net_3104;
	wire new_net_1060;
	wire new_net_5365;
	wire new_net_5932;
	wire new_net_6486;
	wire new_net_6591;
	wire new_net_8135;
	wire new_net_9989;
	wire new_net_9626;
	wire new_net_4822;
	wire new_net_8670;
	wire new_net_7600;
	wire new_net_5096;
	wire new_net_7893;
	wire new_net_7886;
	wire new_net_682;
	wire new_net_730;
	wire new_net_1556;
	wire new_net_2328;
	wire new_net_2655;
	wire new_net_4066;
	wire new_net_4729;
	wire new_net_5251;
	wire new_net_6072;
	wire new_net_6706;
	wire new_net_7397;
	wire new_net_10397;
	wire new_net_7743;
	wire new_net_9928;
	wire new_net_9926;
	wire n_0117_;
	wire n_1125_;
	wire n_0621_;
	wire new_net_2906;
	wire new_net_3288;
	wire new_net_47;
	wire new_net_3146;
	wire new_net_878;
	wire new_net_3782;
	wire new_net_4236;
	wire new_net_7908;
	wire new_net_10525;
	wire new_net_345;
	wire new_net_1177;
	wire new_net_2721;
	wire new_net_3482;
	wire new_net_3366;
	wire new_net_3390;
	wire new_net_4425;
	wire new_net_5749;
	wire new_net_5804;
	wire new_net_8170;
	wire new_net_3858;
	wire new_net_8326;
	wire new_net_6901;
	wire new_net_5576;
	wire new_net_9636;
	wire new_net_7064;
	wire new_net_6312;
	wire new_net_466;
	wire n_0622_;
	wire n_0118_;
	wire n_1126_;
	wire new_net_2033;
	wire new_net_1061;
	wire new_net_3524;
	wire new_net_4642;
	wire new_net_4711;
	wire new_net_5286;
	wire new_net_7157;
	wire new_net_9450;
	wire new_net_9723;
	wire new_net_6744;
	wire new_net_5221;
	wire new_net_4204;
	wire new_net_9612;
	wire new_net_6543;
	wire new_net_9388;
	wire new_net_10680;
	wire n_0590_;
	wire new_net_2656;
	wire new_net_683;
	wire new_net_731;
	wire new_net_1557;
	wire new_net_2465;
	wire new_net_2234;
	wire new_net_2297;
	wire new_net_5765;
	wire new_net_5789;
	wire new_net_7074;
	wire new_net_7672;
	wire new_net_5013;
	wire new_net_8957;
	wire new_net_10105;
	wire new_net_7547;
	wire new_net_6155;
	wire new_net_4219;
	wire new_net_9279;
	wire n_0119_;
	wire n_0623_;
	wire new_net_1144;
	wire new_net_2722;
	wire new_net_3086;
	wire n_1127_;
	wire new_net_48;
	wire new_net_2769;
	wire new_net_3207;
	wire new_net_4021;
	wire new_net_6479;
	wire new_net_6657;
	wire new_net_4440;
	wire new_net_5664;
	wire new_net_4438;
	wire new_net_9487;
	wire new_net_9298;
	wire new_net_1817;
	wire new_net_3105;
	wire new_net_5933;
	wire new_net_7115;
	wire new_net_7139;
	wire new_net_7198;
	wire new_net_5356;
	wire new_net_7447;
	wire new_net_9005;
	wire new_net_9175;
	wire n_0721_;
	wire new_net_10361;
	wire new_net_9980;
	wire new_net_7474;
	wire new_net_4813;
	wire new_net_6679;
	wire new_net_5050;
	wire new_net_7586;
	wire new_net_9045;
	wire new_net_2122;
	wire new_net_467;
	wire n_1128_;
	wire n_0120_;
	wire n_0624_;
	wire new_net_1062;
	wire new_net_4067;
	wire n_1071_;
	wire new_net_4730;
	wire new_net_5198;
	wire new_net_8335;
	wire new_net_9237;
	wire new_net_4748;
	wire new_net_8499;
	wire new_net_8021;
	wire new_net_3147;
	wire new_net_2329;
	wire new_net_732;
	wire new_net_879;
	wire new_net_2907;
	wire new_net_3289;
	wire new_net_3783;
	wire new_net_4237;
	wire new_net_4261;
	wire new_net_4402;
	wire new_net_6238;
	wire new_net_8893;
	wire new_net_3972;
	wire new_net_7780;
	wire new_net_8989;
	wire new_net_8073;
	wire new_net_8609;
	wire new_net_6627;
	wire new_net_9777;
	wire new_net_8937;
	wire new_net_3391;
	wire new_net_3367;
	wire n_0121_;
	wire n_1129_;
	wire n_0625_;
	wire new_net_1178;
	wire new_net_3483;
	wire new_net_346;
	wire new_net_2113;
	wire new_net_2036;
	wire new_net_8328;
	wire new_net_6887;
	wire new_net_10174;
	wire new_net_9185;
	wire new_net_7842;
	wire new_net_5285;
	wire new_net_5278;
	wire new_net_5567;
	wire new_net_5461;
	wire new_net_6303;
	wire new_net_3525;
	wire new_net_2118;
	wire new_net_17;
	wire new_net_1818;
	wire new_net_2116;
	wire new_net_4643;
	wire new_net_4712;
	wire new_net_5159;
	wire new_net_5287;
	wire new_net_8050;
	wire new_net_6443;
	wire new_net_9330;
	wire new_net_9202;
	wire new_net_8230;
	wire new_net_7203;
	wire new_net_684;
	wire new_net_1558;
	wire new_net_2657;
	wire n_0626_;
	wire n_0122_;
	wire n_1130_;
	wire new_net_5199;
	wire new_net_5766;
	wire new_net_5790;
	wire new_net_7075;
	wire n_0166_;
	wire new_net_6923;
	wire new_net_8452;
	wire new_net_9429;
	wire new_net_1994;
	wire new_net_2298;
	wire new_net_49;
	wire new_net_880;
	wire new_net_2723;
	wire new_net_3087;
	wire new_net_2466;
	wire new_net_2235;
	wire new_net_2770;
	wire new_net_4022;
	wire new_net_4263;
	wire new_net_4859;
	wire new_net_10499;
	wire new_net_7927;
	wire new_net_9833;
	wire new_net_5655;
	wire new_net_8678;
	wire new_net_2144;
	wire n_0627_;
	wire n_0123_;
	wire n_1131_;
	wire new_net_1146;
	wire new_net_1179;
	wire new_net_3106;
	wire new_net_347;
	wire new_net_5160;
	wire new_net_5934;
	wire new_net_6568;
	wire new_net_4799;
	wire new_net_4157;
	wire new_net_4154;
	wire new_net_10481;
	wire new_net_7870;
	wire new_net_5235;
	wire new_net_9417;
	wire n_0591_;
	wire new_net_468;
	wire new_net_1063;
	wire new_net_4068;
	wire new_net_4731;
	wire new_net_6074;
	wire new_net_6708;
	wire new_net_7406;
	wire new_net_9223;
	wire new_net_8490;
	wire new_net_7720;
	wire new_net_8668;
	wire new_net_3810;
	wire new_net_4505;
	wire new_net_8545;
	wire new_net_733;
	wire new_net_3148;
	wire new_net_2625;
	wire n_1132_;
	wire n_0628_;
	wire n_0124_;
	wire new_net_685;
	wire new_net_1559;
	wire new_net_2908;
	wire new_net_3290;
	wire new_net_9674;
	wire new_net_4558;
	wire new_net_8059;
	wire new_net_4793;
	wire new_net_4556;
	wire new_net_9768;
	wire new_net_8115;
	wire new_net_4605;
	wire new_net_3392;
	wire new_net_50;
	wire new_net_2330;
	wire new_net_3368;
	wire new_net_4427;
	wire new_net_5806;
	wire new_net_8172;
	wire new_net_8196;
	wire new_net_8859;
	wire new_net_9361;
	wire new_net_9534;
	wire new_net_6878;
	wire new_net_8202;
	wire n_0722_;
	wire new_net_10445;
	wire new_net_7417;
	wire new_net_7410;
	wire new_net_5447;
	wire new_net_7041;
	wire new_net_8874;
	wire new_net_10138;
	wire new_net_3526;
	wire n_1133_;
	wire n_0125_;
	wire n_0629_;
	wire new_net_1819;
	wire new_net_2154;
	wire new_net_1180;
	wire new_net_3276;
	wire new_net_4380;
	wire new_net_4644;
	wire new_net_5503;
	wire new_net_6429;
	wire new_net_4181;
	wire new_net_5922;
	wire new_net_8749;
	wire new_net_9370;
	wire new_net_7649;
	wire new_net_18;
	wire new_net_2658;
	wire new_net_469;
	wire new_net_1064;
	wire new_net_3760;
	wire new_net_5623;
	wire new_net_5767;
	wire new_net_5791;
	wire new_net_7076;
	wire new_net_7242;
	wire new_net_4996;
	wire new_net_7497;
	wire new_net_8438;
	wire new_net_6837;
	wire new_net_7495;
	wire new_net_2771;
	wire new_net_881;
	wire n_0630_;
	wire n_1134_;
	wire n_0126_;
	wire new_net_734;
	wire new_net_2724;
	wire new_net_3088;
	wire new_net_4023;
	wire new_net_5347;
	wire new_net_7007;
	wire new_net_8916;
	wire new_net_5646;
	wire new_net_10652;
	wire new_net_9908;
	wire new_net_10188;
	wire new_net_9275;
	wire new_net_2467;
	wire new_net_2236;
	wire new_net_51;
	wire new_net_348;
	wire new_net_1147;
	wire new_net_2299;
	wire new_net_2160;
	wire new_net_2162;
	wire new_net_5161;
	wire new_net_5333;
	wire new_net_9800;
	wire new_net_10585;
	wire new_net_6046;
	wire new_net_5430;
	wire new_net_7568;
	wire n_0631_;
	wire n_0127_;
	wire n_1135_;
	wire new_net_1008;
	wire new_net_1820;
	wire new_net_2156;
	wire new_net_2102;
	wire new_net_1181;
	wire new_net_4069;
	wire new_net_5179;
	wire new_net_6710;
	wire new_net_9658;
	wire new_net_7536;
	wire new_net_9459;
	wire new_net_9739;
	wire new_net_9901;
	wire new_net_3291;
	wire new_net_3149;
	wire new_net_470;
	wire new_net_686;
	wire new_net_1065;
	wire new_net_2134;
	wire new_net_1560;
	wire new_net_2112;
	wire new_net_2909;
	wire new_net_3761;
	wire new_net_6215;
	wire new_net_7760;
	wire new_net_9952;
	wire new_net_8052;
	wire new_net_9950;
	wire new_net_10293;
	wire new_net_8587;
	wire new_net_8585;
	wire new_net_9754;
	wire new_net_10039;
	wire new_net_10264;
	wire new_net_8305;
	wire new_net_3369;
	wire n_1136_;
	wire n_0632_;
	wire n_0128_;
	wire new_net_882;
	wire new_net_3393;
	wire new_net_735;
	wire new_net_4428;
	wire new_net_5807;
	wire new_net_6088;
	wire new_net_7819;
	wire new_net_10151;
	wire new_net_9066;
	wire new_net_9967;
	wire new_net_9894;
	wire new_net_6280;
	wire new_net_4963;
	wire new_net_5600;
	wire new_net_7457;
	wire new_net_2626;
	wire new_net_3527;
	wire new_net_19;
	wire new_net_349;
	wire new_net_1148;
	wire new_net_2117;
	wire new_net_2331;
	wire new_net_4645;
	wire new_net_4686;
	wire new_net_4714;
	wire new_net_7088;
	wire new_net_7180;
	wire new_net_10453;
	wire new_net_6768;
	wire new_net_10615;
	wire n_1137_;
	wire n_0129_;
	wire n_0633_;
	wire new_net_2659;
	wire new_net_1821;
	wire new_net_4625;
	wire new_net_5768;
	wire new_net_5792;
	wire new_net_7077;
	wire new_net_7243;
	wire new_net_7319;
	wire new_net_5037;
	wire new_net_8228;
	wire new_net_8790;
	wire new_net_9148;
	wire new_net_6828;
	wire new_net_4242;
	wire new_net_2725;
	wire new_net_3089;
	wire new_net_2772;
	wire new_net_471;
	wire new_net_687;
	wire new_net_1066;
	wire new_net_1561;
	wire new_net_1997;
	wire new_net_4024;
	wire new_net_5348;
	wire new_net_9285;
	wire new_net_10095;
	wire new_net_8728;
	wire new_net_8998;
	wire new_net_10250;
	wire new_net_9150;
	wire new_net_4462;
	wire new_net_9511;
	wire new_net_736;
	wire n_0634_;
	wire n_1138_;
	wire n_0130_;
	wire new_net_883;
	wire new_net_4763;
	wire new_net_5162;
	wire new_net_5936;
	wire new_net_6089;
	wire new_net_7118;
	wire new_net_9708;
	wire new_net_10576;
	wire new_net_6608;
	wire new_net_10112;
	wire new_net_7556;
	wire new_net_4749;
	wire new_net_6606;
	wire new_net_6696;
	wire new_net_4482;
	wire new_net_2468;
	wire new_net_1149;
	wire new_net_1182;
	wire new_net_2300;
	wire new_net_2237;
	wire new_net_4520;
	wire new_net_4565;
	wire new_net_5074;
	wire new_net_5625;
	wire new_net_6076;
	wire new_net_8469;
	wire new_net_7407;
	wire new_net_7291;
	wire new_net_9254;
	wire new_net_10407;
	wire new_net_8523;
	wire new_net_2910;
	wire new_net_3292;
	wire n_0635_;
	wire n_1139_;
	wire n_0131_;
	wire new_net_3150;
	wire new_net_1822;
	wire new_net_3762;
	wire new_net_3786;
	wire new_net_4240;
	wire new_net_8399;
	wire new_net_9651;
	wire new_net_10564;
	wire new_net_7261;
	wire new_net_8776;
	wire new_net_5714;
	wire new_net_8296;
	wire new_net_3370;
	wire new_net_688;
	wire new_net_1562;
	wire new_net_4429;
	wire new_net_5808;
	wire new_net_8174;
	wire new_net_4985;
	wire new_net_6855;
	wire new_net_8198;
	wire new_net_8943;
	wire new_net_9438;
	wire new_net_10346;
	wire new_net_9880;
	wire new_net_6911;
	wire new_net_3736;
	wire new_net_5302;
	wire new_net_5591;
	wire new_net_7448;
	wire new_net_9028;
	wire new_net_2091;
	wire new_net_20;
	wire n_0636_;
	wire n_0132_;
	wire n_1140_;
	wire new_net_53;
	wire new_net_350;
	wire new_net_3528;
	wire new_net_884;
	wire new_net_4646;
	wire new_net_8203;
	wire new_net_5049;
	wire new_net_1150;
	wire new_net_1183;
	wire new_net_2332;
	wire new_net_2660;
	wire new_net_4566;
	wire new_net_4626;
	wire new_net_4732;
	wire new_net_5202;
	wire new_net_5769;
	wire new_net_5793;
	wire new_net_10690;
	wire new_net_472;
	wire new_net_1823;
	wire new_net_2726;
	wire new_net_3090;
	wire n_1141_;
	wire n_0637_;
	wire n_0133_;
	wire new_net_1067;
	wire new_net_2773;
	wire new_net_2141;
	wire new_net_5684;
	wire new_net_6947;
	wire new_net_7528;
	wire new_net_10316;
	wire new_net_5521;
	wire new_net_7951;
	wire new_net_10545;
	wire new_net_10125;
	wire new_net_9497;
	wire new_net_3484;
	wire new_net_689;
	wire new_net_737;
	wire new_net_4764;
	wire new_net_5163;
	wire new_net_5937;
	wire new_net_6090;
	wire new_net_7119;
	wire new_net_7143;
	wire new_net_7202;
	wire new_net_5409;
	wire new_net_8379;
	wire new_net_9588;
	wire new_net_6592;
	wire new_net_9990;
	wire new_net_4823;
	wire new_net_4506;
	wire new_net_6077;
	wire new_net_21;
	wire new_net_3108;
	wire n_1142_;
	wire n_0638_;
	wire n_0134_;
	wire new_net_351;
	wire new_net_4733;
	wire new_net_5097;
	wire new_net_5626;
	wire new_net_5880;
	wire new_net_7894;
	wire new_net_9117;
	wire new_net_10506;
	wire new_net_8509;
	wire new_net_10398;
	wire new_net_7744;
	wire new_net_9929;
	wire new_net_2911;
	wire new_net_2469;
	wire new_net_3293;
	wire new_net_2238;
	wire new_net_3151;
	wire new_net_2125;
	wire new_net_2301;
	wire new_net_3763;
	wire new_net_3787;
	wire new_net_4241;
	wire new_net_9927;
	wire new_net_8564;
	wire new_net_6248;
	wire new_net_6186;
	wire new_net_8083;
	wire new_net_10526;
	wire new_net_6968;
	wire new_net_8282;
	wire new_net_8534;
	wire new_net_795;
	wire new_net_6115;
	wire new_net_5750;
	wire new_net_8338;
	wire new_net_6902;
	wire new_net_4350;
	wire new_net_10661;
	wire new_net_5577;
	wire new_net_9637;
	wire new_net_5471;
	wire new_net_7065;
	wire new_net_6313;
	wire new_net_10089;
	wire new_net_902;
	wire new_net_3011;
	wire new_net_524;
	wire n_1185_;
	wire n_0177_;
	wire n_0387_;
	wire n_0891_;
	wire new_net_1200;
	wire n_0681_;
	wire new_net_3664;
	wire new_net_6745;
	wire new_net_9340;
	wire new_net_4205;
	wire new_net_9613;
	wire new_net_9748;
	wire new_net_9389;
	wire new_net_7673;
	wire new_net_8958;
	wire new_net_639;
	wire new_net_789;
	wire new_net_1498;
	wire new_net_1840;
	wire new_net_2602;
	wire new_net_4481;
	wire new_net_5014;
	wire new_net_5073;
	wire new_net_5142;
	wire new_net_7585;
	wire new_net_7548;
	wire new_net_6156;
	wire new_net_6487;
	wire new_net_3552;
	wire new_net_1580;
	wire new_net_2673;
	wire new_net_2859;
	wire n_0892_;
	wire new_net_223;
	wire n_0178_;
	wire n_0388_;
	wire n_0682_;
	wire new_net_265;
	wire new_net_6658;
	wire new_net_5665;
	wire new_net_9574;
	wire new_net_9299;
	wire new_net_2396;
	wire new_net_2693;
	wire new_net_3055;
	wire new_net_368;
	wire new_net_755;
	wire new_net_3250;
	wire new_net_3944;
	wire new_net_3967;
	wire new_net_3991;
	wire new_net_4191;
	wire new_net_5357;
	wire new_net_10362;
	wire new_net_9981;
	wire new_net_6680;
	wire new_net_6389;
	wire new_net_5051;
	wire new_net_7587;
	wire new_net_9046;
	wire n_0683_;
	wire new_net_2105;
	wire new_net_936;
	wire n_0893_;
	wire new_net_2881;
	wire n_0179_;
	wire n_0389_;
	wire new_net_525;
	wire new_net_1201;
	wire n_1187_;
	wire new_net_9238;
	wire new_net_8500;
	wire new_net_7730;
	wire new_net_8022;
	wire new_net_8894;
	wire new_net_2635;
	wire new_net_1382;
	wire new_net_3618;
	wire new_net_640;
	wire new_net_790;
	wire new_net_1349;
	wire new_net_1499;
	wire new_net_3642;
	wire new_net_4439;
	wire new_net_4658;
	wire new_net_6239;
	wire new_net_7781;
	wire new_net_8990;
	wire new_net_8074;
	wire new_net_8610;
	wire new_net_6628;
	wire new_net_9778;
	wire new_net_8329;
	wire n_0684_;
	wire new_net_224;
	wire new_net_3235;
	wire n_0894_;
	wire n_1188_;
	wire n_0180_;
	wire n_0390_;
	wire new_net_266;
	wire new_net_3338;
	wire new_net_5092;
	wire new_net_6888;
	wire new_net_7843;
	wire new_net_9186;
	wire new_net_10175;
	wire new_net_5568;
	wire new_net_6304;
	wire new_net_1963;
	wire new_net_3012;
	wire new_net_2365;
	wire new_net_369;
	wire new_net_903;
	wire new_net_2094;
	wire new_net_2428;
	wire new_net_2197;
	wire new_net_2470;
	wire new_net_3665;
	wire new_net_6736;
	wire new_net_9331;
	wire new_net_6014;
	wire new_net_7204;
	wire new_net_7197;
	wire n_1189_;
	wire new_net_2145;
	wire n_0685_;
	wire new_net_937;
	wire n_0181_;
	wire n_0391_;
	wire n_0895_;
	wire new_net_1841;
	wire new_net_526;
	wire new_net_2603;
	wire new_net_6798;
	wire new_net_8453;
	wire new_net_9430;
	wire new_net_3229;
	wire new_net_2101;
	wire new_net_1350;
	wire new_net_1383;
	wire new_net_2860;
	wire new_net_2674;
	wire new_net_3851;
	wire new_net_4264;
	wire new_net_4580;
	wire new_net_5012;
	wire new_net_7017;
	wire new_net_7928;
	wire new_net_9834;
	wire new_net_5656;
	wire new_net_10402;
	wire new_net_6576;
	wire new_net_9810;
	wire n_1190_;
	wire new_net_3056;
	wire n_0686_;
	wire n_0182_;
	wire n_0392_;
	wire new_net_2694;
	wire n_0896_;
	wire new_net_225;
	wire new_net_267;
	wire new_net_756;
	wire new_net_4158;
	wire new_net_4155;
	wire new_net_7578;
	wire new_net_7871;
	wire new_net_9418;
	wire new_net_9224;
	wire new_net_2505;
	wire new_net_904;
	wire new_net_1202;
	wire new_net_2397;
	wire new_net_2882;
	wire new_net_3317;
	wire new_net_5951;
	wire new_net_6128;
	wire new_net_7216;
	wire new_net_7631;
	wire new_net_9827;
	wire new_net_8134;
	wire new_net_7721;
	wire new_net_8669;
	wire new_net_6339;
	wire n_0929_;
	wire new_net_7229;
	wire new_net_8546;
	wire n_1191_;
	wire new_net_1500;
	wire n_0393_;
	wire new_net_641;
	wire new_net_2636;
	wire n_0687_;
	wire n_0183_;
	wire n_0897_;
	wire new_net_1842;
	wire new_net_527;
	wire new_net_9059;
	wire new_net_9675;
	wire new_net_8116;
	wire new_net_9769;
	wire new_net_5738;
	wire new_net_9535;
	wire new_net_3339;
	wire new_net_2120;
	wire new_net_1582;
	wire new_net_5607;
	wire new_net_6352;
	wire new_net_7340;
	wire new_net_6879;
	wire new_net_7829;
	wire new_net_7876;
	wire new_net_7900;
	wire new_net_8311;
	wire new_net_7418;
	wire new_net_5448;
	wire new_net_7042;
	wire new_net_8875;
	wire new_net_6295;
	wire new_net_10139;
	wire new_net_8532;
	wire new_net_5610;
	wire new_net_4381;
	wire new_net_7140;
	wire new_net_9317;
	wire n_1192_;
	wire new_net_370;
	wire n_0688_;
	wire new_net_3013;
	wire n_0184_;
	wire n_0394_;
	wire n_0898_;
	wire new_net_226;
	wire new_net_268;
	wire new_net_757;
	wire new_net_4182;
	wire new_net_8336;
	wire n_0790_;
	wire new_net_4904;
	wire new_net_8750;
	wire new_net_9371;
	wire new_net_7650;
	wire new_net_1203;
	wire new_net_2198;
	wire new_net_2471;
	wire new_net_2604;
	wire new_net_1728;
	wire new_net_905;
	wire new_net_938;
	wire new_net_2366;
	wire new_net_2429;
	wire new_net_4483;
	wire new_net_5151;
	wire new_net_8439;
	wire new_net_6838;
	wire n_0595_;
	wire new_net_10019;
	wire new_net_792;
	wire new_net_1501;
	wire n_0395_;
	wire n_0689_;
	wire new_net_642;
	wire new_net_3554;
	wire n_0899_;
	wire n_1193_;
	wire n_0185_;
	wire new_net_2861;
	wire new_net_6327;
	wire new_net_8917;
	wire new_net_8839;
	wire new_net_10653;
	wire new_net_5540;
	wire new_net_10189;
	wire new_net_9276;
	wire new_net_5334;
	wire new_net_9801;
	wire new_net_1965;
	wire new_net_1583;
	wire new_net_2695;
	wire new_net_3057;
	wire new_net_3252;
	wire new_net_3946;
	wire new_net_3969;
	wire new_net_3993;
	wire new_net_4193;
	wire new_net_4294;
	wire new_net_5433;
	wire new_net_7100;
	wire new_net_7728;
	wire new_net_10276;
	wire new_net_10586;
	wire new_net_6047;
	wire new_net_7569;
	wire new_net_1009;
	wire new_net_1652;
	wire new_net_6711;
	wire new_net_2584;
	wire n_1194_;
	wire new_net_371;
	wire n_0690_;
	wire n_0186_;
	wire n_0396_;
	wire n_0900_;
	wire new_net_227;
	wire new_net_269;
	wire new_net_5904;
	wire new_net_9460;
	wire new_net_9740;
	wire new_net_9902;
	wire new_net_6330;
	wire new_net_5088;
	wire new_net_8175;
	wire new_net_6216;
	wire new_net_9953;
	wire new_net_1729;
	wire new_net_528;
	wire new_net_906;
	wire new_net_939;
	wire new_net_1843;
	wire new_net_2398;
	wire new_net_3620;
	wire new_net_3644;
	wire new_net_3951;
	wire new_net_4441;
	wire new_net_7761;
	wire new_net_8053;
	wire new_net_8588;
	wire new_net_9951;
	wire new_net_9755;
	wire new_net_10040;
	wire new_net_4592;
	wire new_net_10265;
	wire new_net_8306;
	wire new_net_8938;
	wire new_net_3318;
	wire n_1195_;
	wire new_net_1502;
	wire new_net_2058;
	wire n_0397_;
	wire new_net_643;
	wire new_net_2077;
	wire new_net_3340;
	wire n_0691_;
	wire n_0187_;
	wire new_net_2583;
	wire new_net_6139;
	wire new_net_7820;
	wire new_net_9067;
	wire new_net_9095;
	wire new_net_9968;
	wire new_net_8355;
	wire new_net_5398;
	wire new_net_9895;
	wire new_net_6281;
	wire new_net_5396;
	wire new_net_4964;
	wire new_net_5601;
	wire new_net_7458;
	wire new_net_5495;
	wire new_net_7089;
	wire new_net_758;
	wire new_net_3014;
	wire new_net_1584;
	wire new_net_3667;
	wire new_net_6257;
	wire new_net_6307;
	wire new_net_10418;
	wire new_net_10633;
	wire new_net_7181;
	wire new_net_10618;
	wire new_net_6769;
	wire new_net_9627;
	wire new_net_8436;
	wire new_net_9362;
	wire new_net_10616;
	wire new_net_270;
	wire new_net_1204;
	wire new_net_2605;
	wire n_1196_;
	wire new_net_372;
	wire n_0398_;
	wire n_0692_;
	wire n_0188_;
	wire n_0902_;
	wire new_net_228;
	wire new_net_7917;
	wire new_net_5137;
	wire new_net_7320;
	wire new_net_7984;
	wire new_net_8229;
	wire new_net_6829;
	wire new_net_1844;
	wire new_net_3231;
	wire new_net_2430;
	wire new_net_2199;
	wire new_net_2472;
	wire new_net_1967;
	wire new_net_3555;
	wire new_net_529;
	wire new_net_793;
	wire new_net_907;
	wire new_net_5633;
	wire new_net_10096;
	wire new_net_8729;
	wire new_net_8999;
	wire new_net_7706;
	wire new_net_10251;
	wire new_net_9151;
	wire new_net_9149;
	wire new_net_2696;
	wire new_net_3253;
	wire n_0189_;
	wire new_net_3058;
	wire n_0903_;
	wire n_1197_;
	wire n_0399_;
	wire n_0693_;
	wire new_net_644;
	wire new_net_1353;
	wire new_net_9598;
	wire new_net_10577;
	wire new_net_6609;
	wire new_net_10113;
	wire new_net_6266;
	wire new_net_7557;
	wire new_net_5075;
	wire new_net_6697;
	wire new_net_7359;
	wire new_net_7611;
	wire new_net_8266;
	wire new_net_2507;
	wire new_net_759;
	wire new_net_1585;
	wire new_net_5953;
	wire new_net_5972;
	wire new_net_6130;
	wire new_net_7218;
	wire new_net_8470;
	wire new_net_9025;
	wire new_net_9132;
	wire new_net_8722;
	wire new_net_7408;
	wire new_net_9255;
	wire new_net_10408;
	wire new_net_8524;
	wire new_net_8402;
	wire new_net_9659;
	wire new_net_4326;
	wire new_net_10565;
	wire new_net_229;
	wire new_net_3621;
	wire new_net_271;
	wire n_0190_;
	wire new_net_1205;
	wire new_net_373;
	wire new_net_1730;
	wire n_0904_;
	wire n_1198_;
	wire n_0400_;
	wire new_net_8265;
	wire new_net_8373;
	wire new_net_8777;
	wire new_net_5715;
	wire new_net_8297;
	wire new_net_10430;
	wire new_net_2675;
	wire new_net_2399;
	wire new_net_3319;
	wire new_net_3341;
	wire new_net_794;
	wire new_net_1386;
	wire new_net_1503;
	wire new_net_4210;
	wire new_net_5094;
	wire new_net_5609;
	wire new_net_6856;
	wire new_net_9881;
	wire new_net_4787;
	wire new_net_6912;
	wire new_net_3737;
	wire new_net_4360;
	wire new_net_5592;
	wire new_net_7449;
	wire new_net_6415;
	wire new_net_9029;
	wire new_net_10212;
	wire n_0191_;
	wire n_0695_;
	wire n_0905_;
	wire n_1199_;
	wire n_0401_;
	wire new_net_3015;
	wire new_net_3668;
	wire new_net_6258;
	wire new_net_10419;
	wire new_net_6505;
	wire new_net_7167;
	wire new_net_6503;
	wire new_net_6760;
	wire new_net_10691;
	wire new_net_2606;
	wire new_net_4485;
	wire new_net_5053;
	wire new_net_5077;
	wire new_net_5146;
	wire new_net_5973;
	wire new_net_7589;
	wire new_net_7613;
	wire new_net_7797;
	wire new_net_7683;
	wire new_net_7311;
	wire new_net_6166;
	wire new_net_8896;
	wire new_net_941;
	wire n_0906_;
	wire new_net_230;
	wire new_net_1845;
	wire new_net_3232;
	wire new_net_272;
	wire new_net_530;
	wire n_0192_;
	wire new_net_1206;
	wire n_0696_;
	wire new_net_7529;
	wire new_net_4283;
	wire new_net_5524;
	wire new_net_8895;
	wire new_net_10317;
	wire new_net_5522;
	wire new_net_7952;
	wire new_net_10126;
	wire new_net_9498;
	wire new_net_2106;
	wire new_net_2697;
	wire new_net_3059;
	wire new_net_1354;
	wire new_net_2368;
	wire new_net_2431;
	wire new_net_3254;
	wire new_net_2200;
	wire new_net_2473;
	wire new_net_645;
	wire new_net_5410;
	wire new_net_6031;
	wire new_net_5367;
	wire new_net_4684;
	wire new_net_9991;
	wire new_net_4824;
	wire n_0938_;
	wire new_net_3068;
	wire new_net_9522;
	wire new_net_4507;
	wire new_net_7602;
	wire new_net_5098;
	wire new_net_1586;
	wire new_net_760;
	wire n_0193_;
	wire n_0907_;
	wire n_1201_;
	wire n_0697_;
	wire n_0403_;
	wire new_net_2638;
	wire new_net_5253;
	wire new_net_5881;
	wire new_net_9089;
	wire new_net_10507;
	wire new_net_8980;
	wire new_net_8510;
	wire new_net_10399;
	wire new_net_7745;
	wire new_net_9451;
	wire new_net_9930;
	wire new_net_3622;
	wire new_net_2073;
	wire new_net_3646;
	wire new_net_4443;
	wire new_net_4662;
	wire new_net_5389;
	wire new_net_5413;
	wire new_net_5437;
	wire new_net_5667;
	wire new_net_6034;
	wire new_net_4121;
	wire new_net_6361;
	wire new_net_8565;
	wire new_net_8125;
	wire new_net_10529;
	wire new_net_9823;
	wire new_net_10527;
	wire new_net_909;
	wire new_net_231;
	wire new_net_1846;
	wire new_net_273;
	wire new_net_531;
	wire n_0194_;
	wire new_net_3320;
	wire n_0908_;
	wire n_1202_;
	wire new_net_375;
	wire new_net_6116;
	wire new_net_3860;
	wire new_net_6903;
	wire new_net_10662;
	wire n_0522_;
	wire new_net_164;
	wire new_net_5578;
	wire new_net_5472;
	wire new_net_8679;
	wire new_net_7066;
	wire new_net_6314;
	wire new_net_3016;
	wire new_net_1388;
	wire new_net_2400;
	wire new_net_796;
	wire new_net_646;
	wire new_net_1505;
	wire new_net_3669;
	wire new_net_3994;
	wire new_net_6259;
	wire new_net_8133;
	wire new_net_9452;
	wire new_net_10090;
	wire new_net_9341;
	wire new_net_4880;
	wire new_net_6746;
	wire new_net_4206;
	wire new_net_9614;
	wire new_net_10482;
	wire new_net_6545;
	wire new_net_9390;
	wire n_0405_;
	wire new_net_1587;
	wire new_net_761;
	wire n_0195_;
	wire n_0699_;
	wire n_0909_;
	wire n_1203_;
	wire new_net_2607;
	wire new_net_4486;
	wire new_net_4582;
	wire new_net_7674;
	wire new_net_8959;
	wire new_net_6328;
	wire new_net_374;
	wire new_net_5015;
	wire new_net_7549;
	wire new_net_4340;
	wire new_net_6808;
	wire new_net_4304;
	wire new_net_6157;
	wire new_net_4221;
	wire new_net_6934;
	wire new_net_3557;
	wire new_net_2864;
	wire new_net_3233;
	wire new_net_942;
	wire new_net_1207;
	wire new_net_1732;
	wire new_net_3855;
	wire new_net_5016;
	wire new_net_5264;
	wire new_net_6428;
	wire new_net_6488;
	wire new_net_6481;
	wire new_net_7938;
	wire new_net_6659;
	wire new_net_4442;
	wire new_net_5666;
	wire new_net_9575;
	wire new_net_9300;
	wire n_0406_;
	wire new_net_3255;
	wire new_net_232;
	wire new_net_1847;
	wire new_net_2698;
	wire new_net_3060;
	wire new_net_274;
	wire new_net_532;
	wire n_0196_;
	wire n_0700_;
	wire new_net_1653;
	wire new_net_5358;
	wire new_net_9177;
	wire new_net_10370;
	wire new_net_10363;
	wire new_net_9982;
	wire new_net_4815;
	wire new_net_6681;
	wire new_net_5052;
	wire new_net_7588;
	wire new_net_2639;
	wire new_net_1356;
	wire new_net_2369;
	wire new_net_1389;
	wire new_net_2432;
	wire new_net_2201;
	wire new_net_2474;
	wire new_net_2509;
	wire new_net_1506;
	wire new_net_4583;
	wire new_net_9047;
	wire n_1078_;
	wire new_net_9239;
	wire new_net_8501;
	wire new_net_7731;
	wire new_net_8023;
	wire n_0407_;
	wire new_net_3623;
	wire new_net_762;
	wire n_0911_;
	wire n_0701_;
	wire n_1205_;
	wire n_0197_;
	wire new_net_3647;
	wire new_net_4444;
	wire new_net_4663;
	wire new_net_8556;
	wire new_net_4404;
	wire new_net_6240;
	wire new_net_3974;
	wire new_net_8356;
	wire new_net_8991;
	wire new_net_8075;
	wire new_net_8611;
	wire new_net_9779;
	wire new_net_4618;
	wire new_net_5194;
	wire new_net_1733;
	wire new_net_910;
	wire new_net_943;
	wire new_net_1208;
	wire new_net_3343;
	wire new_net_4212;
	wire new_net_5611;
	wire new_net_6356;
	wire new_net_7344;
	wire new_net_7880;
	wire new_net_8330;
	wire new_net_1504;
	wire new_net_3714;
	wire new_net_6889;
	wire new_net_7844;
	wire new_net_9187;
	wire new_net_7428;
	wire new_net_8738;
	wire new_net_5569;
	wire new_net_8374;
	wire new_net_9909;
	wire new_net_6305;
	wire n_1206_;
	wire new_net_377;
	wire n_0702_;
	wire new_net_647;
	wire new_net_3017;
	wire n_0912_;
	wire new_net_233;
	wire new_net_1848;
	wire new_net_275;
	wire n_0198_;
	wire new_net_10076;
	wire new_net_9332;
	wire new_net_6737;
	wire new_net_4192;
	wire new_net_8597;
	wire new_net_4761;
	wire new_net_9204;
	wire new_net_7205;
	wire new_net_2988;
	wire new_net_1588;
	wire new_net_2401;
	wire new_net_1357;
	wire new_net_2608;
	wire new_net_4487;
	wire new_net_5055;
	wire new_net_5148;
	wire new_net_5975;
	wire new_net_7591;
	wire new_net_7615;
	wire new_net_6799;
	wire n_1323_;
	wire new_net_1779;
	wire new_net_1986;
	wire new_net_7339;
	wire new_net_7508;
	wire n_1207_;
	wire new_net_2059;
	wire new_net_3558;
	wire new_net_2865;
	wire n_0913_;
	wire new_net_3234;
	wire new_net_763;
	wire n_0703_;
	wire n_0199_;
	wire n_0409_;
	wire new_net_5204;
	wire new_net_7018;
	wire new_net_7929;
	wire new_net_5657;
	wire new_net_10267;
	wire new_net_2699;
	wire new_net_2883;
	wire new_net_3061;
	wire new_net_533;
	wire new_net_911;
	wire new_net_944;
	wire new_net_1734;
	wire new_net_3256;
	wire new_net_3950;
	wire new_net_3973;
	wire new_net_6577;
	wire new_net_6570;
	wire new_net_9811;
	wire new_net_4801;
	wire new_net_7579;
	wire new_net_5237;
	wire new_net_9419;
	wire n_1208_;
	wire new_net_378;
	wire new_net_1507;
	wire n_0704_;
	wire new_net_648;
	wire new_net_2640;
	wire n_0914_;
	wire new_net_234;
	wire n_0200_;
	wire n_0410_;
	wire new_net_9225;
	wire new_net_10456;
	wire new_net_4777;
	wire new_net_9828;
	wire new_net_10454;
	wire new_net_7722;
	wire new_net_3812;
	wire new_net_2370;
	wire new_net_3624;
	wire new_net_1589;
	wire new_net_2433;
	wire new_net_2202;
	wire new_net_2475;
	wire new_net_3648;
	wire new_net_4445;
	wire new_net_4664;
	wire new_net_5078;
	wire new_net_7230;
	wire new_net_7553;
	wire new_net_8426;
	wire new_net_8547;
	wire new_net_9060;
	wire new_net_9678;
	wire new_net_9676;
	wire new_net_1055;
	wire new_net_4560;
	wire new_net_8061;
	wire new_net_7281;
	wire new_net_9840;
	wire new_net_8791;
	wire new_net_7610;
	wire new_net_8117;
	wire new_net_1209;
	wire new_net_3344;
	wire n_0705_;
	wire n_0915_;
	wire n_1209_;
	wire n_0201_;
	wire n_0411_;
	wire new_net_4213;
	wire new_net_5612;
	wire new_net_6357;
	wire new_net_9536;
	wire new_net_9851;
	wire new_net_4036;
	wire new_net_7830;
	wire new_net_6880;
	wire new_net_8123;
	wire new_net_7419;
	wire new_net_7412;
	wire new_net_5449;
	wire new_net_8876;
	wire new_net_6296;
	wire new_net_8533;
	wire new_net_1968;
	wire new_net_3018;
	wire new_net_1849;
	wire new_net_2884;
	wire new_net_534;
	wire new_net_945;
	wire new_net_3671;
	wire new_net_4382;
	wire new_net_6261;
	wire new_net_7141;
	wire new_net_6431;
	wire new_net_9318;
	wire new_net_9709;
	wire new_net_8337;
	wire new_net_4183;
	wire new_net_4176;
	wire new_net_6529;
	wire new_net_8751;
	wire new_net_9372;
	wire new_net_799;
	wire new_net_2609;
	wire new_net_379;
	wire new_net_1508;
	wire n_0706_;
	wire new_net_649;
	wire new_net_2103;
	wire new_net_1358;
	wire n_0202_;
	wire n_0412_;
	wire new_net_7358;
	wire new_net_7651;
	wire new_net_8823;
	wire new_net_5152;
	wire new_net_7335;
	wire new_net_4081;
	wire new_net_7499;
	wire new_net_4079;
	wire new_net_8440;
	wire new_net_6839;
	wire new_net_3559;
	wire new_net_2866;
	wire new_net_764;
	wire new_net_2402;
	wire new_net_3857;
	wire new_net_4746;
	wire n_0320_;
	wire new_net_5018;
	wire new_net_5266;
	wire new_net_6430;
	wire new_net_6465;
	wire new_net_10106;
	wire new_net_5648;
	wire new_net_8840;
	wire new_net_5548;
	wire new_net_1391;
	wire new_net_10190;
	wire new_net_9277;
	wire new_net_1210;
	wire new_net_3321;
	wire n_1211_;
	wire new_net_1735;
	wire n_0707_;
	wire new_net_912;
	wire n_0203_;
	wire n_0413_;
	wire new_net_2013;
	wire n_0917_;
	wire new_net_5335;
	wire new_net_7108;
	wire new_net_9802;
	wire new_net_10347;
	wire new_net_10587;
	wire new_net_5434;
	wire new_net_6048;
	wire new_net_5432;
	wire new_net_7570;
	wire new_net_3328;
	wire new_net_2511;
	wire new_net_2641;
	wire new_net_535;
	wire new_net_1850;
	wire new_net_3841;
	wire new_net_5957;
	wire new_net_6134;
	wire new_net_7222;
	wire new_net_10536;
	wire new_net_5905;
	wire new_net_8204;
	wire new_net_9461;
	wire new_net_9741;
	wire new_net_3892;
	wire new_net_6331;
	wire new_net_8347;
	wire new_net_5089;
	wire new_net_8176;
	wire new_net_278;
	wire new_net_800;
	wire n_1212_;
	wire new_net_380;
	wire new_net_1359;
	wire new_net_1590;
	wire n_0708_;
	wire n_0204_;
	wire n_0414_;
	wire new_net_797;
	wire new_net_3670;
	wire new_net_6217;
	wire new_net_7762;
	wire new_net_9954;
	wire new_net_10295;
	wire new_net_8589;
	wire new_net_9756;
	wire new_net_165;
	wire new_net_8384;
	wire new_net_10041;
	wire new_net_10553;
	wire new_net_10266;
	wire new_net_2434;
	wire new_net_2203;
	wire new_net_2476;
	wire new_net_3345;
	wire new_net_765;
	wire new_net_1972;
	wire new_net_2371;
	wire new_net_4214;
	wire new_net_4747;
	wire new_net_5040;
	wire new_net_8939;
	wire new_net_7821;
	wire new_net_6140;
	wire new_net_9096;
	wire new_net_6298;
	wire new_net_9969;
	wire new_net_9896;
	wire new_net_9379;
	wire new_net_6282;
	wire new_net_3322;
	wire n_1213_;
	wire new_net_1736;
	wire n_0415_;
	wire n_0709_;
	wire new_net_913;
	wire new_net_2107;
	wire new_net_3019;
	wire n_0205_;
	wire new_net_946;
	wire new_net_5496;
	wire new_net_7090;
	wire new_net_10619;
	wire new_net_6770;
	wire new_net_9628;
	wire new_net_9363;
	wire new_net_10617;
	wire new_net_2016;
	wire new_net_2610;
	wire new_net_1509;
	wire new_net_650;
	wire new_net_1392;
	wire new_net_4489;
	wire new_net_5057;
	wire new_net_5150;
	wire new_net_5977;
	wire new_net_7593;
	wire new_net_7321;
	wire new_net_7985;
	wire new_net_6830;
	wire new_net_237;
	wire new_net_279;
	wire new_net_381;
	wire n_0416_;
	wire n_0710_;
	wire new_net_3560;
	wire n_0920_;
	wire n_1214_;
	wire n_0206_;
	wire new_net_1360;
	wire new_net_4244;
	wire new_net_4530;
	wire new_net_6629;
	wire new_net_6958;
	wire new_net_10097;
	wire new_net_303;
	wire new_net_5634;
	wire new_net_9000;
	wire n_0460_;
	wire new_net_10176;
	wire new_net_2403;
	wire new_net_2701;
	wire new_net_3063;
	wire new_net_3258;
	wire new_net_766;
	wire new_net_1211;
	wire new_net_3975;
	wire new_net_3998;
	wire new_net_2926;
	wire new_net_4199;
	wire new_net_9599;
	wire new_net_10578;
	wire n_1080_;
	wire new_net_10500;
	wire new_net_6610;
	wire new_net_10114;
	wire new_net_7851;
	wire new_net_7558;
	wire new_net_2855;
	wire new_net_1851;
	wire new_net_2642;
	wire new_net_536;
	wire new_net_1737;
	wire n_0417_;
	wire n_0711_;
	wire new_net_914;
	wire n_0921_;
	wire n_1215_;
	wire n_0207_;
	wire new_net_4484;
	wire new_net_4522;
	wire new_net_5076;
	wire new_net_7612;
	wire new_net_9176;
	wire new_net_8471;
	wire new_net_8007;
	wire new_net_9616;
	wire new_net_9552;
	wire new_net_7293;
	wire new_net_9256;
	wire new_net_10409;
	wire new_net_8525;
	wire new_net_1393;
	wire new_net_3626;
	wire new_net_1510;
	wire new_net_801;
	wire new_net_4447;
	wire new_net_4666;
	wire new_net_5393;
	wire new_net_5417;
	wire new_net_5441;
	wire new_net_5671;
	wire new_net_8403;
	wire new_net_8401;
	wire new_net_8696;
	wire new_net_9653;
	wire new_net_9660;
	wire new_net_10566;
	wire new_net_7263;
	wire new_net_3156;
	wire new_net_5716;
	wire new_net_1361;
	wire n_0418_;
	wire n_0922_;
	wire new_net_238;
	wire new_net_2088;
	wire new_net_280;
	wire new_net_3346;
	wire n_1216_;
	wire new_net_382;
	wire n_0712_;
	wire new_net_6857;
	wire new_net_9440;
	wire new_net_6502;
	wire new_net_9882;
	wire new_net_5593;
	wire new_net_2372;
	wire new_net_2677;
	wire new_net_2435;
	wire new_net_2204;
	wire new_net_2477;
	wire new_net_3323;
	wire new_net_2171;
	wire new_net_767;
	wire new_net_1212;
	wire new_net_3020;
	wire new_net_7450;
	wire new_net_9030;
	wire new_net_10213;
	wire new_net_7168;
	wire new_net_6761;
	wire new_net_948;
	wire n_0923_;
	wire new_net_1852;
	wire new_net_537;
	wire n_0209_;
	wire new_net_1998;
	wire new_net_2611;
	wire n_1217_;
	wire new_net_1738;
	wire n_0419_;
	wire new_net_10692;
	wire new_net_3424;
	wire new_net_6167;
	wire new_net_1592;
	wire new_net_2868;
	wire new_net_1511;
	wire new_net_3561;
	wire new_net_652;
	wire new_net_802;
	wire new_net_1394;
	wire new_net_3859;
	wire new_net_5020;
	wire new_net_5079;
	wire new_net_5686;
	wire new_net_8897;
	wire new_net_7530;
	wire new_net_5525;
	wire new_net_10318;
	wire new_net_5523;
	wire new_net_7953;
	wire new_net_10127;
	wire new_net_9499;
	wire new_net_2678;
	wire new_net_239;
	wire new_net_2702;
	wire new_net_3064;
	wire new_net_3259;
	wire new_net_281;
	wire n_0210_;
	wire new_net_383;
	wire n_0924_;
	wire n_1218_;
	wire n_1186_;
	wire new_net_9590;
	wire new_net_5411;
	wire new_net_6032;
	wire new_net_6594;
	wire new_net_9992;
	wire new_net_4825;
	wire new_net_9523;
	wire new_net_2404;
	wire new_net_2513;
	wire new_net_2643;
	wire new_net_4508;
	wire new_net_5959;
	wire new_net_6136;
	wire new_net_7603;
	wire new_net_9382;
	wire new_net_10514;
	wire new_net_10538;
	wire new_net_7896;
	wire new_net_5882;
	wire new_net_5254;
	wire new_net_10508;
	wire new_net_8511;
	wire new_net_10400;
	wire new_net_949;
	wire new_net_1853;
	wire new_net_3627;
	wire n_0211_;
	wire n_0925_;
	wire n_1219_;
	wire n_0421_;
	wire n_0715_;
	wire new_net_4448;
	wire new_net_4667;
	wire new_net_7746;
	wire new_net_9931;
	wire new_net_8566;
	wire new_net_5239;
	wire new_net_10020;
	wire new_net_6188;
	wire new_net_3142;
	wire new_net_8085;
	wire new_net_10530;
	wire new_net_6972;
	wire new_net_8918;
	wire new_net_10528;
	wire new_net_1987;
	wire new_net_3347;
	wire new_net_1362;
	wire new_net_1395;
	wire new_net_1512;
	wire new_net_1593;
	wire new_net_4216;
	wire new_net_5615;
	wire new_net_6360;
	wire new_net_7884;
	wire new_net_10334;
	wire new_net_9431;
	wire new_net_6117;
	wire new_net_5752;
	wire new_net_6267;
	wire new_net_6904;
	wire new_net_10663;
	wire new_net_5579;
	wire new_net_7069;
	wire new_net_8382;
	wire new_net_3021;
	wire new_net_240;
	wire new_net_282;
	wire new_net_768;
	wire new_net_1213;
	wire new_net_3324;
	wire new_net_384;
	wire n_0422_;
	wire n_0716_;
	wire n_0926_;
	wire new_net_5473;
	wire new_net_6315;
	wire new_net_9453;
	wire new_net_9342;
	wire new_net_6747;
	wire new_net_4207;
	wire new_net_10483;
	wire new_net_6553;
	wire new_net_6546;
	wire new_net_2022;
	wire new_net_2373;
	wire new_net_2436;
	wire new_net_2205;
	wire new_net_2478;
	wire new_net_2612;
	wire new_net_538;
	wire new_net_916;
	wire new_net_1739;
	wire new_net_4491;
	wire n_0322_;
	wire new_net_2791;
	wire new_net_7675;
	wire new_net_8960;
	wire new_net_7550;
	wire new_net_4305;
	wire new_net_3625;
	wire new_net_6158;
	wire n_0942_;
	wire new_net_653;
	wire new_net_2869;
	wire n_0927_;
	wire new_net_1854;
	wire n_0213_;
	wire new_net_803;
	wire new_net_3562;
	wire n_0423_;
	wire n_0717_;
	wire new_net_2081;
	wire new_net_6935;
	wire new_net_6489;
	wire new_net_1347;
	wire new_net_7939;
	wire new_net_6660;
	wire new_net_8758;
	wire new_net_1990;
	wire new_net_2679;
	wire new_net_3260;
	wire new_net_2885;
	wire new_net_3065;
	wire new_net_2703;
	wire new_net_1363;
	wire new_net_1513;
	wire new_net_3977;
	wire new_net_4000;
	wire new_net_9301;
	wire new_net_9576;
	wire new_net_5359;
	wire new_net_10371;
	wire new_net_10364;
	wire new_net_9983;
	wire new_net_6682;
	wire new_net_385;
	wire new_net_2644;
	wire new_net_241;
	wire new_net_283;
	wire new_net_769;
	wire n_0214_;
	wire new_net_1214;
	wire n_0928_;
	wire n_1222_;
	wire n_0424_;
	wire new_net_798;
	wire new_net_9048;
	wire new_net_9240;
	wire new_net_8502;
	wire new_net_7732;
	wire new_net_1740;
	wire new_net_2172;
	wire new_net_2405;
	wire new_net_3628;
	wire new_net_539;
	wire new_net_917;
	wire new_net_950;
	wire new_net_4449;
	wire new_net_4668;
	wire new_net_5395;
	wire new_net_5105;
	wire new_net_8024;
	wire new_net_7240;
	wire new_net_8557;
	wire new_net_6241;
	wire new_net_710;
	wire n_1146_;
	wire new_net_8357;
	wire new_net_8612;
	wire new_net_9782;
	wire n_0425_;
	wire n_0719_;
	wire new_net_654;
	wire new_net_2114;
	wire new_net_1594;
	wire new_net_1396;
	wire new_net_2886;
	wire new_net_3236;
	wire n_0215_;
	wire new_net_804;
	wire new_net_9780;
	wire new_net_3188;
	wire new_net_376;
	wire new_net_3715;
	wire new_net_6890;
	wire new_net_9188;
	wire new_net_742;
	wire new_net_4685;
	wire new_net_5288;
	wire new_net_7429;
	wire new_net_6405;
	wire new_net_8739;
	wire new_net_10654;
	wire new_net_9910;
	wire new_net_5027;
	wire new_net_1514;
	wire new_net_3022;
	wire new_net_3325;
	wire new_net_3651;
	wire new_net_3675;
	wire new_net_6265;
	wire new_net_6306;
	wire new_net_7925;
	wire new_net_9138;
	wire new_net_10094;
	wire new_net_10077;
	wire new_net_9333;
	wire new_net_6738;
	wire new_net_8598;
	wire new_net_9205;
	wire new_net_5038;
	wire new_net_6016;
	wire new_net_7206;
	wire new_net_1417;
	wire new_net_7199;
	wire new_net_2613;
	wire new_net_386;
	wire new_net_242;
	wire new_net_284;
	wire n_0216_;
	wire new_net_1215;
	wire n_0426_;
	wire n_0720_;
	wire n_0930_;
	wire n_1224_;
	wire new_net_4920;
	wire new_net_304;
	wire new_net_7537;
	wire new_net_6800;
	wire new_net_5157;
	wire new_net_9903;
	wire new_net_3563;
	wire new_net_2374;
	wire new_net_2870;
	wire new_net_1855;
	wire new_net_2437;
	wire new_net_2206;
	wire new_net_2479;
	wire new_net_540;
	wire new_net_951;
	wire new_net_3861;
	wire new_net_7509;
	wire new_net_8455;
	wire new_net_8633;
	wire n_1082_;
	wire new_net_7019;
	wire new_net_7930;
	wire new_net_6651;
	wire new_net_5658;
	wire new_net_10268;
	wire n_1225_;
	wire new_net_1973;
	wire new_net_1364;
	wire new_net_1595;
	wire new_net_2680;
	wire n_0931_;
	wire new_net_1397;
	wire new_net_2704;
	wire new_net_3066;
	wire new_net_3237;
	wire new_net_9905;
	wire new_net_10200;
	wire new_net_9572;
	wire new_net_5345;
	wire new_net_6578;
	wire new_net_9812;
	wire new_net_1479;
	wire new_net_4160;
	wire new_net_7580;
	wire new_net_2515;
	wire new_net_1966;
	wire new_net_770;
	wire new_net_5961;
	wire new_net_6138;
	wire new_net_7873;
	wire new_net_8200;
	wire new_net_9420;
	wire new_net_10516;
	wire new_net_10540;
	wire new_net_216;
	wire new_net_6724;
	wire n_0323_;
	wire new_net_9226;
	wire new_net_10457;
	wire new_net_9829;
	wire new_net_10455;
	wire new_net_3909;
	wire new_net_7723;
	wire n_0218_;
	wire new_net_1216;
	wire new_net_387;
	wire new_net_1741;
	wire new_net_918;
	wire new_net_243;
	wire new_net_3629;
	wire new_net_285;
	wire new_net_1977;
	wire n_0932_;
	wire new_net_4102;
	wire new_net_866;
	wire new_net_4100;
	wire new_net_7231;
	wire new_net_8427;
	wire new_net_8548;
	wire new_net_9679;
	wire new_net_3546;
	wire new_net_4561;
	wire new_net_6445;
	wire new_net_9677;
	wire new_net_7282;
	wire new_net_3349;
	wire new_net_2887;
	wire new_net_2406;
	wire new_net_1856;
	wire new_net_541;
	wire new_net_655;
	wire new_net_805;
	wire new_net_4218;
	wire new_net_5617;
	wire new_net_6362;
	wire new_net_8118;
	wire new_net_9852;
	wire new_net_9537;
	wire new_net_7831;
	wire new_net_6881;
	wire new_net_8207;
	wire new_net_7420;
	wire new_net_8730;
	wire new_net_7413;
	wire new_net_5450;
	wire new_net_8877;
	wire new_net_9152;
	wire new_net_6297;
	wire new_net_4383;
	wire new_net_7142;
	wire new_net_9710;
	wire new_net_6432;
	wire new_net_4184;
	wire new_net_4906;
	wire new_net_9373;
	wire new_net_7654;
	wire new_net_9638;
	wire new_net_8267;
	wire n_0975_;
	wire n_0471_;
	wire new_net_1905;
	wire new_net_1872;
	wire new_net_968;
	wire new_net_3687;
	wire new_net_4914;
	wire new_net_5455;
	wire new_net_5821;
	wire new_net_5845;
	wire new_net_8723;
	wire new_net_5153;
	wire new_net_7336;
	wire new_net_7500;
	wire new_net_8441;
	wire new_net_6840;
	wire new_net_102;
	wire new_net_3529;
	wire new_net_1971;
	wire new_net_4134;
	wire new_net_5182;
	wire new_net_4853;
	wire new_net_5303;
	wire new_net_5993;
	wire new_net_6017;
	wire new_net_7632;
	wire new_net_10107;
	wire new_net_8841;
	wire new_net_5549;
	wire new_net_10191;
	wire new_net_9278;
	wire new_net_6169;
	wire new_net_10431;
	wire n_0976_;
	wire n_0472_;
	wire new_net_181;
	wire new_net_1118;
	wire new_net_1613;
	wire new_net_5868;
	wire new_net_5892;
	wire new_net_6641;
	wire new_net_6665;
	wire new_net_6924;
	wire new_net_7102;
	wire new_net_7109;
	wire new_net_10588;
	wire new_net_5435;
	wire new_net_6049;
	wire new_net_7571;
	wire new_net_5809;
	wire new_net_1086;
	wire new_net_1233;
	wire new_net_2438;
	wire new_net_2270;
	wire new_net_1758;
	wire new_net_2333;
	wire new_net_3446;
	wire new_net_3828;
	wire new_net_3873;
	wire new_net_3897;
	wire new_net_5906;
	wire new_net_9462;
	wire new_net_9742;
	wire new_net_10476;
	wire new_net_6332;
	wire new_net_3804;
	wire new_net_5090;
	wire new_net_8177;
	wire n_0977_;
	wire n_0473_;
	wire new_net_1873;
	wire new_net_3466;
	wire new_net_822;
	wire new_net_3034;
	wire new_net_492;
	wire new_net_969;
	wire new_net_5164;
	wire new_net_6989;
	wire new_net_7763;
	wire new_net_9955;
	wire new_net_10296;
	wire new_net_4146;
	wire new_net_8590;
	wire new_net_10044;
	wire new_net_9757;
	wire new_net_10042;
	wire new_net_10554;
	wire new_net_8310;
	wire new_net_8942;
	wire new_net_8308;
	wire new_net_103;
	wire new_net_1268;
	wire new_net_3597;
	wire new_net_4463;
	wire new_net_4834;
	wire new_net_6054;
	wire new_net_7484;
	wire new_net_8467;
	wire new_net_8717;
	wire new_net_7822;
	wire new_net_9099;
	wire new_net_9097;
	wire new_net_6141;
	wire new_net_9736;
	wire new_net_6396;
	wire new_net_9970;
	wire new_net_5400;
	wire new_net_5316;
	wire new_net_6283;
	wire new_net_5603;
	wire new_net_7460;
	wire n_0474_;
	wire n_0978_;
	wire new_net_71;
	wire new_net_2992;
	wire new_net_3194;
	wire new_net_182;
	wire new_net_1119;
	wire new_net_4273;
	wire new_net_4855;
	wire new_net_5497;
	wire new_net_7183;
	wire new_net_4935;
	wire new_net_10620;
	wire new_net_6771;
	wire new_net_6402;
	wire new_net_9629;
	wire new_net_3;
	wire new_net_1234;
	wire new_net_1906;
	wire new_net_2187;
	wire new_net_1759;
	wire new_net_3688;
	wire new_net_4915;
	wire new_net_5456;
	wire new_net_5822;
	wire new_net_5846;
	wire new_net_5139;
	wire new_net_7322;
	wire new_net_10642;
	wire n_0475_;
	wire n_0979_;
	wire new_net_493;
	wire new_net_970;
	wire new_net_823;
	wire new_net_3530;
	wire new_net_5183;
	wire new_net_5304;
	wire new_net_5994;
	wire new_net_6018;
	wire new_net_6959;
	wire new_net_8675;
	wire new_net_9001;
	wire new_net_4208;
	wire new_net_10177;
	wire new_net_1269;
	wire new_net_1614;
	wire new_net_2839;
	wire new_net_5869;
	wire new_net_5893;
	wire new_net_6642;
	wire new_net_6666;
	wire new_net_6925;
	wire new_net_6949;
	wire new_net_6973;
	wire new_net_10579;
	wire new_net_10501;
	wire new_net_6611;
	wire n_0798_;
	wire new_net_7852;
	wire new_net_7559;
	wire new_net_6699;
	wire new_net_7361;
	wire new_net_183;
	wire new_net_1120;
	wire n_0980_;
	wire n_0476_;
	wire new_net_3447;
	wire new_net_2034;
	wire new_net_72;
	wire new_net_1087;
	wire new_net_3829;
	wire new_net_3874;
	wire new_net_8472;
	wire new_net_10091;
	wire new_net_9617;
	wire new_net_9615;
	wire new_net_9257;
	wire new_net_10410;
	wire new_net_8526;
	wire new_net_8404;
	wire new_net_8697;
	wire new_net_2439;
	wire new_net_3035;
	wire new_net_1874;
	wire new_net_1907;
	wire new_net_2517;
	wire new_net_2271;
	wire new_net_3467;
	wire new_net_2334;
	wire new_net_3939;
	wire new_net_5165;
	wire new_net_9661;
	wire new_net_7264;
	wire new_net_6260;
	wire new_net_8138;
	wire new_net_6406;
	wire n_0981_;
	wire new_net_3598;
	wire new_net_494;
	wire new_net_971;
	wire new_net_824;
	wire new_net_2035;
	wire new_net_104;
	wire n_0477_;
	wire new_net_3684;
	wire new_net_4671;
	wire new_net_6127;
	wire new_net_6858;
	wire new_net_9441;
	wire new_net_9883;
	wire new_net_5039;
	wire new_net_9964;
	wire new_net_4362;
	wire new_net_9033;
	wire new_net_7451;
	wire new_net_9031;
	wire new_net_1615;
	wire new_net_2993;
	wire new_net_3195;
	wire new_net_4274;
	wire new_net_4856;
	wire new_net_5537;
	wire new_net_5561;
	wire new_net_6376;
	wire new_net_7304;
	wire new_net_7328;
	wire new_net_6507;
	wire new_net_7169;
	wire new_net_8205;
	wire new_net_6762;
	wire new_net_1088;
	wire n_0478_;
	wire n_0982_;
	wire new_net_184;
	wire new_net_1121;
	wire new_net_1760;
	wire new_net_3689;
	wire new_net_4916;
	wire new_net_5457;
	wire new_net_5823;
	wire new_net_7685;
	wire new_net_7313;
	wire new_net_6168;
	wire new_net_1236;
	wire new_net_1875;
	wire new_net_1908;
	wire new_net_2188;
	wire new_net_3531;
	wire new_net_5184;
	wire new_net_5305;
	wire new_net_5995;
	wire new_net_6019;
	wire new_net_6987;
	wire new_net_7531;
	wire new_net_4285;
	wire new_net_5526;
	wire new_net_10319;
	wire new_net_8657;
	wire new_net_8992;
	wire new_net_7954;
	wire new_net_10128;
	wire new_net_2840;
	wire n_0479_;
	wire n_0983_;
	wire new_net_825;
	wire new_net_1270;
	wire new_net_105;
	wire new_net_5124;
	wire new_net_5870;
	wire new_net_5894;
	wire new_net_6643;
	wire new_net_5412;
	wire new_net_6033;
	wire new_net_9591;
	wire new_net_5369;
	wire new_net_9993;
	wire new_net_8375;
	wire new_net_9524;
	wire new_net_4509;
	wire new_net_7604;
	wire new_net_73;
	wire new_net_3448;
	wire new_net_3830;
	wire new_net_3875;
	wire new_net_3899;
	wire new_net_3922;
	wire new_net_4171;
	wire new_net_5127;
	wire new_net_6197;
	wire new_net_6448;
	wire new_net_5255;
	wire new_net_7897;
	wire new_net_10509;
	wire new_net_8512;
	wire new_net_10401;
	wire new_net_10275;
	wire new_net_7747;
	wire new_net_9932;
	wire new_net_1761;
	wire n_0984_;
	wire n_0480_;
	wire new_net_185;
	wire new_net_3036;
	wire new_net_3468;
	wire new_net_4877;
	wire new_net_5166;
	wire new_net_6991;
	wire new_net_7158;
	wire new_net_8567;
	wire new_net_10294;
	wire new_net_4123;
	wire new_net_6251;
	wire new_net_10021;
	wire new_net_10670;
	wire new_net_8088;
	wire new_net_10531;
	wire new_net_8919;
	wire new_net_10335;
	wire new_net_495;
	wire new_net_972;
	wire new_net_1876;
	wire new_net_2335;
	wire new_net_3599;
	wire new_net_2440;
	wire new_net_2272;
	wire new_net_6056;
	wire new_net_6118;
	wire new_net_7486;
	wire new_net_6905;
	wire new_net_4945;
	wire new_net_5580;
	wire new_net_7070;
	wire new_net_8383;
	wire new_net_5474;
	wire new_net_8681;
	wire new_net_7299;
	wire new_net_106;
	wire n_0481_;
	wire n_0985_;
	wire new_net_3196;
	wire new_net_1271;
	wire new_net_2994;
	wire new_net_1616;
	wire new_net_4135;
	wire new_net_4857;
	wire new_net_5125;
	wire new_net_6316;
	wire new_net_4998;
	wire new_net_9454;
	wire new_net_9343;
	wire new_net_6748;
	wire new_net_9258;
	wire new_net_6554;
	wire new_net_10484;
	wire new_net_6547;
	wire new_net_74;
	wire new_net_1089;
	wire new_net_1122;
	wire new_net_3690;
	wire new_net_4275;
	wire new_net_4917;
	wire new_net_5458;
	wire new_net_5824;
	wire new_net_5848;
	wire new_net_6743;
	wire new_net_8963;
	wire new_net_7676;
	wire new_net_8961;
	wire new_net_5017;
	wire new_net_7551;
	wire new_net_4342;
	wire new_net_6810;
	wire new_net_4306;
	wire new_net_3532;
	wire n_0482_;
	wire n_0986_;
	wire new_net_186;
	wire new_net_1909;
	wire new_net_1237;
	wire new_net_5185;
	wire new_net_5306;
	wire new_net_5996;
	wire new_net_6020;
	wire new_net_6490;
	wire new_net_4271;
	wire new_net_7940;
	wire new_net_9841;
	wire new_net_6661;
	wire new_net_5668;
	wire new_net_8233;
	wire new_net_8759;
	wire new_net_496;
	wire new_net_826;
	wire new_net_973;
	wire new_net_2189;
	wire new_net_5871;
	wire new_net_5895;
	wire new_net_6644;
	wire new_net_6668;
	wire new_net_6927;
	wire new_net_6951;
	wire new_net_9302;
	wire new_net_9577;
	wire new_net_5360;
	wire new_net_10372;
	wire new_net_10365;
	wire new_net_9984;
	wire new_net_6683;
	wire new_net_5054;
	wire new_net_7590;
	wire n_0483_;
	wire n_0987_;
	wire new_net_107;
	wire new_net_1617;
	wire new_net_3278;
	wire new_net_3449;
	wire new_net_3831;
	wire new_net_3876;
	wire new_net_3900;
	wire new_net_3923;
	wire new_net_5833;
	wire new_net_9049;
	wire new_net_9241;
	wire new_net_7733;
	wire new_net_8025;
	wire new_net_1090;
	wire new_net_1762;
	wire new_net_3037;
	wire new_net_2061;
	wire new_net_3469;
	wire new_net_2519;
	wire new_net_5167;
	wire new_net_6992;
	wire new_net_7159;
	wire new_net_7182;
	wire new_net_7241;
	wire new_net_8558;
	wire new_net_3976;
	wire new_net_8358;
	wire new_net_8613;
	wire new_net_9781;
	wire n_0484_;
	wire n_0988_;
	wire new_net_187;
	wire new_net_3600;
	wire new_net_1877;
	wire new_net_1910;
	wire new_net_1238;
	wire new_net_4464;
	wire new_net_4620;
	wire new_net_6057;
	wire new_net_6654;
	wire new_net_8332;
	wire new_net_8843;
	wire new_net_6891;
	wire new_net_4936;
	wire new_net_5289;
	wire new_net_7430;
	wire new_net_8740;
	wire new_net_8136;
	wire new_net_10655;
	wire new_net_9911;
	wire new_net_5465;
	wire new_net_2273;
	wire new_net_827;
	wire new_net_1272;
	wire new_net_2995;
	wire new_net_2336;
	wire new_net_3197;
	wire new_net_2441;
	wire new_net_4858;
	wire new_net_5126;
	wire new_net_5539;
	wire new_net_4986;
	wire new_net_10078;
	wire new_net_9334;
	wire new_net_6739;
	wire new_net_4194;
	wire new_net_8599;
	wire new_net_9206;
	wire new_net_7207;
	wire new_net_5935;
	wire new_net_7200;
	wire n_0989_;
	wire n_0485_;
	wire new_net_75;
	wire new_net_2841;
	wire new_net_1618;
	wire new_net_3691;
	wire new_net_4276;
	wire new_net_4839;
	wire new_net_4918;
	wire new_net_5108;
	wire new_net_4292;
	wire new_net_4209;
	wire new_net_7341;
	wire new_net_9904;
	wire new_net_7510;
	wire new_net_4;
	wire new_net_1091;
	wire new_net_1124;
	wire new_net_1763;
	wire new_net_3533;
	wire new_net_4003;
	wire new_net_4136;
	wire new_net_5186;
	wire new_net_5307;
	wire new_net_5997;
	wire new_net_8456;
	wire new_net_8634;
	wire new_net_7020;
	wire new_net_7931;
	wire new_net_6652;
	wire new_net_5659;
	wire new_net_10269;
	wire new_net_10201;
	wire n_0990_;
	wire new_net_974;
	wire n_0486_;
	wire new_net_188;
	wire new_net_497;
	wire new_net_4465;
	wire new_net_4836;
	wire new_net_5872;
	wire new_net_5896;
	wire new_net_6645;
	wire new_net_8824;
	wire new_net_5346;
	wire new_net_6579;
	wire new_net_9813;
	wire new_net_9069;
	wire new_net_6064;
	wire new_net_6674;
	wire new_net_7581;
	wire new_net_7874;
	wire new_net_3273;
	wire new_net_3450;
	wire new_net_108;
	wire new_net_828;
	wire new_net_1273;
	wire new_net_3832;
	wire new_net_3877;
	wire new_net_3901;
	wire new_net_3924;
	wire new_net_4173;
	wire new_net_6725;
	wire new_net_9421;
	wire new_net_10223;
	wire new_net_9227;
	wire new_net_10458;
	wire new_net_4779;
	wire new_net_7724;
	wire new_net_8672;
	wire new_net_2190;
	wire n_0487_;
	wire n_0991_;
	wire new_net_76;
	wire new_net_3038;
	wire new_net_3470;
	wire new_net_3814;
	wire new_net_4878;
	wire new_net_6993;
	wire new_net_7160;
	wire new_net_7232;
	wire new_net_8549;
	wire new_net_3685;
	wire new_net_4990;
	wire new_net_6228;
	wire new_net_8428;
	wire new_net_4562;
	wire new_net_8063;
	wire new_net_7283;
	wire new_net_8793;
	wire new_net_4606;
	wire new_net_6789;
	wire new_net_8119;
	wire new_net_1911;
	wire new_net_1092;
	wire new_net_1125;
	wire new_net_1239;
	wire new_net_1764;
	wire new_net_3601;
	wire new_net_6058;
	wire new_net_7488;
	wire new_net_8721;
	wire new_net_9492;
	wire new_net_9853;
	wire new_net_9538;
	wire new_net_7832;
	wire new_net_6882;
	wire new_net_7421;
	wire new_net_8731;
	wire new_net_7414;
	wire new_net_5451;
	wire new_net_8878;
	wire new_net_9153;
	wire new_net_3280;
	wire n_0488_;
	wire new_net_2996;
	wire new_net_3198;
	wire new_net_189;
	wire new_net_498;
	wire new_net_975;
	wire n_0992_;
	wire new_net_1879;
	wire new_net_3955;
	wire new_net_4713;
	wire new_net_5613;
	wire new_net_9711;
	wire new_net_9320;
	wire new_net_3953;
	wire new_net_6433;
	wire new_net_8339;
	wire new_net_10115;
	wire new_net_6531;
	wire new_net_9376;
	wire new_net_10630;
	wire new_net_9374;
	wire new_net_9639;
	wire new_net_7655;
	wire new_net_2442;
	wire new_net_109;
	wire new_net_1619;
	wire new_net_2274;
	wire new_net_2093;
	wire new_net_2337;
	wire new_net_3213;
	wire new_net_3692;
	wire new_net_4879;
	wire new_net_4919;
	wire new_net_7653;
	wire new_net_8578;
	wire new_net_4282;
	wire new_net_7337;
	wire new_net_4083;
	wire new_net_7501;
	wire n_0993_;
	wire n_0489_;
	wire new_net_3534;
	wire new_net_4137;
	wire new_net_5187;
	wire new_net_5308;
	wire new_net_5998;
	wire new_net_6022;
	wire new_net_6841;
	wire new_net_7636;
	wire new_net_8442;
	wire n_0327_;
	wire new_net_9391;
	wire new_net_4854;
	wire new_net_7011;
	wire new_net_10108;
	wire new_net_5650;
	wire new_net_8842;
	wire new_net_5550;
	wire new_net_9281;
	wire new_net_10192;
	wire new_net_8250;
	wire new_net_1240;
	wire new_net_1912;
	wire new_net_2842;
	wire new_net_4466;
	wire new_net_5873;
	wire new_net_5897;
	wire new_net_6391;
	wire new_net_6646;
	wire new_net_6670;
	wire new_net_6929;
	wire new_net_10432;
	wire new_net_5337;
	wire new_net_9804;
	wire new_net_10349;
	wire new_net_10589;
	wire new_net_5436;
	wire new_net_8231;
	wire new_net_7572;
	wire new_net_5810;
	wire new_net_1880;
	wire n_0994_;
	wire n_0490_;
	wire new_net_829;
	wire new_net_1274;
	wire new_net_190;
	wire new_net_499;
	wire new_net_976;
	wire new_net_3451;
	wire new_net_3833;
	wire new_net_3843;
	wire new_net_5907;
	wire new_net_9463;
	wire new_net_9743;
	wire new_net_7633;
	wire new_net_6333;
	wire new_net_3471;
	wire new_net_77;
	wire new_net_1620;
	wire new_net_2521;
	wire new_net_3039;
	wire new_net_6994;
	wire new_net_7184;
	wire new_net_3672;
	wire new_net_7208;
	wire new_net_7469;
	wire new_net_7766;
	wire new_net_8178;
	wire new_net_8414;
	wire new_net_8535;
	wire new_net_9956;
	wire new_net_10299;
	wire new_net_7764;
	wire new_net_10297;
	wire new_net_8591;
	wire new_net_10045;
	wire new_net_10043;
	wire new_net_10555;
	wire n_0491_;
	wire n_0995_;
	wire new_net_2011;
	wire new_net_1765;
	wire new_net_1093;
	wire new_net_3602;
	wire new_net_1126;
	wire new_net_6059;
	wire new_net_6392;
	wire new_net_7489;
	wire new_net_8941;
	wire new_net_9100;
	wire new_net_7823;
	wire new_net_6142;
	wire new_net_9098;
	wire new_net_3749;
	wire new_net_4969;
	wire new_net_6284;
	wire new_net_10065;
	wire new_net_2040;
	wire new_net_3279;
	wire new_net_1241;
	wire new_net_1913;
	wire new_net_3199;
	wire new_net_4838;
	wire new_net_4860;
	wire new_net_4967;
	wire new_net_5541;
	wire new_net_5604;
	wire new_net_7461;
	wire new_net_5498;
	wire new_net_6517;
	wire new_net_9122;
	wire new_net_10381;
	wire new_net_10621;
	wire new_net_6772;
	wire new_net_500;
	wire new_net_977;
	wire n_0492_;
	wire n_0996_;
	wire new_net_5;
	wire new_net_830;
	wire new_net_1275;
	wire new_net_191;
	wire new_net_110;
	wire new_net_3693;
	wire new_net_7323;
	wire new_net_10643;
	wire new_net_2443;
	wire new_net_78;
	wire new_net_2191;
	wire new_net_3535;
	wire new_net_2275;
	wire new_net_2338;
	wire new_net_5168;
	wire new_net_5188;
	wire new_net_5309;
	wire new_net_5999;
	wire new_net_6631;
	wire new_net_4532;
	wire new_net_9002;
	wire new_net_10178;
	wire new_net_9512;
	wire new_net_1127;
	wire new_net_2057;
	wire n_0997_;
	wire n_0493_;
	wire new_net_1094;
	wire new_net_2843;
	wire new_net_5874;
	wire new_net_5898;
	wire new_net_6647;
	wire new_net_6671;
	wire new_net_10580;
	wire new_net_10502;
	wire new_net_6612;
	wire new_net_7853;
	wire new_net_10664;
	wire new_net_5801;
	wire new_net_3452;
	wire new_net_1242;
	wire new_net_1881;
	wire new_net_1914;
	wire new_net_3834;
	wire new_net_3879;
	wire new_net_3903;
	wire new_net_3926;
	wire new_net_4277;
	wire new_net_6201;
	wire new_net_7614;
	wire new_net_4524;
	wire new_net_8268;
	wire new_net_8473;
	wire new_net_7995;
	wire new_net_7295;
	wire new_net_10411;
	wire new_net_192;
	wire new_net_3040;
	wire new_net_1621;
	wire n_0998_;
	wire n_0494_;
	wire new_net_3472;
	wire new_net_1276;
	wire new_net_111;
	wire new_net_4278;
	wire new_net_6995;
	wire new_net_8405;
	wire new_net_8698;
	wire new_net_6375;
	wire new_net_9662;
	wire n_0328_;
	wire new_net_7265;
	wire new_net_744;
	wire new_net_10541;
	wire new_net_8378;
	wire new_net_3603;
	wire new_net_5128;
	wire new_net_5169;
	wire new_net_5718;
	wire new_net_6060;
	wire new_net_7490;
	wire new_net_8947;
	wire new_net_6861;
	wire new_net_9494;
	wire new_net_4987;
	wire new_net_6859;
	wire new_net_9442;
	wire new_net_10665;
	wire new_net_9884;
	wire new_net_8862;
	wire new_net_3740;
	wire new_net_4363;
	wire new_net_1095;
	wire new_net_3200;
	wire n_0495_;
	wire n_0999_;
	wire new_net_1767;
	wire new_net_4861;
	wire new_net_5542;
	wire new_net_6381;
	wire new_net_7309;
	wire new_net_7333;
	wire new_net_8686;
	wire new_net_9032;
	wire new_net_10215;
	wire new_net_6508;
	wire new_net_7170;
	wire new_net_8206;
	wire new_net_6763;
	wire new_net_3764;
	wire new_net_501;
	wire new_net_831;
	wire new_net_978;
	wire new_net_1882;
	wire new_net_1243;
	wire new_net_3694;
	wire new_net_4921;
	wire new_net_5462;
	wire new_net_5828;
	wire new_net_5852;
	wire new_net_7314;
	wire new_net_6171;
	wire new_net_8752;
	wire new_net_193;
	wire n_0496_;
	wire n_1000_;
	wire new_net_1622;
	wire new_net_79;
	wire new_net_3536;
	wire new_net_4174;
	wire new_net_5189;
	wire new_net_5310;
	wire new_net_5690;
	wire new_net_6990;
	wire new_net_8899;
	wire new_net_5688;
	wire new_net_4027;
	wire new_net_4025;
	wire new_net_5527;
	wire new_net_10320;
	wire new_net_8658;
	wire new_net_8993;
	wire new_net_7955;
	wire new_net_9783;
	wire new_net_10129;
	wire new_net_2339;
	wire new_net_1128;
	wire new_net_2444;
	wire new_net_2192;
	wire new_net_2276;
	wire new_net_5875;
	wire new_net_5899;
	wire new_net_6648;
	wire new_net_6672;
	wire new_net_6931;
	wire new_net_9592;
	wire new_net_5370;
	wire new_net_6480;
	wire new_net_9994;
	wire new_net_1768;
	wire n_1001_;
	wire n_0497_;
	wire new_net_3453;
	wire new_net_1915;
	wire new_net_6;
	wire new_net_3835;
	wire new_net_3880;
	wire new_net_3904;
	wire new_net_3927;
	wire new_net_4472;
	wire new_net_4510;
	wire new_net_5064;
	wire new_net_7605;
	wire new_net_7898;
	wire new_net_5884;
	wire new_net_8661;
	wire new_net_8513;
	wire new_net_112;
	wire new_net_502;
	wire new_net_832;
	wire new_net_979;
	wire new_net_1277;
	wire new_net_1883;
	wire new_net_3473;
	wire new_net_2523;
	wire new_net_3041;
	wire new_net_6996;
	wire new_net_7748;
	wire new_net_9933;
	wire new_net_8208;
	wire new_net_8568;
	wire new_net_4039;
	wire new_net_6252;
	wire new_net_10022;
	wire new_net_8089;
	wire new_net_6190;
	wire new_net_8087;
	wire new_net_10532;
	wire new_net_6974;
	wire new_net_8920;
	wire new_net_194;
	wire new_net_3604;
	wire n_1002_;
	wire n_0498_;
	wire new_net_1623;
	wire new_net_80;
	wire new_net_5129;
	wire new_net_5170;
	wire new_net_6061;
	wire new_net_6790;
	wire new_net_10336;
	wire new_net_6119;
	wire new_net_5754;
	wire new_net_4946;
	wire new_net_6906;
	wire new_net_4354;
	wire new_net_5581;
	wire new_net_3201;
	wire new_net_1096;
	wire new_net_1129;
	wire new_net_4862;
	wire new_net_5543;
	wire new_net_6382;
	wire new_net_7286;
	wire new_net_5475;
	wire new_net_7310;
	wire new_net_7334;
	wire new_net_8682;
	wire new_net_6317;
	wire new_net_9344;
	wire new_net_9897;
	wire new_net_6555;
	wire new_net_2997;
	wire n_0499_;
	wire n_1003_;
	wire new_net_3214;
	wire new_net_1244;
	wire new_net_3695;
	wire new_net_4175;
	wire new_net_4922;
	wire new_net_5110;
	wire new_net_5463;
	wire new_net_8964;
	wire new_net_7677;
	wire new_net_8962;
	wire new_net_9282;
	wire new_net_4307;
	wire new_net_3537;
	wire new_net_113;
	wire new_net_1278;
	wire new_net_1884;
	wire new_net_1980;
	wire new_net_5190;
	wire new_net_5311;
	wire new_net_6001;
	wire new_net_6025;
	wire new_net_7662;
	wire new_net_9680;
	wire new_net_6491;
	wire new_net_9062;
	wire new_net_7941;
	wire new_net_9842;
	wire new_net_6662;
	wire new_net_5669;
	wire n_0500_;
	wire n_1004_;
	wire new_net_195;
	wire new_net_4467;
	wire new_net_5876;
	wire new_net_5900;
	wire new_net_6393;
	wire new_net_6649;
	wire new_net_6932;
	wire new_net_6956;
	wire new_net_9305;
	wire new_net_5739;
	wire new_net_9578;
	wire new_net_9303;
	wire new_net_10098;
	wire new_net_5361;
	wire new_net_10373;
	wire new_net_7538;
	wire new_net_4680;
	wire new_net_10366;
	wire new_net_9985;
	wire new_net_2277;
	wire new_net_1769;
	wire new_net_2340;
	wire new_net_1097;
	wire new_net_3454;
	wire new_net_2445;
	wire new_net_2193;
	wire new_net_3836;
	wire new_net_3881;
	wire new_net_3905;
	wire new_net_9490;
	wire new_net_5834;
	wire new_net_9050;
	wire new_net_9600;
	wire new_net_10468;
	wire new_net_9242;
	wire n_0803_;
	wire n_0501_;
	wire new_net_3042;
	wire new_net_503;
	wire new_net_980;
	wire n_1005_;
	wire new_net_3474;
	wire new_net_1917;
	wire new_net_833;
	wire new_net_1245;
	wire new_net_6997;
	wire new_net_7734;
	wire new_net_8026;
	wire new_net_8559;
	wire new_net_3979;
	wire new_net_6458;
	wire new_net_8724;
	wire new_net_9259;
	wire new_net_8359;
	wire new_net_5702;
	wire new_net_8614;
	wire new_net_1279;
	wire new_net_2012;
	wire new_net_1624;
	wire new_net_4138;
	wire new_net_5171;
	wire new_net_6062;
	wire new_net_6394;
	wire new_net_6791;
	wire new_net_7492;
	wire new_net_7638;
	wire new_net_7793;
	wire new_net_4621;
	wire new_net_5196;
	wire new_net_7962;
	wire new_net_9863;
	wire new_net_8333;
	wire new_net_8844;
	wire new_net_6892;
	wire new_net_4937;
	wire new_net_5290;
	wire new_net_7431;
	wire new_net_8137;
	wire new_net_6895;
	wire new_net_8741;
	wire new_net_10656;
	wire new_net_3215;
	wire n_0502_;
	wire n_1006_;
	wire new_net_1130;
	wire new_net_3202;
	wire new_net_196;
	wire new_net_4279;
	wire new_net_4863;
	wire new_net_5544;
	wire new_net_6383;
	wire new_net_6308;
	wire new_net_5620;
	wire new_net_10079;
	wire new_net_9335;
	wire new_net_4195;
	wire new_net_9207;
	wire new_net_1770;
	wire new_net_3696;
	wire new_net_4923;
	wire new_net_5464;
	wire new_net_5830;
	wire new_net_5854;
	wire new_net_6749;
	wire new_net_6773;
	wire new_net_7201;
	wire new_net_7947;
	wire new_net_4293;
	wire new_net_6802;
	wire new_net_7342;
	wire new_net_834;
	wire new_net_1246;
	wire new_net_3538;
	wire new_net_114;
	wire n_1007_;
	wire n_0503_;
	wire new_net_504;
	wire new_net_981;
	wire new_net_1885;
	wire new_net_1918;
	wire new_net_7511;
	wire new_net_4004;
	wire new_net_8457;
	wire new_net_8635;
	wire new_net_7021;
	wire new_net_7932;
	wire new_net_5660;
	wire new_net_1625;
	wire new_net_4139;
	wire new_net_5877;
	wire new_net_5901;
	wire new_net_6650;
	wire new_net_6933;
	wire new_net_6957;
	wire new_net_8319;
	wire new_net_8476;
	wire new_net_8516;
	wire new_net_10202;
	wire new_net_8825;
	wire new_net_6580;
	wire new_net_9070;
	wire new_net_9971;
	wire new_net_4162;
	wire new_net_6675;
	wire n_0504_;
	wire n_1008_;
	wire new_net_1098;
	wire new_net_197;
	wire new_net_1131;
	wire new_net_841;
	wire new_net_3837;
	wire new_net_3882;
	wire new_net_3906;
	wire new_net_3929;
	wire new_net_6726;
	wire new_net_10224;
	wire new_net_9228;
	wire new_net_10459;
	wire new_net_2194;
	wire new_net_2525;
	wire new_net_2278;
	wire new_net_2341;
	wire new_net_3043;
	wire new_net_2446;
	wire new_net_4469;
	wire new_net_6343;
	wire new_net_6998;
	wire new_net_7164;
	wire new_net_7725;
	wire new_net_4104;
	wire new_net_8188;
	wire new_net_8429;
	wire new_net_7284;
	wire new_net_8600;
	wire new_net_1247;
	wire new_net_1280;
	wire n_0505_;
	wire n_1009_;
	wire new_net_115;
	wire new_net_982;
	wire new_net_1886;
	wire new_net_3649;
	wire new_net_5172;
	wire new_net_6063;
	wire new_net_8120;
	wire new_net_8794;
	wire new_net_9539;
	wire new_net_7833;
	wire new_net_6883;
	wire new_net_7422;
	wire new_net_8732;
	wire new_net_7415;
	wire new_net_2844;
	wire new_net_3203;
	wire new_net_4280;
	wire new_net_4840;
	wire new_net_4864;
	wire new_net_4881;
	wire new_net_5545;
	wire new_net_6384;
	wire new_net_7288;
	wire new_net_7312;
	wire new_net_8879;
	wire new_net_6299;
	wire new_net_9154;
	wire new_net_5614;
	wire new_net_9321;
	wire new_net_3954;
	wire new_net_6434;
	wire new_net_8340;
	wire new_net_6532;
	wire new_net_7560;
	wire new_net_10631;
	wire n_1010_;
	wire n_0506_;
	wire new_net_1771;
	wire new_net_1099;
	wire new_net_198;
	wire new_net_170;
	wire new_net_3697;
	wire new_net_4468;
	wire new_net_4908;
	wire new_net_4924;
	wire new_net_7656;
	wire new_net_9375;
	wire new_net_3788;
	wire new_net_9640;
	wire new_net_7161;
	wire new_net_9540;
	wire new_net_7338;
	wire new_net_1919;
	wire new_net_505;
	wire new_net_835;
	wire new_net_3539;
	wire new_net_5192;
	wire new_net_5313;
	wire new_net_6003;
	wire new_net_6027;
	wire new_net_6673;
	wire new_net_7640;
	wire new_net_8443;
	wire new_net_6842;
	wire new_net_9392;
	wire new_net_8621;
	wire new_net_5551;
	wire new_net_9012;
	wire new_net_1887;
	wire n_1011_;
	wire n_0507_;
	wire new_net_83;
	wire new_net_1281;
	wire new_net_116;
	wire new_net_2845;
	wire new_net_3216;
	wire new_net_983;
	wire new_net_1626;
	wire new_net_9280;
	wire new_net_10193;
	wire new_net_10433;
	wire new_net_10350;
	wire new_net_10590;
	wire new_net_6051;
	wire new_net_8232;
	wire new_net_1132;
	wire new_net_3838;
	wire new_net_3883;
	wire new_net_3907;
	wire new_net_3930;
	wire new_net_4177;
	wire new_net_5113;
	wire new_net_6456;
	wire new_net_5811;
	wire new_net_8459;
	wire new_net_7374;
	wire new_net_9034;
	wire new_net_9466;
	wire new_net_5908;
	wire new_net_9464;
	wire new_net_9744;
	wire new_net_9652;
	wire new_net_2119;
	wire n_0508_;
	wire n_1012_;
	wire new_net_1772;
	wire new_net_199;
	wire new_net_3044;
	wire new_net_6334;
	wire new_net_6999;
	wire new_net_7165;
	wire new_net_7189;
	wire new_net_8179;
	wire new_net_8536;
	wire new_net_3673;
	wire new_net_7767;
	wire new_net_8415;
	wire new_net_10300;
	wire new_net_9957;
	wire new_net_7765;
	wire new_net_10298;
	wire new_net_4148;
	wire new_net_8592;
	wire new_net_10046;
	wire new_net_3281;
	wire new_net_2447;
	wire new_net_2195;
	wire new_net_506;
	wire new_net_836;
	wire new_net_1248;
	wire new_net_1920;
	wire new_net_2279;
	wire new_net_2342;
	wire new_net_5173;
	wire new_net_10556;
	wire new_net_8312;
	wire new_net_9101;
	wire new_net_7824;
	wire new_net_6143;
	wire new_net_2092;
	wire new_net_1627;
	wire n_1013_;
	wire new_net_1888;
	wire n_0509_;
	wire new_net_84;
	wire new_net_1978;
	wire new_net_3750;
	wire new_net_4281;
	wire new_net_4841;
	wire new_net_4865;
	wire new_net_4970;
	wire new_net_5318;
	wire new_net_6285;
	wire new_net_4968;
	wire new_net_5605;
	wire new_net_7462;
	wire new_net_5499;
	wire new_net_5123;
	wire new_net_6518;
	wire new_net_9123;
	wire new_net_10382;
	wire new_net_7533;
	wire new_net_7185;
	wire new_net_10622;
	wire new_net_1100;
	wire new_net_1133;
	wire new_net_3698;
	wire new_net_4925;
	wire new_net_5466;
	wire new_net_5832;
	wire new_net_6175;
	wire new_net_6751;
	wire new_net_6775;
	wire new_net_6975;
	wire new_net_10510;
	wire new_net_5141;
	wire new_net_7324;
	wire new_net_200;
	wire n_1014_;
	wire n_0510_;
	wire new_net_3540;
	wire new_net_1773;
	wire new_net_5193;
	wire new_net_5314;
	wire new_net_6004;
	wire new_net_6028;
	wire new_net_7641;
	wire new_net_10644;
	wire new_net_3217;
	wire new_net_117;
	wire new_net_507;
	wire new_net_984;
	wire new_net_1249;
	wire new_net_1282;
	wire new_net_2846;
	wire new_net_4141;
	wire new_net_4883;
	wire new_net_5879;
	wire new_net_9513;
	wire new_net_10179;
	wire new_net_10581;
	wire new_net_6613;
	wire new_net_7854;
	wire new_net_1628;
	wire n_1015_;
	wire n_0511_;
	wire new_net_2998;
	wire new_net_3839;
	wire new_net_3884;
	wire new_net_3908;
	wire new_net_3931;
	wire new_net_4178;
	wire new_net_5114;
	wire new_net_5802;
	wire new_net_8387;
	wire new_net_8269;
	wire new_net_8474;
	wire new_net_7996;
	wire new_net_3045;
	wire new_net_1101;
	wire new_net_2527;
	wire new_net_6976;
	wire new_net_7000;
	wire new_net_7166;
	wire new_net_7190;
	wire new_net_7214;
	wire new_net_7296;
	wire new_net_8165;
	wire new_net_10066;
	wire new_net_8406;
	wire new_net_3941;
	wire new_net_9663;
	wire new_net_7266;
	wire new_net_9830;
	wire new_net_3716;
	wire new_net_6262;
	wire new_net_8778;
	wire new_net_201;
	wire n_0512_;
	wire n_1016_;
	wire new_net_1921;
	wire new_net_837;
	wire new_net_2127;
	wire new_net_1774;
	wire new_net_5174;
	wire new_net_5726;
	wire new_net_6065;
	wire new_net_10542;
	wire new_net_9439;
	wire new_net_6862;
	wire new_net_4988;
	wire new_net_6860;
	wire new_net_9443;
	wire new_net_6129;
	wire new_net_8863;
	wire new_net_9885;
	wire new_net_2343;
	wire new_net_1889;
	wire new_net_85;
	wire new_net_118;
	wire new_net_508;
	wire new_net_985;
	wire new_net_1250;
	wire new_net_2196;
	wire new_net_2448;
	wire new_net_1283;
	wire new_net_4364;
	wire new_net_8760;
	wire new_net_6509;
	wire new_net_7171;
	wire new_net_7634;
	wire new_net_5962;
	wire new_net_5504;
	wire new_net_7687;
	wire new_net_9835;
	wire new_net_6172;
	wire new_net_8753;
	wire new_net_6170;
	wire new_net_3507;
	wire n_0765_;
	wire new_net_2947;
	wire n_0555_;
	wire new_net_473;
	wire n_0051_;
	wire n_0261_;
	wire n_1059_;
	wire new_net_557;
	wire n_1269_;
	wire new_net_5689;
	wire new_net_8900;
	wire new_net_4028;
	wire new_net_9690;
	wire new_net_5528;
	wire new_net_10321;
	wire new_net_8659;
	wire new_net_8994;
	wire new_net_7956;
	wire new_net_9784;
	wire new_net_10130;
	wire new_net_2614;
	wire new_net_738;
	wire new_net_1645;
	wire new_net_4092;
	wire new_net_5327;
	wire new_net_7678;
	wire new_net_8006;
	wire new_net_8030;
	wire new_net_10567;
	wire new_net_9593;
	wire new_net_5414;
	wire new_net_6035;
	wire new_net_5371;
	wire new_net_8604;
	wire new_net_4687;
	wire new_net_9995;
	wire new_net_4828;
	wire new_net_9912;
	wire n_1270_;
	wire n_0766_;
	wire new_net_139;
	wire new_net_706;
	wire n_0052_;
	wire n_0262_;
	wire n_0556_;
	wire n_1060_;
	wire new_net_4113;
	wire new_net_5259;
	wire new_net_5885;
	wire new_net_5257;
	wire new_net_2152;
	wire new_net_8514;
	wire new_net_10403;
	wire new_net_3650;
	wire new_net_10277;
	wire new_net_1791;
	wire new_net_3575;
	wire new_net_2135;
	wire new_net_2681;
	wire new_net_2705;
	wire new_net_2727;
	wire new_net_2774;
	wire new_net_2798;
	wire new_net_4525;
	wire new_net_5350;
	wire new_net_7749;
	wire new_net_9934;
	wire new_net_8209;
	wire new_net_8569;
	wire new_net_10023;
	wire new_net_8090;
	wire new_net_6191;
	wire new_net_10533;
	wire new_net_8921;
	wire n_1271_;
	wire new_net_2821;
	wire n_0767_;
	wire new_net_2017;
	wire n_0557_;
	wire new_net_474;
	wire n_0053_;
	wire n_0263_;
	wire new_net_1002;
	wire n_1061_;
	wire new_net_10337;
	wire new_net_6120;
	wire new_net_5755;
	wire new_net_6907;
	wire new_net_4947;
	wire n_0536_;
	wire new_net_1532;
	wire new_net_406;
	wire new_net_739;
	wire new_net_1415;
	wire new_net_4315;
	wire new_net_4339;
	wire new_net_5476;
	wire new_net_6078;
	wire new_net_6318;
	wire new_net_6807;
	wire new_net_8683;
	wire new_net_9814;
	wire new_net_7162;
	wire new_net_9345;
	wire new_net_6750;
	wire new_net_4494;
	wire new_net_6556;
	wire new_net_6549;
	wire new_net_854;
	wire new_net_2968;
	wire new_net_3152;
	wire n_1272_;
	wire new_net_140;
	wire n_0558_;
	wire new_net_707;
	wire n_0054_;
	wire n_0264_;
	wire n_0768_;
	wire new_net_8965;
	wire new_net_5019;
	wire new_net_7472;
	wire new_net_9402;
	wire new_net_6812;
	wire new_net_4308;
	wire new_net_2302;
	wire new_net_1792;
	wire new_net_2159;
	wire new_net_2407;
	wire new_net_2239;
	wire new_net_3508;
	wire new_net_4151;
	wire new_net_5480;
	wire new_net_5914;
	wire new_net_7963;
	wire new_net_9681;
	wire new_net_6492;
	wire new_net_9063;
	wire new_net_8645;
	wire new_net_7942;
	wire new_net_9843;
	wire new_net_4795;
	wire new_net_6663;
	wire new_net_4446;
	wire new_net_5670;
	wire n_1273_;
	wire n_0769_;
	wire n_0559_;
	wire new_net_475;
	wire n_0265_;
	wire n_0055_;
	wire new_net_2108;
	wire new_net_2176;
	wire new_net_1003;
	wire new_net_1646;
	wire new_net_9304;
	wire new_net_9579;
	wire new_net_10099;
	wire new_net_10374;
	wire new_net_7539;
	wire new_net_10367;
	wire new_net_4819;
	wire new_net_6685;
	wire new_net_5056;
	wire new_net_7592;
	wire new_net_1533;
	wire new_net_407;
	wire new_net_740;
	wire new_net_1416;
	wire new_net_4114;
	wire new_net_5691;
	wire new_net_5747;
	wire new_net_6399;
	wire new_net_5835;
	wire new_net_8492;
	wire new_net_8705;
	wire new_net_9051;
	wire new_net_9601;
	wire n_1092_;
	wire new_net_10469;
	wire new_net_9243;
	wire new_net_8852;
	wire new_net_10116;
	wire new_net_3920;
	wire new_net_7735;
	wire new_net_8385;
	wire new_net_3431;
	wire new_net_855;
	wire new_net_1976;
	wire new_net_2799;
	wire n_1274_;
	wire new_net_3576;
	wire n_0770_;
	wire new_net_141;
	wire new_net_3414;
	wire new_net_2775;
	wire new_net_7245;
	wire new_net_7909;
	wire new_net_8027;
	wire new_net_8560;
	wire new_net_10092;
	wire new_net_3980;
	wire new_net_6459;
	wire new_net_3978;
	wire new_net_8725;
	wire new_net_9260;
	wire new_net_8615;
	wire new_net_7794;
	wire new_net_3485;
	wire new_net_2822;
	wire new_net_4090;
	wire new_net_4152;
	wire new_net_5915;
	wire new_net_6092;
	wire new_net_4622;
	wire new_net_7014;
	wire new_net_9864;
	wire new_net_9589;
	wire new_net_8845;
	wire new_net_6893;
	wire new_net_10109;
	wire new_net_7432;
	wire new_net_8742;
	wire new_net_10657;
	wire new_net_8377;
	wire n_1275_;
	wire n_0771_;
	wire n_0057_;
	wire n_0267_;
	wire n_0561_;
	wire new_net_476;
	wire new_net_1004;
	wire new_net_1647;
	wire n_1065_;
	wire new_net_560;
	wire new_net_6309;
	wire new_net_9724;
	wire new_net_10080;
	wire new_net_9336;
	wire new_net_4196;
	wire new_net_6021;
	wire new_net_5939;
	wire new_net_9208;
	wire new_net_7209;
	wire new_net_3133;
	wire new_net_2969;
	wire new_net_3153;
	wire new_net_708;
	wire new_net_2051;
	wire new_net_3765;
	wire new_net_3789;
	wire new_net_3807;
	wire new_net_4361;
	wire new_net_4893;
	wire new_net_4211;
	wire new_net_7343;
	wire new_net_3509;
	wire n_1276_;
	wire new_net_142;
	wire new_net_1793;
	wire new_net_3415;
	wire n_0772_;
	wire n_1066_;
	wire n_0058_;
	wire n_0268_;
	wire n_0562_;
	wire new_net_5208;
	wire new_net_8636;
	wire new_net_7933;
	wire new_net_5661;
	wire new_net_2240;
	wire new_net_2616;
	wire new_net_2303;
	wire new_net_593;
	wire new_net_2041;
	wire new_net_2158;
	wire new_net_2408;
	wire new_net_5203;
	wire new_net_5329;
	wire new_net_7680;
	wire new_net_8944;
	wire new_net_10203;
	wire new_net_6581;
	wire new_net_4884;
	wire new_net_4882;
	wire new_net_9972;
	wire new_net_4805;
	wire new_net_8245;
	wire new_net_7583;
	wire n_1277_;
	wire new_net_408;
	wire new_net_1534;
	wire n_0773_;
	wire n_1067_;
	wire n_0269_;
	wire n_0059_;
	wire n_0563_;
	wire new_net_477;
	wire new_net_741;
	wire new_net_5241;
	wire new_net_10225;
	wire new_net_9229;
	wire new_net_9448;
	wire new_net_10460;
	wire new_net_4781;
	wire new_net_3717;
	wire new_net_7845;
	wire new_net_3911;
	wire new_net_7726;
	wire new_net_986;
	wire new_net_3306;
	wire new_net_3816;
	wire new_net_2776;
	wire new_net_2800;
	wire new_net_3176;
	wire new_net_709;
	wire new_net_856;
	wire new_net_3577;
	wire new_net_2683;
	wire new_net_3432;
	wire new_net_2707;
	wire new_net_2729;
	wire new_net_8189;
	wire new_net_8430;
	wire new_net_4564;
	wire new_net_8601;
	wire new_net_8797;
	wire n_1068_;
	wire n_1278_;
	wire new_net_2823;
	wire n_0564_;
	wire n_0270_;
	wire n_0060_;
	wire n_0774_;
	wire new_net_143;
	wire new_net_2042;
	wire new_net_1794;
	wire new_net_4608;
	wire new_net_8121;
	wire new_net_9855;
	wire new_net_9111;
	wire new_net_7834;
	wire new_net_6884;
	wire new_net_7423;
	wire new_net_8733;
	wire new_net_5453;
	wire new_net_1648;
	wire new_net_3486;
	wire new_net_561;
	wire new_net_594;
	wire new_net_4317;
	wire new_net_4341;
	wire new_net_6080;
	wire new_net_6809;
	wire new_net_4715;
	wire new_net_7223;
	wire new_net_8880;
	wire new_net_9155;
	wire new_net_9322;
	wire new_net_4187;
	wire new_net_10503;
	wire new_net_6533;
	wire new_net_10632;
	wire new_net_4909;
	wire new_net_1418;
	wire n_1069_;
	wire n_0271_;
	wire new_net_3134;
	wire new_net_1974;
	wire new_net_2970;
	wire new_net_3154;
	wire n_1279_;
	wire new_net_409;
	wire new_net_1535;
	wire new_net_7657;
	wire new_net_9641;
	wire new_net_9815;
	wire new_net_7782;
	wire new_net_9541;
	wire new_net_4085;
	wire new_net_3416;
	wire new_net_3510;
	wire new_net_857;
	wire new_net_2155;
	wire new_net_3992;
	wire new_net_4072;
	wire new_net_5482;
	wire new_net_7503;
	wire new_net_7965;
	wire new_net_5197;
	wire new_net_8444;
	wire new_net_8622;
	wire new_net_7905;
	wire new_net_5552;
	wire new_net_9013;
	wire new_net_9283;
	wire n_1070_;
	wire new_net_2617;
	wire new_net_2052;
	wire n_0776_;
	wire n_0062_;
	wire n_0272_;
	wire n_1280_;
	wire new_net_144;
	wire n_0566_;
	wire new_net_4533;
	wire new_net_10194;
	wire new_net_4672;
	wire new_net_10351;
	wire new_net_10591;
	wire new_net_5438;
	wire new_net_8275;
	wire new_net_2409;
	wire new_net_1649;
	wire new_net_2241;
	wire new_net_2948;
	wire new_net_478;
	wire new_net_562;
	wire new_net_595;
	wire new_net_1006;
	wire new_net_2304;
	wire new_net_4116;
	wire new_net_7375;
	wire new_net_9035;
	wire new_net_10216;
	wire new_net_3405;
	wire new_net_9467;
	wire new_net_5909;
	wire new_net_8210;
	wire new_net_9465;
	wire new_net_9745;
	wire new_net_3898;
	wire new_net_3896;
	wire n_0063_;
	wire new_net_743;
	wire new_net_2708;
	wire new_net_1419;
	wire new_net_2730;
	wire new_net_2777;
	wire new_net_2957;
	wire new_net_3578;
	wire new_net_2801;
	wire n_0777_;
	wire new_net_8180;
	wire new_net_8537;
	wire new_net_3674;
	wire new_net_7768;
	wire new_net_8416;
	wire new_net_10301;
	wire new_net_9958;
	wire new_net_4149;
	wire new_net_8201;
	wire new_net_8593;
	wire new_net_172;
	wire new_net_2824;
	wire new_net_1795;
	wire new_net_4527;
	wire new_net_5917;
	wire new_net_6094;
	wire new_net_7016;
	wire new_net_8313;
	wire new_net_9068;
	wire new_net_10557;
	wire new_net_4734;
	wire new_net_9697;
	wire new_net_9102;
	wire new_net_7825;
	wire new_net_6144;
	wire new_net_5403;
	wire new_net_5319;
	wire new_net_2115;
	wire n_0568_;
	wire n_0778_;
	wire n_1072_;
	wire n_0274_;
	wire n_0064_;
	wire n_1282_;
	wire new_net_3177;
	wire new_net_145;
	wire new_net_4093;
	wire new_net_4971;
	wire new_net_7463;
	wire new_net_5500;
	wire n_0056_;
	wire new_net_2706;
	wire new_net_6519;
	wire new_net_9124;
	wire new_net_10383;
	wire new_net_7186;
	wire new_net_10623;
	wire new_net_6774;
	wire new_net_2949;
	wire new_net_3135;
	wire new_net_2971;
	wire new_net_3155;
	wire new_net_410;
	wire new_net_479;
	wire new_net_1007;
	wire new_net_1536;
	wire new_net_3767;
	wire new_net_3809;
	wire new_net_9526;
	wire new_net_7986;
	wire new_net_10511;
	wire new_net_7325;
	wire new_net_5041;
	wire new_net_711;
	wire n_0065_;
	wire n_1073_;
	wire new_net_3487;
	wire new_net_3511;
	wire n_0569_;
	wire n_0275_;
	wire new_net_858;
	wire n_1283_;
	wire n_0779_;
	wire new_net_4842;
	wire new_net_6633;
	wire new_net_5638;
	wire new_net_9004;
	wire new_net_10180;
	wire new_net_9514;
	wire new_net_2618;
	wire new_net_1796;
	wire new_net_4153;
	wire new_net_5205;
	wire new_net_7682;
	wire new_net_8010;
	wire new_net_8034;
	wire new_net_8826;
	wire new_net_4628;
	wire new_net_10582;
	wire new_net_6614;
	wire new_net_7855;
	wire new_net_7441;
	wire new_net_7561;
	wire new_net_10666;
	wire new_net_146;
	wire n_0066_;
	wire new_net_1650;
	wire new_net_563;
	wire n_0276_;
	wire new_net_596;
	wire n_0780_;
	wire n_1074_;
	wire n_0570_;
	wire n_1284_;
	wire new_net_5107;
	wire new_net_5803;
	wire new_net_4488;
	wire new_net_7616;
	wire new_net_8475;
	wire new_net_7997;
	wire new_net_7297;
	wire new_net_2685;
	wire new_net_2305;
	wire new_net_1537;
	wire new_net_2410;
	wire new_net_2709;
	wire new_net_2731;
	wire new_net_3579;
	wire new_net_2242;
	wire new_net_2778;
	wire new_net_1420;
	wire new_net_4659;
	wire new_net_10067;
	wire new_net_8400;
	wire new_net_8407;
	wire new_net_9664;
	wire new_net_6377;
	wire new_net_7269;
	wire new_net_7267;
	wire new_net_9831;
	wire new_net_6263;
	wire new_net_6204;
	wire new_net_8779;
	wire new_net_8100;
	wire new_net_10543;
	wire n_0067_;
	wire n_0277_;
	wire n_0781_;
	wire n_1075_;
	wire n_0571_;
	wire new_net_859;
	wire n_1285_;
	wire new_net_2825;
	wire new_net_4528;
	wire new_net_5720;
	wire new_net_10152;
	wire new_net_6863;
	wire new_net_9886;
	wire new_net_8864;
	wire new_net_2184;
	wire new_net_3178;
	wire new_net_2157;
	wire new_net_4319;
	wire new_net_4343;
	wire new_net_6082;
	wire new_net_6811;
	wire new_net_7366;
	wire new_net_7390;
	wire new_net_7512;
	wire new_net_8688;
	wire new_net_8761;
	wire new_net_6510;
	wire new_net_7172;
	wire new_net_7635;
	wire new_net_147;
	wire n_0572_;
	wire new_net_2044;
	wire n_0068_;
	wire new_net_1651;
	wire new_net_564;
	wire n_0782_;
	wire n_1076_;
	wire n_0278_;
	wire new_net_597;
	wire new_net_3766;
	wire new_net_5963;
	wire new_net_7690;
	wire new_net_8975;
	wire n_0816_;
	wire new_net_9836;
	wire new_net_6173;
	wire new_net_9377;
	wire new_net_712;
	wire new_net_745;
	wire new_net_1421;
	wire new_net_3488;
	wire new_net_412;
	wire new_net_481;
	wire new_net_3512;
	wire new_net_4074;
	wire new_net_4526;
	wire new_net_5484;
	wire new_net_5692;
	wire new_net_8901;
	wire new_net_4029;
	wire new_net_9691;
	wire new_net_5529;
	wire new_net_1715;
	wire new_net_8660;
	wire new_net_7957;
	wire n_1287_;
	wire new_net_1797;
	wire new_net_3434;
	wire n_0069_;
	wire n_0573_;
	wire n_0783_;
	wire n_1077_;
	wire n_0279_;
	wire new_net_2619;
	wire new_net_5206;
	wire new_net_9785;
	wire new_net_10131;
	wire n_1200_;
	wire new_net_10568;
	wire new_net_4750;
	wire new_net_5374;
	wire new_net_5415;
	wire new_net_6036;
	wire new_net_9594;
	wire new_net_5372;
	wire new_net_7846;
	wire new_net_9998;
	wire new_net_9996;
	wire new_net_2168;
	wire new_net_4095;
	wire new_net_3817;
	wire new_net_4118;
	wire new_net_4829;
	wire new_net_5695;
	wire new_net_5751;
	wire new_net_6401;
	wire new_net_7226;
	wire new_net_5066;
	wire new_net_9913;
	wire new_net_4512;
	wire new_net_7607;
	wire n_0670_;
	wire new_net_5260;
	wire new_net_5886;
	wire n_1288_;
	wire new_net_1538;
	wire n_0784_;
	wire new_net_148;
	wire new_net_3417;
	wire new_net_3580;
	wire new_net_2686;
	wire n_0070_;
	wire new_net_2710;
	wire new_net_2732;
	wire new_net_6792;
	wire new_net_7750;
	wire n_1020_;
	wire new_net_6363;
	wire new_net_9935;
	wire new_net_10278;
	wire new_net_8570;
	wire new_net_4041;
	wire new_net_10024;
	wire new_net_8091;
	wire new_net_6192;
	wire new_net_558;
	wire new_net_10534;
	wire new_net_2306;
	wire new_net_2826;
	wire new_net_2411;
	wire new_net_482;
	wire new_net_713;
	wire new_net_860;
	wire new_net_2243;
	wire new_net_4529;
	wire new_net_4930;
	wire new_net_5919;
	wire new_net_10338;
	wire new_net_3862;
	wire new_net_6121;
	wire new_net_5756;
	wire new_net_4948;
	wire new_net_6908;
	wire n_1289_;
	wire new_net_1798;
	wire n_0575_;
	wire n_0071_;
	wire new_net_3179;
	wire n_0785_;
	wire n_1079_;
	wire n_0281_;
	wire new_net_4320;
	wire new_net_4344;
	wire new_net_5479;
	wire new_net_5477;
	wire new_net_8684;
	wire new_net_6319;
	wire new_net_2950;
	wire new_net_7163;
	wire new_net_9346;
	wire new_net_2973;
	wire new_net_3157;
	wire new_net_598;
	wire new_net_2951;
	wire new_net_3769;
	wire new_net_3811;
	wire new_net_4365;
	wire new_net_4938;
	wire new_net_6557;
	wire new_net_7868;
	wire new_net_8966;
	wire new_net_2795;
	wire new_net_7473;
	wire new_net_6813;
	wire new_net_4309;
	wire n_1290_;
	wire new_net_1422;
	wire n_0786_;
	wire new_net_149;
	wire new_net_2015;
	wire new_net_3418;
	wire new_net_1010;
	wire n_0576_;
	wire new_net_1539;
	wire new_net_746;
	wire new_net_3251;
	wire new_net_9682;
	wire new_net_6493;
	wire new_net_9064;
	wire new_net_8646;
	wire new_net_7943;
	wire new_net_9844;
	wire new_net_6664;
	wire new_net_10056;
	wire new_net_2620;
	wire new_net_483;
	wire new_net_714;
	wire new_net_861;
	wire new_net_5207;
	wire new_net_7684;
	wire new_net_7989;
	wire new_net_8012;
	wire new_net_8036;
	wire new_net_8847;
	wire new_net_9307;
	wire new_net_9580;
	wire new_net_10375;
	wire new_net_10368;
	wire new_net_3136;
	wire n_1291_;
	wire n_0787_;
	wire new_net_1799;
	wire n_0073_;
	wire n_0283_;
	wire n_0577_;
	wire n_1081_;
	wire new_net_4096;
	wire new_net_4119;
	wire new_net_6686;
	wire new_net_5836;
	wire new_net_8706;
	wire new_net_9052;
	wire new_net_9602;
	wire new_net_7679;
	wire n_0817_;
	wire new_net_10470;
	wire new_net_8853;
	wire new_net_9244;
	wire new_net_10117;
	wire new_net_2780;
	wire new_net_2804;
	wire new_net_3581;
	wire new_net_2687;
	wire new_net_3435;
	wire new_net_2711;
	wire new_net_599;
	wire new_net_2045;
	wire new_net_2165;
	wire new_net_2733;
	wire new_net_3921;
	wire new_net_7736;
	wire new_net_8386;
	wire new_net_8028;
	wire new_net_7246;
	wire new_net_4406;
	wire new_net_7244;
	wire new_net_8561;
	wire new_net_6460;
	wire new_net_10093;
	wire new_net_9619;
	wire new_net_8726;
	wire new_net_5704;
	wire new_net_8616;
	wire n_1292_;
	wire new_net_414;
	wire new_net_2827;
	wire n_0788_;
	wire new_net_150;
	wire n_0578_;
	wire new_net_747;
	wire n_0074_;
	wire n_0284_;
	wire new_net_1423;
	wire new_net_7795;
	wire new_net_4623;
	wire new_net_8699;
	wire new_net_7964;
	wire new_net_9865;
	wire new_net_9189;
	wire new_net_6894;
	wire new_net_10110;
	wire new_net_4939;
	wire new_net_7433;
	wire new_net_8743;
	wire new_net_10658;
	wire new_net_2244;
	wire new_net_2063;
	wire new_net_2307;
	wire new_net_3180;
	wire new_net_2412;
	wire new_net_4321;
	wire new_net_4345;
	wire new_net_6084;
	wire new_net_6403;
	wire new_net_6407;
	wire new_net_6310;
	wire new_net_10081;
	wire new_net_9337;
	wire new_net_2728;
	wire new_net_9211;
	wire new_net_4197;
	wire new_net_4762;
	wire new_net_5940;
	wire new_net_9209;
	wire new_net_2952;
	wire new_net_3137;
	wire new_net_2974;
	wire new_net_3158;
	wire n_1293_;
	wire new_net_1800;
	wire n_0579_;
	wire n_0789_;
	wire n_1083_;
	wire n_0285_;
	wire new_net_7210;
	wire new_net_10027;
	wire new_net_4295;
	wire new_net_6804;
	wire new_net_3490;
	wire new_net_3514;
	wire new_net_567;
	wire new_net_1011;
	wire new_net_1540;
	wire new_net_1654;
	wire new_net_4076;
	wire new_net_4897;
	wire new_net_5486;
	wire new_net_7969;
	wire new_net_7513;
	wire new_net_4006;
	wire new_net_7025;
	wire new_net_5506;
	wire new_net_4866;
	wire new_net_8637;
	wire new_net_7023;
	wire new_net_7934;
	wire new_net_5662;
	wire new_net_10047;
	wire n_1084_;
	wire new_net_2621;
	wire new_net_862;
	wire new_net_1979;
	wire n_1294_;
	wire new_net_151;
	wire n_0580_;
	wire new_net_484;
	wire new_net_715;
	wire n_0286_;
	wire new_net_8945;
	wire new_net_10204;
	wire new_net_5349;
	wire new_net_6582;
	wire new_net_9973;
	wire new_net_8246;
	wire new_net_2075;
	wire new_net_4097;
	wire new_net_4120;
	wire new_net_4164;
	wire new_net_5697;
	wire new_net_5753;
	wire new_net_7228;
	wire new_net_8376;
	wire new_net_7584;
	wire new_net_8498;
	wire new_net_3230;
	wire new_net_10226;
	wire new_net_9230;
	wire new_net_10461;
	wire n_1085_;
	wire new_net_600;
	wire new_net_2781;
	wire new_net_2805;
	wire n_1295_;
	wire new_net_2734;
	wire n_0791_;
	wire new_net_3582;
	wire new_net_2688;
	wire new_net_3436;
	wire new_net_7727;
	wire new_net_6345;
	wire new_net_6030;
	wire new_net_8190;
	wire new_net_5706;
	wire new_net_6446;
	wire new_net_8431;
	wire new_net_8602;
	wire new_net_1655;
	wire new_net_2828;
	wire new_net_415;
	wire new_net_568;
	wire new_net_748;
	wire new_net_1012;
	wire new_net_1983;
	wire new_net_1541;
	wire new_net_4531;
	wire new_net_5921;
	wire new_net_8798;
	wire new_net_8796;
	wire new_net_10322;
	wire new_net_6105;
	wire new_net_9856;
	wire new_net_9112;
	wire new_net_7835;
	wire new_net_7424;
	wire new_net_8734;
	wire n_1086_;
	wire new_net_863;
	wire new_net_2064;
	wire n_1296_;
	wire new_net_3181;
	wire n_0792_;
	wire new_net_152;
	wire new_net_2018;
	wire n_0078_;
	wire n_0288_;
	wire new_net_4718;
	wire new_net_5454;
	wire new_net_4384;
	wire new_net_5618;
	wire new_net_8881;
	wire new_net_9156;
	wire new_net_5616;
	wire new_net_4188;
	wire new_net_10504;
	wire new_net_6534;
	wire new_net_2245;
	wire new_net_2953;
	wire new_net_2975;
	wire new_net_3159;
	wire new_net_2308;
	wire new_net_1801;
	wire new_net_2173;
	wire new_net_2413;
	wire new_net_3771;
	wire new_net_3813;
	wire new_net_4910;
	wire new_net_7658;
	wire new_net_9642;
	wire new_net_3790;
	wire new_net_9816;
	wire new_net_4999;
	wire new_net_716;
	wire new_net_9542;
	wire new_net_3491;
	wire new_net_601;
	wire new_net_3515;
	wire n_1297_;
	wire n_0793_;
	wire n_1087_;
	wire n_0289_;
	wire n_0079_;
	wire n_0583_;
	wire new_net_4077;
	wire new_net_10415;
	wire new_net_10413;
	wire new_net_8445;
	wire new_net_8623;
	wire new_net_1656;
	wire new_net_2622;
	wire new_net_416;
	wire new_net_749;
	wire new_net_1425;
	wire new_net_5209;
	wire new_net_5546;
	wire new_net_5553;
	wire new_net_7686;
	wire new_net_7991;
	wire new_net_9014;
	wire new_net_9284;
	wire new_net_10195;
	wire new_net_10352;
	wire n_0402_;
	wire new_net_3556;
	wire new_net_7106;
	wire new_net_10592;
	wire new_net_5439;
	wire new_net_4797;
	wire new_net_6053;
	wire new_net_2627;
	wire n_1298_;
	wire new_net_153;
	wire n_0794_;
	wire n_1088_;
	wire n_0290_;
	wire n_0080_;
	wire n_0584_;
	wire new_net_486;
	wire new_net_4098;
	wire new_net_5813;
	wire new_net_9036;
	wire new_net_1020;
	wire new_net_1663;
	wire new_net_10217;
	wire new_net_9468;
	wire new_net_5910;
	wire new_net_9746;
	wire new_net_559;
	wire new_net_2170;
	wire new_net_2713;
	wire new_net_2735;
	wire new_net_2782;
	wire new_net_2806;
	wire new_net_1802;
	wire new_net_3419;
	wire new_net_2689;
	wire new_net_3437;
	wire new_net_3791;
	wire new_net_6336;
	wire new_net_8181;
	wire new_net_3958;
	wire new_net_8417;
	wire new_net_10302;
	wire new_net_1695;
	wire new_net_3120;
	wire new_net_6387;
	wire new_net_9959;
	wire new_net_10234;
	wire n_1097_;
	wire new_net_4150;
	wire new_net_8594;
	wire new_net_1013;
	wire n_1089_;
	wire n_1299_;
	wire new_net_1542;
	wire new_net_2829;
	wire n_0585_;
	wire n_0291_;
	wire n_0081_;
	wire n_0795_;
	wire new_net_591;
	wire new_net_6091;
	wire new_net_8754;
	wire new_net_10558;
	wire new_net_8314;
	wire new_net_4735;
	wire new_net_9103;
	wire new_net_7826;
	wire new_net_7043;
	wire new_net_6145;
	wire new_net_8360;
	wire new_net_1426;
	wire new_net_864;
	wire new_net_2047;
	wire new_net_717;
	wire new_net_750;
	wire new_net_4323;
	wire new_net_5404;
	wire new_net_6086;
	wire new_net_6815;
	wire new_net_5320;
	wire new_net_4972;
	wire new_net_6287;
	wire n_0338_;
	wire new_net_5501;
	wire new_net_2700;
	wire new_net_2972;
	wire new_net_6520;
	wire new_net_7187;
	wire new_net_487;
	wire new_net_2954;
	wire n_1300_;
	wire new_net_3160;
	wire n_0586_;
	wire n_0796_;
	wire n_1090_;
	wire n_0292_;
	wire n_0082_;
	wire new_net_2976;
	wire new_net_10624;
	wire new_net_9527;
	wire new_net_1296;
	wire new_net_7987;
	wire new_net_10512;
	wire new_net_7326;
	wire new_net_2414;
	wire new_net_3492;
	wire new_net_2246;
	wire new_net_3516;
	wire new_net_2309;
	wire new_net_602;
	wire new_net_2019;
	wire new_net_3420;
	wire new_net_4078;
	wire new_net_4899;
	wire new_net_8234;
	wire new_net_1014;
	wire new_net_1657;
	wire n_1091_;
	wire n_1301_;
	wire new_net_417;
	wire new_net_1543;
	wire n_0797_;
	wire n_0587_;
	wire n_0293_;
	wire n_0083_;
	wire new_net_9515;
	wire new_net_9906;
	wire new_net_10181;
	wire new_net_8458;
	wire new_net_9130;
	wire new_net_1427;
	wire new_net_3138;
	wire new_net_2624;
	wire new_net_718;
	wire new_net_751;
	wire new_net_865;
	wire new_net_2862;
	wire new_net_4099;
	wire new_net_4122;
	wire new_net_5699;
	wire new_net_174;
	wire new_net_7362;
	wire new_net_7617;
	wire new_net_6397;
	wire new_net_7998;
	wire new_net_155;
	wire new_net_1803;
	wire n_0588_;
	wire new_net_2690;
	wire n_0084_;
	wire new_net_2714;
	wire new_net_2140;
	wire new_net_2736;
	wire new_net_2807;
	wire new_net_2783;
	wire new_net_7298;
	wire new_net_8167;
	wire new_net_10068;
	wire new_net_4660;
	wire new_net_8408;
	wire new_net_3943;
	wire new_net_6378;
	wire new_net_9665;
	wire new_net_7270;
	wire new_net_4430;
	wire new_net_7268;
	wire new_net_9832;
	wire new_net_6264;
	wire new_net_8780;
	wire new_net_8101;
	wire new_net_603;
	wire new_net_2095;
	wire new_net_2123;
	wire new_net_2830;
	wire new_net_5923;
	wire new_net_6100;
	wire new_net_6408;
	wire new_net_7022;
	wire new_net_8995;
	wire new_net_9088;
	wire new_net_9631;
	wire new_net_5728;
	wire new_net_10544;
	wire new_net_5721;
	wire new_net_10609;
	wire new_net_6864;
	wire new_net_4673;
	wire new_net_6131;
	wire n_0589_;
	wire n_0085_;
	wire new_net_1015;
	wire new_net_1658;
	wire new_net_411;
	wire n_0295_;
	wire n_0799_;
	wire n_1093_;
	wire n_1303_;
	wire new_net_418;
	wire new_net_7120;
	wire new_net_4366;
	wire new_net_8762;
	wire new_net_10100;
	wire new_net_6511;
	wire new_net_7173;
	wire new_net_2955;
	wire new_net_2977;
	wire new_net_3161;
	wire new_net_488;
	wire new_net_3773;
	wire new_net_3815;
	wire new_net_4369;
	wire new_net_4942;
	wire new_net_6404;
	wire new_net_7872;
	wire new_net_5964;
	wire new_net_8460;
	wire new_net_7691;
	wire new_net_8976;
	wire new_net_7689;
	wire new_net_9837;
	wire n_1304_;
	wire n_0800_;
	wire new_net_156;
	wire new_net_1804;
	wire new_net_3421;
	wire new_net_2049;
	wire n_0086_;
	wire n_1094_;
	wire new_net_3493;
	wire n_0296_;
	wire new_net_6174;
	wire new_net_9378;
	wire new_net_5693;
	wire new_net_8902;
	wire new_net_4030;
	wire new_net_7784;
	wire new_net_9692;
	wire new_net_5530;
	wire new_net_2310;
	wire new_net_2415;
	wire new_net_2247;
	wire new_net_604;
	wire new_net_5211;
	wire new_net_7688;
	wire new_net_8016;
	wire new_net_7958;
	wire new_net_8040;
	wire new_net_8996;
	wire new_net_9786;
	wire new_net_10132;
	wire new_net_10569;
	wire new_net_9595;
	wire new_net_4751;
	wire new_net_5375;
	wire new_net_5416;
	wire new_net_6037;
	wire new_net_8846;
	wire new_net_2046;
	wire new_net_5373;
	wire n_1305_;
	wire new_net_419;
	wire n_0801_;
	wire new_net_719;
	wire new_net_2048;
	wire n_0087_;
	wire new_net_752;
	wire new_net_1016;
	wire new_net_1428;
	wire n_1095_;
	wire new_net_9997;
	wire new_net_8381;
	wire new_net_9914;
	wire new_net_3298;
	wire new_net_10473;
	wire new_net_455;
	wire new_net_7608;
	wire new_net_10434;
	wire new_net_5261;
	wire new_net_9725;
	wire new_net_5887;
	wire new_net_2715;
	wire new_net_2020;
	wire new_net_2691;
	wire new_net_2808;
	wire new_net_2737;
	wire new_net_2784;
	wire new_net_489;
	wire new_net_4511;
	wire new_net_3654;
	wire new_net_5336;
	wire new_net_9073;
	wire new_net_10279;
	wire new_net_6793;
	wire new_net_3182;
	wire new_net_6364;
	wire new_net_7751;
	wire new_net_9936;
	wire new_net_10486;
	wire new_net_8571;
	wire new_net_6195;
	wire new_net_10025;
	wire new_net_8092;
	wire n_1306_;
	wire new_net_2831;
	wire new_net_157;
	wire n_0592_;
	wire n_0088_;
	wire n_0298_;
	wire n_0802_;
	wire n_1096_;
	wire new_net_5924;
	wire new_net_6101;
	wire new_net_8923;
	wire new_net_9551;
	wire new_net_10535;
	wire new_net_807;
	wire new_net_10339;
	wire new_net_8855;
	wire new_net_89;
	wire new_net_5757;
	wire new_net_8341;
	wire new_net_1545;
	wire new_net_1659;
	wire new_net_4325;
	wire new_net_4534;
	wire new_net_6817;
	wire new_net_7348;
	wire new_net_4949;
	wire new_net_7372;
	wire new_net_7396;
	wire new_net_7518;
	wire new_net_5478;
	wire new_net_8685;
	wire new_net_5983;
	wire new_net_6320;
	wire new_net_8827;
	wire new_net_2582;
	wire n_1163_;
	wire new_net_867;
	wire n_1307_;
	wire n_0593_;
	wire new_net_720;
	wire new_net_2089;
	wire n_0089_;
	wire new_net_753;
	wire new_net_1429;
	wire new_net_573;
	wire new_net_3162;
	wire new_net_4496;
	wire new_net_5950;
	wire new_net_7215;
	wire new_net_6558;
	wire new_net_6551;
	wire new_net_7895;
	wire n_1204_;
	wire new_net_8967;
	wire n_0061_;
	wire new_net_388;
	wire new_net_5023;
	wire new_net_5021;
	wire new_net_1805;
	wire new_net_3422;
	wire new_net_3494;
	wire new_net_490;
	wire new_net_4080;
	wire new_net_4346;
	wire new_net_4901;
	wire new_net_5490;
	wire new_net_6205;
	wire new_net_6814;
	wire new_net_9683;
	wire n_0404_;
	wire new_net_8647;
	wire n_0300_;
	wire new_net_605;
	wire n_1308_;
	wire new_net_158;
	wire new_net_3583;
	wire n_0090_;
	wire n_0594_;
	wire n_0804_;
	wire n_1098_;
	wire new_net_4156;
	wire new_net_5672;
	wire new_net_7944;
	wire new_net_10057;
	wire new_net_1424;
	wire new_net_10645;
	wire new_net_9308;
	wire n_1024_;
	wire new_net_1021;
	wire new_net_1664;
	wire new_net_9581;
	wire new_net_9306;
	wire new_net_7464;
	wire new_net_311;
	wire new_net_10376;
	wire new_net_10369;
	wire new_net_2248;
	wire new_net_3139;
	wire new_net_1546;
	wire new_net_2311;
	wire new_net_2416;
	wire new_net_1660;
	wire new_net_420;
	wire new_net_1017;
	wire new_net_4101;
	wire new_net_4124;
	wire new_net_6079;
	wire new_net_4821;
	wire new_net_6687;
	wire new_net_5058;
	wire new_net_7594;
	wire new_net_5837;
	wire new_net_5878;
	wire new_net_9053;
	wire new_net_8343;
	wire n_1099_;
	wire new_net_10471;
	wire new_net_9245;
	wire new_net_8854;
	wire n_0301_;
	wire new_net_2785;
	wire new_net_1984;
	wire new_net_2628;
	wire new_net_2809;
	wire n_1309_;
	wire n_0805_;
	wire new_net_2692;
	wire n_0091_;
	wire new_net_2716;
	wire new_net_8151;
	wire new_net_8149;
	wire new_net_592;
	wire new_net_8031;
	wire new_net_7737;
	wire new_net_8029;
	wire new_net_9571;
	wire new_net_7247;
	wire new_net_4407;
	wire new_net_3982;
	wire new_net_6461;
	wire new_net_2832;
	wire new_net_1806;
	wire new_net_491;
	wire new_net_5925;
	wire new_net_6102;
	wire new_net_6504;
	wire new_net_7024;
	wire new_net_8997;
	wire new_net_9620;
	wire new_net_10485;
	wire new_net_8617;
	wire new_net_7796;
	wire new_net_8700;
	wire new_net_9866;
	wire new_net_9190;
	wire n_0302_;
	wire new_net_606;
	wire new_net_1988;
	wire n_1310_;
	wire new_net_159;
	wire new_net_3584;
	wire n_0596_;
	wire n_0092_;
	wire new_net_2050;
	wire n_0806_;
	wire new_net_4940;
	wire new_net_7434;
	wire new_net_8744;
	wire new_net_6311;
	wire new_net_10082;
	wire new_net_1297;
	wire new_net_9338;
	wire new_net_9212;
	wire new_net_2979;
	wire new_net_3163;
	wire new_net_2043;
	wire new_net_2169;
	wire new_net_1018;
	wire new_net_1430;
	wire new_net_421;
	wire new_net_574;
	wire new_net_721;
	wire new_net_754;
	wire new_net_4198;
	wire new_net_6023;
	wire new_net_9210;
	wire new_net_7211;
	wire new_net_9393;
	wire new_net_4296;
	wire new_net_7345;
	wire new_net_7514;
	wire new_net_4007;
	wire new_net_4869;
	wire new_net_5210;
	wire new_net_7026;
	wire new_net_5507;
	wire new_net_8638;
	wire new_net_7935;
	wire new_net_10048;
	wire n_0345_;
	wire n_0849_;
	wire new_net_1034;
	wire new_net_1938;
	wire new_net_3371;
	wire n_1353_;
	wire new_net_1332;
	wire new_net_175;
	wire new_net_3676;
	wire new_net_5109;
	wire new_net_8946;
	wire new_net_10205;
	wire new_net_8270;
	wire new_net_8247;
	wire new_net_4165;
	wire new_net_7875;
	wire new_net_54;
	wire new_net_885;
	wire new_net_1962;
	wire new_net_1678;
	wire new_net_2927;
	wire new_net_2068;
	wire new_net_1300;
	wire new_net_3718;
	wire new_net_4716;
	wire new_net_5981;
	wire new_net_5243;
	wire new_net_7386;
	wire new_net_10227;
	wire new_net_9231;
	wire new_net_9478;
	wire new_net_10462;
	wire new_net_10384;
	wire new_net_3913;
	wire n_0346_;
	wire n_0850_;
	wire new_net_286;
	wire new_net_1184;
	wire n_1354_;
	wire new_net_439;
	wire new_net_2661;
	wire new_net_244;
	wire new_net_1151;
	wire new_net_3308;
	wire new_net_6346;
	wire new_net_10153;
	wire new_net_8191;
	wire new_net_6447;
	wire new_net_8432;
	wire new_net_8603;
	wire new_net_8799;
	wire new_net_10323;
	wire new_net_623;
	wire new_net_2207;
	wire new_net_3238;
	wire new_net_2480;
	wire new_net_2751;
	wire new_net_1824;
	wire new_net_2375;
	wire new_net_3741;
	wire new_net_4002;
	wire new_net_4026;
	wire new_net_4610;
	wire new_net_9857;
	wire new_net_8213;
	wire new_net_9113;
	wire new_net_7836;
	wire new_net_8128;
	wire new_net_7425;
	wire new_net_8735;
	wire n_0347_;
	wire n_0851_;
	wire new_net_1035;
	wire new_net_1447;
	wire new_net_2066;
	wire n_1355_;
	wire new_net_1564;
	wire new_net_4719;
	wire new_net_4765;
	wire new_net_5938;
	wire new_net_7144;
	wire new_net_8882;
	wire new_net_9157;
	wire new_net_9712;
	wire new_net_9324;
	wire n_1100_;
	wire new_net_8342;
	wire new_net_10505;
	wire new_net_10669;
	wire new_net_6535;
	wire new_net_10634;
	wire new_net_10667;
	wire new_net_55;
	wire new_net_319;
	wire new_net_886;
	wire new_net_1964;
	wire new_net_1679;
	wire new_net_3109;
	wire n_0266_;
	wire new_net_1301;
	wire new_net_4048;
	wire new_net_4585;
	wire new_net_7659;
	wire new_net_9817;
	wire new_net_5000;
	wire new_net_9543;
	wire new_net_10416;
	wire n_0348_;
	wire n_0852_;
	wire new_net_245;
	wire new_net_1152;
	wire new_net_287;
	wire new_net_1185;
	wire new_net_2912;
	wire new_net_2591;
	wire new_net_3350;
	wire n_1356_;
	wire new_net_4087;
	wire new_net_7505;
	wire new_net_8446;
	wire new_net_10414;
	wire new_net_8624;
	wire new_net_5554;
	wire new_net_9015;
	wire new_net_5547;
	wire new_net_624;
	wire new_net_1333;
	wire new_net_3372;
	wire new_net_1939;
	wire new_net_2281;
	wire new_net_2344;
	wire new_net_1825;
	wire new_net_3677;
	wire new_net_3719;
	wire new_net_6219;
	wire new_net_10196;
	wire new_net_10353;
	wire new_net_10595;
	wire new_net_7114;
	wire new_net_10593;
	wire new_net_5440;
	wire n_0349_;
	wire n_0853_;
	wire new_net_1448;
	wire n_1357_;
	wire new_net_1565;
	wire new_net_2027;
	wire new_net_4688;
	wire new_net_4717;
	wire new_net_5982;
	wire new_net_7574;
	wire new_net_7377;
	wire new_net_8689;
	wire new_net_9037;
	wire new_net_10218;
	wire new_net_9469;
	wire new_net_5911;
	wire new_net_8008;
	wire new_net_320;
	wire new_net_1680;
	wire new_net_2097;
	wire new_net_2662;
	wire new_net_4568;
	wire new_net_5224;
	wire new_net_5771;
	wire new_net_5795;
	wire new_net_6337;
	wire new_net_6436;
	wire new_net_8182;
	wire new_net_8418;
	wire new_net_10303;
	wire new_net_6388;
	wire new_net_8595;
	wire n_0854_;
	wire n_0350_;
	wire new_net_246;
	wire new_net_1153;
	wire new_net_3239;
	wire new_net_288;
	wire new_net_1186;
	wire new_net_2752;
	wire n_1358_;
	wire new_net_3742;
	wire new_net_8315;
	wire new_net_8755;
	wire new_net_10559;
	wire new_net_9104;
	wire new_net_7827;
	wire new_net_7044;
	wire new_net_10252;
	wire new_net_625;
	wire new_net_1334;
	wire new_net_1826;
	wire new_net_2376;
	wire new_net_2208;
	wire new_net_2481;
	wire new_net_1940;
	wire new_net_2529;
	wire new_net_3394;
	wire new_net_4766;
	wire new_net_4973;
	wire new_net_5502;
	wire new_net_6000;
	wire new_net_6521;
	wire new_net_7188;
	wire new_net_10625;
	wire new_net_4851;
	wire n_0351_;
	wire n_0855_;
	wire new_net_1036;
	wire new_net_1449;
	wire new_net_3110;
	wire new_net_56;
	wire new_net_887;
	wire new_net_1302;
	wire n_1359_;
	wire new_net_4049;
	wire new_net_10436;
	wire new_net_8235;
	wire new_net_321;
	wire new_net_441;
	wire new_net_1999;
	wire new_net_2928;
	wire new_net_3351;
	wire new_net_4220;
	wire new_net_4243;
	wire new_net_4284;
	wire new_net_4547;
	wire new_net_4958;
	wire new_net_9006;
	wire n_1360_;
	wire n_0352_;
	wire n_0856_;
	wire new_net_247;
	wire new_net_1154;
	wire new_net_3373;
	wire new_net_3678;
	wire new_net_6220;
	wire new_net_6244;
	wire new_net_7910;
	wire new_net_9516;
	wire new_net_10182;
	wire new_net_7857;
	wire new_net_2345;
	wire new_net_1335;
	wire new_net_1566;
	wire new_net_1827;
	wire new_net_2592;
	wire new_net_2080;
	wire new_net_2282;
	wire new_net_2863;
	wire new_net_3735;
	wire new_net_4689;
	wire new_net_5805;
	wire new_net_7363;
	wire new_net_4490;
	wire new_net_7618;
	wire new_net_5271;
	wire new_net_8479;
	wire new_net_5902;
	wire new_net_8477;
	wire new_net_7707;
	wire new_net_7999;
	wire n_0353_;
	wire n_0857_;
	wire n_1361_;
	wire new_net_2663;
	wire new_net_2024;
	wire new_net_1450;
	wire new_net_1681;
	wire new_net_57;
	wire new_net_888;
	wire new_net_1303;
	wire new_net_4661;
	wire new_net_8168;
	wire new_net_10069;
	wire new_net_8409;
	wire new_net_6379;
	wire new_net_7271;
	wire new_net_4431;
	wire new_net_8781;
	wire new_net_8102;
	wire new_net_4594;
	wire new_net_289;
	wire new_net_322;
	wire new_net_442;
	wire new_net_1037;
	wire new_net_1187;
	wire new_net_2003;
	wire new_net_3240;
	wire new_net_2753;
	wire new_net_2079;
	wire new_net_3743;
	wire new_net_5722;
	wire new_net_9632;
	wire new_net_10154;
	wire new_net_4106;
	wire new_net_6865;
	wire new_net_6132;
	wire new_net_8866;
	wire n_0858_;
	wire n_0354_;
	wire n_1362_;
	wire new_net_248;
	wire new_net_1155;
	wire new_net_2185;
	wire new_net_1941;
	wire new_net_626;
	wire new_net_3720;
	wire new_net_4367;
	wire new_net_5312;
	wire new_net_7091;
	wire new_net_8211;
	wire new_net_10101;
	wire new_net_7174;
	wire new_net_1567;
	wire new_net_2209;
	wire new_net_2377;
	wire new_net_2482;
	wire new_net_3111;
	wire new_net_4050;
	wire new_net_3768;
	wire new_net_4695;
	wire new_net_4736;
	wire new_net_4800;
	wire new_net_7637;
	wire new_net_7692;
	wire new_net_8977;
	wire new_net_9603;
	wire new_net_3395;
	wire new_net_58;
	wire n_0859_;
	wire n_0355_;
	wire n_1363_;
	wire new_net_2182;
	wire new_net_1961;
	wire new_net_3352;
	wire new_net_1451;
	wire new_net_1682;
	wire n_0546_;
	wire new_net_5694;
	wire new_net_8271;
	wire new_net_8903;
	wire new_net_4031;
	wire new_net_9693;
	wire new_net_5531;
	wire new_net_9262;
	wire new_net_3374;
	wire new_net_290;
	wire new_net_443;
	wire new_net_1188;
	wire new_net_2581;
	wire new_net_3679;
	wire new_net_6221;
	wire new_net_6245;
	wire new_net_7959;
	wire new_net_9319;
	wire new_net_9787;
	wire new_net_10412;
	wire new_net_10570;
	wire new_net_4752;
	wire new_net_5376;
	wire new_net_6038;
	wire new_net_8217;
	wire new_net_9596;
	wire new_net_10464;
	wire new_net_7848;
	wire new_net_10000;
	wire new_net_627;
	wire n_0356_;
	wire n_0860_;
	wire n_1364_;
	wire new_net_1336;
	wire new_net_1828;
	wire new_net_249;
	wire new_net_2593;
	wire new_net_1942;
	wire new_net_3819;
	wire new_net_8673;
	wire new_net_7899;
	wire new_net_4476;
	wire new_net_5068;
	wire new_net_4129;
	wire new_net_5262;
	wire new_net_9726;
	wire new_net_10435;
	wire new_net_5847;
	wire new_net_5888;
	wire new_net_2283;
	wire new_net_889;
	wire new_net_1304;
	wire new_net_2346;
	wire new_net_2664;
	wire new_net_4570;
	wire new_net_5226;
	wire new_net_5773;
	wire new_net_5797;
	wire new_net_6438;
	wire new_net_10280;
	wire new_net_6794;
	wire new_net_7752;
	wire new_net_4536;
	wire new_net_6365;
	wire new_net_9937;
	wire new_net_10487;
	wire new_net_7919;
	wire new_net_8574;
	wire new_net_8572;
	wire new_net_6196;
	wire new_net_10026;
	wire new_net_8093;
	wire new_net_6194;
	wire n_0357_;
	wire n_0861_;
	wire n_1365_;
	wire new_net_3241;
	wire new_net_323;
	wire new_net_1038;
	wire new_net_1683;
	wire new_net_2754;
	wire new_net_3744;
	wire new_net_4005;
	wire new_net_8924;
	wire new_net_8818;
	wire new_net_7806;
	wire new_net_10340;
	wire new_net_8346;
	wire new_net_444;
	wire new_net_1993;
	wire new_net_1156;
	wire new_net_2531;
	wire new_net_3721;
	wire new_net_4358;
	wire new_net_4950;
	wire new_net_5941;
	wire new_net_5481;
	wire new_net_5965;
	wire new_net_480;
	wire new_net_5984;
	wire new_net_6321;
	wire new_net_8828;
	wire new_net_8363;
	wire new_net_9348;
	wire new_net_4497;
	wire new_net_8362;
	wire new_net_1943;
	wire n_0862_;
	wire n_0358_;
	wire n_1366_;
	wire new_net_1337;
	wire new_net_1568;
	wire new_net_1829;
	wire new_net_250;
	wire new_net_3112;
	wire new_net_4051;
	wire new_net_6559;
	wire new_net_6552;
	wire new_net_8968;
	wire new_net_5024;
	wire new_net_5022;
	wire new_net_7475;
	wire new_net_3353;
	wire new_net_59;
	wire new_net_890;
	wire new_net_1305;
	wire new_net_1452;
	wire new_net_2483;
	wire new_net_2378;
	wire new_net_2210;
	wire new_net_4222;
	wire new_net_4245;
	wire new_net_4311;
	wire new_net_8454;
	wire new_net_9684;
	wire new_net_8648;
	wire new_net_8239;
	wire new_net_9500;
	wire new_net_7945;
	wire new_net_9846;
	wire n_0863_;
	wire n_0359_;
	wire new_net_3375;
	wire n_1367_;
	wire new_net_291;
	wire new_net_1189;
	wire new_net_324;
	wire new_net_1039;
	wire new_net_3680;
	wire new_net_5673;
	wire new_net_10058;
	wire new_net_10646;
	wire new_net_9309;
	wire new_net_6595;
	wire new_net_9582;
	wire new_net_7465;
	wire new_net_10377;
	wire new_net_2067;
	wire new_net_445;
	wire new_net_628;
	wire new_net_1157;
	wire new_net_2594;
	wire new_net_4720;
	wire new_net_5985;
	wire new_net_7577;
	wire new_net_7601;
	wire new_net_8671;
	wire new_net_5059;
	wire new_net_7595;
	wire new_net_5838;
	wire new_net_8708;
	wire new_net_9054;
	wire new_net_9872;
	wire new_net_10472;
	wire new_net_9246;
	wire new_net_8152;
	wire new_net_1944;
	wire n_0864_;
	wire n_0360_;
	wire n_1368_;
	wire new_net_1569;
	wire new_net_2665;
	wire new_net_251;
	wire new_net_4571;
	wire new_net_5227;
	wire new_net_5774;
	wire new_net_8032;
	wire new_net_7738;
	wire new_net_10271;
	wire new_net_7248;
	wire new_net_7911;
	wire new_net_3701;
	wire new_net_4408;
	wire new_net_6462;
	wire new_net_9071;
	wire new_net_1453;
	wire new_net_1684;
	wire new_net_2755;
	wire new_net_60;
	wire new_net_2174;
	wire new_net_891;
	wire new_net_2284;
	wire new_net_2347;
	wire new_net_3242;
	wire new_net_3745;
	wire new_net_8618;
	wire new_net_5200;
	wire new_net_8701;
	wire new_net_7966;
	wire new_net_9867;
	wire new_net_9191;
	wire new_net_6896;
	wire new_net_325;
	wire new_net_1040;
	wire n_0361_;
	wire n_0865_;
	wire n_1369_;
	wire new_net_292;
	wire new_net_1190;
	wire new_net_3722;
	wire new_net_4941;
	wire new_net_5942;
	wire new_net_8649;
	wire new_net_8745;
	wire new_net_10083;
	wire n_0408_;
	wire new_net_9339;
	wire new_net_9213;
	wire new_net_6024;
	wire new_net_2929;
	wire new_net_3113;
	wire new_net_629;
	wire new_net_1338;
	wire new_net_1830;
	wire new_net_4052;
	wire new_net_4696;
	wire new_net_4738;
	wire new_net_4802;
	wire new_net_4826;
	wire new_net_7212;
	wire new_net_4297;
	wire new_net_4338;
	wire new_net_6806;
	wire n_0866_;
	wire n_0362_;
	wire new_net_3354;
	wire new_net_1306;
	wire n_1370_;
	wire new_net_252;
	wire new_net_4223;
	wire new_net_4246;
	wire new_net_4550;
	wire new_net_4768;
	wire new_net_6936;
	wire new_net_7346;
	wire new_net_10141;
	wire new_net_7515;
	wire new_net_7027;
	wire new_net_10235;
	wire new_net_5508;
	wire new_net_8639;
	wire new_net_6615;
	wire new_net_7936;
	wire new_net_1685;
	wire new_net_2211;
	wire new_net_2484;
	wire new_net_892;
	wire new_net_3376;
	wire new_net_2379;
	wire new_net_3681;
	wire new_net_6223;
	wire new_net_6247;
	wire new_net_9125;
	wire new_net_10049;
	wire new_net_10206;
	wire new_net_8664;
	wire new_net_326;
	wire new_net_2595;
	wire new_net_2930;
	wire n_0867_;
	wire n_0363_;
	wire n_1371_;
	wire new_net_446;
	wire new_net_1158;
	wire new_net_4166;
	wire new_net_4697;
	wire new_net_7387;
	wire new_net_10228;
	wire new_net_9232;
	wire new_net_10463;
	wire new_net_10385;
	wire new_net_1339;
	wire new_net_1570;
	wire new_net_1831;
	wire new_net_1945;
	wire new_net_2666;
	wire new_net_4572;
	wire new_net_5228;
	wire new_net_5775;
	wire new_net_6440;
	wire new_net_7060;
	wire new_net_7729;
	wire new_net_8380;
	wire new_net_10111;
	wire n_0964_;
	wire new_net_6347;
	wire new_net_4107;
	wire new_net_8192;
	wire new_net_8433;
	wire new_net_10513;
	wire new_net_7285;
	wire new_net_253;
	wire new_net_3243;
	wire n_0868_;
	wire new_net_1454;
	wire new_net_2756;
	wire new_net_61;
	wire n_0364_;
	wire new_net_1307;
	wire new_net_413;
	wire new_net_3746;
	wire new_net_8800;
	wire new_net_10324;
	wire new_net_3847;
	wire new_net_4743;
	wire new_net_9114;
	wire new_net_7837;
	wire new_net_293;
	wire new_net_1041;
	wire new_net_1191;
	wire new_net_2533;
	wire new_net_2285;
	wire new_net_3396;
	wire new_net_2348;
	wire new_net_3723;
	wire new_net_5943;
	wire new_net_5967;
	wire new_net_7426;
	wire new_net_8736;
	wire new_net_8885;
	wire new_net_8883;
	wire new_net_9158;
	wire new_net_9713;
	wire new_net_8344;
	wire new_net_9325;
	wire new_net_9131;
	wire new_net_1159;
	wire n_0869_;
	wire n_0365_;
	wire new_net_3114;
	wire new_net_447;
	wire new_net_4053;
	wire new_net_4739;
	wire new_net_4803;
	wire new_net_4827;
	wire new_net_5632;
	wire new_net_10635;
	wire new_net_10668;
	wire new_net_4912;
	wire new_net_7660;
	wire new_net_9072;
	wire new_net_9818;
	wire new_net_5001;
	wire new_net_4288;
	wire new_net_1571;
	wire new_net_1946;
	wire new_net_4224;
	wire new_net_4247;
	wire new_net_4286;
	wire new_net_4551;
	wire new_net_4690;
	wire new_net_4769;
	wire new_net_4962;
	wire new_net_5505;
	wire new_net_8248;
	wire new_net_8808;
	wire new_net_10417;
	wire new_net_7506;
	wire new_net_8447;
	wire new_net_8625;
	wire new_net_254;
	wire n_0366_;
	wire n_0870_;
	wire new_net_1455;
	wire new_net_62;
	wire new_net_3377;
	wire new_net_893;
	wire new_net_3682;
	wire new_net_5555;
	wire new_net_6224;
	wire new_net_9016;
	wire new_net_9286;
	wire new_net_8674;
	wire new_net_10197;
	wire new_net_5402;
	wire new_net_10354;
	wire new_net_10596;
	wire new_net_10594;
	wire new_net_8237;
	wire new_net_2380;
	wire new_net_294;
	wire new_net_327;
	wire new_net_1042;
	wire new_net_1192;
	wire new_net_2212;
	wire new_net_2485;
	wire new_net_2596;
	wire new_net_2931;
	wire new_net_4698;
	wire new_net_5858;
	wire new_net_8763;
	wire new_net_5815;
	wire new_net_6419;
	wire new_net_7378;
	wire new_net_8690;
	wire new_net_9038;
	wire new_net_10219;
	wire new_net_9470;
	wire new_net_5912;
	wire new_net_1832;
	wire n_0367_;
	wire n_0871_;
	wire new_net_631;
	wire new_net_1340;
	wire new_net_2667;
	wire new_net_4573;
	wire new_net_5229;
	wire new_net_5776;
	wire new_net_6441;
	wire new_net_8009;
	wire new_net_6338;
	wire new_net_8183;
	wire new_net_3960;
	wire new_net_7770;
	wire new_net_8419;
	wire new_net_6617;
	wire new_net_9838;
	wire new_net_2002;
	wire new_net_3244;
	wire new_net_1308;
	wire new_net_2757;
	wire new_net_3747;
	wire new_net_4008;
	wire new_net_4032;
	wire new_net_4185;
	wire new_net_4310;
	wire new_net_4587;
	wire new_net_8756;
	wire new_net_6093;
	wire new_net_8390;
	wire new_net_10560;
	wire new_net_10164;
	wire new_net_8316;
	wire new_net_4737;
	wire new_net_9105;
	wire new_net_7828;
	wire new_net_7045;
	wire new_net_2030;
	wire new_net_255;
	wire n_0368_;
	wire n_0872_;
	wire new_net_1456;
	wire new_net_1687;
	wire new_net_894;
	wire new_net_3724;
	wire new_net_3756;
	wire new_net_5406;
	wire new_net_5322;
	wire new_net_4974;
	wire new_net_6522;
	wire new_net_2349;
	wire new_net_328;
	wire new_net_448;
	wire new_net_1043;
	wire new_net_1160;
	wire new_net_3115;
	wire new_net_2286;
	wire new_net_4054;
	wire new_net_4740;
	wire new_net_4804;
	wire new_net_9917;
	wire new_net_10626;
	wire new_net_9915;
	wire new_net_3778;
	wire new_net_10437;
	wire new_net_1341;
	wire new_net_1572;
	wire new_net_1833;
	wire n_0369_;
	wire n_0873_;
	wire new_net_1947;
	wire new_net_2580;
	wire new_net_3397;
	wire new_net_4225;
	wire new_net_4248;
	wire new_net_6209;
	wire new_net_9139;
	wire new_net_2029;
	wire new_net_63;
	wire new_net_3378;
	wire new_net_1309;
	wire new_net_3683;
	wire new_net_6225;
	wire new_net_6249;
	wire new_net_9007;
	wire new_net_9323;
	wire new_net_9347;
	wire new_net_10183;
	wire new_net_9517;
	wire new_net_5386;
	wire n_0370_;
	wire n_0874_;
	wire new_net_256;
	wire new_net_295;
	wire new_net_1193;
	wire new_net_2597;
	wire new_net_2932;
	wire new_net_895;
	wire new_net_4691;
	wire new_net_4699;
	wire new_net_7858;
	wire new_net_10010;
	wire new_net_7364;
	wire new_net_7619;
	wire new_net_8480;
	wire new_net_4926;
	wire new_net_5903;
	wire new_net_8478;
	wire new_net_2668;
	wire new_net_2381;
	wire new_net_449;
	wire new_net_632;
	wire new_net_1161;
	wire new_net_2213;
	wire new_net_2486;
	wire new_net_4574;
	wire new_net_5230;
	wire new_net_5777;
	wire new_net_7300;
	wire new_net_8000;
	wire new_net_8662;
	wire new_net_8264;
	wire new_net_8169;
	wire new_net_10070;
	wire new_net_8410;
	wire new_net_4546;
	wire n_1210_;
	wire new_net_6380;
	wire new_net_7272;
	wire new_net_4432;
	wire new_net_9758;
	wire new_net_1573;
	wire n_0875_;
	wire n_0371_;
	wire new_net_3245;
	wire new_net_2758;
	wire new_net_1948;
	wire new_net_3748;
	wire new_net_4009;
	wire new_net_4033;
	wire new_net_4186;
	wire new_net_4595;
	wire new_net_8103;
	wire new_net_10546;
	wire new_net_5730;
	wire new_net_10155;
	wire new_net_6866;
	wire new_net_4567;
	wire new_net_5770;
	wire new_net_6133;
	wire new_net_64;
	wire new_net_1457;
	wire new_net_1688;
	wire new_net_2535;
	wire new_net_3725;
	wire new_net_5945;
	wire new_net_5969;
	wire new_net_6122;
	wire new_net_6524;
	wire new_net_7435;
	wire new_net_8867;
	wire new_net_7122;
	wire new_net_4368;
	wire new_net_7092;
	wire new_net_8212;
	wire new_net_10102;
	wire new_net_7175;
	wire new_net_3116;
	wire n_0372_;
	wire n_0876_;
	wire new_net_257;
	wire new_net_296;
	wire new_net_1194;
	wire new_net_329;
	wire new_net_1044;
	wire new_net_2084;
	wire new_net_4055;
	wire new_net_5966;
	wire new_net_7693;
	wire new_net_8978;
	wire new_net_2287;
	wire new_net_3398;
	wire new_net_2350;
	wire new_net_450;
	wire new_net_633;
	wire new_net_1834;
	wire new_net_4226;
	wire new_net_4249;
	wire new_net_4553;
	wire new_net_4589;
	wire new_net_7485;
	wire new_net_10119;
	wire new_net_6176;
	wire new_net_8906;
	wire new_net_8272;
	wire new_net_8904;
	wire new_net_7786;
	wire new_net_9694;
	wire new_net_3379;
	wire new_net_1310;
	wire new_net_1574;
	wire n_0373_;
	wire n_0877_;
	wire new_net_1949;
	wire new_net_4287;
	wire new_net_5532;
	wire new_net_6226;
	wire new_net_6250;
	wire new_net_9263;
	wire new_net_7960;
	wire new_net_9788;
	wire new_net_9597;
	wire new_net_4753;
	wire new_net_5377;
	wire new_net_5418;
	wire new_net_6039;
	wire new_net_8848;
	wire new_net_65;
	wire new_net_896;
	wire new_net_1458;
	wire new_net_1689;
	wire new_net_2933;
	wire new_net_2179;
	wire new_net_2181;
	wire new_net_2598;
	wire new_net_4692;
	wire new_net_4700;
	wire new_net_7849;
	wire new_net_9403;
	wire new_net_10001;
	wire new_net_3820;
	wire new_net_5263;
	wire new_net_8795;
	wire new_net_9727;
	wire new_net_5889;
	wire new_net_3878;
	wire new_net_2669;
	wire n_0374_;
	wire n_0878_;
	wire new_net_258;
	wire new_net_1162;
	wire new_net_1195;
	wire new_net_330;
	wire new_net_1045;
	wire new_net_4575;
	wire new_net_5231;
	wire new_net_3656;
	wire new_net_8042;
	wire new_net_9940;
	wire new_net_10281;
	wire new_net_4537;
	wire new_net_6366;
	wire new_net_7753;
	wire new_net_9938;
	wire new_net_10488;
	wire new_net_8575;
	wire new_net_4423;
	wire new_net_8573;
	wire new_net_451;
	wire new_net_634;
	wire new_net_1343;
	wire new_net_1835;
	wire new_net_2382;
	wire new_net_3246;
	wire new_net_2214;
	wire new_net_2487;
	wire new_net_2759;
	wire new_net_3355;
	wire new_net_8094;
	wire new_net_9553;
	wire new_net_10537;
	wire new_net_8925;
	wire new_net_8819;
	wire new_net_7807;
	wire new_net_10341;
	wire new_net_6124;
	wire new_net_9960;
	wire new_net_1950;
	wire new_net_1311;
	wire n_0879_;
	wire n_0375_;
	wire new_net_3726;
	wire new_net_5946;
	wire new_net_5970;
	wire new_net_6123;
	wire new_net_6525;
	wire new_net_7436;
	wire new_net_4951;
	wire new_net_8388;
	wire new_net_6324;
	wire new_net_6322;
	wire new_net_8829;
	wire new_net_8364;
	wire new_net_66;
	wire new_net_1989;
	wire new_net_297;
	wire new_net_897;
	wire new_net_1459;
	wire new_net_4056;
	wire new_net_4806;
	wire new_net_4830;
	wire new_net_5635;
	wire new_net_4498;
	wire new_net_9349;
	wire new_net_5952;
	wire new_net_7217;
	wire new_net_8770;
	wire new_net_8969;
	wire new_net_5025;
	wire new_net_3399;
	wire n_0880_;
	wire n_0376_;
	wire new_net_2913;
	wire new_net_259;
	wire new_net_1163;
	wire new_net_331;
	wire new_net_1046;
	wire new_net_4227;
	wire new_net_4250;
	wire new_net_6816;
	wire new_net_4312;
	wire new_net_7476;
	wire new_net_9685;
	wire new_net_3356;
	wire new_net_2288;
	wire new_net_3380;
	wire new_net_1344;
	wire new_net_1575;
	wire new_net_2351;
	wire new_net_5042;
	wire new_net_5676;
	wire new_net_6227;
	wire new_net_6236;
	wire new_net_6913;
	wire new_net_7946;
	wire new_net_9501;
	wire new_net_9847;
	wire new_net_4450;
	wire new_net_5674;
	wire new_net_10059;
	wire new_net_9075;
	wire new_net_10647;
	wire new_net_9310;
	wire new_net_9583;
	wire new_net_6596;
	wire new_net_7466;
	wire new_net_9394;
	wire new_net_1690;
	wire new_net_2599;
	wire n_0377_;
	wire n_0881_;
	wire new_net_2934;
	wire new_net_4701;
	wire new_net_4725;
	wire new_net_5990;
	wire new_net_7582;
	wire new_net_7606;
	wire new_net_6081;
	wire new_net_5060;
	wire new_net_7596;
	wire new_net_5839;
	wire new_net_8709;
	wire new_net_9055;
	wire new_net_298;
	wire new_net_898;
	wire new_net_1196;
	wire new_net_2031;
	wire new_net_2670;
	wire new_net_4576;
	wire new_net_4741;
	wire new_net_5232;
	wire new_net_5779;
	wire new_net_6625;
	wire new_net_8153;
	wire new_net_8033;
	wire new_net_7739;
	wire new_net_10272;
	wire new_net_7249;
	wire new_net_7912;
	wire new_net_3984;
	wire new_net_6463;
	wire new_net_332;
	wire new_net_1047;
	wire new_net_2760;
	wire new_net_635;
	wire n_0378_;
	wire new_net_452;
	wire n_0882_;
	wire new_net_1836;
	wire new_net_610;
	wire new_net_260;
	wire new_net_5707;
	wire new_net_8286;
	wire new_net_9544;
	wire new_net_8619;
	wire new_net_7798;
	wire new_net_7974;
	wire new_net_7967;
	wire new_net_9868;
	wire new_net_9192;
	wire new_net_2215;
	wire new_net_2488;
	wire new_net_2537;
	wire new_net_1312;
	wire new_net_1345;
	wire new_net_1576;
	wire new_net_1951;
	wire new_net_2383;
	wire new_net_3713;
	wire new_net_3727;
	wire new_net_10084;
	wire new_net_2919;
	wire new_net_1691;
	wire new_net_67;
	wire n_0883_;
	wire n_0379_;
	wire new_net_4057;
	wire new_net_4200;
	wire new_net_4807;
	wire new_net_4831;
	wire new_net_5636;
	wire new_net_7988;
	wire new_net_9214;
	wire new_net_7213;
	wire new_net_899;
	wire new_net_1164;
	wire new_net_1197;
	wire new_net_3400;
	wire new_net_4228;
	wire new_net_4251;
	wire new_net_4298;
	wire new_net_4555;
	wire new_net_4591;
	wire new_net_4966;
	wire n_0208_;
	wire new_net_4215;
	wire new_net_6937;
	wire new_net_10142;
	wire new_net_7516;
	wire new_net_10304;
	wire new_net_4871;
	wire new_net_5212;
	wire new_net_7028;
	wire new_net_5509;
	wire new_net_10236;
	wire new_net_8640;
	wire new_net_333;
	wire new_net_1048;
	wire new_net_3357;
	wire n_0884_;
	wire n_0380_;
	wire new_net_636;
	wire new_net_3381;
	wire new_net_453;
	wire new_net_1837;
	wire new_net_261;
	wire new_net_7937;
	wire new_net_10050;
	wire n_0551_;
	wire new_net_10207;
	wire new_net_2914;
	wire new_net_2600;
	wire new_net_2935;
	wire new_net_1952;
	wire new_net_1313;
	wire new_net_2289;
	wire new_net_2352;
	wire new_net_4034;
	wire new_net_4702;
	wire new_net_5991;
	wire new_net_10253;
	wire new_net_4167;
	wire new_net_7877;
	wire new_net_5825;
	wire new_net_5245;
	wire new_net_7388;
	wire new_net_9233;
	wire new_net_9480;
	wire new_net_299;
	wire new_net_1461;
	wire new_net_3117;
	wire new_net_68;
	wire n_0885_;
	wire n_0381_;
	wire new_net_2671;
	wire new_net_4577;
	wire new_net_5233;
	wire new_net_5780;
	wire new_net_10386;
	wire new_net_10270;
	wire new_net_6348;
	wire new_net_9529;
	wire new_net_8193;
	wire new_net_6449;
	wire new_net_8434;
	wire new_net_3248;
	wire new_net_2761;
	wire new_net_900;
	wire new_net_1165;
	wire new_net_1198;
	wire new_net_3751;
	wire new_net_4012;
	wire new_net_4189;
	wire new_net_4290;
	wire new_net_4772;
	wire new_net_8605;
	wire new_net_8801;
	wire new_net_10325;
	wire new_net_4612;
	wire new_net_4744;
	wire new_net_9859;
	wire new_net_9115;
	wire new_net_262;
	wire new_net_334;
	wire new_net_1049;
	wire n_0886_;
	wire n_0382_;
	wire new_net_454;
	wire new_net_1838;
	wire new_net_3728;
	wire new_net_5794;
	wire new_net_5948;
	wire new_net_7055;
	wire new_net_7838;
	wire new_net_7427;
	wire new_net_8737;
	wire new_net_10258;
	wire new_net_9161;
	wire new_net_4721;
	wire new_net_8884;
	wire new_net_9159;
	wire new_net_7146;
	wire new_net_9714;
	wire new_net_8345;
	wire new_net_9326;
	wire new_net_2100;
	wire new_net_2216;
	wire new_net_1578;
	wire new_net_1692;
	wire new_net_2384;
	wire new_net_4035;
	wire new_net_4058;
	wire new_net_4808;
	wire new_net_4832;
	wire new_net_5637;
	wire new_net_10671;
	wire new_net_6537;
	wire new_net_10636;
	wire n_0273_;
	wire new_net_7661;
	wire new_net_9819;
	wire new_net_8767;
	wire new_net_4651;
	wire new_net_2001;
	wire new_net_300;
	wire new_net_1462;
	wire new_net_3118;
	wire n_0383_;
	wire new_net_3401;
	wire n_0887_;
	wire new_net_4229;
	wire new_net_4252;
	wire new_net_4289;
	wire new_net_8249;
	wire new_net_4089;
	wire new_net_6470;
	wire new_net_3995;
	wire new_net_7507;
	wire new_net_8448;
	wire new_net_8626;
	wire new_net_637;
	wire new_net_1199;
	wire new_net_3358;
	wire new_net_3382;
	wire new_net_3686;
	wire new_net_6229;
	wire new_net_6253;
	wire new_net_6444;
	wire new_net_9327;
	wire new_net_9351;
	wire new_net_5556;
	wire new_net_9287;
	wire new_net_10198;
	wire new_net_10355;
	wire new_net_10597;
	wire new_net_7116;
	wire new_net_263;
	wire new_net_2915;
	wire new_net_335;
	wire new_net_1050;
	wire new_net_2601;
	wire new_net_2936;
	wire n_0888_;
	wire n_0384_;
	wire new_net_1953;
	wire new_net_1314;
	wire new_net_5442;
	wire new_net_8238;
	wire new_net_8764;
	wire new_net_9039;
	wire new_net_6717;
	wire new_net_7379;
	wire new_net_8691;
	wire new_net_10220;
	wire new_net_1693;
	wire new_net_69;
	wire new_net_2290;
	wire new_net_2353;
	wire new_net_2672;
	wire new_net_4313;
	wire new_net_4578;
	wire new_net_5234;
	wire new_net_5781;
	wire new_net_5913;
	wire new_net_3902;
	wire new_net_8184;
	wire new_net_8064;
	wire new_net_7771;
	wire new_net_8420;
	wire new_net_1166;
	wire new_net_3249;
	wire n_0889_;
	wire n_0385_;
	wire new_net_1463;
	wire new_net_2762;
	wire new_net_901;
	wire new_net_3752;
	wire new_net_4013;
	wire new_net_4190;
	wire new_net_6268;
	wire new_net_6616;
	wire new_net_9839;
	wire new_net_10165;
	wire new_net_8317;
	wire new_net_9106;
	wire new_net_1839;
	wire new_net_638;
	wire new_net_2180;
	wire new_net_2491;
	wire new_net_2539;
	wire new_net_3729;
	wire new_net_5949;
	wire new_net_6126;
	wire new_net_6528;
	wire new_net_7046;
	wire new_net_9621;
	wire new_net_8809;
	wire new_net_5323;
	wire new_net_4975;
	wire new_net_1348;
	wire new_net_1579;
	wire new_net_264;
	wire n_0890_;
	wire n_0386_;
	wire new_net_1954;
	wire new_net_1315;
	wire new_net_4059;
	wire new_net_4314;
	wire new_net_4809;
	wire new_net_6002;
	wire new_net_6523;
	wire new_net_10627;
	wire new_net_3779;
	wire new_net_9916;
	wire new_net_10438;
	wire new_net_2385;
	wire new_net_70;
	wire new_net_301;
	wire new_net_2217;
	wire new_net_3119;
	wire new_net_3402;
	wire new_net_4230;
	wire new_net_4253;
	wire new_net_4557;
	wire new_net_4593;
	wire new_net_5043;
	wire new_net_6914;
	wire new_net_6637;
	wire new_net_9008;
	wire new_net_10184;
	wire new_net_9518;
	wire new_net_4629;
	wire new_net_5387;
	wire new_net_3023;
	wire new_net_1992;
	wire n_0933_;
	wire n_0135_;
	wire n_0429_;
	wire n_1143_;
	wire new_net_3326;
	wire n_0639_;
	wire new_net_3652;
	wire new_net_3699;
	wire new_net_7365;
	wire new_net_8393;
	wire new_net_4492;
	wire new_net_7620;
	wire new_net_8481;
	wire new_net_7709;
	wire new_net_8001;
	wire new_net_8663;
	wire new_net_3605;
	wire new_net_4782;
	wire new_net_7471;
	wire new_net_7621;
	wire new_net_8054;
	wire new_net_7301;
	wire new_net_8076;
	wire new_net_9689;
	wire new_net_10055;
	wire new_net_9082;
	wire new_net_5354;
	wire new_net_10071;
	wire new_net_8411;
	wire new_net_7273;
	wire new_net_9759;
	wire new_net_9126;
	wire new_net_8104;
	wire new_net_919;
	wire new_net_2847;
	wire new_net_202;
	wire new_net_3218;
	wire n_0934_;
	wire n_0136_;
	wire n_0430_;
	wire n_1144_;
	wire new_net_352;
	wire n_0640_;
	wire new_net_3166;
	wire new_net_5731;
	wire new_net_10547;
	wire new_net_10156;
	wire new_net_5724;
	wire new_net_6867;
	wire new_net_9975;
	wire new_net_2312;
	wire new_net_1596;
	wire new_net_3067;
	wire new_net_656;
	wire new_net_806;
	wire new_net_3091;
	wire new_net_3262;
	wire new_net_1710;
	wire new_net_2249;
	wire new_net_3840;
	wire new_net_8868;
	wire new_net_7093;
	wire new_net_6514;
	wire new_net_7176;
	wire new_net_10378;
	wire n_0431_;
	wire new_net_3046;
	wire n_0641_;
	wire n_0935_;
	wire n_0137_;
	wire n_1145_;
	wire new_net_6541;
	wire new_net_7452;
	wire new_net_8817;
	wire new_net_9010;
	wire new_net_3770;
	wire new_net_7694;
	wire new_net_9605;
	wire new_net_10360;
	wire n_0830_;
	wire new_net_8856;
	wire new_net_10120;
	wire new_net_3606;
	wire new_net_22;
	wire n_0560_;
	wire new_net_4451;
	wire new_net_5397;
	wire new_net_5421;
	wire new_net_5675;
	wire new_net_6177;
	wire new_net_6688;
	wire new_net_7350;
	wire new_net_5180;
	wire new_net_8907;
	wire new_net_5696;
	wire new_net_8273;
	wire new_net_8905;
	wire new_net_5533;
	wire new_net_9264;
	wire n_0642_;
	wire new_net_389;
	wire n_0432_;
	wire new_net_920;
	wire new_net_203;
	wire n_0138_;
	wire n_0936_;
	wire new_net_509;
	wire new_net_1857;
	wire new_net_2888;
	wire new_net_7961;
	wire new_net_9789;
	wire new_net_4754;
	wire new_net_5378;
	wire new_net_5419;
	wire new_net_6040;
	wire new_net_9404;
	wire new_net_10104;
	wire new_net_7850;
	wire new_net_3024;
	wire new_net_1597;
	wire new_net_657;
	wire new_net_1069;
	wire new_net_2449;
	wire new_net_2218;
	wire new_net_3277;
	wire new_net_3327;
	wire new_net_3653;
	wire new_net_3700;
	wire new_net_6701;
	wire new_net_8746;
	wire new_net_3821;
	wire new_net_4833;
	wire new_net_7901;
	wire new_net_9728;
	wire new_net_5849;
	wire new_net_5890;
	wire new_net_10243;
	wire n_0643_;
	wire n_0433_;
	wire n_1147_;
	wire n_0139_;
	wire n_0937_;
	wire new_net_4783;
	wire new_net_7287;
	wire new_net_6210;
	wire new_net_7622;
	wire new_net_8055;
	wire new_net_9941;
	wire new_net_10282;
	wire n_1034_;
	wire new_net_4538;
	wire new_net_6367;
	wire new_net_9939;
	wire new_net_8576;
	wire new_net_6198;
	wire new_net_4045;
	wire new_net_10028;
	wire new_net_8095;
	wire new_net_1482;
	wire new_net_3475;
	wire new_net_2848;
	wire new_net_1969;
	wire new_net_3219;
	wire new_net_23;
	wire new_net_353;
	wire new_net_2126;
	wire new_net_3956;
	wire new_net_4143;
	wire new_net_8926;
	wire new_net_9554;
	wire new_net_8820;
	wire new_net_7808;
	wire new_net_10342;
	wire new_net_3866;
	wire new_net_6125;
	wire new_net_9961;
	wire new_net_6269;
	wire new_net_1711;
	wire n_0644_;
	wire new_net_390;
	wire new_net_3263;
	wire new_net_921;
	wire new_net_3092;
	wire n_0140_;
	wire n_0434_;
	wire n_1148_;
	wire new_net_204;
	wire new_net_4952;
	wire new_net_7079;
	wire new_net_5483;
	wire new_net_8389;
	wire new_net_6325;
	wire new_net_8948;
	wire new_net_5986;
	wire new_net_5080;
	wire new_net_6323;
	wire new_net_8830;
	wire new_net_9352;
	wire new_net_10606;
	wire new_net_8365;
	wire new_net_9350;
	wire new_net_2313;
	wire new_net_658;
	wire new_net_1070;
	wire new_net_1598;
	wire new_net_2250;
	wire new_net_3047;
	wire new_net_6542;
	wire new_net_7453;
	wire new_net_9011;
	wire new_net_9479;
	wire new_net_8970;
	wire new_net_10229;
	wire new_net_6819;
	wire new_net_7477;
	wire n_1149_;
	wire new_net_2060;
	wire n_0435_;
	wire n_0645_;
	wire n_0939_;
	wire n_0141_;
	wire new_net_1970;
	wire new_net_3607;
	wire new_net_4265;
	wire new_net_4452;
	wire new_net_6494;
	wire new_net_9686;
	wire new_net_8650;
	wire new_net_9502;
	wire new_net_354;
	wire new_net_1483;
	wire new_net_2889;
	wire new_net_4385;
	wire new_net_4607;
	wire new_net_4844;
	wire new_net_5619;
	wire new_net_6340;
	wire new_net_7292;
	wire new_net_9848;
	wire new_net_9311;
	wire new_net_6597;
	wire new_net_9584;
	wire new_net_7467;
	wire new_net_9395;
	wire new_net_4894;
	wire new_net_808;
	wire n_1150_;
	wire new_net_1712;
	wire new_net_391;
	wire n_0436_;
	wire n_0646_;
	wire n_0940_;
	wire n_0142_;
	wire new_net_205;
	wire new_net_1859;
	wire new_net_8886;
	wire new_net_8710;
	wire n_0831_;
	wire new_net_10474;
	wire new_net_2219;
	wire new_net_2450;
	wire new_net_4266;
	wire new_net_4627;
	wire new_net_4784;
	wire new_net_4316;
	wire new_net_7623;
	wire new_net_7783;
	wire new_net_8078;
	wire new_net_8154;
	wire new_net_8391;
	wire new_net_3925;
	wire new_net_7740;
	wire new_net_10273;
	wire new_net_7250;
	wire new_net_7913;
	wire new_net_3703;
	wire new_net_4410;
	wire n_1151_;
	wire n_0647_;
	wire n_0437_;
	wire n_0143_;
	wire new_net_2849;
	wire new_net_3220;
	wire n_0941_;
	wire new_net_24;
	wire new_net_4144;
	wire new_net_4647;
	wire new_net_5708;
	wire new_net_8620;
	wire new_net_9545;
	wire new_net_7799;
	wire new_net_4624;
	wire new_net_7975;
	wire n_0072_;
	wire new_net_7968;
	wire new_net_9193;
	wire new_net_9869;
	wire new_net_5582;
	wire new_net_3264;
	wire new_net_511;
	wire new_net_922;
	wire new_net_1484;
	wire new_net_2586;
	wire new_net_3069;
	wire new_net_3842;
	wire new_net_3957;
	wire new_net_3981;
	wire new_net_4159;
	wire new_net_4943;
	wire new_net_6409;
	wire new_net_7437;
	wire new_net_10085;
	wire new_net_9630;
	wire new_net_9215;
	wire new_net_545;
	wire n_0648_;
	wire new_net_392;
	wire new_net_659;
	wire n_0438_;
	wire n_1152_;
	wire n_0144_;
	wire new_net_206;
	wire new_net_1599;
	wire new_net_3048;
	wire new_net_5944;
	wire new_net_6026;
	wire new_net_9422;
	wire new_net_10681;
	wire new_net_2251;
	wire new_net_2314;
	wire new_net_1072;
	wire new_net_3608;
	wire new_net_4299;
	wire new_net_4453;
	wire new_net_4648;
	wire new_net_5399;
	wire new_net_5423;
	wire new_net_5677;
	wire new_net_6938;
	wire new_net_10143;
	wire new_net_6427;
	wire new_net_7517;
	wire new_net_4010;
	wire new_net_5512;
	wire new_net_10305;
	wire new_net_7029;
	wire new_net_10237;
	wire new_net_5510;
	wire new_net_10011;
	wire new_net_8641;
	wire new_net_9488;
	wire new_net_2890;
	wire n_1153_;
	wire new_net_355;
	wire new_net_25;
	wire n_0649_;
	wire n_0943_;
	wire n_0439_;
	wire n_0145_;
	wire new_net_3910;
	wire new_net_4386;
	wire new_net_10051;
	wire new_net_9380;
	wire new_net_8757;
	wire new_net_6583;
	wire new_net_10208;
	wire new_net_1713;
	wire new_net_512;
	wire new_net_809;
	wire new_net_923;
	wire new_net_1485;
	wire new_net_3655;
	wire new_net_3702;
	wire new_net_3952;
	wire new_net_4409;
	wire new_net_5812;
	wire new_net_4168;
	wire new_net_7878;
	wire new_net_5826;
	wire new_net_5246;
	wire new_net_7389;
	wire new_net_9234;
	wire new_net_9481;
	wire new_net_10465;
	wire new_net_10387;
	wire new_net_546;
	wire n_1154_;
	wire n_0650_;
	wire n_0944_;
	wire n_0146_;
	wire n_0440_;
	wire new_net_660;
	wire new_net_207;
	wire new_net_1600;
	wire new_net_4267;
	wire new_net_9918;
	wire new_net_6351;
	wire new_net_6349;
	wire new_net_9530;
	wire new_net_4109;
	wire new_net_8194;
	wire new_net_6450;
	wire new_net_8435;
	wire new_net_10517;
	wire new_net_2451;
	wire new_net_2220;
	wire new_net_2850;
	wire new_net_3221;
	wire new_net_4145;
	wire new_net_5002;
	wire new_net_5026;
	wire new_net_5044;
	wire new_net_5250;
	wire new_net_5717;
	wire new_net_8606;
	wire new_net_9140;
	wire new_net_8802;
	wire new_net_10326;
	wire new_net_3850;
	wire new_net_4745;
	wire new_net_9860;
	wire new_net_9116;
	wire new_net_7839;
	wire new_net_2037;
	wire new_net_3070;
	wire n_0147_;
	wire new_net_26;
	wire new_net_3330;
	wire n_1155_;
	wire new_net_356;
	wire new_net_3265;
	wire n_0651_;
	wire n_0945_;
	wire n_0212_;
	wire new_net_9162;
	wire new_net_4722;
	wire new_net_9160;
	wire new_net_6390;
	wire n_0832_;
	wire new_net_3049;
	wire new_net_1861;
	wire new_net_3457;
	wire new_net_1714;
	wire new_net_393;
	wire new_net_513;
	wire new_net_810;
	wire new_net_6538;
	wire new_net_6544;
	wire new_net_7455;
	wire new_net_9133;
	wire new_net_9643;
	wire new_net_10637;
	wire new_net_10672;
	wire new_net_9820;
	wire new_net_5003;
	wire new_net_8768;
	wire new_net_6147;
	wire new_net_4652;
	wire new_net_208;
	wire new_net_3609;
	wire n_0946_;
	wire n_0148_;
	wire new_net_1073;
	wire n_0442_;
	wire n_1156_;
	wire n_0652_;
	wire new_net_4454;
	wire new_net_4649;
	wire new_net_6471;
	wire new_net_3996;
	wire new_net_8449;
	wire new_net_8627;
	wire new_net_8221;
	wire new_net_2891;
	wire new_net_3329;
	wire new_net_2252;
	wire new_net_2315;
	wire new_net_4387;
	wire new_net_4609;
	wire new_net_4846;
	wire new_net_6342;
	wire new_net_7294;
	wire new_net_9618;
	wire new_net_5557;
	wire new_net_9018;
	wire new_net_9288;
	wire new_net_10199;
	wire new_net_10356;
	wire new_net_7117;
	wire n_0947_;
	wire n_0149_;
	wire new_net_27;
	wire new_net_357;
	wire new_net_1486;
	wire n_0443_;
	wire n_1157_;
	wire n_0653_;
	wire new_net_924;
	wire new_net_3025;
	wire new_net_4767;
	wire new_net_5443;
	wire new_net_8765;
	wire new_net_5817;
	wire new_net_9040;
	wire new_net_8692;
	wire new_net_10498;
	wire new_net_10221;
	wire new_net_8491;
	wire new_net_9747;
	wire new_net_9472;
	wire new_net_1601;
	wire new_net_394;
	wire new_net_547;
	wire new_net_661;
	wire new_net_1862;
	wire new_net_4268;
	wire new_net_7625;
	wire new_net_7769;
	wire new_net_7785;
	wire new_net_8011;
	wire new_net_4394;
	wire new_net_6230;
	wire new_net_8185;
	wire new_net_8065;
	wire new_net_7772;
	wire new_net_8421;
	wire new_net_8979;
	wire new_net_6619;
	wire new_net_2851;
	wire new_net_209;
	wire new_net_3222;
	wire n_0150_;
	wire new_net_3476;
	wire new_net_1074;
	wire n_0654_;
	wire n_0948_;
	wire n_0444_;
	wire n_1158_;
	wire new_net_6095;
	wire new_net_10166;
	wire new_net_8318;
	wire new_net_10446;
	wire new_net_9107;
	wire new_net_9695;
	wire new_net_2452;
	wire new_net_3266;
	wire new_net_2221;
	wire new_net_3071;
	wire new_net_3844;
	wire new_net_3912;
	wire new_net_3959;
	wire new_net_3983;
	wire new_net_4161;
	wire new_net_6163;
	wire new_net_9622;
	wire new_net_5408;
	wire new_net_8810;
	wire new_net_5324;
	wire new_net_4976;
	wire new_net_6435;
	wire new_net_510;
	wire new_net_925;
	wire new_net_3026;
	wire new_net_3050;
	wire new_net_3458;
	wire n_0151_;
	wire new_net_811;
	wire n_0655_;
	wire n_0949_;
	wire n_1159_;
	wire new_net_1487;
	wire new_net_10628;
	wire n_1281_;
	wire new_net_542;
	wire new_net_1991;
	wire new_net_3610;
	wire new_net_548;
	wire new_net_662;
	wire new_net_1602;
	wire new_net_4455;
	wire new_net_4650;
	wire new_net_5401;
	wire new_net_5425;
	wire new_net_5679;
	wire new_net_6843;
	wire new_net_6915;
	wire new_net_10489;
	wire new_net_210;
	wire new_net_2892;
	wire n_0152_;
	wire n_0446_;
	wire n_1160_;
	wire n_0656_;
	wire n_0950_;
	wire new_net_1075;
	wire new_net_4388;
	wire new_net_4435;
	wire new_net_9009;
	wire new_net_6416;
	wire new_net_8256;
	wire new_net_10185;
	wire new_net_9519;
	wire new_net_10173;
	wire new_net_2316;
	wire new_net_28;
	wire new_net_358;
	wire new_net_2253;
	wire new_net_3657;
	wire new_net_3704;
	wire new_net_3342;
	wire new_net_4411;
	wire new_net_4433;
	wire new_net_5814;
	wire new_net_7860;
	wire new_net_5111;
	wire new_net_8482;
	wire new_net_4928;
	wire n_0951_;
	wire new_net_515;
	wire new_net_1863;
	wire n_0153_;
	wire new_net_812;
	wire n_0447_;
	wire n_1161_;
	wire n_0657_;
	wire new_net_1716;
	wire new_net_395;
	wire new_net_7710;
	wire new_net_8002;
	wire new_net_7302;
	wire new_net_8171;
	wire new_net_9666;
	wire new_net_8412;
	wire new_net_4548;
	wire new_net_7274;
	wire new_net_4140;
	wire new_net_2852;
	wire new_net_1603;
	wire new_net_3223;
	wire new_net_663;
	wire new_net_4147;
	wire new_net_5004;
	wire new_net_5028;
	wire new_net_5046;
	wire new_net_5252;
	wire new_net_5719;
	wire new_net_8105;
	wire new_net_4597;
	wire new_net_9127;
	wire new_net_6410;
	wire new_net_10548;
	wire new_net_5732;
	wire new_net_10157;
	wire n_0694_;
	wire new_net_6868;
	wire new_net_4569;
	wire new_net_5772;
	wire new_net_6135;
	wire new_net_211;
	wire new_net_3072;
	wire n_0154_;
	wire new_net_3267;
	wire n_0658_;
	wire n_0952_;
	wire n_0448_;
	wire n_1162_;
	wire new_net_1076;
	wire new_net_3845;
	wire new_net_8869;
	wire new_net_4372;
	wire new_net_10060;
	wire new_net_7124;
	wire new_net_4370;
	wire new_net_7094;
	wire new_net_2177;
	wire new_net_3027;
	wire new_net_3051;
	wire new_net_3459;
	wire new_net_2453;
	wire new_net_29;
	wire new_net_359;
	wire new_net_926;
	wire new_net_2222;
	wire new_net_1488;
	wire new_net_6515;
	wire new_net_7177;
	wire new_net_565;
	wire new_net_8258;
	wire new_net_7639;
	wire new_net_5968;
	wire new_net_7695;
	wire new_net_396;
	wire n_0449_;
	wire new_net_1995;
	wire new_net_1864;
	wire new_net_516;
	wire new_net_3611;
	wire n_0155_;
	wire new_net_549;
	wire n_0953_;
	wire n_0659_;
	wire new_net_7487;
	wire new_net_8857;
	wire new_net_10121;
	wire new_net_6178;
	wire new_net_5181;
	wire new_net_8908;
	wire new_net_1604;
	wire new_net_2893;
	wire new_net_3331;
	wire new_net_4389;
	wire new_net_4611;
	wire new_net_4848;
	wire new_net_5534;
	wire new_net_6344;
	wire new_net_6398;
	wire new_net_6417;
	wire new_net_9265;
	wire new_net_9790;
	wire new_net_4400;
	wire new_net_5422;
	wire new_net_4755;
	wire new_net_5379;
	wire new_net_5420;
	wire new_net_6041;
	wire new_net_1077;
	wire n_0660_;
	wire new_net_212;
	wire n_0156_;
	wire n_0450_;
	wire n_1164_;
	wire n_0954_;
	wire new_net_3477;
	wire new_net_3658;
	wire new_net_3705;
	wire new_net_9405;
	wire new_net_10003;
	wire new_net_8747;
	wire new_net_7902;
	wire new_net_3302;
	wire new_net_5265;
	wire new_net_9729;
	wire new_net_5850;
	wire new_net_5891;
	wire new_net_10244;
	wire new_net_1717;
	wire new_net_2254;
	wire new_net_2317;
	wire new_net_30;
	wire new_net_813;
	wire new_net_927;
	wire new_net_1489;
	wire new_net_7627;
	wire new_net_7787;
	wire new_net_8082;
	wire new_net_8044;
	wire new_net_9942;
	wire new_net_10283;
	wire new_net_4539;
	wire new_net_6368;
	wire new_net_8577;
	wire new_net_8214;
	wire n_0661_;
	wire new_net_397;
	wire new_net_664;
	wire new_net_2853;
	wire new_net_3224;
	wire n_0955_;
	wire n_0157_;
	wire n_0451_;
	wire n_1165_;
	wire new_net_550;
	wire new_net_6199;
	wire new_net_8096;
	wire new_net_10029;
	wire new_net_9555;
	wire new_net_10539;
	wire new_net_8927;
	wire new_net_4989;
	wire new_net_9444;
	wire new_net_7809;
	wire new_net_10343;
	wire new_net_9962;
	wire new_net_3268;
	wire new_net_3073;
	wire new_net_3914;
	wire new_net_3961;
	wire new_net_3985;
	wire new_net_4163;
	wire new_net_6165;
	wire new_net_6270;
	wire new_net_6418;
	wire new_net_6464;
	wire new_net_4953;
	wire new_net_7080;
	wire new_net_7078;
	wire new_net_6326;
	wire new_net_10561;
	wire new_net_8949;
	wire new_net_5987;
	wire new_net_8831;
	wire new_net_9353;
	wire new_net_10607;
	wire n_1166_;
	wire new_net_360;
	wire new_net_2098;
	wire n_0452_;
	wire new_net_3028;
	wire new_net_213;
	wire new_net_3052;
	wire new_net_3460;
	wire n_0662_;
	wire n_0956_;
	wire new_net_8366;
	wire new_net_4500;
	wire new_net_5954;
	wire new_net_7219;
	wire new_net_2802;
	wire new_net_8971;
	wire new_net_10230;
	wire n_0075_;
	wire new_net_2223;
	wire new_net_3612;
	wire new_net_517;
	wire new_net_814;
	wire new_net_928;
	wire new_net_1490;
	wire new_net_1718;
	wire new_net_1865;
	wire new_net_2454;
	wire new_net_4457;
	wire new_net_6820;
	wire new_net_7478;
	wire new_net_6818;
	wire new_net_4232;
	wire new_net_6948;
	wire new_net_6495;
	wire new_net_9687;
	wire new_net_3332;
	wire n_1167_;
	wire n_0663_;
	wire new_net_398;
	wire n_0453_;
	wire new_net_665;
	wire new_net_1605;
	wire n_0159_;
	wire n_0957_;
	wire new_net_2894;
	wire new_net_5678;
	wire new_net_8651;
	wire new_net_7948;
	wire new_net_9503;
	wire new_net_9849;
	wire new_net_9312;
	wire new_net_3849;
	wire new_net_6598;
	wire new_net_9585;
	wire new_net_1078;
	wire new_net_3478;
	wire new_net_3659;
	wire new_net_3706;
	wire new_net_4413;
	wire new_net_5816;
	wire new_net_5840;
	wire new_net_6735;
	wire new_net_6759;
	wire new_net_7468;
	wire new_net_9396;
	wire new_net_6083;
	wire new_net_8887;
	wire new_net_7399;
	wire new_net_5841;
	wire new_net_8711;
	wire new_net_8349;
	wire n_1168_;
	wire new_net_361;
	wire n_0664_;
	wire n_0454_;
	wire new_net_214;
	wire n_0160_;
	wire n_0958_;
	wire new_net_31;
	wire new_net_4630;
	wire new_net_7788;
	wire new_net_8515;
	wire new_net_10475;
	wire new_net_8155;
	wire new_net_8392;
	wire new_net_8035;
	wire new_net_7741;
	wire new_net_10274;
	wire new_net_7251;
	wire new_net_7914;
	wire new_net_2255;
	wire new_net_1491;
	wire new_net_2318;
	wire new_net_2854;
	wire new_net_3225;
	wire new_net_518;
	wire new_net_551;
	wire new_net_815;
	wire new_net_929;
	wire new_net_1866;
	wire new_net_3986;
	wire new_net_8288;
	wire new_net_5709;
	wire new_net_9546;
	wire new_net_235;
	wire new_net_7800;
	wire new_net_3455;
	wire new_net_7976;
	wire new_net_9870;
	wire new_net_9194;
	wire n_0665_;
	wire new_net_399;
	wire new_net_1606;
	wire n_0455_;
	wire n_1169_;
	wire n_0161_;
	wire n_0959_;
	wire new_net_3074;
	wire new_net_3915;
	wire new_net_3962;
	wire new_net_5294;
	wire new_net_5583;
	wire new_net_7440;
	wire new_net_8783;
	wire new_net_4944;
	wire new_net_7438;
	wire n_0974_;
	wire new_net_5223;
	wire new_net_276;
	wire new_net_10598;
	wire new_net_3029;
	wire new_net_3053;
	wire new_net_543;
	wire new_net_3461;
	wire new_net_6548;
	wire new_net_7411;
	wire new_net_7459;
	wire new_net_8821;
	wire new_net_8890;
	wire new_net_9017;
	wire new_net_9216;
	wire new_net_4202;
	wire new_net_9423;
	wire new_net_10682;
	wire new_net_32;
	wire n_1170_;
	wire new_net_362;
	wire new_net_1719;
	wire n_0666_;
	wire n_0456_;
	wire new_net_3613;
	wire n_0162_;
	wire new_net_215;
	wire n_0960_;
	wire new_net_4300;
	wire new_net_10002;
	wire new_net_4217;
	wire new_net_6939;
	wire new_net_8257;
	wire new_net_10144;
	wire new_net_7520;
	wire new_net_3247;
	wire new_net_4011;
	wire new_net_5513;
	wire new_net_9607;
	wire new_net_10306;
	wire new_net_4873;
	wire new_net_7030;
	wire new_net_5511;
	wire new_net_1867;
	wire new_net_2895;
	wire new_net_2455;
	wire new_net_2224;
	wire new_net_3333;
	wire new_net_552;
	wire new_net_666;
	wire new_net_4391;
	wire new_net_4613;
	wire new_net_4850;
	wire new_net_8642;
	wire new_net_9489;
	wire n_0565_;
	wire new_net_10052;
	wire new_net_10209;
	wire new_net_6584;
	wire new_net_485;
	wire new_net_3107;
	wire n_1171_;
	wire new_net_400;
	wire n_0457_;
	wire new_net_2096;
	wire n_0667_;
	wire n_0961_;
	wire n_0163_;
	wire new_net_3660;
	wire new_net_3707;
	wire new_net_6069;
	wire new_net_7879;
	wire new_net_5827;
	wire new_net_8702;
	wire n_0076_;
	wire new_net_3093;
	wire new_net_1080;
	wire new_net_4269;
	wire new_net_4631;
	wire new_net_7789;
	wire new_net_8060;
	wire new_net_8084;
	wire new_net_8243;
	wire new_net_9482;
	wire new_net_9604;
	wire new_net_10388;
	wire new_net_10466;
	wire new_net_9919;
	wire new_net_3917;
	wire new_net_6350;
	wire new_net_10439;
	wire new_net_8195;
	wire new_net_6451;
	wire new_net_4675;
	wire n_0962_;
	wire new_net_519;
	wire new_net_816;
	wire n_1172_;
	wire new_net_1492;
	wire new_net_1720;
	wire n_0668_;
	wire n_0458_;
	wire n_0164_;
	wire new_net_930;
	wire new_net_6960;
	wire new_net_8274;
	wire new_net_10518;
	wire new_net_8607;
	wire new_net_9141;
	wire new_net_1432;
	wire new_net_8803;
	wire new_net_10327;
	wire new_net_4614;
	wire new_net_9861;
	wire new_net_1607;
	wire new_net_2587;
	wire new_net_3075;
	wire new_net_2256;
	wire new_net_2319;
	wire new_net_667;
	wire new_net_3916;
	wire new_net_3963;
	wire new_net_317;
	wire new_net_3987;
	wire new_net_7840;
	wire new_net_5796;
	wire new_net_7057;
	wire new_net_566;
	wire new_net_3489;
	wire new_net_9163;
	wire new_net_4723;
	wire new_net_7148;
	wire new_net_9716;
	wire n_0963_;
	wire new_net_3462;
	wire new_net_3094;
	wire n_0669_;
	wire new_net_401;
	wire n_0459_;
	wire n_1173_;
	wire n_0165_;
	wire new_net_3030;
	wire new_net_4436;
	wire new_net_8218;
	wire new_net_10673;
	wire new_net_6539;
	wire new_net_10012;
	wire new_net_10638;
	wire n_0280_;
	wire new_net_2779;
	wire new_net_7663;
	wire new_net_7360;
	wire new_net_3614;
	wire new_net_33;
	wire new_net_363;
	wire new_net_4459;
	wire new_net_4653;
	wire new_net_4654;
	wire new_net_4677;
	wire new_net_5405;
	wire new_net_5429;
	wire new_net_6148;
	wire new_net_4291;
	wire new_net_8667;
	wire new_net_10420;
	wire new_net_6472;
	wire new_net_3997;
	wire new_net_5201;
	wire new_net_8628;
	wire new_net_3334;
	wire n_1174_;
	wire new_net_817;
	wire new_net_520;
	wire new_net_1868;
	wire new_net_2896;
	wire new_net_217;
	wire new_net_553;
	wire new_net_931;
	wire new_net_1493;
	wire new_net_5558;
	wire new_net_9019;
	wire new_net_9289;
	wire n_0000_;
	wire new_net_10357;
	wire new_net_2456;
	wire new_net_2225;
	wire new_net_2178;
	wire new_net_668;
	wire new_net_1608;
	wire new_net_3661;
	wire new_net_3708;
	wire new_net_4415;
	wire new_net_5818;
	wire new_net_5842;
	wire new_net_5444;
	wire new_net_9041;
	wire new_net_6719;
	wire new_net_7381;
	wire new_net_10222;
	wire n_0167_;
	wire new_net_3269;
	wire n_1175_;
	wire new_net_3411;
	wire n_0671_;
	wire n_0965_;
	wire n_0461_;
	wire new_net_4632;
	wire new_net_7629;
	wire new_net_7790;
	wire new_net_9473;
	wire new_net_6231;
	wire new_net_8186;
	wire new_net_8066;
	wire new_net_7773;
	wire new_net_8422;
	wire new_net_2856;
	wire new_net_3227;
	wire new_net_3282;
	wire new_net_34;
	wire new_net_3848;
	wire new_net_4678;
	wire new_net_5008;
	wire new_net_5032;
	wire new_net_5256;
	wire new_net_5723;
	wire new_net_6620;
	wire new_net_9770;
	wire new_net_6096;
	wire new_net_10167;
	wire new_net_10447;
	wire new_net_218;
	wire new_net_3076;
	wire new_net_1869;
	wire n_0168_;
	wire new_net_554;
	wire n_1176_;
	wire new_net_1494;
	wire n_0672_;
	wire n_0966_;
	wire n_0462_;
	wire new_net_4579;
	wire new_net_7048;
	wire new_net_9108;
	wire new_net_9696;
	wire new_net_9623;
	wire new_net_8811;
	wire new_net_4977;
	wire new_net_8424;
	wire new_net_6728;
	wire n_1220_;
	wire new_net_3031;
	wire new_net_3463;
	wire new_net_3095;
	wire n_0077_;
	wire new_net_402;
	wire new_net_2257;
	wire new_net_2712;
	wire new_net_2320;
	wire new_net_6212;
	wire new_net_6550;
	wire new_net_8850;
	wire new_net_10629;
	wire new_net_3615;
	wire new_net_3270;
	wire n_0463_;
	wire n_1177_;
	wire n_0673_;
	wire n_0967_;
	wire n_0169_;
	wire n_0420_;
	wire new_net_4460;
	wire new_net_4655;
	wire new_net_5045;
	wire new_net_6916;
	wire new_net_8240;
	wire new_net_8680;
	wire new_net_6844;
	wire new_net_4256;
	wire n_1040_;
	wire new_net_10490;
	wire new_net_2897;
	wire new_net_3335;
	wire new_net_818;
	wire new_net_932;
	wire new_net_1722;
	wire new_net_4270;
	wire new_net_4615;
	wire new_net_4852;
	wire new_net_5048;
	wire new_net_6207;
	wire new_net_10186;
	wire new_net_9520;
	wire new_net_669;
	wire new_net_219;
	wire n_0968_;
	wire new_net_1495;
	wire n_0464_;
	wire n_1178_;
	wire n_0170_;
	wire n_0674_;
	wire new_net_3662;
	wire new_net_3709;
	wire new_net_7863;
	wire new_net_7861;
	wire new_net_2867;
	wire new_net_7367;
	wire new_net_7624;
	wire new_net_5112;
	wire new_net_1610;
	wire new_net_2457;
	wire new_net_2226;
	wire new_net_403;
	wire new_net_4633;
	wire new_net_7630;
	wire new_net_7791;
	wire new_net_8062;
	wire new_net_8086;
	wire new_net_8483;
	wire new_net_7711;
	wire n_0901_;
	wire new_net_8922;
	wire new_net_8003;
	wire new_net_10584;
	wire new_net_8538;
	wire new_net_9667;
	wire new_net_236;
	wire new_net_4665;
	wire new_net_4549;
	wire new_net_8413;
	wire new_net_3456;
	wire new_net_2857;
	wire n_0171_;
	wire new_net_35;
	wire new_net_365;
	wire n_0675_;
	wire n_0969_;
	wire n_0465_;
	wire n_1179_;
	wire new_net_4679;
	wire new_net_5009;
	wire new_net_7275;
	wire new_net_9761;
	wire new_net_8106;
	wire new_net_3168;
	wire new_net_4598;
	wire new_net_10549;
	wire new_net_5733;
	wire new_net_10158;
	wire n_0001_;
	wire new_net_6869;
	wire new_net_277;
	wire new_net_1870;
	wire new_net_3077;
	wire new_net_522;
	wire new_net_555;
	wire new_net_819;
	wire new_net_933;
	wire new_net_3918;
	wire new_net_3965;
	wire new_net_544;
	wire new_net_3989;
	wire new_net_2142;
	wire new_net_4373;
	wire new_net_8870;
	wire new_net_7132;
	wire new_net_10061;
	wire new_net_4371;
	wire new_net_7095;
	wire new_net_6420;
	wire new_net_4169;
	wire new_net_5740;
	wire new_net_3032;
	wire n_0466_;
	wire new_net_670;
	wire new_net_220;
	wire new_net_3464;
	wire n_0172_;
	wire new_net_3096;
	wire n_0676_;
	wire n_0970_;
	wire n_1180_;
	wire new_net_6516;
	wire new_net_7178;
	wire new_net_10380;
	wire n_0217_;
	wire new_net_3772;
	wire new_net_694;
	wire new_net_5214;
	wire new_net_5143;
	wire new_net_2321;
	wire new_net_2104;
	wire new_net_3616;
	wire new_net_3271;
	wire new_net_1083;
	wire new_net_2258;
	wire new_net_4461;
	wire new_net_4656;
	wire new_net_5407;
	wire new_net_5431;
	wire n_0567_;
	wire new_net_6179;
	wire new_net_4843;
	wire new_net_8909;
	wire new_net_5698;
	wire new_net_366;
	wire new_net_2898;
	wire n_0173_;
	wire new_net_36;
	wire new_net_3336;
	wire n_0467_;
	wire n_1181_;
	wire n_0677_;
	wire n_0971_;
	wire new_net_1726;
	wire new_net_5535;
	wire new_net_6146;
	wire new_net_8665;
	wire new_net_9266;
	wire new_net_9793;
	wire new_net_8253;
	wire new_net_9791;
	wire n_1221_;
	wire new_net_1496;
	wire new_net_1724;
	wire new_net_2099;
	wire new_net_1871;
	wire new_net_523;
	wire new_net_556;
	wire new_net_820;
	wire new_net_934;
	wire new_net_3663;
	wire new_net_3710;
	wire new_net_4756;
	wire new_net_5380;
	wire new_net_8220;
	wire new_net_9406;
	wire new_net_10004;
	wire new_net_8748;
	wire new_net_6703;
	wire new_net_3823;
	wire n_0698_;
	wire new_net_7903;
	wire new_net_5072;
	wire new_net_9730;
	wire n_0678_;
	wire new_net_404;
	wire new_net_671;
	wire new_net_221;
	wire new_net_1611;
	wire new_net_3054;
	wire n_0972_;
	wire n_0174_;
	wire n_0468_;
	wire n_1182_;
	wire new_net_5851;
	wire new_net_10245;
	wire new_net_7990;
	wire new_net_7289;
	wire new_net_1433;
	wire new_net_8045;
	wire new_net_9943;
	wire new_net_10284;
	wire n_1041_;
	wire new_net_1671;
	wire new_net_4540;
	wire new_net_6369;
	wire new_net_1084;
	wire new_net_2858;
	wire new_net_2458;
	wire new_net_908;
	wire new_net_2227;
	wire new_net_5010;
	wire new_net_5034;
	wire new_net_4426;
	wire new_net_5258;
	wire new_net_5725;
	wire new_net_8215;
	wire new_net_10032;
	wire new_net_6200;
	wire new_net_4047;
	wire new_net_10030;
	wire new_net_4586;
	wire new_net_8097;
	wire new_net_8298;
	wire new_net_8930;
	wire new_net_9563;
	wire new_net_9556;
	wire new_net_8928;
	wire new_net_9445;
	wire new_net_7810;
	wire new_net_10344;
	wire new_net_367;
	wire new_net_3078;
	wire n_0175_;
	wire n_0679_;
	wire n_0973_;
	wire n_0469_;
	wire n_1183_;
	wire new_net_3919;
	wire new_net_3966;
	wire new_net_3990;
	wire new_net_940;
	wire new_net_9887;
	wire new_net_2615;
	wire new_net_6271;
	wire new_net_4954;
	wire new_net_7081;
	wire new_net_9381;
	wire n_0282_;
	wire new_net_3513;
	wire new_net_5485;
	wire new_net_10562;
	wire new_net_5988;
	wire new_net_1497;
	wire new_net_1725;
	wire new_net_2129;
	wire new_net_3033;
	wire new_net_3465;
	wire new_net_3097;
	wire new_net_821;
	wire new_net_935;
	wire new_net_2956;
	wire new_net_4788;
	wire new_net_3226;
	wire new_net_8832;
	wire new_net_9354;
	wire new_net_10608;
	wire new_net_8367;
	wire new_net_6335;
	wire new_net_5955;
	wire new_net_7220;
	wire new_net_8058;
	wire new_net_2803;
	wire n_1184_;
	wire new_net_405;
	wire n_0470_;
	wire new_net_672;
	wire new_net_222;
	wire new_net_1612;
	wire new_net_3617;
	wire n_0176_;
	wire new_net_3272;
	wire n_0680_;
	wire new_net_8972;
	wire new_net_10231;
	wire new_net_6698;
	wire new_net_6821;
	wire new_net_7479;
	wire new_net_4233;
	wire new_net_9170;
	wire new_net_9531;
	wire n_0002_;
	wire new_net_6496;
	wire new_net_3337;
	wire new_net_1085;
	wire new_net_2259;
	wire new_net_2322;
	wire new_net_3228;
	wire new_net_2899;
	wire new_net_3257;
	wire new_net_37;
	wire n_1286_;
	wire new_net_4272;
	wire new_net_9688;
	wire new_net_8652;
	wire new_net_9504;
	wire new_net_7949;
	wire new_net_9850;
	wire new_net_1544;
	wire new_net_9701;
	wire new_net_9313;
	input N1;
	input N100;
	input N103;
	input N106;
	input N109;
	input N110;
	input N111;
	input N112;
	input N113;
	input N114;
	input N115;
	input N118;
	input N12;
	input N121;
	input N124;
	input N127;
	input N130;
	input N133;
	input N134;
	input N135;
	input N138;
	input N141;
	input N144;
	input N147;
	input N15;
	input N150;
	input N151;
	input N152;
	input N153;
	input N154;
	input N155;
	input N156;
	input N157;
	input N158;
	input N159;
	input N160;
	input N161;
	input N162;
	input N163;
	input N164;
	input N165;
	input N166;
	input N167;
	input N168;
	input N169;
	input N170;
	input N171;
	input N172;
	input N173;
	input N174;
	input N175;
	input N176;
	input N177;
	input N178;
	input N179;
	input N18;
	input N180;
	input N181;
	input N182;
	input N183;
	input N184;
	input N185;
	input N186;
	input N187;
	input N188;
	input N189;
	input N190;
	input N191;
	input N192;
	input N193;
	input N194;
	input N195;
	input N196;
	input N197;
	input N198;
	input N199;
	input N200;
	input N201;
	input N202;
	input N203;
	input N204;
	input N205;
	input N206;
	input N207;
	input N208;
	input N209;
	input N210;
	input N211;
	input N212;
	input N213;
	input N214;
	input N215;
	input N216;
	input N217;
	input N218;
	input N219;
	input N220;
	input N221;
	input N222;
	input N223;
	input N224;
	input N225;
	input N226;
	input N227;
	input N228;
	input N229;
	input N23;
	input N230;
	input N231;
	input N232;
	input N233;
	input N234;
	input N235;
	input N236;
	input N237;
	input N238;
	input N239;
	input N240;
	input N241_I;
	input N242;
	input N245;
	input N248;
	input N251;
	input N254;
	input N257;
	input N26;
	input N260;
	input N263;
	input N267;
	input N271;
	input N274;
	input N277;
	input N280;
	input N283;
	input N286;
	input N289;
	input N29;
	input N293;
	input N296;
	input N299;
	input N303;
	input N307;
	input N310;
	input N313;
	input N316;
	input N319;
	input N32;
	input N322;
	input N325;
	input N328;
	input N331;
	input N334;
	input N337;
	input N340;
	input N343;
	input N346;
	input N349;
	input N35;
	input N352;
	input N355;
	input N358;
	input N361;
	input N364;
	input N367;
	input N38;
	input N382;
	input N41;
	input N44;
	input N47;
	input N5;
	input N50;
	input N53;
	input N54;
	input N55;
	input N56;
	input N57;
	input N58;
	input N59;
	input N60;
	input N61;
	input N62;
	input N63;
	input N64;
	input N65;
	input N66;
	input N69;
	input N70;
	input N73;
	input N74;
	input N75;
	input N76;
	input N77;
	input N78;
	input N79;
	input N80;
	input N81;
	input N82;
	input N83;
	input N84;
	input N85;
	input N86;
	input N87;
	input N88;
	input N89;
	input N9;
	input N94;
	input N97;
	output N10025;
	output N10101;
	output N10102;
	output N10103;
	output N10104;
	output N10109;
	output N10110;
	output N10111;
	output N10112;
	output N10350;
	output N10351;
	output N10352;
	output N10353;
	output N10574;
	output N10575;
	output N10576;
	output N10628;
	output N10632;
	output N10641;
	output N10704;
	output N10706;
	output N10711;
	output N10712;
	output N10713;
	output N10714;
	output N10715;
	output N10716;
	output N10717;
	output N10718;
	output N10729;
	output N10759;
	output N10760;
	output N10761;
	output N10762;
	output N10763;
	output N10827;
	output N10837;
	output N10838;
	output N10839;
	output N10840;
	output N10868;
	output N10869;
	output N10870;
	output N10871;
	output N10905;
	output N10906;
	output N10907;
	output N10908;
	output N1110;
	output N1111;
	output N1112;
	output N1113;
	output N1114;
	output N11333;
	output N11334;
	output N11340;
	output N11342;
	output N1489;
	output N1490;
	output N1781;
	output N241_O;
	output N387;
	output N388;
	output N478;
	output N482;
	output N484;
	output N486;
	output N489;
	output N492;
	output N501;
	output N505;
	output N507;
	output N509;
	output N511;
	output N513;
	output N515;
	output N517;
	output N519;
	output N535;
	output N537;
	output N539;
	output N541;
	output N543;
	output N545;
	output N547;
	output N549;
	output N551;
	output N553;
	output N556;
	output N559;
	output N561;
	output N563;
	output N565;
	output N567;
	output N569;
	output N571;
	output N573;
	output N582;
	output N643;
	output N707;
	output N813;
	output N881;
	output N882;
	output N883;
	output N884;
	output N885;
	output N889;
	output N945;

	or_bb n_1372_ (
		.a(new_net_826),
		.b(new_net_2183),
		.c(new_net_2562)
	);

	or_ii n_1373_ (
		.a(N184),
		.b(N150),
		.c(n_0653_)
	);

	or_ii n_1374_ (
		.a(N240),
		.b(N228),
		.c(n_0654_)
	);

	or_bb n_1375_ (
		.a(n_0654_),
		.b(n_0653_),
		.c(new_net_1)
	);

	or_ii n_1376_ (
		.a(N152),
		.b(N210),
		.c(n_0655_)
	);

	or_ii n_1377_ (
		.a(N230),
		.b(N218),
		.c(n_0656_)
	);

	or_bb n_1378_ (
		.a(n_0656_),
		.b(n_0655_),
		.c(new_net_0)
	);

	or_ii n_1379_ (
		.a(N182),
		.b(N183),
		.c(n_0657_)
	);

	or_ii n_1380_ (
		.a(N186),
		.b(N185),
		.c(n_0658_)
	);

	or_bb n_1381_ (
		.a(n_0658_),
		.b(n_0657_),
		.c(new_net_3)
	);

	or_ii n_1382_ (
		.a(N172),
		.b(N162),
		.c(n_0659_)
	);

	or_ii n_1383_ (
		.a(N199),
		.b(N188),
		.c(n_0660_)
	);

	or_bb n_1384_ (
		.a(n_0660_),
		.b(n_0659_),
		.c(new_net_2)
	);

	or_bi n_1385_ (
		.a(new_net_827),
		.b(new_net_2184),
		.c(new_net_10)
	);

	inv n_1386_ (
		.din(N15),
		.dout(new_net_11)
	);

	and_bi n_1387_ (
		.a(new_net_2185),
		.b(new_net_828),
		.c(n_0661_)
	);

	or_ii n_1388_ (
		.a(n_0661_),
		.b(new_net_2186),
		.c(new_net_12)
	);

	or_bi n_1389_ (
		.a(new_net_120),
		.b(new_net_1486),
		.c(n_0662_)
	);

	or_bb n_1390_ (
		.a(new_net_641),
		.b(new_net_511),
		.c(n_0663_)
	);

	or_bb n_1391_ (
		.a(new_net_1487),
		.b(new_net_195),
		.c(n_0664_)
	);

	and_bi n_1392_ (
		.a(new_net_512),
		.b(n_0664_),
		.c(n_0665_)
	);

	or_bi n_1393_ (
		.a(new_net_1611),
		.b(new_net_733),
		.c(n_0666_)
	);

	and_bi n_1394_ (
		.a(new_net_960),
		.b(new_net_1059),
		.c(n_0667_)
	);

	inv n_1395_ (
		.din(new_net_962),
		.dout(n_0668_)
	);

	or_ii n_1396_ (
		.a(new_net_1061),
		.b(new_net_1676),
		.c(n_0669_)
	);

	and_bi n_1397_ (
		.a(new_net_2187),
		.b(new_net_1654),
		.c(new_net_2531)
	);

	inv n_1398_ (
		.din(new_net_1078),
		.dout(n_0670_)
	);

	and_bb n_1399_ (
		.a(new_net_2188),
		.b(new_net_196),
		.c(n_0671_)
	);

	and_bi n_1400_ (
		.a(new_net_2189),
		.b(new_net_132),
		.c(n_0672_)
	);

	and_ii n_1401_ (
		.a(new_net_1751),
		.b(new_net_2190),
		.c(n_0673_)
	);

	and_bi n_1402_ (
		.a(new_net_1452),
		.b(new_net_1771),
		.c(n_0674_)
	);

	and_bi n_1403_ (
		.a(new_net_1774),
		.b(new_net_1453),
		.c(n_0675_)
	);

	and_ii n_1404_ (
		.a(new_net_1801),
		.b(new_net_1874),
		.c(n_0676_)
	);

	or_ii n_1405_ (
		.a(new_net_2191),
		.b(new_net_192),
		.c(n_0677_)
	);

	and_bi n_1406_ (
		.a(new_net_2192),
		.b(new_net_125),
		.c(n_0678_)
	);

	and_bi n_1407_ (
		.a(new_net_2193),
		.b(new_net_1889),
		.c(n_0679_)
	);

	or_ii n_1408_ (
		.a(new_net_1911),
		.b(new_net_1386),
		.c(n_0680_)
	);

	or_ii n_1409_ (
		.a(new_net_2194),
		.b(new_net_135),
		.c(n_0681_)
	);

	and_bi n_1410_ (
		.a(new_net_2195),
		.b(new_net_250),
		.c(n_0682_)
	);

	and_bi n_1411_ (
		.a(new_net_2196),
		.b(new_net_1104),
		.c(n_0683_)
	);

	or_ii n_1412_ (
		.a(new_net_1118),
		.b(new_net_1354),
		.c(n_0684_)
	);

	and_ii n_1413_ (
		.a(new_net_1119),
		.b(new_net_1356),
		.c(n_0685_)
	);

	and_bi n_1414_ (
		.a(new_net_353),
		.b(new_net_509),
		.c(n_0686_)
	);

	or_ii n_1415_ (
		.a(new_net_2197),
		.b(new_net_130),
		.c(n_0687_)
	);

	and_bi n_1416_ (
		.a(new_net_2198),
		.b(new_net_246),
		.c(n_0688_)
	);

	or_bi n_1417_ (
		.a(new_net_845),
		.b(new_net_2199),
		.c(n_0689_)
	);

	and_bi n_1418_ (
		.a(new_net_1329),
		.b(new_net_942),
		.c(n_0690_)
	);

	and_bi n_1419_ (
		.a(new_net_943),
		.b(new_net_1330),
		.c(n_0691_)
	);

	or_bb n_1420_ (
		.a(new_net_1259),
		.b(new_net_1063),
		.c(n_0692_)
	);

	or_bb n_1421_ (
		.a(new_net_1282),
		.b(new_net_1062),
		.c(n_0693_)
	);

	and_bi n_1422_ (
		.a(new_net_1171),
		.b(new_net_1338),
		.c(n_0694_)
	);

	or_ii n_1423_ (
		.a(new_net_1454),
		.b(new_net_961),
		.c(n_0695_)
	);

	and_ii n_1424_ (
		.a(new_net_1912),
		.b(new_net_1388),
		.c(n_0696_)
	);

	or_bb n_1425_ (
		.a(new_net_1064),
		.b(new_net_736),
		.c(n_0697_)
	);

	or_bb n_1426_ (
		.a(new_net_1262),
		.b(new_net_510),
		.c(n_0698_)
	);

	and_bi n_1427_ (
		.a(new_net_1762),
		.b(new_net_2200),
		.c(n_0699_)
	);

	and_bi n_1428_ (
		.a(new_net_354),
		.b(n_0699_),
		.c(n_0700_)
	);

	and_ii n_1429_ (
		.a(new_net_1469),
		.b(new_net_1670),
		.c(n_0701_)
	);

	and_bb n_1430_ (
		.a(new_net_360),
		.b(new_net_1352),
		.c(n_0702_)
	);

	and_bi n_1431_ (
		.a(new_net_737),
		.b(n_0702_),
		.c(n_0703_)
	);

	or_ii n_1432_ (
		.a(new_net_1536),
		.b(new_net_104),
		.c(n_0704_)
	);

	and_ii n_1433_ (
		.a(new_net_1537),
		.b(new_net_106),
		.c(n_0705_)
	);

	and_bi n_1434_ (
		.a(n_0704_),
		.b(n_0705_),
		.c(new_net_2568)
	);

	or_bi n_1435_ (
		.a(new_net_1472),
		.b(new_net_1353),
		.c(n_0706_)
	);

	or_bi n_1436_ (
		.a(new_net_1671),
		.b(new_net_738),
		.c(n_0707_)
	);

	or_ii n_1437_ (
		.a(new_net_1075),
		.b(new_net_952),
		.c(n_0708_)
	);

	or_bb n_1438_ (
		.a(new_net_1074),
		.b(new_net_953),
		.c(n_0709_)
	);

	or_ii n_1439_ (
		.a(n_0709_),
		.b(n_0708_),
		.c(new_net_2513)
	);

	and_bi n_1440_ (
		.a(new_net_734),
		.b(new_net_1261),
		.c(n_0710_)
	);

	and_bi n_1441_ (
		.a(new_net_1347),
		.b(new_net_1656),
		.c(n_0711_)
	);

	and_ii n_1442_ (
		.a(n_0711_),
		.b(new_net_1066),
		.c(n_0712_)
	);

	and_bi n_1443_ (
		.a(new_net_1709),
		.b(new_net_1175),
		.c(n_0713_)
	);

	and_bi n_1444_ (
		.a(new_net_1172),
		.b(new_net_1710),
		.c(n_0714_)
	);

	or_bb n_1445_ (
		.a(n_0714_),
		.b(n_0713_),
		.c(new_net_2558)
	);

	and_bi n_1446_ (
		.a(new_net_735),
		.b(new_net_1655),
		.c(n_0715_)
	);

	and_bi n_1447_ (
		.a(new_net_1891),
		.b(new_net_1283),
		.c(n_0716_)
	);

	and_bi n_1448_ (
		.a(new_net_1285),
		.b(new_net_1892),
		.c(n_0717_)
	);

	or_bb n_1449_ (
		.a(n_0717_),
		.b(n_0716_),
		.c(new_net_2507)
	);

	and_bb n_1450_ (
		.a(N9),
		.b(N12),
		.c(n_0718_)
	);

	and_bi n_1451_ (
		.a(new_net_281),
		.b(new_net_2201),
		.c(n_0719_)
	);

	and_ii n_1452_ (
		.a(new_net_517),
		.b(new_net_383),
		.c(n_0720_)
	);

	and_bi n_1453_ (
		.a(new_net_148),
		.b(new_net_2202),
		.c(n_0721_)
	);

	or_ii n_1454_ (
		.a(new_net_1921),
		.b(new_net_647),
		.c(n_0722_)
	);

	and_ii n_1455_ (
		.a(new_net_1922),
		.b(new_net_378),
		.c(n_0723_)
	);

	and_bb n_1456_ (
		.a(new_net_17),
		.b(new_net_518),
		.c(n_0724_)
	);

	and_bi n_1457_ (
		.a(n_0722_),
		.b(n_0724_),
		.c(n_0725_)
	);

	and_bi n_1458_ (
		.a(new_net_224),
		.b(new_net_2203),
		.c(n_0726_)
	);

	and_ii n_1459_ (
		.a(new_net_47),
		.b(new_net_377),
		.c(n_0727_)
	);

	and_bi n_1460_ (
		.a(new_net_119),
		.b(new_net_2204),
		.c(n_0728_)
	);

	and_bb n_1461_ (
		.a(new_net_79),
		.b(new_net_56),
		.c(n_0729_)
	);

	and_ii n_1462_ (
		.a(new_net_80),
		.b(new_net_370),
		.c(n_0730_)
	);

	and_bb n_1463_ (
		.a(new_net_1836),
		.b(new_net_48),
		.c(n_0731_)
	);

	or_bb n_1464_ (
		.a(n_0731_),
		.b(n_0729_),
		.c(n_0732_)
	);

	and_bi n_1465_ (
		.a(new_net_2205),
		.b(new_net_193),
		.c(n_0733_)
	);

	and_bb n_1466_ (
		.a(new_net_2206),
		.b(new_net_126),
		.c(n_0734_)
	);

	and_ii n_1467_ (
		.a(new_net_2207),
		.b(new_net_338),
		.c(n_0735_)
	);

	and_bi n_1468_ (
		.a(new_net_2208),
		.b(new_net_183),
		.c(n_0736_)
	);

	and_bb n_1469_ (
		.a(new_net_2209),
		.b(new_net_136),
		.c(n_0737_)
	);

	and_ii n_1470_ (
		.a(new_net_2210),
		.b(new_net_721),
		.c(n_0738_)
	);

	and_bb n_1471_ (
		.a(new_net_484),
		.b(new_net_615),
		.c(n_0739_)
	);

	and_ii n_1472_ (
		.a(new_net_485),
		.b(new_net_616),
		.c(n_0740_)
	);

	and_ii n_1473_ (
		.a(n_0740_),
		.b(n_0739_),
		.c(n_0741_)
	);

	or_bb n_1474_ (
		.a(new_net_549),
		.b(new_net_297),
		.c(n_0742_)
	);

	and_bb n_1475_ (
		.a(new_net_550),
		.b(new_net_298),
		.c(n_0743_)
	);

	and_bi n_1476_ (
		.a(n_0742_),
		.b(n_0743_),
		.c(n_0744_)
	);

	and_ii n_1477_ (
		.a(new_net_1564),
		.b(new_net_35),
		.c(n_0745_)
	);

	and_bb n_1478_ (
		.a(new_net_1565),
		.b(new_net_36),
		.c(n_0746_)
	);

	and_ii n_1479_ (
		.a(n_0746_),
		.b(n_0745_),
		.c(n_0747_)
	);

	and_bi n_1480_ (
		.a(new_net_2211),
		.b(new_net_184),
		.c(n_0748_)
	);

	and_bb n_1481_ (
		.a(new_net_2212),
		.b(new_net_137),
		.c(n_0749_)
	);

	or_bb n_1482_ (
		.a(new_net_2213),
		.b(new_net_715),
		.c(n_0750_)
	);

	and_bi n_1483_ (
		.a(new_net_164),
		.b(new_net_2214),
		.c(n_0751_)
	);

	and_ii n_1484_ (
		.a(n_0751_),
		.b(new_net_385),
		.c(n_0752_)
	);

	or_bb n_1485_ (
		.a(new_net_793),
		.b(new_net_760),
		.c(n_0753_)
	);

	and_bb n_1486_ (
		.a(new_net_795),
		.b(new_net_761),
		.c(n_0754_)
	);

	and_bi n_1487_ (
		.a(n_0753_),
		.b(n_0754_),
		.c(n_0755_)
	);

	and_bi n_1488_ (
		.a(new_net_2215),
		.b(new_net_247),
		.c(n_0756_)
	);

	and_bb n_1489_ (
		.a(new_net_2216),
		.b(new_net_194),
		.c(n_0757_)
	);

	and_ii n_1490_ (
		.a(new_net_2217),
		.b(new_net_871),
		.c(n_0758_)
	);

	and_bi n_1491_ (
		.a(new_net_2218),
		.b(new_net_238),
		.c(n_0759_)
	);

	and_bb n_1492_ (
		.a(new_net_2219),
		.b(new_net_185),
		.c(n_0760_)
	);

	and_ii n_1493_ (
		.a(new_net_2220),
		.b(new_net_938),
		.c(n_0761_)
	);

	and_ii n_1494_ (
		.a(new_net_988),
		.b(new_net_918),
		.c(n_0762_)
	);

	and_bb n_1495_ (
		.a(new_net_990),
		.b(new_net_919),
		.c(n_0763_)
	);

	or_bb n_1496_ (
		.a(n_0763_),
		.b(n_0762_),
		.c(n_0764_)
	);

	and_ii n_1497_ (
		.a(new_net_1051),
		.b(new_net_862),
		.c(n_0765_)
	);

	and_bb n_1498_ (
		.a(new_net_1052),
		.b(new_net_863),
		.c(n_0766_)
	);

	and_ii n_1499_ (
		.a(n_0766_),
		.b(n_0765_),
		.c(n_0767_)
	);

	and_bb n_1500_ (
		.a(new_net_1116),
		.b(new_net_1849),
		.c(n_0768_)
	);

	and_bi n_1501_ (
		.a(new_net_149),
		.b(new_net_2221),
		.c(n_0769_)
	);

	and_bi n_1502_ (
		.a(new_net_807),
		.b(new_net_374),
		.c(n_0770_)
	);

	and_bi n_1503_ (
		.a(new_net_209),
		.b(new_net_2222),
		.c(n_0771_)
	);

	and_ii n_1504_ (
		.a(new_net_1011),
		.b(new_net_386),
		.c(n_0772_)
	);

	and_bi n_1505_ (
		.a(new_net_258),
		.b(new_net_2223),
		.c(n_0773_)
	);

	and_bb n_1506_ (
		.a(new_net_1191),
		.b(new_net_1193),
		.c(n_0774_)
	);

	and_ii n_1507_ (
		.a(new_net_1192),
		.b(new_net_379),
		.c(n_0775_)
	);

	and_bb n_1508_ (
		.a(new_net_1263),
		.b(new_net_1012),
		.c(n_0776_)
	);

	and_ii n_1509_ (
		.a(n_0776_),
		.b(n_0774_),
		.c(n_0777_)
	);

	or_bi n_1510_ (
		.a(new_net_901),
		.b(new_net_1640),
		.c(n_0778_)
	);

	and_bi n_1511_ (
		.a(new_net_902),
		.b(new_net_1641),
		.c(n_0779_)
	);

	and_bi n_1512_ (
		.a(n_0778_),
		.b(n_0779_),
		.c(n_0780_)
	);

	and_bi n_1513_ (
		.a(new_net_150),
		.b(new_net_2224),
		.c(n_0781_)
	);

	and_ii n_1514_ (
		.a(new_net_1405),
		.b(new_net_375),
		.c(n_0782_)
	);

	and_bi n_1515_ (
		.a(new_net_210),
		.b(new_net_2225),
		.c(n_0783_)
	);

	and_bb n_1516_ (
		.a(new_net_1443),
		.b(new_net_1425),
		.c(n_0784_)
	);

	and_ii n_1517_ (
		.a(new_net_1444),
		.b(new_net_389),
		.c(n_0785_)
	);

	and_bb n_1518_ (
		.a(new_net_1500),
		.b(new_net_1406),
		.c(n_0786_)
	);

	and_ii n_1519_ (
		.a(n_0786_),
		.b(n_0784_),
		.c(n_0787_)
	);

	or_bi n_1520_ (
		.a(new_net_387),
		.b(new_net_151),
		.c(n_0788_)
	);

	and_ii n_1521_ (
		.a(new_net_1032),
		.b(new_net_1057),
		.c(n_0789_)
	);

	and_bb n_1522_ (
		.a(new_net_1033),
		.b(new_net_1058),
		.c(n_0790_)
	);

	or_bb n_1523_ (
		.a(n_0790_),
		.b(n_0789_),
		.c(n_0791_)
	);

	and_ii n_1524_ (
		.a(new_net_2226),
		.b(new_net_1017),
		.c(n_0792_)
	);

	and_bb n_1525_ (
		.a(new_net_1632),
		.b(new_net_910),
		.c(n_0793_)
	);

	and_ii n_1526_ (
		.a(new_net_1633),
		.b(new_net_911),
		.c(n_0794_)
	);

	and_ii n_1527_ (
		.a(n_0794_),
		.b(n_0793_),
		.c(n_0795_)
	);

	or_bi n_1528_ (
		.a(new_net_1382),
		.b(new_net_1745),
		.c(n_0796_)
	);

	and_bi n_1529_ (
		.a(new_net_1383),
		.b(new_net_1746),
		.c(n_0797_)
	);

	and_bi n_1530_ (
		.a(n_0796_),
		.b(n_0797_),
		.c(n_0798_)
	);

	and_ii n_1531_ (
		.a(new_net_1117),
		.b(new_net_1850),
		.c(n_0799_)
	);

	or_bb n_1532_ (
		.a(n_0799_),
		.b(new_net_2227),
		.c(n_0800_)
	);

	or_bb n_1533_ (
		.a(n_0800_),
		.b(new_net_2228),
		.c(n_0801_)
	);

	and_bb n_1534_ (
		.a(new_net_2229),
		.b(new_net_211),
		.c(n_0802_)
	);

	and_bi n_1535_ (
		.a(new_net_2230),
		.b(new_net_143),
		.c(n_0803_)
	);

	and_ii n_1536_ (
		.a(new_net_1843),
		.b(new_net_2231),
		.c(n_0804_)
	);

	and_bb n_1537_ (
		.a(new_net_2232),
		.b(new_net_204),
		.c(n_0805_)
	);

	and_bi n_1538_ (
		.a(new_net_642),
		.b(new_net_2233),
		.c(n_0806_)
	);

	and_bi n_1539_ (
		.a(new_net_912),
		.b(new_net_1937),
		.c(n_0807_)
	);

	and_bi n_1540_ (
		.a(new_net_1938),
		.b(new_net_913),
		.c(n_0808_)
	);

	and_ii n_1541_ (
		.a(n_0808_),
		.b(n_0807_),
		.c(n_0809_)
	);

	and_bb n_1542_ (
		.a(new_net_2234),
		.b(new_net_282),
		.c(n_0810_)
	);

	and_bi n_1543_ (
		.a(new_net_2235),
		.b(new_net_217),
		.c(n_0811_)
	);

	and_ii n_1544_ (
		.a(new_net_1158),
		.b(new_net_2236),
		.c(n_0812_)
	);

	and_bi n_1545_ (
		.a(new_net_1914),
		.b(new_net_1020),
		.c(n_0813_)
	);

	and_bi n_1546_ (
		.a(new_net_1023),
		.b(new_net_1913),
		.c(n_0814_)
	);

	and_ii n_1547_ (
		.a(n_0814_),
		.b(n_0813_),
		.c(n_0815_)
	);

	and_bi n_1548_ (
		.a(new_net_706),
		.b(new_net_1310),
		.c(n_0816_)
	);

	and_bi n_1549_ (
		.a(new_net_1311),
		.b(new_net_707),
		.c(n_0817_)
	);

	or_bb n_1550_ (
		.a(n_0817_),
		.b(n_0816_),
		.c(n_0818_)
	);

	and_bi n_1551_ (
		.a(new_net_1773),
		.b(new_net_1121),
		.c(n_0819_)
	);

	and_bi n_1552_ (
		.a(new_net_1120),
		.b(new_net_1772),
		.c(n_0820_)
	);

	or_bb n_1553_ (
		.a(n_0820_),
		.b(n_0819_),
		.c(n_0821_)
	);

	or_ii n_1554_ (
		.a(new_net_2237),
		.b(new_net_283),
		.c(n_0822_)
	);

	and_bi n_1555_ (
		.a(new_net_2238),
		.b(new_net_218),
		.c(n_0823_)
	);

	and_bi n_1556_ (
		.a(new_net_2239),
		.b(new_net_1413),
		.c(n_0824_)
	);

	or_ii n_1557_ (
		.a(new_net_2240),
		.b(new_net_269),
		.c(n_0825_)
	);

	and_bi n_1558_ (
		.a(new_net_2241),
		.b(new_net_212),
		.c(n_0826_)
	);

	and_bi n_1559_ (
		.a(new_net_2242),
		.b(new_net_710),
		.c(n_0827_)
	);

	and_bi n_1560_ (
		.a(new_net_464),
		.b(new_net_1503),
		.c(n_0828_)
	);

	and_bi n_1561_ (
		.a(new_net_1506),
		.b(new_net_465),
		.c(n_0829_)
	);

	and_ii n_1562_ (
		.a(n_0829_),
		.b(n_0828_),
		.c(n_0830_)
	);

	and_bb n_1563_ (
		.a(new_net_2243),
		.b(new_net_251),
		.c(n_0831_)
	);

	and_bi n_1564_ (
		.a(new_net_2244),
		.b(new_net_197),
		.c(n_0832_)
	);

	and_ii n_1565_ (
		.a(new_net_1316),
		.b(new_net_2245),
		.c(n_0833_)
	);

	and_bi n_1566_ (
		.a(new_net_1614),
		.b(new_net_945),
		.c(n_0834_)
	);

	and_bi n_1567_ (
		.a(new_net_944),
		.b(new_net_1615),
		.c(n_0835_)
	);

	and_ii n_1568_ (
		.a(n_0835_),
		.b(n_0834_),
		.c(n_0836_)
	);

	and_ii n_1569_ (
		.a(new_net_1747),
		.b(new_net_1558),
		.c(n_0837_)
	);

	and_bb n_1570_ (
		.a(new_net_1748),
		.b(new_net_1559),
		.c(n_0838_)
	);

	or_bb n_1571_ (
		.a(n_0838_),
		.b(n_0837_),
		.c(n_0839_)
	);

	and_ii n_1572_ (
		.a(new_net_1739),
		.b(new_net_15),
		.c(n_0840_)
	);

	and_bb n_1573_ (
		.a(new_net_1740),
		.b(new_net_16),
		.c(n_0841_)
	);

	and_ii n_1574_ (
		.a(n_0841_),
		.b(n_0840_),
		.c(n_0842_)
	);

	or_bi n_1575_ (
		.a(new_net_1642),
		.b(new_net_605),
		.c(n_0843_)
	);

	and_bi n_1576_ (
		.a(new_net_1643),
		.b(new_net_606),
		.c(n_0844_)
	);

	and_bi n_1577_ (
		.a(n_0843_),
		.b(n_0844_),
		.c(n_0845_)
	);

	and_bb n_1578_ (
		.a(new_net_2246),
		.b(new_net_284),
		.c(n_0846_)
	);

	and_bi n_1579_ (
		.a(new_net_2247),
		.b(new_net_219),
		.c(n_0847_)
	);

	or_bb n_1580_ (
		.a(new_net_1919),
		.b(new_net_2248),
		.c(n_0848_)
	);

	and_bb n_1581_ (
		.a(new_net_2249),
		.b(new_net_270),
		.c(n_0849_)
	);

	and_bi n_1582_ (
		.a(new_net_2250),
		.b(new_net_213),
		.c(n_0850_)
	);

	and_ii n_1583_ (
		.a(new_net_1619),
		.b(new_net_2251),
		.c(n_0851_)
	);

	or_bb n_1584_ (
		.a(new_net_37),
		.b(new_net_1941),
		.c(n_0852_)
	);

	and_bb n_1585_ (
		.a(new_net_40),
		.b(new_net_1942),
		.c(n_0853_)
	);

	and_bi n_1586_ (
		.a(n_0852_),
		.b(n_0853_),
		.c(n_0854_)
	);

	or_ii n_1587_ (
		.a(new_net_2252),
		.b(new_net_252),
		.c(n_0855_)
	);

	and_bi n_1588_ (
		.a(new_net_2253),
		.b(new_net_198),
		.c(n_0856_)
	);

	and_bi n_1589_ (
		.a(new_net_2254),
		.b(new_net_433),
		.c(n_0857_)
	);

	and_bb n_1590_ (
		.a(new_net_2255),
		.b(new_net_280),
		.c(n_0858_)
	);

	and_bi n_1591_ (
		.a(new_net_2256),
		.b(new_net_220),
		.c(n_0859_)
	);

	and_ii n_1592_ (
		.a(new_net_327),
		.b(new_net_2257),
		.c(n_0860_)
	);

	and_ii n_1593_ (
		.a(new_net_881),
		.b(new_net_563),
		.c(n_0861_)
	);

	and_bb n_1594_ (
		.a(new_net_884),
		.b(new_net_565),
		.c(n_0862_)
	);

	and_ii n_1595_ (
		.a(n_0862_),
		.b(n_0861_),
		.c(n_0863_)
	);

	or_bb n_1596_ (
		.a(new_net_1182),
		.b(new_net_77),
		.c(n_0864_)
	);

	and_bb n_1597_ (
		.a(new_net_1183),
		.b(new_net_78),
		.c(n_0865_)
	);

	and_bi n_1598_ (
		.a(n_0864_),
		.b(n_0865_),
		.c(n_0866_)
	);

	and_bb n_1599_ (
		.a(new_net_2258),
		.b(new_net_248),
		.c(n_0867_)
	);

	and_bi n_1600_ (
		.a(new_net_2259),
		.b(new_net_199),
		.c(n_0868_)
	);

	and_ii n_1601_ (
		.a(new_net_1726),
		.b(new_net_2260),
		.c(n_0869_)
	);

	or_ii n_1602_ (
		.a(new_net_2261),
		.b(new_net_279),
		.c(n_0870_)
	);

	and_bi n_1603_ (
		.a(new_net_2262),
		.b(new_net_221),
		.c(n_0871_)
	);

	and_bi n_1604_ (
		.a(new_net_2263),
		.b(new_net_67),
		.c(n_0872_)
	);

	and_bb n_1605_ (
		.a(new_net_307),
		.b(new_net_598),
		.c(n_0873_)
	);

	and_ii n_1606_ (
		.a(new_net_310),
		.b(new_net_599),
		.c(n_0874_)
	);

	and_ii n_1607_ (
		.a(n_0874_),
		.b(n_0873_),
		.c(n_0875_)
	);

	and_bb n_1608_ (
		.a(new_net_2264),
		.b(new_net_259),
		.c(n_0876_)
	);

	and_bi n_1609_ (
		.a(new_net_2265),
		.b(new_net_205),
		.c(n_0877_)
	);

	and_ii n_1610_ (
		.a(new_net_774),
		.b(new_net_2266),
		.c(n_0878_)
	);

	and_bb n_1611_ (
		.a(new_net_2267),
		.b(new_net_249),
		.c(n_0879_)
	);

	and_bi n_1612_ (
		.a(new_net_2268),
		.b(new_net_200),
		.c(n_0880_)
	);

	and_ii n_1613_ (
		.a(new_net_841),
		.b(new_net_2269),
		.c(n_0881_)
	);

	and_bi n_1614_ (
		.a(new_net_797),
		.b(new_net_1298),
		.c(n_0882_)
	);

	and_bi n_1615_ (
		.a(new_net_1299),
		.b(new_net_799),
		.c(n_0883_)
	);

	and_ii n_1616_ (
		.a(n_0883_),
		.b(n_0882_),
		.c(n_0884_)
	);

	or_ii n_1617_ (
		.a(new_net_2270),
		.b(new_net_271),
		.c(n_0885_)
	);

	and_bi n_1618_ (
		.a(new_net_2271),
		.b(new_net_214),
		.c(n_0886_)
	);

	and_bi n_1619_ (
		.a(new_net_2272),
		.b(new_net_972),
		.c(n_0887_)
	);

	or_ii n_1620_ (
		.a(new_net_2273),
		.b(new_net_260),
		.c(n_0888_)
	);

	and_bi n_1621_ (
		.a(new_net_2274),
		.b(new_net_206),
		.c(n_0889_)
	);

	and_bi n_1622_ (
		.a(new_net_2275),
		.b(new_net_1026),
		.c(n_0890_)
	);

	and_ii n_1623_ (
		.a(new_net_1053),
		.b(new_net_1957),
		.c(n_0891_)
	);

	and_bb n_1624_ (
		.a(new_net_1056),
		.b(new_net_1958),
		.c(n_0892_)
	);

	and_ii n_1625_ (
		.a(n_0892_),
		.b(n_0891_),
		.c(n_0893_)
	);

	and_bi n_1626_ (
		.a(new_net_916),
		.b(new_net_994),
		.c(n_0894_)
	);

	and_bi n_1627_ (
		.a(new_net_995),
		.b(new_net_917),
		.c(n_0895_)
	);

	and_ii n_1628_ (
		.a(n_0895_),
		.b(n_0894_),
		.c(n_0896_)
	);

	and_bi n_1629_ (
		.a(new_net_1272),
		.b(new_net_696),
		.c(n_0897_)
	);

	and_bi n_1630_ (
		.a(new_net_697),
		.b(new_net_1273),
		.c(n_0898_)
	);

	and_ii n_1631_ (
		.a(n_0898_),
		.b(n_0897_),
		.c(n_0899_)
	);

	or_bi n_1632_ (
		.a(new_net_528),
		.b(new_net_1211),
		.c(n_0900_)
	);

	and_bi n_1633_ (
		.a(new_net_529),
		.b(new_net_1212),
		.c(n_0901_)
	);

	and_bi n_1634_ (
		.a(n_0900_),
		.b(n_0901_),
		.c(n_0902_)
	);

	or_bb n_1635_ (
		.a(n_0902_),
		.b(n_0845_),
		.c(n_0903_)
	);

	or_bb n_1636_ (
		.a(n_0903_),
		.b(n_0801_),
		.c(new_net_4)
	);

	or_bi n_1637_ (
		.a(new_net_127),
		.b(new_net_2276),
		.c(n_0904_)
	);

	and_bi n_1638_ (
		.a(new_net_239),
		.b(new_net_847),
		.c(n_0905_)
	);

	and_bi n_1639_ (
		.a(n_0904_),
		.b(n_0905_),
		.c(n_0906_)
	);

	and_bi n_1640_ (
		.a(new_net_2277),
		.b(new_net_152),
		.c(n_0907_)
	);

	and_bi n_1641_ (
		.a(new_net_232),
		.b(new_net_946),
		.c(n_0908_)
	);

	and_ii n_1642_ (
		.a(n_0908_),
		.b(n_0907_),
		.c(n_0909_)
	);

	and_ii n_1643_ (
		.a(new_net_1439),
		.b(new_net_553),
		.c(n_0910_)
	);

	and_bb n_1644_ (
		.a(new_net_1442),
		.b(new_net_554),
		.c(n_0911_)
	);

	and_ii n_1645_ (
		.a(n_0911_),
		.b(n_0910_),
		.c(n_0912_)
	);

	and_bi n_1646_ (
		.a(new_net_2278),
		.b(new_net_133),
		.c(n_0913_)
	);

	and_bi n_1647_ (
		.a(new_net_225),
		.b(new_net_1805),
		.c(n_0914_)
	);

	and_ii n_1648_ (
		.a(n_0914_),
		.b(n_0913_),
		.c(n_0915_)
	);

	or_bi n_1649_ (
		.a(new_net_128),
		.b(new_net_2279),
		.c(n_0916_)
	);

	and_bi n_1650_ (
		.a(new_net_240),
		.b(new_net_1343),
		.c(n_0917_)
	);

	and_bi n_1651_ (
		.a(n_0916_),
		.b(n_0917_),
		.c(n_0918_)
	);

	and_bi n_1652_ (
		.a(new_net_1582),
		.b(new_net_1797),
		.c(n_0919_)
	);

	and_bi n_1653_ (
		.a(new_net_1799),
		.b(new_net_1584),
		.c(n_0920_)
	);

	and_ii n_1654_ (
		.a(n_0920_),
		.b(n_0919_),
		.c(n_0921_)
	);

	and_ii n_1655_ (
		.a(new_net_1700),
		.b(new_net_1522),
		.c(n_0922_)
	);

	and_bb n_1656_ (
		.a(new_net_1701),
		.b(new_net_1523),
		.c(n_0923_)
	);

	or_bb n_1657_ (
		.a(n_0923_),
		.b(n_0922_),
		.c(n_0924_)
	);

	and_bi n_1658_ (
		.a(new_net_2280),
		.b(new_net_134),
		.c(n_0925_)
	);

	and_bi n_1659_ (
		.a(new_net_226),
		.b(new_net_1069),
		.c(n_0926_)
	);

	and_ii n_1660_ (
		.a(n_0926_),
		.b(n_0925_),
		.c(n_0927_)
	);

	and_bi n_1661_ (
		.a(new_net_2281),
		.b(new_net_158),
		.c(n_0928_)
	);

	and_bi n_1662_ (
		.a(new_net_241),
		.b(new_net_1722),
		.c(n_0929_)
	);

	and_ii n_1663_ (
		.a(n_0929_),
		.b(n_0928_),
		.c(n_0930_)
	);

	and_ii n_1664_ (
		.a(new_net_1881),
		.b(new_net_996),
		.c(n_0931_)
	);

	and_bb n_1665_ (
		.a(new_net_1883),
		.b(new_net_998),
		.c(n_0932_)
	);

	and_ii n_1666_ (
		.a(n_0932_),
		.b(n_0931_),
		.c(n_0933_)
	);

	or_bi n_1667_ (
		.a(new_net_1915),
		.b(new_net_1464),
		.c(n_0934_)
	);

	and_bi n_1668_ (
		.a(new_net_1917),
		.b(new_net_1468),
		.c(n_0935_)
	);

	and_bi n_1669_ (
		.a(n_0934_),
		.b(n_0935_),
		.c(n_0936_)
	);

	and_bi n_1670_ (
		.a(new_net_121),
		.b(new_net_2282),
		.c(n_0937_)
	);

	or_bb n_1671_ (
		.a(new_net_1674),
		.b(new_net_1730),
		.c(n_0938_)
	);

	and_bb n_1672_ (
		.a(new_net_1675),
		.b(new_net_1731),
		.c(n_0939_)
	);

	or_bb n_1673_ (
		.a(new_net_1176),
		.b(new_net_159),
		.c(n_0940_)
	);

	and_bi n_1674_ (
		.a(new_net_1169),
		.b(n_0940_),
		.c(n_0941_)
	);

	and_ii n_1675_ (
		.a(n_0941_),
		.b(new_net_2283),
		.c(n_0942_)
	);

	and_ii n_1676_ (
		.a(new_net_1229),
		.b(new_net_1098),
		.c(n_0943_)
	);

	and_bb n_1677_ (
		.a(new_net_1230),
		.b(new_net_1099),
		.c(n_0944_)
	);

	and_ii n_1678_ (
		.a(n_0944_),
		.b(n_0943_),
		.c(n_0945_)
	);

	or_bb n_1679_ (
		.a(new_net_1304),
		.b(new_net_682),
		.c(n_0946_)
	);

	and_bb n_1680_ (
		.a(new_net_1305),
		.b(new_net_683),
		.c(n_0947_)
	);

	and_bi n_1681_ (
		.a(n_0946_),
		.b(n_0947_),
		.c(n_0948_)
	);

	and_bb n_1682_ (
		.a(new_net_122),
		.b(new_net_513),
		.c(n_0949_)
	);

	and_ii n_1683_ (
		.a(new_net_1257),
		.b(new_net_253),
		.c(n_0950_)
	);

	and_ii n_1684_ (
		.a(new_net_1428),
		.b(new_net_2284),
		.c(n_0951_)
	);

	and_bi n_1685_ (
		.a(new_net_2285),
		.b(new_net_160),
		.c(n_0952_)
	);

	and_bi n_1686_ (
		.a(new_net_242),
		.b(new_net_363),
		.c(n_0953_)
	);

	and_ii n_1687_ (
		.a(n_0953_),
		.b(n_0952_),
		.c(n_0954_)
	);

	and_bi n_1688_ (
		.a(new_net_1445),
		.b(new_net_1288),
		.c(n_0955_)
	);

	and_bi n_1689_ (
		.a(new_net_1289),
		.b(new_net_1446),
		.c(n_0956_)
	);

	and_ii n_1690_ (
		.a(n_0956_),
		.b(n_0955_),
		.c(n_0957_)
	);

	and_bi n_1691_ (
		.a(new_net_2286),
		.b(new_net_144),
		.c(n_0958_)
	);

	and_bi n_1692_ (
		.a(new_net_230),
		.b(new_net_1357),
		.c(n_0959_)
	);

	and_ii n_1693_ (
		.a(n_0959_),
		.b(n_0958_),
		.c(n_0960_)
	);

	and_bi n_1694_ (
		.a(new_net_2287),
		.b(new_net_138),
		.c(n_0961_)
	);

	and_bi n_1695_ (
		.a(new_net_227),
		.b(new_net_1332),
		.c(n_0962_)
	);

	and_ii n_1696_ (
		.a(n_0962_),
		.b(n_0961_),
		.c(n_0963_)
	);

	and_ii n_1697_ (
		.a(new_net_422),
		.b(new_net_1947),
		.c(n_0964_)
	);

	and_bb n_1698_ (
		.a(new_net_425),
		.b(new_net_1950),
		.c(n_0965_)
	);

	and_ii n_1699_ (
		.a(n_0965_),
		.b(n_0964_),
		.c(n_0966_)
	);

	and_bi n_1700_ (
		.a(new_net_1588),
		.b(new_net_1749),
		.c(n_0967_)
	);

	and_bi n_1701_ (
		.a(new_net_1750),
		.b(new_net_1589),
		.c(n_0968_)
	);

	or_bb n_1702_ (
		.a(n_0968_),
		.b(n_0967_),
		.c(n_0969_)
	);

	and_bi n_1703_ (
		.a(new_net_2288),
		.b(new_net_145),
		.c(n_0970_)
	);

	and_bi n_1704_ (
		.a(new_net_231),
		.b(new_net_1349),
		.c(n_0971_)
	);

	and_ii n_1705_ (
		.a(n_0971_),
		.b(n_0970_),
		.c(n_0972_)
	);

	and_bi n_1706_ (
		.a(new_net_2289),
		.b(new_net_139),
		.c(n_0973_)
	);

	and_bi n_1707_ (
		.a(new_net_228),
		.b(new_net_1479),
		.c(n_0974_)
	);

	and_ii n_1708_ (
		.a(n_0974_),
		.b(n_0973_),
		.c(n_0975_)
	);

	and_bi n_1709_ (
		.a(new_net_1885),
		.b(new_net_1925),
		.c(n_0976_)
	);

	and_bi n_1710_ (
		.a(new_net_1928),
		.b(new_net_1886),
		.c(n_0977_)
	);

	and_ii n_1711_ (
		.a(n_0977_),
		.b(n_0976_),
		.c(n_0978_)
	);

	and_bi n_1712_ (
		.a(new_net_2290),
		.b(new_net_153),
		.c(n_0979_)
	);

	and_bi n_1713_ (
		.a(new_net_233),
		.b(new_net_1225),
		.c(n_0980_)
	);

	and_ii n_1714_ (
		.a(n_0980_),
		.b(n_0979_),
		.c(n_0981_)
	);

	and_bi n_1715_ (
		.a(new_net_45),
		.b(new_net_764),
		.c(n_0982_)
	);

	and_bi n_1716_ (
		.a(new_net_766),
		.b(new_net_46),
		.c(n_0983_)
	);

	or_bb n_1717_ (
		.a(n_0983_),
		.b(n_0982_),
		.c(n_0984_)
	);

	and_bi n_1718_ (
		.a(new_net_2291),
		.b(new_net_140),
		.c(n_0985_)
	);

	and_bi n_1719_ (
		.a(new_net_229),
		.b(new_net_1389),
		.c(n_0986_)
	);

	and_ii n_1720_ (
		.a(n_0986_),
		.b(n_0985_),
		.c(n_0987_)
	);

	and_bi n_1721_ (
		.a(new_net_2292),
		.b(new_net_161),
		.c(n_0988_)
	);

	and_bi n_1722_ (
		.a(new_net_243),
		.b(new_net_1080),
		.c(n_0989_)
	);

	and_ii n_1723_ (
		.a(n_0989_),
		.b(n_0988_),
		.c(n_0990_)
	);

	and_bi n_1724_ (
		.a(new_net_2293),
		.b(new_net_154),
		.c(n_0991_)
	);

	and_bi n_1725_ (
		.a(new_net_234),
		.b(new_net_1432),
		.c(n_0992_)
	);

	and_ii n_1726_ (
		.a(n_0992_),
		.b(n_0991_),
		.c(n_0993_)
	);

	and_ii n_1727_ (
		.a(new_net_41),
		.b(new_net_488),
		.c(n_0994_)
	);

	and_bb n_1728_ (
		.a(new_net_44),
		.b(new_net_491),
		.c(n_0995_)
	);

	or_bb n_1729_ (
		.a(n_0995_),
		.b(n_0994_),
		.c(n_0996_)
	);

	or_bb n_1730_ (
		.a(new_net_628),
		.b(new_net_1392),
		.c(n_0997_)
	);

	or_ii n_1731_ (
		.a(new_net_629),
		.b(new_net_1395),
		.c(n_0998_)
	);

	and_bb n_1732_ (
		.a(n_0998_),
		.b(n_0997_),
		.c(n_0999_)
	);

	and_bi n_1733_ (
		.a(new_net_694),
		.b(new_net_299),
		.c(n_1000_)
	);

	and_bi n_1734_ (
		.a(new_net_300),
		.b(new_net_695),
		.c(n_1001_)
	);

	and_ii n_1735_ (
		.a(n_1001_),
		.b(n_1000_),
		.c(n_1002_)
	);

	or_bb n_1736_ (
		.a(new_net_754),
		.b(new_net_1803),
		.c(n_1003_)
	);

	and_bb n_1737_ (
		.a(new_net_755),
		.b(new_net_1804),
		.c(n_1004_)
	);

	and_bi n_1738_ (
		.a(n_1003_),
		.b(n_1004_),
		.c(n_1005_)
	);

	or_bb n_1739_ (
		.a(n_1005_),
		.b(new_net_2294),
		.c(n_1006_)
	);

	and_bi n_1740_ (
		.a(new_net_2295),
		.b(new_net_261),
		.c(n_1007_)
	);

	and_bi n_1741_ (
		.a(new_net_168),
		.b(new_net_1607),
		.c(n_1008_)
	);

	and_ii n_1742_ (
		.a(n_1008_),
		.b(n_1007_),
		.c(n_1009_)
	);

	and_bi n_1743_ (
		.a(new_net_2296),
		.b(new_net_254),
		.c(n_1010_)
	);

	and_bi n_1744_ (
		.a(new_net_165),
		.b(new_net_1659),
		.c(n_1011_)
	);

	and_ii n_1745_ (
		.a(n_1011_),
		.b(n_1010_),
		.c(n_1012_)
	);

	or_bb n_1746_ (
		.a(new_net_974),
		.b(new_net_1929),
		.c(n_1013_)
	);

	and_bb n_1747_ (
		.a(new_net_977),
		.b(new_net_1931),
		.c(n_1014_)
	);

	and_bi n_1748_ (
		.a(n_1013_),
		.b(n_1014_),
		.c(n_1015_)
	);

	and_bi n_1749_ (
		.a(new_net_2297),
		.b(new_net_272),
		.c(n_1016_)
	);

	and_bi n_1750_ (
		.a(new_net_174),
		.b(new_net_1719),
		.c(n_1017_)
	);

	and_ii n_1751_ (
		.a(n_1017_),
		.b(n_1016_),
		.c(n_1018_)
	);

	and_bi n_1752_ (
		.a(new_net_2298),
		.b(new_net_262),
		.c(n_1019_)
	);

	and_bi n_1753_ (
		.a(new_net_169),
		.b(new_net_849),
		.c(n_1020_)
	);

	and_ii n_1754_ (
		.a(n_1020_),
		.b(n_1019_),
		.c(n_1021_)
	);

	and_bi n_1755_ (
		.a(new_net_1244),
		.b(new_net_1147),
		.c(n_1022_)
	);

	and_bi n_1756_ (
		.a(new_net_1150),
		.b(new_net_1245),
		.c(n_1023_)
	);

	and_ii n_1757_ (
		.a(n_1023_),
		.b(n_1022_),
		.c(n_1024_)
	);

	or_bi n_1758_ (
		.a(new_net_1024),
		.b(new_net_1900),
		.c(n_1025_)
	);

	and_bi n_1759_ (
		.a(new_net_1025),
		.b(new_net_1901),
		.c(n_1026_)
	);

	and_bi n_1760_ (
		.a(n_1025_),
		.b(n_1026_),
		.c(n_1027_)
	);

	and_bi n_1761_ (
		.a(new_net_2299),
		.b(new_net_273),
		.c(n_1028_)
	);

	and_bi n_1762_ (
		.a(new_net_175),
		.b(new_net_1579),
		.c(n_1029_)
	);

	and_ii n_1763_ (
		.a(n_1029_),
		.b(n_1028_),
		.c(n_1030_)
	);

	and_bi n_1764_ (
		.a(new_net_2300),
		.b(new_net_263),
		.c(n_1031_)
	);

	and_bi n_1765_ (
		.a(new_net_170),
		.b(new_net_1895),
		.c(n_1032_)
	);

	and_ii n_1766_ (
		.a(n_1032_),
		.b(n_1031_),
		.c(n_1033_)
	);

	and_ii n_1767_ (
		.a(new_net_1089),
		.b(new_net_748),
		.c(n_1034_)
	);

	and_bb n_1768_ (
		.a(new_net_1091),
		.b(new_net_749),
		.c(n_1035_)
	);

	and_ii n_1769_ (
		.a(n_1035_),
		.b(n_1034_),
		.c(n_1036_)
	);

	or_bi n_1770_ (
		.a(new_net_402),
		.b(new_net_1371),
		.c(n_1037_)
	);

	and_bi n_1771_ (
		.a(new_net_403),
		.b(new_net_1372),
		.c(n_1038_)
	);

	and_bi n_1772_ (
		.a(n_1037_),
		.b(n_1038_),
		.c(n_1039_)
	);

	and_bi n_1773_ (
		.a(new_net_2301),
		.b(new_net_274),
		.c(n_1040_)
	);

	and_bi n_1774_ (
		.a(new_net_176),
		.b(new_net_519),
		.c(n_1041_)
	);

	and_ii n_1775_ (
		.a(n_1041_),
		.b(n_1040_),
		.c(n_1042_)
	);

	and_bi n_1776_ (
		.a(new_net_2302),
		.b(new_net_264),
		.c(n_1043_)
	);

	and_bi n_1777_ (
		.a(new_net_171),
		.b(new_net_650),
		.c(n_1044_)
	);

	and_ii n_1778_ (
		.a(n_1044_),
		.b(n_1043_),
		.c(n_1045_)
	);

	and_ii n_1779_ (
		.a(new_net_524),
		.b(new_net_1601),
		.c(n_1046_)
	);

	and_bb n_1780_ (
		.a(new_net_527),
		.b(new_net_1602),
		.c(n_1047_)
	);

	and_ii n_1781_ (
		.a(n_1047_),
		.b(n_1046_),
		.c(n_1048_)
	);

	and_bi n_1782_ (
		.a(new_net_2303),
		.b(new_net_285),
		.c(n_1049_)
	);

	and_bi n_1783_ (
		.a(new_net_186),
		.b(new_net_1590),
		.c(n_1050_)
	);

	and_ii n_1784_ (
		.a(n_1050_),
		.b(n_1049_),
		.c(n_1051_)
	);

	and_bi n_1785_ (
		.a(new_net_2304),
		.b(new_net_275),
		.c(n_1052_)
	);

	and_bi n_1786_ (
		.a(new_net_177),
		.b(new_net_1560),
		.c(n_1053_)
	);

	and_ii n_1787_ (
		.a(n_1053_),
		.b(n_1052_),
		.c(n_1054_)
	);

	and_ii n_1788_ (
		.a(new_net_1488),
		.b(new_net_1162),
		.c(n_1055_)
	);

	and_bb n_1789_ (
		.a(new_net_1491),
		.b(new_net_1163),
		.c(n_1056_)
	);

	and_ii n_1790_ (
		.a(n_1056_),
		.b(n_1055_),
		.c(n_1057_)
	);

	and_ii n_1791_ (
		.a(new_net_1780),
		.b(new_net_1713),
		.c(n_1058_)
	);

	and_bb n_1792_ (
		.a(new_net_1781),
		.b(new_net_1714),
		.c(n_1059_)
	);

	and_ii n_1793_ (
		.a(n_1059_),
		.b(n_1058_),
		.c(n_1060_)
	);

	or_bb n_1794_ (
		.a(new_net_1376),
		.b(new_net_1690),
		.c(n_1061_)
	);

	and_bb n_1795_ (
		.a(new_net_1377),
		.b(new_net_1691),
		.c(n_1062_)
	);

	and_bi n_1796_ (
		.a(n_1061_),
		.b(n_1062_),
		.c(n_1063_)
	);

	and_bi n_1797_ (
		.a(new_net_2305),
		.b(new_net_276),
		.c(n_1064_)
	);

	and_bi n_1798_ (
		.a(new_net_178),
		.b(new_net_1457),
		.c(n_1065_)
	);

	and_ii n_1799_ (
		.a(n_1065_),
		.b(n_1064_),
		.c(n_1066_)
	);

	and_bi n_1800_ (
		.a(new_net_2306),
		.b(new_net_265),
		.c(n_1067_)
	);

	and_bi n_1801_ (
		.a(new_net_172),
		.b(new_net_1575),
		.c(n_1068_)
	);

	and_ii n_1802_ (
		.a(n_1068_),
		.b(n_1067_),
		.c(n_1069_)
	);

	or_bb n_1803_ (
		.a(new_net_538),
		.b(new_net_1196),
		.c(n_1070_)
	);

	and_bb n_1804_ (
		.a(new_net_541),
		.b(new_net_1197),
		.c(n_1071_)
	);

	and_bi n_1805_ (
		.a(n_1070_),
		.b(n_1071_),
		.c(n_1072_)
	);

	and_bi n_1806_ (
		.a(new_net_2307),
		.b(new_net_286),
		.c(n_1073_)
	);

	and_bi n_1807_ (
		.a(new_net_187),
		.b(new_net_1233),
		.c(n_1074_)
	);

	and_ii n_1808_ (
		.a(n_1074_),
		.b(n_1073_),
		.c(n_1075_)
	);

	and_bi n_1809_ (
		.a(new_net_2308),
		.b(new_net_277),
		.c(n_1076_)
	);

	and_bi n_1810_ (
		.a(new_net_179),
		.b(new_net_1266),
		.c(n_1077_)
	);

	and_ii n_1811_ (
		.a(n_1077_),
		.b(n_1076_),
		.c(n_1078_)
	);

	or_bi n_1812_ (
		.a(new_net_1492),
		.b(new_net_1409),
		.c(n_1079_)
	);

	and_bi n_1813_ (
		.a(new_net_1495),
		.b(new_net_1410),
		.c(n_1080_)
	);

	and_bi n_1814_ (
		.a(n_1079_),
		.b(n_1080_),
		.c(n_1081_)
	);

	and_ii n_1815_ (
		.a(new_net_1545),
		.b(new_net_864),
		.c(n_1082_)
	);

	and_bb n_1816_ (
		.a(new_net_1546),
		.b(new_net_865),
		.c(n_1083_)
	);

	and_ii n_1817_ (
		.a(n_1083_),
		.b(n_1082_),
		.c(n_1084_)
	);

	and_bi n_1818_ (
		.a(new_net_2309),
		.b(new_net_287),
		.c(n_1085_)
	);

	and_bi n_1819_ (
		.a(new_net_188),
		.b(new_net_1067),
		.c(n_1086_)
	);

	and_ii n_1820_ (
		.a(n_1086_),
		.b(n_1085_),
		.c(n_1087_)
	);

	and_bi n_1821_ (
		.a(new_net_2310),
		.b(new_net_278),
		.c(n_1088_)
	);

	and_bi n_1822_ (
		.a(new_net_180),
		.b(new_net_1144),
		.c(n_1089_)
	);

	and_ii n_1823_ (
		.a(n_1089_),
		.b(n_1088_),
		.c(n_1090_)
	);

	and_bi n_1824_ (
		.a(new_net_1648),
		.b(new_net_980),
		.c(n_1091_)
	);

	and_bi n_1825_ (
		.a(new_net_983),
		.b(new_net_1649),
		.c(n_1092_)
	);

	and_ii n_1826_ (
		.a(n_1092_),
		.b(n_1091_),
		.c(n_1093_)
	);

	and_bi n_1827_ (
		.a(new_net_2311),
		.b(new_net_255),
		.c(n_1094_)
	);

	and_bi n_1828_ (
		.a(new_net_166),
		.b(new_net_1340),
		.c(n_1095_)
	);

	and_ii n_1829_ (
		.a(n_1095_),
		.b(n_1094_),
		.c(n_1096_)
	);

	or_ii n_1830_ (
		.a(new_net_1824),
		.b(new_net_1769),
		.c(n_1097_)
	);

	or_bb n_1831_ (
		.a(new_net_1825),
		.b(new_net_1770),
		.c(n_1098_)
	);

	or_ii n_1832_ (
		.a(n_1098_),
		.b(n_1097_),
		.c(n_1099_)
	);

	and_bi n_1833_ (
		.a(new_net_2312),
		.b(new_net_155),
		.c(n_1100_)
	);

	and_bi n_1834_ (
		.a(new_net_181),
		.b(new_net_1765),
		.c(n_1101_)
	);

	and_ii n_1835_ (
		.a(n_1101_),
		.b(n_1100_),
		.c(n_1102_)
	);

	and_bi n_1836_ (
		.a(new_net_2313),
		.b(new_net_266),
		.c(n_1103_)
	);

	and_bi n_1837_ (
		.a(new_net_173),
		.b(new_net_1877),
		.c(n_1104_)
	);

	and_ii n_1838_ (
		.a(n_1104_),
		.b(n_1103_),
		.c(n_1105_)
	);

	and_bi n_1839_ (
		.a(new_net_637),
		.b(new_net_63),
		.c(n_1106_)
	);

	and_bi n_1840_ (
		.a(new_net_65),
		.b(new_net_638),
		.c(n_1107_)
	);

	and_ii n_1841_ (
		.a(n_1107_),
		.b(n_1106_),
		.c(n_1108_)
	);

	and_bi n_1842_ (
		.a(new_net_2314),
		.b(new_net_288),
		.c(n_1109_)
	);

	and_bi n_1843_ (
		.a(new_net_189),
		.b(new_net_1122),
		.c(n_1110_)
	);

	and_ii n_1844_ (
		.a(n_1110_),
		.b(n_1109_),
		.c(n_1111_)
	);

	or_bb n_1845_ (
		.a(new_net_319),
		.b(new_net_110),
		.c(n_1112_)
	);

	or_ii n_1846_ (
		.a(new_net_322),
		.b(new_net_111),
		.c(n_1113_)
	);

	or_ii n_1847_ (
		.a(n_1113_),
		.b(n_1112_),
		.c(n_1114_)
	);

	and_ii n_1848_ (
		.a(new_net_1872),
		.b(new_net_1909),
		.c(n_1115_)
	);

	and_bb n_1849_ (
		.a(new_net_1873),
		.b(new_net_1910),
		.c(n_1116_)
	);

	and_ii n_1850_ (
		.a(n_1116_),
		.b(n_1115_),
		.c(n_1117_)
	);

	and_bi n_1851_ (
		.a(new_net_358),
		.b(new_net_1599),
		.c(n_1118_)
	);

	and_bi n_1852_ (
		.a(new_net_1600),
		.b(new_net_359),
		.c(n_1119_)
	);

	or_bb n_1853_ (
		.a(n_1119_),
		.b(n_1118_),
		.c(n_1120_)
	);

	or_bb n_1854_ (
		.a(n_1120_),
		.b(n_1063_),
		.c(n_1121_)
	);

	or_bb n_1855_ (
		.a(n_1121_),
		.b(n_1006_),
		.c(new_net_6)
	);

	and_ii n_1856_ (
		.a(new_net_1018),
		.b(new_net_2315),
		.c(n_1122_)
	);

	and_bi n_1857_ (
		.a(new_net_235),
		.b(new_net_2316),
		.c(n_1123_)
	);

	and_ii n_1858_ (
		.a(new_net_659),
		.b(new_net_388),
		.c(n_1124_)
	);

	and_bi n_1859_ (
		.a(new_net_124),
		.b(new_net_2317),
		.c(n_1125_)
	);

	and_bb n_1860_ (
		.a(new_net_684),
		.b(new_net_666),
		.c(n_1126_)
	);

	or_bb n_1861_ (
		.a(new_net_685),
		.b(new_net_384),
		.c(n_1127_)
	);

	and_bi n_1862_ (
		.a(new_net_660),
		.b(new_net_1461),
		.c(n_1128_)
	);

	and_ii n_1863_ (
		.a(n_1128_),
		.b(n_1126_),
		.c(n_1129_)
	);

	and_ii n_1864_ (
		.a(new_net_1672),
		.b(new_net_626),
		.c(n_1130_)
	);

	and_bb n_1865_ (
		.a(new_net_1673),
		.b(new_net_627),
		.c(n_1131_)
	);

	or_bb n_1866_ (
		.a(n_1131_),
		.b(n_1130_),
		.c(n_1132_)
	);

	and_bi n_1867_ (
		.a(new_net_190),
		.b(new_net_2318),
		.c(n_1133_)
	);

	and_ii n_1868_ (
		.a(new_net_856),
		.b(new_net_380),
		.c(n_1134_)
	);

	and_bi n_1869_ (
		.a(new_net_236),
		.b(new_net_2319),
		.c(n_1135_)
	);

	and_bb n_1870_ (
		.a(new_net_515),
		.b(new_net_365),
		.c(n_1136_)
	);

	and_ii n_1871_ (
		.a(new_net_516),
		.b(new_net_371),
		.c(n_1137_)
	);

	and_bb n_1872_ (
		.a(new_net_741),
		.b(new_net_857),
		.c(n_1138_)
	);

	and_ii n_1873_ (
		.a(n_1138_),
		.b(n_1136_),
		.c(n_1139_)
	);

	or_bi n_1874_ (
		.a(new_net_551),
		.b(new_net_1775),
		.c(n_1140_)
	);

	and_bi n_1875_ (
		.a(new_net_552),
		.b(new_net_1776),
		.c(n_1141_)
	);

	and_bi n_1876_ (
		.a(n_1140_),
		.b(n_1141_),
		.c(n_1142_)
	);

	and_ii n_1877_ (
		.a(new_net_2320),
		.b(new_net_1019),
		.c(n_1143_)
	);

	and_bi n_1878_ (
		.a(new_net_954),
		.b(new_net_1549),
		.c(n_1144_)
	);

	and_bi n_1879_ (
		.a(new_net_1550),
		.b(new_net_955),
		.c(n_1145_)
	);

	and_ii n_1880_ (
		.a(n_1145_),
		.b(n_1144_),
		.c(n_1146_)
	);

	or_bb n_1881_ (
		.a(new_net_1834),
		.b(new_net_839),
		.c(n_1147_)
	);

	and_bb n_1882_ (
		.a(new_net_1835),
		.b(new_net_840),
		.c(n_1148_)
	);

	and_bi n_1883_ (
		.a(n_1147_),
		.b(n_1148_),
		.c(n_1149_)
	);

	and_bb n_1884_ (
		.a(new_net_2321),
		.b(new_net_267),
		.c(n_1150_)
	);

	and_ii n_1885_ (
		.a(new_net_2322),
		.b(new_net_434),
		.c(n_1151_)
	);

	and_bb n_1886_ (
		.a(new_net_2323),
		.b(new_net_141),
		.c(n_1152_)
	);

	and_ii n_1887_ (
		.a(new_net_2324),
		.b(new_net_328),
		.c(n_1153_)
	);

	and_ii n_1888_ (
		.a(new_net_822),
		.b(new_net_611),
		.c(n_1154_)
	);

	and_bb n_1889_ (
		.a(new_net_823),
		.b(new_net_613),
		.c(n_1155_)
	);

	and_ii n_1890_ (
		.a(n_1155_),
		.b(n_1154_),
		.c(n_1156_)
	);

	and_bb n_1891_ (
		.a(new_net_2325),
		.b(new_net_222),
		.c(n_1157_)
	);

	and_ii n_1892_ (
		.a(new_net_2326),
		.b(new_net_775),
		.c(n_1158_)
	);

	and_bb n_1893_ (
		.a(new_net_2327),
		.b(new_net_201),
		.c(n_1159_)
	);

	and_ii n_1894_ (
		.a(new_net_2328),
		.b(new_net_842),
		.c(n_1160_)
	);

	and_bi n_1895_ (
		.a(new_net_1320),
		.b(new_net_1551),
		.c(n_1161_)
	);

	and_bi n_1896_ (
		.a(new_net_1553),
		.b(new_net_1323),
		.c(n_1162_)
	);

	and_ii n_1897_ (
		.a(n_1162_),
		.b(n_1161_),
		.c(n_1163_)
	);

	and_bb n_1898_ (
		.a(new_net_2329),
		.b(new_net_142),
		.c(n_1164_)
	);

	and_ii n_1899_ (
		.a(new_net_2330),
		.b(new_net_973),
		.c(n_1165_)
	);

	and_bb n_1900_ (
		.a(new_net_2331),
		.b(new_net_202),
		.c(n_1166_)
	);

	and_ii n_1901_ (
		.a(new_net_2332),
		.b(new_net_1027),
		.c(n_1167_)
	);

	and_ii n_1902_ (
		.a(new_net_497),
		.b(new_net_87),
		.c(n_1168_)
	);

	and_bb n_1903_ (
		.a(new_net_499),
		.b(new_net_88),
		.c(n_1169_)
	);

	and_ii n_1904_ (
		.a(n_1169_),
		.b(n_1168_),
		.c(n_1170_)
	);

	and_bb n_1905_ (
		.a(new_net_829),
		.b(new_net_1839),
		.c(n_1171_)
	);

	and_ii n_1906_ (
		.a(new_net_830),
		.b(new_net_1840),
		.c(n_1172_)
	);

	and_ii n_1907_ (
		.a(n_1172_),
		.b(n_1171_),
		.c(n_1173_)
	);

	and_bi n_1908_ (
		.a(new_net_1130),
		.b(new_net_1132),
		.c(n_1174_)
	);

	and_bi n_1909_ (
		.a(new_net_1133),
		.b(new_net_1131),
		.c(n_1175_)
	);

	and_ii n_1910_ (
		.a(n_1175_),
		.b(n_1174_),
		.c(n_1176_)
	);

	and_bb n_1911_ (
		.a(new_net_2333),
		.b(new_net_256),
		.c(n_1177_)
	);

	and_ii n_1912_ (
		.a(new_net_2334),
		.b(new_net_1920),
		.c(n_1178_)
	);

	and_bb n_1913_ (
		.a(new_net_2335),
		.b(new_net_162),
		.c(n_1179_)
	);

	and_ii n_1914_ (
		.a(new_net_2336),
		.b(new_net_1620),
		.c(n_1180_)
	);

	and_ii n_1915_ (
		.a(new_net_1851),
		.b(new_net_1663),
		.c(n_1181_)
	);

	and_bb n_1916_ (
		.a(new_net_1853),
		.b(new_net_1665),
		.c(n_1182_)
	);

	and_ii n_1917_ (
		.a(n_1182_),
		.b(n_1181_),
		.c(n_1183_)
	);

	and_bb n_1918_ (
		.a(new_net_2337),
		.b(new_net_215),
		.c(n_1184_)
	);

	and_ii n_1919_ (
		.a(new_net_2338),
		.b(new_net_1727),
		.c(n_1185_)
	);

	and_bb n_1920_ (
		.a(new_net_2339),
		.b(new_net_182),
		.c(n_1186_)
	);

	and_ii n_1921_ (
		.a(new_net_2340),
		.b(new_net_68),
		.c(n_1187_)
	);

	and_bb n_1922_ (
		.a(new_net_1845),
		.b(new_net_1096),
		.c(n_1188_)
	);

	and_ii n_1923_ (
		.a(new_net_1847),
		.b(new_net_1097),
		.c(n_1189_)
	);

	and_ii n_1924_ (
		.a(n_1189_),
		.b(n_1188_),
		.c(n_1190_)
	);

	and_bi n_1925_ (
		.a(new_net_342),
		.b(new_net_344),
		.c(n_1191_)
	);

	and_bi n_1926_ (
		.a(new_net_345),
		.b(new_net_343),
		.c(n_1192_)
	);

	and_ii n_1927_ (
		.a(n_1192_),
		.b(n_1191_),
		.c(n_1193_)
	);

	and_bi n_1928_ (
		.a(new_net_1209),
		.b(new_net_1437),
		.c(n_1194_)
	);

	and_bi n_1929_ (
		.a(new_net_1438),
		.b(new_net_1210),
		.c(n_1195_)
	);

	or_bb n_1930_ (
		.a(n_1195_),
		.b(n_1194_),
		.c(n_1196_)
	);

	or_bb n_1931_ (
		.a(n_1196_),
		.b(new_net_2341),
		.c(n_1197_)
	);

	and_bb n_1932_ (
		.a(new_net_2342),
		.b(new_net_131),
		.c(n_1198_)
	);

	and_ii n_1933_ (
		.a(new_net_2343),
		.b(new_net_339),
		.c(n_1199_)
	);

	and_bb n_1934_ (
		.a(new_net_2344),
		.b(new_net_244),
		.c(n_1200_)
	);

	and_ii n_1935_ (
		.a(new_net_2345),
		.b(new_net_722),
		.c(n_1201_)
	);

	and_bi n_1936_ (
		.a(new_net_1364),
		.b(new_net_1401),
		.c(n_1202_)
	);

	and_bi n_1937_ (
		.a(new_net_1402),
		.b(new_net_1365),
		.c(n_1203_)
	);

	or_bb n_1938_ (
		.a(n_1203_),
		.b(n_1202_),
		.c(n_1204_)
	);

	and_bi n_1939_ (
		.a(new_net_191),
		.b(new_net_2346),
		.c(n_1205_)
	);

	and_ii n_1940_ (
		.a(new_net_1507),
		.b(new_net_381),
		.c(n_1206_)
	);

	and_bi n_1941_ (
		.a(new_net_237),
		.b(new_net_2347),
		.c(n_1207_)
	);

	and_bb n_1942_ (
		.a(new_net_346),
		.b(new_net_1515),
		.c(n_1208_)
	);

	and_ii n_1943_ (
		.a(new_net_347),
		.b(new_net_372),
		.c(n_1209_)
	);

	and_bb n_1944_ (
		.a(new_net_617),
		.b(new_net_1508),
		.c(n_1210_)
	);

	and_ii n_1945_ (
		.a(n_1210_),
		.b(n_1208_),
		.c(n_1211_)
	);

	and_bi n_1946_ (
		.a(new_net_123),
		.b(new_net_2348),
		.c(n_1212_)
	);

	and_ii n_1947_ (
		.a(new_net_936),
		.b(new_net_376),
		.c(n_1213_)
	);

	and_bi n_1948_ (
		.a(new_net_167),
		.b(new_net_2349),
		.c(n_1214_)
	);

	and_bb n_1949_ (
		.a(new_net_1142),
		.b(new_net_1041),
		.c(n_1215_)
	);

	and_ii n_1950_ (
		.a(new_net_1143),
		.b(new_net_390),
		.c(n_1216_)
	);

	and_bb n_1951_ (
		.a(new_net_1333),
		.b(new_net_937),
		.c(n_1217_)
	);

	and_ii n_1952_ (
		.a(n_1217_),
		.b(n_1215_),
		.c(n_1218_)
	);

	and_bb n_1953_ (
		.a(new_net_1568),
		.b(new_net_833),
		.c(n_1219_)
	);

	and_ii n_1954_ (
		.a(new_net_1569),
		.b(new_net_834),
		.c(n_1220_)
	);

	or_bb n_1955_ (
		.a(n_1220_),
		.b(n_1219_),
		.c(n_1221_)
	);

	and_ii n_1956_ (
		.a(new_net_1863),
		.b(new_net_1855),
		.c(n_1222_)
	);

	and_bb n_1957_ (
		.a(new_net_1864),
		.b(new_net_1856),
		.c(n_1223_)
	);

	and_ii n_1958_ (
		.a(n_1223_),
		.b(n_1222_),
		.c(n_1224_)
	);

	and_bb n_1959_ (
		.a(new_net_2350),
		.b(new_net_257),
		.c(n_1225_)
	);

	and_ii n_1960_ (
		.a(new_net_2351),
		.b(new_net_716),
		.c(n_1226_)
	);

	and_bi n_1961_ (
		.a(new_net_129),
		.b(new_net_2352),
		.c(n_1227_)
	);

	and_ii n_1962_ (
		.a(n_1227_),
		.b(new_net_391),
		.c(n_1228_)
	);

	and_ii n_1963_ (
		.a(new_net_1013),
		.b(new_net_622),
		.c(n_1229_)
	);

	and_bb n_1964_ (
		.a(new_net_1014),
		.b(new_net_625),
		.c(n_1230_)
	);

	and_ii n_1965_ (
		.a(n_1230_),
		.b(n_1229_),
		.c(n_1231_)
	);

	and_bb n_1966_ (
		.a(new_net_2353),
		.b(new_net_216),
		.c(n_1232_)
	);

	and_ii n_1967_ (
		.a(new_net_2354),
		.b(new_net_872),
		.c(n_1233_)
	);

	and_bb n_1968_ (
		.a(new_net_2355),
		.b(new_net_268),
		.c(n_1234_)
	);

	and_ii n_1969_ (
		.a(new_net_2356),
		.b(new_net_939),
		.c(n_1235_)
	);

	and_ii n_1970_ (
		.a(new_net_1741),
		.b(new_net_94),
		.c(n_1236_)
	);

	and_bb n_1971_ (
		.a(new_net_1742),
		.b(new_net_97),
		.c(n_1237_)
	);

	and_ii n_1972_ (
		.a(n_1237_),
		.b(n_1236_),
		.c(n_1238_)
	);

	and_bi n_1973_ (
		.a(new_net_73),
		.b(new_net_54),
		.c(n_1239_)
	);

	and_bi n_1974_ (
		.a(new_net_55),
		.b(new_net_74),
		.c(n_1240_)
	);

	and_ii n_1975_ (
		.a(n_1240_),
		.b(n_1239_),
		.c(n_1241_)
	);

	and_bi n_1976_ (
		.a(new_net_348),
		.b(new_net_591),
		.c(n_1242_)
	);

	and_bi n_1977_ (
		.a(new_net_592),
		.b(new_net_349),
		.c(n_1243_)
	);

	or_bb n_1978_ (
		.a(n_1243_),
		.b(n_1242_),
		.c(n_1244_)
	);

	and_bb n_1979_ (
		.a(new_net_2357),
		.b(new_net_146),
		.c(n_1245_)
	);

	and_ii n_1980_ (
		.a(new_net_2358),
		.b(new_net_1317),
		.c(n_1246_)
	);

	and_bb n_1981_ (
		.a(new_net_2359),
		.b(new_net_207),
		.c(n_1247_)
	);

	and_bi n_1982_ (
		.a(new_net_643),
		.b(new_net_2360),
		.c(n_1248_)
	);

	and_bb n_1983_ (
		.a(new_net_1312),
		.b(new_net_1126),
		.c(n_1249_)
	);

	and_ii n_1984_ (
		.a(new_net_1313),
		.b(new_net_1127),
		.c(n_1250_)
	);

	and_ii n_1985_ (
		.a(n_1250_),
		.b(n_1249_),
		.c(n_1251_)
	);

	and_bb n_1986_ (
		.a(new_net_2361),
		.b(new_net_223),
		.c(n_1252_)
	);

	and_ii n_1987_ (
		.a(new_net_2362),
		.b(new_net_846),
		.c(n_1253_)
	);

	and_bb n_1988_ (
		.a(new_net_2363),
		.b(new_net_156),
		.c(n_1254_)
	);

	and_ii n_1989_ (
		.a(new_net_2364),
		.b(new_net_1105),
		.c(n_1255_)
	);

	and_ii n_1990_ (
		.a(new_net_770),
		.b(new_net_729),
		.c(n_1256_)
	);

	and_bb n_1991_ (
		.a(new_net_771),
		.b(new_net_731),
		.c(n_1257_)
	);

	and_ii n_1992_ (
		.a(n_1257_),
		.b(n_1256_),
		.c(n_1258_)
	);

	and_bb n_1993_ (
		.a(new_net_2365),
		.b(new_net_208),
		.c(n_1259_)
	);

	and_ii n_1994_ (
		.a(new_net_2366),
		.b(new_net_1890),
		.c(n_1260_)
	);

	and_bb n_1995_ (
		.a(new_net_2367),
		.b(new_net_163),
		.c(n_1261_)
	);

	and_ii n_1996_ (
		.a(new_net_2368),
		.b(new_net_1752),
		.c(n_1262_)
	);

	and_bi n_1997_ (
		.a(new_net_818),
		.b(new_net_926),
		.c(n_1263_)
	);

	and_bi n_1998_ (
		.a(new_net_929),
		.b(new_net_819),
		.c(n_1264_)
	);

	and_ii n_1999_ (
		.a(n_1264_),
		.b(n_1263_),
		.c(n_1265_)
	);

	and_bi n_2000_ (
		.a(new_net_992),
		.b(new_net_837),
		.c(n_1266_)
	);

	and_bi n_2001_ (
		.a(new_net_838),
		.b(new_net_993),
		.c(n_1267_)
	);

	and_ii n_2002_ (
		.a(n_1267_),
		.b(n_1266_),
		.c(n_1268_)
	);

	and_ii n_2003_ (
		.a(new_net_1646),
		.b(new_net_1644),
		.c(n_1269_)
	);

	and_bb n_2004_ (
		.a(new_net_1647),
		.b(new_net_1645),
		.c(n_1270_)
	);

	and_ii n_2005_ (
		.a(n_1270_),
		.b(n_1269_),
		.c(n_1271_)
	);

	and_bb n_2006_ (
		.a(new_net_2369),
		.b(new_net_245),
		.c(n_1272_)
	);

	and_ii n_2007_ (
		.a(new_net_2370),
		.b(new_net_1844),
		.c(n_1273_)
	);

	and_bb n_2008_ (
		.a(new_net_2371),
		.b(new_net_203),
		.c(n_1274_)
	);

	and_ii n_2009_ (
		.a(new_net_2372),
		.b(new_net_1159),
		.c(n_1275_)
	);

	and_bi n_2010_ (
		.a(new_net_557),
		.b(new_net_1178),
		.c(n_1276_)
	);

	and_bi n_2011_ (
		.a(new_net_1179),
		.b(new_net_560),
		.c(n_1277_)
	);

	and_ii n_2012_ (
		.a(n_1277_),
		.b(n_1276_),
		.c(n_1278_)
	);

	and_bb n_2013_ (
		.a(new_net_2373),
		.b(new_net_157),
		.c(n_1279_)
	);

	and_ii n_2014_ (
		.a(new_net_2374),
		.b(new_net_1414),
		.c(n_1280_)
	);

	and_bb n_2015_ (
		.a(new_net_2375),
		.b(new_net_147),
		.c(n_1281_)
	);

	and_ii n_2016_ (
		.a(new_net_2376),
		.b(new_net_711),
		.c(n_1282_)
	);

	and_ii n_2017_ (
		.a(new_net_1526),
		.b(new_net_1290),
		.c(n_1283_)
	);

	and_bb n_2018_ (
		.a(new_net_1527),
		.b(new_net_1292),
		.c(n_1284_)
	);

	and_ii n_2019_ (
		.a(n_1284_),
		.b(n_1283_),
		.c(n_1285_)
	);

	and_bi n_2020_ (
		.a(new_net_1231),
		.b(new_net_1407),
		.c(n_1286_)
	);

	and_bi n_2021_ (
		.a(new_net_1408),
		.b(new_net_1232),
		.c(n_1287_)
	);

	and_ii n_2022_ (
		.a(n_1287_),
		.b(n_1286_),
		.c(n_1288_)
	);

	and_bb n_2023_ (
		.a(new_net_1475),
		.b(new_net_295),
		.c(n_1289_)
	);

	and_ii n_2024_ (
		.a(new_net_1476),
		.b(new_net_296),
		.c(n_1290_)
	);

	or_bb n_2025_ (
		.a(n_1290_),
		.b(n_1289_),
		.c(n_1291_)
	);

	or_bb n_2026_ (
		.a(n_1291_),
		.b(n_1244_),
		.c(n_1292_)
	);

	or_bb n_2027_ (
		.a(n_1292_),
		.b(n_1197_),
		.c(new_net_5)
	);

	inv n_2028_ (
		.din(new_net_1146),
		.dout(n_1293_)
	);

	and_bi n_2029_ (
		.a(new_net_885),
		.b(new_net_487),
		.c(n_1294_)
	);

	and_bi n_2030_ (
		.a(new_net_486),
		.b(new_net_886),
		.c(n_1295_)
	);

	and_ii n_2031_ (
		.a(new_net_1108),
		.b(new_net_1002),
		.c(n_1296_)
	);

	inv n_2032_ (
		.din(new_net_850),
		.dout(n_1297_)
	);

	and_bi n_2033_ (
		.a(new_net_1294),
		.b(new_net_1300),
		.c(n_1298_)
	);

	and_bi n_2034_ (
		.a(new_net_1301),
		.b(new_net_1295),
		.c(n_1299_)
	);

	inv n_2035_ (
		.din(new_net_1720),
		.dout(n_1300_)
	);

	and_bi n_2036_ (
		.a(new_net_798),
		.b(new_net_1624),
		.c(n_1301_)
	);

	and_bi n_2037_ (
		.a(new_net_1625),
		.b(new_net_800),
		.c(n_1302_)
	);

	inv n_2038_ (
		.din(new_net_1815),
		.dout(n_1303_)
	);

	inv n_2039_ (
		.din(new_net_652),
		.dout(n_1304_)
	);

	and_bi n_2040_ (
		.a(new_net_1055),
		.b(new_net_1785),
		.c(n_1305_)
	);

	and_bi n_2041_ (
		.a(new_net_1786),
		.b(new_net_1054),
		.c(n_1306_)
	);

	inv n_2042_ (
		.din(new_net_520),
		.dout(n_1307_)
	);

	and_bi n_2043_ (
		.a(new_net_582),
		.b(new_net_1960),
		.c(n_1308_)
	);

	and_ii n_2044_ (
		.a(new_net_698),
		.b(new_net_448),
		.c(n_1309_)
	);

	and_ii n_2045_ (
		.a(new_net_803),
		.b(new_net_311),
		.c(n_1310_)
	);

	and_bi n_2046_ (
		.a(new_net_1953),
		.b(new_net_889),
		.c(n_1311_)
	);

	or_bb n_2047_ (
		.a(n_1311_),
		.b(new_net_1732),
		.c(n_1312_)
	);

	inv n_2048_ (
		.din(new_net_1733),
		.dout(n_1313_)
	);

	and_ii n_2049_ (
		.a(new_net_449),
		.b(new_net_312),
		.c(n_1314_)
	);

	and_bi n_2050_ (
		.a(new_net_1959),
		.b(new_net_583),
		.c(n_1315_)
	);

	or_bb n_2051_ (
		.a(new_net_1151),
		.b(new_net_699),
		.c(n_1316_)
	);

	and_bi n_2052_ (
		.a(new_net_1136),
		.b(new_net_1166),
		.c(n_1317_)
	);

	or_ii n_2053_ (
		.a(new_net_887),
		.b(new_net_446),
		.c(n_1318_)
	);

	or_ii n_2054_ (
		.a(new_net_2377),
		.b(new_net_1106),
		.c(n_1319_)
	);

	or_bb n_2055_ (
		.a(new_net_309),
		.b(new_net_1561),
		.c(n_1320_)
	);

	inv n_2056_ (
		.din(new_net_1580),
		.dout(n_1321_)
	);

	and_bi n_2057_ (
		.a(new_net_564),
		.b(new_net_1296),
		.c(n_1322_)
	);

	and_bi n_2058_ (
		.a(new_net_1240),
		.b(new_net_1417),
		.c(n_1323_)
	);

	and_bb n_2059_ (
		.a(new_net_308),
		.b(new_net_1562),
		.c(n_1324_)
	);

	and_bi n_2060_ (
		.a(new_net_1297),
		.b(new_net_566),
		.c(n_1325_)
	);

	and_ii n_2061_ (
		.a(new_net_1358),
		.b(new_net_1626),
		.c(n_1326_)
	);

	and_bb n_2062_ (
		.a(new_net_1817),
		.b(new_net_1532),
		.c(n_1327_)
	);

	and_bi n_2063_ (
		.a(new_net_1608),
		.b(new_net_1944),
		.c(n_1328_)
	);

	and_bi n_2064_ (
		.a(new_net_1943),
		.b(new_net_1610),
		.c(n_1329_)
	);

	and_ii n_2065_ (
		.a(new_net_317),
		.b(new_net_69),
		.c(n_1330_)
	);

	inv n_2066_ (
		.din(new_net_1896),
		.dout(n_1331_)
	);

	and_bi n_2067_ (
		.a(new_net_882),
		.b(new_net_584),
		.c(n_1332_)
	);

	and_bi n_2068_ (
		.a(new_net_585),
		.b(new_net_883),
		.c(n_1333_)
	);

	and_ii n_2069_ (
		.a(new_net_1542),
		.b(new_net_1518),
		.c(n_1334_)
	);

	or_ii n_2070_ (
		.a(new_net_899),
		.b(new_net_456),
		.c(n_1335_)
	);

	or_bi n_2071_ (
		.a(new_net_1009),
		.b(new_net_1955),
		.c(n_1336_)
	);

	and_ii n_2072_ (
		.a(new_net_39),
		.b(new_net_1660),
		.c(n_1337_)
	);

	and_bb n_2073_ (
		.a(new_net_38),
		.b(new_net_1662),
		.c(n_1338_)
	);

	or_bb n_2074_ (
		.a(new_net_1302),
		.b(new_net_1189),
		.c(n_1339_)
	);

	and_ii n_2075_ (
		.a(new_net_1422),
		.b(new_net_1596),
		.c(n_1340_)
	);

	inv n_2076_ (
		.din(new_net_1480),
		.dout(n_1341_)
	);

	and_bi n_2077_ (
		.a(new_net_1021),
		.b(new_net_1696),
		.c(n_1342_)
	);

	and_bi n_2078_ (
		.a(new_net_1697),
		.b(new_net_1022),
		.c(n_1343_)
	);

	inv n_2079_ (
		.din(new_net_1350),
		.dout(n_1344_)
	);

	and_bi n_2080_ (
		.a(new_net_915),
		.b(new_net_13),
		.c(n_1345_)
	);

	inv n_2081_ (
		.din(new_net_71),
		.dout(n_1346_)
	);

	and_bi n_2082_ (
		.a(new_net_14),
		.b(new_net_914),
		.c(n_1347_)
	);

	and_bb n_2083_ (
		.a(new_net_1504),
		.b(new_net_1227),
		.c(n_1348_)
	);

	or_bb n_2084_ (
		.a(new_net_1505),
		.b(new_net_1228),
		.c(n_1349_)
	);

	inv n_2085_ (
		.din(new_net_1433),
		.dout(n_1350_)
	);

	and_bi n_2086_ (
		.a(new_net_809),
		.b(new_net_466),
		.c(n_1351_)
	);

	and_bi n_2087_ (
		.a(new_net_702),
		.b(new_net_903),
		.c(n_1352_)
	);

	and_ii n_2088_ (
		.a(n_1352_),
		.b(new_net_586),
		.c(n_1353_)
	);

	and_ii n_2089_ (
		.a(new_net_1274),
		.b(new_net_460),
		.c(n_1354_)
	);

	and_bi n_2090_ (
		.a(new_net_2378),
		.b(n_1354_),
		.c(n_1355_)
	);

	and_ii n_2091_ (
		.a(new_net_1509),
		.b(new_net_1830),
		.c(n_1356_)
	);

	or_bb n_2092_ (
		.a(n_1356_),
		.b(new_net_1717),
		.c(n_1357_)
	);

	inv n_2093_ (
		.din(new_net_1802),
		.dout(n_1358_)
	);

	or_bi n_2094_ (
		.a(new_net_361),
		.b(new_net_740),
		.c(n_1359_)
	);

	and_bi n_2095_ (
		.a(new_net_85),
		.b(new_net_1935),
		.c(n_1360_)
	);

	or_bb n_2096_ (
		.a(n_1360_),
		.b(new_net_1875),
		.c(n_1361_)
	);

	and_bi n_2097_ (
		.a(new_net_1678),
		.b(new_net_291),
		.c(n_1362_)
	);

	and_bi n_2098_ (
		.a(new_net_1456),
		.b(new_net_1076),
		.c(n_1363_)
	);

	and_bi n_2099_ (
		.a(new_net_1936),
		.b(new_net_2379),
		.c(n_1364_)
	);

	and_bi n_2100_ (
		.a(new_net_86),
		.b(new_net_679),
		.c(n_1365_)
	);

	or_bb n_2101_ (
		.a(n_1365_),
		.b(new_net_1876),
		.c(n_1366_)
	);

	and_bi n_2102_ (
		.a(new_net_410),
		.b(new_net_420),
		.c(n_1367_)
	);

	and_bi n_2103_ (
		.a(new_net_703),
		.b(new_net_588),
		.c(n_1368_)
	);

	and_bi n_2104_ (
		.a(new_net_467),
		.b(new_net_810),
		.c(n_1369_)
	);

	and_ii n_2105_ (
		.a(new_net_505),
		.b(new_net_904),
		.c(n_1370_)
	);

	or_ii n_2106_ (
		.a(new_net_1277),
		.b(new_net_468),
		.c(n_1371_)
	);

	and_ii n_2107_ (
		.a(new_net_461),
		.b(new_net_72),
		.c(n_0000_)
	);

	and_ii n_2108_ (
		.a(new_net_1831),
		.b(new_net_1718),
		.c(n_0001_)
	);

	or_ii n_2109_ (
		.a(new_net_1811),
		.b(new_net_1753),
		.c(n_0002_)
	);

	or_bb n_2110_ (
		.a(new_net_1951),
		.b(new_net_1398),
		.c(n_0003_)
	);

	and_bi n_2111_ (
		.a(new_net_441),
		.b(new_net_2380),
		.c(n_0004_)
	);

	and_bi n_2112_ (
		.a(new_net_2381),
		.b(n_0004_),
		.c(n_0005_)
	);

	or_bi n_2113_ (
		.a(new_net_426),
		.b(new_net_1534),
		.c(n_0006_)
	);

	and_bi n_2114_ (
		.a(new_net_1243),
		.b(new_net_1359),
		.c(n_0007_)
	);

	or_bb n_2115_ (
		.a(n_0007_),
		.b(new_net_1419),
		.c(n_0008_)
	);

	and_ii n_2116_ (
		.a(new_net_788),
		.b(new_net_1519),
		.c(n_0009_)
	);

	and_ii n_2117_ (
		.a(new_net_20),
		.b(new_net_1543),
		.c(n_0010_)
	);

	and_ii n_2118_ (
		.a(new_net_28),
		.b(new_net_70),
		.c(n_0011_)
	);

	and_ii n_2119_ (
		.a(n_0011_),
		.b(new_net_318),
		.c(n_0012_)
	);

	and_ii n_2120_ (
		.a(new_net_49),
		.b(new_net_1303),
		.c(n_0013_)
	);

	or_bb n_2121_ (
		.a(n_0013_),
		.b(new_net_1190),
		.c(n_0014_)
	);

	or_bi n_2122_ (
		.a(new_net_2382),
		.b(new_net_561),
		.c(n_0015_)
	);

	and_bi n_2123_ (
		.a(new_net_1107),
		.b(new_net_395),
		.c(n_0016_)
	);

	or_bi n_2124_ (
		.a(n_0016_),
		.b(new_net_1217),
		.c(n_0017_)
	);

	and_ii n_2125_ (
		.a(new_net_114),
		.b(new_net_1530),
		.c(n_0018_)
	);

	and_ii n_2126_ (
		.a(n_0018_),
		.b(new_net_1684),
		.c(n_0019_)
	);

	and_bi n_2127_ (
		.a(new_net_1634),
		.b(new_net_329),
		.c(n_0020_)
	);

	or_bi n_2128_ (
		.a(new_net_1636),
		.b(new_net_333),
		.c(n_0021_)
	);

	and_bi n_2129_ (
		.a(new_net_2383),
		.b(new_net_958),
		.c(new_net_2578)
	);

	and_ii n_2130_ (
		.a(new_net_808),
		.b(new_net_392),
		.c(n_0022_)
	);

	and_bi n_2131_ (
		.a(new_net_406),
		.b(new_net_949),
		.c(n_0023_)
	);

	and_bi n_2132_ (
		.a(new_net_948),
		.b(new_net_407),
		.c(n_0024_)
	);

	and_ii n_2133_ (
		.a(new_net_1368),
		.b(new_net_435),
		.c(n_0025_)
	);

	and_bi n_2134_ (
		.a(new_net_1269),
		.b(new_net_18),
		.c(n_0026_)
	);

	and_bi n_2135_ (
		.a(new_net_19),
		.b(new_net_1268),
		.c(n_0027_)
	);

	and_bi n_2136_ (
		.a(new_net_1234),
		.b(new_net_648),
		.c(n_0028_)
	);

	and_bi n_2137_ (
		.a(new_net_649),
		.b(new_net_1236),
		.c(n_0029_)
	);

	and_bi n_2138_ (
		.a(new_net_1880),
		.b(new_net_1838),
		.c(n_0030_)
	);

	and_bi n_2139_ (
		.a(new_net_1837),
		.b(new_net_1879),
		.c(n_0031_)
	);

	and_bi n_2140_ (
		.a(new_net_57),
		.b(new_net_1768),
		.c(n_0032_)
	);

	and_ii n_2141_ (
		.a(new_net_676),
		.b(new_net_655),
		.c(n_0033_)
	);

	and_ii n_2142_ (
		.a(new_net_522),
		.b(new_net_632),
		.c(n_0034_)
	);

	and_ii n_2143_ (
		.a(new_net_712),
		.b(new_net_596),
		.c(n_0035_)
	);

	or_bb n_2144_ (
		.a(new_net_725),
		.b(new_net_1777),
		.c(n_0036_)
	);

	and_bi n_2145_ (
		.a(new_net_1767),
		.b(new_net_58),
		.c(n_0037_)
	);

	and_ii n_2146_ (
		.a(new_net_784),
		.b(new_net_633),
		.c(n_0038_)
	);

	and_bb n_2147_ (
		.a(new_net_523),
		.b(new_net_1093),
		.c(n_0039_)
	);

	and_ii n_2148_ (
		.a(new_net_597),
		.b(new_net_1778),
		.c(n_0040_)
	);

	inv n_2149_ (
		.din(new_net_1248),
		.dout(n_0041_)
	);

	and_bi n_2150_ (
		.a(new_net_813),
		.b(new_net_1373),
		.c(n_0042_)
	);

	and_bi n_2151_ (
		.a(new_net_854),
		.b(new_net_2384),
		.c(n_0043_)
	);

	and_bi n_2152_ (
		.a(new_net_1576),
		.b(new_net_794),
		.c(n_0044_)
	);

	and_bi n_2153_ (
		.a(new_net_796),
		.b(new_net_1578),
		.c(n_0045_)
	);

	and_bi n_2154_ (
		.a(new_net_1459),
		.b(new_net_762),
		.c(n_0046_)
	);

	and_bi n_2155_ (
		.a(new_net_763),
		.b(new_net_1458),
		.c(n_0047_)
	);

	inv n_2156_ (
		.din(new_net_1341),
		.dout(n_0048_)
	);

	and_bi n_2157_ (
		.a(new_net_1000),
		.b(new_net_989),
		.c(n_0049_)
	);

	inv n_2158_ (
		.din(new_net_1030),
		.dout(n_0050_)
	);

	and_bi n_2159_ (
		.a(new_net_991),
		.b(new_net_1001),
		.c(n_0051_)
	);

	and_ii n_2160_ (
		.a(new_net_920),
		.b(new_net_1124),
		.c(n_0052_)
	);

	and_bb n_2161_ (
		.a(new_net_921),
		.b(new_net_1125),
		.c(n_0053_)
	);

	and_bi n_2162_ (
		.a(new_net_1005),
		.b(new_net_1038),
		.c(n_0054_)
	);

	and_ii n_2163_ (
		.a(new_net_1140),
		.b(new_net_932),
		.c(n_0055_)
	);

	and_ii n_2164_ (
		.a(new_net_1220),
		.b(new_net_831),
		.c(n_0056_)
	);

	and_bi n_2165_ (
		.a(new_net_2385),
		.b(n_0056_),
		.c(n_0057_)
	);

	or_bi n_2166_ (
		.a(new_net_984),
		.b(new_net_1449),
		.c(n_0058_)
	);

	and_bi n_2167_ (
		.a(n_0058_),
		.b(new_net_1904),
		.c(n_0059_)
	);

	and_ii n_2168_ (
		.a(new_net_1213),
		.b(new_net_940),
		.c(n_0060_)
	);

	and_ii n_2169_ (
		.a(new_net_1040),
		.b(new_net_933),
		.c(n_0061_)
	);

	and_bb n_2170_ (
		.a(new_net_1857),
		.b(new_net_1637),
		.c(n_0062_)
	);

	and_ii n_2171_ (
		.a(new_net_985),
		.b(new_net_1905),
		.c(n_0063_)
	);

	and_ii n_2172_ (
		.a(new_net_832),
		.b(new_net_1031),
		.c(n_0064_)
	);

	and_bb n_2173_ (
		.a(new_net_1326),
		.b(new_net_91),
		.c(n_0065_)
	);

	and_bb n_2174_ (
		.a(new_net_501),
		.b(new_net_24),
		.c(n_0066_)
	);

	or_bi n_2175_ (
		.a(new_net_620),
		.b(new_net_1756),
		.c(n_0067_)
	);

	and_bi n_2176_ (
		.a(n_0067_),
		.b(new_net_1692),
		.c(n_0068_)
	);

	and_bb n_2177_ (
		.a(new_net_1757),
		.b(new_net_330),
		.c(n_0069_)
	);

	and_bi n_2178_ (
		.a(new_net_2386),
		.b(n_0069_),
		.c(n_0070_)
	);

	and_bi n_2179_ (
		.a(new_net_855),
		.b(new_net_1044),
		.c(n_0071_)
	);

	and_ii n_2180_ (
		.a(n_0071_),
		.b(new_net_873),
		.c(n_0072_)
	);

	and_ii n_2181_ (
		.a(new_net_1222),
		.b(new_net_1688),
		.c(n_0073_)
	);

	or_bb n_2182_ (
		.a(new_net_1336),
		.b(new_net_530),
		.c(n_0074_)
	);

	and_bi n_2183_ (
		.a(new_net_1482),
		.b(new_net_1555),
		.c(n_0075_)
	);

	and_ii n_2184_ (
		.a(new_net_1337),
		.b(new_net_532),
		.c(n_0076_)
	);

	or_bb n_2185_ (
		.a(new_net_1667),
		.b(new_net_1485),
		.c(n_0077_)
	);

	and_bi n_2186_ (
		.a(new_net_2387),
		.b(new_net_1570),
		.c(new_net_2545)
	);

	and_ii n_2187_ (
		.a(new_net_941),
		.b(new_net_1693),
		.c(n_0078_)
	);

	inv n_2188_ (
		.din(new_net_1865),
		.dout(n_0079_)
	);

	inv n_2189_ (
		.din(new_net_92),
		.dout(n_0080_)
	);

	inv n_2190_ (
		.din(new_net_1327),
		.dout(n_0081_)
	);

	and_bi n_2191_ (
		.a(new_net_25),
		.b(new_net_1702),
		.c(n_0082_)
	);

	and_bi n_2192_ (
		.a(new_net_1715),
		.b(new_net_332),
		.c(n_0083_)
	);

	and_bi n_2193_ (
		.a(new_net_635),
		.b(new_net_1681),
		.c(n_0084_)
	);

	and_ii n_2194_ (
		.a(n_0084_),
		.b(new_net_1216),
		.c(n_0085_)
	);

	and_bi n_2195_ (
		.a(new_net_843),
		.b(new_net_1650),
		.c(n_0086_)
	);

	and_bi n_2196_ (
		.a(new_net_1653),
		.b(new_net_844),
		.c(n_0087_)
	);

	or_bb n_2197_ (
		.a(n_0087_),
		.b(n_0086_),
		.c(new_net_2505)
	);

	and_bi n_2198_ (
		.a(new_net_1451),
		.b(new_net_636),
		.c(n_0088_)
	);

	and_bi n_2199_ (
		.a(new_net_1828),
		.b(new_net_1683),
		.c(n_0089_)
	);

	and_bi n_2200_ (
		.a(new_net_1682),
		.b(new_net_1829),
		.c(n_0090_)
	);

	or_bb n_2201_ (
		.a(n_0090_),
		.b(n_0089_),
		.c(new_net_2517)
	);

	and_bi n_2202_ (
		.a(new_net_27),
		.b(new_net_331),
		.c(n_0091_)
	);

	and_bi n_2203_ (
		.a(new_net_1221),
		.b(n_0091_),
		.c(n_0092_)
	);

	and_bi n_2204_ (
		.a(new_net_1704),
		.b(new_net_1939),
		.c(n_0093_)
	);

	and_bi n_2205_ (
		.a(new_net_1940),
		.b(new_net_1703),
		.c(n_0094_)
	);

	or_bb n_2206_ (
		.a(n_0094_),
		.b(n_0093_),
		.c(new_net_2564)
	);

	and_ii n_2207_ (
		.a(new_net_959),
		.b(new_net_1003),
		.c(n_0095_)
	);

	or_ii n_2208_ (
		.a(new_net_75),
		.b(new_net_1858),
		.c(n_0096_)
	);

	or_bb n_2209_ (
		.a(new_net_76),
		.b(new_net_1859),
		.c(n_0097_)
	);

	or_ii n_2210_ (
		.a(n_0097_),
		.b(n_0096_),
		.c(new_net_2495)
	);

	and_bi n_2211_ (
		.a(new_net_1194),
		.b(new_net_1807),
		.c(n_0098_)
	);

	and_bi n_2212_ (
		.a(new_net_1806),
		.b(new_net_1195),
		.c(n_0099_)
	);

	and_bi n_2213_ (
		.a(new_net_1502),
		.b(new_net_1724),
		.c(n_0100_)
	);

	inv n_2214_ (
		.din(new_net_811),
		.dout(n_0101_)
	);

	and_bi n_2215_ (
		.a(new_net_1725),
		.b(new_net_1501),
		.c(n_0102_)
	);

	and_bi n_2216_ (
		.a(new_net_1070),
		.b(new_net_1427),
		.c(n_0103_)
	);

	and_bi n_2217_ (
		.a(new_net_1426),
		.b(new_net_1072),
		.c(n_0104_)
	);

	and_ii n_2218_ (
		.a(new_net_1204),
		.b(new_net_436),
		.c(n_0105_)
	);

	or_bb n_2219_ (
		.a(new_net_1314),
		.b(new_net_323),
		.c(n_0106_)
	);

	and_ii n_2220_ (
		.a(new_net_413),
		.b(new_net_301),
		.c(n_0107_)
	);

	and_bi n_2221_ (
		.a(new_net_2388),
		.b(n_0107_),
		.c(n_0108_)
	);

	and_ii n_2222_ (
		.a(new_net_480),
		.b(new_net_100),
		.c(n_0109_)
	);

	and_ii n_2223_ (
		.a(n_0109_),
		.b(new_net_593),
		.c(n_0110_)
	);

	and_ii n_2224_ (
		.a(new_net_302),
		.b(new_net_812),
		.c(n_0111_)
	);

	and_ii n_2225_ (
		.a(new_net_324),
		.b(new_net_1206),
		.c(n_0112_)
	);

	or_ii n_2226_ (
		.a(new_net_574),
		.b(new_net_1483),
		.c(n_0113_)
	);

	and_bi n_2227_ (
		.a(new_net_542),
		.b(new_net_602),
		.c(n_0114_)
	);

	and_bi n_2228_ (
		.a(new_net_492),
		.b(new_net_1556),
		.c(n_0115_)
	);

	and_ii n_2229_ (
		.a(new_net_101),
		.b(new_net_595),
		.c(n_0116_)
	);

	or_ii n_2230_ (
		.a(new_net_671),
		.b(new_net_661),
		.c(n_0117_)
	);

	or_ii n_2231_ (
		.a(n_0117_),
		.b(new_net_533),
		.c(n_0118_)
	);

	and_bi n_2232_ (
		.a(new_net_1265),
		.b(new_net_1345),
		.c(n_0119_)
	);

	and_bi n_2233_ (
		.a(new_net_1344),
		.b(new_net_1264),
		.c(n_0120_)
	);

	and_ii n_2234_ (
		.a(new_net_758),
		.b(new_net_1034),
		.c(n_0121_)
	);

	and_bi n_2235_ (
		.a(new_net_776),
		.b(new_net_717),
		.c(n_0122_)
	);

	and_bi n_2236_ (
		.a(new_net_718),
		.b(new_net_779),
		.c(n_0123_)
	);

	or_bb n_2237_ (
		.a(n_0123_),
		.b(n_0122_),
		.c(new_net_2556)
	);

	or_bi n_2238_ (
		.a(new_net_662),
		.b(new_net_482),
		.c(n_0124_)
	);

	and_bi n_2239_ (
		.a(new_net_1547),
		.b(new_net_669),
		.c(n_0125_)
	);

	and_bi n_2240_ (
		.a(new_net_672),
		.b(new_net_1548),
		.c(n_0126_)
	);

	or_bb n_2241_ (
		.a(n_0126_),
		.b(n_0125_),
		.c(new_net_2497)
	);

	and_bi n_2242_ (
		.a(new_net_1669),
		.b(new_net_603),
		.c(n_0127_)
	);

	or_bi n_2243_ (
		.a(n_0127_),
		.b(new_net_414),
		.c(n_0128_)
	);

	and_bi n_2244_ (
		.a(new_net_924),
		.b(new_net_545),
		.c(n_0129_)
	);

	and_bi n_2245_ (
		.a(new_net_544),
		.b(new_net_925),
		.c(n_0130_)
	);

	or_bb n_2246_ (
		.a(n_0130_),
		.b(n_0129_),
		.c(new_net_2537)
	);

	and_ii n_2247_ (
		.a(new_net_1571),
		.b(new_net_438),
		.c(n_0131_)
	);

	and_bi n_2248_ (
		.a(new_net_495),
		.b(new_net_576),
		.c(n_0132_)
	);

	and_bi n_2249_ (
		.a(new_net_575),
		.b(new_net_496),
		.c(n_0133_)
	);

	and_ii n_2250_ (
		.a(n_0133_),
		.b(n_0132_),
		.c(new_net_2572)
	);

	or_bb n_2251_ (
		.a(new_net_1687),
		.b(new_net_1391),
		.c(n_0134_)
	);

	or_bb n_2252_ (
		.a(new_net_1934),
		.b(new_net_53),
		.c(n_0135_)
	);

	or_bb n_2253_ (
		.a(n_0135_),
		.b(n_0134_),
		.c(n_0136_)
	);

	or_bb n_2254_ (
		.a(new_net_2389),
		.b(new_net_463),
		.c(n_0137_)
	);

	or_bb n_2255_ (
		.a(new_net_631),
		.b(new_net_724),
		.c(n_0138_)
	);

	or_bb n_2256_ (
		.a(n_0138_),
		.b(n_0137_),
		.c(new_net_2560)
	);

	and_bi n_2257_ (
		.a(new_net_1239),
		.b(new_net_1629),
		.c(n_0139_)
	);

	and_bi n_2258_ (
		.a(new_net_1156),
		.b(new_net_430),
		.c(n_0140_)
	);

	and_bi n_2259_ (
		.a(new_net_427),
		.b(new_net_1157),
		.c(n_0141_)
	);

	and_ii n_2260_ (
		.a(new_net_2390),
		.b(new_net_1621),
		.c(new_net_2525)
	);

	or_bb n_2261_ (
		.a(new_net_428),
		.b(new_net_1598),
		.c(n_0142_)
	);

	and_ii n_2262_ (
		.a(new_net_50),
		.b(new_net_1424),
		.c(n_0143_)
	);

	and_bb n_2263_ (
		.a(new_net_51),
		.b(new_net_1423),
		.c(n_0144_)
	);

	and_ii n_2264_ (
		.a(n_0144_),
		.b(n_0143_),
		.c(n_0145_)
	);

	and_bi n_2265_ (
		.a(n_0142_),
		.b(new_net_303),
		.c(n_0146_)
	);

	and_bi n_2266_ (
		.a(new_net_562),
		.b(n_0146_),
		.c(new_net_2543)
	);

	and_bb n_2267_ (
		.a(new_net_898),
		.b(new_net_1956),
		.c(n_0147_)
	);

	and_bi n_2268_ (
		.a(new_net_580),
		.b(new_net_431),
		.c(n_0148_)
	);

	and_bi n_2269_ (
		.a(new_net_29),
		.b(n_0148_),
		.c(n_0149_)
	);

	or_ii n_2270_ (
		.a(new_net_801),
		.b(new_net_457),
		.c(n_0150_)
	);

	or_bb n_2271_ (
		.a(new_net_802),
		.b(new_net_459),
		.c(n_0151_)
	);

	or_ii n_2272_ (
		.a(n_0151_),
		.b(n_0150_),
		.c(new_net_2511)
	);

	and_ii n_2273_ (
		.a(new_net_1361),
		.b(new_net_1418),
		.c(n_0152_)
	);

	inv n_2274_ (
		.din(new_net_1111),
		.dout(n_0153_)
	);

	and_bi n_2275_ (
		.a(new_net_1623),
		.b(new_net_1184),
		.c(n_0154_)
	);

	or_bi n_2276_ (
		.a(n_0154_),
		.b(new_net_790),
		.c(n_0155_)
	);

	and_bi n_2277_ (
		.a(new_net_1415),
		.b(new_net_896),
		.c(n_0156_)
	);

	and_bi n_2278_ (
		.a(new_net_900),
		.b(new_net_1416),
		.c(n_0157_)
	);

	or_bb n_2279_ (
		.a(n_0157_),
		.b(n_0156_),
		.c(new_net_2523)
	);

	and_bi n_2280_ (
		.a(new_net_1242),
		.b(new_net_1622),
		.c(n_0158_)
	);

	and_bi n_2281_ (
		.a(new_net_1728),
		.b(new_net_1186),
		.c(n_0159_)
	);

	and_bi n_2282_ (
		.a(new_net_1185),
		.b(new_net_1729),
		.c(n_0160_)
	);

	or_bb n_2283_ (
		.a(n_0160_),
		.b(n_0159_),
		.c(new_net_2547)
	);

	and_bb n_2284_ (
		.a(new_net_573),
		.b(new_net_2391),
		.c(new_net_2499)
	);

	inv n_2285_ (
		.din(new_net_1083),
		.dout(n_0161_)
	);

	and_bb n_2286_ (
		.a(new_net_1787),
		.b(new_net_1918),
		.c(n_0162_)
	);

	or_ii n_2287_ (
		.a(new_net_313),
		.b(new_net_1616),
		.c(n_0163_)
	);

	and_bb n_2288_ (
		.a(new_net_314),
		.b(new_net_1467),
		.c(n_0164_)
	);

	and_bi n_2289_ (
		.a(new_net_1086),
		.b(n_0164_),
		.c(n_0165_)
	);

	and_bb n_2290_ (
		.a(new_net_1789),
		.b(new_net_1466),
		.c(n_0166_)
	);

	and_bi n_2291_ (
		.a(new_net_805),
		.b(new_net_1618),
		.c(n_0167_)
	);

	and_bi n_2292_ (
		.a(new_net_1617),
		.b(new_net_806),
		.c(n_0168_)
	);

	and_ii n_2293_ (
		.a(new_net_1006),
		.b(new_net_893),
		.c(n_0169_)
	);

	and_bi n_2294_ (
		.a(new_net_594),
		.b(new_net_759),
		.c(n_0170_)
	);

	and_ii n_2295_ (
		.a(n_0170_),
		.b(new_net_1035),
		.c(n_0171_)
	);

	or_ii n_2296_ (
		.a(new_net_781),
		.b(new_net_673),
		.c(n_0172_)
	);

	and_ii n_2297_ (
		.a(new_net_1420),
		.b(new_net_479),
		.c(n_0173_)
	);

	and_bi n_2298_ (
		.a(new_net_2392),
		.b(n_0173_),
		.c(n_0174_)
	);

	and_bi n_2299_ (
		.a(new_net_663),
		.b(new_net_1421),
		.c(n_0175_)
	);

	and_bi n_2300_ (
		.a(new_net_2393),
		.b(n_0175_),
		.c(n_0176_)
	);

	or_bb n_2301_ (
		.a(new_net_1819),
		.b(new_net_1114),
		.c(n_0177_)
	);

	and_bi n_2302_ (
		.a(new_net_1187),
		.b(new_net_2394),
		.c(n_0178_)
	);

	and_bi n_2303_ (
		.a(new_net_452),
		.b(new_net_1100),
		.c(new_net_2489)
	);

	or_bi n_2304_ (
		.a(new_net_1085),
		.b(new_net_1788),
		.c(n_0179_)
	);

	or_bb n_2305_ (
		.a(new_net_2395),
		.b(new_net_1177),
		.c(n_0180_)
	);

	and_bb n_2306_ (
		.a(new_net_1291),
		.b(new_net_43),
		.c(n_0181_)
	);

	or_bb n_2307_ (
		.a(new_net_927),
		.b(new_net_490),
		.c(n_0182_)
	);

	and_ii n_2308_ (
		.a(new_net_732),
		.b(new_net_423),
		.c(n_0183_)
	);

	or_bb n_2309_ (
		.a(new_net_1430),
		.b(new_net_1258),
		.c(n_0184_)
	);

	and_bi n_2310_ (
		.a(new_net_2396),
		.b(new_net_644),
		.c(n_0185_)
	);

	and_bi n_2311_ (
		.a(new_net_1431),
		.b(new_net_1429),
		.c(n_0186_)
	);

	or_bb n_2312_ (
		.a(n_0186_),
		.b(n_0185_),
		.c(n_0187_)
	);

	or_bb n_2313_ (
		.a(new_net_2397),
		.b(n_0183_),
		.c(n_0188_)
	);

	and_bb n_2314_ (
		.a(new_net_773),
		.b(new_net_1948),
		.c(n_0189_)
	);

	and_bb n_2315_ (
		.a(new_net_730),
		.b(new_net_424),
		.c(n_0190_)
	);

	or_bb n_2316_ (
		.a(n_0190_),
		.b(n_0189_),
		.c(n_0191_)
	);

	and_bi n_2317_ (
		.a(n_0188_),
		.b(n_0191_),
		.c(n_0192_)
	);

	and_ii n_2318_ (
		.a(new_net_772),
		.b(new_net_1949),
		.c(n_0193_)
	);

	and_ii n_2319_ (
		.a(new_net_820),
		.b(new_net_1394),
		.c(n_0194_)
	);

	or_bb n_2320_ (
		.a(n_0194_),
		.b(n_0193_),
		.c(n_0195_)
	);

	or_bb n_2321_ (
		.a(new_net_2398),
		.b(n_0192_),
		.c(n_0196_)
	);

	and_bb n_2322_ (
		.a(new_net_928),
		.b(new_net_489),
		.c(n_0197_)
	);

	and_bb n_2323_ (
		.a(new_net_821),
		.b(new_net_1393),
		.c(n_0198_)
	);

	or_bb n_2324_ (
		.a(n_0198_),
		.b(n_0197_),
		.c(n_0199_)
	);

	and_bi n_2325_ (
		.a(n_0196_),
		.b(new_net_2399),
		.c(n_0200_)
	);

	and_bi n_2326_ (
		.a(new_net_2400),
		.b(n_0200_),
		.c(n_0201_)
	);

	and_ii n_2327_ (
		.a(n_0201_),
		.b(new_net_2401),
		.c(n_0202_)
	);

	and_ii n_2328_ (
		.a(new_net_1528),
		.b(new_net_767),
		.c(n_0203_)
	);

	and_ii n_2329_ (
		.a(new_net_1293),
		.b(new_net_42),
		.c(n_0204_)
	);

	or_bb n_2330_ (
		.a(n_0204_),
		.b(n_0203_),
		.c(n_0205_)
	);

	and_ii n_2331_ (
		.a(new_net_2402),
		.b(n_0202_),
		.c(n_0206_)
	);

	and_bb n_2332_ (
		.a(new_net_1181),
		.b(new_net_1927),
		.c(n_0207_)
	);

	and_ii n_2333_ (
		.a(new_net_559),
		.b(new_net_1888),
		.c(n_0208_)
	);

	or_bb n_2334_ (
		.a(new_net_908),
		.b(new_net_1698),
		.c(n_0209_)
	);

	and_bb n_2335_ (
		.a(new_net_1529),
		.b(new_net_765),
		.c(n_0210_)
	);

	and_bb n_2336_ (
		.a(new_net_558),
		.b(new_net_1887),
		.c(n_0211_)
	);

	or_bb n_2337_ (
		.a(n_0211_),
		.b(n_0210_),
		.c(n_0212_)
	);

	or_bb n_2338_ (
		.a(new_net_2403),
		.b(n_0209_),
		.c(n_0213_)
	);

	and_ii n_2339_ (
		.a(new_net_2404),
		.b(n_0206_),
		.c(n_0214_)
	);

	and_bi n_2340_ (
		.a(new_net_909),
		.b(new_net_1699),
		.c(n_0215_)
	);

	and_ii n_2341_ (
		.a(new_net_1180),
		.b(new_net_1926),
		.c(n_0216_)
	);

	and_ii n_2342_ (
		.a(new_net_1848),
		.b(new_net_1489),
		.c(n_0217_)
	);

	or_bb n_2343_ (
		.a(n_0217_),
		.b(n_0216_),
		.c(n_0218_)
	);

	or_bb n_2344_ (
		.a(new_net_2405),
		.b(n_0215_),
		.c(n_0219_)
	);

	and_ii n_2345_ (
		.a(new_net_2406),
		.b(n_0214_),
		.c(n_0220_)
	);

	and_ii n_2346_ (
		.a(new_net_1664),
		.b(new_net_1932),
		.c(n_0221_)
	);

	and_ii n_2347_ (
		.a(new_net_1854),
		.b(new_net_975),
		.c(n_0222_)
	);

	or_bb n_2348_ (
		.a(n_0222_),
		.b(n_0221_),
		.c(n_0223_)
	);

	and_bb n_2349_ (
		.a(new_net_824),
		.b(new_net_1092),
		.c(n_0224_)
	);

	and_bb n_2350_ (
		.a(new_net_1666),
		.b(new_net_1930),
		.c(n_0225_)
	);

	and_bb n_2351_ (
		.a(new_net_1852),
		.b(new_net_976),
		.c(n_0226_)
	);

	or_bb n_2352_ (
		.a(new_net_108),
		.b(new_net_2407),
		.c(n_0227_)
	);

	or_bb n_2353_ (
		.a(n_0227_),
		.b(new_net_2408),
		.c(n_0228_)
	);

	and_ii n_2354_ (
		.a(n_0228_),
		.b(new_net_61),
		.c(n_0229_)
	);

	and_ii n_2355_ (
		.a(new_net_612),
		.b(new_net_751),
		.c(n_0230_)
	);

	and_ii n_2356_ (
		.a(new_net_825),
		.b(new_net_1090),
		.c(n_0231_)
	);

	and_ii n_2357_ (
		.a(n_0231_),
		.b(n_0230_),
		.c(n_0232_)
	);

	and_bb n_2358_ (
		.a(new_net_1846),
		.b(new_net_1490),
		.c(n_0233_)
	);

	and_bb n_2359_ (
		.a(new_net_614),
		.b(new_net_750),
		.c(n_0234_)
	);

	and_ii n_2360_ (
		.a(n_0234_),
		.b(n_0233_),
		.c(n_0235_)
	);

	and_bb n_2361_ (
		.a(new_net_2409),
		.b(new_net_1809),
		.c(n_0236_)
	);

	or_ii n_2362_ (
		.a(new_net_2410),
		.b(new_net_1524),
		.c(n_0237_)
	);

	and_ii n_2363_ (
		.a(new_net_2411),
		.b(n_0220_),
		.c(n_0238_)
	);

	and_bi n_2364_ (
		.a(new_net_1525),
		.b(new_net_1810),
		.c(n_0239_)
	);

	and_bi n_2365_ (
		.a(new_net_62),
		.b(new_net_109),
		.c(n_0240_)
	);

	or_bb n_2366_ (
		.a(new_net_2412),
		.b(n_0239_),
		.c(n_0241_)
	);

	and_ii n_2367_ (
		.a(new_net_2413),
		.b(n_0238_),
		.c(n_0242_)
	);

	and_bb n_2368_ (
		.a(new_net_1554),
		.b(new_net_1149),
		.c(n_0243_)
	);

	and_ii n_2369_ (
		.a(new_net_1322),
		.b(new_net_1247),
		.c(n_0244_)
	);

	and_ii n_2370_ (
		.a(new_net_719),
		.b(new_net_692),
		.c(n_0245_)
	);

	and_ii n_2371_ (
		.a(new_net_1552),
		.b(new_net_1148),
		.c(n_0246_)
	);

	and_bb n_2372_ (
		.a(new_net_1321),
		.b(new_net_1246),
		.c(n_0247_)
	);

	or_bb n_2373_ (
		.a(new_net_2414),
		.b(new_net_752),
		.c(n_0248_)
	);

	and_bi n_2374_ (
		.a(n_0245_),
		.b(n_0248_),
		.c(n_0249_)
	);

	and_ii n_2375_ (
		.a(new_net_498),
		.b(new_net_526),
		.c(n_0250_)
	);

	and_ii n_2376_ (
		.a(new_net_89),
		.b(new_net_1604),
		.c(n_0251_)
	);

	and_ii n_2377_ (
		.a(n_0251_),
		.b(n_0250_),
		.c(n_0252_)
	);

	and_bb n_2378_ (
		.a(new_net_500),
		.b(new_net_525),
		.c(n_0253_)
	);

	and_bb n_2379_ (
		.a(new_net_90),
		.b(new_net_1603),
		.c(n_0254_)
	);

	and_ii n_2380_ (
		.a(new_net_2415),
		.b(new_net_879),
		.c(n_0255_)
	);

	and_bb n_2381_ (
		.a(n_0255_),
		.b(new_net_866),
		.c(n_0256_)
	);

	or_ii n_2382_ (
		.a(new_net_2416),
		.b(new_net_816),
		.c(n_0257_)
	);

	and_ii n_2383_ (
		.a(new_net_2417),
		.b(n_0242_),
		.c(n_0258_)
	);

	or_bb n_2384_ (
		.a(new_net_880),
		.b(new_net_867),
		.c(n_0259_)
	);

	and_bi n_2385_ (
		.a(new_net_817),
		.b(new_net_2418),
		.c(n_0260_)
	);

	and_bi n_2386_ (
		.a(new_net_720),
		.b(new_net_693),
		.c(n_0261_)
	);

	or_bb n_2387_ (
		.a(n_0261_),
		.b(new_net_753),
		.c(n_0262_)
	);

	or_bb n_2388_ (
		.a(new_net_2419),
		.b(n_0260_),
		.c(n_0263_)
	);

	and_ii n_2389_ (
		.a(new_net_2420),
		.b(n_0258_),
		.c(n_0264_)
	);

	and_bi n_2390_ (
		.a(new_net_1016),
		.b(new_net_540),
		.c(n_0265_)
	);

	and_ii n_2391_ (
		.a(new_net_623),
		.b(new_net_1198),
		.c(n_0266_)
	);

	or_bb n_2392_ (
		.a(n_0266_),
		.b(new_net_2421),
		.c(n_0267_)
	);

	and_bi n_2393_ (
		.a(new_net_539),
		.b(new_net_1015),
		.c(n_0268_)
	);

	and_bb n_2394_ (
		.a(new_net_624),
		.b(new_net_1199),
		.c(n_0269_)
	);

	or_bb n_2395_ (
		.a(n_0269_),
		.b(new_net_1200),
		.c(n_0270_)
	);

	and_ii n_2396_ (
		.a(new_net_2422),
		.b(new_net_112),
		.c(n_0271_)
	);

	and_ii n_2397_ (
		.a(new_net_1743),
		.b(new_net_1826),
		.c(n_0272_)
	);

	and_ii n_2398_ (
		.a(new_net_95),
		.b(new_net_321),
		.c(n_0273_)
	);

	and_ii n_2399_ (
		.a(n_0273_),
		.b(n_0272_),
		.c(n_0274_)
	);

	and_bb n_2400_ (
		.a(new_net_1744),
		.b(new_net_1827),
		.c(n_0275_)
	);

	and_bb n_2401_ (
		.a(new_net_96),
		.b(new_net_320),
		.c(n_0276_)
	);

	and_ii n_2402_ (
		.a(new_net_2423),
		.b(new_net_1366),
		.c(n_0277_)
	);

	or_ii n_2403_ (
		.a(n_0277_),
		.b(new_net_1324),
		.c(n_0278_)
	);

	and_bi n_2404_ (
		.a(new_net_768),
		.b(new_net_2424),
		.c(n_0279_)
	);

	and_ii n_2405_ (
		.a(new_net_1403),
		.b(new_net_982),
		.c(n_0280_)
	);

	and_bb n_2406_ (
		.a(new_net_1404),
		.b(new_net_981),
		.c(n_0281_)
	);

	and_ii n_2407_ (
		.a(new_net_2425),
		.b(new_net_1705),
		.c(n_0282_)
	);

	or_ii n_2408_ (
		.a(new_net_2426),
		.b(new_net_1435),
		.c(n_0283_)
	);

	or_bb n_2409_ (
		.a(new_net_2427),
		.b(new_net_1793),
		.c(n_0284_)
	);

	and_bb n_2410_ (
		.a(new_net_1706),
		.b(new_net_1436),
		.c(n_0285_)
	);

	or_bb n_2411_ (
		.a(new_net_1367),
		.b(new_net_1325),
		.c(n_0286_)
	);

	and_bi n_2412_ (
		.a(new_net_769),
		.b(new_net_2428),
		.c(n_0287_)
	);

	and_bi n_2413_ (
		.a(new_net_113),
		.b(new_net_1201),
		.c(n_0288_)
	);

	or_bb n_2414_ (
		.a(new_net_2429),
		.b(n_0287_),
		.c(n_0289_)
	);

	or_bb n_2415_ (
		.a(new_net_2430),
		.b(n_0285_),
		.c(n_0290_)
	);

	and_bi n_2416_ (
		.a(n_0284_),
		.b(new_net_2431),
		.c(n_0291_)
	);

	and_bi n_2417_ (
		.a(new_net_1516),
		.b(new_net_1412),
		.c(n_0292_)
	);

	and_bi n_2418_ (
		.a(new_net_619),
		.b(new_net_1493),
		.c(n_0293_)
	);

	or_bb n_2419_ (
		.a(n_0293_),
		.b(n_0292_),
		.c(n_0294_)
	);

	and_bi n_2420_ (
		.a(new_net_1411),
		.b(new_net_1517),
		.c(n_0295_)
	);

	and_bi n_2421_ (
		.a(new_net_1494),
		.b(new_net_618),
		.c(n_0296_)
	);

	and_ii n_2422_ (
		.a(new_net_1605),
		.b(new_net_2432),
		.c(n_0297_)
	);

	and_bi n_2423_ (
		.a(n_0297_),
		.b(new_net_1396),
		.c(n_0298_)
	);

	and_bi n_2424_ (
		.a(new_net_1334),
		.b(new_net_66),
		.c(n_0299_)
	);

	and_bi n_2425_ (
		.a(new_net_1043),
		.b(new_net_639),
		.c(n_0300_)
	);

	and_ii n_2426_ (
		.a(n_0300_),
		.b(n_0299_),
		.c(n_0301_)
	);

	and_bi n_2427_ (
		.a(new_net_64),
		.b(new_net_1335),
		.c(n_0302_)
	);

	and_bi n_2428_ (
		.a(new_net_640),
		.b(new_net_1042),
		.c(n_0303_)
	);

	and_ii n_2429_ (
		.a(new_net_2433),
		.b(new_net_404),
		.c(n_0304_)
	);

	and_bb n_2430_ (
		.a(n_0304_),
		.b(new_net_1923),
		.c(n_0305_)
	);

	or_ii n_2431_ (
		.a(new_net_2434),
		.b(new_net_1795),
		.c(n_0306_)
	);

	or_bb n_2432_ (
		.a(new_net_2435),
		.b(n_0291_),
		.c(n_0307_)
	);

	or_bb n_2433_ (
		.a(new_net_405),
		.b(new_net_1924),
		.c(n_0308_)
	);

	and_bi n_2434_ (
		.a(new_net_1796),
		.b(new_net_2436),
		.c(n_0309_)
	);

	and_bi n_2435_ (
		.a(new_net_1397),
		.b(new_net_1606),
		.c(n_0310_)
	);

	or_bb n_2436_ (
		.a(new_net_2437),
		.b(n_0309_),
		.c(n_0311_)
	);

	and_bi n_2437_ (
		.a(n_0307_),
		.b(new_net_2438),
		.c(n_0312_)
	);

	and_bi n_2438_ (
		.a(new_net_1882),
		.b(new_net_743),
		.c(n_0313_)
	);

	and_bb n_2439_ (
		.a(new_net_1463),
		.b(new_net_1800),
		.c(n_0314_)
	);

	and_ii n_2440_ (
		.a(new_net_1462),
		.b(new_net_1798),
		.c(n_0315_)
	);

	or_bb n_2441_ (
		.a(new_net_1306),
		.b(new_net_986),
		.c(n_0316_)
	);

	and_bi n_2442_ (
		.a(new_net_668),
		.b(new_net_1583),
		.c(n_0317_)
	);

	and_bi n_2443_ (
		.a(new_net_1585),
		.b(new_net_667),
		.c(n_0318_)
	);

	or_bb n_2444_ (
		.a(new_net_2439),
		.b(new_net_1362),
		.c(n_0319_)
	);

	or_bb n_2445_ (
		.a(n_0319_),
		.b(n_0316_),
		.c(n_0320_)
	);

	and_ii n_2446_ (
		.a(n_0320_),
		.b(new_net_2440),
		.c(n_0321_)
	);

	and_ii n_2447_ (
		.a(new_net_1440),
		.b(new_net_382),
		.c(n_0322_)
	);

	and_bi n_2448_ (
		.a(new_net_367),
		.b(new_net_999),
		.c(n_0323_)
	);

	or_bb n_2449_ (
		.a(n_0323_),
		.b(new_net_2441),
		.c(n_0324_)
	);

	and_bb n_2450_ (
		.a(new_net_1441),
		.b(new_net_373),
		.c(n_0325_)
	);

	and_bi n_2451_ (
		.a(new_net_742),
		.b(new_net_1884),
		.c(n_0326_)
	);

	and_bi n_2452_ (
		.a(new_net_997),
		.b(new_net_366),
		.c(n_0327_)
	);

	or_bb n_2453_ (
		.a(new_net_1586),
		.b(new_net_415),
		.c(n_0328_)
	);

	or_bb n_2454_ (
		.a(n_0328_),
		.b(new_net_2442),
		.c(n_0329_)
	);

	and_ii n_2455_ (
		.a(n_0329_),
		.b(new_net_1520),
		.c(n_0330_)
	);

	or_ii n_2456_ (
		.a(new_net_2443),
		.b(new_net_1707),
		.c(n_0331_)
	);

	or_bb n_2457_ (
		.a(new_net_2444),
		.b(n_0312_),
		.c(n_0332_)
	);

	or_bi n_2458_ (
		.a(new_net_1587),
		.b(new_net_1521),
		.c(n_0333_)
	);

	and_bi n_2459_ (
		.a(n_0333_),
		.b(new_net_416),
		.c(n_0334_)
	);

	and_bi n_2460_ (
		.a(new_net_1708),
		.b(new_net_2445),
		.c(n_0335_)
	);

	and_bi n_2461_ (
		.a(new_net_1790),
		.b(new_net_1170),
		.c(n_0336_)
	);

	and_bi n_2462_ (
		.a(new_net_1084),
		.b(n_0336_),
		.c(n_0337_)
	);

	or_bb n_2463_ (
		.a(new_net_1363),
		.b(new_net_1307),
		.c(n_0338_)
	);

	and_bi n_2464_ (
		.a(n_0338_),
		.b(new_net_987),
		.c(n_0339_)
	);

	or_bb n_2465_ (
		.a(n_0339_),
		.b(new_net_2446),
		.c(n_0340_)
	);

	or_bb n_2466_ (
		.a(new_net_2447),
		.b(n_0335_),
		.c(n_0341_)
	);

	and_bi n_2467_ (
		.a(n_0332_),
		.b(new_net_2448),
		.c(n_0342_)
	);

	and_bi n_2468_ (
		.a(new_net_1134),
		.b(new_net_293),
		.c(new_net_7)
	);

	inv n_2469_ (
		.din(new_net_1755),
		.dout(n_0343_)
	);

	or_bb n_2470_ (
		.a(new_net_417),
		.b(new_net_1400),
		.c(n_0344_)
	);

	or_bi n_2471_ (
		.a(new_net_555),
		.b(new_net_444),
		.c(n_0345_)
	);

	and_bi n_2472_ (
		.a(n_0345_),
		.b(new_net_1511),
		.c(n_0346_)
	);

	or_ii n_2473_ (
		.a(new_net_31),
		.b(new_net_1814),
		.c(n_0347_)
	);

	or_bb n_2474_ (
		.a(new_net_32),
		.b(new_net_1812),
		.c(n_0348_)
	);

	or_ii n_2475_ (
		.a(n_0348_),
		.b(n_0347_),
		.c(new_net_2501)
	);

	and_bi n_2476_ (
		.a(new_net_442),
		.b(new_net_506),
		.c(n_0349_)
	);

	or_ii n_2477_ (
		.a(new_net_59),
		.b(new_net_469),
		.c(n_0350_)
	);

	and_bi n_2478_ (
		.a(n_0350_),
		.b(new_net_1276),
		.c(n_0351_)
	);

	and_bi n_2479_ (
		.a(new_net_102),
		.b(new_net_419),
		.c(n_0352_)
	);

	and_bi n_2480_ (
		.a(new_net_418),
		.b(new_net_103),
		.c(n_0353_)
	);

	or_bb n_2481_ (
		.a(n_0353_),
		.b(n_0352_),
		.c(new_net_2515)
	);

	inv n_2482_ (
		.din(new_net_470),
		.dout(n_0354_)
	);

	and_ii n_2483_ (
		.a(new_net_60),
		.b(new_net_907),
		.c(n_0355_)
	);

	and_bi n_2484_ (
		.a(new_net_336),
		.b(new_net_1782),
		.c(n_0356_)
	);

	and_bi n_2485_ (
		.a(new_net_1783),
		.b(new_net_337),
		.c(n_0357_)
	);

	or_bb n_2486_ (
		.a(n_0357_),
		.b(n_0356_),
		.c(new_net_2535)
	);

	and_bi n_2487_ (
		.a(new_net_445),
		.b(new_net_1278),
		.c(n_0358_)
	);

	and_bi n_2488_ (
		.a(new_net_1279),
		.b(new_net_443),
		.c(n_0359_)
	);

	or_bb n_2489_ (
		.a(n_0359_),
		.b(n_0358_),
		.c(new_net_2493)
	);

	inv n_2490_ (
		.din(new_net_1794),
		.dout(new_net_2570)
	);

	and_ii n_2491_ (
		.a(new_net_1689),
		.b(new_net_531),
		.c(n_0360_)
	);

	and_bi n_2492_ (
		.a(new_net_1223),
		.b(new_net_472),
		.c(n_0361_)
	);

	and_bi n_2493_ (
		.a(new_net_475),
		.b(new_net_1224),
		.c(n_0362_)
	);

	or_bb n_2494_ (
		.a(n_0362_),
		.b(n_0361_),
		.c(new_net_2491)
	);

	and_bb n_2495_ (
		.a(new_net_1047),
		.b(new_net_814),
		.c(n_0363_)
	);

	and_ii n_2496_ (
		.a(n_0363_),
		.b(new_net_714),
		.c(n_0364_)
	);

	and_bi n_2497_ (
		.a(new_net_567),
		.b(new_net_1374),
		.c(n_0365_)
	);

	and_bi n_2498_ (
		.a(new_net_1375),
		.b(new_net_568),
		.c(n_0366_)
	);

	or_bb n_2499_ (
		.a(n_0366_),
		.b(n_0365_),
		.c(new_net_2521)
	);

	and_ii n_2500_ (
		.a(new_net_658),
		.b(new_net_634),
		.c(n_0367_)
	);

	and_bi n_2501_ (
		.a(new_net_1048),
		.b(new_net_786),
		.c(n_0368_)
	);

	or_bb n_2502_ (
		.a(n_0368_),
		.b(new_net_677),
		.c(n_0369_)
	);

	or_ii n_2503_ (
		.a(new_net_690),
		.b(new_net_1378),
		.c(n_0370_)
	);

	and_ii n_2504_ (
		.a(new_net_691),
		.b(new_net_1380),
		.c(n_0371_)
	);

	and_bi n_2505_ (
		.a(n_0370_),
		.b(n_0371_),
		.c(new_net_2566)
	);

	and_ii n_2506_ (
		.a(new_net_678),
		.b(new_net_783),
		.c(n_0372_)
	);

	or_ii n_2507_ (
		.a(new_net_1049),
		.b(new_net_1906),
		.c(n_0373_)
	);

	and_ii n_2508_ (
		.a(new_net_1045),
		.b(new_net_1908),
		.c(n_0374_)
	);

	and_bi n_2509_ (
		.a(n_0373_),
		.b(n_0374_),
		.c(new_net_2549)
	);

	or_ii n_2510_ (
		.a(new_net_1820),
		.b(new_net_895),
		.c(n_0375_)
	);

	and_bi n_2511_ (
		.a(new_net_1007),
		.b(new_net_1822),
		.c(n_0376_)
	);

	and_bi n_2512_ (
		.a(n_0375_),
		.b(n_0376_),
		.c(n_0377_)
	);

	or_ii n_2513_ (
		.a(new_net_664),
		.b(new_net_316),
		.c(n_0378_)
	);

	inv n_2514_ (
		.din(new_net_315),
		.dout(n_0379_)
	);

	and_bi n_2515_ (
		.a(new_net_876),
		.b(new_net_665),
		.c(n_0380_)
	);

	and_bi n_2516_ (
		.a(n_0378_),
		.b(n_0380_),
		.c(new_net_8)
	);

	and_bb n_2517_ (
		.a(new_net_1823),
		.b(new_net_1115),
		.c(n_0381_)
	);

	and_bi n_2518_ (
		.a(new_net_1188),
		.b(new_net_2449),
		.c(new_net_9)
	);

	and_ii n_2519_ (
		.a(new_net_1685),
		.b(new_net_1531),
		.c(n_0382_)
	);

	or_bi n_2520_ (
		.a(new_net_966),
		.b(new_net_115),
		.c(n_0383_)
	);

	and_bi n_2521_ (
		.a(new_net_970),
		.b(new_net_116),
		.c(n_0384_)
	);

	and_bi n_2522_ (
		.a(n_0383_),
		.b(n_0384_),
		.c(new_net_2509)
	);

	and_ii n_2523_ (
		.a(new_net_1734),
		.b(new_net_1816),
		.c(n_0385_)
	);

	and_bb n_2524_ (
		.a(new_net_397),
		.b(new_net_888),
		.c(n_0386_)
	);

	and_ii n_2525_ (
		.a(n_0386_),
		.b(new_net_890),
		.c(n_0387_)
	);

	or_ii n_2526_ (
		.a(new_net_1870),
		.b(new_net_1496),
		.c(n_0388_)
	);

	or_bb n_2527_ (
		.a(new_net_1871),
		.b(new_net_1499),
		.c(n_0389_)
	);

	or_ii n_2528_ (
		.a(n_0389_),
		.b(n_0388_),
		.c(new_net_2503)
	);

	inv n_2529_ (
		.din(new_net_1137),
		.dout(n_0390_)
	);

	and_ii n_2530_ (
		.a(new_net_396),
		.b(new_net_700),
		.c(n_0391_)
	);

	or_bb n_2531_ (
		.a(n_0391_),
		.b(new_net_1155),
		.c(n_0392_)
	);

	or_ii n_2532_ (
		.a(new_net_645),
		.b(new_net_355),
		.c(n_0393_)
	);

	and_bi n_2533_ (
		.a(new_net_1139),
		.b(new_net_646),
		.c(n_0394_)
	);

	and_bi n_2534_ (
		.a(n_0393_),
		.b(n_0394_),
		.c(new_net_2574)
	);

	or_bi n_2535_ (
		.a(new_net_1168),
		.b(new_net_400),
		.c(n_0395_)
	);

	and_bi n_2536_ (
		.a(new_net_1167),
		.b(new_net_398),
		.c(n_0396_)
	);

	and_bi n_2537_ (
		.a(n_0395_),
		.b(n_0396_),
		.c(new_net_2576)
	);

	and_ii n_2538_ (
		.a(new_net_1860),
		.b(new_net_1635),
		.c(n_0397_)
	);

	or_bb n_2539_ (
		.a(new_net_2450),
		.b(new_net_26),
		.c(n_0398_)
	);

	and_bi n_2540_ (
		.a(new_net_1215),
		.b(new_net_1286),
		.c(n_0399_)
	);

	and_bi n_2541_ (
		.a(new_net_1287),
		.b(new_net_1214),
		.c(n_0400_)
	);

	and_ii n_2542_ (
		.a(n_0400_),
		.b(n_0399_),
		.c(n_0401_)
	);

	and_ii n_2543_ (
		.a(new_net_1572),
		.b(new_net_621),
		.c(n_0402_)
	);

	and_bi n_2544_ (
		.a(new_net_1447),
		.b(new_net_1716),
		.c(n_0403_)
	);

	and_bi n_2545_ (
		.a(new_net_1110),
		.b(new_net_935),
		.c(n_0404_)
	);

	and_ii n_2546_ (
		.a(new_net_1039),
		.b(new_net_1109),
		.c(n_0405_)
	);

	and_ii n_2547_ (
		.a(n_0405_),
		.b(n_0404_),
		.c(n_0406_)
	);

	and_bi n_2548_ (
		.a(new_net_1866),
		.b(new_net_1473),
		.c(n_0407_)
	);

	and_bi n_2549_ (
		.a(new_net_1474),
		.b(new_net_1867),
		.c(n_0408_)
	);

	and_ii n_2550_ (
		.a(n_0408_),
		.b(n_0407_),
		.c(n_0409_)
	);

	and_bb n_2551_ (
		.a(new_net_1538),
		.b(new_net_1760),
		.c(n_0410_)
	);

	and_ii n_2552_ (
		.a(new_net_1539),
		.b(new_net_1761),
		.c(n_0411_)
	);

	or_bb n_2553_ (
		.a(n_0411_),
		.b(n_0410_),
		.c(n_0412_)
	);

	or_bb n_2554_ (
		.a(new_net_950),
		.b(new_net_1384),
		.c(n_0413_)
	);

	and_bb n_2555_ (
		.a(new_net_951),
		.b(new_net_1385),
		.c(n_0414_)
	);

	and_bi n_2556_ (
		.a(n_0413_),
		.b(n_0414_),
		.c(n_0415_)
	);

	or_bb n_2557_ (
		.a(new_net_2451),
		.b(new_net_334),
		.c(n_0416_)
	);

	and_ii n_2558_ (
		.a(new_net_934),
		.b(new_net_1004),
		.c(n_0417_)
	);

	and_ii n_2559_ (
		.a(new_net_2452),
		.b(new_net_1141),
		.c(n_0418_)
	);

	and_bi n_2560_ (
		.a(new_net_1711),
		.b(new_net_1651),
		.c(n_0419_)
	);

	and_bi n_2561_ (
		.a(new_net_1652),
		.b(new_net_1712),
		.c(n_0420_)
	);

	and_ii n_2562_ (
		.a(n_0420_),
		.b(n_0419_),
		.c(n_0421_)
	);

	and_bi n_2563_ (
		.a(new_net_1450),
		.b(new_net_1893),
		.c(n_0422_)
	);

	and_bi n_2564_ (
		.a(new_net_1894),
		.b(new_net_1448),
		.c(n_0423_)
	);

	and_ii n_2565_ (
		.a(n_0423_),
		.b(n_0422_),
		.c(n_0424_)
	);

	and_bb n_2566_ (
		.a(new_net_393),
		.b(new_net_1573),
		.c(n_0425_)
	);

	and_ii n_2567_ (
		.a(new_net_394),
		.b(new_net_1574),
		.c(n_0426_)
	);

	or_bb n_2568_ (
		.a(n_0426_),
		.b(n_0425_),
		.c(n_0427_)
	);

	and_bi n_2569_ (
		.a(new_net_335),
		.b(new_net_2453),
		.c(n_0428_)
	);

	and_bi n_2570_ (
		.a(n_0416_),
		.b(n_0428_),
		.c(n_0429_)
	);

	and_ii n_2571_ (
		.a(new_net_1328),
		.b(new_net_93),
		.c(n_0430_)
	);

	or_bb n_2572_ (
		.a(new_net_2454),
		.b(new_net_502),
		.c(n_0431_)
	);

	or_bi n_2573_ (
		.a(new_net_33),
		.b(new_net_368),
		.c(n_0432_)
	);

	and_bi n_2574_ (
		.a(new_net_34),
		.b(new_net_369),
		.c(n_0433_)
	);

	and_bi n_2575_ (
		.a(n_0432_),
		.b(n_0433_),
		.c(n_0434_)
	);

	and_bi n_2576_ (
		.a(new_net_713),
		.b(new_net_1779),
		.c(n_0435_)
	);

	and_ii n_2577_ (
		.a(new_net_2455),
		.b(new_net_726),
		.c(n_0436_)
	);

	and_bi n_2578_ (
		.a(new_net_1094),
		.b(new_net_656),
		.c(n_0437_)
	);

	and_bi n_2579_ (
		.a(new_net_785),
		.b(new_net_1381),
		.c(n_0438_)
	);

	or_bb n_2580_ (
		.a(n_0438_),
		.b(n_0437_),
		.c(n_0439_)
	);

	and_bi n_2581_ (
		.a(new_net_476),
		.b(new_net_1251),
		.c(n_0440_)
	);

	and_bi n_2582_ (
		.a(new_net_1250),
		.b(new_net_474),
		.c(n_0441_)
	);

	or_bb n_2583_ (
		.a(n_0441_),
		.b(n_0440_),
		.c(n_0442_)
	);

	and_ii n_2584_ (
		.a(new_net_1592),
		.b(new_net_1270),
		.c(n_0443_)
	);

	and_bb n_2585_ (
		.a(new_net_1593),
		.b(new_net_1271),
		.c(n_0444_)
	);

	and_ii n_2586_ (
		.a(n_0444_),
		.b(n_0443_),
		.c(n_0445_)
	);

	and_bi n_2587_ (
		.a(new_net_1898),
		.b(new_net_956),
		.c(n_0446_)
	);

	and_bi n_2588_ (
		.a(new_net_957),
		.b(new_net_1899),
		.c(n_0447_)
	);

	or_bb n_2589_ (
		.a(n_0447_),
		.b(n_0446_),
		.c(n_0448_)
	);

	and_ii n_2590_ (
		.a(new_net_2456),
		.b(new_net_1046),
		.c(n_0449_)
	);

	and_bi n_2591_ (
		.a(new_net_787),
		.b(new_net_657),
		.c(n_0450_)
	);

	and_ii n_2592_ (
		.a(new_net_2457),
		.b(new_net_1095),
		.c(n_0451_)
	);

	and_bi n_2593_ (
		.a(new_net_746),
		.b(new_net_1252),
		.c(n_0452_)
	);

	and_bi n_2594_ (
		.a(new_net_1249),
		.b(new_net_747),
		.c(n_0453_)
	);

	and_ii n_2595_ (
		.a(n_0453_),
		.b(n_0452_),
		.c(n_0454_)
	);

	and_ii n_2596_ (
		.a(new_net_1907),
		.b(new_net_1379),
		.c(n_0455_)
	);

	and_ii n_2597_ (
		.a(new_net_2458),
		.b(new_net_815),
		.c(n_0456_)
	);

	or_ii n_2598_ (
		.a(new_net_1630),
		.b(new_net_473),
		.c(n_0457_)
	);

	and_ii n_2599_ (
		.a(new_net_1631),
		.b(new_net_477),
		.c(n_0458_)
	);

	and_bi n_2600_ (
		.a(n_0457_),
		.b(n_0458_),
		.c(n_0459_)
	);

	and_ii n_2601_ (
		.a(new_net_1594),
		.b(new_net_874),
		.c(n_0460_)
	);

	and_bb n_2602_ (
		.a(new_net_1595),
		.b(new_net_875),
		.c(n_0461_)
	);

	and_ii n_2603_ (
		.a(n_0461_),
		.b(n_0460_),
		.c(n_0462_)
	);

	and_bi n_2604_ (
		.a(new_net_1902),
		.b(new_net_1087),
		.c(n_0463_)
	);

	and_bi n_2605_ (
		.a(new_net_1088),
		.b(new_net_1903),
		.c(n_0464_)
	);

	or_bb n_2606_ (
		.a(n_0464_),
		.b(n_0463_),
		.c(n_0465_)
	);

	and_bi n_2607_ (
		.a(new_net_1050),
		.b(new_net_2459),
		.c(n_0466_)
	);

	and_ii n_2608_ (
		.a(n_0466_),
		.b(n_0449_),
		.c(n_0467_)
	);

	or_bi n_2609_ (
		.a(new_net_744),
		.b(new_net_1841),
		.c(n_0468_)
	);

	and_bi n_2610_ (
		.a(new_net_745),
		.b(new_net_1842),
		.c(n_0469_)
	);

	and_bi n_2611_ (
		.a(n_0468_),
		.b(n_0469_),
		.c(new_net_2527)
	);

	and_bi n_2612_ (
		.a(new_net_1821),
		.b(new_net_1008),
		.c(n_0470_)
	);

	or_bb n_2613_ (
		.a(n_0470_),
		.b(new_net_894),
		.c(n_0471_)
	);

	and_bi n_2614_ (
		.a(new_net_543),
		.b(new_net_670),
		.c(n_0472_)
	);

	and_bi n_2615_ (
		.a(new_net_674),
		.b(new_net_546),
		.c(n_0473_)
	);

	and_ii n_2616_ (
		.a(n_0473_),
		.b(n_0472_),
		.c(n_0474_)
	);

	and_bi n_2617_ (
		.a(new_net_878),
		.b(new_net_1566),
		.c(n_0475_)
	);

	and_bi n_2618_ (
		.a(new_net_1567),
		.b(new_net_877),
		.c(n_0476_)
	);

	or_bb n_2619_ (
		.a(n_0476_),
		.b(n_0475_),
		.c(n_0477_)
	);

	and_ii n_2620_ (
		.a(new_net_577),
		.b(new_net_1484),
		.c(n_0478_)
	);

	and_bi n_2621_ (
		.a(new_net_604),
		.b(new_net_2460),
		.c(n_0479_)
	);

	and_bi n_2622_ (
		.a(new_net_535),
		.b(new_net_289),
		.c(n_0480_)
	);

	and_bi n_2623_ (
		.a(new_net_290),
		.b(new_net_534),
		.c(n_0481_)
	);

	and_ii n_2624_ (
		.a(n_0481_),
		.b(n_0480_),
		.c(n_0482_)
	);

	and_bb n_2625_ (
		.a(new_net_675),
		.b(new_net_493),
		.c(n_0483_)
	);

	and_ii n_2626_ (
		.a(new_net_2461),
		.b(new_net_350),
		.c(n_0484_)
	);

	and_bi n_2627_ (
		.a(new_net_481),
		.b(new_net_494),
		.c(n_0485_)
	);

	and_ii n_2628_ (
		.a(new_net_326),
		.b(new_net_1369),
		.c(n_0486_)
	);

	and_bi n_2629_ (
		.a(new_net_1370),
		.b(new_net_1205),
		.c(n_0487_)
	);

	or_bb n_2630_ (
		.a(n_0487_),
		.b(n_0486_),
		.c(n_0488_)
	);

	and_bi n_2631_ (
		.a(new_net_780),
		.b(new_net_536),
		.c(n_0489_)
	);

	and_bi n_2632_ (
		.a(new_net_537),
		.b(new_net_777),
		.c(n_0490_)
	);

	or_bb n_2633_ (
		.a(n_0490_),
		.b(n_0489_),
		.c(n_0491_)
	);

	and_ii n_2634_ (
		.a(new_net_600),
		.b(new_net_439),
		.c(n_0492_)
	);

	and_bb n_2635_ (
		.a(new_net_601),
		.b(new_net_440),
		.c(n_0493_)
	);

	and_ii n_2636_ (
		.a(n_0493_),
		.b(n_0492_),
		.c(n_0494_)
	);

	and_bb n_2637_ (
		.a(new_net_1861),
		.b(new_net_408),
		.c(n_0495_)
	);

	and_ii n_2638_ (
		.a(new_net_1862),
		.b(new_net_409),
		.c(n_0496_)
	);

	or_bb n_2639_ (
		.a(n_0496_),
		.b(n_0495_),
		.c(n_0497_)
	);

	and_bi n_2640_ (
		.a(new_net_1668),
		.b(new_net_2462),
		.c(n_0498_)
	);

	and_bi n_2641_ (
		.a(new_net_437),
		.b(new_net_325),
		.c(n_0499_)
	);

	and_ii n_2642_ (
		.a(new_net_1315),
		.b(new_net_2463),
		.c(n_0500_)
	);

	and_bi n_2643_ (
		.a(new_net_791),
		.b(new_net_782),
		.c(n_0501_)
	);

	and_bi n_2644_ (
		.a(new_net_778),
		.b(new_net_792),
		.c(n_0502_)
	);

	and_ii n_2645_ (
		.a(n_0502_),
		.b(n_0501_),
		.c(n_0503_)
	);

	and_bi n_2646_ (
		.a(new_net_858),
		.b(new_net_478),
		.c(n_0504_)
	);

	and_bi n_2647_ (
		.a(new_net_483),
		.b(new_net_859),
		.c(n_0505_)
	);

	and_ii n_2648_ (
		.a(n_0505_),
		.b(n_0504_),
		.c(n_0506_)
	);

	and_bi n_2649_ (
		.a(new_net_922),
		.b(new_net_351),
		.c(n_0507_)
	);

	and_bi n_2650_ (
		.a(new_net_352),
		.b(new_net_923),
		.c(n_0508_)
	);

	or_bb n_2651_ (
		.a(n_0508_),
		.b(n_0507_),
		.c(n_0509_)
	);

	and_bi n_2652_ (
		.a(new_net_1557),
		.b(new_net_2464),
		.c(n_0510_)
	);

	or_bb n_2653_ (
		.a(n_0510_),
		.b(n_0498_),
		.c(n_0511_)
	);

	or_bb n_2654_ (
		.a(new_net_1868),
		.b(new_net_98),
		.c(n_0512_)
	);

	and_bb n_2655_ (
		.a(new_net_1869),
		.b(new_net_99),
		.c(n_0513_)
	);

	and_bi n_2656_ (
		.a(n_0512_),
		.b(n_0513_),
		.c(n_0514_)
	);

	or_bi n_2657_ (
		.a(new_net_22),
		.b(new_net_589),
		.c(n_0515_)
	);

	and_bi n_2658_ (
		.a(new_net_23),
		.b(new_net_590),
		.c(n_0516_)
	);

	and_bi n_2659_ (
		.a(n_0515_),
		.b(n_0516_),
		.c(new_net_2529)
	);

	and_bb n_2660_ (
		.a(new_net_701),
		.b(new_net_451),
		.c(n_0517_)
	);

	and_ii n_2661_ (
		.a(new_net_2465),
		.b(new_net_804),
		.c(n_0518_)
	);

	and_bb n_2662_ (
		.a(new_net_1152),
		.b(new_net_1138),
		.c(n_0519_)
	);

	or_bb n_2663_ (
		.a(n_0519_),
		.b(n_0518_),
		.c(n_0520_)
	);

	and_bi n_2664_ (
		.a(new_net_968),
		.b(new_net_1497),
		.c(n_0521_)
	);

	and_bi n_2665_ (
		.a(new_net_1498),
		.b(new_net_969),
		.c(n_0522_)
	);

	and_ii n_2666_ (
		.a(n_0522_),
		.b(n_0521_),
		.c(n_0523_)
	);

	and_bb n_2667_ (
		.a(new_net_1255),
		.b(new_net_1202),
		.c(n_0524_)
	);

	and_ii n_2668_ (
		.a(new_net_1256),
		.b(new_net_1203),
		.c(n_0525_)
	);

	and_ii n_2669_ (
		.a(n_0525_),
		.b(n_0524_),
		.c(n_0526_)
	);

	or_bb n_2670_ (
		.a(new_net_1832),
		.b(new_net_1218),
		.c(n_0527_)
	);

	and_bb n_2671_ (
		.a(new_net_1833),
		.b(new_net_1219),
		.c(n_0528_)
	);

	and_bi n_2672_ (
		.a(n_0527_),
		.b(n_0528_),
		.c(n_0529_)
	);

	and_bi n_2673_ (
		.a(new_net_401),
		.b(new_net_2466),
		.c(n_0530_)
	);

	and_bi n_2674_ (
		.a(new_net_447),
		.b(new_net_891),
		.c(n_0531_)
	);

	and_bi n_2675_ (
		.a(new_net_1954),
		.b(n_0531_),
		.c(n_0532_)
	);

	and_bi n_2676_ (
		.a(new_net_357),
		.b(new_net_708),
		.c(n_0533_)
	);

	and_bi n_2677_ (
		.a(new_net_709),
		.b(new_net_356),
		.c(n_0534_)
	);

	or_bb n_2678_ (
		.a(n_0534_),
		.b(n_0533_),
		.c(n_0535_)
	);

	and_bi n_2679_ (
		.a(new_net_892),
		.b(new_net_1154),
		.c(n_0536_)
	);

	and_bi n_2680_ (
		.a(new_net_1153),
		.b(new_net_450),
		.c(n_0537_)
	);

	and_ii n_2681_ (
		.a(new_net_2467),
		.b(n_0536_),
		.c(n_0538_)
	);

	and_bi n_2682_ (
		.a(new_net_1318),
		.b(new_net_967),
		.c(n_0539_)
	);

	and_bi n_2683_ (
		.a(new_net_971),
		.b(new_net_1319),
		.c(n_0540_)
	);

	and_ii n_2684_ (
		.a(n_0540_),
		.b(n_0539_),
		.c(n_0541_)
	);

	or_bi n_2685_ (
		.a(new_net_1540),
		.b(new_net_1657),
		.c(n_0542_)
	);

	and_bi n_2686_ (
		.a(new_net_1541),
		.b(new_net_1658),
		.c(n_0543_)
	);

	or_bi n_2687_ (
		.a(n_0543_),
		.b(n_0542_),
		.c(n_0544_)
	);

	and_bi n_2688_ (
		.a(new_net_2468),
		.b(new_net_399),
		.c(n_0545_)
	);

	and_ii n_2689_ (
		.a(n_0545_),
		.b(n_0530_),
		.c(n_0546_)
	);

	and_bi n_2690_ (
		.a(new_net_789),
		.b(new_net_1544),
		.c(n_0547_)
	);

	and_ii n_2691_ (
		.a(new_net_2469),
		.b(new_net_21),
		.c(n_0548_)
	);

	and_bi n_2692_ (
		.a(new_net_1112),
		.b(new_net_1627),
		.c(n_0549_)
	);

	and_bi n_2693_ (
		.a(new_net_1628),
		.b(new_net_1113),
		.c(n_0550_)
	);

	and_ii n_2694_ (
		.a(n_0550_),
		.b(n_0549_),
		.c(n_0551_)
	);

	and_bb n_2695_ (
		.a(new_net_930),
		.b(new_net_607),
		.c(n_0552_)
	);

	and_ii n_2696_ (
		.a(new_net_931),
		.b(new_net_608),
		.c(n_0553_)
	);

	and_ii n_2697_ (
		.a(n_0553_),
		.b(n_0552_),
		.c(n_0554_)
	);

	and_bi n_2698_ (
		.a(new_net_304),
		.b(new_net_1945),
		.c(n_0555_)
	);

	and_bi n_2699_ (
		.a(new_net_1946),
		.b(new_net_306),
		.c(n_0556_)
	);

	and_ii n_2700_ (
		.a(n_0556_),
		.b(n_0555_),
		.c(n_0557_)
	);

	and_bi n_2701_ (
		.a(new_net_432),
		.b(new_net_2470),
		.c(n_0558_)
	);

	and_bi n_2702_ (
		.a(new_net_1597),
		.b(new_net_305),
		.c(n_0559_)
	);

	or_bb n_2703_ (
		.a(n_0559_),
		.b(new_net_1535),
		.c(n_0560_)
	);

	and_bi n_2704_ (
		.a(new_net_30),
		.b(new_net_581),
		.c(n_0561_)
	);

	and_ii n_2705_ (
		.a(new_net_1360),
		.b(new_net_1241),
		.c(n_0562_)
	);

	and_bi n_2706_ (
		.a(new_net_1533),
		.b(new_net_1818),
		.c(n_0563_)
	);

	or_bb n_2707_ (
		.a(n_0563_),
		.b(new_net_2471),
		.c(n_0564_)
	);

	and_ii n_2708_ (
		.a(new_net_1237),
		.b(new_net_1207),
		.c(n_0565_)
	);

	and_bb n_2709_ (
		.a(new_net_1238),
		.b(new_net_1208),
		.c(n_0566_)
	);

	and_ii n_2710_ (
		.a(n_0566_),
		.b(n_0565_),
		.c(n_0567_)
	);

	or_bb n_2711_ (
		.a(new_net_1308),
		.b(new_net_1164),
		.c(n_0568_)
	);

	and_bb n_2712_ (
		.a(new_net_1309),
		.b(new_net_1165),
		.c(n_0569_)
	);

	or_bi n_2713_ (
		.a(n_0569_),
		.b(n_0568_),
		.c(n_0570_)
	);

	and_bi n_2714_ (
		.a(new_net_2472),
		.b(new_net_429),
		.c(n_0571_)
	);

	and_ii n_2715_ (
		.a(n_0571_),
		.b(n_0558_),
		.c(n_0572_)
	);

	and_ii n_2716_ (
		.a(new_net_897),
		.b(new_net_458),
		.c(n_0573_)
	);

	or_bi n_2717_ (
		.a(new_net_2473),
		.b(new_net_1010),
		.c(n_0574_)
	);

	and_bb n_2718_ (
		.a(new_net_1477),
		.b(new_net_609),
		.c(n_0575_)
	);

	and_ii n_2719_ (
		.a(new_net_1478),
		.b(new_net_610),
		.c(n_0576_)
	);

	and_ii n_2720_ (
		.a(n_0576_),
		.b(n_0575_),
		.c(n_0577_)
	);

	and_ii n_2721_ (
		.a(new_net_1128),
		.b(new_net_340),
		.c(n_0578_)
	);

	and_bb n_2722_ (
		.a(new_net_1129),
		.b(new_net_341),
		.c(n_0579_)
	);

	or_bb n_2723_ (
		.a(n_0579_),
		.b(n_0578_),
		.c(new_net_2539)
	);

	and_ii n_2724_ (
		.a(new_net_508),
		.b(new_net_1275),
		.c(n_0580_)
	);

	and_bi n_2725_ (
		.a(new_net_507),
		.b(new_net_704),
		.c(n_0581_)
	);

	and_ii n_2726_ (
		.a(new_net_2474),
		.b(n_0580_),
		.c(n_0582_)
	);

	and_ii n_2727_ (
		.a(new_net_1638),
		.b(new_net_1513),
		.c(n_0583_)
	);

	and_bb n_2728_ (
		.a(new_net_1639),
		.b(new_net_1510),
		.c(n_0584_)
	);

	or_bb n_2729_ (
		.a(n_0584_),
		.b(n_0583_),
		.c(n_0585_)
	);

	and_ii n_2730_ (
		.a(new_net_1813),
		.b(new_net_1754),
		.c(n_0586_)
	);

	and_bi n_2731_ (
		.a(new_net_1952),
		.b(new_net_2475),
		.c(n_0587_)
	);

	or_bb n_2732_ (
		.a(new_net_1735),
		.b(new_net_471),
		.c(n_0588_)
	);

	and_bi n_2733_ (
		.a(new_net_1738),
		.b(new_net_1784),
		.c(n_0589_)
	);

	and_bi n_2734_ (
		.a(n_0588_),
		.b(n_0589_),
		.c(n_0590_)
	);

	and_ii n_2735_ (
		.a(new_net_1791),
		.b(new_net_1694),
		.c(n_0591_)
	);

	and_bb n_2736_ (
		.a(new_net_1792),
		.b(new_net_1695),
		.c(n_0592_)
	);

	and_ii n_2737_ (
		.a(n_0592_),
		.b(n_0591_),
		.c(n_0593_)
	);

	or_bb n_2738_ (
		.a(new_net_1036),
		.b(new_net_412),
		.c(n_0594_)
	);

	and_bi n_2739_ (
		.a(new_net_587),
		.b(new_net_906),
		.c(n_0595_)
	);

	and_bi n_2740_ (
		.a(new_net_905),
		.b(new_net_705),
		.c(n_0596_)
	);

	or_bb n_2741_ (
		.a(n_0596_),
		.b(n_0595_),
		.c(n_0597_)
	);

	or_bi n_2742_ (
		.a(new_net_2476),
		.b(new_net_1399),
		.c(n_0598_)
	);

	and_bi n_2743_ (
		.a(new_net_1512),
		.b(new_net_852),
		.c(n_0599_)
	);

	and_bb n_2744_ (
		.a(new_net_853),
		.b(new_net_556),
		.c(n_0600_)
	);

	and_bi n_2745_ (
		.a(new_net_2477),
		.b(new_net_1514),
		.c(n_0601_)
	);

	and_ii n_2746_ (
		.a(n_0601_),
		.b(new_net_2478),
		.c(n_0602_)
	);

	and_ii n_2747_ (
		.a(new_net_83),
		.b(new_net_1736),
		.c(n_0603_)
	);

	and_bb n_2748_ (
		.a(new_net_84),
		.b(new_net_1737),
		.c(n_0604_)
	);

	or_bb n_2749_ (
		.a(n_0604_),
		.b(n_0603_),
		.c(n_0605_)
	);

	and_bi n_2750_ (
		.a(new_net_411),
		.b(new_net_117),
		.c(n_0606_)
	);

	or_bb n_2751_ (
		.a(n_0606_),
		.b(new_net_1680),
		.c(n_0607_)
	);

	and_bi n_2752_ (
		.a(new_net_2479),
		.b(n_0607_),
		.c(n_0608_)
	);

	and_bb n_2753_ (
		.a(new_net_1037),
		.b(new_net_421),
		.c(n_0609_)
	);

	or_ii n_2754_ (
		.a(new_net_292),
		.b(new_net_1677),
		.c(n_0610_)
	);

	and_bi n_2755_ (
		.a(new_net_118),
		.b(new_net_2480),
		.c(n_0611_)
	);

	or_bb n_2756_ (
		.a(n_0611_),
		.b(new_net_2481),
		.c(n_0612_)
	);

	or_bb n_2757_ (
		.a(new_net_2482),
		.b(n_0608_),
		.c(n_0613_)
	);

	and_bb n_2758_ (
		.a(new_net_1470),
		.b(new_net_739),
		.c(n_0614_)
	);

	or_bb n_2759_ (
		.a(new_net_2483),
		.b(new_net_362),
		.c(n_0615_)
	);

	and_bi n_2760_ (
		.a(new_net_1764),
		.b(new_net_1348),
		.c(n_0616_)
	);

	and_bb n_2761_ (
		.a(new_net_1284),
		.b(new_net_1060),
		.c(n_0617_)
	);

	and_bi n_2762_ (
		.a(new_net_1339),
		.b(new_net_2484),
		.c(n_0618_)
	);

	and_bi n_2763_ (
		.a(new_net_1160),
		.b(new_net_105),
		.c(n_0619_)
	);

	and_bi n_2764_ (
		.a(new_net_107),
		.b(new_net_1161),
		.c(n_0620_)
	);

	and_ii n_2765_ (
		.a(n_0620_),
		.b(n_0619_),
		.c(n_0621_)
	);

	and_bi n_2766_ (
		.a(new_net_686),
		.b(new_net_964),
		.c(n_0622_)
	);

	and_bi n_2767_ (
		.a(new_net_965),
		.b(new_net_689),
		.c(n_0623_)
	);

	or_bb n_2768_ (
		.a(n_0623_),
		.b(n_0622_),
		.c(n_0624_)
	);

	and_ii n_2769_ (
		.a(new_net_756),
		.b(new_net_547),
		.c(n_0625_)
	);

	and_bb n_2770_ (
		.a(new_net_757),
		.b(new_net_548),
		.c(n_0626_)
	);

	or_bb n_2771_ (
		.a(n_0626_),
		.b(new_net_963),
		.c(n_0627_)
	);

	or_bb n_2772_ (
		.a(n_0627_),
		.b(new_net_2485),
		.c(n_0628_)
	);

	and_ii n_2773_ (
		.a(new_net_1471),
		.b(new_net_1455),
		.c(n_0629_)
	);

	and_ii n_2774_ (
		.a(new_net_1065),
		.b(new_net_1613),
		.c(n_0630_)
	);

	or_bi n_2775_ (
		.a(new_net_1260),
		.b(new_net_1763),
		.c(n_0631_)
	);

	and_bi n_2776_ (
		.a(new_net_1612),
		.b(n_0631_),
		.c(n_0632_)
	);

	and_ii n_2777_ (
		.a(n_0632_),
		.b(new_net_2486),
		.c(n_0633_)
	);

	or_bi n_2778_ (
		.a(new_net_860),
		.b(new_net_978),
		.c(n_0634_)
	);

	and_bi n_2779_ (
		.a(new_net_861),
		.b(new_net_979),
		.c(n_0635_)
	);

	and_bi n_2780_ (
		.a(n_0634_),
		.b(n_0635_),
		.c(n_0636_)
	);

	and_bi n_2781_ (
		.a(new_net_681),
		.b(new_net_687),
		.c(n_0637_)
	);

	and_bi n_2782_ (
		.a(new_net_688),
		.b(new_net_680),
		.c(n_0638_)
	);

	or_bb n_2783_ (
		.a(n_0638_),
		.b(n_0637_),
		.c(n_0639_)
	);

	or_bi n_2784_ (
		.a(new_net_1253),
		.b(new_net_1758),
		.c(n_0640_)
	);

	and_bi n_2785_ (
		.a(new_net_1254),
		.b(new_net_1759),
		.c(n_0641_)
	);

	or_bb n_2786_ (
		.a(n_0641_),
		.b(new_net_1679),
		.c(n_0642_)
	);

	and_bi n_2787_ (
		.a(new_net_2487),
		.b(n_0642_),
		.c(n_0643_)
	);

	and_bi n_2788_ (
		.a(new_net_2488),
		.b(n_0643_),
		.c(n_0644_)
	);

	or_bi n_2789_ (
		.a(new_net_1174),
		.b(new_net_1077),
		.c(n_0645_)
	);

	and_bi n_2790_ (
		.a(new_net_1173),
		.b(new_net_1073),
		.c(n_0646_)
	);

	and_bi n_2791_ (
		.a(n_0645_),
		.b(n_0646_),
		.c(n_0647_)
	);

	and_ii n_2792_ (
		.a(new_net_835),
		.b(new_net_503),
		.c(n_0648_)
	);

	and_bb n_2793_ (
		.a(new_net_836),
		.b(new_net_504),
		.c(n_0649_)
	);

	and_ii n_2794_ (
		.a(n_0649_),
		.b(n_0648_),
		.c(n_0650_)
	);

	or_bb n_2795_ (
		.a(new_net_1280),
		.b(new_net_653),
		.c(n_0651_)
	);

	and_bb n_2796_ (
		.a(new_net_1281),
		.b(new_net_654),
		.c(n_0652_)
	);

	and_bi n_2797_ (
		.a(n_0651_),
		.b(n_0652_),
		.c(new_net_2541)
	);

	and_bi n_2798_ (
		.a(new_net_453),
		.b(new_net_1102),
		.c(new_net_2554)
	);

	and_bi n_2799_ (
		.a(new_net_1135),
		.b(new_net_294),
		.c(new_net_2533)
	);

	and_bi n_2800_ (
		.a(new_net_455),
		.b(new_net_1101),
		.c(new_net_2552)
	);

	and_bi n_2801_ (
		.a(new_net_454),
		.b(new_net_1103),
		.c(new_net_2519)
	);

	spl2 new_net_8_v_fanout (
		.a(new_net_8),
		.b(N10838),
		.c(N10837)
	);

	bfr new_net_2580_bfr_after (
		.din(new_net_9),
		.dout(new_net_2580)
	);

	bfr new_net_2581_bfr_after (
		.din(new_net_2580),
		.dout(new_net_2581)
	);

	spl2 new_net_9_v_fanout (
		.a(new_net_2581),
		.b(N10840),
		.c(N10839)
	);

	spl4L n_0178__v_fanout (
		.a(n_0178_),
		.b(new_net_1102),
		.c(new_net_1103),
		.d(new_net_1101),
		.e(new_net_1100)
	);

	spl2 n_0471__v_fanout (
		.a(n_0471_),
		.b(new_net_23),
		.c(new_net_22)
	);

	spl2 n_0377__v_fanout (
		.a(n_0377_),
		.b(new_net_665),
		.c(new_net_664)
	);

	spl2 n_0177__v_fanout (
		.a(n_0177_),
		.b(new_net_1188),
		.c(new_net_1187)
	);

	spl4L new_net_2182_v_fanout (
		.a(new_net_2182),
		.b(new_net_1822),
		.c(new_net_1820),
		.d(new_net_1823),
		.e(new_net_1821)
	);

	bfr new_net_2582_bfr_after (
		.din(n_0514_),
		.dout(new_net_2582)
	);

	bfr new_net_2583_bfr_after (
		.din(new_net_2582),
		.dout(new_net_2583)
	);

	bfr new_net_2584_bfr_after (
		.din(new_net_2583),
		.dout(new_net_2584)
	);

	spl2 n_0514__v_fanout (
		.a(new_net_2584),
		.b(new_net_590),
		.c(new_net_589)
	);

	spl2 n_0118__v_fanout (
		.a(n_0118_),
		.b(new_net_718),
		.c(new_net_717)
	);

	bfr new_net_2585_bfr_before (
		.din(new_net_2585),
		.dout(new_net_1819)
	);

	spl2 n_0176__v_fanout (
		.a(n_0176_),
		.b(new_net_2182),
		.c(new_net_2585)
	);

	spl2 n_0124__v_fanout (
		.a(n_0124_),
		.b(new_net_1548),
		.c(new_net_1547)
	);

	spl2 n_0131__v_fanout (
		.a(n_0131_),
		.b(new_net_496),
		.c(new_net_495)
	);

	spl2 n_0511__v_fanout (
		.a(n_0511_),
		.b(new_net_1869),
		.c(new_net_1868)
	);

	spl4L new_net_1961_v_fanout (
		.a(new_net_1961),
		.b(N388),
		.c(N889),
		.d(N1490),
		.e(N387)
	);

	spl2 n_0128__v_fanout (
		.a(n_0128_),
		.b(new_net_925),
		.c(new_net_924)
	);

	spl3L n_0115__v_fanout (
		.a(n_0115_),
		.b(new_net_663),
		.c(new_net_661),
		.d(new_net_662)
	);

	spl2 n_0075__v_fanout (
		.a(n_0075_),
		.b(new_net_1571),
		.c(new_net_1570)
	);

	spl3L n_0074__v_fanout (
		.a(n_0074_),
		.b(new_net_1557),
		.c(new_net_1555),
		.d(new_net_1556)
	);

	spl2 new_net_2068_v_fanout (
		.a(new_net_2068),
		.b(new_net_1007),
		.c(new_net_1008)
	);

	spl2 new_net_2133_v_fanout (
		.a(new_net_2133),
		.b(new_net_779),
		.c(new_net_776)
	);

	spl3L n_0076__v_fanout (
		.a(n_0076_),
		.b(new_net_1669),
		.c(new_net_1667),
		.d(new_net_1668)
	);

	bfr new_net_2586_bfr_before (
		.din(new_net_2586),
		.dout(new_net_894)
	);

	spl2 new_net_2067_v_fanout (
		.a(new_net_2067),
		.b(new_net_2586),
		.c(new_net_895)
	);

	spl2 new_net_2127_v_fanout (
		.a(new_net_2127),
		.b(new_net_576),
		.c(new_net_575)
	);

	spl2 new_net_2130_v_fanout (
		.a(new_net_2130),
		.b(new_net_672),
		.c(new_net_669)
	);

	spl2 new_net_2126_v_fanout (
		.a(new_net_2126),
		.b(new_net_544),
		.c(new_net_545)
	);

	spl2 n_0073__v_fanout (
		.a(n_0073_),
		.b(new_net_1337),
		.c(new_net_1336)
	);

	bfr new_net_2587_bfr_before (
		.din(new_net_2587),
		.dout(new_net_2130)
	);

	spl2 new_net_2129_v_fanout (
		.a(new_net_2129),
		.b(new_net_2587),
		.c(new_net_671)
	);

	spl2 n_0369__v_fanout (
		.a(n_0369_),
		.b(new_net_691),
		.c(new_net_690)
	);

	spl2 n_0467__v_fanout (
		.a(n_0467_),
		.b(new_net_1842),
		.c(new_net_1841)
	);

	spl3L n_0072__v_fanout (
		.a(n_0072_),
		.b(new_net_1223),
		.c(new_net_1222),
		.d(new_net_1224)
	);

	spl2 n_0364__v_fanout (
		.a(n_0364_),
		.b(new_net_568),
		.c(new_net_567)
	);

	spl2 new_net_2122_v_fanout (
		.a(new_net_2122),
		.b(new_net_1485),
		.c(new_net_1482)
	);

	bfr new_net_2588_bfr_after (
		.din(n_0434_),
		.dout(new_net_2588)
	);

	spl2 n_0434__v_fanout (
		.a(new_net_2588),
		.b(new_net_745),
		.c(new_net_744)
	);

	spl2 n_0085__v_fanout (
		.a(n_0085_),
		.b(new_net_844),
		.c(new_net_843)
	);

	spl2 new_net_2102_v_fanout (
		.a(new_net_2102),
		.b(new_net_532),
		.c(new_net_530)
	);

	spl3L new_net_2180_v_fanout (
		.a(new_net_2180),
		.b(new_net_1046),
		.c(new_net_1044),
		.d(new_net_1047)
	);

	spl2 n_0088__v_fanout (
		.a(n_0088_),
		.b(new_net_1829),
		.c(new_net_1828)
	);

	spl2 n_0095__v_fanout (
		.a(n_0095_),
		.b(new_net_76),
		.c(new_net_75)
	);

	spl4L new_net_2181_v_fanout (
		.a(new_net_2181),
		.b(new_net_1050),
		.c(new_net_1048),
		.d(new_net_1049),
		.e(new_net_1045)
	);

	spl2 n_0070__v_fanout (
		.a(n_0070_),
		.b(new_net_2181),
		.c(new_net_2180)
	);

	spl2 n_0092__v_fanout (
		.a(n_0092_),
		.b(new_net_1940),
		.c(new_net_1939)
	);

	spl2 n_0429__v_fanout (
		.a(n_0429_),
		.b(new_net_34),
		.c(new_net_33)
	);

	spl2 n_0083__v_fanout (
		.a(n_0083_),
		.b(new_net_636),
		.c(new_net_635)
	);

	spl2 new_net_2135_v_fanout (
		.a(new_net_2135),
		.b(new_net_475),
		.c(new_net_472)
	);

	spl2 new_net_2136_v_fanout (
		.a(new_net_2136),
		.b(new_net_1380),
		.c(new_net_1378)
	);

	spl2 new_net_2157_v_fanout (
		.a(new_net_2157),
		.b(new_net_1374),
		.c(new_net_1375)
	);

	spl2 n_0020__v_fanout (
		.a(n_0020_),
		.b(new_net_959),
		.c(new_net_958)
	);

	spl2 new_net_2155_v_fanout (
		.a(new_net_2155),
		.b(new_net_1653),
		.c(new_net_1650)
	);

	spl2 new_net_2124_v_fanout (
		.a(new_net_2124),
		.b(new_net_1858),
		.c(new_net_1859)
	);

	spl2 new_net_2158_v_fanout (
		.a(new_net_2158),
		.b(new_net_1682),
		.c(new_net_1683)
	);

	spl3L new_net_2178_v_fanout (
		.a(new_net_2178),
		.b(new_net_331),
		.c(new_net_329),
		.d(new_net_332)
	);

	spl4L new_net_2179_v_fanout (
		.a(new_net_2179),
		.b(new_net_335),
		.c(new_net_333),
		.d(new_net_334),
		.e(new_net_330)
	);

	spl2 new_net_2137_v_fanout (
		.a(new_net_2137),
		.b(new_net_1908),
		.c(new_net_1906)
	);

	spl2 n_0019__v_fanout (
		.a(n_0019_),
		.b(new_net_2179),
		.c(new_net_2178)
	);

	spl2 new_net_2159_v_fanout (
		.a(new_net_2159),
		.b(new_net_1704),
		.c(new_net_1703)
	);

	spl2 new_net_2147_v_fanout (
		.a(new_net_2147),
		.b(new_net_1636),
		.c(new_net_1634)
	);

	spl3L n_0017__v_fanout (
		.a(n_0017_),
		.b(new_net_116),
		.c(new_net_114),
		.d(new_net_115)
	);

	spl2 n_0387__v_fanout (
		.a(n_0387_),
		.b(new_net_1871),
		.c(new_net_1870)
	);

	spl2 n_0392__v_fanout (
		.a(n_0392_),
		.b(new_net_646),
		.c(new_net_645)
	);

	spl2 n_0546__v_fanout (
		.a(n_0546_),
		.b(new_net_341),
		.c(new_net_340)
	);

	bfr new_net_2589_bfr_after (
		.din(n_0577_),
		.dout(new_net_2589)
	);

	bfr new_net_2590_bfr_after (
		.din(new_net_2589),
		.dout(new_net_2590)
	);

	spl2 n_0577__v_fanout (
		.a(new_net_2590),
		.b(new_net_1129),
		.c(new_net_1128)
	);

	spl2 new_net_2139_v_fanout (
		.a(new_net_2139),
		.b(new_net_970),
		.c(new_net_966)
	);

	spl2 n_0155__v_fanout (
		.a(n_0155_),
		.b(new_net_1416),
		.c(new_net_1415)
	);

	spl2 new_net_2140_v_fanout (
		.a(new_net_2140),
		.b(new_net_1499),
		.c(new_net_1496)
	);

	spl4L new_net_2177_v_fanout (
		.a(new_net_2177),
		.b(new_net_400),
		.c(new_net_397),
		.d(new_net_401),
		.e(new_net_398)
	);

	spl3L new_net_2176_v_fanout (
		.a(new_net_2176),
		.b(new_net_399),
		.c(new_net_395),
		.d(new_net_396)
	);

	spl2 n_0015__v_fanout (
		.a(n_0015_),
		.b(new_net_2177),
		.c(new_net_2176)
	);

	spl2 n_0158__v_fanout (
		.a(n_0158_),
		.b(new_net_1729),
		.c(new_net_1728)
	);

	spl2 new_net_2160_v_fanout (
		.a(new_net_2160),
		.b(new_net_1185),
		.c(new_net_1186)
	);

	spl2 n_0572__v_fanout (
		.a(n_0572_),
		.b(new_net_610),
		.c(new_net_609)
	);

	spl2 n_0149__v_fanout (
		.a(n_0149_),
		.b(new_net_802),
		.c(new_net_801)
	);

	spl2 new_net_2151_v_fanout (
		.a(new_net_2151),
		.b(new_net_900),
		.c(new_net_896)
	);

	spl2 n_0006__v_fanout (
		.a(n_0006_),
		.b(new_net_562),
		.c(new_net_561)
	);

	spl2 new_net_2148_v_fanout (
		.a(new_net_2148),
		.b(new_net_1167),
		.c(new_net_1168)
	);

	spl3L n_0140__v_fanout (
		.a(n_0140_),
		.b(new_net_1622),
		.c(new_net_1621),
		.d(new_net_1623)
	);

	spl2 n_0650__v_fanout (
		.a(n_0650_),
		.b(new_net_1281),
		.c(new_net_1280)
	);

	spl2 new_net_2149_v_fanout (
		.a(new_net_2149),
		.b(new_net_457),
		.c(new_net_459)
	);

	bfr new_net_2591_bfr_after (
		.din(new_net_7),
		.dout(new_net_2591)
	);

	bfr new_net_2592_bfr_after (
		.din(new_net_2591),
		.dout(new_net_2592)
	);

	bfr new_net_2593_bfr_after (
		.din(new_net_2592),
		.dout(new_net_2593)
	);

	bfr new_net_2594_bfr_after (
		.din(new_net_2593),
		.dout(new_net_2594)
	);

	bfr new_net_2595_bfr_after (
		.din(new_net_2594),
		.dout(new_net_2595)
	);

	bfr new_net_2596_bfr_after (
		.din(new_net_2595),
		.dout(new_net_2596)
	);

	bfr new_net_2597_bfr_after (
		.din(new_net_2596),
		.dout(new_net_2597)
	);

	bfr new_net_2598_bfr_after (
		.din(new_net_2597),
		.dout(new_net_2598)
	);

	bfr new_net_2599_bfr_after (
		.din(new_net_2598),
		.dout(new_net_2599)
	);

	bfr new_net_2600_bfr_after (
		.din(new_net_2599),
		.dout(new_net_2600)
	);

	bfr new_net_2601_bfr_after (
		.din(new_net_2600),
		.dout(new_net_2601)
	);

	bfr new_net_2602_bfr_after (
		.din(new_net_2601),
		.dout(new_net_2602)
	);

	bfr new_net_2603_bfr_after (
		.din(new_net_2602),
		.dout(new_net_2603)
	);

	bfr new_net_2604_bfr_after (
		.din(new_net_2603),
		.dout(new_net_2604)
	);

	bfr new_net_2605_bfr_after (
		.din(new_net_2604),
		.dout(new_net_2605)
	);

	bfr new_net_2606_bfr_after (
		.din(new_net_2605),
		.dout(new_net_2606)
	);

	bfr new_net_2607_bfr_after (
		.din(new_net_2606),
		.dout(new_net_2607)
	);

	bfr new_net_2608_bfr_after (
		.din(new_net_2607),
		.dout(new_net_2608)
	);

	bfr new_net_2609_bfr_after (
		.din(new_net_2608),
		.dout(new_net_2609)
	);

	bfr new_net_2610_bfr_after (
		.din(new_net_2609),
		.dout(new_net_2610)
	);

	bfr new_net_2611_bfr_after (
		.din(new_net_2610),
		.dout(new_net_2611)
	);

	bfr new_net_2612_bfr_after (
		.din(new_net_2611),
		.dout(new_net_2612)
	);

	bfr new_net_2613_bfr_after (
		.din(new_net_2612),
		.dout(new_net_2613)
	);

	bfr new_net_2614_bfr_after (
		.din(new_net_2613),
		.dout(new_net_2614)
	);

	bfr new_net_2615_bfr_after (
		.din(new_net_2614),
		.dout(new_net_2615)
	);

	bfr new_net_2616_bfr_after (
		.din(new_net_2615),
		.dout(new_net_2616)
	);

	bfr new_net_2617_bfr_after (
		.din(new_net_2616),
		.dout(new_net_2617)
	);

	bfr new_net_2618_bfr_after (
		.din(new_net_2617),
		.dout(new_net_2618)
	);

	bfr new_net_2619_bfr_after (
		.din(new_net_2618),
		.dout(new_net_2619)
	);

	bfr new_net_2620_bfr_after (
		.din(new_net_2619),
		.dout(new_net_2620)
	);

	bfr new_net_2621_bfr_after (
		.din(new_net_2620),
		.dout(new_net_2621)
	);

	bfr new_net_2622_bfr_after (
		.din(new_net_2621),
		.dout(new_net_2622)
	);

	bfr new_net_2623_bfr_after (
		.din(new_net_2622),
		.dout(new_net_2623)
	);

	bfr new_net_2624_bfr_after (
		.din(new_net_2623),
		.dout(new_net_2624)
	);

	spl2 new_net_7_v_fanout (
		.a(new_net_2624),
		.b(N10103),
		.c(N10102)
	);

	spl2 n_0351__v_fanout (
		.a(n_0351_),
		.b(new_net_103),
		.c(new_net_102)
	);

	spl3L new_net_2174_v_fanout (
		.a(new_net_2174),
		.b(new_net_430),
		.c(new_net_426),
		.d(new_net_427)
	);

	spl2 n_0355__v_fanout (
		.a(n_0355_),
		.b(new_net_337),
		.c(new_net_336)
	);

	spl4L new_net_2175_v_fanout (
		.a(new_net_2175),
		.b(new_net_428),
		.c(new_net_432),
		.d(new_net_431),
		.e(new_net_429)
	);

	spl2 new_net_2162_v_fanout (
		.a(new_net_2162),
		.b(new_net_1783),
		.c(new_net_1782)
	);

	spl2 new_net_2161_v_fanout (
		.a(new_net_2161),
		.b(new_net_418),
		.c(new_net_419)
	);

	spl2 n_0346__v_fanout (
		.a(n_0346_),
		.b(new_net_32),
		.c(new_net_31)
	);

	spl2 n_0342__v_fanout (
		.a(n_0342_),
		.b(new_net_294),
		.c(new_net_293)
	);

	spl2 n_0005__v_fanout (
		.a(n_0005_),
		.b(new_net_2175),
		.c(new_net_2174)
	);

	bfr new_net_2625_bfr_after (
		.din(n_0613_),
		.dout(new_net_2625)
	);

	bfr new_net_2626_bfr_after (
		.din(new_net_2625),
		.dout(new_net_2626)
	);

	spl2 n_0613__v_fanout (
		.a(new_net_2626),
		.b(new_net_654),
		.c(new_net_653)
	);

	spl2 n_0644__v_fanout (
		.a(n_0644_),
		.b(new_net_504),
		.c(new_net_503)
	);

	spl2 new_net_2121_v_fanout (
		.a(new_net_2121),
		.b(new_net_1812),
		.c(new_net_1814)
	);

	spl2 n_0349__v_fanout (
		.a(n_0349_),
		.b(new_net_60),
		.c(new_net_59)
	);

	spl2 n_0560__v_fanout (
		.a(n_0560_),
		.b(new_net_1165),
		.c(new_net_1164)
	);

	spl4L new_net_2173_v_fanout (
		.a(new_net_2173),
		.b(new_net_442),
		.c(new_net_444),
		.d(new_net_443),
		.e(new_net_445)
	);

	spl2 n_0402__v_fanout (
		.a(n_0402_),
		.b(new_net_1385),
		.c(new_net_1384)
	);

	spl2 new_net_2156_v_fanout (
		.a(new_net_2156),
		.b(new_net_1278),
		.c(new_net_1279)
	);

	bfr new_net_2627_bfr_before (
		.din(new_net_2627),
		.dout(new_net_441)
	);

	spl2 n_1367__v_fanout (
		.a(n_1367_),
		.b(new_net_2173),
		.c(new_net_2627)
	);

	spl2 n_0484__v_fanout (
		.a(n_0484_),
		.b(new_net_409),
		.c(new_net_408)
	);

	spl2 n_0605__v_fanout (
		.a(n_0605_),
		.b(new_net_118),
		.c(new_net_117)
	);

	bfr new_net_2628_bfr_before (
		.din(new_net_2628),
		.dout(new_net_1680)
	);

	spl2 new_net_2066_v_fanout (
		.a(new_net_2066),
		.b(new_net_1679),
		.c(new_net_2628)
	);

	spl2 n_0593__v_fanout (
		.a(n_0593_),
		.b(new_net_1037),
		.c(new_net_1036)
	);

	spl3L n_0482__v_fanout (
		.a(n_0482_),
		.b(new_net_352),
		.c(new_net_350),
		.d(new_net_351)
	);

	spl3L n_0401__v_fanout (
		.a(n_0401_),
		.b(new_net_1574),
		.c(new_net_1572),
		.d(new_net_1573)
	);

	bfr new_net_2629_bfr_before (
		.din(new_net_2629),
		.dout(new_net_411)
	);

	spl3L n_1366__v_fanout (
		.a(n_1366_),
		.b(new_net_412),
		.c(new_net_410),
		.d(new_net_2629)
	);

	bfr new_net_2630_bfr_before (
		.din(new_net_2630),
		.dout(new_net_1598)
	);

	bfr new_net_2631_bfr_before (
		.din(new_net_2631),
		.dout(new_net_2630)
	);

	bfr new_net_2632_bfr_before (
		.din(new_net_2632),
		.dout(new_net_2631)
	);

	bfr new_net_2633_bfr_before (
		.din(new_net_2633),
		.dout(new_net_2632)
	);

	bfr new_net_2634_bfr_before (
		.din(new_net_2634),
		.dout(new_net_2633)
	);

	bfr new_net_2635_bfr_before (
		.din(new_net_2635),
		.dout(new_net_2634)
	);

	bfr new_net_2636_bfr_before (
		.din(new_net_2636),
		.dout(new_net_2635)
	);

	spl2 new_net_2169_v_fanout (
		.a(new_net_2169),
		.b(new_net_2636),
		.c(new_net_1597)
	);

	bfr new_net_2637_bfr_before (
		.din(new_net_2637),
		.dout(new_net_303)
	);

	bfr new_net_2638_bfr_before (
		.din(new_net_2638),
		.dout(new_net_2637)
	);

	bfr new_net_2639_bfr_before (
		.din(new_net_2639),
		.dout(new_net_2638)
	);

	bfr new_net_2640_bfr_before (
		.din(new_net_2640),
		.dout(new_net_2639)
	);

	bfr new_net_2641_bfr_before (
		.din(new_net_2641),
		.dout(new_net_2640)
	);

	bfr new_net_2642_bfr_before (
		.din(new_net_2642),
		.dout(new_net_2641)
	);

	bfr new_net_2643_bfr_before (
		.din(new_net_2643),
		.dout(new_net_2642)
	);

	bfr new_net_2644_bfr_before (
		.din(new_net_2644),
		.dout(new_net_2643)
	);

	spl4L n_0145__v_fanout (
		.a(n_0145_),
		.b(new_net_304),
		.c(new_net_305),
		.d(new_net_306),
		.e(new_net_2644)
	);

	spl2 n_1362__v_fanout (
		.a(n_1362_),
		.b(new_net_421),
		.c(new_net_420)
	);

	spl2 n_0639__v_fanout (
		.a(n_0639_),
		.b(new_net_1759),
		.c(new_net_1758)
	);

	spl2 n_0462__v_fanout (
		.a(n_0462_),
		.b(new_net_1903),
		.c(new_net_1902)
	);

	spl2 n_0264__v_fanout (
		.a(n_0264_),
		.b(new_net_1794),
		.c(new_net_1793)
	);

	bfr new_net_2645_bfr_after (
		.din(n_0567_),
		.dout(new_net_2645)
	);

	bfr new_net_2646_bfr_after (
		.din(new_net_2645),
		.dout(new_net_2646)
	);

	bfr new_net_2647_bfr_after (
		.din(new_net_2646),
		.dout(new_net_2647)
	);

	bfr new_net_2648_bfr_after (
		.din(new_net_2647),
		.dout(new_net_2648)
	);

	spl2 n_0567__v_fanout (
		.a(new_net_2648),
		.b(new_net_1309),
		.c(new_net_1308)
	);

	bfr new_net_2649_bfr_after (
		.din(n_0412_),
		.dout(new_net_2649)
	);

	bfr new_net_2650_bfr_after (
		.din(new_net_2649),
		.dout(new_net_2650)
	);

	bfr new_net_2651_bfr_after (
		.din(new_net_2650),
		.dout(new_net_2651)
	);

	spl2 n_0412__v_fanout (
		.a(new_net_2651),
		.b(new_net_951),
		.c(new_net_950)
	);

	bfr new_net_2652_bfr_after (
		.din(n_0494_),
		.dout(new_net_2652)
	);

	bfr new_net_2653_bfr_after (
		.din(new_net_2652),
		.dout(new_net_2653)
	);

	bfr new_net_2654_bfr_after (
		.din(new_net_2653),
		.dout(new_net_2654)
	);

	spl2 n_0494__v_fanout (
		.a(new_net_2654),
		.b(new_net_1862),
		.c(new_net_1861)
	);

	bfr new_net_2655_bfr_before (
		.din(new_net_2655),
		.dout(new_net_1757)
	);

	bfr new_net_2656_bfr_before (
		.din(new_net_2656),
		.dout(new_net_2655)
	);

	bfr new_net_2657_bfr_before (
		.din(new_net_2657),
		.dout(new_net_2656)
	);

	bfr new_net_2658_bfr_before (
		.din(new_net_2658),
		.dout(new_net_2657)
	);

	bfr new_net_2659_bfr_before (
		.din(new_net_2659),
		.dout(new_net_2658)
	);

	bfr new_net_2660_bfr_before (
		.din(new_net_2660),
		.dout(new_net_2659)
	);

	bfr new_net_2661_bfr_before (
		.din(new_net_2661),
		.dout(new_net_2660)
	);

	bfr new_net_2662_bfr_before (
		.din(new_net_2662),
		.dout(new_net_2661)
	);

	bfr new_net_2663_bfr_before (
		.din(new_net_2663),
		.dout(new_net_2662)
	);

	bfr new_net_2664_bfr_before (
		.din(new_net_2664),
		.dout(new_net_2663)
	);

	bfr new_net_2665_bfr_before (
		.din(new_net_2665),
		.dout(new_net_2664)
	);

	bfr new_net_2666_bfr_before (
		.din(new_net_2666),
		.dout(new_net_2665)
	);

	bfr new_net_2667_bfr_before (
		.din(new_net_2667),
		.dout(new_net_2666)
	);

	bfr new_net_2668_bfr_before (
		.din(new_net_2668),
		.dout(new_net_2667)
	);

	bfr new_net_2669_bfr_before (
		.din(new_net_2669),
		.dout(new_net_2668)
	);

	bfr new_net_2670_bfr_before (
		.din(new_net_2670),
		.dout(new_net_2669)
	);

	bfr new_net_2671_bfr_before (
		.din(new_net_2671),
		.dout(new_net_2670)
	);

	bfr new_net_2672_bfr_before (
		.din(new_net_2672),
		.dout(new_net_2671)
	);

	bfr new_net_2673_bfr_before (
		.din(new_net_2673),
		.dout(new_net_2672)
	);

	bfr new_net_2674_bfr_before (
		.din(new_net_2674),
		.dout(new_net_2673)
	);

	spl2 n_0060__v_fanout (
		.a(n_0060_),
		.b(new_net_2674),
		.c(new_net_1756)
	);

	bfr new_net_2675_bfr_before (
		.din(new_net_2675),
		.dout(new_net_2066)
	);

	bfr new_net_2676_bfr_before (
		.din(new_net_2676),
		.dout(new_net_2675)
	);

	spl3L new_net_2065_v_fanout (
		.a(new_net_2065),
		.b(new_net_1677),
		.c(new_net_1678),
		.d(new_net_2676)
	);

	spl2 n_0624__v_fanout (
		.a(n_0624_),
		.b(new_net_757),
		.c(new_net_756)
	);

	spl2 n_0602__v_fanout (
		.a(n_0602_),
		.b(new_net_84),
		.c(new_net_83)
	);

	bfr new_net_2677_bfr_before (
		.din(new_net_2677),
		.dout(N10574)
	);

	bfr new_net_2678_bfr_before (
		.din(new_net_2678),
		.dout(new_net_2677)
	);

	bfr new_net_2679_bfr_before (
		.din(new_net_2679),
		.dout(new_net_2678)
	);

	bfr new_net_2680_bfr_before (
		.din(new_net_2680),
		.dout(new_net_2679)
	);

	bfr new_net_2681_bfr_before (
		.din(new_net_2681),
		.dout(new_net_2680)
	);

	bfr new_net_2682_bfr_before (
		.din(new_net_2682),
		.dout(new_net_2681)
	);

	bfr new_net_2683_bfr_before (
		.din(new_net_2683),
		.dout(new_net_2682)
	);

	bfr new_net_2684_bfr_before (
		.din(new_net_2684),
		.dout(new_net_2683)
	);

	bfr new_net_2685_bfr_before (
		.din(new_net_2685),
		.dout(new_net_2684)
	);

	bfr new_net_2686_bfr_before (
		.din(new_net_2686),
		.dout(new_net_2685)
	);

	bfr new_net_2687_bfr_before (
		.din(new_net_2687),
		.dout(new_net_2686)
	);

	bfr new_net_2688_bfr_before (
		.din(new_net_2688),
		.dout(new_net_2687)
	);

	bfr new_net_2689_bfr_before (
		.din(new_net_2689),
		.dout(new_net_2688)
	);

	bfr new_net_2690_bfr_before (
		.din(new_net_2690),
		.dout(new_net_2689)
	);

	bfr new_net_2691_bfr_before (
		.din(new_net_2691),
		.dout(new_net_2690)
	);

	bfr new_net_2692_bfr_before (
		.din(new_net_2692),
		.dout(new_net_2691)
	);

	bfr new_net_2693_bfr_before (
		.din(new_net_2693),
		.dout(new_net_2692)
	);

	bfr new_net_2694_bfr_before (
		.din(new_net_2694),
		.dout(new_net_2693)
	);

	bfr new_net_2695_bfr_before (
		.din(new_net_2695),
		.dout(new_net_2694)
	);

	bfr new_net_2696_bfr_before (
		.din(new_net_2696),
		.dout(new_net_2695)
	);

	bfr new_net_2697_bfr_before (
		.din(new_net_2697),
		.dout(new_net_2696)
	);

	bfr new_net_2698_bfr_before (
		.din(new_net_2698),
		.dout(new_net_2697)
	);

	bfr new_net_2699_bfr_before (
		.din(new_net_2699),
		.dout(new_net_2698)
	);

	bfr new_net_2700_bfr_before (
		.din(new_net_2700),
		.dout(new_net_2699)
	);

	bfr new_net_2701_bfr_before (
		.din(new_net_2701),
		.dout(new_net_2700)
	);

	bfr new_net_2702_bfr_before (
		.din(new_net_2702),
		.dout(new_net_2701)
	);

	bfr new_net_2703_bfr_before (
		.din(new_net_2703),
		.dout(new_net_2702)
	);

	bfr new_net_2704_bfr_before (
		.din(new_net_2704),
		.dout(new_net_2703)
	);

	bfr new_net_2705_bfr_before (
		.din(new_net_2705),
		.dout(new_net_2704)
	);

	bfr new_net_2706_bfr_before (
		.din(new_net_2706),
		.dout(new_net_2705)
	);

	bfr new_net_2707_bfr_before (
		.din(new_net_2707),
		.dout(new_net_2706)
	);

	bfr new_net_2708_bfr_before (
		.din(new_net_2708),
		.dout(new_net_2707)
	);

	bfr new_net_2709_bfr_before (
		.din(new_net_2709),
		.dout(new_net_2708)
	);

	bfr new_net_2710_bfr_before (
		.din(new_net_2710),
		.dout(new_net_2709)
	);

	bfr new_net_2711_bfr_before (
		.din(new_net_2711),
		.dout(new_net_2710)
	);

	bfr new_net_2712_bfr_before (
		.din(new_net_2712),
		.dout(new_net_2711)
	);

	bfr new_net_2713_bfr_before (
		.din(new_net_2713),
		.dout(new_net_2712)
	);

	bfr new_net_2714_bfr_before (
		.din(new_net_2714),
		.dout(new_net_2713)
	);

	bfr new_net_2715_bfr_before (
		.din(new_net_2715),
		.dout(new_net_2714)
	);

	bfr new_net_2716_bfr_before (
		.din(new_net_2716),
		.dout(new_net_2715)
	);

	bfr new_net_2717_bfr_before (
		.din(new_net_2717),
		.dout(new_net_2716)
	);

	bfr new_net_2718_bfr_before (
		.din(new_net_2718),
		.dout(new_net_2717)
	);

	bfr new_net_2719_bfr_before (
		.din(new_net_2719),
		.dout(new_net_2718)
	);

	bfr new_net_2720_bfr_before (
		.din(new_net_2720),
		.dout(new_net_2719)
	);

	spl2 new_net_4_v_fanout (
		.a(new_net_4),
		.b(new_net_463),
		.c(new_net_2720)
	);

	spl2 n_1361__v_fanout (
		.a(n_1361_),
		.b(new_net_292),
		.c(new_net_291)
	);

	bfr new_net_2721_bfr_before (
		.din(new_net_2721),
		.dout(N10576)
	);

	bfr new_net_2722_bfr_before (
		.din(new_net_2722),
		.dout(new_net_2721)
	);

	bfr new_net_2723_bfr_before (
		.din(new_net_2723),
		.dout(new_net_2722)
	);

	bfr new_net_2724_bfr_before (
		.din(new_net_2724),
		.dout(new_net_2723)
	);

	bfr new_net_2725_bfr_before (
		.din(new_net_2725),
		.dout(new_net_2724)
	);

	bfr new_net_2726_bfr_before (
		.din(new_net_2726),
		.dout(new_net_2725)
	);

	bfr new_net_2727_bfr_before (
		.din(new_net_2727),
		.dout(new_net_2726)
	);

	bfr new_net_2728_bfr_before (
		.din(new_net_2728),
		.dout(new_net_2727)
	);

	bfr new_net_2729_bfr_before (
		.din(new_net_2729),
		.dout(new_net_2728)
	);

	bfr new_net_2730_bfr_before (
		.din(new_net_2730),
		.dout(new_net_2729)
	);

	bfr new_net_2731_bfr_before (
		.din(new_net_2731),
		.dout(new_net_2730)
	);

	bfr new_net_2732_bfr_before (
		.din(new_net_2732),
		.dout(new_net_2731)
	);

	bfr new_net_2733_bfr_before (
		.din(new_net_2733),
		.dout(new_net_2732)
	);

	bfr new_net_2734_bfr_before (
		.din(new_net_2734),
		.dout(new_net_2733)
	);

	bfr new_net_2735_bfr_before (
		.din(new_net_2735),
		.dout(new_net_2734)
	);

	bfr new_net_2736_bfr_before (
		.din(new_net_2736),
		.dout(new_net_2735)
	);

	bfr new_net_2737_bfr_before (
		.din(new_net_2737),
		.dout(new_net_2736)
	);

	bfr new_net_2738_bfr_before (
		.din(new_net_2738),
		.dout(new_net_2737)
	);

	bfr new_net_2739_bfr_before (
		.din(new_net_2739),
		.dout(new_net_2738)
	);

	bfr new_net_2740_bfr_before (
		.din(new_net_2740),
		.dout(new_net_2739)
	);

	bfr new_net_2741_bfr_before (
		.din(new_net_2741),
		.dout(new_net_2740)
	);

	bfr new_net_2742_bfr_before (
		.din(new_net_2742),
		.dout(new_net_2741)
	);

	bfr new_net_2743_bfr_before (
		.din(new_net_2743),
		.dout(new_net_2742)
	);

	bfr new_net_2744_bfr_before (
		.din(new_net_2744),
		.dout(new_net_2743)
	);

	bfr new_net_2745_bfr_before (
		.din(new_net_2745),
		.dout(new_net_2744)
	);

	bfr new_net_2746_bfr_before (
		.din(new_net_2746),
		.dout(new_net_2745)
	);

	bfr new_net_2747_bfr_before (
		.din(new_net_2747),
		.dout(new_net_2746)
	);

	bfr new_net_2748_bfr_before (
		.din(new_net_2748),
		.dout(new_net_2747)
	);

	bfr new_net_2749_bfr_before (
		.din(new_net_2749),
		.dout(new_net_2748)
	);

	bfr new_net_2750_bfr_before (
		.din(new_net_2750),
		.dout(new_net_2749)
	);

	bfr new_net_2751_bfr_before (
		.din(new_net_2751),
		.dout(new_net_2750)
	);

	bfr new_net_2752_bfr_before (
		.din(new_net_2752),
		.dout(new_net_2751)
	);

	bfr new_net_2753_bfr_before (
		.din(new_net_2753),
		.dout(new_net_2752)
	);

	bfr new_net_2754_bfr_before (
		.din(new_net_2754),
		.dout(new_net_2753)
	);

	bfr new_net_2755_bfr_before (
		.din(new_net_2755),
		.dout(new_net_2754)
	);

	bfr new_net_2756_bfr_before (
		.din(new_net_2756),
		.dout(new_net_2755)
	);

	bfr new_net_2757_bfr_before (
		.din(new_net_2757),
		.dout(new_net_2756)
	);

	bfr new_net_2758_bfr_before (
		.din(new_net_2758),
		.dout(new_net_2757)
	);

	bfr new_net_2759_bfr_before (
		.din(new_net_2759),
		.dout(new_net_2758)
	);

	bfr new_net_2760_bfr_before (
		.din(new_net_2760),
		.dout(new_net_2759)
	);

	bfr new_net_2761_bfr_before (
		.din(new_net_2761),
		.dout(new_net_2760)
	);

	bfr new_net_2762_bfr_before (
		.din(new_net_2762),
		.dout(new_net_2761)
	);

	bfr new_net_2763_bfr_before (
		.din(new_net_2763),
		.dout(new_net_2762)
	);

	bfr new_net_2764_bfr_before (
		.din(new_net_2764),
		.dout(new_net_2763)
	);

	spl2 new_net_5_v_fanout (
		.a(new_net_5),
		.b(new_net_631),
		.c(new_net_2764)
	);

	bfr new_net_2765_bfr_after (
		.din(new_net_6),
		.dout(new_net_2765)
	);

	bfr new_net_2766_bfr_before (
		.din(new_net_2766),
		.dout(N10575)
	);

	bfr new_net_2767_bfr_before (
		.din(new_net_2767),
		.dout(new_net_2766)
	);

	bfr new_net_2768_bfr_before (
		.din(new_net_2768),
		.dout(new_net_2767)
	);

	bfr new_net_2769_bfr_before (
		.din(new_net_2769),
		.dout(new_net_2768)
	);

	bfr new_net_2770_bfr_before (
		.din(new_net_2770),
		.dout(new_net_2769)
	);

	bfr new_net_2771_bfr_before (
		.din(new_net_2771),
		.dout(new_net_2770)
	);

	bfr new_net_2772_bfr_before (
		.din(new_net_2772),
		.dout(new_net_2771)
	);

	bfr new_net_2773_bfr_before (
		.din(new_net_2773),
		.dout(new_net_2772)
	);

	bfr new_net_2774_bfr_before (
		.din(new_net_2774),
		.dout(new_net_2773)
	);

	bfr new_net_2775_bfr_before (
		.din(new_net_2775),
		.dout(new_net_2774)
	);

	bfr new_net_2776_bfr_before (
		.din(new_net_2776),
		.dout(new_net_2775)
	);

	bfr new_net_2777_bfr_before (
		.din(new_net_2777),
		.dout(new_net_2776)
	);

	bfr new_net_2778_bfr_before (
		.din(new_net_2778),
		.dout(new_net_2777)
	);

	bfr new_net_2779_bfr_before (
		.din(new_net_2779),
		.dout(new_net_2778)
	);

	bfr new_net_2780_bfr_before (
		.din(new_net_2780),
		.dout(new_net_2779)
	);

	bfr new_net_2781_bfr_before (
		.din(new_net_2781),
		.dout(new_net_2780)
	);

	bfr new_net_2782_bfr_before (
		.din(new_net_2782),
		.dout(new_net_2781)
	);

	bfr new_net_2783_bfr_before (
		.din(new_net_2783),
		.dout(new_net_2782)
	);

	bfr new_net_2784_bfr_before (
		.din(new_net_2784),
		.dout(new_net_2783)
	);

	bfr new_net_2785_bfr_before (
		.din(new_net_2785),
		.dout(new_net_2784)
	);

	bfr new_net_2786_bfr_before (
		.din(new_net_2786),
		.dout(new_net_2785)
	);

	bfr new_net_2787_bfr_before (
		.din(new_net_2787),
		.dout(new_net_2786)
	);

	bfr new_net_2788_bfr_before (
		.din(new_net_2788),
		.dout(new_net_2787)
	);

	bfr new_net_2789_bfr_before (
		.din(new_net_2789),
		.dout(new_net_2788)
	);

	bfr new_net_2790_bfr_before (
		.din(new_net_2790),
		.dout(new_net_2789)
	);

	bfr new_net_2791_bfr_before (
		.din(new_net_2791),
		.dout(new_net_2790)
	);

	bfr new_net_2792_bfr_before (
		.din(new_net_2792),
		.dout(new_net_2791)
	);

	bfr new_net_2793_bfr_before (
		.din(new_net_2793),
		.dout(new_net_2792)
	);

	bfr new_net_2794_bfr_before (
		.din(new_net_2794),
		.dout(new_net_2793)
	);

	bfr new_net_2795_bfr_before (
		.din(new_net_2795),
		.dout(new_net_2794)
	);

	bfr new_net_2796_bfr_before (
		.din(new_net_2796),
		.dout(new_net_2795)
	);

	bfr new_net_2797_bfr_before (
		.din(new_net_2797),
		.dout(new_net_2796)
	);

	bfr new_net_2798_bfr_before (
		.din(new_net_2798),
		.dout(new_net_2797)
	);

	bfr new_net_2799_bfr_before (
		.din(new_net_2799),
		.dout(new_net_2798)
	);

	bfr new_net_2800_bfr_before (
		.din(new_net_2800),
		.dout(new_net_2799)
	);

	bfr new_net_2801_bfr_before (
		.din(new_net_2801),
		.dout(new_net_2800)
	);

	bfr new_net_2802_bfr_before (
		.din(new_net_2802),
		.dout(new_net_2801)
	);

	bfr new_net_2803_bfr_before (
		.din(new_net_2803),
		.dout(new_net_2802)
	);

	bfr new_net_2804_bfr_before (
		.din(new_net_2804),
		.dout(new_net_2803)
	);

	bfr new_net_2805_bfr_before (
		.din(new_net_2805),
		.dout(new_net_2804)
	);

	bfr new_net_2806_bfr_before (
		.din(new_net_2806),
		.dout(new_net_2805)
	);

	bfr new_net_2807_bfr_before (
		.din(new_net_2807),
		.dout(new_net_2806)
	);

	bfr new_net_2808_bfr_before (
		.din(new_net_2808),
		.dout(new_net_2807)
	);

	bfr new_net_2809_bfr_before (
		.din(new_net_2809),
		.dout(new_net_2808)
	);

	spl2 new_net_6_v_fanout (
		.a(new_net_2765),
		.b(new_net_724),
		.c(new_net_2809)
	);

	bfr new_net_2810_bfr_before (
		.din(new_net_2810),
		.dout(new_net_1216)
	);

	bfr new_net_2811_bfr_before (
		.din(new_net_2811),
		.dout(new_net_2810)
	);

	bfr new_net_2812_bfr_before (
		.din(new_net_2812),
		.dout(new_net_2811)
	);

	bfr new_net_2813_bfr_before (
		.din(new_net_2813),
		.dout(new_net_2812)
	);

	bfr new_net_2814_bfr_before (
		.din(new_net_2814),
		.dout(new_net_2813)
	);

	bfr new_net_2815_bfr_before (
		.din(new_net_2815),
		.dout(new_net_2814)
	);

	bfr new_net_2816_bfr_before (
		.din(new_net_2816),
		.dout(new_net_2815)
	);

	bfr new_net_2817_bfr_before (
		.din(new_net_2817),
		.dout(new_net_2816)
	);

	bfr new_net_2818_bfr_before (
		.din(new_net_2818),
		.dout(new_net_2817)
	);

	bfr new_net_2819_bfr_before (
		.din(new_net_2819),
		.dout(new_net_2818)
	);

	bfr new_net_2820_bfr_before (
		.din(new_net_2820),
		.dout(new_net_2819)
	);

	bfr new_net_2821_bfr_before (
		.din(new_net_2821),
		.dout(new_net_2820)
	);

	bfr new_net_2822_bfr_before (
		.din(new_net_2822),
		.dout(new_net_2821)
	);

	bfr new_net_2823_bfr_before (
		.din(new_net_2823),
		.dout(new_net_2822)
	);

	bfr new_net_2824_bfr_before (
		.din(new_net_2824),
		.dout(new_net_2823)
	);

	bfr new_net_2825_bfr_before (
		.din(new_net_2825),
		.dout(new_net_2824)
	);

	bfr new_net_2826_bfr_before (
		.din(new_net_2826),
		.dout(new_net_2825)
	);

	bfr new_net_2827_bfr_before (
		.din(new_net_2827),
		.dout(new_net_2826)
	);

	bfr new_net_2828_bfr_before (
		.din(new_net_2828),
		.dout(new_net_2827)
	);

	bfr new_net_2829_bfr_before (
		.din(new_net_2829),
		.dout(new_net_2828)
	);

	bfr new_net_2830_bfr_before (
		.din(new_net_2830),
		.dout(new_net_2829)
	);

	bfr new_net_2831_bfr_before (
		.din(new_net_2831),
		.dout(new_net_2830)
	);

	bfr new_net_2832_bfr_before (
		.din(new_net_2832),
		.dout(new_net_2831)
	);

	bfr new_net_2833_bfr_before (
		.din(new_net_2833),
		.dout(new_net_2832)
	);

	bfr new_net_2834_bfr_before (
		.din(new_net_2834),
		.dout(new_net_2833)
	);

	spl4L n_0059__v_fanout (
		.a(n_0059_),
		.b(new_net_1215),
		.c(new_net_2834),
		.d(new_net_1214),
		.e(new_net_1213)
	);

	spl2 new_net_2172_v_fanout (
		.a(new_net_2172),
		.b(new_net_687),
		.c(new_net_688)
	);

	spl2 new_net_2165_v_fanout (
		.a(new_net_2165),
		.b(new_net_1737),
		.c(new_net_1736)
	);

	bfr new_net_2835_bfr_after (
		.din(n_0636_),
		.dout(new_net_2835)
	);

	bfr new_net_2836_bfr_after (
		.din(new_net_2835),
		.dout(new_net_2836)
	);

	bfr new_net_2837_bfr_after (
		.din(new_net_2836),
		.dout(new_net_2837)
	);

	spl2 n_0636__v_fanout (
		.a(new_net_2837),
		.b(new_net_1254),
		.c(new_net_1253)
	);

	spl2 n_0585__v_fanout (
		.a(n_0585_),
		.b(new_net_1695),
		.c(new_net_1694)
	);

	spl3L n_0012__v_fanout (
		.a(n_0012_),
		.b(new_net_51),
		.c(new_net_49),
		.d(new_net_50)
	);

	bfr new_net_2838_bfr_after (
		.din(n_0424_),
		.dout(new_net_2838)
	);

	bfr new_net_2839_bfr_after (
		.din(new_net_2838),
		.dout(new_net_2839)
	);

	bfr new_net_2840_bfr_after (
		.din(new_net_2839),
		.dout(new_net_2840)
	);

	spl2 n_0424__v_fanout (
		.a(new_net_2840),
		.b(new_net_394),
		.c(new_net_393)
	);

	bfr new_net_2841_bfr_after (
		.din(n_0506_),
		.dout(new_net_2841)
	);

	bfr new_net_2842_bfr_after (
		.din(new_net_2841),
		.dout(new_net_2842)
	);

	bfr new_net_2843_bfr_after (
		.din(new_net_2842),
		.dout(new_net_2843)
	);

	spl2 n_0506__v_fanout (
		.a(new_net_2843),
		.b(new_net_923),
		.c(new_net_922)
	);

	spl2 new_net_2141_v_fanout (
		.a(new_net_2141),
		.b(new_net_106),
		.c(new_net_104)
	);

	bfr new_net_2844_bfr_before (
		.din(new_net_2844),
		.dout(new_net_533)
	);

	bfr new_net_2845_bfr_before (
		.din(new_net_2845),
		.dout(new_net_2844)
	);

	bfr new_net_2846_bfr_before (
		.din(new_net_2846),
		.dout(new_net_2845)
	);

	bfr new_net_2847_bfr_before (
		.din(new_net_2847),
		.dout(new_net_2846)
	);

	bfr new_net_2848_bfr_before (
		.din(new_net_2848),
		.dout(new_net_2847)
	);

	bfr new_net_2849_bfr_before (
		.din(new_net_2849),
		.dout(new_net_2848)
	);

	bfr new_net_2850_bfr_before (
		.din(new_net_2850),
		.dout(new_net_2849)
	);

	bfr new_net_2851_bfr_before (
		.din(new_net_2851),
		.dout(new_net_2850)
	);

	bfr new_net_2852_bfr_before (
		.din(new_net_2852),
		.dout(new_net_2851)
	);

	bfr new_net_2853_bfr_before (
		.din(new_net_2853),
		.dout(new_net_2852)
	);

	bfr new_net_2854_bfr_before (
		.din(new_net_2854),
		.dout(new_net_2853)
	);

	bfr new_net_2855_bfr_before (
		.din(new_net_2855),
		.dout(new_net_2854)
	);

	bfr new_net_2856_bfr_before (
		.din(new_net_2856),
		.dout(new_net_2855)
	);

	bfr new_net_2857_bfr_before (
		.din(new_net_2857),
		.dout(new_net_2856)
	);

	bfr new_net_2858_bfr_before (
		.din(new_net_2858),
		.dout(new_net_2857)
	);

	bfr new_net_2859_bfr_before (
		.din(new_net_2859),
		.dout(new_net_2858)
	);

	bfr new_net_2860_bfr_before (
		.din(new_net_2860),
		.dout(new_net_2859)
	);

	bfr new_net_2861_bfr_before (
		.din(new_net_2861),
		.dout(new_net_2860)
	);

	bfr new_net_2862_bfr_before (
		.din(new_net_2862),
		.dout(new_net_2861)
	);

	bfr new_net_2863_bfr_before (
		.din(new_net_2863),
		.dout(new_net_2862)
	);

	bfr new_net_2864_bfr_before (
		.din(new_net_2864),
		.dout(new_net_2863)
	);

	bfr new_net_2865_bfr_before (
		.din(new_net_2865),
		.dout(new_net_2864)
	);

	bfr new_net_2866_bfr_before (
		.din(new_net_2866),
		.dout(new_net_2865)
	);

	bfr new_net_2867_bfr_before (
		.din(new_net_2867),
		.dout(new_net_2866)
	);

	bfr new_net_2868_bfr_before (
		.din(new_net_2868),
		.dout(new_net_2867)
	);

	bfr new_net_2869_bfr_before (
		.din(new_net_2869),
		.dout(new_net_2868)
	);

	bfr new_net_2870_bfr_before (
		.din(new_net_2870),
		.dout(new_net_2869)
	);

	bfr new_net_2871_bfr_before (
		.din(new_net_2871),
		.dout(new_net_2870)
	);

	bfr new_net_2872_bfr_before (
		.din(new_net_2872),
		.dout(new_net_2871)
	);

	bfr new_net_2873_bfr_before (
		.din(new_net_2873),
		.dout(new_net_2872)
	);

	bfr new_net_2874_bfr_before (
		.din(new_net_2874),
		.dout(new_net_2873)
	);

	bfr new_net_2875_bfr_before (
		.din(new_net_2875),
		.dout(new_net_2874)
	);

	bfr new_net_2876_bfr_before (
		.din(new_net_2876),
		.dout(new_net_2875)
	);

	bfr new_net_2877_bfr_before (
		.din(new_net_2877),
		.dout(new_net_2876)
	);

	bfr new_net_2878_bfr_before (
		.din(new_net_2878),
		.dout(new_net_2877)
	);

	bfr new_net_2879_bfr_before (
		.din(new_net_2879),
		.dout(new_net_2878)
	);

	spl3L n_0110__v_fanout (
		.a(n_0110_),
		.b(new_net_535),
		.c(new_net_2879),
		.d(new_net_534)
	);

	spl2 new_net_2152_v_fanout (
		.a(new_net_2152),
		.b(new_net_1423),
		.c(new_net_1424)
	);

	bfr new_net_2880_bfr_after (
		.din(n_0554_),
		.dout(new_net_2880)
	);

	bfr new_net_2881_bfr_after (
		.din(new_net_2880),
		.dout(new_net_2881)
	);

	bfr new_net_2882_bfr_after (
		.din(new_net_2881),
		.dout(new_net_2882)
	);

	spl2 n_0554__v_fanout (
		.a(new_net_2882),
		.b(new_net_1946),
		.c(new_net_1945)
	);

	spl3L n_1364__v_fanout (
		.a(n_1364_),
		.b(new_net_681),
		.c(new_net_679),
		.d(new_net_680)
	);

	spl2 n_0703__v_fanout (
		.a(n_0703_),
		.b(new_net_1537),
		.c(new_net_1536)
	);

	bfr new_net_2883_bfr_before (
		.din(new_net_2883),
		.dout(new_net_1876)
	);

	bfr new_net_2884_bfr_before (
		.din(new_net_2884),
		.dout(new_net_2883)
	);

	spl2 new_net_2106_v_fanout (
		.a(new_net_2106),
		.b(new_net_2884),
		.c(new_net_1875)
	);

	spl2 n_0541__v_fanout (
		.a(n_0541_),
		.b(new_net_1658),
		.c(new_net_1657)
	);

	bfr new_net_2885_bfr_before (
		.din(new_net_2885),
		.dout(new_net_873)
	);

	bfr new_net_2886_bfr_before (
		.din(new_net_2886),
		.dout(new_net_2885)
	);

	bfr new_net_2887_bfr_before (
		.din(new_net_2887),
		.dout(new_net_2886)
	);

	bfr new_net_2888_bfr_before (
		.din(new_net_2888),
		.dout(new_net_2887)
	);

	bfr new_net_2889_bfr_before (
		.din(new_net_2889),
		.dout(new_net_2888)
	);

	bfr new_net_2890_bfr_before (
		.din(new_net_2890),
		.dout(new_net_2889)
	);

	bfr new_net_2891_bfr_before (
		.din(new_net_2891),
		.dout(new_net_2890)
	);

	bfr new_net_2892_bfr_before (
		.din(new_net_2892),
		.dout(new_net_2891)
	);

	bfr new_net_2893_bfr_before (
		.din(new_net_2893),
		.dout(new_net_2892)
	);

	bfr new_net_2894_bfr_before (
		.din(new_net_2894),
		.dout(new_net_2893)
	);

	bfr new_net_2895_bfr_before (
		.din(new_net_2895),
		.dout(new_net_2894)
	);

	bfr new_net_2896_bfr_before (
		.din(new_net_2896),
		.dout(new_net_2895)
	);

	bfr new_net_2897_bfr_before (
		.din(new_net_2897),
		.dout(new_net_2896)
	);

	bfr new_net_2898_bfr_before (
		.din(new_net_2898),
		.dout(new_net_2897)
	);

	bfr new_net_2899_bfr_before (
		.din(new_net_2899),
		.dout(new_net_2898)
	);

	bfr new_net_2900_bfr_before (
		.din(new_net_2900),
		.dout(new_net_2899)
	);

	bfr new_net_2901_bfr_before (
		.din(new_net_2901),
		.dout(new_net_2900)
	);

	bfr new_net_2902_bfr_before (
		.din(new_net_2902),
		.dout(new_net_2901)
	);

	bfr new_net_2903_bfr_before (
		.din(new_net_2903),
		.dout(new_net_2902)
	);

	bfr new_net_2904_bfr_before (
		.din(new_net_2904),
		.dout(new_net_2903)
	);

	bfr new_net_2905_bfr_before (
		.din(new_net_2905),
		.dout(new_net_2904)
	);

	bfr new_net_2906_bfr_before (
		.din(new_net_2906),
		.dout(new_net_2905)
	);

	bfr new_net_2907_bfr_before (
		.din(new_net_2907),
		.dout(new_net_2906)
	);

	bfr new_net_2908_bfr_before (
		.din(new_net_2908),
		.dout(new_net_2907)
	);

	bfr new_net_2909_bfr_before (
		.din(new_net_2909),
		.dout(new_net_2908)
	);

	bfr new_net_2910_bfr_before (
		.din(new_net_2910),
		.dout(new_net_2909)
	);

	bfr new_net_2911_bfr_before (
		.din(new_net_2911),
		.dout(new_net_2910)
	);

	bfr new_net_2912_bfr_before (
		.din(new_net_2912),
		.dout(new_net_2911)
	);

	spl3L n_0043__v_fanout (
		.a(n_0043_),
		.b(new_net_874),
		.c(new_net_2912),
		.d(new_net_875)
	);

	spl2 new_net_2146_v_fanout (
		.a(new_net_2146),
		.b(new_net_1074),
		.c(new_net_1075)
	);

	spl2 n_0535__v_fanout (
		.a(n_0535_),
		.b(new_net_1541),
		.c(new_net_1540)
	);

	spl2 n_0403__v_fanout (
		.a(n_0403_),
		.b(new_net_1761),
		.c(new_net_1760)
	);

	spl2 n_0485__v_fanout (
		.a(n_0485_),
		.b(new_net_440),
		.c(new_net_439)
	);

	spl2 n_0706__v_fanout (
		.a(n_0706_),
		.b(new_net_953),
		.c(new_net_952)
	);

	spl2 n_0561__v_fanout (
		.a(n_0561_),
		.b(new_net_1208),
		.c(new_net_1207)
	);

	bfr new_net_2913_bfr_after (
		.din(n_1340_),
		.dout(new_net_2913)
	);

	bfr new_net_2914_bfr_after (
		.din(new_net_2913),
		.dout(new_net_2914)
	);

	bfr new_net_2915_bfr_after (
		.din(new_net_2914),
		.dout(new_net_2915)
	);

	bfr new_net_2916_bfr_after (
		.din(new_net_2915),
		.dout(new_net_2916)
	);

	bfr new_net_2917_bfr_after (
		.din(new_net_2916),
		.dout(new_net_2917)
	);

	bfr new_net_2918_bfr_after (
		.din(new_net_2917),
		.dout(new_net_2918)
	);

	bfr new_net_2919_bfr_before (
		.din(new_net_2919),
		.dout(new_net_1534)
	);

	bfr new_net_2920_bfr_before (
		.din(new_net_2920),
		.dout(new_net_2919)
	);

	bfr new_net_2921_bfr_before (
		.din(new_net_2921),
		.dout(new_net_2920)
	);

	bfr new_net_2922_bfr_before (
		.din(new_net_2922),
		.dout(new_net_2921)
	);

	bfr new_net_2923_bfr_before (
		.din(new_net_2923),
		.dout(new_net_2922)
	);

	bfr new_net_2924_bfr_before (
		.din(new_net_2924),
		.dout(new_net_2923)
	);

	spl2 n_1340__v_fanout (
		.a(new_net_2918),
		.b(new_net_1535),
		.c(new_net_2924)
	);

	bfr new_net_2925_bfr_after (
		.din(n_0615_),
		.dout(new_net_2925)
	);

	bfr new_net_2926_bfr_after (
		.din(new_net_2925),
		.dout(new_net_2926)
	);

	bfr new_net_2927_bfr_after (
		.din(new_net_2926),
		.dout(new_net_2927)
	);

	spl2 n_0615__v_fanout (
		.a(new_net_2927),
		.b(new_net_548),
		.c(new_net_547)
	);

	bfr new_net_2928_bfr_after (
		.din(n_0459_),
		.dout(new_net_2928)
	);

	spl2 n_0459__v_fanout (
		.a(new_net_2928),
		.b(new_net_1595),
		.c(new_net_1594)
	);

	bfr new_net_2929_bfr_before (
		.din(new_net_2929),
		.dout(new_net_1217)
	);

	bfr new_net_2930_bfr_before (
		.din(new_net_2930),
		.dout(new_net_2929)
	);

	bfr new_net_2931_bfr_before (
		.din(new_net_2931),
		.dout(new_net_2930)
	);

	bfr new_net_2932_bfr_before (
		.din(new_net_2932),
		.dout(new_net_2931)
	);

	bfr new_net_2933_bfr_before (
		.din(new_net_2933),
		.dout(new_net_2932)
	);

	bfr new_net_2934_bfr_before (
		.din(new_net_2934),
		.dout(new_net_2933)
	);

	bfr new_net_2935_bfr_before (
		.din(new_net_2935),
		.dout(new_net_2934)
	);

	bfr new_net_2936_bfr_before (
		.din(new_net_2936),
		.dout(new_net_2935)
	);

	bfr new_net_2937_bfr_before (
		.din(new_net_2937),
		.dout(new_net_2936)
	);

	bfr new_net_2938_bfr_before (
		.din(new_net_2938),
		.dout(new_net_2937)
	);

	bfr new_net_2939_bfr_before (
		.din(new_net_2939),
		.dout(new_net_2938)
	);

	bfr new_net_2940_bfr_before (
		.din(new_net_2940),
		.dout(new_net_2939)
	);

	bfr new_net_2941_bfr_before (
		.din(new_net_2941),
		.dout(new_net_2940)
	);

	bfr new_net_2942_bfr_before (
		.din(new_net_2942),
		.dout(new_net_2941)
	);

	bfr new_net_2943_bfr_before (
		.din(new_net_2943),
		.dout(new_net_2942)
	);

	bfr new_net_2944_bfr_before (
		.din(new_net_2944),
		.dout(new_net_2943)
	);

	bfr new_net_2945_bfr_before (
		.din(new_net_2945),
		.dout(new_net_2944)
	);

	bfr new_net_2946_bfr_before (
		.din(new_net_2946),
		.dout(new_net_2945)
	);

	spl3L n_1319__v_fanout (
		.a(n_1319_),
		.b(new_net_1219),
		.c(new_net_2946),
		.d(new_net_1218)
	);

	bfr new_net_2947_bfr_before (
		.din(new_net_2947),
		.dout(new_net_2172)
	);

	spl3L n_0621__v_fanout (
		.a(n_0621_),
		.b(new_net_2947),
		.c(new_net_686),
		.d(new_net_689)
	);

	spl2 n_1359__v_fanout (
		.a(n_1359_),
		.b(new_net_1936),
		.c(new_net_1935)
	);

	bfr new_net_2948_bfr_before (
		.din(new_net_2948),
		.dout(new_net_1511)
	);

	bfr new_net_2949_bfr_before (
		.din(new_net_2949),
		.dout(new_net_2948)
	);

	bfr new_net_2950_bfr_before (
		.din(new_net_2950),
		.dout(new_net_2949)
	);

	bfr new_net_2951_bfr_before (
		.din(new_net_2951),
		.dout(new_net_2950)
	);

	bfr new_net_2952_bfr_before (
		.din(new_net_2952),
		.dout(new_net_2951)
	);

	bfr new_net_2953_bfr_before (
		.din(new_net_2953),
		.dout(new_net_2952)
	);

	bfr new_net_2954_bfr_before (
		.din(new_net_2954),
		.dout(new_net_2953)
	);

	bfr new_net_2955_bfr_before (
		.din(new_net_2955),
		.dout(new_net_2954)
	);

	bfr new_net_2956_bfr_before (
		.din(new_net_2956),
		.dout(new_net_2955)
	);

	spl2 new_net_2171_v_fanout (
		.a(new_net_2171),
		.b(new_net_2956),
		.c(new_net_1514)
	);

	bfr new_net_2957_bfr_after (
		.din(n_0590_),
		.dout(new_net_2957)
	);

	bfr new_net_2958_bfr_after (
		.din(new_net_2957),
		.dout(new_net_2958)
	);

	spl2 n_0590__v_fanout (
		.a(new_net_2958),
		.b(new_net_1792),
		.c(new_net_1791)
	);

	bfr new_net_2959_bfr_before (
		.din(new_net_2959),
		.dout(new_net_482)
	);

	bfr new_net_2960_bfr_before (
		.din(new_net_2960),
		.dout(new_net_2959)
	);

	bfr new_net_2961_bfr_before (
		.din(new_net_2961),
		.dout(new_net_2960)
	);

	bfr new_net_2962_bfr_before (
		.din(new_net_2962),
		.dout(new_net_2961)
	);

	bfr new_net_2963_bfr_before (
		.din(new_net_2963),
		.dout(new_net_2962)
	);

	bfr new_net_2964_bfr_before (
		.din(new_net_2964),
		.dout(new_net_2963)
	);

	bfr new_net_2965_bfr_before (
		.din(new_net_2965),
		.dout(new_net_2964)
	);

	bfr new_net_2966_bfr_before (
		.din(new_net_2966),
		.dout(new_net_2965)
	);

	bfr new_net_2967_bfr_before (
		.din(new_net_2967),
		.dout(new_net_2966)
	);

	bfr new_net_2968_bfr_before (
		.din(new_net_2968),
		.dout(new_net_2967)
	);

	bfr new_net_2969_bfr_before (
		.din(new_net_2969),
		.dout(new_net_2968)
	);

	bfr new_net_2970_bfr_before (
		.din(new_net_2970),
		.dout(new_net_2969)
	);

	bfr new_net_2971_bfr_before (
		.din(new_net_2971),
		.dout(new_net_2970)
	);

	bfr new_net_2972_bfr_before (
		.din(new_net_2972),
		.dout(new_net_2971)
	);

	bfr new_net_2973_bfr_before (
		.din(new_net_2973),
		.dout(new_net_2972)
	);

	bfr new_net_2974_bfr_before (
		.din(new_net_2974),
		.dout(new_net_2973)
	);

	bfr new_net_2975_bfr_before (
		.din(new_net_2975),
		.dout(new_net_2974)
	);

	bfr new_net_2976_bfr_before (
		.din(new_net_2976),
		.dout(new_net_2975)
	);

	bfr new_net_2977_bfr_before (
		.din(new_net_2977),
		.dout(new_net_2976)
	);

	bfr new_net_2978_bfr_before (
		.din(new_net_2978),
		.dout(new_net_2977)
	);

	bfr new_net_2979_bfr_before (
		.din(new_net_2979),
		.dout(new_net_2978)
	);

	bfr new_net_2980_bfr_before (
		.din(new_net_2980),
		.dout(new_net_2979)
	);

	bfr new_net_2981_bfr_before (
		.din(new_net_2981),
		.dout(new_net_2980)
	);

	bfr new_net_2982_bfr_before (
		.din(new_net_2982),
		.dout(new_net_2981)
	);

	bfr new_net_2983_bfr_before (
		.din(new_net_2983),
		.dout(new_net_2982)
	);

	bfr new_net_2984_bfr_before (
		.din(new_net_2984),
		.dout(new_net_2983)
	);

	bfr new_net_2985_bfr_before (
		.din(new_net_2985),
		.dout(new_net_2984)
	);

	bfr new_net_2986_bfr_before (
		.din(new_net_2986),
		.dout(new_net_2985)
	);

	bfr new_net_2987_bfr_before (
		.din(new_net_2987),
		.dout(new_net_2986)
	);

	bfr new_net_2988_bfr_before (
		.din(new_net_2988),
		.dout(new_net_2987)
	);

	bfr new_net_2989_bfr_before (
		.din(new_net_2989),
		.dout(new_net_2988)
	);

	bfr new_net_2990_bfr_before (
		.din(new_net_2990),
		.dout(new_net_2989)
	);

	bfr new_net_2991_bfr_before (
		.din(new_net_2991),
		.dout(new_net_2990)
	);

	bfr new_net_2992_bfr_before (
		.din(new_net_2992),
		.dout(new_net_2991)
	);

	bfr new_net_2993_bfr_before (
		.din(new_net_2993),
		.dout(new_net_2992)
	);

	bfr new_net_2994_bfr_before (
		.din(new_net_2994),
		.dout(new_net_2993)
	);

	bfr new_net_2995_bfr_before (
		.din(new_net_2995),
		.dout(new_net_2994)
	);

	bfr new_net_2996_bfr_before (
		.din(new_net_2996),
		.dout(new_net_2995)
	);

	spl4L new_net_2168_v_fanout (
		.a(new_net_2168),
		.b(new_net_483),
		.c(new_net_479),
		.d(new_net_2996),
		.e(new_net_480)
	);

	spl4L new_net_2170_v_fanout (
		.a(new_net_2170),
		.b(new_net_1512),
		.c(new_net_1510),
		.d(new_net_2171),
		.e(new_net_1513)
	);

	bfr new_net_2997_bfr_after (
		.din(n_0526_),
		.dout(new_net_2997)
	);

	spl2 n_0526__v_fanout (
		.a(new_net_2997),
		.b(new_net_1833),
		.c(new_net_1832)
	);

	bfr new_net_2998_bfr_before (
		.din(new_net_2998),
		.dout(new_net_1451)
	);

	bfr new_net_2999_bfr_before (
		.din(new_net_2999),
		.dout(new_net_2998)
	);

	bfr new_net_3000_bfr_before (
		.din(new_net_3000),
		.dout(new_net_2999)
	);

	bfr new_net_3001_bfr_before (
		.din(new_net_3001),
		.dout(new_net_3000)
	);

	bfr new_net_3002_bfr_before (
		.din(new_net_3002),
		.dout(new_net_3001)
	);

	bfr new_net_3003_bfr_before (
		.din(new_net_3003),
		.dout(new_net_3002)
	);

	bfr new_net_3004_bfr_before (
		.din(new_net_3004),
		.dout(new_net_3003)
	);

	bfr new_net_3005_bfr_before (
		.din(new_net_3005),
		.dout(new_net_3004)
	);

	bfr new_net_3006_bfr_before (
		.din(new_net_3006),
		.dout(new_net_3005)
	);

	bfr new_net_3007_bfr_before (
		.din(new_net_3007),
		.dout(new_net_3006)
	);

	bfr new_net_3008_bfr_before (
		.din(new_net_3008),
		.dout(new_net_3007)
	);

	bfr new_net_3009_bfr_before (
		.din(new_net_3009),
		.dout(new_net_3008)
	);

	bfr new_net_3010_bfr_before (
		.din(new_net_3010),
		.dout(new_net_3009)
	);

	bfr new_net_3011_bfr_before (
		.din(new_net_3011),
		.dout(new_net_3010)
	);

	bfr new_net_3012_bfr_before (
		.din(new_net_3012),
		.dout(new_net_3011)
	);

	bfr new_net_3013_bfr_before (
		.din(new_net_3013),
		.dout(new_net_3012)
	);

	bfr new_net_3014_bfr_before (
		.din(new_net_3014),
		.dout(new_net_3013)
	);

	bfr new_net_3015_bfr_before (
		.din(new_net_3015),
		.dout(new_net_3014)
	);

	bfr new_net_3016_bfr_before (
		.din(new_net_3016),
		.dout(new_net_3015)
	);

	bfr new_net_3017_bfr_before (
		.din(new_net_3017),
		.dout(new_net_3016)
	);

	bfr new_net_3018_bfr_before (
		.din(new_net_3018),
		.dout(new_net_3017)
	);

	bfr new_net_3019_bfr_before (
		.din(new_net_3019),
		.dout(new_net_3018)
	);

	bfr new_net_3020_bfr_before (
		.din(new_net_3020),
		.dout(new_net_3019)
	);

	bfr new_net_3021_bfr_before (
		.din(new_net_3021),
		.dout(new_net_3020)
	);

	bfr new_net_3022_bfr_before (
		.din(new_net_3022),
		.dout(new_net_3021)
	);

	bfr new_net_3023_bfr_before (
		.din(new_net_3023),
		.dout(new_net_3022)
	);

	bfr new_net_3024_bfr_before (
		.din(new_net_3024),
		.dout(new_net_3023)
	);

	spl4L new_net_2166_v_fanout (
		.a(new_net_2166),
		.b(new_net_1448),
		.c(new_net_3024),
		.d(new_net_1450),
		.e(new_net_1449)
	);

	bfr new_net_3025_bfr_before (
		.din(new_net_3025),
		.dout(new_net_855)
	);

	bfr new_net_3026_bfr_before (
		.din(new_net_3026),
		.dout(new_net_3025)
	);

	bfr new_net_3027_bfr_before (
		.din(new_net_3027),
		.dout(new_net_3026)
	);

	bfr new_net_3028_bfr_before (
		.din(new_net_3028),
		.dout(new_net_3027)
	);

	bfr new_net_3029_bfr_before (
		.din(new_net_3029),
		.dout(new_net_3028)
	);

	bfr new_net_3030_bfr_before (
		.din(new_net_3030),
		.dout(new_net_3029)
	);

	bfr new_net_3031_bfr_before (
		.din(new_net_3031),
		.dout(new_net_3030)
	);

	bfr new_net_3032_bfr_before (
		.din(new_net_3032),
		.dout(new_net_3031)
	);

	bfr new_net_3033_bfr_before (
		.din(new_net_3033),
		.dout(new_net_3032)
	);

	bfr new_net_3034_bfr_before (
		.din(new_net_3034),
		.dout(new_net_3033)
	);

	bfr new_net_3035_bfr_before (
		.din(new_net_3035),
		.dout(new_net_3034)
	);

	bfr new_net_3036_bfr_before (
		.din(new_net_3036),
		.dout(new_net_3035)
	);

	bfr new_net_3037_bfr_before (
		.din(new_net_3037),
		.dout(new_net_3036)
	);

	bfr new_net_3038_bfr_before (
		.din(new_net_3038),
		.dout(new_net_3037)
	);

	bfr new_net_3039_bfr_before (
		.din(new_net_3039),
		.dout(new_net_3038)
	);

	bfr new_net_3040_bfr_before (
		.din(new_net_3040),
		.dout(new_net_3039)
	);

	bfr new_net_3041_bfr_before (
		.din(new_net_3041),
		.dout(new_net_3040)
	);

	bfr new_net_3042_bfr_before (
		.din(new_net_3042),
		.dout(new_net_3041)
	);

	bfr new_net_3043_bfr_before (
		.din(new_net_3043),
		.dout(new_net_3042)
	);

	bfr new_net_3044_bfr_before (
		.din(new_net_3044),
		.dout(new_net_3043)
	);

	bfr new_net_3045_bfr_before (
		.din(new_net_3045),
		.dout(new_net_3044)
	);

	bfr new_net_3046_bfr_before (
		.din(new_net_3046),
		.dout(new_net_3045)
	);

	bfr new_net_3047_bfr_before (
		.din(new_net_3047),
		.dout(new_net_3046)
	);

	bfr new_net_3048_bfr_before (
		.din(new_net_3048),
		.dout(new_net_3047)
	);

	bfr new_net_3049_bfr_before (
		.din(new_net_3049),
		.dout(new_net_3048)
	);

	bfr new_net_3050_bfr_before (
		.din(new_net_3050),
		.dout(new_net_3049)
	);

	bfr new_net_3051_bfr_before (
		.din(new_net_3051),
		.dout(new_net_3050)
	);

	bfr new_net_3052_bfr_before (
		.din(new_net_3052),
		.dout(new_net_3051)
	);

	bfr new_net_3053_bfr_before (
		.din(new_net_3053),
		.dout(new_net_3052)
	);

	spl2 n_0036__v_fanout (
		.a(n_0036_),
		.b(new_net_3053),
		.c(new_net_854)
	);

	spl2 n_0695__v_fanout (
		.a(n_0695_),
		.b(new_net_1353),
		.c(new_net_1352)
	);

	spl2 new_net_2167_v_fanout (
		.a(new_net_2167),
		.b(new_net_481),
		.c(new_net_478)
	);

	bfr new_net_3054_bfr_after (
		.din(n_0477_),
		.dout(new_net_3054)
	);

	bfr new_net_3055_bfr_after (
		.din(new_net_3054),
		.dout(new_net_3055)
	);

	bfr new_net_3056_bfr_after (
		.din(new_net_3055),
		.dout(new_net_3056)
	);

	bfr new_net_3057_bfr_after (
		.din(new_net_3056),
		.dout(new_net_3057)
	);

	bfr new_net_3058_bfr_after (
		.din(new_net_3057),
		.dout(new_net_3058)
	);

	bfr new_net_3059_bfr_after (
		.din(new_net_3058),
		.dout(new_net_3059)
	);

	bfr new_net_3060_bfr_after (
		.din(new_net_3059),
		.dout(new_net_3060)
	);

	bfr new_net_3061_bfr_after (
		.din(new_net_3060),
		.dout(new_net_3061)
	);

	bfr new_net_3062_bfr_after (
		.din(new_net_3061),
		.dout(new_net_3062)
	);

	bfr new_net_3063_bfr_after (
		.din(new_net_3062),
		.dout(new_net_3063)
	);

	bfr new_net_3064_bfr_after (
		.din(new_net_3063),
		.dout(new_net_3064)
	);

	bfr new_net_3065_bfr_after (
		.din(new_net_3064),
		.dout(new_net_3065)
	);

	bfr new_net_3066_bfr_after (
		.din(new_net_3065),
		.dout(new_net_3066)
	);

	bfr new_net_3067_bfr_after (
		.din(new_net_3066),
		.dout(new_net_3067)
	);

	bfr new_net_3068_bfr_after (
		.din(new_net_3067),
		.dout(new_net_3068)
	);

	bfr new_net_3069_bfr_after (
		.din(new_net_3068),
		.dout(new_net_3069)
	);

	bfr new_net_3070_bfr_after (
		.din(new_net_3069),
		.dout(new_net_3070)
	);

	bfr new_net_3071_bfr_after (
		.din(new_net_3070),
		.dout(new_net_3071)
	);

	bfr new_net_3072_bfr_after (
		.din(new_net_3071),
		.dout(new_net_3072)
	);

	bfr new_net_3073_bfr_after (
		.din(new_net_3072),
		.dout(new_net_3073)
	);

	bfr new_net_3074_bfr_after (
		.din(new_net_3073),
		.dout(new_net_3074)
	);

	bfr new_net_3075_bfr_after (
		.din(new_net_3074),
		.dout(new_net_3075)
	);

	bfr new_net_3076_bfr_after (
		.din(new_net_3075),
		.dout(new_net_3076)
	);

	bfr new_net_3077_bfr_after (
		.din(new_net_3076),
		.dout(new_net_3077)
	);

	bfr new_net_3078_bfr_after (
		.din(new_net_3077),
		.dout(new_net_3078)
	);

	bfr new_net_3079_bfr_after (
		.din(new_net_3078),
		.dout(new_net_3079)
	);

	bfr new_net_3080_bfr_after (
		.din(new_net_3079),
		.dout(new_net_3080)
	);

	bfr new_net_3081_bfr_after (
		.din(new_net_3080),
		.dout(new_net_3081)
	);

	bfr new_net_3082_bfr_after (
		.din(new_net_3081),
		.dout(new_net_3082)
	);

	bfr new_net_3083_bfr_after (
		.din(new_net_3082),
		.dout(new_net_3083)
	);

	bfr new_net_3084_bfr_after (
		.din(new_net_3083),
		.dout(new_net_3084)
	);

	bfr new_net_3085_bfr_after (
		.din(new_net_3084),
		.dout(new_net_3085)
	);

	bfr new_net_3086_bfr_after (
		.din(new_net_3085),
		.dout(new_net_3086)
	);

	bfr new_net_3087_bfr_after (
		.din(new_net_3086),
		.dout(new_net_3087)
	);

	bfr new_net_3088_bfr_after (
		.din(new_net_3087),
		.dout(new_net_3088)
	);

	bfr new_net_3089_bfr_after (
		.din(new_net_3088),
		.dout(new_net_3089)
	);

	bfr new_net_3090_bfr_after (
		.din(new_net_3089),
		.dout(new_net_3090)
	);

	bfr new_net_3091_bfr_after (
		.din(new_net_3090),
		.dout(new_net_3091)
	);

	bfr new_net_3092_bfr_after (
		.din(new_net_3091),
		.dout(new_net_3092)
	);

	spl2 n_0477__v_fanout (
		.a(new_net_3092),
		.b(new_net_99),
		.c(new_net_98)
	);

	spl2 n_0436__v_fanout (
		.a(n_0436_),
		.b(new_net_957),
		.c(new_net_956)
	);

	spl2 n_0445__v_fanout (
		.a(n_0445_),
		.b(new_net_1899),
		.c(new_net_1898)
	);

	spl2 n_0548__v_fanout (
		.a(n_0548_),
		.b(new_net_608),
		.c(new_net_607)
	);

	spl2 n_0629__v_fanout (
		.a(n_0629_),
		.b(new_net_861),
		.c(new_net_860)
	);

	bfr new_net_3093_bfr_before (
		.din(new_net_3093),
		.dout(new_net_29)
	);

	bfr new_net_3094_bfr_before (
		.din(new_net_3094),
		.dout(new_net_3093)
	);

	bfr new_net_3095_bfr_before (
		.din(new_net_3095),
		.dout(new_net_3094)
	);

	bfr new_net_3096_bfr_before (
		.din(new_net_3096),
		.dout(new_net_3095)
	);

	bfr new_net_3097_bfr_before (
		.din(new_net_3097),
		.dout(new_net_3096)
	);

	bfr new_net_3098_bfr_before (
		.din(new_net_3098),
		.dout(new_net_3097)
	);

	bfr new_net_3099_bfr_before (
		.din(new_net_3099),
		.dout(new_net_3098)
	);

	bfr new_net_3100_bfr_before (
		.din(new_net_3100),
		.dout(new_net_3099)
	);

	bfr new_net_3101_bfr_before (
		.din(new_net_3101),
		.dout(new_net_3100)
	);

	bfr new_net_3102_bfr_before (
		.din(new_net_3102),
		.dout(new_net_3101)
	);

	bfr new_net_3103_bfr_before (
		.din(new_net_3103),
		.dout(new_net_3102)
	);

	bfr new_net_3104_bfr_before (
		.din(new_net_3104),
		.dout(new_net_3103)
	);

	bfr new_net_3105_bfr_before (
		.din(new_net_3105),
		.dout(new_net_3104)
	);

	bfr new_net_3106_bfr_before (
		.din(new_net_3106),
		.dout(new_net_3105)
	);

	spl3L n_0010__v_fanout (
		.a(n_0010_),
		.b(new_net_30),
		.c(new_net_28),
		.d(new_net_3106)
	);

	bfr new_net_3107_bfr_before (
		.din(new_net_3107),
		.dout(new_net_555)
	);

	bfr new_net_3108_bfr_before (
		.din(new_net_3108),
		.dout(new_net_3107)
	);

	bfr new_net_3109_bfr_before (
		.din(new_net_3109),
		.dout(new_net_3108)
	);

	bfr new_net_3110_bfr_before (
		.din(new_net_3110),
		.dout(new_net_3109)
	);

	bfr new_net_3111_bfr_before (
		.din(new_net_3111),
		.dout(new_net_3110)
	);

	bfr new_net_3112_bfr_before (
		.din(new_net_3112),
		.dout(new_net_3111)
	);

	bfr new_net_3113_bfr_before (
		.din(new_net_3113),
		.dout(new_net_3112)
	);

	bfr new_net_3114_bfr_before (
		.din(new_net_3114),
		.dout(new_net_3113)
	);

	bfr new_net_3115_bfr_before (
		.din(new_net_3115),
		.dout(new_net_3114)
	);

	bfr new_net_3116_bfr_before (
		.din(new_net_3116),
		.dout(new_net_3115)
	);

	spl2 n_0344__v_fanout (
		.a(n_0344_),
		.b(new_net_556),
		.c(new_net_3116)
	);

	bfr new_net_3117_bfr_before (
		.din(new_net_3117),
		.dout(new_net_1107)
	);

	bfr new_net_3118_bfr_before (
		.din(new_net_3118),
		.dout(new_net_3117)
	);

	bfr new_net_3119_bfr_before (
		.din(new_net_3119),
		.dout(new_net_3118)
	);

	bfr new_net_3120_bfr_before (
		.din(new_net_3120),
		.dout(new_net_3119)
	);

	bfr new_net_3121_bfr_before (
		.din(new_net_3121),
		.dout(new_net_3120)
	);

	bfr new_net_3122_bfr_before (
		.din(new_net_3122),
		.dout(new_net_3121)
	);

	bfr new_net_3123_bfr_before (
		.din(new_net_3123),
		.dout(new_net_3122)
	);

	bfr new_net_3124_bfr_before (
		.din(new_net_3124),
		.dout(new_net_3123)
	);

	bfr new_net_3125_bfr_before (
		.din(new_net_3125),
		.dout(new_net_3124)
	);

	bfr new_net_3126_bfr_before (
		.din(new_net_3126),
		.dout(new_net_3125)
	);

	bfr new_net_3127_bfr_before (
		.din(new_net_3127),
		.dout(new_net_3126)
	);

	bfr new_net_3128_bfr_before (
		.din(new_net_3128),
		.dout(new_net_3127)
	);

	bfr new_net_3129_bfr_before (
		.din(new_net_3129),
		.dout(new_net_3128)
	);

	bfr new_net_3130_bfr_before (
		.din(new_net_3130),
		.dout(new_net_3129)
	);

	bfr new_net_3131_bfr_before (
		.din(new_net_3131),
		.dout(new_net_3130)
	);

	bfr new_net_3132_bfr_before (
		.din(new_net_3132),
		.dout(new_net_3131)
	);

	bfr new_net_3133_bfr_before (
		.din(new_net_3133),
		.dout(new_net_3132)
	);

	bfr new_net_3134_bfr_before (
		.din(new_net_3134),
		.dout(new_net_3133)
	);

	bfr new_net_3135_bfr_before (
		.din(new_net_3135),
		.dout(new_net_3134)
	);

	spl2 n_1312__v_fanout (
		.a(n_1312_),
		.b(new_net_3135),
		.c(new_net_1106)
	);

	bfr new_net_3136_bfr_before (
		.din(new_net_3136),
		.dout(new_net_737)
	);

	bfr new_net_3137_bfr_before (
		.din(new_net_3137),
		.dout(new_net_3136)
	);

	spl2 new_net_2108_v_fanout (
		.a(new_net_2108),
		.b(new_net_3137),
		.c(new_net_740)
	);

	bfr new_net_3138_bfr_before (
		.din(new_net_3138),
		.dout(new_net_1447)
	);

	spl2 n_0057__v_fanout (
		.a(n_0057_),
		.b(new_net_2166),
		.c(new_net_3138)
	);

	bfr new_net_3139_bfr_before (
		.din(new_net_3139),
		.dout(new_net_852)
	);

	spl2 n_0598__v_fanout (
		.a(n_0598_),
		.b(new_net_853),
		.c(new_net_3139)
	);

	bfr new_net_3140_bfr_before (
		.din(new_net_3140),
		.dout(new_net_492)
	);

	bfr new_net_3141_bfr_before (
		.din(new_net_3141),
		.dout(new_net_3140)
	);

	bfr new_net_3142_bfr_before (
		.din(new_net_3142),
		.dout(new_net_3141)
	);

	bfr new_net_3143_bfr_before (
		.din(new_net_3143),
		.dout(new_net_3142)
	);

	bfr new_net_3144_bfr_before (
		.din(new_net_3144),
		.dout(new_net_3143)
	);

	bfr new_net_3145_bfr_before (
		.din(new_net_3145),
		.dout(new_net_3144)
	);

	bfr new_net_3146_bfr_before (
		.din(new_net_3146),
		.dout(new_net_3145)
	);

	bfr new_net_3147_bfr_before (
		.din(new_net_3147),
		.dout(new_net_3146)
	);

	bfr new_net_3148_bfr_before (
		.din(new_net_3148),
		.dout(new_net_3147)
	);

	bfr new_net_3149_bfr_before (
		.din(new_net_3149),
		.dout(new_net_3148)
	);

	bfr new_net_3150_bfr_before (
		.din(new_net_3150),
		.dout(new_net_3149)
	);

	bfr new_net_3151_bfr_before (
		.din(new_net_3151),
		.dout(new_net_3150)
	);

	bfr new_net_3152_bfr_before (
		.din(new_net_3152),
		.dout(new_net_3151)
	);

	bfr new_net_3153_bfr_before (
		.din(new_net_3153),
		.dout(new_net_3152)
	);

	bfr new_net_3154_bfr_before (
		.din(new_net_3154),
		.dout(new_net_3153)
	);

	bfr new_net_3155_bfr_before (
		.din(new_net_3155),
		.dout(new_net_3154)
	);

	bfr new_net_3156_bfr_before (
		.din(new_net_3156),
		.dout(new_net_3155)
	);

	bfr new_net_3157_bfr_before (
		.din(new_net_3157),
		.dout(new_net_3156)
	);

	bfr new_net_3158_bfr_before (
		.din(new_net_3158),
		.dout(new_net_3157)
	);

	bfr new_net_3159_bfr_before (
		.din(new_net_3159),
		.dout(new_net_3158)
	);

	bfr new_net_3160_bfr_before (
		.din(new_net_3160),
		.dout(new_net_3159)
	);

	bfr new_net_3161_bfr_before (
		.din(new_net_3161),
		.dout(new_net_3160)
	);

	bfr new_net_3162_bfr_before (
		.din(new_net_3162),
		.dout(new_net_3161)
	);

	bfr new_net_3163_bfr_before (
		.din(new_net_3163),
		.dout(new_net_3162)
	);

	bfr new_net_3164_bfr_before (
		.din(new_net_3164),
		.dout(new_net_3163)
	);

	bfr new_net_3165_bfr_before (
		.din(new_net_3165),
		.dout(new_net_3164)
	);

	bfr new_net_3166_bfr_before (
		.din(new_net_3166),
		.dout(new_net_3165)
	);

	bfr new_net_3167_bfr_before (
		.din(new_net_3167),
		.dout(new_net_3166)
	);

	bfr new_net_3168_bfr_before (
		.din(new_net_3168),
		.dout(new_net_3167)
	);

	bfr new_net_3169_bfr_before (
		.din(new_net_3169),
		.dout(new_net_3168)
	);

	bfr new_net_3170_bfr_before (
		.din(new_net_3170),
		.dout(new_net_3169)
	);

	bfr new_net_3171_bfr_before (
		.din(new_net_3171),
		.dout(new_net_3170)
	);

	bfr new_net_3172_bfr_before (
		.din(new_net_3172),
		.dout(new_net_3171)
	);

	bfr new_net_3173_bfr_before (
		.din(new_net_3173),
		.dout(new_net_3172)
	);

	bfr new_net_3174_bfr_before (
		.din(new_net_3174),
		.dout(new_net_3173)
	);

	bfr new_net_3175_bfr_before (
		.din(new_net_3175),
		.dout(new_net_3174)
	);

	spl2 new_net_2164_v_fanout (
		.a(new_net_2164),
		.b(new_net_3175),
		.c(new_net_494)
	);

	spl2 n_1224__v_fanout (
		.a(n_1224_),
		.b(new_net_349),
		.c(new_net_348)
	);

	bfr new_net_3176_bfr_after (
		.din(n_0454_),
		.dout(new_net_3176)
	);

	bfr new_net_3177_bfr_after (
		.din(new_net_3176),
		.dout(new_net_3177)
	);

	bfr new_net_3178_bfr_after (
		.din(new_net_3177),
		.dout(new_net_3178)
	);

	bfr new_net_3179_bfr_after (
		.din(new_net_3178),
		.dout(new_net_3179)
	);

	bfr new_net_3180_bfr_after (
		.din(new_net_3179),
		.dout(new_net_3180)
	);

	bfr new_net_3181_bfr_after (
		.din(new_net_3180),
		.dout(new_net_3181)
	);

	spl2 n_0454__v_fanout (
		.a(new_net_3181),
		.b(new_net_1088),
		.c(new_net_1087)
	);

	bfr new_net_3182_bfr_after (
		.din(n_0582_),
		.dout(new_net_3182)
	);

	spl2 n_0582__v_fanout (
		.a(new_net_3182),
		.b(new_net_1639),
		.c(new_net_1638)
	);

	spl2 n_1271__v_fanout (
		.a(n_1271_),
		.b(new_net_296),
		.c(new_net_295)
	);

	spl2 n_0747__v_fanout (
		.a(n_0747_),
		.b(new_net_1850),
		.c(new_net_1849)
	);

	bfr new_net_3183_bfr_before (
		.din(new_net_3183),
		.dout(new_net_2139)
	);

	bfr new_net_3184_bfr_before (
		.din(new_net_3184),
		.dout(new_net_3183)
	);

	bfr new_net_3185_bfr_before (
		.din(new_net_3185),
		.dout(new_net_3184)
	);

	bfr new_net_3186_bfr_before (
		.din(new_net_3186),
		.dout(new_net_3185)
	);

	bfr new_net_3187_bfr_before (
		.din(new_net_3187),
		.dout(new_net_3186)
	);

	bfr new_net_3188_bfr_before (
		.din(new_net_3188),
		.dout(new_net_3187)
	);

	bfr new_net_3189_bfr_before (
		.din(new_net_3189),
		.dout(new_net_3188)
	);

	bfr new_net_3190_bfr_before (
		.din(new_net_3190),
		.dout(new_net_3189)
	);

	bfr new_net_3191_bfr_before (
		.din(new_net_3191),
		.dout(new_net_3190)
	);

	bfr new_net_3192_bfr_before (
		.din(new_net_3192),
		.dout(new_net_3191)
	);

	bfr new_net_3193_bfr_before (
		.din(new_net_3193),
		.dout(new_net_3192)
	);

	bfr new_net_3194_bfr_before (
		.din(new_net_3194),
		.dout(new_net_3193)
	);

	bfr new_net_3195_bfr_before (
		.din(new_net_3195),
		.dout(new_net_3194)
	);

	bfr new_net_3196_bfr_before (
		.din(new_net_3196),
		.dout(new_net_3195)
	);

	bfr new_net_3197_bfr_before (
		.din(new_net_3197),
		.dout(new_net_3196)
	);

	bfr new_net_3198_bfr_before (
		.din(new_net_3198),
		.dout(new_net_3197)
	);

	bfr new_net_3199_bfr_before (
		.din(new_net_3199),
		.dout(new_net_3198)
	);

	bfr new_net_3200_bfr_before (
		.din(new_net_3200),
		.dout(new_net_3199)
	);

	bfr new_net_3201_bfr_before (
		.din(new_net_3201),
		.dout(new_net_3200)
	);

	bfr new_net_3202_bfr_before (
		.din(new_net_3202),
		.dout(new_net_3201)
	);

	bfr new_net_3203_bfr_before (
		.din(new_net_3203),
		.dout(new_net_3202)
	);

	spl3L new_net_2138_v_fanout (
		.a(new_net_2138),
		.b(new_net_3203),
		.c(new_net_967),
		.d(new_net_971)
	);

	bfr new_net_3204_bfr_before (
		.din(new_net_3204),
		.dout(new_net_2169)
	);

	bfr new_net_3205_bfr_before (
		.din(new_net_3205),
		.dout(new_net_3204)
	);

	bfr new_net_3206_bfr_before (
		.din(new_net_3206),
		.dout(new_net_3205)
	);

	bfr new_net_3207_bfr_before (
		.din(new_net_3207),
		.dout(new_net_3206)
	);

	bfr new_net_3208_bfr_before (
		.din(new_net_3208),
		.dout(new_net_3207)
	);

	bfr new_net_3209_bfr_before (
		.din(new_net_3209),
		.dout(new_net_3208)
	);

	spl2 n_1336__v_fanout (
		.a(n_1336_),
		.b(new_net_3209),
		.c(new_net_1596)
	);

	spl2 n_0899__v_fanout (
		.a(n_0899_),
		.b(new_net_1212),
		.c(new_net_1211)
	);

	bfr new_net_3210_bfr_before (
		.din(new_net_3210),
		.dout(new_net_1509)
	);

	spl2 n_1355__v_fanout (
		.a(n_1355_),
		.b(new_net_2170),
		.c(new_net_3210)
	);

	bfr new_net_3211_bfr_before (
		.din(new_net_3211),
		.dout(new_net_360)
	);

	spl3L n_0701__v_fanout (
		.a(n_0701_),
		.b(new_net_361),
		.c(new_net_3211),
		.d(new_net_362)
	);

	bfr new_net_3212_bfr_after (
		.din(n_0503_),
		.dout(new_net_3212)
	);

	spl2 n_0503__v_fanout (
		.a(new_net_3212),
		.b(new_net_859),
		.c(new_net_858)
	);

	spl2 n_0108__v_fanout (
		.a(n_0108_),
		.b(new_net_2168),
		.c(new_net_2167)
	);

	spl2 n_0842__v_fanout (
		.a(n_0842_),
		.b(new_net_606),
		.c(new_net_605)
	);

	spl2 n_1176__v_fanout (
		.a(n_1176_),
		.b(new_net_1438),
		.c(new_net_1437)
	);

	bfr new_net_3213_bfr_after (
		.din(n_0421_),
		.dout(new_net_3213)
	);

	spl2 n_0421__v_fanout (
		.a(new_net_3213),
		.b(new_net_1894),
		.c(new_net_1893)
	);

	spl2 n_0538__v_fanout (
		.a(n_0538_),
		.b(new_net_1319),
		.c(new_net_1318)
	);

	bfr new_net_3214_bfr_after (
		.din(n_0147_),
		.dout(new_net_3214)
	);

	bfr new_net_3215_bfr_before (
		.din(new_net_3215),
		.dout(new_net_580)
	);

	bfr new_net_3216_bfr_before (
		.din(new_net_3216),
		.dout(new_net_3215)
	);

	bfr new_net_3217_bfr_before (
		.din(new_net_3217),
		.dout(new_net_3216)
	);

	bfr new_net_3218_bfr_before (
		.din(new_net_3218),
		.dout(new_net_3217)
	);

	bfr new_net_3219_bfr_before (
		.din(new_net_3219),
		.dout(new_net_3218)
	);

	bfr new_net_3220_bfr_before (
		.din(new_net_3220),
		.dout(new_net_3219)
	);

	bfr new_net_3221_bfr_before (
		.din(new_net_3221),
		.dout(new_net_3220)
	);

	bfr new_net_3222_bfr_before (
		.din(new_net_3222),
		.dout(new_net_3221)
	);

	bfr new_net_3223_bfr_before (
		.din(new_net_3223),
		.dout(new_net_3222)
	);

	bfr new_net_3224_bfr_before (
		.din(new_net_3224),
		.dout(new_net_3223)
	);

	bfr new_net_3225_bfr_before (
		.din(new_net_3225),
		.dout(new_net_3224)
	);

	bfr new_net_3226_bfr_before (
		.din(new_net_3226),
		.dout(new_net_3225)
	);

	bfr new_net_3227_bfr_before (
		.din(new_net_3227),
		.dout(new_net_3226)
	);

	spl2 n_0147__v_fanout (
		.a(new_net_3214),
		.b(new_net_581),
		.c(new_net_3227)
	);

	spl2 n_0532__v_fanout (
		.a(n_0532_),
		.b(new_net_709),
		.c(new_net_708)
	);

	bfr new_net_3228_bfr_after (
		.din(n_0066_),
		.dout(new_net_3228)
	);

	bfr new_net_3229_bfr_after (
		.din(new_net_3228),
		.dout(new_net_3229)
	);

	bfr new_net_3230_bfr_after (
		.din(new_net_3229),
		.dout(new_net_3230)
	);

	bfr new_net_3231_bfr_after (
		.din(new_net_3230),
		.dout(new_net_3231)
	);

	bfr new_net_3232_bfr_after (
		.din(new_net_3231),
		.dout(new_net_3232)
	);

	bfr new_net_3233_bfr_after (
		.din(new_net_3232),
		.dout(new_net_3233)
	);

	bfr new_net_3234_bfr_after (
		.din(new_net_3233),
		.dout(new_net_3234)
	);

	bfr new_net_3235_bfr_before (
		.din(new_net_3235),
		.dout(new_net_621)
	);

	spl2 n_0066__v_fanout (
		.a(new_net_3234),
		.b(new_net_3235),
		.c(new_net_620)
	);

	spl2 n_1117__v_fanout (
		.a(n_1117_),
		.b(new_net_359),
		.c(new_net_358)
	);

	bfr new_net_3236_bfr_before (
		.din(new_net_3236),
		.dout(new_net_2135)
	);

	bfr new_net_3237_bfr_before (
		.din(new_net_3237),
		.dout(new_net_3236)
	);

	bfr new_net_3238_bfr_before (
		.din(new_net_3238),
		.dout(new_net_3237)
	);

	bfr new_net_3239_bfr_before (
		.din(new_net_3239),
		.dout(new_net_3238)
	);

	bfr new_net_3240_bfr_before (
		.din(new_net_3240),
		.dout(new_net_3239)
	);

	bfr new_net_3241_bfr_before (
		.din(new_net_3241),
		.dout(new_net_3240)
	);

	bfr new_net_3242_bfr_before (
		.din(new_net_3242),
		.dout(new_net_3241)
	);

	bfr new_net_3243_bfr_before (
		.din(new_net_3243),
		.dout(new_net_3242)
	);

	bfr new_net_3244_bfr_before (
		.din(new_net_3244),
		.dout(new_net_3243)
	);

	bfr new_net_3245_bfr_before (
		.din(new_net_3245),
		.dout(new_net_3244)
	);

	bfr new_net_3246_bfr_before (
		.din(new_net_3246),
		.dout(new_net_3245)
	);

	bfr new_net_3247_bfr_before (
		.din(new_net_3247),
		.dout(new_net_3246)
	);

	bfr new_net_3248_bfr_before (
		.din(new_net_3248),
		.dout(new_net_3247)
	);

	bfr new_net_3249_bfr_before (
		.din(new_net_3249),
		.dout(new_net_3248)
	);

	bfr new_net_3250_bfr_before (
		.din(new_net_3250),
		.dout(new_net_3249)
	);

	bfr new_net_3251_bfr_before (
		.din(new_net_3251),
		.dout(new_net_3250)
	);

	bfr new_net_3252_bfr_before (
		.din(new_net_3252),
		.dout(new_net_3251)
	);

	bfr new_net_3253_bfr_before (
		.din(new_net_3253),
		.dout(new_net_3252)
	);

	bfr new_net_3254_bfr_before (
		.din(new_net_3254),
		.dout(new_net_3253)
	);

	bfr new_net_3255_bfr_before (
		.din(new_net_3255),
		.dout(new_net_3254)
	);

	bfr new_net_3256_bfr_before (
		.din(new_net_3256),
		.dout(new_net_3255)
	);

	bfr new_net_3257_bfr_before (
		.din(new_net_3257),
		.dout(new_net_3256)
	);

	bfr new_net_3258_bfr_before (
		.din(new_net_3258),
		.dout(new_net_3257)
	);

	bfr new_net_3259_bfr_before (
		.din(new_net_3259),
		.dout(new_net_3258)
	);

	bfr new_net_3260_bfr_before (
		.din(new_net_3260),
		.dout(new_net_3259)
	);

	bfr new_net_3261_bfr_before (
		.din(new_net_3261),
		.dout(new_net_3260)
	);

	bfr new_net_3262_bfr_before (
		.din(new_net_3262),
		.dout(new_net_3261)
	);

	bfr new_net_3263_bfr_before (
		.din(new_net_3263),
		.dout(new_net_3262)
	);

	bfr new_net_3264_bfr_before (
		.din(new_net_3264),
		.dout(new_net_3263)
	);

	bfr new_net_3265_bfr_before (
		.din(new_net_3265),
		.dout(new_net_3264)
	);

	bfr new_net_3266_bfr_before (
		.din(new_net_3266),
		.dout(new_net_3265)
	);

	bfr new_net_3267_bfr_before (
		.din(new_net_3267),
		.dout(new_net_3266)
	);

	bfr new_net_3268_bfr_before (
		.din(new_net_3268),
		.dout(new_net_3267)
	);

	spl3L new_net_2134_v_fanout (
		.a(new_net_2134),
		.b(new_net_3268),
		.c(new_net_473),
		.d(new_net_477)
	);

	bfr new_net_3269_bfr_before (
		.din(new_net_3269),
		.dout(new_net_469)
	);

	bfr new_net_3270_bfr_before (
		.din(new_net_3270),
		.dout(new_net_3269)
	);

	bfr new_net_3271_bfr_before (
		.din(new_net_3271),
		.dout(new_net_3270)
	);

	bfr new_net_3272_bfr_before (
		.din(new_net_3272),
		.dout(new_net_3271)
	);

	bfr new_net_3273_bfr_before (
		.din(new_net_3273),
		.dout(new_net_3272)
	);

	bfr new_net_3274_bfr_before (
		.din(new_net_3274),
		.dout(new_net_3273)
	);

	bfr new_net_3275_bfr_before (
		.din(new_net_3275),
		.dout(new_net_3274)
	);

	bfr new_net_3276_bfr_before (
		.din(new_net_3276),
		.dout(new_net_3275)
	);

	bfr new_net_3277_bfr_before (
		.din(new_net_3277),
		.dout(new_net_3276)
	);

	bfr new_net_3278_bfr_before (
		.din(new_net_3278),
		.dout(new_net_3277)
	);

	bfr new_net_3279_bfr_before (
		.din(new_net_3279),
		.dout(new_net_3278)
	);

	bfr new_net_3280_bfr_before (
		.din(new_net_3280),
		.dout(new_net_3279)
	);

	bfr new_net_3281_bfr_before (
		.din(new_net_3281),
		.dout(new_net_3280)
	);

	spl2 new_net_2154_v_fanout (
		.a(new_net_2154),
		.b(new_net_3281),
		.c(new_net_471)
	);

	bfr new_net_3282_bfr_after (
		.din(n_0431_),
		.dout(new_net_3282)
	);

	bfr new_net_3283_bfr_after (
		.din(new_net_3282),
		.dout(new_net_3283)
	);

	bfr new_net_3284_bfr_after (
		.din(new_net_3283),
		.dout(new_net_3284)
	);

	bfr new_net_3285_bfr_after (
		.din(new_net_3284),
		.dout(new_net_3285)
	);

	bfr new_net_3286_bfr_after (
		.din(new_net_3285),
		.dout(new_net_3286)
	);

	bfr new_net_3287_bfr_after (
		.din(new_net_3286),
		.dout(new_net_3287)
	);

	bfr new_net_3288_bfr_after (
		.din(new_net_3287),
		.dout(new_net_3288)
	);

	bfr new_net_3289_bfr_after (
		.din(new_net_3288),
		.dout(new_net_3289)
	);

	bfr new_net_3290_bfr_after (
		.din(new_net_3289),
		.dout(new_net_3290)
	);

	bfr new_net_3291_bfr_after (
		.din(new_net_3290),
		.dout(new_net_3291)
	);

	bfr new_net_3292_bfr_after (
		.din(new_net_3291),
		.dout(new_net_3292)
	);

	bfr new_net_3293_bfr_after (
		.din(new_net_3292),
		.dout(new_net_3293)
	);

	bfr new_net_3294_bfr_after (
		.din(new_net_3293),
		.dout(new_net_3294)
	);

	bfr new_net_3295_bfr_after (
		.din(new_net_3294),
		.dout(new_net_3295)
	);

	bfr new_net_3296_bfr_after (
		.din(new_net_3295),
		.dout(new_net_3296)
	);

	bfr new_net_3297_bfr_after (
		.din(new_net_3296),
		.dout(new_net_3297)
	);

	bfr new_net_3298_bfr_after (
		.din(new_net_3297),
		.dout(new_net_3298)
	);

	bfr new_net_3299_bfr_after (
		.din(new_net_3298),
		.dout(new_net_3299)
	);

	bfr new_net_3300_bfr_after (
		.din(new_net_3299),
		.dout(new_net_3300)
	);

	bfr new_net_3301_bfr_after (
		.din(new_net_3300),
		.dout(new_net_3301)
	);

	bfr new_net_3302_bfr_after (
		.din(new_net_3301),
		.dout(new_net_3302)
	);

	bfr new_net_3303_bfr_after (
		.din(new_net_3302),
		.dout(new_net_3303)
	);

	bfr new_net_3304_bfr_after (
		.din(new_net_3303),
		.dout(new_net_3304)
	);

	bfr new_net_3305_bfr_after (
		.din(new_net_3304),
		.dout(new_net_3305)
	);

	bfr new_net_3306_bfr_after (
		.din(new_net_3305),
		.dout(new_net_3306)
	);

	bfr new_net_3307_bfr_after (
		.din(new_net_3306),
		.dout(new_net_3307)
	);

	bfr new_net_3308_bfr_after (
		.din(new_net_3307),
		.dout(new_net_3308)
	);

	bfr new_net_3309_bfr_after (
		.din(new_net_3308),
		.dout(new_net_3309)
	);

	bfr new_net_3310_bfr_after (
		.din(new_net_3309),
		.dout(new_net_3310)
	);

	bfr new_net_3311_bfr_after (
		.din(new_net_3310),
		.dout(new_net_3311)
	);

	spl2 n_0431__v_fanout (
		.a(new_net_3311),
		.b(new_net_369),
		.c(new_net_368)
	);

	bfr new_net_3312_bfr_after (
		.din(n_0479_),
		.dout(new_net_3312)
	);

	bfr new_net_3313_bfr_after (
		.din(new_net_3312),
		.dout(new_net_3313)
	);

	bfr new_net_3314_bfr_after (
		.din(new_net_3313),
		.dout(new_net_3314)
	);

	bfr new_net_3315_bfr_after (
		.din(new_net_3314),
		.dout(new_net_3315)
	);

	bfr new_net_3316_bfr_after (
		.din(new_net_3315),
		.dout(new_net_3316)
	);

	spl2 n_0479__v_fanout (
		.a(new_net_3316),
		.b(new_net_290),
		.c(new_net_289)
	);

	bfr new_net_3317_bfr_after (
		.din(n_0564_),
		.dout(new_net_3317)
	);

	bfr new_net_3318_bfr_after (
		.din(new_net_3317),
		.dout(new_net_3318)
	);

	bfr new_net_3319_bfr_after (
		.din(new_net_3318),
		.dout(new_net_3319)
	);

	bfr new_net_3320_bfr_after (
		.din(new_net_3319),
		.dout(new_net_3320)
	);

	spl2 n_0564__v_fanout (
		.a(new_net_3320),
		.b(new_net_1238),
		.c(new_net_1237)
	);

	bfr new_net_3321_bfr_before (
		.din(new_net_3321),
		.dout(new_net_963)
	);

	bfr new_net_3322_bfr_before (
		.din(new_net_3322),
		.dout(new_net_3321)
	);

	bfr new_net_3323_bfr_before (
		.din(new_net_3323),
		.dout(new_net_3322)
	);

	bfr new_net_3324_bfr_before (
		.din(new_net_3324),
		.dout(new_net_3323)
	);

	bfr new_net_3325_bfr_before (
		.din(new_net_3325),
		.dout(new_net_3324)
	);

	bfr new_net_3326_bfr_before (
		.din(new_net_3326),
		.dout(new_net_3325)
	);

	bfr new_net_3327_bfr_before (
		.din(new_net_3327),
		.dout(new_net_3326)
	);

	spl2 new_net_2055_v_fanout (
		.a(new_net_2055),
		.b(new_net_3327),
		.c(new_net_961)
	);

	bfr new_net_3328_bfr_after (
		.din(n_0082_),
		.dout(new_net_3328)
	);

	bfr new_net_3329_bfr_after (
		.din(new_net_3328),
		.dout(new_net_3329)
	);

	bfr new_net_3330_bfr_before (
		.din(new_net_3330),
		.dout(new_net_1715)
	);

	bfr new_net_3331_bfr_before (
		.din(new_net_3331),
		.dout(new_net_3330)
	);

	bfr new_net_3332_bfr_before (
		.din(new_net_3332),
		.dout(new_net_3331)
	);

	bfr new_net_3333_bfr_before (
		.din(new_net_3333),
		.dout(new_net_3332)
	);

	bfr new_net_3334_bfr_before (
		.din(new_net_3334),
		.dout(new_net_3333)
	);

	bfr new_net_3335_bfr_before (
		.din(new_net_3335),
		.dout(new_net_3334)
	);

	bfr new_net_3336_bfr_before (
		.din(new_net_3336),
		.dout(new_net_3335)
	);

	bfr new_net_3337_bfr_before (
		.din(new_net_3337),
		.dout(new_net_3336)
	);

	bfr new_net_3338_bfr_before (
		.din(new_net_3338),
		.dout(new_net_3337)
	);

	bfr new_net_3339_bfr_before (
		.din(new_net_3339),
		.dout(new_net_3338)
	);

	bfr new_net_3340_bfr_before (
		.din(new_net_3340),
		.dout(new_net_3339)
	);

	bfr new_net_3341_bfr_before (
		.din(new_net_3341),
		.dout(new_net_3340)
	);

	bfr new_net_3342_bfr_before (
		.din(new_net_3342),
		.dout(new_net_3341)
	);

	bfr new_net_3343_bfr_before (
		.din(new_net_3343),
		.dout(new_net_3342)
	);

	bfr new_net_3344_bfr_before (
		.din(new_net_3344),
		.dout(new_net_3343)
	);

	bfr new_net_3345_bfr_before (
		.din(new_net_3345),
		.dout(new_net_3344)
	);

	bfr new_net_3346_bfr_before (
		.din(new_net_3346),
		.dout(new_net_3345)
	);

	bfr new_net_3347_bfr_before (
		.din(new_net_3347),
		.dout(new_net_3346)
	);

	bfr new_net_3348_bfr_before (
		.din(new_net_3348),
		.dout(new_net_3347)
	);

	bfr new_net_3349_bfr_before (
		.din(new_net_3349),
		.dout(new_net_3348)
	);

	bfr new_net_3350_bfr_before (
		.din(new_net_3350),
		.dout(new_net_3349)
	);

	bfr new_net_3351_bfr_before (
		.din(new_net_3351),
		.dout(new_net_3350)
	);

	bfr new_net_3352_bfr_before (
		.din(new_net_3352),
		.dout(new_net_3351)
	);

	bfr new_net_3353_bfr_before (
		.din(new_net_3353),
		.dout(new_net_3352)
	);

	bfr new_net_3354_bfr_before (
		.din(new_net_3354),
		.dout(new_net_3353)
	);

	spl2 n_0082__v_fanout (
		.a(new_net_3329),
		.b(new_net_1716),
		.c(new_net_3354)
	);

	spl2 n_1039__v_fanout (
		.a(n_1039_),
		.b(new_net_1691),
		.c(new_net_1690)
	);

	bfr new_net_3355_bfr_before (
		.din(new_net_3355),
		.dout(new_net_2129)
	);

	bfr new_net_3356_bfr_before (
		.din(new_net_3356),
		.dout(new_net_3355)
	);

	bfr new_net_3357_bfr_before (
		.din(new_net_3357),
		.dout(new_net_3356)
	);

	bfr new_net_3358_bfr_before (
		.din(new_net_3358),
		.dout(new_net_3357)
	);

	bfr new_net_3359_bfr_before (
		.din(new_net_3359),
		.dout(new_net_3358)
	);

	bfr new_net_3360_bfr_before (
		.din(new_net_3360),
		.dout(new_net_3359)
	);

	bfr new_net_3361_bfr_before (
		.din(new_net_3361),
		.dout(new_net_3360)
	);

	bfr new_net_3362_bfr_before (
		.din(new_net_3362),
		.dout(new_net_3361)
	);

	bfr new_net_3363_bfr_before (
		.din(new_net_3363),
		.dout(new_net_3362)
	);

	bfr new_net_3364_bfr_before (
		.din(new_net_3364),
		.dout(new_net_3363)
	);

	bfr new_net_3365_bfr_before (
		.din(new_net_3365),
		.dout(new_net_3364)
	);

	bfr new_net_3366_bfr_before (
		.din(new_net_3366),
		.dout(new_net_3365)
	);

	bfr new_net_3367_bfr_before (
		.din(new_net_3367),
		.dout(new_net_3366)
	);

	bfr new_net_3368_bfr_before (
		.din(new_net_3368),
		.dout(new_net_3367)
	);

	bfr new_net_3369_bfr_before (
		.din(new_net_3369),
		.dout(new_net_3368)
	);

	bfr new_net_3370_bfr_before (
		.din(new_net_3370),
		.dout(new_net_3369)
	);

	bfr new_net_3371_bfr_before (
		.din(new_net_3371),
		.dout(new_net_3370)
	);

	bfr new_net_3372_bfr_before (
		.din(new_net_3372),
		.dout(new_net_3371)
	);

	bfr new_net_3373_bfr_before (
		.din(new_net_3373),
		.dout(new_net_3372)
	);

	bfr new_net_3374_bfr_before (
		.din(new_net_3374),
		.dout(new_net_3373)
	);

	bfr new_net_3375_bfr_before (
		.din(new_net_3375),
		.dout(new_net_3374)
	);

	bfr new_net_3376_bfr_before (
		.din(new_net_3376),
		.dout(new_net_3375)
	);

	bfr new_net_3377_bfr_before (
		.din(new_net_3377),
		.dout(new_net_3376)
	);

	bfr new_net_3378_bfr_before (
		.din(new_net_3378),
		.dout(new_net_3377)
	);

	bfr new_net_3379_bfr_before (
		.din(new_net_3379),
		.dout(new_net_3378)
	);

	bfr new_net_3380_bfr_before (
		.din(new_net_3380),
		.dout(new_net_3379)
	);

	bfr new_net_3381_bfr_before (
		.din(new_net_3381),
		.dout(new_net_3380)
	);

	bfr new_net_3382_bfr_before (
		.din(new_net_3382),
		.dout(new_net_3381)
	);

	bfr new_net_3383_bfr_before (
		.din(new_net_3383),
		.dout(new_net_3382)
	);

	bfr new_net_3384_bfr_before (
		.din(new_net_3384),
		.dout(new_net_3383)
	);

	bfr new_net_3385_bfr_before (
		.din(new_net_3385),
		.dout(new_net_3384)
	);

	bfr new_net_3386_bfr_before (
		.din(new_net_3386),
		.dout(new_net_3385)
	);

	bfr new_net_3387_bfr_before (
		.din(new_net_3387),
		.dout(new_net_3386)
	);

	bfr new_net_3388_bfr_before (
		.din(new_net_3388),
		.dout(new_net_3387)
	);

	bfr new_net_3389_bfr_before (
		.din(new_net_3389),
		.dout(new_net_3388)
	);

	bfr new_net_3390_bfr_before (
		.din(new_net_3390),
		.dout(new_net_3389)
	);

	bfr new_net_3391_bfr_before (
		.din(new_net_3391),
		.dout(new_net_3390)
	);

	bfr new_net_3392_bfr_before (
		.din(new_net_3392),
		.dout(new_net_3391)
	);

	bfr new_net_3393_bfr_before (
		.din(new_net_3393),
		.dout(new_net_3392)
	);

	spl2 new_net_2128_v_fanout (
		.a(new_net_2128),
		.b(new_net_3393),
		.c(new_net_675)
	);

	spl2 n_0618__v_fanout (
		.a(n_0618_),
		.b(new_net_1161),
		.c(new_net_1160)
	);

	spl2 n_1002__v_fanout (
		.a(n_1002_),
		.b(new_net_755),
		.c(new_net_754)
	);

	bfr new_net_3394_bfr_after (
		.din(n_0633_),
		.dout(new_net_3394)
	);

	bfr new_net_3395_bfr_after (
		.din(new_net_3394),
		.dout(new_net_3395)
	);

	spl2 n_0633__v_fanout (
		.a(new_net_3395),
		.b(new_net_979),
		.c(new_net_978)
	);

	spl2 n_0009__v_fanout (
		.a(n_0009_),
		.b(new_net_21),
		.c(new_net_20)
	);

	bfr new_net_3396_bfr_after (
		.din(n_0574_),
		.dout(new_net_3396)
	);

	bfr new_net_3397_bfr_after (
		.din(new_net_3396),
		.dout(new_net_3397)
	);

	bfr new_net_3398_bfr_after (
		.din(new_net_3397),
		.dout(new_net_3398)
	);

	bfr new_net_3399_bfr_after (
		.din(new_net_3398),
		.dout(new_net_3399)
	);

	bfr new_net_3400_bfr_after (
		.din(new_net_3399),
		.dout(new_net_3400)
	);

	bfr new_net_3401_bfr_after (
		.din(new_net_3400),
		.dout(new_net_3401)
	);

	bfr new_net_3402_bfr_after (
		.din(new_net_3401),
		.dout(new_net_3402)
	);

	bfr new_net_3403_bfr_after (
		.din(new_net_3402),
		.dout(new_net_3403)
	);

	bfr new_net_3404_bfr_after (
		.din(new_net_3403),
		.dout(new_net_3404)
	);

	bfr new_net_3405_bfr_after (
		.din(new_net_3404),
		.dout(new_net_3405)
	);

	bfr new_net_3406_bfr_after (
		.din(new_net_3405),
		.dout(new_net_3406)
	);

	bfr new_net_3407_bfr_after (
		.din(new_net_3406),
		.dout(new_net_3407)
	);

	bfr new_net_3408_bfr_after (
		.din(new_net_3407),
		.dout(new_net_3408)
	);

	bfr new_net_3409_bfr_after (
		.din(new_net_3408),
		.dout(new_net_3409)
	);

	bfr new_net_3410_bfr_after (
		.din(new_net_3409),
		.dout(new_net_3410)
	);

	bfr new_net_3411_bfr_after (
		.din(new_net_3410),
		.dout(new_net_3411)
	);

	bfr new_net_3412_bfr_after (
		.din(new_net_3411),
		.dout(new_net_3412)
	);

	bfr new_net_3413_bfr_after (
		.din(new_net_3412),
		.dout(new_net_3413)
	);

	spl2 n_0574__v_fanout (
		.a(new_net_3413),
		.b(new_net_1478),
		.c(new_net_1477)
	);

	bfr new_net_3414_bfr_before (
		.din(new_net_3414),
		.dout(new_net_2146)
	);

	bfr new_net_3415_bfr_before (
		.din(new_net_3415),
		.dout(new_net_3414)
	);

	bfr new_net_3416_bfr_before (
		.din(new_net_3416),
		.dout(new_net_3415)
	);

	spl2 new_net_2145_v_fanout (
		.a(new_net_2145),
		.b(new_net_3416),
		.c(new_net_1076)
	);

	bfr new_net_3417_bfr_before (
		.din(new_net_3417),
		.dout(new_net_1472)
	);

	bfr new_net_3418_bfr_before (
		.din(new_net_3418),
		.dout(new_net_3417)
	);

	spl2 new_net_2163_v_fanout (
		.a(new_net_2163),
		.b(new_net_3418),
		.c(new_net_1471)
	);

	bfr new_net_3419_bfr_before (
		.din(new_net_3419),
		.dout(new_net_2165)
	);

	bfr new_net_3420_bfr_before (
		.din(new_net_3420),
		.dout(new_net_3419)
	);

	bfr new_net_3421_bfr_before (
		.din(new_net_3421),
		.dout(new_net_3420)
	);

	bfr new_net_3422_bfr_before (
		.din(new_net_3422),
		.dout(new_net_3421)
	);

	bfr new_net_3423_bfr_before (
		.din(new_net_3423),
		.dout(new_net_3422)
	);

	spl3L n_0587__v_fanout (
		.a(n_0587_),
		.b(new_net_3423),
		.c(new_net_1735),
		.d(new_net_1738)
	);

	bfr new_net_3424_bfr_before (
		.din(new_net_3424),
		.dout(new_net_2164)
	);

	spl2 n_0114__v_fanout (
		.a(n_0114_),
		.b(new_net_493),
		.c(new_net_3424)
	);

	spl3L n_0694__v_fanout (
		.a(n_0694_),
		.b(new_net_1456),
		.c(new_net_1454),
		.d(new_net_1455)
	);

	spl2 n_0456__v_fanout (
		.a(n_0456_),
		.b(new_net_1631),
		.c(new_net_1630)
	);

	bfr new_net_3425_bfr_after (
		.din(n_0398_),
		.dout(new_net_3425)
	);

	bfr new_net_3426_bfr_after (
		.din(new_net_3425),
		.dout(new_net_3426)
	);

	bfr new_net_3427_bfr_after (
		.din(new_net_3426),
		.dout(new_net_3427)
	);

	bfr new_net_3428_bfr_after (
		.din(new_net_3427),
		.dout(new_net_3428)
	);

	bfr new_net_3429_bfr_after (
		.din(new_net_3428),
		.dout(new_net_3429)
	);

	spl2 n_0398__v_fanout (
		.a(new_net_3429),
		.b(new_net_1287),
		.c(new_net_1286)
	);

	bfr new_net_3430_bfr_after (
		.din(n_0409_),
		.dout(new_net_3430)
	);

	bfr new_net_3431_bfr_after (
		.din(new_net_3430),
		.dout(new_net_3431)
	);

	bfr new_net_3432_bfr_after (
		.din(new_net_3431),
		.dout(new_net_3432)
	);

	bfr new_net_3433_bfr_after (
		.din(new_net_3432),
		.dout(new_net_3433)
	);

	spl2 n_0409__v_fanout (
		.a(new_net_3433),
		.b(new_net_1539),
		.c(new_net_1538)
	);

	bfr new_net_3434_bfr_after (
		.din(n_0491_),
		.dout(new_net_3434)
	);

	bfr new_net_3435_bfr_after (
		.din(new_net_3434),
		.dout(new_net_3435)
	);

	bfr new_net_3436_bfr_after (
		.din(new_net_3435),
		.dout(new_net_3436)
	);

	bfr new_net_3437_bfr_after (
		.din(new_net_3436),
		.dout(new_net_3437)
	);

	spl2 n_0491__v_fanout (
		.a(new_net_3437),
		.b(new_net_601),
		.c(new_net_600)
	);

	spl2 n_0035__v_fanout (
		.a(n_0035_),
		.b(new_net_726),
		.c(new_net_725)
	);

	spl2 n_0442__v_fanout (
		.a(n_0442_),
		.b(new_net_1593),
		.c(new_net_1592)
	);

	spl2 n_1327__v_fanout (
		.a(n_1327_),
		.b(new_net_1956),
		.c(new_net_1955)
	);

	spl2 n_0712__v_fanout (
		.a(n_0712_),
		.b(new_net_1710),
		.c(new_net_1709)
	);

	spl2 n_0523__v_fanout (
		.a(n_0523_),
		.b(new_net_1256),
		.c(new_net_1255)
	);

	bfr new_net_3438_bfr_after (
		.din(n_0551_),
		.dout(new_net_3438)
	);

	bfr new_net_3439_bfr_after (
		.din(new_net_3438),
		.dout(new_net_3439)
	);

	bfr new_net_3440_bfr_after (
		.din(new_net_3439),
		.dout(new_net_3440)
	);

	spl2 n_0551__v_fanout (
		.a(new_net_3440),
		.b(new_net_931),
		.c(new_net_930)
	);

	bfr new_net_3441_bfr_after (
		.din(n_0647_),
		.dout(new_net_3441)
	);

	bfr new_net_3442_bfr_after (
		.din(new_net_3441),
		.dout(new_net_3442)
	);

	bfr new_net_3443_bfr_after (
		.din(new_net_3442),
		.dout(new_net_3443)
	);

	bfr new_net_3444_bfr_after (
		.din(new_net_3443),
		.dout(new_net_3444)
	);

	bfr new_net_3445_bfr_after (
		.din(new_net_3444),
		.dout(new_net_3445)
	);

	bfr new_net_3446_bfr_after (
		.din(new_net_3445),
		.dout(new_net_3446)
	);

	bfr new_net_3447_bfr_after (
		.din(new_net_3446),
		.dout(new_net_3447)
	);

	bfr new_net_3448_bfr_after (
		.din(new_net_3447),
		.dout(new_net_3448)
	);

	bfr new_net_3449_bfr_after (
		.din(new_net_3448),
		.dout(new_net_3449)
	);

	bfr new_net_3450_bfr_after (
		.din(new_net_3449),
		.dout(new_net_3450)
	);

	bfr new_net_3451_bfr_after (
		.din(new_net_3450),
		.dout(new_net_3451)
	);

	bfr new_net_3452_bfr_after (
		.din(new_net_3451),
		.dout(new_net_3452)
	);

	bfr new_net_3453_bfr_after (
		.din(new_net_3452),
		.dout(new_net_3453)
	);

	bfr new_net_3454_bfr_after (
		.din(new_net_3453),
		.dout(new_net_3454)
	);

	spl2 n_0647__v_fanout (
		.a(new_net_3454),
		.b(new_net_836),
		.c(new_net_835)
	);

	spl2 n_0279__v_fanout (
		.a(n_0279_),
		.b(new_net_1436),
		.c(new_net_1435)
	);

	spl2 n_0439__v_fanout (
		.a(n_0439_),
		.b(new_net_1271),
		.c(new_net_1270)
	);

	spl2 n_0520__v_fanout (
		.a(n_0520_),
		.b(new_net_1203),
		.c(new_net_1202)
	);

	bfr new_net_3455_bfr_before (
		.din(new_net_3455),
		.dout(new_net_2151)
	);

	bfr new_net_3456_bfr_before (
		.din(new_net_3456),
		.dout(new_net_3455)
	);

	bfr new_net_3457_bfr_before (
		.din(new_net_3457),
		.dout(new_net_3456)
	);

	bfr new_net_3458_bfr_before (
		.din(new_net_3458),
		.dout(new_net_3457)
	);

	bfr new_net_3459_bfr_before (
		.din(new_net_3459),
		.dout(new_net_3458)
	);

	bfr new_net_3460_bfr_before (
		.din(new_net_3460),
		.dout(new_net_3459)
	);

	bfr new_net_3461_bfr_before (
		.din(new_net_3461),
		.dout(new_net_3460)
	);

	bfr new_net_3462_bfr_before (
		.din(new_net_3462),
		.dout(new_net_3461)
	);

	bfr new_net_3463_bfr_before (
		.din(new_net_3463),
		.dout(new_net_3462)
	);

	bfr new_net_3464_bfr_before (
		.din(new_net_3464),
		.dout(new_net_3463)
	);

	bfr new_net_3465_bfr_before (
		.din(new_net_3465),
		.dout(new_net_3464)
	);

	bfr new_net_3466_bfr_before (
		.din(new_net_3466),
		.dout(new_net_3465)
	);

	bfr new_net_3467_bfr_before (
		.din(new_net_3467),
		.dout(new_net_3466)
	);

	bfr new_net_3468_bfr_before (
		.din(new_net_3468),
		.dout(new_net_3467)
	);

	bfr new_net_3469_bfr_before (
		.din(new_net_3469),
		.dout(new_net_3468)
	);

	bfr new_net_3470_bfr_before (
		.din(new_net_3470),
		.dout(new_net_3469)
	);

	bfr new_net_3471_bfr_before (
		.din(new_net_3471),
		.dout(new_net_3470)
	);

	bfr new_net_3472_bfr_before (
		.din(new_net_3472),
		.dout(new_net_3471)
	);

	bfr new_net_3473_bfr_before (
		.din(new_net_3473),
		.dout(new_net_3472)
	);

	bfr new_net_3474_bfr_before (
		.din(new_net_3474),
		.dout(new_net_3473)
	);

	spl2 new_net_2150_v_fanout (
		.a(new_net_2150),
		.b(new_net_3474),
		.c(new_net_898)
	);

	spl2 n_0474__v_fanout (
		.a(n_0474_),
		.b(new_net_1567),
		.c(new_net_1566)
	);

	spl3L n_0700__v_fanout (
		.a(n_0700_),
		.b(new_net_2163),
		.c(new_net_1469),
		.d(new_net_1470)
	);

	bfr new_net_3475_bfr_before (
		.din(new_net_3475),
		.dout(new_net_2108)
	);

	spl2 new_net_2107_v_fanout (
		.a(new_net_2107),
		.b(new_net_3475),
		.c(new_net_739)
	);

	spl2 new_net_2143_v_fanout (
		.a(new_net_2143),
		.b(new_net_1175),
		.c(new_net_1172)
	);

	spl3L n_1371__v_fanout (
		.a(n_1371_),
		.b(new_net_1399),
		.c(new_net_1398),
		.d(new_net_1400)
	);

	bfr new_net_3476_bfr_after (
		.din(n_1241_),
		.dout(new_net_3476)
	);

	bfr new_net_3477_bfr_after (
		.din(new_net_3476),
		.dout(new_net_3477)
	);

	bfr new_net_3478_bfr_after (
		.din(new_net_3477),
		.dout(new_net_3478)
	);

	spl2 n_1241__v_fanout (
		.a(new_net_3478),
		.b(new_net_592),
		.c(new_net_591)
	);

	spl2 n_0065__v_fanout (
		.a(n_0065_),
		.b(new_net_502),
		.c(new_net_501)
	);

	spl2 n_0744__v_fanout (
		.a(n_0744_),
		.b(new_net_1565),
		.c(new_net_1564)
	);

	spl2 n_0795__v_fanout (
		.a(n_0795_),
		.b(new_net_1746),
		.c(new_net_1745)
	);

	spl2 n_0229__v_fanout (
		.a(n_0229_),
		.b(new_net_1525),
		.c(new_net_1524)
	);

	spl2 new_net_2144_v_fanout (
		.a(new_net_2144),
		.b(new_net_1285),
		.c(new_net_1283)
	);

	spl2 n_0500__v_fanout (
		.a(n_0500_),
		.b(new_net_792),
		.c(new_net_791)
	);

	spl2 n_0839__v_fanout (
		.a(n_0839_),
		.b(new_net_1740),
		.c(new_net_1739)
	);

	bfr new_net_3479_bfr_after (
		.din(n_0616_),
		.dout(new_net_3479)
	);

	bfr new_net_3480_bfr_after (
		.din(new_net_3479),
		.dout(new_net_3480)
	);

	bfr new_net_3481_bfr_after (
		.din(new_net_3480),
		.dout(new_net_3481)
	);

	bfr new_net_3482_bfr_after (
		.din(new_net_3481),
		.dout(new_net_3482)
	);

	bfr new_net_3483_bfr_after (
		.din(new_net_3482),
		.dout(new_net_3483)
	);

	spl2 n_0616__v_fanout (
		.a(new_net_3483),
		.b(new_net_965),
		.c(new_net_964)
	);

	spl2 n_1268__v_fanout (
		.a(n_1268_),
		.b(new_net_1647),
		.c(new_net_1646)
	);

	bfr new_net_3484_bfr_before (
		.din(new_net_3484),
		.dout(new_net_1009)
	);

	spl2 n_1335__v_fanout (
		.a(n_1335_),
		.b(new_net_1010),
		.c(new_net_3484)
	);

	bfr new_net_3485_bfr_before (
		.din(new_net_3485),
		.dout(new_net_1951)
	);

	spl2 n_0002__v_fanout (
		.a(n_0002_),
		.b(new_net_1952),
		.c(new_net_3485)
	);

	bfr new_net_3486_bfr_after (
		.din(n_0080_),
		.dout(new_net_3486)
	);

	bfr new_net_3487_bfr_after (
		.din(new_net_3486),
		.dout(new_net_3487)
	);

	bfr new_net_3488_bfr_after (
		.din(new_net_3487),
		.dout(new_net_3488)
	);

	bfr new_net_3489_bfr_after (
		.din(new_net_3488),
		.dout(new_net_3489)
	);

	bfr new_net_3490_bfr_after (
		.din(new_net_3489),
		.dout(new_net_3490)
	);

	bfr new_net_3491_bfr_after (
		.din(new_net_3490),
		.dout(new_net_3491)
	);

	bfr new_net_3492_bfr_after (
		.din(new_net_3491),
		.dout(new_net_3492)
	);

	bfr new_net_3493_bfr_after (
		.din(new_net_3492),
		.dout(new_net_3493)
	);

	bfr new_net_3494_bfr_after (
		.din(new_net_3493),
		.dout(new_net_3494)
	);

	bfr new_net_3495_bfr_after (
		.din(new_net_3494),
		.dout(new_net_3495)
	);

	bfr new_net_3496_bfr_after (
		.din(new_net_3495),
		.dout(new_net_3496)
	);

	bfr new_net_3497_bfr_after (
		.din(new_net_3496),
		.dout(new_net_3497)
	);

	bfr new_net_3498_bfr_after (
		.din(new_net_3497),
		.dout(new_net_3498)
	);

	bfr new_net_3499_bfr_after (
		.din(new_net_3498),
		.dout(new_net_3499)
	);

	bfr new_net_3500_bfr_after (
		.din(new_net_3499),
		.dout(new_net_3500)
	);

	bfr new_net_3501_bfr_after (
		.din(new_net_3500),
		.dout(new_net_3501)
	);

	bfr new_net_3502_bfr_after (
		.din(new_net_3501),
		.dout(new_net_3502)
	);

	bfr new_net_3503_bfr_after (
		.din(new_net_3502),
		.dout(new_net_3503)
	);

	bfr new_net_3504_bfr_after (
		.din(new_net_3503),
		.dout(new_net_3504)
	);

	bfr new_net_3505_bfr_after (
		.din(new_net_3504),
		.dout(new_net_3505)
	);

	bfr new_net_3506_bfr_after (
		.din(new_net_3505),
		.dout(new_net_3506)
	);

	bfr new_net_3507_bfr_after (
		.din(new_net_3506),
		.dout(new_net_3507)
	);

	bfr new_net_3508_bfr_after (
		.din(new_net_3507),
		.dout(new_net_3508)
	);

	bfr new_net_3509_bfr_after (
		.din(new_net_3508),
		.dout(new_net_3509)
	);

	bfr new_net_3510_bfr_after (
		.din(new_net_3509),
		.dout(new_net_3510)
	);

	bfr new_net_3511_bfr_after (
		.din(new_net_3510),
		.dout(new_net_3511)
	);

	bfr new_net_3512_bfr_after (
		.din(new_net_3511),
		.dout(new_net_3512)
	);

	bfr new_net_3513_bfr_after (
		.din(new_net_3512),
		.dout(new_net_3513)
	);

	bfr new_net_3514_bfr_after (
		.din(new_net_3513),
		.dout(new_net_3514)
	);

	bfr new_net_3515_bfr_after (
		.din(new_net_3514),
		.dout(new_net_3515)
	);

	bfr new_net_3516_bfr_after (
		.din(new_net_3515),
		.dout(new_net_3516)
	);

	bfr new_net_3517_bfr_before (
		.din(new_net_3517),
		.dout(new_net_2158)
	);

	spl2 n_0080__v_fanout (
		.a(new_net_3516),
		.b(new_net_3517),
		.c(new_net_1681)
	);

	spl2 n_0321__v_fanout (
		.a(n_0321_),
		.b(new_net_1708),
		.c(new_net_1707)
	);

	bfr new_net_3518_bfr_before (
		.din(new_net_3518),
		.dout(new_net_814)
	);

	bfr new_net_3519_bfr_before (
		.din(new_net_3519),
		.dout(new_net_3518)
	);

	bfr new_net_3520_bfr_before (
		.din(new_net_3520),
		.dout(new_net_3519)
	);

	bfr new_net_3521_bfr_before (
		.din(new_net_3521),
		.dout(new_net_3520)
	);

	bfr new_net_3522_bfr_before (
		.din(new_net_3522),
		.dout(new_net_3521)
	);

	bfr new_net_3523_bfr_before (
		.din(new_net_3523),
		.dout(new_net_3522)
	);

	bfr new_net_3524_bfr_before (
		.din(new_net_3524),
		.dout(new_net_3523)
	);

	bfr new_net_3525_bfr_before (
		.din(new_net_3525),
		.dout(new_net_3524)
	);

	bfr new_net_3526_bfr_before (
		.din(new_net_3526),
		.dout(new_net_3525)
	);

	bfr new_net_3527_bfr_before (
		.din(new_net_3527),
		.dout(new_net_3526)
	);

	bfr new_net_3528_bfr_before (
		.din(new_net_3528),
		.dout(new_net_3527)
	);

	bfr new_net_3529_bfr_before (
		.din(new_net_3529),
		.dout(new_net_3528)
	);

	bfr new_net_3530_bfr_before (
		.din(new_net_3530),
		.dout(new_net_3529)
	);

	bfr new_net_3531_bfr_before (
		.din(new_net_3531),
		.dout(new_net_3530)
	);

	bfr new_net_3532_bfr_before (
		.din(new_net_3532),
		.dout(new_net_3531)
	);

	bfr new_net_3533_bfr_before (
		.din(new_net_3533),
		.dout(new_net_3532)
	);

	bfr new_net_3534_bfr_before (
		.din(new_net_3534),
		.dout(new_net_3533)
	);

	bfr new_net_3535_bfr_before (
		.din(new_net_3535),
		.dout(new_net_3534)
	);

	bfr new_net_3536_bfr_before (
		.din(new_net_3536),
		.dout(new_net_3535)
	);

	bfr new_net_3537_bfr_before (
		.din(new_net_3537),
		.dout(new_net_3536)
	);

	bfr new_net_3538_bfr_before (
		.din(new_net_3538),
		.dout(new_net_3537)
	);

	bfr new_net_3539_bfr_before (
		.din(new_net_3539),
		.dout(new_net_3538)
	);

	bfr new_net_3540_bfr_before (
		.din(new_net_3540),
		.dout(new_net_3539)
	);

	bfr new_net_3541_bfr_before (
		.din(new_net_3541),
		.dout(new_net_3540)
	);

	bfr new_net_3542_bfr_before (
		.din(new_net_3542),
		.dout(new_net_3541)
	);

	bfr new_net_3543_bfr_before (
		.din(new_net_3543),
		.dout(new_net_3542)
	);

	bfr new_net_3544_bfr_before (
		.din(new_net_3544),
		.dout(new_net_3543)
	);

	bfr new_net_3545_bfr_before (
		.din(new_net_3545),
		.dout(new_net_3544)
	);

	bfr new_net_3546_bfr_before (
		.din(new_net_3546),
		.dout(new_net_3545)
	);

	bfr new_net_3547_bfr_before (
		.din(new_net_3547),
		.dout(new_net_3546)
	);

	bfr new_net_3548_bfr_before (
		.din(new_net_3548),
		.dout(new_net_3547)
	);

	bfr new_net_3549_bfr_before (
		.din(new_net_3549),
		.dout(new_net_3548)
	);

	bfr new_net_3550_bfr_before (
		.din(new_net_3550),
		.dout(new_net_3549)
	);

	spl3L n_0039__v_fanout (
		.a(n_0039_),
		.b(new_net_815),
		.c(new_net_813),
		.d(new_net_3550)
	);

	bfr new_net_3551_bfr_after (
		.din(n_0354_),
		.dout(new_net_3551)
	);

	bfr new_net_3552_bfr_after (
		.din(new_net_3551),
		.dout(new_net_3552)
	);

	bfr new_net_3553_bfr_before (
		.din(new_net_3553),
		.dout(new_net_2162)
	);

	bfr new_net_3554_bfr_before (
		.din(new_net_3554),
		.dout(new_net_3553)
	);

	bfr new_net_3555_bfr_before (
		.din(new_net_3555),
		.dout(new_net_3554)
	);

	bfr new_net_3556_bfr_before (
		.din(new_net_3556),
		.dout(new_net_3555)
	);

	bfr new_net_3557_bfr_before (
		.din(new_net_3557),
		.dout(new_net_3556)
	);

	bfr new_net_3558_bfr_before (
		.din(new_net_3558),
		.dout(new_net_3557)
	);

	bfr new_net_3559_bfr_before (
		.din(new_net_3559),
		.dout(new_net_3558)
	);

	bfr new_net_3560_bfr_before (
		.din(new_net_3560),
		.dout(new_net_3559)
	);

	bfr new_net_3561_bfr_before (
		.din(new_net_3561),
		.dout(new_net_3560)
	);

	bfr new_net_3562_bfr_before (
		.din(new_net_3562),
		.dout(new_net_3561)
	);

	bfr new_net_3563_bfr_before (
		.din(new_net_3563),
		.dout(new_net_3562)
	);

	bfr new_net_3564_bfr_before (
		.din(new_net_3564),
		.dout(new_net_3563)
	);

	bfr new_net_3565_bfr_before (
		.din(new_net_3565),
		.dout(new_net_3564)
	);

	bfr new_net_3566_bfr_before (
		.din(new_net_3566),
		.dout(new_net_3565)
	);

	spl2 n_0354__v_fanout (
		.a(new_net_3552),
		.b(new_net_1784),
		.c(new_net_3566)
	);

	bfr new_net_3567_bfr_before (
		.din(new_net_3567),
		.dout(new_net_1276)
	);

	bfr new_net_3568_bfr_before (
		.din(new_net_3568),
		.dout(new_net_3567)
	);

	bfr new_net_3569_bfr_before (
		.din(new_net_3569),
		.dout(new_net_3568)
	);

	bfr new_net_3570_bfr_before (
		.din(new_net_3570),
		.dout(new_net_3569)
	);

	bfr new_net_3571_bfr_before (
		.din(new_net_3571),
		.dout(new_net_3570)
	);

	bfr new_net_3572_bfr_before (
		.din(new_net_3572),
		.dout(new_net_3571)
	);

	bfr new_net_3573_bfr_before (
		.din(new_net_3573),
		.dout(new_net_3572)
	);

	bfr new_net_3574_bfr_before (
		.din(new_net_3574),
		.dout(new_net_3573)
	);

	bfr new_net_3575_bfr_before (
		.din(new_net_3575),
		.dout(new_net_3574)
	);

	bfr new_net_3576_bfr_before (
		.din(new_net_3576),
		.dout(new_net_3575)
	);

	bfr new_net_3577_bfr_before (
		.din(new_net_3577),
		.dout(new_net_3576)
	);

	bfr new_net_3578_bfr_before (
		.din(new_net_3578),
		.dout(new_net_3577)
	);

	bfr new_net_3579_bfr_before (
		.din(new_net_3579),
		.dout(new_net_3578)
	);

	bfr new_net_3580_bfr_before (
		.din(new_net_3580),
		.dout(new_net_3579)
	);

	bfr new_net_3581_bfr_before (
		.din(new_net_3581),
		.dout(new_net_3580)
	);

	bfr new_net_3582_bfr_before (
		.din(new_net_3582),
		.dout(new_net_3581)
	);

	spl3L n_1353__v_fanout (
		.a(n_1353_),
		.b(new_net_3582),
		.c(new_net_1274),
		.d(new_net_1275)
	);

	spl2 new_net_2142_v_fanout (
		.a(new_net_2142),
		.b(new_net_2143),
		.c(new_net_1171)
	);

	bfr new_net_3583_bfr_before (
		.din(new_net_3583),
		.dout(new_net_888)
	);

	bfr new_net_3584_bfr_before (
		.din(new_net_3584),
		.dout(new_net_3583)
	);

	bfr new_net_3585_bfr_before (
		.din(new_net_3585),
		.dout(new_net_3584)
	);

	bfr new_net_3586_bfr_before (
		.din(new_net_3586),
		.dout(new_net_3585)
	);

	bfr new_net_3587_bfr_before (
		.din(new_net_3587),
		.dout(new_net_3586)
	);

	bfr new_net_3588_bfr_before (
		.din(new_net_3588),
		.dout(new_net_3587)
	);

	bfr new_net_3589_bfr_before (
		.din(new_net_3589),
		.dout(new_net_3588)
	);

	bfr new_net_3590_bfr_before (
		.din(new_net_3590),
		.dout(new_net_3589)
	);

	bfr new_net_3591_bfr_before (
		.din(new_net_3591),
		.dout(new_net_3590)
	);

	bfr new_net_3592_bfr_before (
		.din(new_net_3592),
		.dout(new_net_3591)
	);

	bfr new_net_3593_bfr_before (
		.din(new_net_3593),
		.dout(new_net_3592)
	);

	bfr new_net_3594_bfr_before (
		.din(new_net_3594),
		.dout(new_net_3593)
	);

	bfr new_net_3595_bfr_before (
		.din(new_net_3595),
		.dout(new_net_3594)
	);

	bfr new_net_3596_bfr_before (
		.din(new_net_3596),
		.dout(new_net_3595)
	);

	bfr new_net_3597_bfr_before (
		.din(new_net_3597),
		.dout(new_net_3596)
	);

	bfr new_net_3598_bfr_before (
		.din(new_net_3598),
		.dout(new_net_3597)
	);

	bfr new_net_3599_bfr_before (
		.din(new_net_3599),
		.dout(new_net_3598)
	);

	bfr new_net_3600_bfr_before (
		.din(new_net_3600),
		.dout(new_net_3599)
	);

	bfr new_net_3601_bfr_before (
		.din(new_net_3601),
		.dout(new_net_3600)
	);

	bfr new_net_3602_bfr_before (
		.din(new_net_3602),
		.dout(new_net_3601)
	);

	bfr new_net_3603_bfr_before (
		.din(new_net_3603),
		.dout(new_net_3602)
	);

	bfr new_net_3604_bfr_before (
		.din(new_net_3604),
		.dout(new_net_3603)
	);

	spl2 n_1317__v_fanout (
		.a(n_1317_),
		.b(new_net_3604),
		.c(new_net_887)
	);

	spl2 n_1221__v_fanout (
		.a(n_1221_),
		.b(new_net_1864),
		.c(new_net_1863)
	);

	spl2 n_0780__v_fanout (
		.a(n_0780_),
		.b(new_net_1383),
		.c(new_net_1382)
	);

	bfr new_net_3605_bfr_before (
		.din(new_net_3605),
		.dout(new_net_2133)
	);

	bfr new_net_3606_bfr_before (
		.din(new_net_3606),
		.dout(new_net_3605)
	);

	bfr new_net_3607_bfr_before (
		.din(new_net_3607),
		.dout(new_net_3606)
	);

	bfr new_net_3608_bfr_before (
		.din(new_net_3608),
		.dout(new_net_3607)
	);

	bfr new_net_3609_bfr_before (
		.din(new_net_3609),
		.dout(new_net_3608)
	);

	bfr new_net_3610_bfr_before (
		.din(new_net_3610),
		.dout(new_net_3609)
	);

	bfr new_net_3611_bfr_before (
		.din(new_net_3611),
		.dout(new_net_3610)
	);

	bfr new_net_3612_bfr_before (
		.din(new_net_3612),
		.dout(new_net_3611)
	);

	bfr new_net_3613_bfr_before (
		.din(new_net_3613),
		.dout(new_net_3612)
	);

	bfr new_net_3614_bfr_before (
		.din(new_net_3614),
		.dout(new_net_3613)
	);

	bfr new_net_3615_bfr_before (
		.din(new_net_3615),
		.dout(new_net_3614)
	);

	bfr new_net_3616_bfr_before (
		.din(new_net_3616),
		.dout(new_net_3615)
	);

	bfr new_net_3617_bfr_before (
		.din(new_net_3617),
		.dout(new_net_3616)
	);

	bfr new_net_3618_bfr_before (
		.din(new_net_3618),
		.dout(new_net_3617)
	);

	bfr new_net_3619_bfr_before (
		.din(new_net_3619),
		.dout(new_net_3618)
	);

	bfr new_net_3620_bfr_before (
		.din(new_net_3620),
		.dout(new_net_3619)
	);

	bfr new_net_3621_bfr_before (
		.din(new_net_3621),
		.dout(new_net_3620)
	);

	bfr new_net_3622_bfr_before (
		.din(new_net_3622),
		.dout(new_net_3621)
	);

	bfr new_net_3623_bfr_before (
		.din(new_net_3623),
		.dout(new_net_3622)
	);

	bfr new_net_3624_bfr_before (
		.din(new_net_3624),
		.dout(new_net_3623)
	);

	bfr new_net_3625_bfr_before (
		.din(new_net_3625),
		.dout(new_net_3624)
	);

	bfr new_net_3626_bfr_before (
		.din(new_net_3626),
		.dout(new_net_3625)
	);

	bfr new_net_3627_bfr_before (
		.din(new_net_3627),
		.dout(new_net_3626)
	);

	bfr new_net_3628_bfr_before (
		.din(new_net_3628),
		.dout(new_net_3627)
	);

	bfr new_net_3629_bfr_before (
		.din(new_net_3629),
		.dout(new_net_3628)
	);

	bfr new_net_3630_bfr_before (
		.din(new_net_3630),
		.dout(new_net_3629)
	);

	bfr new_net_3631_bfr_before (
		.din(new_net_3631),
		.dout(new_net_3630)
	);

	bfr new_net_3632_bfr_before (
		.din(new_net_3632),
		.dout(new_net_3631)
	);

	bfr new_net_3633_bfr_before (
		.din(new_net_3633),
		.dout(new_net_3632)
	);

	bfr new_net_3634_bfr_before (
		.din(new_net_3634),
		.dout(new_net_3633)
	);

	bfr new_net_3635_bfr_before (
		.din(new_net_3635),
		.dout(new_net_3634)
	);

	bfr new_net_3636_bfr_before (
		.din(new_net_3636),
		.dout(new_net_3635)
	);

	bfr new_net_3637_bfr_before (
		.din(new_net_3637),
		.dout(new_net_3636)
	);

	bfr new_net_3638_bfr_before (
		.din(new_net_3638),
		.dout(new_net_3637)
	);

	bfr new_net_3639_bfr_before (
		.din(new_net_3639),
		.dout(new_net_3638)
	);

	bfr new_net_3640_bfr_before (
		.din(new_net_3640),
		.dout(new_net_3639)
	);

	bfr new_net_3641_bfr_before (
		.din(new_net_3641),
		.dout(new_net_3640)
	);

	bfr new_net_3642_bfr_before (
		.din(new_net_3642),
		.dout(new_net_3641)
	);

	bfr new_net_3643_bfr_before (
		.din(new_net_3643),
		.dout(new_net_3642)
	);

	bfr new_net_3644_bfr_before (
		.din(new_net_3644),
		.dout(new_net_3643)
	);

	bfr new_net_3645_bfr_before (
		.din(new_net_3645),
		.dout(new_net_3644)
	);

	bfr new_net_3646_bfr_before (
		.din(new_net_3646),
		.dout(new_net_3645)
	);

	bfr new_net_3647_bfr_before (
		.din(new_net_3647),
		.dout(new_net_3646)
	);

	bfr new_net_3648_bfr_before (
		.din(new_net_3648),
		.dout(new_net_3647)
	);

	spl3L new_net_2132_v_fanout (
		.a(new_net_2132),
		.b(new_net_3648),
		.c(new_net_778),
		.d(new_net_782)
	);

	bfr new_net_3649_bfr_before (
		.din(new_net_3649),
		.dout(new_net_2157)
	);

	bfr new_net_3650_bfr_before (
		.din(new_net_3650),
		.dout(new_net_3649)
	);

	bfr new_net_3651_bfr_before (
		.din(new_net_3651),
		.dout(new_net_3650)
	);

	bfr new_net_3652_bfr_before (
		.din(new_net_3652),
		.dout(new_net_3651)
	);

	bfr new_net_3653_bfr_before (
		.din(new_net_3653),
		.dout(new_net_3652)
	);

	bfr new_net_3654_bfr_before (
		.din(new_net_3654),
		.dout(new_net_3653)
	);

	bfr new_net_3655_bfr_before (
		.din(new_net_3655),
		.dout(new_net_3654)
	);

	bfr new_net_3656_bfr_before (
		.din(new_net_3656),
		.dout(new_net_3655)
	);

	bfr new_net_3657_bfr_before (
		.din(new_net_3657),
		.dout(new_net_3656)
	);

	bfr new_net_3658_bfr_before (
		.din(new_net_3658),
		.dout(new_net_3657)
	);

	bfr new_net_3659_bfr_before (
		.din(new_net_3659),
		.dout(new_net_3658)
	);

	bfr new_net_3660_bfr_before (
		.din(new_net_3660),
		.dout(new_net_3659)
	);

	bfr new_net_3661_bfr_before (
		.din(new_net_3661),
		.dout(new_net_3660)
	);

	bfr new_net_3662_bfr_before (
		.din(new_net_3662),
		.dout(new_net_3661)
	);

	bfr new_net_3663_bfr_before (
		.din(new_net_3663),
		.dout(new_net_3662)
	);

	bfr new_net_3664_bfr_before (
		.din(new_net_3664),
		.dout(new_net_3663)
	);

	bfr new_net_3665_bfr_before (
		.din(new_net_3665),
		.dout(new_net_3664)
	);

	bfr new_net_3666_bfr_before (
		.din(new_net_3666),
		.dout(new_net_3665)
	);

	bfr new_net_3667_bfr_before (
		.din(new_net_3667),
		.dout(new_net_3666)
	);

	bfr new_net_3668_bfr_before (
		.din(new_net_3668),
		.dout(new_net_3667)
	);

	bfr new_net_3669_bfr_before (
		.din(new_net_3669),
		.dout(new_net_3668)
	);

	bfr new_net_3670_bfr_before (
		.din(new_net_3670),
		.dout(new_net_3669)
	);

	bfr new_net_3671_bfr_before (
		.din(new_net_3671),
		.dout(new_net_3670)
	);

	bfr new_net_3672_bfr_before (
		.din(new_net_3672),
		.dout(new_net_3671)
	);

	bfr new_net_3673_bfr_before (
		.din(new_net_3673),
		.dout(new_net_3672)
	);

	bfr new_net_3674_bfr_before (
		.din(new_net_3674),
		.dout(new_net_3673)
	);

	bfr new_net_3675_bfr_before (
		.din(new_net_3675),
		.dout(new_net_3674)
	);

	bfr new_net_3676_bfr_before (
		.din(new_net_3676),
		.dout(new_net_3675)
	);

	bfr new_net_3677_bfr_before (
		.din(new_net_3677),
		.dout(new_net_3676)
	);

	bfr new_net_3678_bfr_before (
		.din(new_net_3678),
		.dout(new_net_3677)
	);

	bfr new_net_3679_bfr_before (
		.din(new_net_3679),
		.dout(new_net_3678)
	);

	bfr new_net_3680_bfr_before (
		.din(new_net_3680),
		.dout(new_net_3679)
	);

	bfr new_net_3681_bfr_before (
		.din(new_net_3681),
		.dout(new_net_3680)
	);

	bfr new_net_3682_bfr_before (
		.din(new_net_3682),
		.dout(new_net_3681)
	);

	bfr new_net_3683_bfr_before (
		.din(new_net_3683),
		.dout(new_net_3682)
	);

	spl2 n_0041__v_fanout (
		.a(n_0041_),
		.b(new_net_3683),
		.c(new_net_1373)
	);

	bfr new_net_3684_bfr_before (
		.din(new_net_3684),
		.dout(new_net_27)
	);

	bfr new_net_3685_bfr_before (
		.din(new_net_3685),
		.dout(new_net_3684)
	);

	bfr new_net_3686_bfr_before (
		.din(new_net_3686),
		.dout(new_net_3685)
	);

	bfr new_net_3687_bfr_before (
		.din(new_net_3687),
		.dout(new_net_3686)
	);

	bfr new_net_3688_bfr_before (
		.din(new_net_3688),
		.dout(new_net_3687)
	);

	bfr new_net_3689_bfr_before (
		.din(new_net_3689),
		.dout(new_net_3688)
	);

	bfr new_net_3690_bfr_before (
		.din(new_net_3690),
		.dout(new_net_3689)
	);

	bfr new_net_3691_bfr_before (
		.din(new_net_3691),
		.dout(new_net_3690)
	);

	bfr new_net_3692_bfr_before (
		.din(new_net_3692),
		.dout(new_net_3691)
	);

	bfr new_net_3693_bfr_before (
		.din(new_net_3693),
		.dout(new_net_3692)
	);

	bfr new_net_3694_bfr_before (
		.din(new_net_3694),
		.dout(new_net_3693)
	);

	bfr new_net_3695_bfr_before (
		.din(new_net_3695),
		.dout(new_net_3694)
	);

	bfr new_net_3696_bfr_before (
		.din(new_net_3696),
		.dout(new_net_3695)
	);

	bfr new_net_3697_bfr_before (
		.din(new_net_3697),
		.dout(new_net_3696)
	);

	bfr new_net_3698_bfr_before (
		.din(new_net_3698),
		.dout(new_net_3697)
	);

	bfr new_net_3699_bfr_before (
		.din(new_net_3699),
		.dout(new_net_3698)
	);

	bfr new_net_3700_bfr_before (
		.din(new_net_3700),
		.dout(new_net_3699)
	);

	bfr new_net_3701_bfr_before (
		.din(new_net_3701),
		.dout(new_net_3700)
	);

	bfr new_net_3702_bfr_before (
		.din(new_net_3702),
		.dout(new_net_3701)
	);

	bfr new_net_3703_bfr_before (
		.din(new_net_3703),
		.dout(new_net_3702)
	);

	bfr new_net_3704_bfr_before (
		.din(new_net_3704),
		.dout(new_net_3703)
	);

	bfr new_net_3705_bfr_before (
		.din(new_net_3705),
		.dout(new_net_3704)
	);

	bfr new_net_3706_bfr_before (
		.din(new_net_3706),
		.dout(new_net_3705)
	);

	bfr new_net_3707_bfr_before (
		.din(new_net_3707),
		.dout(new_net_3706)
	);

	bfr new_net_3708_bfr_before (
		.din(new_net_3708),
		.dout(new_net_3707)
	);

	bfr new_net_3709_bfr_before (
		.din(new_net_3709),
		.dout(new_net_3708)
	);

	bfr new_net_3710_bfr_before (
		.din(new_net_3710),
		.dout(new_net_3709)
	);

	bfr new_net_3711_bfr_before (
		.din(new_net_3711),
		.dout(new_net_3710)
	);

	bfr new_net_3712_bfr_before (
		.din(new_net_3712),
		.dout(new_net_3711)
	);

	spl4L n_0062__v_fanout (
		.a(n_0062_),
		.b(new_net_25),
		.c(new_net_26),
		.d(new_net_3712),
		.e(new_net_24)
	);

	bfr new_net_3713_bfr_after (
		.din(n_1288_),
		.dout(new_net_3713)
	);

	bfr new_net_3714_bfr_after (
		.din(new_net_3713),
		.dout(new_net_3714)
	);

	bfr new_net_3715_bfr_after (
		.din(new_net_3714),
		.dout(new_net_3715)
	);

	spl2 n_1288__v_fanout (
		.a(new_net_3715),
		.b(new_net_1476),
		.c(new_net_1475)
	);

	bfr new_net_3716_bfr_before (
		.din(new_net_3716),
		.dout(new_net_1777)
	);

	bfr new_net_3717_bfr_before (
		.din(new_net_3717),
		.dout(new_net_3716)
	);

	spl2 new_net_2103_v_fanout (
		.a(new_net_2103),
		.b(new_net_3717),
		.c(new_net_1779)
	);

	spl2 new_net_2123_v_fanout (
		.a(new_net_2123),
		.b(new_net_1249),
		.c(new_net_1252)
	);

	spl2 n_0693__v_fanout (
		.a(n_0693_),
		.b(new_net_1339),
		.c(new_net_1338)
	);

	bfr new_net_3718_bfr_after (
		.din(n_0343_),
		.dout(new_net_3718)
	);

	bfr new_net_3719_bfr_before (
		.din(new_net_3719),
		.dout(new_net_2161)
	);

	bfr new_net_3720_bfr_before (
		.din(new_net_3720),
		.dout(new_net_3719)
	);

	bfr new_net_3721_bfr_before (
		.din(new_net_3721),
		.dout(new_net_3720)
	);

	bfr new_net_3722_bfr_before (
		.din(new_net_3722),
		.dout(new_net_3721)
	);

	bfr new_net_3723_bfr_before (
		.din(new_net_3723),
		.dout(new_net_3722)
	);

	bfr new_net_3724_bfr_before (
		.din(new_net_3724),
		.dout(new_net_3723)
	);

	bfr new_net_3725_bfr_before (
		.din(new_net_3725),
		.dout(new_net_3724)
	);

	bfr new_net_3726_bfr_before (
		.din(new_net_3726),
		.dout(new_net_3725)
	);

	bfr new_net_3727_bfr_before (
		.din(new_net_3727),
		.dout(new_net_3726)
	);

	bfr new_net_3728_bfr_before (
		.din(new_net_3728),
		.dout(new_net_3727)
	);

	bfr new_net_3729_bfr_before (
		.din(new_net_3729),
		.dout(new_net_3728)
	);

	bfr new_net_3730_bfr_before (
		.din(new_net_3730),
		.dout(new_net_3729)
	);

	bfr new_net_3731_bfr_before (
		.din(new_net_3731),
		.dout(new_net_3730)
	);

	bfr new_net_3732_bfr_before (
		.din(new_net_3732),
		.dout(new_net_3731)
	);

	bfr new_net_3733_bfr_before (
		.din(new_net_3733),
		.dout(new_net_3732)
	);

	bfr new_net_3734_bfr_before (
		.din(new_net_3734),
		.dout(new_net_3733)
	);

	spl2 n_0343__v_fanout (
		.a(new_net_3718),
		.b(new_net_3734),
		.c(new_net_417)
	);

	bfr new_net_3735_bfr_after (
		.din(n_0390_),
		.dout(new_net_3735)
	);

	bfr new_net_3736_bfr_after (
		.din(new_net_3735),
		.dout(new_net_3736)
	);

	bfr new_net_3737_bfr_after (
		.din(new_net_3736),
		.dout(new_net_3737)
	);

	bfr new_net_3738_bfr_before (
		.din(new_net_3738),
		.dout(new_net_355)
	);

	bfr new_net_3739_bfr_before (
		.din(new_net_3739),
		.dout(new_net_3738)
	);

	bfr new_net_3740_bfr_before (
		.din(new_net_3740),
		.dout(new_net_3739)
	);

	bfr new_net_3741_bfr_before (
		.din(new_net_3741),
		.dout(new_net_3740)
	);

	bfr new_net_3742_bfr_before (
		.din(new_net_3742),
		.dout(new_net_3741)
	);

	bfr new_net_3743_bfr_before (
		.din(new_net_3743),
		.dout(new_net_3742)
	);

	bfr new_net_3744_bfr_before (
		.din(new_net_3744),
		.dout(new_net_3743)
	);

	bfr new_net_3745_bfr_before (
		.din(new_net_3745),
		.dout(new_net_3744)
	);

	bfr new_net_3746_bfr_before (
		.din(new_net_3746),
		.dout(new_net_3745)
	);

	bfr new_net_3747_bfr_before (
		.din(new_net_3747),
		.dout(new_net_3746)
	);

	bfr new_net_3748_bfr_before (
		.din(new_net_3748),
		.dout(new_net_3747)
	);

	bfr new_net_3749_bfr_before (
		.din(new_net_3749),
		.dout(new_net_3748)
	);

	bfr new_net_3750_bfr_before (
		.din(new_net_3750),
		.dout(new_net_3749)
	);

	bfr new_net_3751_bfr_before (
		.din(new_net_3751),
		.dout(new_net_3750)
	);

	bfr new_net_3752_bfr_before (
		.din(new_net_3752),
		.dout(new_net_3751)
	);

	bfr new_net_3753_bfr_before (
		.din(new_net_3753),
		.dout(new_net_3752)
	);

	bfr new_net_3754_bfr_before (
		.din(new_net_3754),
		.dout(new_net_3753)
	);

	bfr new_net_3755_bfr_before (
		.din(new_net_3755),
		.dout(new_net_3754)
	);

	bfr new_net_3756_bfr_before (
		.din(new_net_3756),
		.dout(new_net_3755)
	);

	bfr new_net_3757_bfr_before (
		.din(new_net_3757),
		.dout(new_net_3756)
	);

	bfr new_net_3758_bfr_before (
		.din(new_net_3758),
		.dout(new_net_3757)
	);

	bfr new_net_3759_bfr_before (
		.din(new_net_3759),
		.dout(new_net_3758)
	);

	spl3L n_0390__v_fanout (
		.a(new_net_3737),
		.b(new_net_356),
		.c(new_net_3759),
		.d(new_net_357)
	);

	bfr new_net_3760_bfr_before (
		.din(new_net_3760),
		.dout(new_net_2159)
	);

	bfr new_net_3761_bfr_before (
		.din(new_net_3761),
		.dout(new_net_3760)
	);

	bfr new_net_3762_bfr_before (
		.din(new_net_3762),
		.dout(new_net_3761)
	);

	bfr new_net_3763_bfr_before (
		.din(new_net_3763),
		.dout(new_net_3762)
	);

	bfr new_net_3764_bfr_before (
		.din(new_net_3764),
		.dout(new_net_3763)
	);

	bfr new_net_3765_bfr_before (
		.din(new_net_3765),
		.dout(new_net_3764)
	);

	bfr new_net_3766_bfr_before (
		.din(new_net_3766),
		.dout(new_net_3765)
	);

	bfr new_net_3767_bfr_before (
		.din(new_net_3767),
		.dout(new_net_3766)
	);

	bfr new_net_3768_bfr_before (
		.din(new_net_3768),
		.dout(new_net_3767)
	);

	bfr new_net_3769_bfr_before (
		.din(new_net_3769),
		.dout(new_net_3768)
	);

	bfr new_net_3770_bfr_before (
		.din(new_net_3770),
		.dout(new_net_3769)
	);

	bfr new_net_3771_bfr_before (
		.din(new_net_3771),
		.dout(new_net_3770)
	);

	bfr new_net_3772_bfr_before (
		.din(new_net_3772),
		.dout(new_net_3771)
	);

	bfr new_net_3773_bfr_before (
		.din(new_net_3773),
		.dout(new_net_3772)
	);

	bfr new_net_3774_bfr_before (
		.din(new_net_3774),
		.dout(new_net_3773)
	);

	bfr new_net_3775_bfr_before (
		.din(new_net_3775),
		.dout(new_net_3774)
	);

	bfr new_net_3776_bfr_before (
		.din(new_net_3776),
		.dout(new_net_3775)
	);

	bfr new_net_3777_bfr_before (
		.din(new_net_3777),
		.dout(new_net_3776)
	);

	bfr new_net_3778_bfr_before (
		.din(new_net_3778),
		.dout(new_net_3777)
	);

	bfr new_net_3779_bfr_before (
		.din(new_net_3779),
		.dout(new_net_3778)
	);

	bfr new_net_3780_bfr_before (
		.din(new_net_3780),
		.dout(new_net_3779)
	);

	bfr new_net_3781_bfr_before (
		.din(new_net_3781),
		.dout(new_net_3780)
	);

	bfr new_net_3782_bfr_before (
		.din(new_net_3782),
		.dout(new_net_3781)
	);

	bfr new_net_3783_bfr_before (
		.din(new_net_3783),
		.dout(new_net_3782)
	);

	bfr new_net_3784_bfr_before (
		.din(new_net_3784),
		.dout(new_net_3783)
	);

	bfr new_net_3785_bfr_before (
		.din(new_net_3785),
		.dout(new_net_3784)
	);

	bfr new_net_3786_bfr_before (
		.din(new_net_3786),
		.dout(new_net_3785)
	);

	bfr new_net_3787_bfr_before (
		.din(new_net_3787),
		.dout(new_net_3786)
	);

	bfr new_net_3788_bfr_before (
		.din(new_net_3788),
		.dout(new_net_3787)
	);

	bfr new_net_3789_bfr_before (
		.din(new_net_3789),
		.dout(new_net_3788)
	);

	bfr new_net_3790_bfr_before (
		.din(new_net_3790),
		.dout(new_net_3789)
	);

	spl2 n_0081__v_fanout (
		.a(n_0081_),
		.b(new_net_3790),
		.c(new_net_1702)
	);

	spl2 n_0715__v_fanout (
		.a(n_0715_),
		.b(new_net_1892),
		.c(new_net_1891)
	);

	spl2 n_0451__v_fanout (
		.a(n_0451_),
		.b(new_net_747),
		.c(new_net_746)
	);

	spl2 n_0896__v_fanout (
		.a(n_0896_),
		.b(new_net_1273),
		.c(new_net_1272)
	);

	spl2 n_1173__v_fanout (
		.a(n_1173_),
		.b(new_net_1133),
		.c(new_net_1132)
	);

	bfr new_net_3791_bfr_after (
		.din(n_0969_),
		.dout(new_net_3791)
	);

	bfr new_net_3792_bfr_after (
		.din(new_net_3791),
		.dout(new_net_3792)
	);

	spl2 n_0969__v_fanout (
		.a(new_net_3792),
		.b(new_net_1804),
		.c(new_net_1803)
	);

	bfr new_net_3793_bfr_before (
		.din(new_net_3793),
		.dout(new_net_890)
	);

	bfr new_net_3794_bfr_before (
		.din(new_net_3794),
		.dout(new_net_3793)
	);

	bfr new_net_3795_bfr_before (
		.din(new_net_3795),
		.dout(new_net_3794)
	);

	bfr new_net_3796_bfr_before (
		.din(new_net_3796),
		.dout(new_net_3795)
	);

	bfr new_net_3797_bfr_before (
		.din(new_net_3797),
		.dout(new_net_3796)
	);

	bfr new_net_3798_bfr_before (
		.din(new_net_3798),
		.dout(new_net_3797)
	);

	bfr new_net_3799_bfr_before (
		.din(new_net_3799),
		.dout(new_net_3798)
	);

	bfr new_net_3800_bfr_before (
		.din(new_net_3800),
		.dout(new_net_3799)
	);

	bfr new_net_3801_bfr_before (
		.din(new_net_3801),
		.dout(new_net_3800)
	);

	bfr new_net_3802_bfr_before (
		.din(new_net_3802),
		.dout(new_net_3801)
	);

	bfr new_net_3803_bfr_before (
		.din(new_net_3803),
		.dout(new_net_3802)
	);

	bfr new_net_3804_bfr_before (
		.din(new_net_3804),
		.dout(new_net_3803)
	);

	bfr new_net_3805_bfr_before (
		.din(new_net_3805),
		.dout(new_net_3804)
	);

	bfr new_net_3806_bfr_before (
		.din(new_net_3806),
		.dout(new_net_3805)
	);

	bfr new_net_3807_bfr_before (
		.din(new_net_3807),
		.dout(new_net_3806)
	);

	bfr new_net_3808_bfr_before (
		.din(new_net_3808),
		.dout(new_net_3807)
	);

	bfr new_net_3809_bfr_before (
		.din(new_net_3809),
		.dout(new_net_3808)
	);

	bfr new_net_3810_bfr_before (
		.din(new_net_3810),
		.dout(new_net_3809)
	);

	bfr new_net_3811_bfr_before (
		.din(new_net_3811),
		.dout(new_net_3810)
	);

	bfr new_net_3812_bfr_before (
		.din(new_net_3812),
		.dout(new_net_3811)
	);

	bfr new_net_3813_bfr_before (
		.din(new_net_3813),
		.dout(new_net_3812)
	);

	bfr new_net_3814_bfr_before (
		.din(new_net_3814),
		.dout(new_net_3813)
	);

	bfr new_net_3815_bfr_before (
		.din(new_net_3815),
		.dout(new_net_3814)
	);

	spl4L n_1310__v_fanout (
		.a(n_1310_),
		.b(new_net_891),
		.c(new_net_892),
		.d(new_net_3815),
		.e(new_net_889)
	);

	bfr new_net_3816_bfr_before (
		.din(new_net_3816),
		.dout(new_net_1221)
	);

	bfr new_net_3817_bfr_before (
		.din(new_net_3817),
		.dout(new_net_3816)
	);

	bfr new_net_3818_bfr_before (
		.din(new_net_3818),
		.dout(new_net_3817)
	);

	bfr new_net_3819_bfr_before (
		.din(new_net_3819),
		.dout(new_net_3818)
	);

	bfr new_net_3820_bfr_before (
		.din(new_net_3820),
		.dout(new_net_3819)
	);

	bfr new_net_3821_bfr_before (
		.din(new_net_3821),
		.dout(new_net_3820)
	);

	bfr new_net_3822_bfr_before (
		.din(new_net_3822),
		.dout(new_net_3821)
	);

	bfr new_net_3823_bfr_before (
		.din(new_net_3823),
		.dout(new_net_3822)
	);

	bfr new_net_3824_bfr_before (
		.din(new_net_3824),
		.dout(new_net_3823)
	);

	bfr new_net_3825_bfr_before (
		.din(new_net_3825),
		.dout(new_net_3824)
	);

	bfr new_net_3826_bfr_before (
		.din(new_net_3826),
		.dout(new_net_3825)
	);

	bfr new_net_3827_bfr_before (
		.din(new_net_3827),
		.dout(new_net_3826)
	);

	bfr new_net_3828_bfr_before (
		.din(new_net_3828),
		.dout(new_net_3827)
	);

	bfr new_net_3829_bfr_before (
		.din(new_net_3829),
		.dout(new_net_3828)
	);

	bfr new_net_3830_bfr_before (
		.din(new_net_3830),
		.dout(new_net_3829)
	);

	bfr new_net_3831_bfr_before (
		.din(new_net_3831),
		.dout(new_net_3830)
	);

	bfr new_net_3832_bfr_before (
		.din(new_net_3832),
		.dout(new_net_3831)
	);

	bfr new_net_3833_bfr_before (
		.din(new_net_3833),
		.dout(new_net_3832)
	);

	bfr new_net_3834_bfr_before (
		.din(new_net_3834),
		.dout(new_net_3833)
	);

	bfr new_net_3835_bfr_before (
		.din(new_net_3835),
		.dout(new_net_3834)
	);

	bfr new_net_3836_bfr_before (
		.din(new_net_3836),
		.dout(new_net_3835)
	);

	bfr new_net_3837_bfr_before (
		.din(new_net_3837),
		.dout(new_net_3836)
	);

	bfr new_net_3838_bfr_before (
		.din(new_net_3838),
		.dout(new_net_3837)
	);

	bfr new_net_3839_bfr_before (
		.din(new_net_3839),
		.dout(new_net_3838)
	);

	bfr new_net_3840_bfr_before (
		.din(new_net_3840),
		.dout(new_net_3839)
	);

	bfr new_net_3841_bfr_before (
		.din(new_net_3841),
		.dout(new_net_3840)
	);

	bfr new_net_3842_bfr_before (
		.din(new_net_3842),
		.dout(new_net_3841)
	);

	bfr new_net_3843_bfr_before (
		.din(new_net_3843),
		.dout(new_net_3842)
	);

	bfr new_net_3844_bfr_before (
		.din(new_net_3844),
		.dout(new_net_3843)
	);

	bfr new_net_3845_bfr_before (
		.din(new_net_3845),
		.dout(new_net_3844)
	);

	spl2 n_0055__v_fanout (
		.a(n_0055_),
		.b(new_net_3845),
		.c(new_net_1220)
	);

	bfr new_net_3846_bfr_after (
		.din(n_0866_),
		.dout(new_net_3846)
	);

	bfr new_net_3847_bfr_after (
		.din(new_net_3846),
		.dout(new_net_3847)
	);

	bfr new_net_3848_bfr_after (
		.din(new_net_3847),
		.dout(new_net_3848)
	);

	spl2 n_0866__v_fanout (
		.a(new_net_3848),
		.b(new_net_529),
		.c(new_net_528)
	);

	bfr new_net_3849_bfr_after (
		.din(n_0153_),
		.dout(new_net_3849)
	);

	bfr new_net_3850_bfr_after (
		.din(new_net_3849),
		.dout(new_net_3850)
	);

	bfr new_net_3851_bfr_after (
		.din(new_net_3850),
		.dout(new_net_3851)
	);

	bfr new_net_3852_bfr_after (
		.din(new_net_3851),
		.dout(new_net_3852)
	);

	bfr new_net_3853_bfr_after (
		.din(new_net_3852),
		.dout(new_net_3853)
	);

	bfr new_net_3854_bfr_after (
		.din(new_net_3853),
		.dout(new_net_3854)
	);

	bfr new_net_3855_bfr_after (
		.din(new_net_3854),
		.dout(new_net_3855)
	);

	bfr new_net_3856_bfr_after (
		.din(new_net_3855),
		.dout(new_net_3856)
	);

	bfr new_net_3857_bfr_after (
		.din(new_net_3856),
		.dout(new_net_3857)
	);

	bfr new_net_3858_bfr_after (
		.din(new_net_3857),
		.dout(new_net_3858)
	);

	bfr new_net_3859_bfr_after (
		.din(new_net_3858),
		.dout(new_net_3859)
	);

	bfr new_net_3860_bfr_after (
		.din(new_net_3859),
		.dout(new_net_3860)
	);

	bfr new_net_3861_bfr_after (
		.din(new_net_3860),
		.dout(new_net_3861)
	);

	bfr new_net_3862_bfr_after (
		.din(new_net_3861),
		.dout(new_net_3862)
	);

	bfr new_net_3863_bfr_after (
		.din(new_net_3862),
		.dout(new_net_3863)
	);

	bfr new_net_3864_bfr_after (
		.din(new_net_3863),
		.dout(new_net_3864)
	);

	bfr new_net_3865_bfr_after (
		.din(new_net_3864),
		.dout(new_net_3865)
	);

	bfr new_net_3866_bfr_after (
		.din(new_net_3865),
		.dout(new_net_3866)
	);

	bfr new_net_3867_bfr_after (
		.din(new_net_3866),
		.dout(new_net_3867)
	);

	bfr new_net_3868_bfr_before (
		.din(new_net_3868),
		.dout(new_net_2160)
	);

	spl2 n_0153__v_fanout (
		.a(new_net_3867),
		.b(new_net_3868),
		.c(new_net_1184)
	);

	bfr new_net_3869_bfr_before (
		.din(new_net_3869),
		.dout(new_net_414)
	);

	bfr new_net_3870_bfr_before (
		.din(new_net_3870),
		.dout(new_net_3869)
	);

	bfr new_net_3871_bfr_before (
		.din(new_net_3871),
		.dout(new_net_3870)
	);

	bfr new_net_3872_bfr_before (
		.din(new_net_3872),
		.dout(new_net_3871)
	);

	bfr new_net_3873_bfr_before (
		.din(new_net_3873),
		.dout(new_net_3872)
	);

	bfr new_net_3874_bfr_before (
		.din(new_net_3874),
		.dout(new_net_3873)
	);

	bfr new_net_3875_bfr_before (
		.din(new_net_3875),
		.dout(new_net_3874)
	);

	bfr new_net_3876_bfr_before (
		.din(new_net_3876),
		.dout(new_net_3875)
	);

	bfr new_net_3877_bfr_before (
		.din(new_net_3877),
		.dout(new_net_3876)
	);

	bfr new_net_3878_bfr_before (
		.din(new_net_3878),
		.dout(new_net_3877)
	);

	bfr new_net_3879_bfr_before (
		.din(new_net_3879),
		.dout(new_net_3878)
	);

	bfr new_net_3880_bfr_before (
		.din(new_net_3880),
		.dout(new_net_3879)
	);

	bfr new_net_3881_bfr_before (
		.din(new_net_3881),
		.dout(new_net_3880)
	);

	bfr new_net_3882_bfr_before (
		.din(new_net_3882),
		.dout(new_net_3881)
	);

	bfr new_net_3883_bfr_before (
		.din(new_net_3883),
		.dout(new_net_3882)
	);

	bfr new_net_3884_bfr_before (
		.din(new_net_3884),
		.dout(new_net_3883)
	);

	bfr new_net_3885_bfr_before (
		.din(new_net_3885),
		.dout(new_net_3884)
	);

	bfr new_net_3886_bfr_before (
		.din(new_net_3886),
		.dout(new_net_3885)
	);

	bfr new_net_3887_bfr_before (
		.din(new_net_3887),
		.dout(new_net_3886)
	);

	bfr new_net_3888_bfr_before (
		.din(new_net_3888),
		.dout(new_net_3887)
	);

	bfr new_net_3889_bfr_before (
		.din(new_net_3889),
		.dout(new_net_3888)
	);

	bfr new_net_3890_bfr_before (
		.din(new_net_3890),
		.dout(new_net_3889)
	);

	bfr new_net_3891_bfr_before (
		.din(new_net_3891),
		.dout(new_net_3890)
	);

	bfr new_net_3892_bfr_before (
		.din(new_net_3892),
		.dout(new_net_3891)
	);

	bfr new_net_3893_bfr_before (
		.din(new_net_3893),
		.dout(new_net_3892)
	);

	bfr new_net_3894_bfr_before (
		.din(new_net_3894),
		.dout(new_net_3893)
	);

	bfr new_net_3895_bfr_before (
		.din(new_net_3895),
		.dout(new_net_3894)
	);

	bfr new_net_3896_bfr_before (
		.din(new_net_3896),
		.dout(new_net_3895)
	);

	bfr new_net_3897_bfr_before (
		.din(new_net_3897),
		.dout(new_net_3896)
	);

	bfr new_net_3898_bfr_before (
		.din(new_net_3898),
		.dout(new_net_3897)
	);

	bfr new_net_3899_bfr_before (
		.din(new_net_3899),
		.dout(new_net_3898)
	);

	bfr new_net_3900_bfr_before (
		.din(new_net_3900),
		.dout(new_net_3899)
	);

	bfr new_net_3901_bfr_before (
		.din(new_net_3901),
		.dout(new_net_3900)
	);

	bfr new_net_3902_bfr_before (
		.din(new_net_3902),
		.dout(new_net_3901)
	);

	bfr new_net_3903_bfr_before (
		.din(new_net_3903),
		.dout(new_net_3902)
	);

	bfr new_net_3904_bfr_before (
		.din(new_net_3904),
		.dout(new_net_3903)
	);

	bfr new_net_3905_bfr_before (
		.din(new_net_3905),
		.dout(new_net_3904)
	);

	bfr new_net_3906_bfr_before (
		.din(new_net_3906),
		.dout(new_net_3905)
	);

	bfr new_net_3907_bfr_before (
		.din(new_net_3907),
		.dout(new_net_3906)
	);

	bfr new_net_3908_bfr_before (
		.din(new_net_3908),
		.dout(new_net_3907)
	);

	bfr new_net_3909_bfr_before (
		.din(new_net_3909),
		.dout(new_net_3908)
	);

	spl2 n_0106__v_fanout (
		.a(n_0106_),
		.b(new_net_3909),
		.c(new_net_413)
	);

	bfr new_net_3910_bfr_before (
		.din(new_net_3910),
		.dout(new_net_2126)
	);

	bfr new_net_3911_bfr_before (
		.din(new_net_3911),
		.dout(new_net_3910)
	);

	bfr new_net_3912_bfr_before (
		.din(new_net_3912),
		.dout(new_net_3911)
	);

	bfr new_net_3913_bfr_before (
		.din(new_net_3913),
		.dout(new_net_3912)
	);

	bfr new_net_3914_bfr_before (
		.din(new_net_3914),
		.dout(new_net_3913)
	);

	bfr new_net_3915_bfr_before (
		.din(new_net_3915),
		.dout(new_net_3914)
	);

	bfr new_net_3916_bfr_before (
		.din(new_net_3916),
		.dout(new_net_3915)
	);

	bfr new_net_3917_bfr_before (
		.din(new_net_3917),
		.dout(new_net_3916)
	);

	bfr new_net_3918_bfr_before (
		.din(new_net_3918),
		.dout(new_net_3917)
	);

	bfr new_net_3919_bfr_before (
		.din(new_net_3919),
		.dout(new_net_3918)
	);

	bfr new_net_3920_bfr_before (
		.din(new_net_3920),
		.dout(new_net_3919)
	);

	bfr new_net_3921_bfr_before (
		.din(new_net_3921),
		.dout(new_net_3920)
	);

	bfr new_net_3922_bfr_before (
		.din(new_net_3922),
		.dout(new_net_3921)
	);

	bfr new_net_3923_bfr_before (
		.din(new_net_3923),
		.dout(new_net_3922)
	);

	bfr new_net_3924_bfr_before (
		.din(new_net_3924),
		.dout(new_net_3923)
	);

	bfr new_net_3925_bfr_before (
		.din(new_net_3925),
		.dout(new_net_3924)
	);

	bfr new_net_3926_bfr_before (
		.din(new_net_3926),
		.dout(new_net_3925)
	);

	bfr new_net_3927_bfr_before (
		.din(new_net_3927),
		.dout(new_net_3926)
	);

	bfr new_net_3928_bfr_before (
		.din(new_net_3928),
		.dout(new_net_3927)
	);

	bfr new_net_3929_bfr_before (
		.din(new_net_3929),
		.dout(new_net_3928)
	);

	bfr new_net_3930_bfr_before (
		.din(new_net_3930),
		.dout(new_net_3929)
	);

	bfr new_net_3931_bfr_before (
		.din(new_net_3931),
		.dout(new_net_3930)
	);

	bfr new_net_3932_bfr_before (
		.din(new_net_3932),
		.dout(new_net_3931)
	);

	bfr new_net_3933_bfr_before (
		.din(new_net_3933),
		.dout(new_net_3932)
	);

	bfr new_net_3934_bfr_before (
		.din(new_net_3934),
		.dout(new_net_3933)
	);

	bfr new_net_3935_bfr_before (
		.din(new_net_3935),
		.dout(new_net_3934)
	);

	bfr new_net_3936_bfr_before (
		.din(new_net_3936),
		.dout(new_net_3935)
	);

	bfr new_net_3937_bfr_before (
		.din(new_net_3937),
		.dout(new_net_3936)
	);

	bfr new_net_3938_bfr_before (
		.din(new_net_3938),
		.dout(new_net_3937)
	);

	bfr new_net_3939_bfr_before (
		.din(new_net_3939),
		.dout(new_net_3938)
	);

	bfr new_net_3940_bfr_before (
		.din(new_net_3940),
		.dout(new_net_3939)
	);

	bfr new_net_3941_bfr_before (
		.din(new_net_3941),
		.dout(new_net_3940)
	);

	bfr new_net_3942_bfr_before (
		.din(new_net_3942),
		.dout(new_net_3941)
	);

	bfr new_net_3943_bfr_before (
		.din(new_net_3943),
		.dout(new_net_3942)
	);

	bfr new_net_3944_bfr_before (
		.din(new_net_3944),
		.dout(new_net_3943)
	);

	bfr new_net_3945_bfr_before (
		.din(new_net_3945),
		.dout(new_net_3944)
	);

	bfr new_net_3946_bfr_before (
		.din(new_net_3946),
		.dout(new_net_3945)
	);

	bfr new_net_3947_bfr_before (
		.din(new_net_3947),
		.dout(new_net_3946)
	);

	bfr new_net_3948_bfr_before (
		.din(new_net_3948),
		.dout(new_net_3947)
	);

	bfr new_net_3949_bfr_before (
		.din(new_net_3949),
		.dout(new_net_3948)
	);

	bfr new_net_3950_bfr_before (
		.din(new_net_3950),
		.dout(new_net_3949)
	);

	bfr new_net_3951_bfr_before (
		.din(new_net_3951),
		.dout(new_net_3950)
	);

	spl2 new_net_2125_v_fanout (
		.a(new_net_2125),
		.b(new_net_3951),
		.c(new_net_542)
	);

	bfr new_net_3952_bfr_after (
		.din(n_0172_),
		.dout(new_net_3952)
	);

	bfr new_net_3953_bfr_after (
		.din(new_net_3952),
		.dout(new_net_3953)
	);

	bfr new_net_3954_bfr_after (
		.din(new_net_3953),
		.dout(new_net_3954)
	);

	bfr new_net_3955_bfr_after (
		.din(new_net_3954),
		.dout(new_net_3955)
	);

	bfr new_net_3956_bfr_before (
		.din(new_net_3956),
		.dout(new_net_1421)
	);

	bfr new_net_3957_bfr_before (
		.din(new_net_3957),
		.dout(new_net_3956)
	);

	bfr new_net_3958_bfr_before (
		.din(new_net_3958),
		.dout(new_net_3957)
	);

	bfr new_net_3959_bfr_before (
		.din(new_net_3959),
		.dout(new_net_3958)
	);

	bfr new_net_3960_bfr_before (
		.din(new_net_3960),
		.dout(new_net_3959)
	);

	bfr new_net_3961_bfr_before (
		.din(new_net_3961),
		.dout(new_net_3960)
	);

	bfr new_net_3962_bfr_before (
		.din(new_net_3962),
		.dout(new_net_3961)
	);

	bfr new_net_3963_bfr_before (
		.din(new_net_3963),
		.dout(new_net_3962)
	);

	bfr new_net_3964_bfr_before (
		.din(new_net_3964),
		.dout(new_net_3963)
	);

	bfr new_net_3965_bfr_before (
		.din(new_net_3965),
		.dout(new_net_3964)
	);

	bfr new_net_3966_bfr_before (
		.din(new_net_3966),
		.dout(new_net_3965)
	);

	bfr new_net_3967_bfr_before (
		.din(new_net_3967),
		.dout(new_net_3966)
	);

	bfr new_net_3968_bfr_before (
		.din(new_net_3968),
		.dout(new_net_3967)
	);

	bfr new_net_3969_bfr_before (
		.din(new_net_3969),
		.dout(new_net_3968)
	);

	bfr new_net_3970_bfr_before (
		.din(new_net_3970),
		.dout(new_net_3969)
	);

	bfr new_net_3971_bfr_before (
		.din(new_net_3971),
		.dout(new_net_3970)
	);

	bfr new_net_3972_bfr_before (
		.din(new_net_3972),
		.dout(new_net_3971)
	);

	bfr new_net_3973_bfr_before (
		.din(new_net_3973),
		.dout(new_net_3972)
	);

	bfr new_net_3974_bfr_before (
		.din(new_net_3974),
		.dout(new_net_3973)
	);

	bfr new_net_3975_bfr_before (
		.din(new_net_3975),
		.dout(new_net_3974)
	);

	bfr new_net_3976_bfr_before (
		.din(new_net_3976),
		.dout(new_net_3975)
	);

	bfr new_net_3977_bfr_before (
		.din(new_net_3977),
		.dout(new_net_3976)
	);

	bfr new_net_3978_bfr_before (
		.din(new_net_3978),
		.dout(new_net_3977)
	);

	bfr new_net_3979_bfr_before (
		.din(new_net_3979),
		.dout(new_net_3978)
	);

	bfr new_net_3980_bfr_before (
		.din(new_net_3980),
		.dout(new_net_3979)
	);

	bfr new_net_3981_bfr_before (
		.din(new_net_3981),
		.dout(new_net_3980)
	);

	bfr new_net_3982_bfr_before (
		.din(new_net_3982),
		.dout(new_net_3981)
	);

	bfr new_net_3983_bfr_before (
		.din(new_net_3983),
		.dout(new_net_3982)
	);

	bfr new_net_3984_bfr_before (
		.din(new_net_3984),
		.dout(new_net_3983)
	);

	bfr new_net_3985_bfr_before (
		.din(new_net_3985),
		.dout(new_net_3984)
	);

	bfr new_net_3986_bfr_before (
		.din(new_net_3986),
		.dout(new_net_3985)
	);

	bfr new_net_3987_bfr_before (
		.din(new_net_3987),
		.dout(new_net_3986)
	);

	bfr new_net_3988_bfr_before (
		.din(new_net_3988),
		.dout(new_net_3987)
	);

	bfr new_net_3989_bfr_before (
		.din(new_net_3989),
		.dout(new_net_3988)
	);

	bfr new_net_3990_bfr_before (
		.din(new_net_3990),
		.dout(new_net_3989)
	);

	bfr new_net_3991_bfr_before (
		.din(new_net_3991),
		.dout(new_net_3990)
	);

	bfr new_net_3992_bfr_before (
		.din(new_net_3992),
		.dout(new_net_3991)
	);

	bfr new_net_3993_bfr_before (
		.din(new_net_3993),
		.dout(new_net_3992)
	);

	spl2 n_0172__v_fanout (
		.a(new_net_3955),
		.b(new_net_3993),
		.c(new_net_1420)
	);

	bfr new_net_3994_bfr_before (
		.din(new_net_3994),
		.dout(new_net_603)
	);

	bfr new_net_3995_bfr_before (
		.din(new_net_3995),
		.dout(new_net_3994)
	);

	bfr new_net_3996_bfr_before (
		.din(new_net_3996),
		.dout(new_net_3995)
	);

	bfr new_net_3997_bfr_before (
		.din(new_net_3997),
		.dout(new_net_3996)
	);

	bfr new_net_3998_bfr_before (
		.din(new_net_3998),
		.dout(new_net_3997)
	);

	bfr new_net_3999_bfr_before (
		.din(new_net_3999),
		.dout(new_net_3998)
	);

	bfr new_net_4000_bfr_before (
		.din(new_net_4000),
		.dout(new_net_3999)
	);

	bfr new_net_4001_bfr_before (
		.din(new_net_4001),
		.dout(new_net_4000)
	);

	bfr new_net_4002_bfr_before (
		.din(new_net_4002),
		.dout(new_net_4001)
	);

	bfr new_net_4003_bfr_before (
		.din(new_net_4003),
		.dout(new_net_4002)
	);

	bfr new_net_4004_bfr_before (
		.din(new_net_4004),
		.dout(new_net_4003)
	);

	bfr new_net_4005_bfr_before (
		.din(new_net_4005),
		.dout(new_net_4004)
	);

	bfr new_net_4006_bfr_before (
		.din(new_net_4006),
		.dout(new_net_4005)
	);

	bfr new_net_4007_bfr_before (
		.din(new_net_4007),
		.dout(new_net_4006)
	);

	bfr new_net_4008_bfr_before (
		.din(new_net_4008),
		.dout(new_net_4007)
	);

	bfr new_net_4009_bfr_before (
		.din(new_net_4009),
		.dout(new_net_4008)
	);

	bfr new_net_4010_bfr_before (
		.din(new_net_4010),
		.dout(new_net_4009)
	);

	bfr new_net_4011_bfr_before (
		.din(new_net_4011),
		.dout(new_net_4010)
	);

	bfr new_net_4012_bfr_before (
		.din(new_net_4012),
		.dout(new_net_4011)
	);

	bfr new_net_4013_bfr_before (
		.din(new_net_4013),
		.dout(new_net_4012)
	);

	bfr new_net_4014_bfr_before (
		.din(new_net_4014),
		.dout(new_net_4013)
	);

	bfr new_net_4015_bfr_before (
		.din(new_net_4015),
		.dout(new_net_4014)
	);

	bfr new_net_4016_bfr_before (
		.din(new_net_4016),
		.dout(new_net_4015)
	);

	bfr new_net_4017_bfr_before (
		.din(new_net_4017),
		.dout(new_net_4016)
	);

	bfr new_net_4018_bfr_before (
		.din(new_net_4018),
		.dout(new_net_4017)
	);

	bfr new_net_4019_bfr_before (
		.din(new_net_4019),
		.dout(new_net_4018)
	);

	bfr new_net_4020_bfr_before (
		.din(new_net_4020),
		.dout(new_net_4019)
	);

	bfr new_net_4021_bfr_before (
		.din(new_net_4021),
		.dout(new_net_4020)
	);

	bfr new_net_4022_bfr_before (
		.din(new_net_4022),
		.dout(new_net_4021)
	);

	bfr new_net_4023_bfr_before (
		.din(new_net_4023),
		.dout(new_net_4022)
	);

	bfr new_net_4024_bfr_before (
		.din(new_net_4024),
		.dout(new_net_4023)
	);

	bfr new_net_4025_bfr_before (
		.din(new_net_4025),
		.dout(new_net_4024)
	);

	bfr new_net_4026_bfr_before (
		.din(new_net_4026),
		.dout(new_net_4025)
	);

	bfr new_net_4027_bfr_before (
		.din(new_net_4027),
		.dout(new_net_4026)
	);

	bfr new_net_4028_bfr_before (
		.din(new_net_4028),
		.dout(new_net_4027)
	);

	bfr new_net_4029_bfr_before (
		.din(new_net_4029),
		.dout(new_net_4028)
	);

	bfr new_net_4030_bfr_before (
		.din(new_net_4030),
		.dout(new_net_4029)
	);

	bfr new_net_4031_bfr_before (
		.din(new_net_4031),
		.dout(new_net_4030)
	);

	bfr new_net_4032_bfr_before (
		.din(new_net_4032),
		.dout(new_net_4031)
	);

	bfr new_net_4033_bfr_before (
		.din(new_net_4033),
		.dout(new_net_4032)
	);

	spl3L n_0113__v_fanout (
		.a(n_0113_),
		.b(new_net_604),
		.c(new_net_602),
		.d(new_net_4033)
	);

	bfr new_net_4034_bfr_before (
		.din(new_net_4034),
		.dout(new_net_1543)
	);

	bfr new_net_4035_bfr_before (
		.din(new_net_4035),
		.dout(new_net_4034)
	);

	spl2 new_net_2116_v_fanout (
		.a(new_net_2116),
		.b(new_net_4035),
		.c(new_net_1544)
	);

	bfr new_net_4036_bfr_before (
		.din(new_net_4036),
		.dout(new_net_714)
	);

	bfr new_net_4037_bfr_before (
		.din(new_net_4037),
		.dout(new_net_4036)
	);

	bfr new_net_4038_bfr_before (
		.din(new_net_4038),
		.dout(new_net_4037)
	);

	bfr new_net_4039_bfr_before (
		.din(new_net_4039),
		.dout(new_net_4038)
	);

	bfr new_net_4040_bfr_before (
		.din(new_net_4040),
		.dout(new_net_4039)
	);

	bfr new_net_4041_bfr_before (
		.din(new_net_4041),
		.dout(new_net_4040)
	);

	bfr new_net_4042_bfr_before (
		.din(new_net_4042),
		.dout(new_net_4041)
	);

	bfr new_net_4043_bfr_before (
		.din(new_net_4043),
		.dout(new_net_4042)
	);

	bfr new_net_4044_bfr_before (
		.din(new_net_4044),
		.dout(new_net_4043)
	);

	bfr new_net_4045_bfr_before (
		.din(new_net_4045),
		.dout(new_net_4044)
	);

	bfr new_net_4046_bfr_before (
		.din(new_net_4046),
		.dout(new_net_4045)
	);

	bfr new_net_4047_bfr_before (
		.din(new_net_4047),
		.dout(new_net_4046)
	);

	bfr new_net_4048_bfr_before (
		.din(new_net_4048),
		.dout(new_net_4047)
	);

	bfr new_net_4049_bfr_before (
		.din(new_net_4049),
		.dout(new_net_4048)
	);

	bfr new_net_4050_bfr_before (
		.din(new_net_4050),
		.dout(new_net_4049)
	);

	bfr new_net_4051_bfr_before (
		.din(new_net_4051),
		.dout(new_net_4050)
	);

	bfr new_net_4052_bfr_before (
		.din(new_net_4052),
		.dout(new_net_4051)
	);

	bfr new_net_4053_bfr_before (
		.din(new_net_4053),
		.dout(new_net_4052)
	);

	bfr new_net_4054_bfr_before (
		.din(new_net_4054),
		.dout(new_net_4053)
	);

	bfr new_net_4055_bfr_before (
		.din(new_net_4055),
		.dout(new_net_4054)
	);

	bfr new_net_4056_bfr_before (
		.din(new_net_4056),
		.dout(new_net_4055)
	);

	bfr new_net_4057_bfr_before (
		.din(new_net_4057),
		.dout(new_net_4056)
	);

	bfr new_net_4058_bfr_before (
		.din(new_net_4058),
		.dout(new_net_4057)
	);

	bfr new_net_4059_bfr_before (
		.din(new_net_4059),
		.dout(new_net_4058)
	);

	bfr new_net_4060_bfr_before (
		.din(new_net_4060),
		.dout(new_net_4059)
	);

	bfr new_net_4061_bfr_before (
		.din(new_net_4061),
		.dout(new_net_4060)
	);

	bfr new_net_4062_bfr_before (
		.din(new_net_4062),
		.dout(new_net_4061)
	);

	bfr new_net_4063_bfr_before (
		.din(new_net_4063),
		.dout(new_net_4062)
	);

	bfr new_net_4064_bfr_before (
		.din(new_net_4064),
		.dout(new_net_4063)
	);

	bfr new_net_4065_bfr_before (
		.din(new_net_4065),
		.dout(new_net_4064)
	);

	bfr new_net_4066_bfr_before (
		.din(new_net_4066),
		.dout(new_net_4065)
	);

	bfr new_net_4067_bfr_before (
		.din(new_net_4067),
		.dout(new_net_4066)
	);

	bfr new_net_4068_bfr_before (
		.din(new_net_4068),
		.dout(new_net_4067)
	);

	bfr new_net_4069_bfr_before (
		.din(new_net_4069),
		.dout(new_net_4068)
	);

	spl3L n_0034__v_fanout (
		.a(n_0034_),
		.b(new_net_4069),
		.c(new_net_712),
		.d(new_net_713)
	);

	spl2 n_1146__v_fanout (
		.a(n_1146_),
		.b(new_net_1835),
		.c(new_net_1834)
	);

	bfr new_net_4070_bfr_before (
		.din(new_net_4070),
		.dout(new_net_790)
	);

	bfr new_net_4071_bfr_before (
		.din(new_net_4071),
		.dout(new_net_4070)
	);

	bfr new_net_4072_bfr_before (
		.din(new_net_4072),
		.dout(new_net_4071)
	);

	bfr new_net_4073_bfr_before (
		.din(new_net_4073),
		.dout(new_net_4072)
	);

	bfr new_net_4074_bfr_before (
		.din(new_net_4074),
		.dout(new_net_4073)
	);

	bfr new_net_4075_bfr_before (
		.din(new_net_4075),
		.dout(new_net_4074)
	);

	bfr new_net_4076_bfr_before (
		.din(new_net_4076),
		.dout(new_net_4075)
	);

	bfr new_net_4077_bfr_before (
		.din(new_net_4077),
		.dout(new_net_4076)
	);

	bfr new_net_4078_bfr_before (
		.din(new_net_4078),
		.dout(new_net_4077)
	);

	bfr new_net_4079_bfr_before (
		.din(new_net_4079),
		.dout(new_net_4078)
	);

	bfr new_net_4080_bfr_before (
		.din(new_net_4080),
		.dout(new_net_4079)
	);

	bfr new_net_4081_bfr_before (
		.din(new_net_4081),
		.dout(new_net_4080)
	);

	bfr new_net_4082_bfr_before (
		.din(new_net_4082),
		.dout(new_net_4081)
	);

	bfr new_net_4083_bfr_before (
		.din(new_net_4083),
		.dout(new_net_4082)
	);

	bfr new_net_4084_bfr_before (
		.din(new_net_4084),
		.dout(new_net_4083)
	);

	bfr new_net_4085_bfr_before (
		.din(new_net_4085),
		.dout(new_net_4084)
	);

	bfr new_net_4086_bfr_before (
		.din(new_net_4086),
		.dout(new_net_4085)
	);

	bfr new_net_4087_bfr_before (
		.din(new_net_4087),
		.dout(new_net_4086)
	);

	bfr new_net_4088_bfr_before (
		.din(new_net_4088),
		.dout(new_net_4087)
	);

	bfr new_net_4089_bfr_before (
		.din(new_net_4089),
		.dout(new_net_4088)
	);

	spl3L n_0008__v_fanout (
		.a(n_0008_),
		.b(new_net_4089),
		.c(new_net_788),
		.d(new_net_789)
	);

	bfr new_net_4090_bfr_after (
		.din(n_0767_),
		.dout(new_net_4090)
	);

	bfr new_net_4091_bfr_after (
		.din(new_net_4090),
		.dout(new_net_4091)
	);

	bfr new_net_4092_bfr_after (
		.din(new_net_4091),
		.dout(new_net_4092)
	);

	spl2 n_0767__v_fanout (
		.a(new_net_4092),
		.b(new_net_1117),
		.c(new_net_1116)
	);

	spl2 n_0418__v_fanout (
		.a(n_0418_),
		.b(new_net_1712),
		.c(new_net_1711)
	);

	bfr new_net_4093_bfr_before (
		.din(new_net_4093),
		.dout(new_net_506)
	);

	bfr new_net_4094_bfr_before (
		.din(new_net_4094),
		.dout(new_net_4093)
	);

	bfr new_net_4095_bfr_before (
		.din(new_net_4095),
		.dout(new_net_4094)
	);

	bfr new_net_4096_bfr_before (
		.din(new_net_4096),
		.dout(new_net_4095)
	);

	bfr new_net_4097_bfr_before (
		.din(new_net_4097),
		.dout(new_net_4096)
	);

	bfr new_net_4098_bfr_before (
		.din(new_net_4098),
		.dout(new_net_4097)
	);

	bfr new_net_4099_bfr_before (
		.din(new_net_4099),
		.dout(new_net_4098)
	);

	bfr new_net_4100_bfr_before (
		.din(new_net_4100),
		.dout(new_net_4099)
	);

	bfr new_net_4101_bfr_before (
		.din(new_net_4101),
		.dout(new_net_4100)
	);

	bfr new_net_4102_bfr_before (
		.din(new_net_4102),
		.dout(new_net_4101)
	);

	bfr new_net_4103_bfr_before (
		.din(new_net_4103),
		.dout(new_net_4102)
	);

	bfr new_net_4104_bfr_before (
		.din(new_net_4104),
		.dout(new_net_4103)
	);

	bfr new_net_4105_bfr_before (
		.din(new_net_4105),
		.dout(new_net_4104)
	);

	spl2 new_net_2119_v_fanout (
		.a(new_net_2119),
		.b(new_net_4105),
		.c(new_net_508)
	);

	bfr new_net_4106_bfr_before (
		.din(new_net_4106),
		.dout(new_net_1155)
	);

	bfr new_net_4107_bfr_before (
		.din(new_net_4107),
		.dout(new_net_4106)
	);

	bfr new_net_4108_bfr_before (
		.din(new_net_4108),
		.dout(new_net_4107)
	);

	bfr new_net_4109_bfr_before (
		.din(new_net_4109),
		.dout(new_net_4108)
	);

	bfr new_net_4110_bfr_before (
		.din(new_net_4110),
		.dout(new_net_4109)
	);

	bfr new_net_4111_bfr_before (
		.din(new_net_4111),
		.dout(new_net_4110)
	);

	bfr new_net_4112_bfr_before (
		.din(new_net_4112),
		.dout(new_net_4111)
	);

	bfr new_net_4113_bfr_before (
		.din(new_net_4113),
		.dout(new_net_4112)
	);

	bfr new_net_4114_bfr_before (
		.din(new_net_4114),
		.dout(new_net_4113)
	);

	bfr new_net_4115_bfr_before (
		.din(new_net_4115),
		.dout(new_net_4114)
	);

	bfr new_net_4116_bfr_before (
		.din(new_net_4116),
		.dout(new_net_4115)
	);

	bfr new_net_4117_bfr_before (
		.din(new_net_4117),
		.dout(new_net_4116)
	);

	bfr new_net_4118_bfr_before (
		.din(new_net_4118),
		.dout(new_net_4117)
	);

	bfr new_net_4119_bfr_before (
		.din(new_net_4119),
		.dout(new_net_4118)
	);

	bfr new_net_4120_bfr_before (
		.din(new_net_4120),
		.dout(new_net_4119)
	);

	bfr new_net_4121_bfr_before (
		.din(new_net_4121),
		.dout(new_net_4120)
	);

	bfr new_net_4122_bfr_before (
		.din(new_net_4122),
		.dout(new_net_4121)
	);

	bfr new_net_4123_bfr_before (
		.din(new_net_4123),
		.dout(new_net_4122)
	);

	bfr new_net_4124_bfr_before (
		.din(new_net_4124),
		.dout(new_net_4123)
	);

	bfr new_net_4125_bfr_before (
		.din(new_net_4125),
		.dout(new_net_4124)
	);

	bfr new_net_4126_bfr_before (
		.din(new_net_4126),
		.dout(new_net_4125)
	);

	bfr new_net_4127_bfr_before (
		.din(new_net_4127),
		.dout(new_net_4126)
	);

	bfr new_net_4128_bfr_before (
		.din(new_net_4128),
		.dout(new_net_4127)
	);

	spl2 new_net_2110_v_fanout (
		.a(new_net_2110),
		.b(new_net_4128),
		.c(new_net_1154)
	);

	bfr new_net_4129_bfr_after (
		.din(n_1193_),
		.dout(new_net_4129)
	);

	bfr new_net_4130_bfr_after (
		.din(new_net_4129),
		.dout(new_net_4130)
	);

	bfr new_net_4131_bfr_after (
		.din(new_net_4130),
		.dout(new_net_4131)
	);

	spl2 n_1193__v_fanout (
		.a(new_net_4131),
		.b(new_net_1210),
		.c(new_net_1209)
	);

	spl2 n_1132__v_fanout (
		.a(n_1132_),
		.b(new_net_840),
		.c(new_net_839)
	);

	bfr new_net_4132_bfr_after (
		.din(n_0818_),
		.dout(new_net_4132)
	);

	bfr new_net_4133_bfr_after (
		.din(new_net_4132),
		.dout(new_net_4133)
	);

	bfr new_net_4134_bfr_after (
		.din(new_net_4133),
		.dout(new_net_4134)
	);

	spl2 n_0818__v_fanout (
		.a(new_net_4134),
		.b(new_net_1643),
		.c(new_net_1642)
	);

	spl2 n_0984__v_fanout (
		.a(n_0984_),
		.b(new_net_300),
		.c(new_net_299)
	);

	bfr new_net_4135_bfr_after (
		.din(n_1084_),
		.dout(new_net_4135)
	);

	bfr new_net_4136_bfr_after (
		.din(new_net_4135),
		.dout(new_net_4136)
	);

	bfr new_net_4137_bfr_after (
		.din(new_net_4136),
		.dout(new_net_4137)
	);

	spl2 n_1084__v_fanout (
		.a(new_net_4137),
		.b(new_net_1600),
		.c(new_net_1599)
	);

	spl2 new_net_2120_v_fanout (
		.a(new_net_2120),
		.b(new_net_1867),
		.c(new_net_1866)
	);

	bfr new_net_4138_bfr_before (
		.din(new_net_4138),
		.dout(new_net_2156)
	);

	bfr new_net_4139_bfr_before (
		.din(new_net_4139),
		.dout(new_net_4138)
	);

	bfr new_net_4140_bfr_before (
		.din(new_net_4140),
		.dout(new_net_4139)
	);

	bfr new_net_4141_bfr_before (
		.din(new_net_4141),
		.dout(new_net_4140)
	);

	bfr new_net_4142_bfr_before (
		.din(new_net_4142),
		.dout(new_net_4141)
	);

	bfr new_net_4143_bfr_before (
		.din(new_net_4143),
		.dout(new_net_4142)
	);

	bfr new_net_4144_bfr_before (
		.din(new_net_4144),
		.dout(new_net_4143)
	);

	bfr new_net_4145_bfr_before (
		.din(new_net_4145),
		.dout(new_net_4144)
	);

	bfr new_net_4146_bfr_before (
		.din(new_net_4146),
		.dout(new_net_4145)
	);

	bfr new_net_4147_bfr_before (
		.din(new_net_4147),
		.dout(new_net_4146)
	);

	bfr new_net_4148_bfr_before (
		.din(new_net_4148),
		.dout(new_net_4147)
	);

	bfr new_net_4149_bfr_before (
		.din(new_net_4149),
		.dout(new_net_4148)
	);

	bfr new_net_4150_bfr_before (
		.din(new_net_4150),
		.dout(new_net_4149)
	);

	spl2 n_1370__v_fanout (
		.a(n_1370_),
		.b(new_net_4150),
		.c(new_net_1277)
	);

	spl2 n_1323__v_fanout (
		.a(n_1323_),
		.b(new_net_1533),
		.c(new_net_1532)
	);

	spl3L new_net_2131_v_fanout (
		.a(new_net_2131),
		.b(new_net_780),
		.c(new_net_777),
		.d(new_net_2132)
	);

	bfr new_net_4151_bfr_before (
		.din(new_net_4151),
		.dout(new_net_2154)
	);

	bfr new_net_4152_bfr_before (
		.din(new_net_4152),
		.dout(new_net_4151)
	);

	spl2 new_net_2153_v_fanout (
		.a(new_net_2153),
		.b(new_net_4152),
		.c(new_net_468)
	);

	spl2 n_1099__v_fanout (
		.a(n_1099_),
		.b(new_net_1910),
		.c(new_net_1909)
	);

	bfr new_net_4153_bfr_after (
		.din(n_1060_),
		.dout(new_net_4153)
	);

	bfr new_net_4154_bfr_after (
		.din(new_net_4153),
		.dout(new_net_4154)
	);

	bfr new_net_4155_bfr_after (
		.din(new_net_4154),
		.dout(new_net_4155)
	);

	spl2 n_1060__v_fanout (
		.a(new_net_4155),
		.b(new_net_1377),
		.c(new_net_1376)
	);

	spl2 n_1114__v_fanout (
		.a(n_1114_),
		.b(new_net_1873),
		.c(new_net_1872)
	);

	spl2 n_1027__v_fanout (
		.a(n_1027_),
		.b(new_net_403),
		.c(new_net_402)
	);

	spl2 n_0249__v_fanout (
		.a(n_0249_),
		.b(new_net_817),
		.c(new_net_816)
	);

	bfr new_net_4156_bfr_after (
		.din(n_0139_),
		.dout(new_net_4156)
	);

	bfr new_net_4157_bfr_after (
		.din(new_net_4156),
		.dout(new_net_4157)
	);

	bfr new_net_4158_bfr_after (
		.din(new_net_4157),
		.dout(new_net_4158)
	);

	bfr new_net_4159_bfr_after (
		.din(new_net_4158),
		.dout(new_net_4159)
	);

	bfr new_net_4160_bfr_after (
		.din(new_net_4159),
		.dout(new_net_4160)
	);

	bfr new_net_4161_bfr_after (
		.din(new_net_4160),
		.dout(new_net_4161)
	);

	bfr new_net_4162_bfr_after (
		.din(new_net_4161),
		.dout(new_net_4162)
	);

	bfr new_net_4163_bfr_after (
		.din(new_net_4162),
		.dout(new_net_4163)
	);

	bfr new_net_4164_bfr_after (
		.din(new_net_4163),
		.dout(new_net_4164)
	);

	bfr new_net_4165_bfr_after (
		.din(new_net_4164),
		.dout(new_net_4165)
	);

	bfr new_net_4166_bfr_after (
		.din(new_net_4165),
		.dout(new_net_4166)
	);

	bfr new_net_4167_bfr_after (
		.din(new_net_4166),
		.dout(new_net_4167)
	);

	bfr new_net_4168_bfr_after (
		.din(new_net_4167),
		.dout(new_net_4168)
	);

	bfr new_net_4169_bfr_after (
		.din(new_net_4168),
		.dout(new_net_4169)
	);

	bfr new_net_4170_bfr_after (
		.din(new_net_4169),
		.dout(new_net_4170)
	);

	bfr new_net_4171_bfr_after (
		.din(new_net_4170),
		.dout(new_net_4171)
	);

	bfr new_net_4172_bfr_after (
		.din(new_net_4171),
		.dout(new_net_4172)
	);

	bfr new_net_4173_bfr_after (
		.din(new_net_4172),
		.dout(new_net_4173)
	);

	spl2 n_0139__v_fanout (
		.a(new_net_4173),
		.b(new_net_1157),
		.c(new_net_1156)
	);

	spl2 n_0488__v_fanout (
		.a(n_0488_),
		.b(new_net_537),
		.c(new_net_536)
	);

	bfr new_net_4174_bfr_after (
		.din(n_0079_),
		.dout(new_net_4174)
	);

	bfr new_net_4175_bfr_before (
		.din(new_net_4175),
		.dout(new_net_2155)
	);

	bfr new_net_4176_bfr_before (
		.din(new_net_4176),
		.dout(new_net_4175)
	);

	bfr new_net_4177_bfr_before (
		.din(new_net_4177),
		.dout(new_net_4176)
	);

	bfr new_net_4178_bfr_before (
		.din(new_net_4178),
		.dout(new_net_4177)
	);

	bfr new_net_4179_bfr_before (
		.din(new_net_4179),
		.dout(new_net_4178)
	);

	bfr new_net_4180_bfr_before (
		.din(new_net_4180),
		.dout(new_net_4179)
	);

	bfr new_net_4181_bfr_before (
		.din(new_net_4181),
		.dout(new_net_4180)
	);

	bfr new_net_4182_bfr_before (
		.din(new_net_4182),
		.dout(new_net_4181)
	);

	bfr new_net_4183_bfr_before (
		.din(new_net_4183),
		.dout(new_net_4182)
	);

	bfr new_net_4184_bfr_before (
		.din(new_net_4184),
		.dout(new_net_4183)
	);

	bfr new_net_4185_bfr_before (
		.din(new_net_4185),
		.dout(new_net_4184)
	);

	bfr new_net_4186_bfr_before (
		.din(new_net_4186),
		.dout(new_net_4185)
	);

	bfr new_net_4187_bfr_before (
		.din(new_net_4187),
		.dout(new_net_4186)
	);

	bfr new_net_4188_bfr_before (
		.din(new_net_4188),
		.dout(new_net_4187)
	);

	bfr new_net_4189_bfr_before (
		.din(new_net_4189),
		.dout(new_net_4188)
	);

	bfr new_net_4190_bfr_before (
		.din(new_net_4190),
		.dout(new_net_4189)
	);

	bfr new_net_4191_bfr_before (
		.din(new_net_4191),
		.dout(new_net_4190)
	);

	bfr new_net_4192_bfr_before (
		.din(new_net_4192),
		.dout(new_net_4191)
	);

	bfr new_net_4193_bfr_before (
		.din(new_net_4193),
		.dout(new_net_4192)
	);

	bfr new_net_4194_bfr_before (
		.din(new_net_4194),
		.dout(new_net_4193)
	);

	bfr new_net_4195_bfr_before (
		.din(new_net_4195),
		.dout(new_net_4194)
	);

	bfr new_net_4196_bfr_before (
		.din(new_net_4196),
		.dout(new_net_4195)
	);

	bfr new_net_4197_bfr_before (
		.din(new_net_4197),
		.dout(new_net_4196)
	);

	bfr new_net_4198_bfr_before (
		.din(new_net_4198),
		.dout(new_net_4197)
	);

	bfr new_net_4199_bfr_before (
		.din(new_net_4199),
		.dout(new_net_4198)
	);

	bfr new_net_4200_bfr_before (
		.din(new_net_4200),
		.dout(new_net_4199)
	);

	bfr new_net_4201_bfr_before (
		.din(new_net_4201),
		.dout(new_net_4200)
	);

	bfr new_net_4202_bfr_before (
		.din(new_net_4202),
		.dout(new_net_4201)
	);

	bfr new_net_4203_bfr_before (
		.din(new_net_4203),
		.dout(new_net_4202)
	);

	bfr new_net_4204_bfr_before (
		.din(new_net_4204),
		.dout(new_net_4203)
	);

	bfr new_net_4205_bfr_before (
		.din(new_net_4205),
		.dout(new_net_4204)
	);

	bfr new_net_4206_bfr_before (
		.din(new_net_4206),
		.dout(new_net_4205)
	);

	bfr new_net_4207_bfr_before (
		.din(new_net_4207),
		.dout(new_net_4206)
	);

	spl3L n_0079__v_fanout (
		.a(new_net_4174),
		.b(new_net_1651),
		.c(new_net_4207),
		.d(new_net_1652)
	);

	spl2 n_0999__v_fanout (
		.a(n_0999_),
		.b(new_net_695),
		.c(new_net_694)
	);

	spl2 n_0924__v_fanout (
		.a(n_0924_),
		.b(new_net_683),
		.c(new_net_682)
	);

	spl2 n_0945__v_fanout (
		.a(n_0945_),
		.b(new_net_1305),
		.c(new_net_1304)
	);

	spl2 n_0406__v_fanout (
		.a(n_0406_),
		.b(new_net_1474),
		.c(new_net_1473)
	);

	spl2 n_0298__v_fanout (
		.a(n_0298_),
		.b(new_net_1796),
		.c(new_net_1795)
	);

	spl2 n_0271__v_fanout (
		.a(n_0271_),
		.b(new_net_769),
		.c(new_net_768)
	);

	spl2 n_0054__v_fanout (
		.a(n_0054_),
		.b(new_net_1141),
		.c(new_net_1140)
	);

	bfr new_net_4208_bfr_before (
		.din(new_net_4208),
		.dout(new_net_2148)
	);

	bfr new_net_4209_bfr_before (
		.din(new_net_4209),
		.dout(new_net_4208)
	);

	bfr new_net_4210_bfr_before (
		.din(new_net_4210),
		.dout(new_net_4209)
	);

	bfr new_net_4211_bfr_before (
		.din(new_net_4211),
		.dout(new_net_4210)
	);

	bfr new_net_4212_bfr_before (
		.din(new_net_4212),
		.dout(new_net_4211)
	);

	bfr new_net_4213_bfr_before (
		.din(new_net_4213),
		.dout(new_net_4212)
	);

	bfr new_net_4214_bfr_before (
		.din(new_net_4214),
		.dout(new_net_4213)
	);

	bfr new_net_4215_bfr_before (
		.din(new_net_4215),
		.dout(new_net_4214)
	);

	bfr new_net_4216_bfr_before (
		.din(new_net_4216),
		.dout(new_net_4215)
	);

	bfr new_net_4217_bfr_before (
		.din(new_net_4217),
		.dout(new_net_4216)
	);

	bfr new_net_4218_bfr_before (
		.din(new_net_4218),
		.dout(new_net_4217)
	);

	bfr new_net_4219_bfr_before (
		.din(new_net_4219),
		.dout(new_net_4218)
	);

	bfr new_net_4220_bfr_before (
		.din(new_net_4220),
		.dout(new_net_4219)
	);

	bfr new_net_4221_bfr_before (
		.din(new_net_4221),
		.dout(new_net_4220)
	);

	bfr new_net_4222_bfr_before (
		.din(new_net_4222),
		.dout(new_net_4221)
	);

	bfr new_net_4223_bfr_before (
		.din(new_net_4223),
		.dout(new_net_4222)
	);

	bfr new_net_4224_bfr_before (
		.din(new_net_4224),
		.dout(new_net_4223)
	);

	bfr new_net_4225_bfr_before (
		.din(new_net_4225),
		.dout(new_net_4224)
	);

	bfr new_net_4226_bfr_before (
		.din(new_net_4226),
		.dout(new_net_4225)
	);

	bfr new_net_4227_bfr_before (
		.din(new_net_4227),
		.dout(new_net_4226)
	);

	bfr new_net_4228_bfr_before (
		.din(new_net_4228),
		.dout(new_net_4227)
	);

	bfr new_net_4229_bfr_before (
		.din(new_net_4229),
		.dout(new_net_4228)
	);

	bfr new_net_4230_bfr_before (
		.din(new_net_4230),
		.dout(new_net_4229)
	);

	spl2 n_1316__v_fanout (
		.a(n_1316_),
		.b(new_net_4230),
		.c(new_net_1166)
	);

	bfr new_net_4231_bfr_before (
		.din(new_net_4231),
		.dout(new_net_2124)
	);

	bfr new_net_4232_bfr_before (
		.din(new_net_4232),
		.dout(new_net_4231)
	);

	bfr new_net_4233_bfr_before (
		.din(new_net_4233),
		.dout(new_net_4232)
	);

	bfr new_net_4234_bfr_before (
		.din(new_net_4234),
		.dout(new_net_4233)
	);

	bfr new_net_4235_bfr_before (
		.din(new_net_4235),
		.dout(new_net_4234)
	);

	bfr new_net_4236_bfr_before (
		.din(new_net_4236),
		.dout(new_net_4235)
	);

	bfr new_net_4237_bfr_before (
		.din(new_net_4237),
		.dout(new_net_4236)
	);

	bfr new_net_4238_bfr_before (
		.din(new_net_4238),
		.dout(new_net_4237)
	);

	bfr new_net_4239_bfr_before (
		.din(new_net_4239),
		.dout(new_net_4238)
	);

	bfr new_net_4240_bfr_before (
		.din(new_net_4240),
		.dout(new_net_4239)
	);

	bfr new_net_4241_bfr_before (
		.din(new_net_4241),
		.dout(new_net_4240)
	);

	bfr new_net_4242_bfr_before (
		.din(new_net_4242),
		.dout(new_net_4241)
	);

	bfr new_net_4243_bfr_before (
		.din(new_net_4243),
		.dout(new_net_4242)
	);

	bfr new_net_4244_bfr_before (
		.din(new_net_4244),
		.dout(new_net_4243)
	);

	bfr new_net_4245_bfr_before (
		.din(new_net_4245),
		.dout(new_net_4244)
	);

	bfr new_net_4246_bfr_before (
		.din(new_net_4246),
		.dout(new_net_4245)
	);

	bfr new_net_4247_bfr_before (
		.din(new_net_4247),
		.dout(new_net_4246)
	);

	bfr new_net_4248_bfr_before (
		.din(new_net_4248),
		.dout(new_net_4247)
	);

	bfr new_net_4249_bfr_before (
		.din(new_net_4249),
		.dout(new_net_4248)
	);

	bfr new_net_4250_bfr_before (
		.din(new_net_4250),
		.dout(new_net_4249)
	);

	bfr new_net_4251_bfr_before (
		.din(new_net_4251),
		.dout(new_net_4250)
	);

	bfr new_net_4252_bfr_before (
		.din(new_net_4252),
		.dout(new_net_4251)
	);

	bfr new_net_4253_bfr_before (
		.din(new_net_4253),
		.dout(new_net_4252)
	);

	bfr new_net_4254_bfr_before (
		.din(new_net_4254),
		.dout(new_net_4253)
	);

	bfr new_net_4255_bfr_before (
		.din(new_net_4255),
		.dout(new_net_4254)
	);

	bfr new_net_4256_bfr_before (
		.din(new_net_4256),
		.dout(new_net_4255)
	);

	bfr new_net_4257_bfr_before (
		.din(new_net_4257),
		.dout(new_net_4256)
	);

	bfr new_net_4258_bfr_before (
		.din(new_net_4258),
		.dout(new_net_4257)
	);

	bfr new_net_4259_bfr_before (
		.din(new_net_4259),
		.dout(new_net_4258)
	);

	bfr new_net_4260_bfr_before (
		.din(new_net_4260),
		.dout(new_net_4259)
	);

	bfr new_net_4261_bfr_before (
		.din(new_net_4261),
		.dout(new_net_4260)
	);

	bfr new_net_4262_bfr_before (
		.din(new_net_4262),
		.dout(new_net_4261)
	);

	bfr new_net_4263_bfr_before (
		.din(new_net_4263),
		.dout(new_net_4262)
	);

	bfr new_net_4264_bfr_before (
		.din(new_net_4264),
		.dout(new_net_4263)
	);

	spl3L n_0061__v_fanout (
		.a(n_0061_),
		.b(new_net_1860),
		.c(new_net_1857),
		.d(new_net_4264)
	);

	bfr new_net_4265_bfr_before (
		.din(new_net_4265),
		.dout(new_net_2138)
	);

	bfr new_net_4266_bfr_before (
		.din(new_net_4266),
		.dout(new_net_4265)
	);

	bfr new_net_4267_bfr_before (
		.din(new_net_4267),
		.dout(new_net_4266)
	);

	bfr new_net_4268_bfr_before (
		.din(new_net_4268),
		.dout(new_net_4267)
	);

	spl3L n_0382__v_fanout (
		.a(n_0382_),
		.b(new_net_968),
		.c(new_net_969),
		.d(new_net_4268)
	);

	spl3L n_0000__v_fanout (
		.a(n_0000_),
		.b(new_net_1755),
		.c(new_net_1753),
		.d(new_net_1754)
	);

	spl3L n_0697__v_fanout (
		.a(n_0697_),
		.b(new_net_1763),
		.c(new_net_1762),
		.d(new_net_1764)
	);

	bfr new_net_4269_bfr_after (
		.din(n_1339_),
		.dout(new_net_4269)
	);

	bfr new_net_4270_bfr_after (
		.din(new_net_4269),
		.dout(new_net_4270)
	);

	bfr new_net_4271_bfr_after (
		.din(new_net_4270),
		.dout(new_net_4271)
	);

	bfr new_net_4272_bfr_after (
		.din(new_net_4271),
		.dout(new_net_4272)
	);

	bfr new_net_4273_bfr_after (
		.din(new_net_4272),
		.dout(new_net_4273)
	);

	bfr new_net_4274_bfr_before (
		.din(new_net_4274),
		.dout(new_net_2152)
	);

	bfr new_net_4275_bfr_before (
		.din(new_net_4275),
		.dout(new_net_4274)
	);

	bfr new_net_4276_bfr_before (
		.din(new_net_4276),
		.dout(new_net_4275)
	);

	spl2 n_1339__v_fanout (
		.a(new_net_4273),
		.b(new_net_4276),
		.c(new_net_1422)
	);

	bfr new_net_4277_bfr_before (
		.din(new_net_4277),
		.dout(new_net_2110)
	);

	spl2 new_net_2109_v_fanout (
		.a(new_net_2109),
		.b(new_net_4277),
		.c(new_net_1152)
	);

	bfr new_net_4278_bfr_after (
		.din(n_0676_),
		.dout(new_net_4278)
	);

	bfr new_net_4279_bfr_after (
		.din(new_net_4278),
		.dout(new_net_4279)
	);

	bfr new_net_4280_bfr_after (
		.din(new_net_4279),
		.dout(new_net_4280)
	);

	bfr new_net_4281_bfr_after (
		.din(new_net_4280),
		.dout(new_net_4281)
	);

	bfr new_net_4282_bfr_before (
		.din(new_net_4282),
		.dout(new_net_2141)
	);

	bfr new_net_4283_bfr_before (
		.din(new_net_4283),
		.dout(new_net_4282)
	);

	bfr new_net_4284_bfr_before (
		.din(new_net_4284),
		.dout(new_net_4283)
	);

	bfr new_net_4285_bfr_before (
		.din(new_net_4285),
		.dout(new_net_4284)
	);

	spl3L n_0676__v_fanout (
		.a(new_net_4281),
		.b(new_net_107),
		.c(new_net_4285),
		.d(new_net_105)
	);

	bfr new_net_4286_bfr_before (
		.din(new_net_4286),
		.dout(new_net_2144)
	);

	spl3L n_0692__v_fanout (
		.a(n_0692_),
		.b(new_net_1284),
		.c(new_net_1282),
		.d(new_net_4286)
	);

	bfr new_net_4287_bfr_before (
		.din(new_net_4287),
		.dout(new_net_2140)
	);

	bfr new_net_4288_bfr_before (
		.din(new_net_4288),
		.dout(new_net_4287)
	);

	bfr new_net_4289_bfr_before (
		.din(new_net_4289),
		.dout(new_net_4288)
	);

	bfr new_net_4290_bfr_before (
		.din(new_net_4290),
		.dout(new_net_4289)
	);

	bfr new_net_4291_bfr_before (
		.din(new_net_4291),
		.dout(new_net_4290)
	);

	bfr new_net_4292_bfr_before (
		.din(new_net_4292),
		.dout(new_net_4291)
	);

	bfr new_net_4293_bfr_before (
		.din(new_net_4293),
		.dout(new_net_4292)
	);

	bfr new_net_4294_bfr_before (
		.din(new_net_4294),
		.dout(new_net_4293)
	);

	bfr new_net_4295_bfr_before (
		.din(new_net_4295),
		.dout(new_net_4294)
	);

	bfr new_net_4296_bfr_before (
		.din(new_net_4296),
		.dout(new_net_4295)
	);

	bfr new_net_4297_bfr_before (
		.din(new_net_4297),
		.dout(new_net_4296)
	);

	bfr new_net_4298_bfr_before (
		.din(new_net_4298),
		.dout(new_net_4297)
	);

	bfr new_net_4299_bfr_before (
		.din(new_net_4299),
		.dout(new_net_4298)
	);

	bfr new_net_4300_bfr_before (
		.din(new_net_4300),
		.dout(new_net_4299)
	);

	bfr new_net_4301_bfr_before (
		.din(new_net_4301),
		.dout(new_net_4300)
	);

	bfr new_net_4302_bfr_before (
		.din(new_net_4302),
		.dout(new_net_4301)
	);

	bfr new_net_4303_bfr_before (
		.din(new_net_4303),
		.dout(new_net_4302)
	);

	bfr new_net_4304_bfr_before (
		.din(new_net_4304),
		.dout(new_net_4303)
	);

	bfr new_net_4305_bfr_before (
		.din(new_net_4305),
		.dout(new_net_4304)
	);

	bfr new_net_4306_bfr_before (
		.din(new_net_4306),
		.dout(new_net_4305)
	);

	bfr new_net_4307_bfr_before (
		.din(new_net_4307),
		.dout(new_net_4306)
	);

	bfr new_net_4308_bfr_before (
		.din(new_net_4308),
		.dout(new_net_4307)
	);

	bfr new_net_4309_bfr_before (
		.din(new_net_4309),
		.dout(new_net_4308)
	);

	bfr new_net_4310_bfr_before (
		.din(new_net_4310),
		.dout(new_net_4309)
	);

	bfr new_net_4311_bfr_before (
		.din(new_net_4311),
		.dout(new_net_4310)
	);

	bfr new_net_4312_bfr_before (
		.din(new_net_4312),
		.dout(new_net_4311)
	);

	spl3L n_0385__v_fanout (
		.a(n_0385_),
		.b(new_net_1498),
		.c(new_net_4312),
		.d(new_net_1497)
	);

	bfr new_net_4313_bfr_before (
		.din(new_net_4313),
		.dout(new_net_2137)
	);

	bfr new_net_4314_bfr_before (
		.din(new_net_4314),
		.dout(new_net_4313)
	);

	bfr new_net_4315_bfr_before (
		.din(new_net_4315),
		.dout(new_net_4314)
	);

	bfr new_net_4316_bfr_before (
		.din(new_net_4316),
		.dout(new_net_4315)
	);

	bfr new_net_4317_bfr_before (
		.din(new_net_4317),
		.dout(new_net_4316)
	);

	bfr new_net_4318_bfr_before (
		.din(new_net_4318),
		.dout(new_net_4317)
	);

	bfr new_net_4319_bfr_before (
		.din(new_net_4319),
		.dout(new_net_4318)
	);

	bfr new_net_4320_bfr_before (
		.din(new_net_4320),
		.dout(new_net_4319)
	);

	bfr new_net_4321_bfr_before (
		.din(new_net_4321),
		.dout(new_net_4320)
	);

	bfr new_net_4322_bfr_before (
		.din(new_net_4322),
		.dout(new_net_4321)
	);

	bfr new_net_4323_bfr_before (
		.din(new_net_4323),
		.dout(new_net_4322)
	);

	bfr new_net_4324_bfr_before (
		.din(new_net_4324),
		.dout(new_net_4323)
	);

	bfr new_net_4325_bfr_before (
		.din(new_net_4325),
		.dout(new_net_4324)
	);

	bfr new_net_4326_bfr_before (
		.din(new_net_4326),
		.dout(new_net_4325)
	);

	bfr new_net_4327_bfr_before (
		.din(new_net_4327),
		.dout(new_net_4326)
	);

	bfr new_net_4328_bfr_before (
		.din(new_net_4328),
		.dout(new_net_4327)
	);

	bfr new_net_4329_bfr_before (
		.din(new_net_4329),
		.dout(new_net_4328)
	);

	bfr new_net_4330_bfr_before (
		.din(new_net_4330),
		.dout(new_net_4329)
	);

	bfr new_net_4331_bfr_before (
		.din(new_net_4331),
		.dout(new_net_4330)
	);

	bfr new_net_4332_bfr_before (
		.din(new_net_4332),
		.dout(new_net_4331)
	);

	bfr new_net_4333_bfr_before (
		.din(new_net_4333),
		.dout(new_net_4332)
	);

	bfr new_net_4334_bfr_before (
		.din(new_net_4334),
		.dout(new_net_4333)
	);

	bfr new_net_4335_bfr_before (
		.din(new_net_4335),
		.dout(new_net_4334)
	);

	bfr new_net_4336_bfr_before (
		.din(new_net_4336),
		.dout(new_net_4335)
	);

	bfr new_net_4337_bfr_before (
		.din(new_net_4337),
		.dout(new_net_4336)
	);

	bfr new_net_4338_bfr_before (
		.din(new_net_4338),
		.dout(new_net_4337)
	);

	bfr new_net_4339_bfr_before (
		.din(new_net_4339),
		.dout(new_net_4338)
	);

	bfr new_net_4340_bfr_before (
		.din(new_net_4340),
		.dout(new_net_4339)
	);

	bfr new_net_4341_bfr_before (
		.din(new_net_4341),
		.dout(new_net_4340)
	);

	bfr new_net_4342_bfr_before (
		.din(new_net_4342),
		.dout(new_net_4341)
	);

	bfr new_net_4343_bfr_before (
		.din(new_net_4343),
		.dout(new_net_4342)
	);

	bfr new_net_4344_bfr_before (
		.din(new_net_4344),
		.dout(new_net_4343)
	);

	bfr new_net_4345_bfr_before (
		.din(new_net_4345),
		.dout(new_net_4344)
	);

	bfr new_net_4346_bfr_before (
		.din(new_net_4346),
		.dout(new_net_4345)
	);

	spl2 n_0372__v_fanout (
		.a(n_0372_),
		.b(new_net_1907),
		.c(new_net_4346)
	);

	spl2 n_0033__v_fanout (
		.a(n_0033_),
		.b(new_net_523),
		.c(new_net_522)
	);

	spl2 new_net_2105_v_fanout (
		.a(new_net_2105),
		.b(new_net_1062),
		.c(new_net_1060)
	);

	bfr new_net_4347_bfr_before (
		.din(new_net_4347),
		.dout(new_net_2127)
	);

	bfr new_net_4348_bfr_before (
		.din(new_net_4348),
		.dout(new_net_4347)
	);

	bfr new_net_4349_bfr_before (
		.din(new_net_4349),
		.dout(new_net_4348)
	);

	bfr new_net_4350_bfr_before (
		.din(new_net_4350),
		.dout(new_net_4349)
	);

	bfr new_net_4351_bfr_before (
		.din(new_net_4351),
		.dout(new_net_4350)
	);

	bfr new_net_4352_bfr_before (
		.din(new_net_4352),
		.dout(new_net_4351)
	);

	bfr new_net_4353_bfr_before (
		.din(new_net_4353),
		.dout(new_net_4352)
	);

	bfr new_net_4354_bfr_before (
		.din(new_net_4354),
		.dout(new_net_4353)
	);

	bfr new_net_4355_bfr_before (
		.din(new_net_4355),
		.dout(new_net_4354)
	);

	bfr new_net_4356_bfr_before (
		.din(new_net_4356),
		.dout(new_net_4355)
	);

	bfr new_net_4357_bfr_before (
		.din(new_net_4357),
		.dout(new_net_4356)
	);

	bfr new_net_4358_bfr_before (
		.din(new_net_4358),
		.dout(new_net_4357)
	);

	bfr new_net_4359_bfr_before (
		.din(new_net_4359),
		.dout(new_net_4358)
	);

	bfr new_net_4360_bfr_before (
		.din(new_net_4360),
		.dout(new_net_4359)
	);

	bfr new_net_4361_bfr_before (
		.din(new_net_4361),
		.dout(new_net_4360)
	);

	bfr new_net_4362_bfr_before (
		.din(new_net_4362),
		.dout(new_net_4361)
	);

	bfr new_net_4363_bfr_before (
		.din(new_net_4363),
		.dout(new_net_4362)
	);

	bfr new_net_4364_bfr_before (
		.din(new_net_4364),
		.dout(new_net_4363)
	);

	bfr new_net_4365_bfr_before (
		.din(new_net_4365),
		.dout(new_net_4364)
	);

	bfr new_net_4366_bfr_before (
		.din(new_net_4366),
		.dout(new_net_4365)
	);

	bfr new_net_4367_bfr_before (
		.din(new_net_4367),
		.dout(new_net_4366)
	);

	bfr new_net_4368_bfr_before (
		.din(new_net_4368),
		.dout(new_net_4367)
	);

	bfr new_net_4369_bfr_before (
		.din(new_net_4369),
		.dout(new_net_4368)
	);

	bfr new_net_4370_bfr_before (
		.din(new_net_4370),
		.dout(new_net_4369)
	);

	bfr new_net_4371_bfr_before (
		.din(new_net_4371),
		.dout(new_net_4370)
	);

	bfr new_net_4372_bfr_before (
		.din(new_net_4372),
		.dout(new_net_4371)
	);

	bfr new_net_4373_bfr_before (
		.din(new_net_4373),
		.dout(new_net_4372)
	);

	bfr new_net_4374_bfr_before (
		.din(new_net_4374),
		.dout(new_net_4373)
	);

	bfr new_net_4375_bfr_before (
		.din(new_net_4375),
		.dout(new_net_4374)
	);

	bfr new_net_4376_bfr_before (
		.din(new_net_4376),
		.dout(new_net_4375)
	);

	bfr new_net_4377_bfr_before (
		.din(new_net_4377),
		.dout(new_net_4376)
	);

	bfr new_net_4378_bfr_before (
		.din(new_net_4378),
		.dout(new_net_4377)
	);

	bfr new_net_4379_bfr_before (
		.din(new_net_4379),
		.dout(new_net_4378)
	);

	bfr new_net_4380_bfr_before (
		.din(new_net_4380),
		.dout(new_net_4379)
	);

	bfr new_net_4381_bfr_before (
		.din(new_net_4381),
		.dout(new_net_4380)
	);

	bfr new_net_4382_bfr_before (
		.din(new_net_4382),
		.dout(new_net_4381)
	);

	bfr new_net_4383_bfr_before (
		.din(new_net_4383),
		.dout(new_net_4382)
	);

	bfr new_net_4384_bfr_before (
		.din(new_net_4384),
		.dout(new_net_4383)
	);

	bfr new_net_4385_bfr_before (
		.din(new_net_4385),
		.dout(new_net_4384)
	);

	bfr new_net_4386_bfr_before (
		.din(new_net_4386),
		.dout(new_net_4385)
	);

	bfr new_net_4387_bfr_before (
		.din(new_net_4387),
		.dout(new_net_4386)
	);

	bfr new_net_4388_bfr_before (
		.din(new_net_4388),
		.dout(new_net_4387)
	);

	bfr new_net_4389_bfr_before (
		.din(new_net_4389),
		.dout(new_net_4388)
	);

	bfr new_net_4390_bfr_before (
		.din(new_net_4390),
		.dout(new_net_4389)
	);

	bfr new_net_4391_bfr_before (
		.din(new_net_4391),
		.dout(new_net_4390)
	);

	spl3L n_0112__v_fanout (
		.a(n_0112_),
		.b(new_net_4391),
		.c(new_net_574),
		.d(new_net_577)
	);

	bfr new_net_4392_bfr_before (
		.din(new_net_4392),
		.dout(new_net_2122)
	);

	bfr new_net_4393_bfr_before (
		.din(new_net_4393),
		.dout(new_net_4392)
	);

	bfr new_net_4394_bfr_before (
		.din(new_net_4394),
		.dout(new_net_4393)
	);

	bfr new_net_4395_bfr_before (
		.din(new_net_4395),
		.dout(new_net_4394)
	);

	bfr new_net_4396_bfr_before (
		.din(new_net_4396),
		.dout(new_net_4395)
	);

	bfr new_net_4397_bfr_before (
		.din(new_net_4397),
		.dout(new_net_4396)
	);

	bfr new_net_4398_bfr_before (
		.din(new_net_4398),
		.dout(new_net_4397)
	);

	bfr new_net_4399_bfr_before (
		.din(new_net_4399),
		.dout(new_net_4398)
	);

	bfr new_net_4400_bfr_before (
		.din(new_net_4400),
		.dout(new_net_4399)
	);

	bfr new_net_4401_bfr_before (
		.din(new_net_4401),
		.dout(new_net_4400)
	);

	bfr new_net_4402_bfr_before (
		.din(new_net_4402),
		.dout(new_net_4401)
	);

	bfr new_net_4403_bfr_before (
		.din(new_net_4403),
		.dout(new_net_4402)
	);

	bfr new_net_4404_bfr_before (
		.din(new_net_4404),
		.dout(new_net_4403)
	);

	bfr new_net_4405_bfr_before (
		.din(new_net_4405),
		.dout(new_net_4404)
	);

	bfr new_net_4406_bfr_before (
		.din(new_net_4406),
		.dout(new_net_4405)
	);

	bfr new_net_4407_bfr_before (
		.din(new_net_4407),
		.dout(new_net_4406)
	);

	bfr new_net_4408_bfr_before (
		.din(new_net_4408),
		.dout(new_net_4407)
	);

	bfr new_net_4409_bfr_before (
		.din(new_net_4409),
		.dout(new_net_4408)
	);

	bfr new_net_4410_bfr_before (
		.din(new_net_4410),
		.dout(new_net_4409)
	);

	bfr new_net_4411_bfr_before (
		.din(new_net_4411),
		.dout(new_net_4410)
	);

	bfr new_net_4412_bfr_before (
		.din(new_net_4412),
		.dout(new_net_4411)
	);

	bfr new_net_4413_bfr_before (
		.din(new_net_4413),
		.dout(new_net_4412)
	);

	bfr new_net_4414_bfr_before (
		.din(new_net_4414),
		.dout(new_net_4413)
	);

	bfr new_net_4415_bfr_before (
		.din(new_net_4415),
		.dout(new_net_4414)
	);

	bfr new_net_4416_bfr_before (
		.din(new_net_4416),
		.dout(new_net_4415)
	);

	bfr new_net_4417_bfr_before (
		.din(new_net_4417),
		.dout(new_net_4416)
	);

	bfr new_net_4418_bfr_before (
		.din(new_net_4418),
		.dout(new_net_4417)
	);

	bfr new_net_4419_bfr_before (
		.din(new_net_4419),
		.dout(new_net_4418)
	);

	bfr new_net_4420_bfr_before (
		.din(new_net_4420),
		.dout(new_net_4419)
	);

	bfr new_net_4421_bfr_before (
		.din(new_net_4421),
		.dout(new_net_4420)
	);

	bfr new_net_4422_bfr_before (
		.din(new_net_4422),
		.dout(new_net_4421)
	);

	bfr new_net_4423_bfr_before (
		.din(new_net_4423),
		.dout(new_net_4422)
	);

	bfr new_net_4424_bfr_before (
		.din(new_net_4424),
		.dout(new_net_4423)
	);

	bfr new_net_4425_bfr_before (
		.din(new_net_4425),
		.dout(new_net_4424)
	);

	bfr new_net_4426_bfr_before (
		.din(new_net_4426),
		.dout(new_net_4425)
	);

	bfr new_net_4427_bfr_before (
		.din(new_net_4427),
		.dout(new_net_4426)
	);

	bfr new_net_4428_bfr_before (
		.din(new_net_4428),
		.dout(new_net_4427)
	);

	bfr new_net_4429_bfr_before (
		.din(new_net_4429),
		.dout(new_net_4428)
	);

	bfr new_net_4430_bfr_before (
		.din(new_net_4430),
		.dout(new_net_4429)
	);

	bfr new_net_4431_bfr_before (
		.din(new_net_4431),
		.dout(new_net_4430)
	);

	bfr new_net_4432_bfr_before (
		.din(new_net_4432),
		.dout(new_net_4431)
	);

	spl3L n_0025__v_fanout (
		.a(n_0025_),
		.b(new_net_1483),
		.c(new_net_4432),
		.d(new_net_1484)
	);

	bfr new_net_4433_bfr_before (
		.din(new_net_4433),
		.dout(new_net_2150)
	);

	bfr new_net_4434_bfr_before (
		.din(new_net_4434),
		.dout(new_net_4433)
	);

	spl3L n_1334__v_fanout (
		.a(n_1334_),
		.b(new_net_899),
		.c(new_net_897),
		.d(new_net_4434)
	);

	bfr new_net_4435_bfr_after (
		.din(n_1313_),
		.dout(new_net_4435)
	);

	bfr new_net_4436_bfr_after (
		.din(new_net_4435),
		.dout(new_net_4436)
	);

	spl2 n_1313__v_fanout (
		.a(new_net_4436),
		.b(new_net_447),
		.c(new_net_446)
	);

	bfr new_net_4437_bfr_before (
		.din(new_net_4437),
		.dout(new_net_1139)
	);

	bfr new_net_4438_bfr_before (
		.din(new_net_4438),
		.dout(new_net_4437)
	);

	bfr new_net_4439_bfr_before (
		.din(new_net_4439),
		.dout(new_net_4438)
	);

	bfr new_net_4440_bfr_before (
		.din(new_net_4440),
		.dout(new_net_4439)
	);

	bfr new_net_4441_bfr_before (
		.din(new_net_4441),
		.dout(new_net_4440)
	);

	bfr new_net_4442_bfr_before (
		.din(new_net_4442),
		.dout(new_net_4441)
	);

	bfr new_net_4443_bfr_before (
		.din(new_net_4443),
		.dout(new_net_4442)
	);

	bfr new_net_4444_bfr_before (
		.din(new_net_4444),
		.dout(new_net_4443)
	);

	bfr new_net_4445_bfr_before (
		.din(new_net_4445),
		.dout(new_net_4444)
	);

	bfr new_net_4446_bfr_before (
		.din(new_net_4446),
		.dout(new_net_4445)
	);

	bfr new_net_4447_bfr_before (
		.din(new_net_4447),
		.dout(new_net_4446)
	);

	bfr new_net_4448_bfr_before (
		.din(new_net_4448),
		.dout(new_net_4447)
	);

	bfr new_net_4449_bfr_before (
		.din(new_net_4449),
		.dout(new_net_4448)
	);

	bfr new_net_4450_bfr_before (
		.din(new_net_4450),
		.dout(new_net_4449)
	);

	bfr new_net_4451_bfr_before (
		.din(new_net_4451),
		.dout(new_net_4450)
	);

	bfr new_net_4452_bfr_before (
		.din(new_net_4452),
		.dout(new_net_4451)
	);

	bfr new_net_4453_bfr_before (
		.din(new_net_4453),
		.dout(new_net_4452)
	);

	bfr new_net_4454_bfr_before (
		.din(new_net_4454),
		.dout(new_net_4453)
	);

	bfr new_net_4455_bfr_before (
		.din(new_net_4455),
		.dout(new_net_4454)
	);

	bfr new_net_4456_bfr_before (
		.din(new_net_4456),
		.dout(new_net_4455)
	);

	bfr new_net_4457_bfr_before (
		.din(new_net_4457),
		.dout(new_net_4456)
	);

	bfr new_net_4458_bfr_before (
		.din(new_net_4458),
		.dout(new_net_4457)
	);

	bfr new_net_4459_bfr_before (
		.din(new_net_4459),
		.dout(new_net_4458)
	);

	bfr new_net_4460_bfr_before (
		.din(new_net_4460),
		.dout(new_net_4459)
	);

	bfr new_net_4461_bfr_before (
		.din(new_net_4461),
		.dout(new_net_4460)
	);

	bfr new_net_4462_bfr_before (
		.din(new_net_4462),
		.dout(new_net_4461)
	);

	bfr new_net_4463_bfr_before (
		.din(new_net_4463),
		.dout(new_net_4462)
	);

	spl4L n_1314__v_fanout (
		.a(n_1314_),
		.b(new_net_1138),
		.c(new_net_4463),
		.d(new_net_1137),
		.e(new_net_1136)
	);

	bfr new_net_4464_bfr_before (
		.din(new_net_4464),
		.dout(new_net_2128)
	);

	bfr new_net_4465_bfr_before (
		.din(new_net_4465),
		.dout(new_net_4464)
	);

	bfr new_net_4466_bfr_before (
		.din(new_net_4466),
		.dout(new_net_4465)
	);

	spl4L n_0116__v_fanout (
		.a(n_0116_),
		.b(new_net_674),
		.c(new_net_670),
		.d(new_net_4466),
		.e(new_net_673)
	);

	spl3L n_0063__v_fanout (
		.a(n_0063_),
		.b(new_net_93),
		.c(new_net_91),
		.d(new_net_92)
	);

	bfr new_net_4467_bfr_after (
		.din(n_1303_),
		.dout(new_net_4467)
	);

	bfr new_net_4468_bfr_after (
		.din(new_net_4467),
		.dout(new_net_4468)
	);

	bfr new_net_4469_bfr_before (
		.din(new_net_4469),
		.dout(new_net_1954)
	);

	spl2 n_1303__v_fanout (
		.a(new_net_4468),
		.b(new_net_4469),
		.c(new_net_1953)
	);

	bfr new_net_4470_bfr_before (
		.din(new_net_4470),
		.dout(new_net_786)
	);

	bfr new_net_4471_bfr_before (
		.din(new_net_4471),
		.dout(new_net_4470)
	);

	bfr new_net_4472_bfr_before (
		.din(new_net_4472),
		.dout(new_net_4471)
	);

	bfr new_net_4473_bfr_before (
		.din(new_net_4473),
		.dout(new_net_4472)
	);

	bfr new_net_4474_bfr_before (
		.din(new_net_4474),
		.dout(new_net_4473)
	);

	bfr new_net_4475_bfr_before (
		.din(new_net_4475),
		.dout(new_net_4474)
	);

	bfr new_net_4476_bfr_before (
		.din(new_net_4476),
		.dout(new_net_4475)
	);

	bfr new_net_4477_bfr_before (
		.din(new_net_4477),
		.dout(new_net_4476)
	);

	bfr new_net_4478_bfr_before (
		.din(new_net_4478),
		.dout(new_net_4477)
	);

	bfr new_net_4479_bfr_before (
		.din(new_net_4479),
		.dout(new_net_4478)
	);

	bfr new_net_4480_bfr_before (
		.din(new_net_4480),
		.dout(new_net_4479)
	);

	bfr new_net_4481_bfr_before (
		.din(new_net_4481),
		.dout(new_net_4480)
	);

	bfr new_net_4482_bfr_before (
		.din(new_net_4482),
		.dout(new_net_4481)
	);

	bfr new_net_4483_bfr_before (
		.din(new_net_4483),
		.dout(new_net_4482)
	);

	bfr new_net_4484_bfr_before (
		.din(new_net_4484),
		.dout(new_net_4483)
	);

	bfr new_net_4485_bfr_before (
		.din(new_net_4485),
		.dout(new_net_4484)
	);

	bfr new_net_4486_bfr_before (
		.din(new_net_4486),
		.dout(new_net_4485)
	);

	bfr new_net_4487_bfr_before (
		.din(new_net_4487),
		.dout(new_net_4486)
	);

	bfr new_net_4488_bfr_before (
		.din(new_net_4488),
		.dout(new_net_4487)
	);

	bfr new_net_4489_bfr_before (
		.din(new_net_4489),
		.dout(new_net_4488)
	);

	bfr new_net_4490_bfr_before (
		.din(new_net_4490),
		.dout(new_net_4489)
	);

	bfr new_net_4491_bfr_before (
		.din(new_net_4491),
		.dout(new_net_4490)
	);

	bfr new_net_4492_bfr_before (
		.din(new_net_4492),
		.dout(new_net_4491)
	);

	bfr new_net_4493_bfr_before (
		.din(new_net_4493),
		.dout(new_net_4492)
	);

	bfr new_net_4494_bfr_before (
		.din(new_net_4494),
		.dout(new_net_4493)
	);

	bfr new_net_4495_bfr_before (
		.din(new_net_4495),
		.dout(new_net_4494)
	);

	bfr new_net_4496_bfr_before (
		.din(new_net_4496),
		.dout(new_net_4495)
	);

	bfr new_net_4497_bfr_before (
		.din(new_net_4497),
		.dout(new_net_4496)
	);

	bfr new_net_4498_bfr_before (
		.din(new_net_4498),
		.dout(new_net_4497)
	);

	bfr new_net_4499_bfr_before (
		.din(new_net_4499),
		.dout(new_net_4498)
	);

	bfr new_net_4500_bfr_before (
		.din(new_net_4500),
		.dout(new_net_4499)
	);

	bfr new_net_4501_bfr_before (
		.din(new_net_4501),
		.dout(new_net_4500)
	);

	bfr new_net_4502_bfr_before (
		.din(new_net_4502),
		.dout(new_net_4501)
	);

	bfr new_net_4503_bfr_before (
		.din(new_net_4503),
		.dout(new_net_4502)
	);

	bfr new_net_4504_bfr_before (
		.din(new_net_4504),
		.dout(new_net_4503)
	);

	spl2 new_net_2104_v_fanout (
		.a(new_net_2104),
		.b(new_net_4504),
		.c(new_net_785)
	);

	spl2 n_0105__v_fanout (
		.a(n_0105_),
		.b(new_net_1315),
		.c(new_net_1314)
	);

	spl3L n_0152__v_fanout (
		.a(n_0152_),
		.b(new_net_1113),
		.c(new_net_1111),
		.d(new_net_1112)
	);

	spl2 n_0121__v_fanout (
		.a(n_0121_),
		.b(new_net_2131),
		.c(new_net_781)
	);

	bfr new_net_4505_bfr_before (
		.din(new_net_4505),
		.dout(new_net_2149)
	);

	bfr new_net_4506_bfr_before (
		.din(new_net_4506),
		.dout(new_net_4505)
	);

	bfr new_net_4507_bfr_before (
		.din(new_net_4507),
		.dout(new_net_4506)
	);

	bfr new_net_4508_bfr_before (
		.din(new_net_4508),
		.dout(new_net_4507)
	);

	bfr new_net_4509_bfr_before (
		.din(new_net_4509),
		.dout(new_net_4508)
	);

	bfr new_net_4510_bfr_before (
		.din(new_net_4510),
		.dout(new_net_4509)
	);

	bfr new_net_4511_bfr_before (
		.din(new_net_4511),
		.dout(new_net_4510)
	);

	bfr new_net_4512_bfr_before (
		.din(new_net_4512),
		.dout(new_net_4511)
	);

	bfr new_net_4513_bfr_before (
		.din(new_net_4513),
		.dout(new_net_4512)
	);

	bfr new_net_4514_bfr_before (
		.din(new_net_4514),
		.dout(new_net_4513)
	);

	bfr new_net_4515_bfr_before (
		.din(new_net_4515),
		.dout(new_net_4514)
	);

	bfr new_net_4516_bfr_before (
		.din(new_net_4516),
		.dout(new_net_4515)
	);

	bfr new_net_4517_bfr_before (
		.din(new_net_4517),
		.dout(new_net_4516)
	);

	bfr new_net_4518_bfr_before (
		.din(new_net_4518),
		.dout(new_net_4517)
	);

	bfr new_net_4519_bfr_before (
		.din(new_net_4519),
		.dout(new_net_4518)
	);

	bfr new_net_4520_bfr_before (
		.din(new_net_4520),
		.dout(new_net_4519)
	);

	bfr new_net_4521_bfr_before (
		.din(new_net_4521),
		.dout(new_net_4520)
	);

	bfr new_net_4522_bfr_before (
		.din(new_net_4522),
		.dout(new_net_4521)
	);

	bfr new_net_4523_bfr_before (
		.din(new_net_4523),
		.dout(new_net_4522)
	);

	bfr new_net_4524_bfr_before (
		.din(new_net_4524),
		.dout(new_net_4523)
	);

	bfr new_net_4525_bfr_before (
		.din(new_net_4525),
		.dout(new_net_4524)
	);

	spl3L n_1330__v_fanout (
		.a(n_1330_),
		.b(new_net_4525),
		.c(new_net_456),
		.d(new_net_458)
	);

	bfr new_net_4526_bfr_after (
		.din(n_1358_),
		.dout(new_net_4526)
	);

	bfr new_net_4527_bfr_after (
		.din(new_net_4526),
		.dout(new_net_4527)
	);

	bfr new_net_4528_bfr_after (
		.din(new_net_4527),
		.dout(new_net_4528)
	);

	bfr new_net_4529_bfr_after (
		.din(new_net_4528),
		.dout(new_net_4529)
	);

	bfr new_net_4530_bfr_after (
		.din(new_net_4529),
		.dout(new_net_4530)
	);

	bfr new_net_4531_bfr_after (
		.din(new_net_4530),
		.dout(new_net_4531)
	);

	bfr new_net_4532_bfr_after (
		.din(new_net_4531),
		.dout(new_net_4532)
	);

	bfr new_net_4533_bfr_before (
		.din(new_net_4533),
		.dout(new_net_86)
	);

	bfr new_net_4534_bfr_before (
		.din(new_net_4534),
		.dout(new_net_4533)
	);

	spl2 n_1358__v_fanout (
		.a(new_net_4532),
		.b(new_net_4534),
		.c(new_net_85)
	);

	spl3L n_0064__v_fanout (
		.a(n_0064_),
		.b(new_net_1327),
		.c(new_net_1326),
		.d(new_net_1328)
	);

	bfr new_net_4535_bfr_before (
		.din(new_net_4535),
		.dout(new_net_2147)
	);

	bfr new_net_4536_bfr_before (
		.din(new_net_4536),
		.dout(new_net_4535)
	);

	bfr new_net_4537_bfr_before (
		.din(new_net_4537),
		.dout(new_net_4536)
	);

	bfr new_net_4538_bfr_before (
		.din(new_net_4538),
		.dout(new_net_4537)
	);

	bfr new_net_4539_bfr_before (
		.din(new_net_4539),
		.dout(new_net_4538)
	);

	bfr new_net_4540_bfr_before (
		.din(new_net_4540),
		.dout(new_net_4539)
	);

	bfr new_net_4541_bfr_before (
		.din(new_net_4541),
		.dout(new_net_4540)
	);

	bfr new_net_4542_bfr_before (
		.din(new_net_4542),
		.dout(new_net_4541)
	);

	bfr new_net_4543_bfr_before (
		.din(new_net_4543),
		.dout(new_net_4542)
	);

	bfr new_net_4544_bfr_before (
		.din(new_net_4544),
		.dout(new_net_4543)
	);

	bfr new_net_4545_bfr_before (
		.din(new_net_4545),
		.dout(new_net_4544)
	);

	bfr new_net_4546_bfr_before (
		.din(new_net_4546),
		.dout(new_net_4545)
	);

	bfr new_net_4547_bfr_before (
		.din(new_net_4547),
		.dout(new_net_4546)
	);

	bfr new_net_4548_bfr_before (
		.din(new_net_4548),
		.dout(new_net_4547)
	);

	bfr new_net_4549_bfr_before (
		.din(new_net_4549),
		.dout(new_net_4548)
	);

	bfr new_net_4550_bfr_before (
		.din(new_net_4550),
		.dout(new_net_4549)
	);

	bfr new_net_4551_bfr_before (
		.din(new_net_4551),
		.dout(new_net_4550)
	);

	bfr new_net_4552_bfr_before (
		.din(new_net_4552),
		.dout(new_net_4551)
	);

	bfr new_net_4553_bfr_before (
		.din(new_net_4553),
		.dout(new_net_4552)
	);

	bfr new_net_4554_bfr_before (
		.din(new_net_4554),
		.dout(new_net_4553)
	);

	bfr new_net_4555_bfr_before (
		.din(new_net_4555),
		.dout(new_net_4554)
	);

	bfr new_net_4556_bfr_before (
		.din(new_net_4556),
		.dout(new_net_4555)
	);

	bfr new_net_4557_bfr_before (
		.din(new_net_4557),
		.dout(new_net_4556)
	);

	bfr new_net_4558_bfr_before (
		.din(new_net_4558),
		.dout(new_net_4557)
	);

	bfr new_net_4559_bfr_before (
		.din(new_net_4559),
		.dout(new_net_4558)
	);

	bfr new_net_4560_bfr_before (
		.din(new_net_4560),
		.dout(new_net_4559)
	);

	bfr new_net_4561_bfr_before (
		.din(new_net_4561),
		.dout(new_net_4560)
	);

	bfr new_net_4562_bfr_before (
		.din(new_net_4562),
		.dout(new_net_4561)
	);

	bfr new_net_4563_bfr_before (
		.din(new_net_4563),
		.dout(new_net_4562)
	);

	bfr new_net_4564_bfr_before (
		.din(new_net_4564),
		.dout(new_net_4563)
	);

	spl3L n_1296__v_fanout (
		.a(n_1296_),
		.b(new_net_1637),
		.c(new_net_4564),
		.d(new_net_1635)
	);

	spl2 new_net_2114_v_fanout (
		.a(new_net_2114),
		.b(new_net_1628),
		.c(new_net_1627)
	);

	bfr new_net_4565_bfr_before (
		.din(new_net_4565),
		.dout(new_net_2121)
	);

	bfr new_net_4566_bfr_before (
		.din(new_net_4566),
		.dout(new_net_4565)
	);

	bfr new_net_4567_bfr_before (
		.din(new_net_4567),
		.dout(new_net_4566)
	);

	bfr new_net_4568_bfr_before (
		.din(new_net_4568),
		.dout(new_net_4567)
	);

	bfr new_net_4569_bfr_before (
		.din(new_net_4569),
		.dout(new_net_4568)
	);

	bfr new_net_4570_bfr_before (
		.din(new_net_4570),
		.dout(new_net_4569)
	);

	bfr new_net_4571_bfr_before (
		.din(new_net_4571),
		.dout(new_net_4570)
	);

	bfr new_net_4572_bfr_before (
		.din(new_net_4572),
		.dout(new_net_4571)
	);

	bfr new_net_4573_bfr_before (
		.din(new_net_4573),
		.dout(new_net_4572)
	);

	bfr new_net_4574_bfr_before (
		.din(new_net_4574),
		.dout(new_net_4573)
	);

	bfr new_net_4575_bfr_before (
		.din(new_net_4575),
		.dout(new_net_4574)
	);

	bfr new_net_4576_bfr_before (
		.din(new_net_4576),
		.dout(new_net_4575)
	);

	bfr new_net_4577_bfr_before (
		.din(new_net_4577),
		.dout(new_net_4576)
	);

	bfr new_net_4578_bfr_before (
		.din(new_net_4578),
		.dout(new_net_4577)
	);

	bfr new_net_4579_bfr_before (
		.din(new_net_4579),
		.dout(new_net_4578)
	);

	bfr new_net_4580_bfr_before (
		.din(new_net_4580),
		.dout(new_net_4579)
	);

	bfr new_net_4581_bfr_before (
		.din(new_net_4581),
		.dout(new_net_4580)
	);

	spl3L n_0001__v_fanout (
		.a(n_0001_),
		.b(new_net_4581),
		.c(new_net_1811),
		.d(new_net_1813)
	);

	bfr new_net_4582_bfr_before (
		.din(new_net_4582),
		.dout(new_net_2145)
	);

	bfr new_net_4583_bfr_before (
		.din(new_net_4583),
		.dout(new_net_4582)
	);

	bfr new_net_4584_bfr_before (
		.din(new_net_4584),
		.dout(new_net_4583)
	);

	spl3L n_0707__v_fanout (
		.a(n_0707_),
		.b(new_net_1077),
		.c(new_net_1073),
		.d(new_net_4584)
	);

	spl2 n_1309__v_fanout (
		.a(n_1309_),
		.b(new_net_804),
		.c(new_net_803)
	);

	spl3L n_0038__v_fanout (
		.a(n_0038_),
		.b(new_net_1094),
		.c(new_net_1093),
		.d(new_net_1095)
	);

	spl2 n_1368__v_fanout (
		.a(n_1368_),
		.b(new_net_2153),
		.c(new_net_470)
	);

	bfr new_net_4585_bfr_before (
		.din(new_net_4585),
		.dout(new_net_2142)
	);

	spl3L n_0686__v_fanout (
		.a(n_0686_),
		.b(new_net_1173),
		.c(new_net_1174),
		.d(new_net_4585)
	);

	bfr new_net_4586_bfr_before (
		.din(new_net_4586),
		.dout(new_net_2125)
	);

	spl3L n_0111__v_fanout (
		.a(n_0111_),
		.b(new_net_543),
		.c(new_net_4586),
		.d(new_net_546)
	);

	spl3L n_0667__v_fanout (
		.a(n_0667_),
		.b(new_net_1656),
		.c(new_net_1654),
		.d(new_net_1655)
	);

	bfr new_net_4587_bfr_before (
		.din(new_net_4587),
		.dout(new_net_2136)
	);

	bfr new_net_4588_bfr_before (
		.din(new_net_4588),
		.dout(new_net_4587)
	);

	bfr new_net_4589_bfr_before (
		.din(new_net_4589),
		.dout(new_net_4588)
	);

	bfr new_net_4590_bfr_before (
		.din(new_net_4590),
		.dout(new_net_4589)
	);

	bfr new_net_4591_bfr_before (
		.din(new_net_4591),
		.dout(new_net_4590)
	);

	bfr new_net_4592_bfr_before (
		.din(new_net_4592),
		.dout(new_net_4591)
	);

	bfr new_net_4593_bfr_before (
		.din(new_net_4593),
		.dout(new_net_4592)
	);

	bfr new_net_4594_bfr_before (
		.din(new_net_4594),
		.dout(new_net_4593)
	);

	bfr new_net_4595_bfr_before (
		.din(new_net_4595),
		.dout(new_net_4594)
	);

	bfr new_net_4596_bfr_before (
		.din(new_net_4596),
		.dout(new_net_4595)
	);

	bfr new_net_4597_bfr_before (
		.din(new_net_4597),
		.dout(new_net_4596)
	);

	bfr new_net_4598_bfr_before (
		.din(new_net_4598),
		.dout(new_net_4597)
	);

	bfr new_net_4599_bfr_before (
		.din(new_net_4599),
		.dout(new_net_4598)
	);

	bfr new_net_4600_bfr_before (
		.din(new_net_4600),
		.dout(new_net_4599)
	);

	bfr new_net_4601_bfr_before (
		.din(new_net_4601),
		.dout(new_net_4600)
	);

	bfr new_net_4602_bfr_before (
		.din(new_net_4602),
		.dout(new_net_4601)
	);

	bfr new_net_4603_bfr_before (
		.din(new_net_4603),
		.dout(new_net_4602)
	);

	bfr new_net_4604_bfr_before (
		.din(new_net_4604),
		.dout(new_net_4603)
	);

	bfr new_net_4605_bfr_before (
		.din(new_net_4605),
		.dout(new_net_4604)
	);

	bfr new_net_4606_bfr_before (
		.din(new_net_4606),
		.dout(new_net_4605)
	);

	bfr new_net_4607_bfr_before (
		.din(new_net_4607),
		.dout(new_net_4606)
	);

	bfr new_net_4608_bfr_before (
		.din(new_net_4608),
		.dout(new_net_4607)
	);

	bfr new_net_4609_bfr_before (
		.din(new_net_4609),
		.dout(new_net_4608)
	);

	bfr new_net_4610_bfr_before (
		.din(new_net_4610),
		.dout(new_net_4609)
	);

	bfr new_net_4611_bfr_before (
		.din(new_net_4611),
		.dout(new_net_4610)
	);

	bfr new_net_4612_bfr_before (
		.din(new_net_4612),
		.dout(new_net_4611)
	);

	bfr new_net_4613_bfr_before (
		.din(new_net_4613),
		.dout(new_net_4612)
	);

	bfr new_net_4614_bfr_before (
		.din(new_net_4614),
		.dout(new_net_4613)
	);

	bfr new_net_4615_bfr_before (
		.din(new_net_4615),
		.dout(new_net_4614)
	);

	bfr new_net_4616_bfr_before (
		.din(new_net_4616),
		.dout(new_net_4615)
	);

	bfr new_net_4617_bfr_before (
		.din(new_net_4617),
		.dout(new_net_4616)
	);

	bfr new_net_4618_bfr_before (
		.din(new_net_4618),
		.dout(new_net_4617)
	);

	bfr new_net_4619_bfr_before (
		.din(new_net_4619),
		.dout(new_net_4618)
	);

	bfr new_net_4620_bfr_before (
		.din(new_net_4620),
		.dout(new_net_4619)
	);

	bfr new_net_4621_bfr_before (
		.din(new_net_4621),
		.dout(new_net_4620)
	);

	bfr new_net_4622_bfr_before (
		.din(new_net_4622),
		.dout(new_net_4621)
	);

	bfr new_net_4623_bfr_before (
		.din(new_net_4623),
		.dout(new_net_4622)
	);

	spl3L n_0367__v_fanout (
		.a(n_0367_),
		.b(new_net_1381),
		.c(new_net_4623),
		.d(new_net_1379)
	);

	spl2 n_0710__v_fanout (
		.a(n_0710_),
		.b(new_net_1348),
		.c(new_net_1347)
	);

	bfr new_net_4624_bfr_before (
		.din(new_net_4624),
		.dout(new_net_2134)
	);

	bfr new_net_4625_bfr_before (
		.din(new_net_4625),
		.dout(new_net_4624)
	);

	bfr new_net_4626_bfr_before (
		.din(new_net_4626),
		.dout(new_net_4625)
	);

	spl3L n_0360__v_fanout (
		.a(n_0360_),
		.b(new_net_476),
		.c(new_net_474),
		.d(new_net_4626)
	);

	bfr new_net_4627_bfr_before (
		.din(new_net_4627),
		.dout(new_net_2123)
	);

	spl4L n_0040__v_fanout (
		.a(n_0040_),
		.b(new_net_4627),
		.c(new_net_1251),
		.d(new_net_1250),
		.e(new_net_1248)
	);

	bfr new_net_4628_bfr_after (
		.din(n_1326_),
		.dout(new_net_4628)
	);

	spl2 n_1326__v_fanout (
		.a(new_net_4628),
		.b(new_net_1818),
		.c(new_net_1817)
	);

	bfr new_net_4629_bfr_before (
		.din(new_net_4629),
		.dout(new_net_907)
	);

	bfr new_net_4630_bfr_before (
		.din(new_net_4630),
		.dout(new_net_4629)
	);

	bfr new_net_4631_bfr_before (
		.din(new_net_4631),
		.dout(new_net_4630)
	);

	bfr new_net_4632_bfr_before (
		.din(new_net_4632),
		.dout(new_net_4631)
	);

	bfr new_net_4633_bfr_before (
		.din(new_net_4633),
		.dout(new_net_4632)
	);

	bfr new_net_4634_bfr_before (
		.din(new_net_4634),
		.dout(new_net_4633)
	);

	bfr new_net_4635_bfr_before (
		.din(new_net_4635),
		.dout(new_net_4634)
	);

	bfr new_net_4636_bfr_before (
		.din(new_net_4636),
		.dout(new_net_4635)
	);

	bfr new_net_4637_bfr_before (
		.din(new_net_4637),
		.dout(new_net_4636)
	);

	bfr new_net_4638_bfr_before (
		.din(new_net_4638),
		.dout(new_net_4637)
	);

	bfr new_net_4639_bfr_before (
		.din(new_net_4639),
		.dout(new_net_4638)
	);

	bfr new_net_4640_bfr_before (
		.din(new_net_4640),
		.dout(new_net_4639)
	);

	bfr new_net_4641_bfr_before (
		.din(new_net_4641),
		.dout(new_net_4640)
	);

	bfr new_net_4642_bfr_before (
		.din(new_net_4642),
		.dout(new_net_4641)
	);

	bfr new_net_4643_bfr_before (
		.din(new_net_4643),
		.dout(new_net_4642)
	);

	bfr new_net_4644_bfr_before (
		.din(new_net_4644),
		.dout(new_net_4643)
	);

	bfr new_net_4645_bfr_before (
		.din(new_net_4645),
		.dout(new_net_4644)
	);

	bfr new_net_4646_bfr_before (
		.din(new_net_4646),
		.dout(new_net_4645)
	);

	spl4L new_net_2117_v_fanout (
		.a(new_net_2117),
		.b(new_net_905),
		.c(new_net_4646),
		.d(new_net_904),
		.e(new_net_906)
	);

	bfr new_net_4647_bfr_before (
		.din(new_net_4647),
		.dout(new_net_1242)
	);

	bfr new_net_4648_bfr_before (
		.din(new_net_4648),
		.dout(new_net_4647)
	);

	bfr new_net_4649_bfr_before (
		.din(new_net_4649),
		.dout(new_net_4648)
	);

	bfr new_net_4650_bfr_before (
		.din(new_net_4650),
		.dout(new_net_4649)
	);

	bfr new_net_4651_bfr_before (
		.din(new_net_4651),
		.dout(new_net_4650)
	);

	bfr new_net_4652_bfr_before (
		.din(new_net_4652),
		.dout(new_net_4651)
	);

	bfr new_net_4653_bfr_before (
		.din(new_net_4653),
		.dout(new_net_4652)
	);

	bfr new_net_4654_bfr_before (
		.din(new_net_4654),
		.dout(new_net_4653)
	);

	bfr new_net_4655_bfr_before (
		.din(new_net_4655),
		.dout(new_net_4654)
	);

	bfr new_net_4656_bfr_before (
		.din(new_net_4656),
		.dout(new_net_4655)
	);

	bfr new_net_4657_bfr_before (
		.din(new_net_4657),
		.dout(new_net_4656)
	);

	bfr new_net_4658_bfr_before (
		.din(new_net_4658),
		.dout(new_net_4657)
	);

	bfr new_net_4659_bfr_before (
		.din(new_net_4659),
		.dout(new_net_4658)
	);

	bfr new_net_4660_bfr_before (
		.din(new_net_4660),
		.dout(new_net_4659)
	);

	bfr new_net_4661_bfr_before (
		.din(new_net_4661),
		.dout(new_net_4660)
	);

	bfr new_net_4662_bfr_before (
		.din(new_net_4662),
		.dout(new_net_4661)
	);

	bfr new_net_4663_bfr_before (
		.din(new_net_4663),
		.dout(new_net_4662)
	);

	bfr new_net_4664_bfr_before (
		.din(new_net_4664),
		.dout(new_net_4663)
	);

	bfr new_net_4665_bfr_before (
		.din(new_net_4665),
		.dout(new_net_4664)
	);

	bfr new_net_4666_bfr_before (
		.din(new_net_4666),
		.dout(new_net_4665)
	);

	bfr new_net_4667_bfr_before (
		.din(new_net_4667),
		.dout(new_net_4666)
	);

	bfr new_net_4668_bfr_before (
		.din(new_net_4668),
		.dout(new_net_4667)
	);

	spl4L new_net_2111_v_fanout (
		.a(new_net_2111),
		.b(new_net_4668),
		.c(new_net_1243),
		.d(new_net_1240),
		.e(new_net_1241)
	);

	bfr new_net_4669_bfr_after (
		.din(n_0875_),
		.dout(new_net_4669)
	);

	bfr new_net_4670_bfr_after (
		.din(new_net_4669),
		.dout(new_net_4670)
	);

	bfr new_net_4671_bfr_after (
		.din(new_net_4670),
		.dout(new_net_4671)
	);

	spl2 n_0875__v_fanout (
		.a(new_net_4671),
		.b(new_net_697),
		.c(new_net_696)
	);

	spl2 n_0252__v_fanout (
		.a(n_0252_),
		.b(new_net_867),
		.c(new_net_866)
	);

	bfr new_net_4672_bfr_after (
		.din(n_1251_),
		.dout(new_net_4672)
	);

	bfr new_net_4673_bfr_after (
		.din(new_net_4672),
		.dout(new_net_4673)
	);

	bfr new_net_4674_bfr_after (
		.din(new_net_4673),
		.dout(new_net_4674)
	);

	spl2 n_1251__v_fanout (
		.a(new_net_4674),
		.b(new_net_1645),
		.c(new_net_1644)
	);

	spl2 n_0809__v_fanout (
		.a(n_0809_),
		.b(new_net_707),
		.c(new_net_706)
	);

	bfr new_net_4675_bfr_before (
		.din(new_net_4675),
		.dout(new_net_1419)
	);

	spl2 new_net_2112_v_fanout (
		.a(new_net_2112),
		.b(new_net_4675),
		.c(new_net_1417)
	);

	spl2 n_1129__v_fanout (
		.a(n_1129_),
		.b(new_net_1673),
		.c(new_net_1672)
	);

	spl2 n_1258__v_fanout (
		.a(n_1258_),
		.b(new_net_838),
		.c(new_net_837)
	);

	spl2 n_1218__v_fanout (
		.a(n_1218_),
		.b(new_net_1569),
		.c(new_net_1568)
	);

	spl2 n_0301__v_fanout (
		.a(n_0301_),
		.b(new_net_1924),
		.c(new_net_1923)
	);

	spl2 n_1238__v_fanout (
		.a(n_1238_),
		.b(new_net_74),
		.c(new_net_73)
	);

	spl2 n_1190__v_fanout (
		.a(n_1190_),
		.b(new_net_343),
		.c(new_net_342)
	);

	spl2 n_1139__v_fanout (
		.a(n_1139_),
		.b(new_net_955),
		.c(new_net_954)
	);

	spl2 n_0863__v_fanout (
		.a(n_0863_),
		.b(new_net_1183),
		.c(new_net_1182)
	);

	spl2 n_0267__v_fanout (
		.a(n_0267_),
		.b(new_net_113),
		.c(new_net_112)
	);

	spl2 n_1278__v_fanout (
		.a(n_1278_),
		.b(new_net_1232),
		.c(new_net_1231)
	);

	spl2 n_0777__v_fanout (
		.a(n_0777_),
		.b(new_net_1641),
		.c(new_net_1640)
	);

	spl2 n_1183__v_fanout (
		.a(n_1183_),
		.b(new_net_345),
		.c(new_net_344)
	);

	bfr new_net_4676_bfr_before (
		.din(new_net_4676),
		.dout(new_net_61)
	);

	spl2 n_0223__v_fanout (
		.a(n_0223_),
		.b(new_net_62),
		.c(new_net_4676)
	);

	spl2 n_1285__v_fanout (
		.a(n_1285_),
		.b(new_net_1408),
		.c(new_net_1407)
	);

	spl2 n_1211__v_fanout (
		.a(n_1211_),
		.b(new_net_834),
		.c(new_net_833)
	);

	spl2 n_0294__v_fanout (
		.a(n_0294_),
		.b(new_net_1397),
		.c(new_net_1396)
	);

	spl2 new_net_2113_v_fanout (
		.a(new_net_2113),
		.b(new_net_2114),
		.c(new_net_1629)
	);

	spl2 n_1265__v_fanout (
		.a(n_1265_),
		.b(new_net_993),
		.c(new_net_992)
	);

	bfr new_net_4677_bfr_before (
		.din(new_net_4677),
		.dout(new_net_1810)
	);

	bfr new_net_4678_bfr_before (
		.din(new_net_4678),
		.dout(new_net_4677)
	);

	bfr new_net_4679_bfr_before (
		.din(new_net_4679),
		.dout(new_net_4678)
	);

	spl2 n_0232__v_fanout (
		.a(n_0232_),
		.b(new_net_4679),
		.c(new_net_1809)
	);

	bfr new_net_4680_bfr_after (
		.din(n_1204_),
		.dout(new_net_4680)
	);

	bfr new_net_4681_bfr_after (
		.din(new_net_4680),
		.dout(new_net_4681)
	);

	bfr new_net_4682_bfr_after (
		.din(new_net_4681),
		.dout(new_net_4682)
	);

	spl2 n_1204__v_fanout (
		.a(new_net_4682),
		.b(new_net_1856),
		.c(new_net_1855)
	);

	bfr new_net_4683_bfr_before (
		.din(new_net_4683),
		.dout(new_net_1520)
	);

	spl2 n_0324__v_fanout (
		.a(n_0324_),
		.b(new_net_1521),
		.c(new_net_4683)
	);

	spl2 n_1170__v_fanout (
		.a(n_1170_),
		.b(new_net_830),
		.c(new_net_829)
	);

	spl2 n_0764__v_fanout (
		.a(n_0764_),
		.b(new_net_1052),
		.c(new_net_1051)
	);

	bfr new_net_4684_bfr_after (
		.din(n_0821_),
		.dout(new_net_4684)
	);

	bfr new_net_4685_bfr_after (
		.din(new_net_4684),
		.dout(new_net_4685)
	);

	bfr new_net_4686_bfr_after (
		.din(new_net_4685),
		.dout(new_net_4686)
	);

	spl2 n_0821__v_fanout (
		.a(new_net_4686),
		.b(new_net_16),
		.c(new_net_15)
	);

	bfr new_net_4687_bfr_after (
		.din(n_0725_),
		.dout(new_net_4687)
	);

	bfr new_net_4688_bfr_after (
		.din(new_net_4687),
		.dout(new_net_4688)
	);

	bfr new_net_4689_bfr_after (
		.din(new_net_4688),
		.dout(new_net_4689)
	);

	spl2 n_0725__v_fanout (
		.a(new_net_4689),
		.b(new_net_36),
		.c(new_net_35)
	);

	spl2 n_0884__v_fanout (
		.a(n_0884_),
		.b(new_net_917),
		.c(new_net_916)
	);

	spl2 n_0836__v_fanout (
		.a(n_0836_),
		.b(new_net_1748),
		.c(new_net_1747)
	);

	bfr new_net_4690_bfr_after (
		.din(n_1156_),
		.dout(new_net_4690)
	);

	bfr new_net_4691_bfr_after (
		.din(new_net_4690),
		.dout(new_net_4691)
	);

	bfr new_net_4692_bfr_after (
		.din(new_net_4691),
		.dout(new_net_4692)
	);

	spl2 n_1156__v_fanout (
		.a(new_net_4692),
		.b(new_net_1131),
		.c(new_net_1130)
	);

	spl2 n_0957__v_fanout (
		.a(n_0957_),
		.b(new_net_1589),
		.c(new_net_1588)
	);

	spl2 n_0830__v_fanout (
		.a(n_0830_),
		.b(new_net_1559),
		.c(new_net_1558)
	);

	spl2 n_0755__v_fanout (
		.a(n_0755_),
		.b(new_net_863),
		.c(new_net_862)
	);

	spl2 n_1231__v_fanout (
		.a(n_1231_),
		.b(new_net_55),
		.c(new_net_54)
	);

	bfr new_net_4693_bfr_before (
		.din(new_net_4693),
		.dout(new_net_2119)
	);

	bfr new_net_4694_bfr_before (
		.din(new_net_4694),
		.dout(new_net_4693)
	);

	spl2 new_net_2118_v_fanout (
		.a(new_net_2118),
		.b(new_net_4694),
		.c(new_net_505)
	);

	spl2 n_1163__v_fanout (
		.a(n_1163_),
		.b(new_net_1840),
		.c(new_net_1839)
	);

	spl2 n_0274__v_fanout (
		.a(n_0274_),
		.b(new_net_1325),
		.c(new_net_1324)
	);

	spl2 new_net_2115_v_fanout (
		.a(new_net_2115),
		.b(new_net_1359),
		.c(new_net_1360)
	);

	spl2 n_0854__v_fanout (
		.a(n_0854_),
		.b(new_net_78),
		.c(new_net_77)
	);

	spl2 n_0815__v_fanout (
		.a(n_0815_),
		.b(new_net_1311),
		.c(new_net_1310)
	);

	spl2 n_0732__v_fanout (
		.a(n_0732_),
		.b(new_net_298),
		.c(new_net_297)
	);

	spl2 n_0741__v_fanout (
		.a(n_0741_),
		.b(new_net_550),
		.c(new_net_549)
	);

	spl2 n_0787__v_fanout (
		.a(n_0787_),
		.b(new_net_911),
		.c(new_net_910)
	);

	spl2 n_0893__v_fanout (
		.a(n_0893_),
		.b(new_net_995),
		.c(new_net_994)
	);

	bfr new_net_4695_bfr_before (
		.din(new_net_4695),
		.dout(new_net_2120)
	);

	spl2 n_0078__v_fanout (
		.a(n_0078_),
		.b(new_net_4695),
		.c(new_net_1865)
	);

	bfr new_net_4696_bfr_before (
		.din(new_net_4696),
		.dout(new_net_1684)
	);

	bfr new_net_4697_bfr_before (
		.din(new_net_4697),
		.dout(new_net_4696)
	);

	bfr new_net_4698_bfr_before (
		.din(new_net_4698),
		.dout(new_net_4697)
	);

	bfr new_net_4699_bfr_before (
		.din(new_net_4699),
		.dout(new_net_4698)
	);

	bfr new_net_4700_bfr_before (
		.din(new_net_4700),
		.dout(new_net_4699)
	);

	bfr new_net_4701_bfr_before (
		.din(new_net_4701),
		.dout(new_net_4700)
	);

	bfr new_net_4702_bfr_before (
		.din(new_net_4702),
		.dout(new_net_4701)
	);

	bfr new_net_4703_bfr_before (
		.din(new_net_4703),
		.dout(new_net_4702)
	);

	bfr new_net_4704_bfr_before (
		.din(new_net_4704),
		.dout(new_net_4703)
	);

	bfr new_net_4705_bfr_before (
		.din(new_net_4705),
		.dout(new_net_4704)
	);

	bfr new_net_4706_bfr_before (
		.din(new_net_4706),
		.dout(new_net_4705)
	);

	bfr new_net_4707_bfr_before (
		.din(new_net_4707),
		.dout(new_net_4706)
	);

	bfr new_net_4708_bfr_before (
		.din(new_net_4708),
		.dout(new_net_4707)
	);

	bfr new_net_4709_bfr_before (
		.din(new_net_4709),
		.dout(new_net_4708)
	);

	bfr new_net_4710_bfr_before (
		.din(new_net_4710),
		.dout(new_net_4709)
	);

	bfr new_net_4711_bfr_before (
		.din(new_net_4711),
		.dout(new_net_4710)
	);

	bfr new_net_4712_bfr_before (
		.din(new_net_4712),
		.dout(new_net_4711)
	);

	bfr new_net_4713_bfr_before (
		.din(new_net_4713),
		.dout(new_net_4712)
	);

	bfr new_net_4714_bfr_before (
		.din(new_net_4714),
		.dout(new_net_4713)
	);

	bfr new_net_4715_bfr_before (
		.din(new_net_4715),
		.dout(new_net_4714)
	);

	bfr new_net_4716_bfr_before (
		.din(new_net_4716),
		.dout(new_net_4715)
	);

	bfr new_net_4717_bfr_before (
		.din(new_net_4717),
		.dout(new_net_4716)
	);

	bfr new_net_4718_bfr_before (
		.din(new_net_4718),
		.dout(new_net_4717)
	);

	bfr new_net_4719_bfr_before (
		.din(new_net_4719),
		.dout(new_net_4718)
	);

	bfr new_net_4720_bfr_before (
		.din(new_net_4720),
		.dout(new_net_4719)
	);

	bfr new_net_4721_bfr_before (
		.din(new_net_4721),
		.dout(new_net_4720)
	);

	bfr new_net_4722_bfr_before (
		.din(new_net_4722),
		.dout(new_net_4721)
	);

	bfr new_net_4723_bfr_before (
		.din(new_net_4723),
		.dout(new_net_4722)
	);

	bfr new_net_4724_bfr_before (
		.din(new_net_4724),
		.dout(new_net_4723)
	);

	bfr new_net_4725_bfr_before (
		.din(new_net_4725),
		.dout(new_net_4724)
	);

	spl2 n_1298__v_fanout (
		.a(n_1298_),
		.b(new_net_1685),
		.c(new_net_4725)
	);

	bfr new_net_4726_bfr_before (
		.din(new_net_4726),
		.dout(new_net_2105)
	);

	spl3L n_0666__v_fanout (
		.a(n_0666_),
		.b(new_net_1061),
		.c(new_net_1059),
		.d(new_net_4726)
	);

	spl3L n_1295__v_fanout (
		.a(n_1295_),
		.b(new_net_1110),
		.c(new_net_1108),
		.d(new_net_1109)
	);

	spl2 n_1324__v_fanout (
		.a(n_1324_),
		.b(new_net_2113),
		.c(new_net_1626)
	);

	bfr new_net_4727_bfr_before (
		.din(new_net_4727),
		.dout(new_net_405)
	);

	spl2 n_0302__v_fanout (
		.a(n_0302_),
		.b(new_net_4727),
		.c(new_net_404)
	);

	bfr new_net_4728_bfr_before (
		.din(new_net_4728),
		.dout(new_net_831)
	);

	bfr new_net_4729_bfr_before (
		.din(new_net_4729),
		.dout(new_net_4728)
	);

	bfr new_net_4730_bfr_before (
		.din(new_net_4730),
		.dout(new_net_4729)
	);

	bfr new_net_4731_bfr_before (
		.din(new_net_4731),
		.dout(new_net_4730)
	);

	spl2 n_0051__v_fanout (
		.a(n_0051_),
		.b(new_net_832),
		.c(new_net_4731)
	);

	bfr new_net_4732_bfr_before (
		.din(new_net_4732),
		.dout(new_net_1904)
	);

	bfr new_net_4733_bfr_before (
		.din(new_net_4733),
		.dout(new_net_4732)
	);

	bfr new_net_4734_bfr_before (
		.din(new_net_4734),
		.dout(new_net_4733)
	);

	bfr new_net_4735_bfr_before (
		.din(new_net_4735),
		.dout(new_net_4734)
	);

	bfr new_net_4736_bfr_before (
		.din(new_net_4736),
		.dout(new_net_4735)
	);

	bfr new_net_4737_bfr_before (
		.din(new_net_4737),
		.dout(new_net_4736)
	);

	bfr new_net_4738_bfr_before (
		.din(new_net_4738),
		.dout(new_net_4737)
	);

	bfr new_net_4739_bfr_before (
		.din(new_net_4739),
		.dout(new_net_4738)
	);

	bfr new_net_4740_bfr_before (
		.din(new_net_4740),
		.dout(new_net_4739)
	);

	spl2 n_0046__v_fanout (
		.a(n_0046_),
		.b(new_net_1905),
		.c(new_net_4740)
	);

	bfr new_net_4741_bfr_before (
		.din(new_net_4741),
		.dout(new_net_109)
	);

	spl2 n_0226__v_fanout (
		.a(n_0226_),
		.b(new_net_4741),
		.c(new_net_108)
	);

	spl2 n_0207__v_fanout (
		.a(n_0207_),
		.b(new_net_1699),
		.c(new_net_1698)
	);

	bfr new_net_4742_bfr_before (
		.din(new_net_4742),
		.dout(new_net_596)
	);

	bfr new_net_4743_bfr_before (
		.din(new_net_4743),
		.dout(new_net_4742)
	);

	bfr new_net_4744_bfr_before (
		.din(new_net_4744),
		.dout(new_net_4743)
	);

	bfr new_net_4745_bfr_before (
		.din(new_net_4745),
		.dout(new_net_4744)
	);

	spl2 n_0029__v_fanout (
		.a(n_0029_),
		.b(new_net_597),
		.c(new_net_4745)
	);

	spl2 n_0933__v_fanout (
		.a(n_0933_),
		.b(new_net_1099),
		.c(new_net_1098)
	);

	spl2 n_1072__v_fanout (
		.a(n_1072_),
		.b(new_net_865),
		.c(new_net_864)
	);

	bfr new_net_4746_bfr_before (
		.din(new_net_4746),
		.dout(new_net_1260)
	);

	bfr new_net_4747_bfr_before (
		.din(new_net_4747),
		.dout(new_net_4746)
	);

	spl4L n_0691__v_fanout (
		.a(n_0691_),
		.b(new_net_1261),
		.c(new_net_4747),
		.d(new_net_1262),
		.e(new_net_1259)
	);

	bfr new_net_4748_bfr_before (
		.din(new_net_4748),
		.dout(new_net_1190)
	);

	bfr new_net_4749_bfr_before (
		.din(new_net_4749),
		.dout(new_net_4748)
	);

	bfr new_net_4750_bfr_before (
		.din(new_net_4750),
		.dout(new_net_4749)
	);

	bfr new_net_4751_bfr_before (
		.din(new_net_4751),
		.dout(new_net_4750)
	);

	bfr new_net_4752_bfr_before (
		.din(new_net_4752),
		.dout(new_net_4751)
	);

	bfr new_net_4753_bfr_before (
		.din(new_net_4753),
		.dout(new_net_4752)
	);

	bfr new_net_4754_bfr_before (
		.din(new_net_4754),
		.dout(new_net_4753)
	);

	bfr new_net_4755_bfr_before (
		.din(new_net_4755),
		.dout(new_net_4754)
	);

	bfr new_net_4756_bfr_before (
		.din(new_net_4756),
		.dout(new_net_4755)
	);

	bfr new_net_4757_bfr_before (
		.din(new_net_4757),
		.dout(new_net_4756)
	);

	bfr new_net_4758_bfr_before (
		.din(new_net_4758),
		.dout(new_net_4757)
	);

	bfr new_net_4759_bfr_before (
		.din(new_net_4759),
		.dout(new_net_4758)
	);

	spl2 n_1337__v_fanout (
		.a(n_1337_),
		.b(new_net_4759),
		.c(new_net_1189)
	);

	bfr new_net_4760_bfr_before (
		.din(new_net_4760),
		.dout(new_net_2109)
	);

	spl3L n_1315__v_fanout (
		.a(n_1315_),
		.b(new_net_1153),
		.c(new_net_1151),
		.d(new_net_4760)
	);

	spl2 n_0675__v_fanout (
		.a(n_0675_),
		.b(new_net_1802),
		.c(new_net_1801)
	);

	spl2 n_1015__v_fanout (
		.a(n_1015_),
		.b(new_net_1025),
		.c(new_net_1024)
	);

	spl2 n_0244__v_fanout (
		.a(n_0244_),
		.b(new_net_720),
		.c(new_net_719)
	);

	bfr new_net_4761_bfr_before (
		.din(new_net_4761),
		.dout(new_net_1367)
	);

	spl2 n_0275__v_fanout (
		.a(n_0275_),
		.b(new_net_4761),
		.c(new_net_1366)
	);

	spl2 n_1081__v_fanout (
		.a(n_1081_),
		.b(new_net_1546),
		.c(new_net_1545)
	);

	spl2 n_0912__v_fanout (
		.a(n_0912_),
		.b(new_net_1523),
		.c(new_net_1522)
	);

	spl2 n_0942__v_fanout (
		.a(n_0942_),
		.b(new_net_1230),
		.c(new_net_1229)
	);

	bfr new_net_4762_bfr_before (
		.din(new_net_4762),
		.dout(new_net_1732)
	);

	bfr new_net_4763_bfr_before (
		.din(new_net_4763),
		.dout(new_net_4762)
	);

	bfr new_net_4764_bfr_before (
		.din(new_net_4764),
		.dout(new_net_4763)
	);

	bfr new_net_4765_bfr_before (
		.din(new_net_4765),
		.dout(new_net_4764)
	);

	bfr new_net_4766_bfr_before (
		.din(new_net_4766),
		.dout(new_net_4765)
	);

	spl3L n_1301__v_fanout (
		.a(n_1301_),
		.b(new_net_1734),
		.c(new_net_4766),
		.d(new_net_1733)
	);

	bfr new_net_4767_bfr_before (
		.din(new_net_4767),
		.dout(new_net_1670)
	);

	bfr new_net_4768_bfr_before (
		.din(new_net_4768),
		.dout(new_net_4767)
	);

	bfr new_net_4769_bfr_before (
		.din(new_net_4769),
		.dout(new_net_4768)
	);

	bfr new_net_4770_bfr_before (
		.din(new_net_4770),
		.dout(new_net_4769)
	);

	bfr new_net_4771_bfr_before (
		.din(new_net_4771),
		.dout(new_net_4770)
	);

	spl2 n_0696__v_fanout (
		.a(n_0696_),
		.b(new_net_1671),
		.c(new_net_4771)
	);

	bfr new_net_4772_bfr_before (
		.din(new_net_4772),
		.dout(new_net_586)
	);

	bfr new_net_4773_bfr_before (
		.din(new_net_4773),
		.dout(new_net_4772)
	);

	bfr new_net_4774_bfr_before (
		.din(new_net_4774),
		.dout(new_net_587)
	);

	spl3L n_1348__v_fanout (
		.a(n_1348_),
		.b(new_net_4774),
		.c(new_net_4773),
		.d(new_net_588)
	);

	spl2 n_0049__v_fanout (
		.a(n_0049_),
		.b(new_net_1031),
		.c(new_net_1030)
	);

	spl2 n_1024__v_fanout (
		.a(n_1024_),
		.b(new_net_1901),
		.c(new_net_1900)
	);

	bfr new_net_4775_bfr_before (
		.din(new_net_4775),
		.dout(new_net_903)
	);

	spl2 n_1351__v_fanout (
		.a(n_1351_),
		.b(new_net_2117),
		.c(new_net_4775)
	);

	bfr new_net_4776_bfr_before (
		.din(new_net_4776),
		.dout(new_net_593)
	);

	bfr new_net_4777_bfr_before (
		.din(new_net_4777),
		.dout(new_net_4776)
	);

	bfr new_net_4778_bfr_before (
		.din(new_net_4778),
		.dout(new_net_4777)
	);

	bfr new_net_4779_bfr_before (
		.din(new_net_4779),
		.dout(new_net_4778)
	);

	bfr new_net_4780_bfr_before (
		.din(new_net_4780),
		.dout(new_net_4779)
	);

	bfr new_net_4781_bfr_before (
		.din(new_net_4781),
		.dout(new_net_4780)
	);

	bfr new_net_4782_bfr_before (
		.din(new_net_4782),
		.dout(new_net_4781)
	);

	bfr new_net_4783_bfr_before (
		.din(new_net_4783),
		.dout(new_net_4782)
	);

	bfr new_net_4784_bfr_before (
		.din(new_net_4784),
		.dout(new_net_4783)
	);

	spl3L n_0098__v_fanout (
		.a(n_0098_),
		.b(new_net_594),
		.c(new_net_4784),
		.d(new_net_595)
	);

	spl2 n_1369__v_fanout (
		.a(n_1369_),
		.b(new_net_507),
		.c(new_net_2118)
	);

	spl2 n_1048__v_fanout (
		.a(n_1048_),
		.b(new_net_1714),
		.c(new_net_1713)
	);

	spl2 n_1302__v_fanout (
		.a(n_1302_),
		.b(new_net_1816),
		.c(new_net_1815)
	);

	bfr new_net_4785_bfr_before (
		.din(new_net_4785),
		.dout(new_net_311)
	);

	bfr new_net_4786_bfr_before (
		.din(new_net_4786),
		.dout(new_net_4785)
	);

	spl2 n_1305__v_fanout (
		.a(n_1305_),
		.b(new_net_312),
		.c(new_net_4786)
	);

	bfr new_net_4787_bfr_before (
		.din(new_net_4787),
		.dout(new_net_70)
	);

	bfr new_net_4788_bfr_before (
		.din(new_net_4788),
		.dout(new_net_4787)
	);

	bfr new_net_4789_bfr_before (
		.din(new_net_4789),
		.dout(new_net_4788)
	);

	bfr new_net_4790_bfr_before (
		.din(new_net_4790),
		.dout(new_net_4789)
	);

	bfr new_net_4791_bfr_before (
		.din(new_net_4791),
		.dout(new_net_4790)
	);

	bfr new_net_4792_bfr_before (
		.din(new_net_4792),
		.dout(new_net_4791)
	);

	bfr new_net_4793_bfr_before (
		.din(new_net_4793),
		.dout(new_net_4792)
	);

	bfr new_net_4794_bfr_before (
		.din(new_net_4794),
		.dout(new_net_4793)
	);

	spl2 n_1328__v_fanout (
		.a(n_1328_),
		.b(new_net_4794),
		.c(new_net_69)
	);

	spl3L n_0024__v_fanout (
		.a(n_0024_),
		.b(new_net_1370),
		.c(new_net_1368),
		.d(new_net_1369)
	);

	spl2 n_0996__v_fanout (
		.a(n_0996_),
		.b(new_net_629),
		.c(new_net_628)
	);

	bfr new_net_4795_bfr_before (
		.din(new_net_4795),
		.dout(new_net_2102)
	);

	bfr new_net_4796_bfr_before (
		.din(new_net_4796),
		.dout(new_net_4795)
	);

	bfr new_net_4797_bfr_before (
		.din(new_net_4797),
		.dout(new_net_4796)
	);

	bfr new_net_4798_bfr_before (
		.din(new_net_4798),
		.dout(new_net_4797)
	);

	bfr new_net_4799_bfr_before (
		.din(new_net_4799),
		.dout(new_net_4798)
	);

	bfr new_net_4800_bfr_before (
		.din(new_net_4800),
		.dout(new_net_4799)
	);

	bfr new_net_4801_bfr_before (
		.din(new_net_4801),
		.dout(new_net_4800)
	);

	bfr new_net_4802_bfr_before (
		.din(new_net_4802),
		.dout(new_net_4801)
	);

	bfr new_net_4803_bfr_before (
		.din(new_net_4803),
		.dout(new_net_4802)
	);

	bfr new_net_4804_bfr_before (
		.din(new_net_4804),
		.dout(new_net_4803)
	);

	bfr new_net_4805_bfr_before (
		.din(new_net_4805),
		.dout(new_net_4804)
	);

	bfr new_net_4806_bfr_before (
		.din(new_net_4806),
		.dout(new_net_4805)
	);

	bfr new_net_4807_bfr_before (
		.din(new_net_4807),
		.dout(new_net_4806)
	);

	bfr new_net_4808_bfr_before (
		.din(new_net_4808),
		.dout(new_net_4807)
	);

	bfr new_net_4809_bfr_before (
		.din(new_net_4809),
		.dout(new_net_4808)
	);

	bfr new_net_4810_bfr_before (
		.din(new_net_4810),
		.dout(new_net_4809)
	);

	bfr new_net_4811_bfr_before (
		.din(new_net_4811),
		.dout(new_net_4810)
	);

	bfr new_net_4812_bfr_before (
		.din(new_net_4812),
		.dout(new_net_4811)
	);

	bfr new_net_4813_bfr_before (
		.din(new_net_4813),
		.dout(new_net_4812)
	);

	bfr new_net_4814_bfr_before (
		.din(new_net_4814),
		.dout(new_net_4813)
	);

	bfr new_net_4815_bfr_before (
		.din(new_net_4815),
		.dout(new_net_4814)
	);

	bfr new_net_4816_bfr_before (
		.din(new_net_4816),
		.dout(new_net_4815)
	);

	bfr new_net_4817_bfr_before (
		.din(new_net_4817),
		.dout(new_net_4816)
	);

	bfr new_net_4818_bfr_before (
		.din(new_net_4818),
		.dout(new_net_4817)
	);

	bfr new_net_4819_bfr_before (
		.din(new_net_4819),
		.dout(new_net_4818)
	);

	bfr new_net_4820_bfr_before (
		.din(new_net_4820),
		.dout(new_net_4819)
	);

	bfr new_net_4821_bfr_before (
		.din(new_net_4821),
		.dout(new_net_4820)
	);

	bfr new_net_4822_bfr_before (
		.din(new_net_4822),
		.dout(new_net_4821)
	);

	bfr new_net_4823_bfr_before (
		.din(new_net_4823),
		.dout(new_net_4822)
	);

	bfr new_net_4824_bfr_before (
		.din(new_net_4824),
		.dout(new_net_4823)
	);

	bfr new_net_4825_bfr_before (
		.din(new_net_4825),
		.dout(new_net_4824)
	);

	bfr new_net_4826_bfr_before (
		.din(new_net_4826),
		.dout(new_net_4825)
	);

	bfr new_net_4827_bfr_before (
		.din(new_net_4827),
		.dout(new_net_4826)
	);

	bfr new_net_4828_bfr_before (
		.din(new_net_4828),
		.dout(new_net_4827)
	);

	bfr new_net_4829_bfr_before (
		.din(new_net_4829),
		.dout(new_net_4828)
	);

	bfr new_net_4830_bfr_before (
		.din(new_net_4830),
		.dout(new_net_4829)
	);

	bfr new_net_4831_bfr_before (
		.din(new_net_4831),
		.dout(new_net_4830)
	);

	bfr new_net_4832_bfr_before (
		.din(new_net_4832),
		.dout(new_net_4831)
	);

	bfr new_net_4833_bfr_before (
		.din(new_net_4833),
		.dout(new_net_4832)
	);

	bfr new_net_4834_bfr_before (
		.din(new_net_4834),
		.dout(new_net_4833)
	);

	bfr new_net_4835_bfr_before (
		.din(new_net_4835),
		.dout(new_net_4834)
	);

	spl2 n_0026__v_fanout (
		.a(n_0026_),
		.b(new_net_531),
		.c(new_net_4835)
	);

	bfr new_net_4836_bfr_before (
		.din(new_net_4836),
		.dout(new_net_2116)
	);

	bfr new_net_4837_bfr_before (
		.din(new_net_4837),
		.dout(new_net_4836)
	);

	bfr new_net_4838_bfr_before (
		.din(new_net_4838),
		.dout(new_net_4837)
	);

	spl2 n_1333__v_fanout (
		.a(n_1333_),
		.b(new_net_4838),
		.c(new_net_1542)
	);

	spl2 n_0120__v_fanout (
		.a(n_0120_),
		.b(new_net_759),
		.c(new_net_758)
	);

	bfr new_net_4839_bfr_before (
		.din(new_net_4839),
		.dout(new_net_677)
	);

	bfr new_net_4840_bfr_before (
		.din(new_net_4840),
		.dout(new_net_4839)
	);

	bfr new_net_4841_bfr_before (
		.din(new_net_4841),
		.dout(new_net_4840)
	);

	bfr new_net_4842_bfr_before (
		.din(new_net_4842),
		.dout(new_net_4841)
	);

	bfr new_net_4843_bfr_before (
		.din(new_net_4843),
		.dout(new_net_4842)
	);

	bfr new_net_4844_bfr_before (
		.din(new_net_4844),
		.dout(new_net_4843)
	);

	bfr new_net_4845_bfr_before (
		.din(new_net_4845),
		.dout(new_net_4844)
	);

	bfr new_net_4846_bfr_before (
		.din(new_net_4846),
		.dout(new_net_4845)
	);

	bfr new_net_4847_bfr_before (
		.din(new_net_4847),
		.dout(new_net_4846)
	);

	bfr new_net_4848_bfr_before (
		.din(new_net_4848),
		.dout(new_net_4847)
	);

	bfr new_net_4849_bfr_before (
		.din(new_net_4849),
		.dout(new_net_4848)
	);

	bfr new_net_4850_bfr_before (
		.din(new_net_4850),
		.dout(new_net_4849)
	);

	bfr new_net_4851_bfr_before (
		.din(new_net_4851),
		.dout(new_net_4850)
	);

	bfr new_net_4852_bfr_before (
		.din(new_net_4852),
		.dout(new_net_4851)
	);

	bfr new_net_4853_bfr_before (
		.din(new_net_4853),
		.dout(new_net_4852)
	);

	bfr new_net_4854_bfr_before (
		.din(new_net_4854),
		.dout(new_net_4853)
	);

	bfr new_net_4855_bfr_before (
		.din(new_net_4855),
		.dout(new_net_4854)
	);

	bfr new_net_4856_bfr_before (
		.din(new_net_4856),
		.dout(new_net_4855)
	);

	bfr new_net_4857_bfr_before (
		.din(new_net_4857),
		.dout(new_net_4856)
	);

	bfr new_net_4858_bfr_before (
		.din(new_net_4858),
		.dout(new_net_4857)
	);

	bfr new_net_4859_bfr_before (
		.din(new_net_4859),
		.dout(new_net_4858)
	);

	bfr new_net_4860_bfr_before (
		.din(new_net_4860),
		.dout(new_net_4859)
	);

	bfr new_net_4861_bfr_before (
		.din(new_net_4861),
		.dout(new_net_4860)
	);

	bfr new_net_4862_bfr_before (
		.din(new_net_4862),
		.dout(new_net_4861)
	);

	bfr new_net_4863_bfr_before (
		.din(new_net_4863),
		.dout(new_net_4862)
	);

	bfr new_net_4864_bfr_before (
		.din(new_net_4864),
		.dout(new_net_4863)
	);

	bfr new_net_4865_bfr_before (
		.din(new_net_4865),
		.dout(new_net_4864)
	);

	bfr new_net_4866_bfr_before (
		.din(new_net_4866),
		.dout(new_net_4865)
	);

	bfr new_net_4867_bfr_before (
		.din(new_net_4867),
		.dout(new_net_4866)
	);

	bfr new_net_4868_bfr_before (
		.din(new_net_4868),
		.dout(new_net_4867)
	);

	bfr new_net_4869_bfr_before (
		.din(new_net_4869),
		.dout(new_net_4868)
	);

	bfr new_net_4870_bfr_before (
		.din(new_net_4870),
		.dout(new_net_4869)
	);

	bfr new_net_4871_bfr_before (
		.din(new_net_4871),
		.dout(new_net_4870)
	);

	bfr new_net_4872_bfr_before (
		.din(new_net_4872),
		.dout(new_net_4871)
	);

	bfr new_net_4873_bfr_before (
		.din(new_net_4873),
		.dout(new_net_4872)
	);

	bfr new_net_4874_bfr_before (
		.din(new_net_4874),
		.dout(new_net_4873)
	);

	bfr new_net_4875_bfr_before (
		.din(new_net_4875),
		.dout(new_net_4874)
	);

	bfr new_net_4876_bfr_before (
		.din(new_net_4876),
		.dout(new_net_4875)
	);

	spl3L n_0032__v_fanout (
		.a(n_0032_),
		.b(new_net_678),
		.c(new_net_676),
		.d(new_net_4876)
	);

	spl2 n_1057__v_fanout (
		.a(n_1057_),
		.b(new_net_1781),
		.c(new_net_1780)
	);

	spl2 n_1345__v_fanout (
		.a(n_1345_),
		.b(new_net_72),
		.c(new_net_71)
	);

	bfr new_net_4877_bfr_before (
		.din(new_net_4877),
		.dout(new_net_753)
	);

	spl2 n_0246__v_fanout (
		.a(n_0246_),
		.b(new_net_4877),
		.c(new_net_752)
	);

	bfr new_net_4878_bfr_before (
		.din(new_net_4878),
		.dout(new_net_2103)
	);

	bfr new_net_4879_bfr_before (
		.din(new_net_4879),
		.dout(new_net_4878)
	);

	bfr new_net_4880_bfr_before (
		.din(new_net_4880),
		.dout(new_net_4879)
	);

	spl2 n_0028__v_fanout (
		.a(n_0028_),
		.b(new_net_1778),
		.c(new_net_4880)
	);

	spl3L n_0053__v_fanout (
		.a(n_0053_),
		.b(new_net_1039),
		.c(new_net_1038),
		.d(new_net_1040)
	);

	bfr new_net_4881_bfr_before (
		.din(new_net_4881),
		.dout(new_net_1830)
	);

	bfr new_net_4882_bfr_before (
		.din(new_net_4882),
		.dout(new_net_4881)
	);

	bfr new_net_4883_bfr_before (
		.din(new_net_4883),
		.dout(new_net_4882)
	);

	bfr new_net_4884_bfr_before (
		.din(new_net_4884),
		.dout(new_net_4883)
	);

	bfr new_net_4885_bfr_before (
		.din(new_net_4885),
		.dout(new_net_4884)
	);

	bfr new_net_4886_bfr_before (
		.din(new_net_4886),
		.dout(new_net_4885)
	);

	bfr new_net_4887_bfr_before (
		.din(new_net_4887),
		.dout(new_net_4886)
	);

	bfr new_net_4888_bfr_before (
		.din(new_net_4888),
		.dout(new_net_4887)
	);

	spl2 n_1343__v_fanout (
		.a(n_1343_),
		.b(new_net_1831),
		.c(new_net_4888)
	);

	spl2 n_0100__v_fanout (
		.a(n_0100_),
		.b(new_net_812),
		.c(new_net_811)
	);

	bfr new_net_4889_bfr_before (
		.din(new_net_4889),
		.dout(new_net_1612)
	);

	bfr new_net_4890_bfr_before (
		.din(new_net_4890),
		.dout(new_net_4889)
	);

	bfr new_net_4891_bfr_before (
		.din(new_net_4891),
		.dout(new_net_4890)
	);

	spl2 new_net_2069_v_fanout (
		.a(new_net_2069),
		.b(new_net_4891),
		.c(new_net_1613)
	);

	bfr new_net_4892_bfr_before (
		.din(new_net_4892),
		.dout(new_net_1606)
	);

	spl2 n_0296__v_fanout (
		.a(n_0296_),
		.b(new_net_4892),
		.c(new_net_1605)
	);

	bfr new_net_4893_bfr_before (
		.din(new_net_4893),
		.dout(new_net_702)
	);

	bfr new_net_4894_bfr_before (
		.din(new_net_4894),
		.dout(new_net_705)
	);

	spl4L n_1349__v_fanout (
		.a(n_1349_),
		.b(new_net_704),
		.c(new_net_4894),
		.d(new_net_703),
		.e(new_net_4893)
	);

	bfr new_net_4895_bfr_before (
		.din(new_net_4895),
		.dout(new_net_1003)
	);

	bfr new_net_4896_bfr_before (
		.din(new_net_4896),
		.dout(new_net_4895)
	);

	bfr new_net_4897_bfr_before (
		.din(new_net_4897),
		.dout(new_net_4896)
	);

	bfr new_net_4898_bfr_before (
		.din(new_net_4898),
		.dout(new_net_4897)
	);

	bfr new_net_4899_bfr_before (
		.din(new_net_4899),
		.dout(new_net_4898)
	);

	bfr new_net_4900_bfr_before (
		.din(new_net_4900),
		.dout(new_net_4899)
	);

	bfr new_net_4901_bfr_before (
		.din(new_net_4901),
		.dout(new_net_4900)
	);

	bfr new_net_4902_bfr_before (
		.din(new_net_4902),
		.dout(new_net_4901)
	);

	bfr new_net_4903_bfr_before (
		.din(new_net_4903),
		.dout(new_net_4902)
	);

	bfr new_net_4904_bfr_before (
		.din(new_net_4904),
		.dout(new_net_4903)
	);

	bfr new_net_4905_bfr_before (
		.din(new_net_4905),
		.dout(new_net_4904)
	);

	bfr new_net_4906_bfr_before (
		.din(new_net_4906),
		.dout(new_net_4905)
	);

	bfr new_net_4907_bfr_before (
		.din(new_net_4907),
		.dout(new_net_4906)
	);

	bfr new_net_4908_bfr_before (
		.din(new_net_4908),
		.dout(new_net_4907)
	);

	bfr new_net_4909_bfr_before (
		.din(new_net_4909),
		.dout(new_net_4908)
	);

	bfr new_net_4910_bfr_before (
		.din(new_net_4910),
		.dout(new_net_4909)
	);

	bfr new_net_4911_bfr_before (
		.din(new_net_4911),
		.dout(new_net_4910)
	);

	bfr new_net_4912_bfr_before (
		.din(new_net_4912),
		.dout(new_net_4911)
	);

	bfr new_net_4913_bfr_before (
		.din(new_net_4913),
		.dout(new_net_4912)
	);

	bfr new_net_4914_bfr_before (
		.din(new_net_4914),
		.dout(new_net_4913)
	);

	bfr new_net_4915_bfr_before (
		.din(new_net_4915),
		.dout(new_net_4914)
	);

	bfr new_net_4916_bfr_before (
		.din(new_net_4916),
		.dout(new_net_4915)
	);

	bfr new_net_4917_bfr_before (
		.din(new_net_4917),
		.dout(new_net_4916)
	);

	bfr new_net_4918_bfr_before (
		.din(new_net_4918),
		.dout(new_net_4917)
	);

	bfr new_net_4919_bfr_before (
		.din(new_net_4919),
		.dout(new_net_4918)
	);

	bfr new_net_4920_bfr_before (
		.din(new_net_4920),
		.dout(new_net_4919)
	);

	bfr new_net_4921_bfr_before (
		.din(new_net_4921),
		.dout(new_net_4920)
	);

	bfr new_net_4922_bfr_before (
		.din(new_net_4922),
		.dout(new_net_4921)
	);

	bfr new_net_4923_bfr_before (
		.din(new_net_4923),
		.dout(new_net_4922)
	);

	bfr new_net_4924_bfr_before (
		.din(new_net_4924),
		.dout(new_net_4923)
	);

	bfr new_net_4925_bfr_before (
		.din(new_net_4925),
		.dout(new_net_4924)
	);

	bfr new_net_4926_bfr_before (
		.din(new_net_4926),
		.dout(new_net_4925)
	);

	bfr new_net_4927_bfr_before (
		.din(new_net_4927),
		.dout(new_net_4926)
	);

	bfr new_net_4928_bfr_before (
		.din(new_net_4928),
		.dout(new_net_4927)
	);

	bfr new_net_4929_bfr_before (
		.din(new_net_4929),
		.dout(new_net_4928)
	);

	spl4L n_1294__v_fanout (
		.a(n_1294_),
		.b(new_net_1004),
		.c(new_net_4929),
		.d(new_net_1005),
		.e(new_net_1002)
	);

	bfr new_net_4930_bfr_before (
		.din(new_net_4930),
		.dout(new_net_460)
	);

	bfr new_net_4931_bfr_before (
		.din(new_net_4931),
		.dout(new_net_4930)
	);

	bfr new_net_4932_bfr_before (
		.din(new_net_4932),
		.dout(new_net_4931)
	);

	bfr new_net_4933_bfr_before (
		.din(new_net_4933),
		.dout(new_net_4932)
	);

	spl2 n_1347__v_fanout (
		.a(n_1347_),
		.b(new_net_461),
		.c(new_net_4933)
	);

	bfr new_net_4934_bfr_before (
		.din(new_net_4934),
		.dout(new_net_1239)
	);

	spl2 n_1320__v_fanout (
		.a(n_1320_),
		.b(new_net_2111),
		.c(new_net_4934)
	);

	spl2 new_net_2099_v_fanout (
		.a(new_net_2099),
		.b(new_net_322),
		.c(new_net_319)
	);

	spl3L n_0104__v_fanout (
		.a(n_0104_),
		.b(new_net_1206),
		.c(new_net_1204),
		.d(new_net_1205)
	);

	bfr new_net_4935_bfr_before (
		.din(new_net_4935),
		.dout(new_net_438)
	);

	bfr new_net_4936_bfr_before (
		.din(new_net_4936),
		.dout(new_net_4935)
	);

	bfr new_net_4937_bfr_before (
		.din(new_net_4937),
		.dout(new_net_4936)
	);

	bfr new_net_4938_bfr_before (
		.din(new_net_4938),
		.dout(new_net_4937)
	);

	bfr new_net_4939_bfr_before (
		.din(new_net_4939),
		.dout(new_net_4938)
	);

	bfr new_net_4940_bfr_before (
		.din(new_net_4940),
		.dout(new_net_4939)
	);

	bfr new_net_4941_bfr_before (
		.din(new_net_4941),
		.dout(new_net_4940)
	);

	bfr new_net_4942_bfr_before (
		.din(new_net_4942),
		.dout(new_net_4941)
	);

	bfr new_net_4943_bfr_before (
		.din(new_net_4943),
		.dout(new_net_4942)
	);

	bfr new_net_4944_bfr_before (
		.din(new_net_4944),
		.dout(new_net_4943)
	);

	bfr new_net_4945_bfr_before (
		.din(new_net_4945),
		.dout(new_net_4944)
	);

	bfr new_net_4946_bfr_before (
		.din(new_net_4946),
		.dout(new_net_4945)
	);

	bfr new_net_4947_bfr_before (
		.din(new_net_4947),
		.dout(new_net_4946)
	);

	bfr new_net_4948_bfr_before (
		.din(new_net_4948),
		.dout(new_net_4947)
	);

	bfr new_net_4949_bfr_before (
		.din(new_net_4949),
		.dout(new_net_4948)
	);

	bfr new_net_4950_bfr_before (
		.din(new_net_4950),
		.dout(new_net_4949)
	);

	bfr new_net_4951_bfr_before (
		.din(new_net_4951),
		.dout(new_net_4950)
	);

	bfr new_net_4952_bfr_before (
		.din(new_net_4952),
		.dout(new_net_4951)
	);

	bfr new_net_4953_bfr_before (
		.din(new_net_4953),
		.dout(new_net_4952)
	);

	bfr new_net_4954_bfr_before (
		.din(new_net_4954),
		.dout(new_net_4953)
	);

	bfr new_net_4955_bfr_before (
		.din(new_net_4955),
		.dout(new_net_4954)
	);

	bfr new_net_4956_bfr_before (
		.din(new_net_4956),
		.dout(new_net_4955)
	);

	bfr new_net_4957_bfr_before (
		.din(new_net_4957),
		.dout(new_net_4956)
	);

	bfr new_net_4958_bfr_before (
		.din(new_net_4958),
		.dout(new_net_4957)
	);

	bfr new_net_4959_bfr_before (
		.din(new_net_4959),
		.dout(new_net_4958)
	);

	bfr new_net_4960_bfr_before (
		.din(new_net_4960),
		.dout(new_net_4959)
	);

	bfr new_net_4961_bfr_before (
		.din(new_net_4961),
		.dout(new_net_4960)
	);

	bfr new_net_4962_bfr_before (
		.din(new_net_4962),
		.dout(new_net_4961)
	);

	bfr new_net_4963_bfr_before (
		.din(new_net_4963),
		.dout(new_net_4962)
	);

	bfr new_net_4964_bfr_before (
		.din(new_net_4964),
		.dout(new_net_4963)
	);

	bfr new_net_4965_bfr_before (
		.din(new_net_4965),
		.dout(new_net_4964)
	);

	bfr new_net_4966_bfr_before (
		.din(new_net_4966),
		.dout(new_net_4965)
	);

	bfr new_net_4967_bfr_before (
		.din(new_net_4967),
		.dout(new_net_4966)
	);

	bfr new_net_4968_bfr_before (
		.din(new_net_4968),
		.dout(new_net_4967)
	);

	bfr new_net_4969_bfr_before (
		.din(new_net_4969),
		.dout(new_net_4968)
	);

	bfr new_net_4970_bfr_before (
		.din(new_net_4970),
		.dout(new_net_4969)
	);

	bfr new_net_4971_bfr_before (
		.din(new_net_4971),
		.dout(new_net_4970)
	);

	bfr new_net_4972_bfr_before (
		.din(new_net_4972),
		.dout(new_net_4971)
	);

	bfr new_net_4973_bfr_before (
		.din(new_net_4973),
		.dout(new_net_4972)
	);

	bfr new_net_4974_bfr_before (
		.din(new_net_4974),
		.dout(new_net_4973)
	);

	bfr new_net_4975_bfr_before (
		.din(new_net_4975),
		.dout(new_net_4974)
	);

	bfr new_net_4976_bfr_before (
		.din(new_net_4976),
		.dout(new_net_4975)
	);

	bfr new_net_4977_bfr_before (
		.din(new_net_4977),
		.dout(new_net_4976)
	);

	bfr new_net_4978_bfr_before (
		.din(new_net_4978),
		.dout(new_net_4977)
	);

	bfr new_net_4979_bfr_before (
		.din(new_net_4979),
		.dout(new_net_4978)
	);

	bfr new_net_4980_bfr_before (
		.din(new_net_4980),
		.dout(new_net_4979)
	);

	spl4L n_0023__v_fanout (
		.a(n_0023_),
		.b(new_net_436),
		.c(new_net_4980),
		.d(new_net_437),
		.e(new_net_435)
	);

	bfr new_net_4981_bfr_before (
		.din(new_net_4981),
		.dout(new_net_2055)
	);

	bfr new_net_4982_bfr_before (
		.din(new_net_4982),
		.dout(new_net_4981)
	);

	bfr new_net_4983_bfr_before (
		.din(new_net_4983),
		.dout(new_net_4982)
	);

	bfr new_net_4984_bfr_before (
		.din(new_net_4984),
		.dout(new_net_4983)
	);

	bfr new_net_4985_bfr_before (
		.din(new_net_4985),
		.dout(new_net_4984)
	);

	spl2 new_net_2054_v_fanout (
		.a(new_net_2054),
		.b(new_net_4985),
		.c(new_net_960)
	);

	spl2 new_net_2096_v_fanout (
		.a(new_net_2096),
		.b(new_net_1825),
		.c(new_net_1824)
	);

	bfr new_net_4986_bfr_before (
		.din(new_net_4986),
		.dout(new_net_1519)
	);

	bfr new_net_4987_bfr_before (
		.din(new_net_4987),
		.dout(new_net_4986)
	);

	bfr new_net_4988_bfr_before (
		.din(new_net_4988),
		.dout(new_net_4987)
	);

	bfr new_net_4989_bfr_before (
		.din(new_net_4989),
		.dout(new_net_4988)
	);

	spl2 n_1332__v_fanout (
		.a(n_1332_),
		.b(new_net_4989),
		.c(new_net_1518)
	);

	bfr new_net_4990_bfr_before (
		.din(new_net_4990),
		.dout(new_net_100)
	);

	bfr new_net_4991_bfr_before (
		.din(new_net_4991),
		.dout(new_net_4990)
	);

	bfr new_net_4992_bfr_before (
		.din(new_net_4992),
		.dout(new_net_4991)
	);

	bfr new_net_4993_bfr_before (
		.din(new_net_4993),
		.dout(new_net_4992)
	);

	bfr new_net_4994_bfr_before (
		.din(new_net_4994),
		.dout(new_net_4993)
	);

	bfr new_net_4995_bfr_before (
		.din(new_net_4995),
		.dout(new_net_4994)
	);

	bfr new_net_4996_bfr_before (
		.din(new_net_4996),
		.dout(new_net_4995)
	);

	bfr new_net_4997_bfr_before (
		.din(new_net_4997),
		.dout(new_net_4996)
	);

	spl2 n_0099__v_fanout (
		.a(n_0099_),
		.b(new_net_101),
		.c(new_net_4997)
	);

	bfr new_net_4998_bfr_before (
		.din(new_net_4998),
		.dout(new_net_1688)
	);

	bfr new_net_4999_bfr_before (
		.din(new_net_4999),
		.dout(new_net_4998)
	);

	bfr new_net_5000_bfr_before (
		.din(new_net_5000),
		.dout(new_net_4999)
	);

	bfr new_net_5001_bfr_before (
		.din(new_net_5001),
		.dout(new_net_5000)
	);

	bfr new_net_5002_bfr_before (
		.din(new_net_5002),
		.dout(new_net_5001)
	);

	bfr new_net_5003_bfr_before (
		.din(new_net_5003),
		.dout(new_net_5002)
	);

	bfr new_net_5004_bfr_before (
		.din(new_net_5004),
		.dout(new_net_5003)
	);

	bfr new_net_5005_bfr_before (
		.din(new_net_5005),
		.dout(new_net_5004)
	);

	bfr new_net_5006_bfr_before (
		.din(new_net_5006),
		.dout(new_net_5005)
	);

	bfr new_net_5007_bfr_before (
		.din(new_net_5007),
		.dout(new_net_5006)
	);

	bfr new_net_5008_bfr_before (
		.din(new_net_5008),
		.dout(new_net_5007)
	);

	bfr new_net_5009_bfr_before (
		.din(new_net_5009),
		.dout(new_net_5008)
	);

	bfr new_net_5010_bfr_before (
		.din(new_net_5010),
		.dout(new_net_5009)
	);

	bfr new_net_5011_bfr_before (
		.din(new_net_5011),
		.dout(new_net_5010)
	);

	bfr new_net_5012_bfr_before (
		.din(new_net_5012),
		.dout(new_net_5011)
	);

	bfr new_net_5013_bfr_before (
		.din(new_net_5013),
		.dout(new_net_5012)
	);

	bfr new_net_5014_bfr_before (
		.din(new_net_5014),
		.dout(new_net_5013)
	);

	bfr new_net_5015_bfr_before (
		.din(new_net_5015),
		.dout(new_net_5014)
	);

	bfr new_net_5016_bfr_before (
		.din(new_net_5016),
		.dout(new_net_5015)
	);

	bfr new_net_5017_bfr_before (
		.din(new_net_5017),
		.dout(new_net_5016)
	);

	bfr new_net_5018_bfr_before (
		.din(new_net_5018),
		.dout(new_net_5017)
	);

	bfr new_net_5019_bfr_before (
		.din(new_net_5019),
		.dout(new_net_5018)
	);

	bfr new_net_5020_bfr_before (
		.din(new_net_5020),
		.dout(new_net_5019)
	);

	bfr new_net_5021_bfr_before (
		.din(new_net_5021),
		.dout(new_net_5020)
	);

	bfr new_net_5022_bfr_before (
		.din(new_net_5022),
		.dout(new_net_5021)
	);

	bfr new_net_5023_bfr_before (
		.din(new_net_5023),
		.dout(new_net_5022)
	);

	bfr new_net_5024_bfr_before (
		.din(new_net_5024),
		.dout(new_net_5023)
	);

	bfr new_net_5025_bfr_before (
		.din(new_net_5025),
		.dout(new_net_5024)
	);

	bfr new_net_5026_bfr_before (
		.din(new_net_5026),
		.dout(new_net_5025)
	);

	bfr new_net_5027_bfr_before (
		.din(new_net_5027),
		.dout(new_net_5026)
	);

	bfr new_net_5028_bfr_before (
		.din(new_net_5028),
		.dout(new_net_5027)
	);

	bfr new_net_5029_bfr_before (
		.din(new_net_5029),
		.dout(new_net_5028)
	);

	bfr new_net_5030_bfr_before (
		.din(new_net_5030),
		.dout(new_net_5029)
	);

	bfr new_net_5031_bfr_before (
		.din(new_net_5031),
		.dout(new_net_5030)
	);

	bfr new_net_5032_bfr_before (
		.din(new_net_5032),
		.dout(new_net_5031)
	);

	bfr new_net_5033_bfr_before (
		.din(new_net_5033),
		.dout(new_net_5032)
	);

	bfr new_net_5034_bfr_before (
		.din(new_net_5034),
		.dout(new_net_5033)
	);

	bfr new_net_5035_bfr_before (
		.din(new_net_5035),
		.dout(new_net_5034)
	);

	bfr new_net_5036_bfr_before (
		.din(new_net_5036),
		.dout(new_net_5035)
	);

	bfr new_net_5037_bfr_before (
		.din(new_net_5037),
		.dout(new_net_5036)
	);

	spl2 n_0027__v_fanout (
		.a(n_0027_),
		.b(new_net_1689),
		.c(new_net_5037)
	);

	bfr new_net_5038_bfr_before (
		.din(new_net_5038),
		.dout(new_net_416)
	);

	bfr new_net_5039_bfr_before (
		.din(new_net_5039),
		.dout(new_net_5038)
	);

	spl2 n_0326__v_fanout (
		.a(n_0326_),
		.b(new_net_5039),
		.c(new_net_415)
	);

	bfr new_net_5040_bfr_before (
		.din(new_net_5040),
		.dout(new_net_932)
	);

	bfr new_net_5041_bfr_before (
		.din(new_net_5041),
		.dout(new_net_5040)
	);

	spl4L n_0052__v_fanout (
		.a(n_0052_),
		.b(new_net_933),
		.c(new_net_934),
		.d(new_net_935),
		.e(new_net_5041)
	);

	spl2 n_1093__v_fanout (
		.a(n_1093_),
		.b(new_net_1770),
		.c(new_net_1769)
	);

	spl3L n_1325__v_fanout (
		.a(n_1325_),
		.b(new_net_1361),
		.c(new_net_1358),
		.d(new_net_2115)
	);

	bfr new_net_5042_bfr_before (
		.din(new_net_5042),
		.dout(new_net_1706)
	);

	bfr new_net_5043_bfr_before (
		.din(new_net_5043),
		.dout(new_net_5042)
	);

	bfr new_net_5044_bfr_before (
		.din(new_net_5044),
		.dout(new_net_5043)
	);

	bfr new_net_5045_bfr_before (
		.din(new_net_5045),
		.dout(new_net_5044)
	);

	bfr new_net_5046_bfr_before (
		.din(new_net_5046),
		.dout(new_net_5045)
	);

	spl2 n_0280__v_fanout (
		.a(n_0280_),
		.b(new_net_5046),
		.c(new_net_1705)
	);

	bfr new_net_5047_bfr_before (
		.din(new_net_5047),
		.dout(new_net_880)
	);

	spl2 n_0253__v_fanout (
		.a(n_0253_),
		.b(new_net_5047),
		.c(new_net_879)
	);

	spl2 n_0243__v_fanout (
		.a(n_0243_),
		.b(new_net_693),
		.c(new_net_692)
	);

	bfr new_net_5048_bfr_after (
		.din(n_0966_),
		.dout(new_net_5048)
	);

	spl2 n_0966__v_fanout (
		.a(new_net_5048),
		.b(new_net_1750),
		.c(new_net_1749)
	);

	bfr new_net_5049_bfr_before (
		.din(new_net_5049),
		.dout(new_net_1530)
	);

	bfr new_net_5050_bfr_before (
		.din(new_net_5050),
		.dout(new_net_5049)
	);

	bfr new_net_5051_bfr_before (
		.din(new_net_5051),
		.dout(new_net_5050)
	);

	bfr new_net_5052_bfr_before (
		.din(new_net_5052),
		.dout(new_net_5051)
	);

	bfr new_net_5053_bfr_before (
		.din(new_net_5053),
		.dout(new_net_5052)
	);

	bfr new_net_5054_bfr_before (
		.din(new_net_5054),
		.dout(new_net_5053)
	);

	bfr new_net_5055_bfr_before (
		.din(new_net_5055),
		.dout(new_net_5054)
	);

	bfr new_net_5056_bfr_before (
		.din(new_net_5056),
		.dout(new_net_5055)
	);

	bfr new_net_5057_bfr_before (
		.din(new_net_5057),
		.dout(new_net_5056)
	);

	bfr new_net_5058_bfr_before (
		.din(new_net_5058),
		.dout(new_net_5057)
	);

	bfr new_net_5059_bfr_before (
		.din(new_net_5059),
		.dout(new_net_5058)
	);

	bfr new_net_5060_bfr_before (
		.din(new_net_5060),
		.dout(new_net_5059)
	);

	bfr new_net_5061_bfr_before (
		.din(new_net_5061),
		.dout(new_net_5060)
	);

	bfr new_net_5062_bfr_before (
		.din(new_net_5062),
		.dout(new_net_5061)
	);

	bfr new_net_5063_bfr_before (
		.din(new_net_5063),
		.dout(new_net_5062)
	);

	bfr new_net_5064_bfr_before (
		.din(new_net_5064),
		.dout(new_net_5063)
	);

	bfr new_net_5065_bfr_before (
		.din(new_net_5065),
		.dout(new_net_5064)
	);

	bfr new_net_5066_bfr_before (
		.din(new_net_5066),
		.dout(new_net_5065)
	);

	bfr new_net_5067_bfr_before (
		.din(new_net_5067),
		.dout(new_net_5066)
	);

	bfr new_net_5068_bfr_before (
		.din(new_net_5068),
		.dout(new_net_5067)
	);

	bfr new_net_5069_bfr_before (
		.din(new_net_5069),
		.dout(new_net_5068)
	);

	bfr new_net_5070_bfr_before (
		.din(new_net_5070),
		.dout(new_net_5069)
	);

	bfr new_net_5071_bfr_before (
		.din(new_net_5071),
		.dout(new_net_5070)
	);

	bfr new_net_5072_bfr_before (
		.din(new_net_5072),
		.dout(new_net_5071)
	);

	bfr new_net_5073_bfr_before (
		.din(new_net_5073),
		.dout(new_net_5072)
	);

	bfr new_net_5074_bfr_before (
		.din(new_net_5074),
		.dout(new_net_5073)
	);

	bfr new_net_5075_bfr_before (
		.din(new_net_5075),
		.dout(new_net_5074)
	);

	bfr new_net_5076_bfr_before (
		.din(new_net_5076),
		.dout(new_net_5075)
	);

	bfr new_net_5077_bfr_before (
		.din(new_net_5077),
		.dout(new_net_5076)
	);

	spl2 n_1299__v_fanout (
		.a(n_1299_),
		.b(new_net_1531),
		.c(new_net_5077)
	);

	bfr new_net_5078_bfr_before (
		.din(new_net_5078),
		.dout(new_net_2104)
	);

	spl4L n_0037__v_fanout (
		.a(n_0037_),
		.b(new_net_787),
		.c(new_net_784),
		.d(new_net_5078),
		.e(new_net_783)
	);

	bfr new_net_5079_bfr_before (
		.din(new_net_5079),
		.dout(new_net_1587)
	);

	spl2 n_0327__v_fanout (
		.a(n_0327_),
		.b(new_net_5079),
		.c(new_net_1586)
	);

	spl2 n_1108__v_fanout (
		.a(n_1108_),
		.b(new_net_111),
		.c(new_net_110)
	);

	bfr new_net_5080_bfr_before (
		.din(new_net_5080),
		.dout(new_net_2107)
	);

	bfr new_net_5081_bfr_before (
		.din(new_net_5081),
		.dout(new_net_5080)
	);

	bfr new_net_5082_bfr_before (
		.din(new_net_5082),
		.dout(new_net_5081)
	);

	bfr new_net_5083_bfr_before (
		.din(new_net_5083),
		.dout(new_net_5082)
	);

	spl2 n_0680__v_fanout (
		.a(n_0680_),
		.b(new_net_738),
		.c(new_net_5083)
	);

	bfr new_net_5084_bfr_before (
		.din(new_net_5084),
		.dout(new_net_2106)
	);

	bfr new_net_5085_bfr_before (
		.din(new_net_5085),
		.dout(new_net_5084)
	);

	bfr new_net_5086_bfr_before (
		.din(new_net_5086),
		.dout(new_net_5085)
	);

	bfr new_net_5087_bfr_before (
		.din(new_net_5087),
		.dout(new_net_5086)
	);

	bfr new_net_5088_bfr_before (
		.din(new_net_5088),
		.dout(new_net_5087)
	);

	bfr new_net_5089_bfr_before (
		.din(new_net_5089),
		.dout(new_net_5088)
	);

	bfr new_net_5090_bfr_before (
		.din(new_net_5090),
		.dout(new_net_5089)
	);

	bfr new_net_5091_bfr_before (
		.din(new_net_5091),
		.dout(new_net_5090)
	);

	bfr new_net_5092_bfr_before (
		.din(new_net_5092),
		.dout(new_net_5091)
	);

	spl2 n_0674__v_fanout (
		.a(n_0674_),
		.b(new_net_5092),
		.c(new_net_1874)
	);

	bfr new_net_5093_bfr_before (
		.din(new_net_5093),
		.dout(new_net_656)
	);

	bfr new_net_5094_bfr_before (
		.din(new_net_5094),
		.dout(new_net_5093)
	);

	spl4L n_0031__v_fanout (
		.a(n_0031_),
		.b(new_net_657),
		.c(new_net_5094),
		.d(new_net_658),
		.e(new_net_655)
	);

	spl2 new_net_2080_v_fanout (
		.a(new_net_2080),
		.b(new_net_1395),
		.c(new_net_1392)
	);

	spl2 n_0208__v_fanout (
		.a(n_0208_),
		.b(new_net_909),
		.c(new_net_908)
	);

	bfr new_net_5095_bfr_before (
		.din(new_net_5095),
		.dout(new_net_318)
	);

	bfr new_net_5096_bfr_before (
		.din(new_net_5096),
		.dout(new_net_5095)
	);

	bfr new_net_5097_bfr_before (
		.din(new_net_5097),
		.dout(new_net_5096)
	);

	bfr new_net_5098_bfr_before (
		.din(new_net_5098),
		.dout(new_net_5097)
	);

	bfr new_net_5099_bfr_before (
		.din(new_net_5099),
		.dout(new_net_5098)
	);

	bfr new_net_5100_bfr_before (
		.din(new_net_5100),
		.dout(new_net_5099)
	);

	bfr new_net_5101_bfr_before (
		.din(new_net_5101),
		.dout(new_net_5100)
	);

	bfr new_net_5102_bfr_before (
		.din(new_net_5102),
		.dout(new_net_5101)
	);

	bfr new_net_5103_bfr_before (
		.din(new_net_5103),
		.dout(new_net_5102)
	);

	spl2 n_1329__v_fanout (
		.a(n_1329_),
		.b(new_net_5103),
		.c(new_net_317)
	);

	spl2 n_0317__v_fanout (
		.a(n_0317_),
		.b(new_net_1363),
		.c(new_net_1362)
	);

	bfr new_net_5104_bfr_before (
		.din(new_net_5104),
		.dout(new_net_987)
	);

	spl2 n_0314__v_fanout (
		.a(n_0314_),
		.b(new_net_5104),
		.c(new_net_986)
	);

	bfr new_net_5105_bfr_before (
		.din(new_net_5105),
		.dout(new_net_323)
	);

	bfr new_net_5106_bfr_before (
		.din(new_net_5106),
		.dout(new_net_5105)
	);

	spl4L n_0103__v_fanout (
		.a(n_0103_),
		.b(new_net_326),
		.c(new_net_324),
		.d(new_net_325),
		.e(new_net_5106)
	);

	spl2 n_1322__v_fanout (
		.a(n_1322_),
		.b(new_net_1418),
		.c(new_net_2112)
	);

	spl2 new_net_2079_v_fanout (
		.a(new_net_2079),
		.b(new_net_766),
		.c(new_net_764)
	);

	bfr new_net_5107_bfr_before (
		.din(new_net_5107),
		.dout(new_net_1066)
	);

	bfr new_net_5108_bfr_before (
		.din(new_net_5108),
		.dout(new_net_5107)
	);

	bfr new_net_5109_bfr_before (
		.din(new_net_5109),
		.dout(new_net_5108)
	);

	spl4L n_0690__v_fanout (
		.a(n_0690_),
		.b(new_net_1065),
		.c(new_net_5109),
		.d(new_net_1064),
		.e(new_net_1063)
	);

	bfr new_net_5110_bfr_before (
		.din(new_net_5110),
		.dout(new_net_984)
	);

	bfr new_net_5111_bfr_before (
		.din(new_net_5111),
		.dout(new_net_5110)
	);

	bfr new_net_5112_bfr_before (
		.din(new_net_5112),
		.dout(new_net_5111)
	);

	bfr new_net_5113_bfr_before (
		.din(new_net_5113),
		.dout(new_net_5112)
	);

	bfr new_net_5114_bfr_before (
		.din(new_net_5114),
		.dout(new_net_5113)
	);

	bfr new_net_5115_bfr_before (
		.din(new_net_5115),
		.dout(new_net_5114)
	);

	bfr new_net_5116_bfr_before (
		.din(new_net_5116),
		.dout(new_net_5115)
	);

	bfr new_net_5117_bfr_before (
		.din(new_net_5117),
		.dout(new_net_5116)
	);

	spl2 n_0047__v_fanout (
		.a(n_0047_),
		.b(new_net_985),
		.c(new_net_5117)
	);

	bfr new_net_5118_bfr_before (
		.din(new_net_5118),
		.dout(new_net_632)
	);

	bfr new_net_5119_bfr_before (
		.din(new_net_5119),
		.dout(new_net_5118)
	);

	spl3L n_0030__v_fanout (
		.a(n_0030_),
		.b(new_net_633),
		.c(new_net_5119),
		.d(new_net_634)
	);

	spl2 n_0921__v_fanout (
		.a(n_0921_),
		.b(new_net_1701),
		.c(new_net_1700)
	);

	bfr new_net_5120_bfr_before (
		.din(new_net_5120),
		.dout(new_net_301)
	);

	bfr new_net_5121_bfr_before (
		.din(new_net_5121),
		.dout(new_net_5120)
	);

	bfr new_net_5122_bfr_before (
		.din(new_net_5122),
		.dout(new_net_5121)
	);

	bfr new_net_5123_bfr_before (
		.din(new_net_5123),
		.dout(new_net_5122)
	);

	spl2 n_0102__v_fanout (
		.a(n_0102_),
		.b(new_net_302),
		.c(new_net_5123)
	);

	bfr new_net_5124_bfr_before (
		.din(new_net_5124),
		.dout(new_net_354)
	);

	bfr new_net_5125_bfr_before (
		.din(new_net_5125),
		.dout(new_net_5124)
	);

	bfr new_net_5126_bfr_before (
		.din(new_net_5126),
		.dout(new_net_5125)
	);

	spl2 n_0684__v_fanout (
		.a(n_0684_),
		.b(new_net_5126),
		.c(new_net_353)
	);

	bfr new_net_5127_bfr_after (
		.din(n_1036_),
		.dout(new_net_5127)
	);

	bfr new_net_5128_bfr_after (
		.din(new_net_5127),
		.dout(new_net_5128)
	);

	bfr new_net_5129_bfr_after (
		.din(new_net_5128),
		.dout(new_net_5129)
	);

	spl2 n_1036__v_fanout (
		.a(new_net_5129),
		.b(new_net_1372),
		.c(new_net_1371)
	);

	bfr new_net_5130_bfr_before (
		.din(new_net_5130),
		.dout(new_net_735)
	);

	bfr new_net_5131_bfr_before (
		.din(new_net_5131),
		.dout(new_net_5130)
	);

	spl3L new_net_2101_v_fanout (
		.a(new_net_2101),
		.b(new_net_5131),
		.c(new_net_734),
		.d(new_net_736)
	);

	spl2 n_0978__v_fanout (
		.a(n_0978_),
		.b(new_net_46),
		.c(new_net_45)
	);

	bfr new_net_5132_bfr_before (
		.din(new_net_5132),
		.dout(new_net_700)
	);

	bfr new_net_5133_bfr_before (
		.din(new_net_5133),
		.dout(new_net_5132)
	);

	bfr new_net_5134_bfr_before (
		.din(new_net_5134),
		.dout(new_net_5133)
	);

	bfr new_net_5135_bfr_before (
		.din(new_net_5135),
		.dout(new_net_5134)
	);

	bfr new_net_5136_bfr_before (
		.din(new_net_5136),
		.dout(new_net_5135)
	);

	bfr new_net_5137_bfr_before (
		.din(new_net_5137),
		.dout(new_net_5136)
	);

	bfr new_net_5138_bfr_before (
		.din(new_net_5138),
		.dout(new_net_5137)
	);

	bfr new_net_5139_bfr_before (
		.din(new_net_5139),
		.dout(new_net_5138)
	);

	bfr new_net_5140_bfr_before (
		.din(new_net_5140),
		.dout(new_net_5139)
	);

	bfr new_net_5141_bfr_before (
		.din(new_net_5141),
		.dout(new_net_5140)
	);

	bfr new_net_5142_bfr_before (
		.din(new_net_5142),
		.dout(new_net_5141)
	);

	bfr new_net_5143_bfr_before (
		.din(new_net_5143),
		.dout(new_net_5142)
	);

	bfr new_net_5144_bfr_before (
		.din(new_net_5144),
		.dout(new_net_5143)
	);

	bfr new_net_5145_bfr_before (
		.din(new_net_5145),
		.dout(new_net_5144)
	);

	bfr new_net_5146_bfr_before (
		.din(new_net_5146),
		.dout(new_net_5145)
	);

	bfr new_net_5147_bfr_before (
		.din(new_net_5147),
		.dout(new_net_5146)
	);

	bfr new_net_5148_bfr_before (
		.din(new_net_5148),
		.dout(new_net_5147)
	);

	bfr new_net_5149_bfr_before (
		.din(new_net_5149),
		.dout(new_net_5148)
	);

	bfr new_net_5150_bfr_before (
		.din(new_net_5150),
		.dout(new_net_5149)
	);

	bfr new_net_5151_bfr_before (
		.din(new_net_5151),
		.dout(new_net_5150)
	);

	bfr new_net_5152_bfr_before (
		.din(new_net_5152),
		.dout(new_net_5151)
	);

	bfr new_net_5153_bfr_before (
		.din(new_net_5153),
		.dout(new_net_5152)
	);

	bfr new_net_5154_bfr_before (
		.din(new_net_5154),
		.dout(new_net_5153)
	);

	bfr new_net_5155_bfr_before (
		.din(new_net_5155),
		.dout(new_net_5154)
	);

	bfr new_net_5156_bfr_before (
		.din(new_net_5156),
		.dout(new_net_5155)
	);

	bfr new_net_5157_bfr_before (
		.din(new_net_5157),
		.dout(new_net_5156)
	);

	spl4L n_1308__v_fanout (
		.a(n_1308_),
		.b(new_net_699),
		.c(new_net_5157),
		.d(new_net_701),
		.e(new_net_698)
	);

	bfr new_net_5158_bfr_before (
		.din(new_net_5158),
		.dout(new_net_1035)
	);

	spl2 n_0119__v_fanout (
		.a(n_0119_),
		.b(new_net_5158),
		.c(new_net_1034)
	);

	bfr new_net_5159_bfr_before (
		.din(new_net_5159),
		.dout(new_net_1717)
	);

	bfr new_net_5160_bfr_before (
		.din(new_net_5160),
		.dout(new_net_5159)
	);

	bfr new_net_5161_bfr_before (
		.din(new_net_5161),
		.dout(new_net_5160)
	);

	bfr new_net_5162_bfr_before (
		.din(new_net_5162),
		.dout(new_net_5161)
	);

	bfr new_net_5163_bfr_before (
		.din(new_net_5163),
		.dout(new_net_5162)
	);

	bfr new_net_5164_bfr_before (
		.din(new_net_5164),
		.dout(new_net_5163)
	);

	bfr new_net_5165_bfr_before (
		.din(new_net_5165),
		.dout(new_net_5164)
	);

	bfr new_net_5166_bfr_before (
		.din(new_net_5166),
		.dout(new_net_5165)
	);

	bfr new_net_5167_bfr_before (
		.din(new_net_5167),
		.dout(new_net_5166)
	);

	spl2 n_1342__v_fanout (
		.a(n_1342_),
		.b(new_net_1718),
		.c(new_net_5167)
	);

	bfr new_net_5168_bfr_before (
		.din(new_net_5168),
		.dout(new_net_1303)
	);

	bfr new_net_5169_bfr_before (
		.din(new_net_5169),
		.dout(new_net_5168)
	);

	bfr new_net_5170_bfr_before (
		.din(new_net_5170),
		.dout(new_net_5169)
	);

	bfr new_net_5171_bfr_before (
		.din(new_net_5171),
		.dout(new_net_5170)
	);

	bfr new_net_5172_bfr_before (
		.din(new_net_5172),
		.dout(new_net_5171)
	);

	bfr new_net_5173_bfr_before (
		.din(new_net_5173),
		.dout(new_net_5172)
	);

	bfr new_net_5174_bfr_before (
		.din(new_net_5174),
		.dout(new_net_5173)
	);

	bfr new_net_5175_bfr_before (
		.din(new_net_5175),
		.dout(new_net_5174)
	);

	bfr new_net_5176_bfr_before (
		.din(new_net_5176),
		.dout(new_net_5175)
	);

	bfr new_net_5177_bfr_before (
		.din(new_net_5177),
		.dout(new_net_5176)
	);

	bfr new_net_5178_bfr_before (
		.din(new_net_5178),
		.dout(new_net_5177)
	);

	spl2 n_1338__v_fanout (
		.a(n_1338_),
		.b(new_net_5178),
		.c(new_net_1302)
	);

	spl2 n_0315__v_fanout (
		.a(n_0315_),
		.b(new_net_1307),
		.c(new_net_1306)
	);

	spl4L n_1306__v_fanout (
		.a(n_1306_),
		.b(new_net_450),
		.c(new_net_449),
		.d(new_net_451),
		.e(new_net_448)
	);

	spl2 n_0685__v_fanout (
		.a(n_0685_),
		.b(new_net_510),
		.c(new_net_509)
	);

	bfr new_net_5179_bfr_before (
		.din(new_net_5179),
		.dout(new_net_1692)
	);

	bfr new_net_5180_bfr_before (
		.din(new_net_5180),
		.dout(new_net_5179)
	);

	bfr new_net_5181_bfr_before (
		.din(new_net_5181),
		.dout(new_net_5180)
	);

	bfr new_net_5182_bfr_before (
		.din(new_net_5182),
		.dout(new_net_5181)
	);

	bfr new_net_5183_bfr_before (
		.din(new_net_5183),
		.dout(new_net_5182)
	);

	bfr new_net_5184_bfr_before (
		.din(new_net_5184),
		.dout(new_net_5183)
	);

	bfr new_net_5185_bfr_before (
		.din(new_net_5185),
		.dout(new_net_5184)
	);

	bfr new_net_5186_bfr_before (
		.din(new_net_5186),
		.dout(new_net_5185)
	);

	bfr new_net_5187_bfr_before (
		.din(new_net_5187),
		.dout(new_net_5186)
	);

	bfr new_net_5188_bfr_before (
		.din(new_net_5188),
		.dout(new_net_5187)
	);

	bfr new_net_5189_bfr_before (
		.din(new_net_5189),
		.dout(new_net_5188)
	);

	bfr new_net_5190_bfr_before (
		.din(new_net_5190),
		.dout(new_net_5189)
	);

	bfr new_net_5191_bfr_before (
		.din(new_net_5191),
		.dout(new_net_5190)
	);

	bfr new_net_5192_bfr_before (
		.din(new_net_5192),
		.dout(new_net_5191)
	);

	bfr new_net_5193_bfr_before (
		.din(new_net_5193),
		.dout(new_net_5192)
	);

	spl2 n_0044__v_fanout (
		.a(n_0044_),
		.b(new_net_1693),
		.c(new_net_5193)
	);

	bfr new_net_5194_bfr_after (
		.din(n_0792_),
		.dout(new_net_5194)
	);

	bfr new_net_5195_bfr_after (
		.din(new_net_5194),
		.dout(new_net_5195)
	);

	spl2 n_0792__v_fanout (
		.a(new_net_5195),
		.b(new_net_1633),
		.c(new_net_1632)
	);

	bfr new_net_5196_bfr_after (
		.din(n_1143_),
		.dout(new_net_5196)
	);

	bfr new_net_5197_bfr_after (
		.din(new_net_5196),
		.dout(new_net_5197)
	);

	spl2 n_1143__v_fanout (
		.a(new_net_5197),
		.b(new_net_1550),
		.c(new_net_1549)
	);

	bfr new_net_5198_bfr_before (
		.din(new_net_5198),
		.dout(new_net_1201)
	);

	bfr new_net_5199_bfr_before (
		.din(new_net_5199),
		.dout(new_net_5198)
	);

	spl2 n_0268__v_fanout (
		.a(n_0268_),
		.b(new_net_5199),
		.c(new_net_1200)
	);

	bfr new_net_5200_bfr_after (
		.din(n_1122_),
		.dout(new_net_5200)
	);

	bfr new_net_5201_bfr_after (
		.din(new_net_5200),
		.dout(new_net_5201)
	);

	spl2 n_1122__v_fanout (
		.a(new_net_5201),
		.b(new_net_627),
		.c(new_net_626)
	);

	bfr new_net_5202_bfr_before (
		.din(new_net_5202),
		.dout(new_net_940)
	);

	bfr new_net_5203_bfr_before (
		.din(new_net_5203),
		.dout(new_net_5202)
	);

	bfr new_net_5204_bfr_before (
		.din(new_net_5204),
		.dout(new_net_5203)
	);

	bfr new_net_5205_bfr_before (
		.din(new_net_5205),
		.dout(new_net_5204)
	);

	bfr new_net_5206_bfr_before (
		.din(new_net_5206),
		.dout(new_net_5205)
	);

	bfr new_net_5207_bfr_before (
		.din(new_net_5207),
		.dout(new_net_5206)
	);

	bfr new_net_5208_bfr_before (
		.din(new_net_5208),
		.dout(new_net_5207)
	);

	bfr new_net_5209_bfr_before (
		.din(new_net_5209),
		.dout(new_net_5208)
	);

	bfr new_net_5210_bfr_before (
		.din(new_net_5210),
		.dout(new_net_5209)
	);

	bfr new_net_5211_bfr_before (
		.din(new_net_5211),
		.dout(new_net_5210)
	);

	bfr new_net_5212_bfr_before (
		.din(new_net_5212),
		.dout(new_net_5211)
	);

	bfr new_net_5213_bfr_before (
		.din(new_net_5213),
		.dout(new_net_5212)
	);

	spl2 n_0045__v_fanout (
		.a(n_0045_),
		.b(new_net_941),
		.c(new_net_5213)
	);

	spl2 n_0022__v_fanout (
		.a(n_0022_),
		.b(new_net_407),
		.c(new_net_406)
	);

	bfr new_net_5214_bfr_before (
		.din(new_net_5214),
		.dout(N519)
	);

	bfr new_net_5215_bfr_before (
		.din(new_net_5215),
		.dout(new_net_5214)
	);

	bfr new_net_5216_bfr_before (
		.din(new_net_5216),
		.dout(new_net_5215)
	);

	bfr new_net_5217_bfr_before (
		.din(new_net_5217),
		.dout(new_net_5216)
	);

	bfr new_net_5218_bfr_before (
		.din(new_net_5218),
		.dout(new_net_5217)
	);

	bfr new_net_5219_bfr_before (
		.din(new_net_5219),
		.dout(new_net_5218)
	);

	bfr new_net_5220_bfr_before (
		.din(new_net_5220),
		.dout(new_net_5219)
	);

	bfr new_net_5221_bfr_before (
		.din(new_net_5221),
		.dout(new_net_5220)
	);

	bfr new_net_5222_bfr_before (
		.din(new_net_5222),
		.dout(new_net_5221)
	);

	bfr new_net_5223_bfr_before (
		.din(new_net_5223),
		.dout(new_net_5222)
	);

	bfr new_net_5224_bfr_before (
		.din(new_net_5224),
		.dout(new_net_5223)
	);

	bfr new_net_5225_bfr_before (
		.din(new_net_5225),
		.dout(new_net_5224)
	);

	bfr new_net_5226_bfr_before (
		.din(new_net_5226),
		.dout(new_net_5225)
	);

	bfr new_net_5227_bfr_before (
		.din(new_net_5227),
		.dout(new_net_5226)
	);

	bfr new_net_5228_bfr_before (
		.din(new_net_5228),
		.dout(new_net_5227)
	);

	bfr new_net_5229_bfr_before (
		.din(new_net_5229),
		.dout(new_net_5228)
	);

	bfr new_net_5230_bfr_before (
		.din(new_net_5230),
		.dout(new_net_5229)
	);

	bfr new_net_5231_bfr_before (
		.din(new_net_5231),
		.dout(new_net_5230)
	);

	bfr new_net_5232_bfr_before (
		.din(new_net_5232),
		.dout(new_net_5231)
	);

	bfr new_net_5233_bfr_before (
		.din(new_net_5233),
		.dout(new_net_5232)
	);

	bfr new_net_5234_bfr_before (
		.din(new_net_5234),
		.dout(new_net_5233)
	);

	bfr new_net_5235_bfr_before (
		.din(new_net_5235),
		.dout(new_net_5234)
	);

	bfr new_net_5236_bfr_before (
		.din(new_net_5236),
		.dout(new_net_5235)
	);

	bfr new_net_5237_bfr_before (
		.din(new_net_5237),
		.dout(new_net_5236)
	);

	bfr new_net_5238_bfr_before (
		.din(new_net_5238),
		.dout(new_net_5237)
	);

	bfr new_net_5239_bfr_before (
		.din(new_net_5239),
		.dout(new_net_5238)
	);

	bfr new_net_5240_bfr_before (
		.din(new_net_5240),
		.dout(new_net_5239)
	);

	bfr new_net_5241_bfr_before (
		.din(new_net_5241),
		.dout(new_net_5240)
	);

	bfr new_net_5242_bfr_before (
		.din(new_net_5242),
		.dout(new_net_5241)
	);

	bfr new_net_5243_bfr_before (
		.din(new_net_5243),
		.dout(new_net_5242)
	);

	bfr new_net_5244_bfr_before (
		.din(new_net_5244),
		.dout(new_net_5243)
	);

	bfr new_net_5245_bfr_before (
		.din(new_net_5245),
		.dout(new_net_5244)
	);

	bfr new_net_5246_bfr_before (
		.din(new_net_5246),
		.dout(new_net_5245)
	);

	bfr new_net_5247_bfr_before (
		.din(new_net_5247),
		.dout(new_net_5246)
	);

	bfr new_net_5248_bfr_before (
		.din(new_net_5248),
		.dout(new_net_5247)
	);

	bfr new_net_5249_bfr_before (
		.din(new_net_5249),
		.dout(new_net_5248)
	);

	bfr new_net_5250_bfr_before (
		.din(new_net_5250),
		.dout(new_net_5249)
	);

	bfr new_net_5251_bfr_before (
		.din(new_net_5251),
		.dout(new_net_5250)
	);

	bfr new_net_5252_bfr_before (
		.din(new_net_5252),
		.dout(new_net_5251)
	);

	bfr new_net_5253_bfr_before (
		.din(new_net_5253),
		.dout(new_net_5252)
	);

	bfr new_net_5254_bfr_before (
		.din(new_net_5254),
		.dout(new_net_5253)
	);

	bfr new_net_5255_bfr_before (
		.din(new_net_5255),
		.dout(new_net_5254)
	);

	bfr new_net_5256_bfr_before (
		.din(new_net_5256),
		.dout(new_net_5255)
	);

	bfr new_net_5257_bfr_before (
		.din(new_net_5257),
		.dout(new_net_5256)
	);

	bfr new_net_5258_bfr_before (
		.din(new_net_5258),
		.dout(new_net_5257)
	);

	bfr new_net_5259_bfr_before (
		.din(new_net_5259),
		.dout(new_net_5258)
	);

	bfr new_net_5260_bfr_before (
		.din(new_net_5260),
		.dout(new_net_5259)
	);

	bfr new_net_5261_bfr_before (
		.din(new_net_5261),
		.dout(new_net_5260)
	);

	bfr new_net_5262_bfr_before (
		.din(new_net_5262),
		.dout(new_net_5261)
	);

	bfr new_net_5263_bfr_before (
		.din(new_net_5263),
		.dout(new_net_5262)
	);

	bfr new_net_5264_bfr_before (
		.din(new_net_5264),
		.dout(new_net_5263)
	);

	bfr new_net_5265_bfr_before (
		.din(new_net_5265),
		.dout(new_net_5264)
	);

	bfr new_net_5266_bfr_before (
		.din(new_net_5266),
		.dout(new_net_5265)
	);

	bfr new_net_5267_bfr_before (
		.din(new_net_5267),
		.dout(new_net_5266)
	);

	bfr new_net_5268_bfr_before (
		.din(new_net_5268),
		.dout(new_net_5267)
	);

	bfr new_net_5269_bfr_before (
		.din(new_net_5269),
		.dout(new_net_5268)
	);

	bfr new_net_5270_bfr_before (
		.din(new_net_5270),
		.dout(new_net_5269)
	);

	bfr new_net_5271_bfr_before (
		.din(new_net_5271),
		.dout(new_net_5270)
	);

	spl3L new_net_2034_v_fanout (
		.a(new_net_2034),
		.b(new_net_5271),
		.c(new_net_1269),
		.d(new_net_1268)
	);

	spl4L n_0860__v_fanout (
		.a(n_0860_),
		.b(new_net_883),
		.c(new_net_884),
		.d(new_net_882),
		.e(new_net_881)
	);

	spl2 new_net_2071_v_fanout (
		.a(new_net_2071),
		.b(new_net_1583),
		.c(new_net_1585)
	);

	bfr new_net_5272_bfr_before (
		.din(new_net_5272),
		.dout(N541)
	);

	bfr new_net_5273_bfr_before (
		.din(new_net_5273),
		.dout(new_net_5272)
	);

	bfr new_net_5274_bfr_before (
		.din(new_net_5274),
		.dout(new_net_5273)
	);

	bfr new_net_5275_bfr_before (
		.din(new_net_5275),
		.dout(new_net_5274)
	);

	bfr new_net_5276_bfr_before (
		.din(new_net_5276),
		.dout(new_net_5275)
	);

	bfr new_net_5277_bfr_before (
		.din(new_net_5277),
		.dout(new_net_5276)
	);

	bfr new_net_5278_bfr_before (
		.din(new_net_5278),
		.dout(new_net_5277)
	);

	bfr new_net_5279_bfr_before (
		.din(new_net_5279),
		.dout(new_net_5278)
	);

	bfr new_net_5280_bfr_before (
		.din(new_net_5280),
		.dout(new_net_5279)
	);

	bfr new_net_5281_bfr_before (
		.din(new_net_5281),
		.dout(new_net_5280)
	);

	bfr new_net_5282_bfr_before (
		.din(new_net_5282),
		.dout(new_net_5281)
	);

	bfr new_net_5283_bfr_before (
		.din(new_net_5283),
		.dout(new_net_5282)
	);

	bfr new_net_5284_bfr_before (
		.din(new_net_5284),
		.dout(new_net_5283)
	);

	bfr new_net_5285_bfr_before (
		.din(new_net_5285),
		.dout(new_net_5284)
	);

	bfr new_net_5286_bfr_before (
		.din(new_net_5286),
		.dout(new_net_5285)
	);

	bfr new_net_5287_bfr_before (
		.din(new_net_5287),
		.dout(new_net_5286)
	);

	bfr new_net_5288_bfr_before (
		.din(new_net_5288),
		.dout(new_net_5287)
	);

	bfr new_net_5289_bfr_before (
		.din(new_net_5289),
		.dout(new_net_5288)
	);

	bfr new_net_5290_bfr_before (
		.din(new_net_5290),
		.dout(new_net_5289)
	);

	bfr new_net_5291_bfr_before (
		.din(new_net_5291),
		.dout(new_net_5290)
	);

	bfr new_net_5292_bfr_before (
		.din(new_net_5292),
		.dout(new_net_5291)
	);

	bfr new_net_5293_bfr_before (
		.din(new_net_5293),
		.dout(new_net_5292)
	);

	bfr new_net_5294_bfr_before (
		.din(new_net_5294),
		.dout(new_net_5293)
	);

	bfr new_net_5295_bfr_before (
		.din(new_net_5295),
		.dout(new_net_5294)
	);

	bfr new_net_5296_bfr_before (
		.din(new_net_5296),
		.dout(new_net_5295)
	);

	bfr new_net_5297_bfr_before (
		.din(new_net_5297),
		.dout(new_net_5296)
	);

	bfr new_net_5298_bfr_before (
		.din(new_net_5298),
		.dout(new_net_5297)
	);

	bfr new_net_5299_bfr_before (
		.din(new_net_5299),
		.dout(new_net_5298)
	);

	bfr new_net_5300_bfr_before (
		.din(new_net_5300),
		.dout(new_net_5299)
	);

	bfr new_net_5301_bfr_before (
		.din(new_net_5301),
		.dout(new_net_5300)
	);

	bfr new_net_5302_bfr_before (
		.din(new_net_5302),
		.dout(new_net_5301)
	);

	bfr new_net_5303_bfr_before (
		.din(new_net_5303),
		.dout(new_net_5302)
	);

	bfr new_net_5304_bfr_before (
		.din(new_net_5304),
		.dout(new_net_5303)
	);

	bfr new_net_5305_bfr_before (
		.din(new_net_5305),
		.dout(new_net_5304)
	);

	bfr new_net_5306_bfr_before (
		.din(new_net_5306),
		.dout(new_net_5305)
	);

	bfr new_net_5307_bfr_before (
		.din(new_net_5307),
		.dout(new_net_5306)
	);

	bfr new_net_5308_bfr_before (
		.din(new_net_5308),
		.dout(new_net_5307)
	);

	bfr new_net_5309_bfr_before (
		.din(new_net_5309),
		.dout(new_net_5308)
	);

	bfr new_net_5310_bfr_before (
		.din(new_net_5310),
		.dout(new_net_5309)
	);

	bfr new_net_5311_bfr_before (
		.din(new_net_5311),
		.dout(new_net_5310)
	);

	bfr new_net_5312_bfr_before (
		.din(new_net_5312),
		.dout(new_net_5311)
	);

	bfr new_net_5313_bfr_before (
		.din(new_net_5313),
		.dout(new_net_5312)
	);

	bfr new_net_5314_bfr_before (
		.din(new_net_5314),
		.dout(new_net_5313)
	);

	bfr new_net_5315_bfr_before (
		.din(new_net_5315),
		.dout(new_net_5314)
	);

	bfr new_net_5316_bfr_before (
		.din(new_net_5316),
		.dout(new_net_5315)
	);

	bfr new_net_5317_bfr_before (
		.din(new_net_5317),
		.dout(new_net_5316)
	);

	bfr new_net_5318_bfr_before (
		.din(new_net_5318),
		.dout(new_net_5317)
	);

	bfr new_net_5319_bfr_before (
		.din(new_net_5319),
		.dout(new_net_5318)
	);

	bfr new_net_5320_bfr_before (
		.din(new_net_5320),
		.dout(new_net_5319)
	);

	bfr new_net_5321_bfr_before (
		.din(new_net_5321),
		.dout(new_net_5320)
	);

	bfr new_net_5322_bfr_before (
		.din(new_net_5322),
		.dout(new_net_5321)
	);

	bfr new_net_5323_bfr_before (
		.din(new_net_5323),
		.dout(new_net_5322)
	);

	bfr new_net_5324_bfr_before (
		.din(new_net_5324),
		.dout(new_net_5323)
	);

	bfr new_net_5325_bfr_before (
		.din(new_net_5325),
		.dout(new_net_5324)
	);

	bfr new_net_5326_bfr_before (
		.din(new_net_5326),
		.dout(new_net_5325)
	);

	bfr new_net_5327_bfr_before (
		.din(new_net_5327),
		.dout(new_net_5326)
	);

	bfr new_net_5328_bfr_before (
		.din(new_net_5328),
		.dout(new_net_5327)
	);

	bfr new_net_5329_bfr_before (
		.din(new_net_5329),
		.dout(new_net_5328)
	);

	spl3L new_net_2038_v_fanout (
		.a(new_net_2038),
		.b(new_net_1356),
		.c(new_net_1354),
		.d(new_net_5329)
	);

	bfr new_net_5330_bfr_before (
		.din(new_net_5330),
		.dout(N482)
	);

	bfr new_net_5331_bfr_before (
		.din(new_net_5331),
		.dout(new_net_5330)
	);

	bfr new_net_5332_bfr_before (
		.din(new_net_5332),
		.dout(new_net_5331)
	);

	bfr new_net_5333_bfr_before (
		.din(new_net_5333),
		.dout(new_net_5332)
	);

	bfr new_net_5334_bfr_before (
		.din(new_net_5334),
		.dout(new_net_5333)
	);

	bfr new_net_5335_bfr_before (
		.din(new_net_5335),
		.dout(new_net_5334)
	);

	bfr new_net_5336_bfr_before (
		.din(new_net_5336),
		.dout(new_net_5335)
	);

	bfr new_net_5337_bfr_before (
		.din(new_net_5337),
		.dout(new_net_5336)
	);

	bfr new_net_5338_bfr_before (
		.din(new_net_5338),
		.dout(new_net_5337)
	);

	bfr new_net_5339_bfr_before (
		.din(new_net_5339),
		.dout(new_net_5338)
	);

	bfr new_net_5340_bfr_before (
		.din(new_net_5340),
		.dout(new_net_5339)
	);

	bfr new_net_5341_bfr_before (
		.din(new_net_5341),
		.dout(new_net_5340)
	);

	bfr new_net_5342_bfr_before (
		.din(new_net_5342),
		.dout(new_net_5341)
	);

	bfr new_net_5343_bfr_before (
		.din(new_net_5343),
		.dout(new_net_5342)
	);

	bfr new_net_5344_bfr_before (
		.din(new_net_5344),
		.dout(new_net_5343)
	);

	bfr new_net_5345_bfr_before (
		.din(new_net_5345),
		.dout(new_net_5344)
	);

	bfr new_net_5346_bfr_before (
		.din(new_net_5346),
		.dout(new_net_5345)
	);

	bfr new_net_5347_bfr_before (
		.din(new_net_5347),
		.dout(new_net_5346)
	);

	bfr new_net_5348_bfr_before (
		.din(new_net_5348),
		.dout(new_net_5347)
	);

	bfr new_net_5349_bfr_before (
		.din(new_net_5349),
		.dout(new_net_5348)
	);

	bfr new_net_5350_bfr_before (
		.din(new_net_5350),
		.dout(new_net_5349)
	);

	bfr new_net_5351_bfr_before (
		.din(new_net_5351),
		.dout(new_net_5350)
	);

	bfr new_net_5352_bfr_before (
		.din(new_net_5352),
		.dout(new_net_5351)
	);

	bfr new_net_5353_bfr_before (
		.din(new_net_5353),
		.dout(new_net_5352)
	);

	bfr new_net_5354_bfr_before (
		.din(new_net_5354),
		.dout(new_net_5353)
	);

	bfr new_net_5355_bfr_before (
		.din(new_net_5355),
		.dout(new_net_5354)
	);

	bfr new_net_5356_bfr_before (
		.din(new_net_5356),
		.dout(new_net_5355)
	);

	bfr new_net_5357_bfr_before (
		.din(new_net_5357),
		.dout(new_net_5356)
	);

	bfr new_net_5358_bfr_before (
		.din(new_net_5358),
		.dout(new_net_5357)
	);

	bfr new_net_5359_bfr_before (
		.din(new_net_5359),
		.dout(new_net_5358)
	);

	bfr new_net_5360_bfr_before (
		.din(new_net_5360),
		.dout(new_net_5359)
	);

	bfr new_net_5361_bfr_before (
		.din(new_net_5361),
		.dout(new_net_5360)
	);

	bfr new_net_5362_bfr_before (
		.din(new_net_5362),
		.dout(new_net_5361)
	);

	bfr new_net_5363_bfr_before (
		.din(new_net_5363),
		.dout(new_net_5362)
	);

	bfr new_net_5364_bfr_before (
		.din(new_net_5364),
		.dout(new_net_5363)
	);

	bfr new_net_5365_bfr_before (
		.din(new_net_5365),
		.dout(new_net_5364)
	);

	bfr new_net_5366_bfr_before (
		.din(new_net_5366),
		.dout(new_net_5365)
	);

	bfr new_net_5367_bfr_before (
		.din(new_net_5367),
		.dout(new_net_5366)
	);

	bfr new_net_5368_bfr_before (
		.din(new_net_5368),
		.dout(new_net_5367)
	);

	bfr new_net_5369_bfr_before (
		.din(new_net_5369),
		.dout(new_net_5368)
	);

	bfr new_net_5370_bfr_before (
		.din(new_net_5370),
		.dout(new_net_5369)
	);

	bfr new_net_5371_bfr_before (
		.din(new_net_5371),
		.dout(new_net_5370)
	);

	bfr new_net_5372_bfr_before (
		.din(new_net_5372),
		.dout(new_net_5371)
	);

	bfr new_net_5373_bfr_before (
		.din(new_net_5373),
		.dout(new_net_5372)
	);

	bfr new_net_5374_bfr_before (
		.din(new_net_5374),
		.dout(new_net_5373)
	);

	bfr new_net_5375_bfr_before (
		.din(new_net_5375),
		.dout(new_net_5374)
	);

	bfr new_net_5376_bfr_before (
		.din(new_net_5376),
		.dout(new_net_5375)
	);

	bfr new_net_5377_bfr_before (
		.din(new_net_5377),
		.dout(new_net_5376)
	);

	bfr new_net_5378_bfr_before (
		.din(new_net_5378),
		.dout(new_net_5377)
	);

	bfr new_net_5379_bfr_before (
		.din(new_net_5379),
		.dout(new_net_5378)
	);

	bfr new_net_5380_bfr_before (
		.din(new_net_5380),
		.dout(new_net_5379)
	);

	bfr new_net_5381_bfr_before (
		.din(new_net_5381),
		.dout(new_net_5380)
	);

	bfr new_net_5382_bfr_before (
		.din(new_net_5382),
		.dout(new_net_5381)
	);

	bfr new_net_5383_bfr_before (
		.din(new_net_5383),
		.dout(new_net_5382)
	);

	bfr new_net_5384_bfr_before (
		.din(new_net_5384),
		.dout(new_net_5383)
	);

	bfr new_net_5385_bfr_before (
		.din(new_net_5385),
		.dout(new_net_5384)
	);

	bfr new_net_5386_bfr_before (
		.din(new_net_5386),
		.dout(new_net_5385)
	);

	bfr new_net_5387_bfr_before (
		.din(new_net_5387),
		.dout(new_net_5386)
	);

	spl3L new_net_2022_v_fanout (
		.a(new_net_2022),
		.b(new_net_5387),
		.c(new_net_1072),
		.d(new_net_1070)
	);

	bfr new_net_5388_bfr_before (
		.din(new_net_5388),
		.dout(N563)
	);

	bfr new_net_5389_bfr_before (
		.din(new_net_5389),
		.dout(new_net_5388)
	);

	bfr new_net_5390_bfr_before (
		.din(new_net_5390),
		.dout(new_net_5389)
	);

	bfr new_net_5391_bfr_before (
		.din(new_net_5391),
		.dout(new_net_5390)
	);

	bfr new_net_5392_bfr_before (
		.din(new_net_5392),
		.dout(new_net_5391)
	);

	bfr new_net_5393_bfr_before (
		.din(new_net_5393),
		.dout(new_net_5392)
	);

	bfr new_net_5394_bfr_before (
		.din(new_net_5394),
		.dout(new_net_5393)
	);

	bfr new_net_5395_bfr_before (
		.din(new_net_5395),
		.dout(new_net_5394)
	);

	bfr new_net_5396_bfr_before (
		.din(new_net_5396),
		.dout(new_net_5395)
	);

	bfr new_net_5397_bfr_before (
		.din(new_net_5397),
		.dout(new_net_5396)
	);

	bfr new_net_5398_bfr_before (
		.din(new_net_5398),
		.dout(new_net_5397)
	);

	bfr new_net_5399_bfr_before (
		.din(new_net_5399),
		.dout(new_net_5398)
	);

	bfr new_net_5400_bfr_before (
		.din(new_net_5400),
		.dout(new_net_5399)
	);

	bfr new_net_5401_bfr_before (
		.din(new_net_5401),
		.dout(new_net_5400)
	);

	bfr new_net_5402_bfr_before (
		.din(new_net_5402),
		.dout(new_net_5401)
	);

	bfr new_net_5403_bfr_before (
		.din(new_net_5403),
		.dout(new_net_5402)
	);

	bfr new_net_5404_bfr_before (
		.din(new_net_5404),
		.dout(new_net_5403)
	);

	bfr new_net_5405_bfr_before (
		.din(new_net_5405),
		.dout(new_net_5404)
	);

	bfr new_net_5406_bfr_before (
		.din(new_net_5406),
		.dout(new_net_5405)
	);

	bfr new_net_5407_bfr_before (
		.din(new_net_5407),
		.dout(new_net_5406)
	);

	bfr new_net_5408_bfr_before (
		.din(new_net_5408),
		.dout(new_net_5407)
	);

	bfr new_net_5409_bfr_before (
		.din(new_net_5409),
		.dout(new_net_5408)
	);

	bfr new_net_5410_bfr_before (
		.din(new_net_5410),
		.dout(new_net_5409)
	);

	bfr new_net_5411_bfr_before (
		.din(new_net_5411),
		.dout(new_net_5410)
	);

	bfr new_net_5412_bfr_before (
		.din(new_net_5412),
		.dout(new_net_5411)
	);

	bfr new_net_5413_bfr_before (
		.din(new_net_5413),
		.dout(new_net_5412)
	);

	bfr new_net_5414_bfr_before (
		.din(new_net_5414),
		.dout(new_net_5413)
	);

	bfr new_net_5415_bfr_before (
		.din(new_net_5415),
		.dout(new_net_5414)
	);

	bfr new_net_5416_bfr_before (
		.din(new_net_5416),
		.dout(new_net_5415)
	);

	bfr new_net_5417_bfr_before (
		.din(new_net_5417),
		.dout(new_net_5416)
	);

	bfr new_net_5418_bfr_before (
		.din(new_net_5418),
		.dout(new_net_5417)
	);

	bfr new_net_5419_bfr_before (
		.din(new_net_5419),
		.dout(new_net_5418)
	);

	bfr new_net_5420_bfr_before (
		.din(new_net_5420),
		.dout(new_net_5419)
	);

	bfr new_net_5421_bfr_before (
		.din(new_net_5421),
		.dout(new_net_5420)
	);

	bfr new_net_5422_bfr_before (
		.din(new_net_5422),
		.dout(new_net_5421)
	);

	bfr new_net_5423_bfr_before (
		.din(new_net_5423),
		.dout(new_net_5422)
	);

	bfr new_net_5424_bfr_before (
		.din(new_net_5424),
		.dout(new_net_5423)
	);

	bfr new_net_5425_bfr_before (
		.din(new_net_5425),
		.dout(new_net_5424)
	);

	bfr new_net_5426_bfr_before (
		.din(new_net_5426),
		.dout(new_net_5425)
	);

	bfr new_net_5427_bfr_before (
		.din(new_net_5427),
		.dout(new_net_5426)
	);

	bfr new_net_5428_bfr_before (
		.din(new_net_5428),
		.dout(new_net_5427)
	);

	bfr new_net_5429_bfr_before (
		.din(new_net_5429),
		.dout(new_net_5428)
	);

	bfr new_net_5430_bfr_before (
		.din(new_net_5430),
		.dout(new_net_5429)
	);

	bfr new_net_5431_bfr_before (
		.din(new_net_5431),
		.dout(new_net_5430)
	);

	bfr new_net_5432_bfr_before (
		.din(new_net_5432),
		.dout(new_net_5431)
	);

	bfr new_net_5433_bfr_before (
		.din(new_net_5433),
		.dout(new_net_5432)
	);

	bfr new_net_5434_bfr_before (
		.din(new_net_5434),
		.dout(new_net_5433)
	);

	bfr new_net_5435_bfr_before (
		.din(new_net_5435),
		.dout(new_net_5434)
	);

	bfr new_net_5436_bfr_before (
		.din(new_net_5436),
		.dout(new_net_5435)
	);

	bfr new_net_5437_bfr_before (
		.din(new_net_5437),
		.dout(new_net_5436)
	);

	bfr new_net_5438_bfr_before (
		.din(new_net_5438),
		.dout(new_net_5437)
	);

	bfr new_net_5439_bfr_before (
		.din(new_net_5439),
		.dout(new_net_5438)
	);

	bfr new_net_5440_bfr_before (
		.din(new_net_5440),
		.dout(new_net_5439)
	);

	bfr new_net_5441_bfr_before (
		.din(new_net_5441),
		.dout(new_net_5440)
	);

	bfr new_net_5442_bfr_before (
		.din(new_net_5442),
		.dout(new_net_5441)
	);

	bfr new_net_5443_bfr_before (
		.din(new_net_5443),
		.dout(new_net_5442)
	);

	bfr new_net_5444_bfr_before (
		.din(new_net_5444),
		.dout(new_net_5443)
	);

	bfr new_net_5445_bfr_before (
		.din(new_net_5445),
		.dout(new_net_5444)
	);

	spl3L new_net_2048_v_fanout (
		.a(new_net_2048),
		.b(new_net_1610),
		.c(new_net_1608),
		.d(new_net_5445)
	);

	bfr new_net_5446_bfr_before (
		.din(new_net_5446),
		.dout(N643)
	);

	bfr new_net_5447_bfr_before (
		.din(new_net_5447),
		.dout(new_net_5446)
	);

	bfr new_net_5448_bfr_before (
		.din(new_net_5448),
		.dout(new_net_5447)
	);

	bfr new_net_5449_bfr_before (
		.din(new_net_5449),
		.dout(new_net_5448)
	);

	bfr new_net_5450_bfr_before (
		.din(new_net_5450),
		.dout(new_net_5449)
	);

	bfr new_net_5451_bfr_before (
		.din(new_net_5451),
		.dout(new_net_5450)
	);

	bfr new_net_5452_bfr_before (
		.din(new_net_5452),
		.dout(new_net_5451)
	);

	bfr new_net_5453_bfr_before (
		.din(new_net_5453),
		.dout(new_net_5452)
	);

	bfr new_net_5454_bfr_before (
		.din(new_net_5454),
		.dout(new_net_5453)
	);

	bfr new_net_5455_bfr_before (
		.din(new_net_5455),
		.dout(new_net_5454)
	);

	bfr new_net_5456_bfr_before (
		.din(new_net_5456),
		.dout(new_net_5455)
	);

	bfr new_net_5457_bfr_before (
		.din(new_net_5457),
		.dout(new_net_5456)
	);

	bfr new_net_5458_bfr_before (
		.din(new_net_5458),
		.dout(new_net_5457)
	);

	bfr new_net_5459_bfr_before (
		.din(new_net_5459),
		.dout(new_net_5458)
	);

	bfr new_net_5460_bfr_before (
		.din(new_net_5460),
		.dout(new_net_5459)
	);

	bfr new_net_5461_bfr_before (
		.din(new_net_5461),
		.dout(new_net_5460)
	);

	bfr new_net_5462_bfr_before (
		.din(new_net_5462),
		.dout(new_net_5461)
	);

	bfr new_net_5463_bfr_before (
		.din(new_net_5463),
		.dout(new_net_5462)
	);

	bfr new_net_5464_bfr_before (
		.din(new_net_5464),
		.dout(new_net_5463)
	);

	bfr new_net_5465_bfr_before (
		.din(new_net_5465),
		.dout(new_net_5464)
	);

	bfr new_net_5466_bfr_before (
		.din(new_net_5466),
		.dout(new_net_5465)
	);

	bfr new_net_5467_bfr_before (
		.din(new_net_5467),
		.dout(new_net_5466)
	);

	bfr new_net_5468_bfr_before (
		.din(new_net_5468),
		.dout(new_net_5467)
	);

	bfr new_net_5469_bfr_before (
		.din(new_net_5469),
		.dout(new_net_5468)
	);

	bfr new_net_5470_bfr_before (
		.din(new_net_5470),
		.dout(new_net_5469)
	);

	bfr new_net_5471_bfr_before (
		.din(new_net_5471),
		.dout(new_net_5470)
	);

	bfr new_net_5472_bfr_before (
		.din(new_net_5472),
		.dout(new_net_5471)
	);

	bfr new_net_5473_bfr_before (
		.din(new_net_5473),
		.dout(new_net_5472)
	);

	bfr new_net_5474_bfr_before (
		.din(new_net_5474),
		.dout(new_net_5473)
	);

	bfr new_net_5475_bfr_before (
		.din(new_net_5475),
		.dout(new_net_5474)
	);

	bfr new_net_5476_bfr_before (
		.din(new_net_5476),
		.dout(new_net_5475)
	);

	bfr new_net_5477_bfr_before (
		.din(new_net_5477),
		.dout(new_net_5476)
	);

	bfr new_net_5478_bfr_before (
		.din(new_net_5478),
		.dout(new_net_5477)
	);

	bfr new_net_5479_bfr_before (
		.din(new_net_5479),
		.dout(new_net_5478)
	);

	bfr new_net_5480_bfr_before (
		.din(new_net_5480),
		.dout(new_net_5479)
	);

	bfr new_net_5481_bfr_before (
		.din(new_net_5481),
		.dout(new_net_5480)
	);

	bfr new_net_5482_bfr_before (
		.din(new_net_5482),
		.dout(new_net_5481)
	);

	bfr new_net_5483_bfr_before (
		.din(new_net_5483),
		.dout(new_net_5482)
	);

	bfr new_net_5484_bfr_before (
		.din(new_net_5484),
		.dout(new_net_5483)
	);

	bfr new_net_5485_bfr_before (
		.din(new_net_5485),
		.dout(new_net_5484)
	);

	bfr new_net_5486_bfr_before (
		.din(new_net_5486),
		.dout(new_net_5485)
	);

	bfr new_net_5487_bfr_before (
		.din(new_net_5487),
		.dout(new_net_5486)
	);

	bfr new_net_5488_bfr_before (
		.din(new_net_5488),
		.dout(new_net_5487)
	);

	bfr new_net_5489_bfr_before (
		.din(new_net_5489),
		.dout(new_net_5488)
	);

	bfr new_net_5490_bfr_before (
		.din(new_net_5490),
		.dout(new_net_5489)
	);

	bfr new_net_5491_bfr_before (
		.din(new_net_5491),
		.dout(new_net_5490)
	);

	bfr new_net_5492_bfr_before (
		.din(new_net_5492),
		.dout(new_net_5491)
	);

	bfr new_net_5493_bfr_before (
		.din(new_net_5493),
		.dout(new_net_5492)
	);

	bfr new_net_5494_bfr_before (
		.din(new_net_5494),
		.dout(new_net_5493)
	);

	bfr new_net_5495_bfr_before (
		.din(new_net_5495),
		.dout(new_net_5494)
	);

	bfr new_net_5496_bfr_before (
		.din(new_net_5496),
		.dout(new_net_5495)
	);

	bfr new_net_5497_bfr_before (
		.din(new_net_5497),
		.dout(new_net_5496)
	);

	bfr new_net_5498_bfr_before (
		.din(new_net_5498),
		.dout(new_net_5497)
	);

	bfr new_net_5499_bfr_before (
		.din(new_net_5499),
		.dout(new_net_5498)
	);

	bfr new_net_5500_bfr_before (
		.din(new_net_5500),
		.dout(new_net_5499)
	);

	bfr new_net_5501_bfr_before (
		.din(new_net_5501),
		.dout(new_net_5500)
	);

	bfr new_net_5502_bfr_before (
		.din(new_net_5502),
		.dout(new_net_5501)
	);

	bfr new_net_5503_bfr_before (
		.din(new_net_5503),
		.dout(new_net_5502)
	);

	spl3L new_net_2021_v_fanout (
		.a(new_net_2021),
		.b(new_net_5503),
		.c(new_net_949),
		.d(new_net_948)
	);

	spl4L n_0857__v_fanout (
		.a(n_0857_),
		.b(new_net_566),
		.c(new_net_564),
		.d(new_net_565),
		.e(new_net_563)
	);

	spl2 n_0869__v_fanout (
		.a(n_0869_),
		.b(new_net_599),
		.c(new_net_598)
	);

	bfr new_net_5504_bfr_before (
		.din(new_net_5504),
		.dout(N517)
	);

	bfr new_net_5505_bfr_before (
		.din(new_net_5505),
		.dout(new_net_5504)
	);

	bfr new_net_5506_bfr_before (
		.din(new_net_5506),
		.dout(new_net_5505)
	);

	bfr new_net_5507_bfr_before (
		.din(new_net_5507),
		.dout(new_net_5506)
	);

	bfr new_net_5508_bfr_before (
		.din(new_net_5508),
		.dout(new_net_5507)
	);

	bfr new_net_5509_bfr_before (
		.din(new_net_5509),
		.dout(new_net_5508)
	);

	bfr new_net_5510_bfr_before (
		.din(new_net_5510),
		.dout(new_net_5509)
	);

	bfr new_net_5511_bfr_before (
		.din(new_net_5511),
		.dout(new_net_5510)
	);

	bfr new_net_5512_bfr_before (
		.din(new_net_5512),
		.dout(new_net_5511)
	);

	bfr new_net_5513_bfr_before (
		.din(new_net_5513),
		.dout(new_net_5512)
	);

	bfr new_net_5514_bfr_before (
		.din(new_net_5514),
		.dout(new_net_5513)
	);

	bfr new_net_5515_bfr_before (
		.din(new_net_5515),
		.dout(new_net_5514)
	);

	bfr new_net_5516_bfr_before (
		.din(new_net_5516),
		.dout(new_net_5515)
	);

	bfr new_net_5517_bfr_before (
		.din(new_net_5517),
		.dout(new_net_5516)
	);

	bfr new_net_5518_bfr_before (
		.din(new_net_5518),
		.dout(new_net_5517)
	);

	bfr new_net_5519_bfr_before (
		.din(new_net_5519),
		.dout(new_net_5518)
	);

	bfr new_net_5520_bfr_before (
		.din(new_net_5520),
		.dout(new_net_5519)
	);

	bfr new_net_5521_bfr_before (
		.din(new_net_5521),
		.dout(new_net_5520)
	);

	bfr new_net_5522_bfr_before (
		.din(new_net_5522),
		.dout(new_net_5521)
	);

	bfr new_net_5523_bfr_before (
		.din(new_net_5523),
		.dout(new_net_5522)
	);

	bfr new_net_5524_bfr_before (
		.din(new_net_5524),
		.dout(new_net_5523)
	);

	bfr new_net_5525_bfr_before (
		.din(new_net_5525),
		.dout(new_net_5524)
	);

	bfr new_net_5526_bfr_before (
		.din(new_net_5526),
		.dout(new_net_5525)
	);

	bfr new_net_5527_bfr_before (
		.din(new_net_5527),
		.dout(new_net_5526)
	);

	bfr new_net_5528_bfr_before (
		.din(new_net_5528),
		.dout(new_net_5527)
	);

	bfr new_net_5529_bfr_before (
		.din(new_net_5529),
		.dout(new_net_5528)
	);

	bfr new_net_5530_bfr_before (
		.din(new_net_5530),
		.dout(new_net_5529)
	);

	bfr new_net_5531_bfr_before (
		.din(new_net_5531),
		.dout(new_net_5530)
	);

	bfr new_net_5532_bfr_before (
		.din(new_net_5532),
		.dout(new_net_5531)
	);

	bfr new_net_5533_bfr_before (
		.din(new_net_5533),
		.dout(new_net_5532)
	);

	bfr new_net_5534_bfr_before (
		.din(new_net_5534),
		.dout(new_net_5533)
	);

	bfr new_net_5535_bfr_before (
		.din(new_net_5535),
		.dout(new_net_5534)
	);

	bfr new_net_5536_bfr_before (
		.din(new_net_5536),
		.dout(new_net_5535)
	);

	bfr new_net_5537_bfr_before (
		.din(new_net_5537),
		.dout(new_net_5536)
	);

	bfr new_net_5538_bfr_before (
		.din(new_net_5538),
		.dout(new_net_5537)
	);

	bfr new_net_5539_bfr_before (
		.din(new_net_5539),
		.dout(new_net_5538)
	);

	bfr new_net_5540_bfr_before (
		.din(new_net_5540),
		.dout(new_net_5539)
	);

	bfr new_net_5541_bfr_before (
		.din(new_net_5541),
		.dout(new_net_5540)
	);

	bfr new_net_5542_bfr_before (
		.din(new_net_5542),
		.dout(new_net_5541)
	);

	bfr new_net_5543_bfr_before (
		.din(new_net_5543),
		.dout(new_net_5542)
	);

	bfr new_net_5544_bfr_before (
		.din(new_net_5544),
		.dout(new_net_5543)
	);

	bfr new_net_5545_bfr_before (
		.din(new_net_5545),
		.dout(new_net_5544)
	);

	bfr new_net_5546_bfr_before (
		.din(new_net_5546),
		.dout(new_net_5545)
	);

	bfr new_net_5547_bfr_before (
		.din(new_net_5547),
		.dout(new_net_5546)
	);

	bfr new_net_5548_bfr_before (
		.din(new_net_5548),
		.dout(new_net_5547)
	);

	bfr new_net_5549_bfr_before (
		.din(new_net_5549),
		.dout(new_net_5548)
	);

	bfr new_net_5550_bfr_before (
		.din(new_net_5550),
		.dout(new_net_5549)
	);

	bfr new_net_5551_bfr_before (
		.din(new_net_5551),
		.dout(new_net_5550)
	);

	bfr new_net_5552_bfr_before (
		.din(new_net_5552),
		.dout(new_net_5551)
	);

	bfr new_net_5553_bfr_before (
		.din(new_net_5553),
		.dout(new_net_5552)
	);

	bfr new_net_5554_bfr_before (
		.din(new_net_5554),
		.dout(new_net_5553)
	);

	bfr new_net_5555_bfr_before (
		.din(new_net_5555),
		.dout(new_net_5554)
	);

	bfr new_net_5556_bfr_before (
		.din(new_net_5556),
		.dout(new_net_5555)
	);

	bfr new_net_5557_bfr_before (
		.din(new_net_5557),
		.dout(new_net_5556)
	);

	bfr new_net_5558_bfr_before (
		.din(new_net_5558),
		.dout(new_net_5557)
	);

	bfr new_net_5559_bfr_before (
		.din(new_net_5559),
		.dout(new_net_5558)
	);

	bfr new_net_5560_bfr_before (
		.din(new_net_5560),
		.dout(new_net_5559)
	);

	bfr new_net_5561_bfr_before (
		.din(new_net_5561),
		.dout(new_net_5560)
	);

	spl3L new_net_2033_v_fanout (
		.a(new_net_2033),
		.b(new_net_1236),
		.c(new_net_1234),
		.d(new_net_5561)
	);

	spl4L n_1233__v_fanout (
		.a(n_1233_),
		.b(new_net_96),
		.c(new_net_97),
		.d(new_net_95),
		.e(new_net_94)
	);

	spl3L n_1137__v_fanout (
		.a(n_1137_),
		.b(new_net_743),
		.c(new_net_741),
		.d(new_net_742)
	);

	spl2 new_net_2097_v_fanout (
		.a(new_net_2097),
		.b(new_net_640),
		.c(new_net_639)
	);

	spl2 new_net_2084_v_fanout (
		.a(new_net_2084),
		.b(new_net_976),
		.c(new_net_975)
	);

	spl2 new_net_2082_v_fanout (
		.a(new_net_2082),
		.b(new_net_42),
		.c(new_net_43)
	);

	spl2 new_net_2095_v_fanout (
		.a(new_net_2095),
		.b(new_net_981),
		.c(new_net_982)
	);

	spl4L n_1160__v_fanout (
		.a(n_1160_),
		.b(new_net_1554),
		.c(new_net_1552),
		.d(new_net_1553),
		.e(new_net_1551)
	);

	spl4L n_1178__v_fanout (
		.a(n_1178_),
		.b(new_net_1664),
		.c(new_net_1665),
		.d(new_net_1666),
		.e(new_net_1663)
	);

	spl4L n_1275__v_fanout (
		.a(n_1275_),
		.b(new_net_1181),
		.c(new_net_1179),
		.d(new_net_1180),
		.e(new_net_1178)
	);

	spl2 new_net_2070_v_fanout (
		.a(new_net_2070),
		.b(new_net_795),
		.c(new_net_793)
	);

	spl2 n_1185__v_fanout (
		.a(n_1185_),
		.b(new_net_1097),
		.c(new_net_1096)
	);

	spl4L n_0738__v_fanout (
		.a(n_0738_),
		.b(new_net_486),
		.c(new_net_487),
		.d(new_net_485),
		.e(new_net_484)
	);

	spl4L n_0827__v_fanout (
		.a(n_0827_),
		.b(new_net_1504),
		.c(new_net_1505),
		.d(new_net_1506),
		.e(new_net_1503)
	);

	spl4L n_1280__v_fanout (
		.a(n_1280_),
		.b(new_net_1293),
		.c(new_net_1291),
		.d(new_net_1292),
		.e(new_net_1290)
	);

	spl2 n_0735__v_fanout (
		.a(n_0735_),
		.b(new_net_616),
		.c(new_net_615)
	);

	spl4L n_0878__v_fanout (
		.a(n_0878_),
		.b(new_net_798),
		.c(new_net_799),
		.d(new_net_800),
		.e(new_net_797)
	);

	spl4L n_0851__v_fanout (
		.a(n_0851_),
		.b(new_net_38),
		.c(new_net_39),
		.d(new_net_40),
		.e(new_net_37)
	);

	spl2 n_0806__v_fanout (
		.a(n_0806_),
		.b(new_net_1938),
		.c(new_net_1937)
	);

	spl3L n_0772__v_fanout (
		.a(n_0772_),
		.b(new_net_1195),
		.c(new_net_1193),
		.d(new_net_1194)
	);

	bfr new_net_5562_bfr_before (
		.din(new_net_5562),
		.dout(N505)
	);

	bfr new_net_5563_bfr_before (
		.din(new_net_5563),
		.dout(new_net_5562)
	);

	bfr new_net_5564_bfr_before (
		.din(new_net_5564),
		.dout(new_net_5563)
	);

	bfr new_net_5565_bfr_before (
		.din(new_net_5565),
		.dout(new_net_5564)
	);

	bfr new_net_5566_bfr_before (
		.din(new_net_5566),
		.dout(new_net_5565)
	);

	bfr new_net_5567_bfr_before (
		.din(new_net_5567),
		.dout(new_net_5566)
	);

	bfr new_net_5568_bfr_before (
		.din(new_net_5568),
		.dout(new_net_5567)
	);

	bfr new_net_5569_bfr_before (
		.din(new_net_5569),
		.dout(new_net_5568)
	);

	bfr new_net_5570_bfr_before (
		.din(new_net_5570),
		.dout(new_net_5569)
	);

	bfr new_net_5571_bfr_before (
		.din(new_net_5571),
		.dout(new_net_5570)
	);

	bfr new_net_5572_bfr_before (
		.din(new_net_5572),
		.dout(new_net_5571)
	);

	bfr new_net_5573_bfr_before (
		.din(new_net_5573),
		.dout(new_net_5572)
	);

	bfr new_net_5574_bfr_before (
		.din(new_net_5574),
		.dout(new_net_5573)
	);

	bfr new_net_5575_bfr_before (
		.din(new_net_5575),
		.dout(new_net_5574)
	);

	bfr new_net_5576_bfr_before (
		.din(new_net_5576),
		.dout(new_net_5575)
	);

	bfr new_net_5577_bfr_before (
		.din(new_net_5577),
		.dout(new_net_5576)
	);

	bfr new_net_5578_bfr_before (
		.din(new_net_5578),
		.dout(new_net_5577)
	);

	bfr new_net_5579_bfr_before (
		.din(new_net_5579),
		.dout(new_net_5578)
	);

	bfr new_net_5580_bfr_before (
		.din(new_net_5580),
		.dout(new_net_5579)
	);

	bfr new_net_5581_bfr_before (
		.din(new_net_5581),
		.dout(new_net_5580)
	);

	bfr new_net_5582_bfr_before (
		.din(new_net_5582),
		.dout(new_net_5581)
	);

	bfr new_net_5583_bfr_before (
		.din(new_net_5583),
		.dout(new_net_5582)
	);

	bfr new_net_5584_bfr_before (
		.din(new_net_5584),
		.dout(new_net_5583)
	);

	bfr new_net_5585_bfr_before (
		.din(new_net_5585),
		.dout(new_net_5584)
	);

	bfr new_net_5586_bfr_before (
		.din(new_net_5586),
		.dout(new_net_5585)
	);

	bfr new_net_5587_bfr_before (
		.din(new_net_5587),
		.dout(new_net_5586)
	);

	bfr new_net_5588_bfr_before (
		.din(new_net_5588),
		.dout(new_net_5587)
	);

	bfr new_net_5589_bfr_before (
		.din(new_net_5589),
		.dout(new_net_5588)
	);

	bfr new_net_5590_bfr_before (
		.din(new_net_5590),
		.dout(new_net_5589)
	);

	bfr new_net_5591_bfr_before (
		.din(new_net_5591),
		.dout(new_net_5590)
	);

	bfr new_net_5592_bfr_before (
		.din(new_net_5592),
		.dout(new_net_5591)
	);

	bfr new_net_5593_bfr_before (
		.din(new_net_5593),
		.dout(new_net_5592)
	);

	bfr new_net_5594_bfr_before (
		.din(new_net_5594),
		.dout(new_net_5593)
	);

	bfr new_net_5595_bfr_before (
		.din(new_net_5595),
		.dout(new_net_5594)
	);

	bfr new_net_5596_bfr_before (
		.din(new_net_5596),
		.dout(new_net_5595)
	);

	bfr new_net_5597_bfr_before (
		.din(new_net_5597),
		.dout(new_net_5596)
	);

	bfr new_net_5598_bfr_before (
		.din(new_net_5598),
		.dout(new_net_5597)
	);

	bfr new_net_5599_bfr_before (
		.din(new_net_5599),
		.dout(new_net_5598)
	);

	bfr new_net_5600_bfr_before (
		.din(new_net_5600),
		.dout(new_net_5599)
	);

	bfr new_net_5601_bfr_before (
		.din(new_net_5601),
		.dout(new_net_5600)
	);

	bfr new_net_5602_bfr_before (
		.din(new_net_5602),
		.dout(new_net_5601)
	);

	bfr new_net_5603_bfr_before (
		.din(new_net_5603),
		.dout(new_net_5602)
	);

	bfr new_net_5604_bfr_before (
		.din(new_net_5604),
		.dout(new_net_5603)
	);

	bfr new_net_5605_bfr_before (
		.din(new_net_5605),
		.dout(new_net_5604)
	);

	bfr new_net_5606_bfr_before (
		.din(new_net_5606),
		.dout(new_net_5605)
	);

	bfr new_net_5607_bfr_before (
		.din(new_net_5607),
		.dout(new_net_5606)
	);

	bfr new_net_5608_bfr_before (
		.din(new_net_5608),
		.dout(new_net_5607)
	);

	bfr new_net_5609_bfr_before (
		.din(new_net_5609),
		.dout(new_net_5608)
	);

	bfr new_net_5610_bfr_before (
		.din(new_net_5610),
		.dout(new_net_5609)
	);

	bfr new_net_5611_bfr_before (
		.din(new_net_5611),
		.dout(new_net_5610)
	);

	bfr new_net_5612_bfr_before (
		.din(new_net_5612),
		.dout(new_net_5611)
	);

	bfr new_net_5613_bfr_before (
		.din(new_net_5613),
		.dout(new_net_5612)
	);

	bfr new_net_5614_bfr_before (
		.din(new_net_5614),
		.dout(new_net_5613)
	);

	bfr new_net_5615_bfr_before (
		.din(new_net_5615),
		.dout(new_net_5614)
	);

	bfr new_net_5616_bfr_before (
		.din(new_net_5616),
		.dout(new_net_5615)
	);

	bfr new_net_5617_bfr_before (
		.din(new_net_5617),
		.dout(new_net_5616)
	);

	bfr new_net_5618_bfr_before (
		.din(new_net_5618),
		.dout(new_net_5617)
	);

	bfr new_net_5619_bfr_before (
		.din(new_net_5619),
		.dout(new_net_5618)
	);

	spl3L new_net_2027_v_fanout (
		.a(new_net_2027),
		.b(new_net_5619),
		.c(new_net_1124),
		.d(new_net_1125)
	);

	spl3L n_0782__v_fanout (
		.a(n_0782_),
		.b(new_net_1426),
		.c(new_net_1425),
		.d(new_net_1427)
	);

	spl3L n_1209__v_fanout (
		.a(n_1209_),
		.b(new_net_618),
		.c(new_net_617),
		.d(new_net_619)
	);

	spl2 new_net_2088_v_fanout (
		.a(new_net_2088),
		.b(new_net_1092),
		.c(new_net_1090)
	);

	spl2 new_net_2091_v_fanout (
		.a(new_net_2091),
		.b(new_net_1489),
		.c(new_net_1490)
	);

	spl2 new_net_2100_v_fanout (
		.a(new_net_2100),
		.b(new_net_1014),
		.c(new_net_1013)
	);

	spl2 new_net_2072_v_fanout (
		.a(new_net_2072),
		.b(new_net_1800),
		.c(new_net_1798)
	);

	spl4L n_0812__v_fanout (
		.a(n_0812_),
		.b(new_net_1021),
		.c(new_net_1022),
		.d(new_net_1023),
		.e(new_net_1020)
	);

	spl4L n_1187__v_fanout (
		.a(n_1187_),
		.b(new_net_1848),
		.c(new_net_1846),
		.d(new_net_1847),
		.e(new_net_1845)
	);

	bfr new_net_5620_bfr_after (
		.din(n_0770_),
		.dout(new_net_5620)
	);

	bfr new_net_5621_bfr_after (
		.din(new_net_5620),
		.dout(new_net_5621)
	);

	bfr new_net_5622_bfr_after (
		.din(new_net_5621),
		.dout(new_net_5622)
	);

	spl2 n_0770__v_fanout (
		.a(new_net_5622),
		.b(new_net_902),
		.c(new_net_901)
	);

	spl3L n_0727__v_fanout (
		.a(n_0727_),
		.b(new_net_58),
		.c(new_net_56),
		.d(new_net_57)
	);

	spl4L n_1167__v_fanout (
		.a(n_1167_),
		.b(new_net_500),
		.c(new_net_498),
		.d(new_net_499),
		.e(new_net_497)
	);

	bfr new_net_5623_bfr_before (
		.din(new_net_5623),
		.dout(N549)
	);

	bfr new_net_5624_bfr_before (
		.din(new_net_5624),
		.dout(new_net_5623)
	);

	bfr new_net_5625_bfr_before (
		.din(new_net_5625),
		.dout(new_net_5624)
	);

	bfr new_net_5626_bfr_before (
		.din(new_net_5626),
		.dout(new_net_5625)
	);

	bfr new_net_5627_bfr_before (
		.din(new_net_5627),
		.dout(new_net_5626)
	);

	bfr new_net_5628_bfr_before (
		.din(new_net_5628),
		.dout(new_net_5627)
	);

	bfr new_net_5629_bfr_before (
		.din(new_net_5629),
		.dout(new_net_5628)
	);

	bfr new_net_5630_bfr_before (
		.din(new_net_5630),
		.dout(new_net_5629)
	);

	bfr new_net_5631_bfr_before (
		.din(new_net_5631),
		.dout(new_net_5630)
	);

	bfr new_net_5632_bfr_before (
		.din(new_net_5632),
		.dout(new_net_5631)
	);

	bfr new_net_5633_bfr_before (
		.din(new_net_5633),
		.dout(new_net_5632)
	);

	bfr new_net_5634_bfr_before (
		.din(new_net_5634),
		.dout(new_net_5633)
	);

	bfr new_net_5635_bfr_before (
		.din(new_net_5635),
		.dout(new_net_5634)
	);

	bfr new_net_5636_bfr_before (
		.din(new_net_5636),
		.dout(new_net_5635)
	);

	bfr new_net_5637_bfr_before (
		.din(new_net_5637),
		.dout(new_net_5636)
	);

	bfr new_net_5638_bfr_before (
		.din(new_net_5638),
		.dout(new_net_5637)
	);

	bfr new_net_5639_bfr_before (
		.din(new_net_5639),
		.dout(new_net_5638)
	);

	bfr new_net_5640_bfr_before (
		.din(new_net_5640),
		.dout(new_net_5639)
	);

	bfr new_net_5641_bfr_before (
		.din(new_net_5641),
		.dout(new_net_5640)
	);

	bfr new_net_5642_bfr_before (
		.din(new_net_5642),
		.dout(new_net_5641)
	);

	bfr new_net_5643_bfr_before (
		.din(new_net_5643),
		.dout(new_net_5642)
	);

	bfr new_net_5644_bfr_before (
		.din(new_net_5644),
		.dout(new_net_5643)
	);

	bfr new_net_5645_bfr_before (
		.din(new_net_5645),
		.dout(new_net_5644)
	);

	bfr new_net_5646_bfr_before (
		.din(new_net_5646),
		.dout(new_net_5645)
	);

	bfr new_net_5647_bfr_before (
		.din(new_net_5647),
		.dout(new_net_5646)
	);

	bfr new_net_5648_bfr_before (
		.din(new_net_5648),
		.dout(new_net_5647)
	);

	bfr new_net_5649_bfr_before (
		.din(new_net_5649),
		.dout(new_net_5648)
	);

	bfr new_net_5650_bfr_before (
		.din(new_net_5650),
		.dout(new_net_5649)
	);

	bfr new_net_5651_bfr_before (
		.din(new_net_5651),
		.dout(new_net_5650)
	);

	bfr new_net_5652_bfr_before (
		.din(new_net_5652),
		.dout(new_net_5651)
	);

	bfr new_net_5653_bfr_before (
		.din(new_net_5653),
		.dout(new_net_5652)
	);

	bfr new_net_5654_bfr_before (
		.din(new_net_5654),
		.dout(new_net_5653)
	);

	bfr new_net_5655_bfr_before (
		.din(new_net_5655),
		.dout(new_net_5654)
	);

	bfr new_net_5656_bfr_before (
		.din(new_net_5656),
		.dout(new_net_5655)
	);

	bfr new_net_5657_bfr_before (
		.din(new_net_5657),
		.dout(new_net_5656)
	);

	bfr new_net_5658_bfr_before (
		.din(new_net_5658),
		.dout(new_net_5657)
	);

	bfr new_net_5659_bfr_before (
		.din(new_net_5659),
		.dout(new_net_5658)
	);

	bfr new_net_5660_bfr_before (
		.din(new_net_5660),
		.dout(new_net_5659)
	);

	bfr new_net_5661_bfr_before (
		.din(new_net_5661),
		.dout(new_net_5660)
	);

	bfr new_net_5662_bfr_before (
		.din(new_net_5662),
		.dout(new_net_5661)
	);

	bfr new_net_5663_bfr_before (
		.din(new_net_5663),
		.dout(new_net_5662)
	);

	bfr new_net_5664_bfr_before (
		.din(new_net_5664),
		.dout(new_net_5663)
	);

	bfr new_net_5665_bfr_before (
		.din(new_net_5665),
		.dout(new_net_5664)
	);

	bfr new_net_5666_bfr_before (
		.din(new_net_5666),
		.dout(new_net_5665)
	);

	bfr new_net_5667_bfr_before (
		.din(new_net_5667),
		.dout(new_net_5666)
	);

	bfr new_net_5668_bfr_before (
		.din(new_net_5668),
		.dout(new_net_5667)
	);

	bfr new_net_5669_bfr_before (
		.din(new_net_5669),
		.dout(new_net_5668)
	);

	bfr new_net_5670_bfr_before (
		.din(new_net_5670),
		.dout(new_net_5669)
	);

	bfr new_net_5671_bfr_before (
		.din(new_net_5671),
		.dout(new_net_5670)
	);

	bfr new_net_5672_bfr_before (
		.din(new_net_5672),
		.dout(new_net_5671)
	);

	bfr new_net_5673_bfr_before (
		.din(new_net_5673),
		.dout(new_net_5672)
	);

	bfr new_net_5674_bfr_before (
		.din(new_net_5674),
		.dout(new_net_5673)
	);

	bfr new_net_5675_bfr_before (
		.din(new_net_5675),
		.dout(new_net_5674)
	);

	bfr new_net_5676_bfr_before (
		.din(new_net_5676),
		.dout(new_net_5675)
	);

	bfr new_net_5677_bfr_before (
		.din(new_net_5677),
		.dout(new_net_5676)
	);

	bfr new_net_5678_bfr_before (
		.din(new_net_5678),
		.dout(new_net_5677)
	);

	bfr new_net_5679_bfr_before (
		.din(new_net_5679),
		.dout(new_net_5678)
	);

	bfr new_net_5680_bfr_before (
		.din(new_net_5680),
		.dout(new_net_5679)
	);

	spl3L new_net_2042_v_fanout (
		.a(new_net_2042),
		.b(new_net_1227),
		.c(new_net_1228),
		.d(new_net_5680)
	);

	spl4L n_0848__v_fanout (
		.a(n_0848_),
		.b(new_net_1943),
		.c(new_net_1944),
		.d(new_net_1942),
		.e(new_net_1941)
	);

	spl4L n_1273__v_fanout (
		.a(n_1273_),
		.b(new_net_558),
		.c(new_net_559),
		.d(new_net_560),
		.e(new_net_557)
	);

	spl2 n_1199__v_fanout (
		.a(n_1199_),
		.b(new_net_1365),
		.c(new_net_1364)
	);

	spl4L n_0804__v_fanout (
		.a(n_0804_),
		.b(new_net_915),
		.c(new_net_913),
		.d(new_net_914),
		.e(new_net_912)
	);

	spl2 new_net_2089_v_fanout (
		.a(new_net_2089),
		.b(new_net_1603),
		.c(new_net_1604)
	);

	spl4L n_1235__v_fanout (
		.a(n_1235_),
		.b(new_net_1744),
		.c(new_net_1742),
		.d(new_net_1743),
		.e(new_net_1741)
	);

	spl4L n_1260__v_fanout (
		.a(n_1260_),
		.b(new_net_819),
		.c(new_net_820),
		.d(new_net_821),
		.e(new_net_818)
	);

	spl4L n_0750__v_fanout (
		.a(n_0750_),
		.b(new_net_761),
		.c(new_net_762),
		.d(new_net_763),
		.e(new_net_760)
	);

	spl2 new_net_2073_v_fanout (
		.a(new_net_2073),
		.b(new_net_999),
		.c(new_net_997)
	);

	spl4L n_0890__v_fanout (
		.a(n_0890_),
		.b(new_net_1055),
		.c(new_net_1056),
		.d(new_net_1054),
		.e(new_net_1053)
	);

	spl2 new_net_2078_v_fanout (
		.a(new_net_2078),
		.b(new_net_1927),
		.c(new_net_1926)
	);

	spl2 new_net_2098_v_fanout (
		.a(new_net_2098),
		.b(new_net_64),
		.c(new_net_66)
	);

	spl3L n_0785__v_fanout (
		.a(n_0785_),
		.b(new_net_1502),
		.c(new_net_1500),
		.d(new_net_1501)
	);

	spl2 new_net_2087_v_fanout (
		.a(new_net_2087),
		.b(new_net_751),
		.c(new_net_750)
	);

	spl2 n_1248__v_fanout (
		.a(n_1248_),
		.b(new_net_1313),
		.c(new_net_1312)
	);

	spl3L n_1206__v_fanout (
		.a(n_1206_),
		.b(new_net_1517),
		.c(new_net_1515),
		.d(new_net_1516)
	);

	spl4L n_1255__v_fanout (
		.a(n_1255_),
		.b(new_net_772),
		.c(new_net_773),
		.d(new_net_771),
		.e(new_net_770)
	);

	spl4L n_1151__v_fanout (
		.a(n_1151_),
		.b(new_net_612),
		.c(new_net_613),
		.d(new_net_614),
		.e(new_net_611)
	);

	spl4L n_0887__v_fanout (
		.a(n_0887_),
		.b(new_net_1958),
		.c(new_net_1959),
		.d(new_net_1960),
		.e(new_net_1957)
	);

	spl4L n_0761__v_fanout (
		.a(n_0761_),
		.b(new_net_990),
		.c(new_net_991),
		.d(new_net_989),
		.e(new_net_988)
	);

	spl4L n_0679__v_fanout (
		.a(n_0679_),
		.b(new_net_1913),
		.c(new_net_1914),
		.d(new_net_1912),
		.e(new_net_1911)
	);

	spl3L n_1216__v_fanout (
		.a(n_1216_),
		.b(new_net_1335),
		.c(new_net_1333),
		.d(new_net_1334)
	);

	spl4L n_0673__v_fanout (
		.a(n_0673_),
		.b(new_net_1774),
		.c(new_net_1773),
		.d(new_net_1772),
		.e(new_net_1771)
	);

	bfr new_net_5681_bfr_before (
		.din(new_net_5681),
		.dout(N486)
	);

	bfr new_net_5682_bfr_before (
		.din(new_net_5682),
		.dout(new_net_5681)
	);

	bfr new_net_5683_bfr_before (
		.din(new_net_5683),
		.dout(new_net_5682)
	);

	bfr new_net_5684_bfr_before (
		.din(new_net_5684),
		.dout(new_net_5683)
	);

	bfr new_net_5685_bfr_before (
		.din(new_net_5685),
		.dout(new_net_5684)
	);

	bfr new_net_5686_bfr_before (
		.din(new_net_5686),
		.dout(new_net_5685)
	);

	bfr new_net_5687_bfr_before (
		.din(new_net_5687),
		.dout(new_net_5686)
	);

	bfr new_net_5688_bfr_before (
		.din(new_net_5688),
		.dout(new_net_5687)
	);

	bfr new_net_5689_bfr_before (
		.din(new_net_5689),
		.dout(new_net_5688)
	);

	bfr new_net_5690_bfr_before (
		.din(new_net_5690),
		.dout(new_net_5689)
	);

	bfr new_net_5691_bfr_before (
		.din(new_net_5691),
		.dout(new_net_5690)
	);

	bfr new_net_5692_bfr_before (
		.din(new_net_5692),
		.dout(new_net_5691)
	);

	bfr new_net_5693_bfr_before (
		.din(new_net_5693),
		.dout(new_net_5692)
	);

	bfr new_net_5694_bfr_before (
		.din(new_net_5694),
		.dout(new_net_5693)
	);

	bfr new_net_5695_bfr_before (
		.din(new_net_5695),
		.dout(new_net_5694)
	);

	bfr new_net_5696_bfr_before (
		.din(new_net_5696),
		.dout(new_net_5695)
	);

	bfr new_net_5697_bfr_before (
		.din(new_net_5697),
		.dout(new_net_5696)
	);

	bfr new_net_5698_bfr_before (
		.din(new_net_5698),
		.dout(new_net_5697)
	);

	bfr new_net_5699_bfr_before (
		.din(new_net_5699),
		.dout(new_net_5698)
	);

	bfr new_net_5700_bfr_before (
		.din(new_net_5700),
		.dout(new_net_5699)
	);

	bfr new_net_5701_bfr_before (
		.din(new_net_5701),
		.dout(new_net_5700)
	);

	bfr new_net_5702_bfr_before (
		.din(new_net_5702),
		.dout(new_net_5701)
	);

	bfr new_net_5703_bfr_before (
		.din(new_net_5703),
		.dout(new_net_5702)
	);

	bfr new_net_5704_bfr_before (
		.din(new_net_5704),
		.dout(new_net_5703)
	);

	bfr new_net_5705_bfr_before (
		.din(new_net_5705),
		.dout(new_net_5704)
	);

	bfr new_net_5706_bfr_before (
		.din(new_net_5706),
		.dout(new_net_5705)
	);

	bfr new_net_5707_bfr_before (
		.din(new_net_5707),
		.dout(new_net_5706)
	);

	bfr new_net_5708_bfr_before (
		.din(new_net_5708),
		.dout(new_net_5707)
	);

	bfr new_net_5709_bfr_before (
		.din(new_net_5709),
		.dout(new_net_5708)
	);

	bfr new_net_5710_bfr_before (
		.din(new_net_5710),
		.dout(new_net_5709)
	);

	bfr new_net_5711_bfr_before (
		.din(new_net_5711),
		.dout(new_net_5710)
	);

	bfr new_net_5712_bfr_before (
		.din(new_net_5712),
		.dout(new_net_5711)
	);

	bfr new_net_5713_bfr_before (
		.din(new_net_5713),
		.dout(new_net_5712)
	);

	bfr new_net_5714_bfr_before (
		.din(new_net_5714),
		.dout(new_net_5713)
	);

	bfr new_net_5715_bfr_before (
		.din(new_net_5715),
		.dout(new_net_5714)
	);

	bfr new_net_5716_bfr_before (
		.din(new_net_5716),
		.dout(new_net_5715)
	);

	bfr new_net_5717_bfr_before (
		.din(new_net_5717),
		.dout(new_net_5716)
	);

	bfr new_net_5718_bfr_before (
		.din(new_net_5718),
		.dout(new_net_5717)
	);

	bfr new_net_5719_bfr_before (
		.din(new_net_5719),
		.dout(new_net_5718)
	);

	bfr new_net_5720_bfr_before (
		.din(new_net_5720),
		.dout(new_net_5719)
	);

	bfr new_net_5721_bfr_before (
		.din(new_net_5721),
		.dout(new_net_5720)
	);

	bfr new_net_5722_bfr_before (
		.din(new_net_5722),
		.dout(new_net_5721)
	);

	bfr new_net_5723_bfr_before (
		.din(new_net_5723),
		.dout(new_net_5722)
	);

	bfr new_net_5724_bfr_before (
		.din(new_net_5724),
		.dout(new_net_5723)
	);

	bfr new_net_5725_bfr_before (
		.din(new_net_5725),
		.dout(new_net_5724)
	);

	bfr new_net_5726_bfr_before (
		.din(new_net_5726),
		.dout(new_net_5725)
	);

	bfr new_net_5727_bfr_before (
		.din(new_net_5727),
		.dout(new_net_5726)
	);

	bfr new_net_5728_bfr_before (
		.din(new_net_5728),
		.dout(new_net_5727)
	);

	bfr new_net_5729_bfr_before (
		.din(new_net_5729),
		.dout(new_net_5728)
	);

	bfr new_net_5730_bfr_before (
		.din(new_net_5730),
		.dout(new_net_5729)
	);

	bfr new_net_5731_bfr_before (
		.din(new_net_5731),
		.dout(new_net_5730)
	);

	bfr new_net_5732_bfr_before (
		.din(new_net_5732),
		.dout(new_net_5731)
	);

	bfr new_net_5733_bfr_before (
		.din(new_net_5733),
		.dout(new_net_5732)
	);

	bfr new_net_5734_bfr_before (
		.din(new_net_5734),
		.dout(new_net_5733)
	);

	bfr new_net_5735_bfr_before (
		.din(new_net_5735),
		.dout(new_net_5734)
	);

	bfr new_net_5736_bfr_before (
		.din(new_net_5736),
		.dout(new_net_5735)
	);

	bfr new_net_5737_bfr_before (
		.din(new_net_5737),
		.dout(new_net_5736)
	);

	bfr new_net_5738_bfr_before (
		.din(new_net_5738),
		.dout(new_net_5737)
	);

	spl3L new_net_2024_v_fanout (
		.a(new_net_2024),
		.b(new_net_5738),
		.c(new_net_1345),
		.d(new_net_1344)
	);

	spl2 new_net_2081_v_fanout (
		.a(new_net_2081),
		.b(new_net_489),
		.c(new_net_490)
	);

	bfr new_net_5739_bfr_before (
		.din(new_net_5739),
		.dout(new_net_2101)
	);

	spl2 n_0663__v_fanout (
		.a(n_0663_),
		.b(new_net_5739),
		.c(new_net_733)
	);

	spl3L n_0723__v_fanout (
		.a(n_0723_),
		.b(new_net_18),
		.c(new_net_17),
		.d(new_net_19)
	);

	spl4L n_0824__v_fanout (
		.a(n_0824_),
		.b(new_net_465),
		.c(new_net_466),
		.d(new_net_467),
		.e(new_net_464)
	);

	spl3L n_1134__v_fanout (
		.a(n_1134_),
		.b(new_net_366),
		.c(new_net_365),
		.d(new_net_367)
	);

	spl4L n_1282__v_fanout (
		.a(n_1282_),
		.b(new_net_1527),
		.c(new_net_1528),
		.d(new_net_1529),
		.e(new_net_1526)
	);

	spl4L n_1262__v_fanout (
		.a(n_1262_),
		.b(new_net_928),
		.c(new_net_929),
		.d(new_net_927),
		.e(new_net_926)
	);

	spl3L n_0775__v_fanout (
		.a(n_0775_),
		.b(new_net_1265),
		.c(new_net_1263),
		.d(new_net_1264)
	);

	spl4L n_0758__v_fanout (
		.a(n_0758_),
		.b(new_net_921),
		.c(new_net_919),
		.d(new_net_920),
		.e(new_net_918)
	);

	spl2 new_net_2090_v_fanout (
		.a(new_net_2090),
		.b(new_net_525),
		.c(new_net_526)
	);

	spl4L n_1201__v_fanout (
		.a(n_1201_),
		.b(new_net_1403),
		.c(new_net_1404),
		.d(new_net_1402),
		.e(new_net_1401)
	);

	bfr new_net_5740_bfr_before (
		.din(new_net_5740),
		.dout(N513)
	);

	bfr new_net_5741_bfr_before (
		.din(new_net_5741),
		.dout(new_net_5740)
	);

	bfr new_net_5742_bfr_before (
		.din(new_net_5742),
		.dout(new_net_5741)
	);

	bfr new_net_5743_bfr_before (
		.din(new_net_5743),
		.dout(new_net_5742)
	);

	bfr new_net_5744_bfr_before (
		.din(new_net_5744),
		.dout(new_net_5743)
	);

	bfr new_net_5745_bfr_before (
		.din(new_net_5745),
		.dout(new_net_5744)
	);

	bfr new_net_5746_bfr_before (
		.din(new_net_5746),
		.dout(new_net_5745)
	);

	bfr new_net_5747_bfr_before (
		.din(new_net_5747),
		.dout(new_net_5746)
	);

	bfr new_net_5748_bfr_before (
		.din(new_net_5748),
		.dout(new_net_5747)
	);

	bfr new_net_5749_bfr_before (
		.din(new_net_5749),
		.dout(new_net_5748)
	);

	bfr new_net_5750_bfr_before (
		.din(new_net_5750),
		.dout(new_net_5749)
	);

	bfr new_net_5751_bfr_before (
		.din(new_net_5751),
		.dout(new_net_5750)
	);

	bfr new_net_5752_bfr_before (
		.din(new_net_5752),
		.dout(new_net_5751)
	);

	bfr new_net_5753_bfr_before (
		.din(new_net_5753),
		.dout(new_net_5752)
	);

	bfr new_net_5754_bfr_before (
		.din(new_net_5754),
		.dout(new_net_5753)
	);

	bfr new_net_5755_bfr_before (
		.din(new_net_5755),
		.dout(new_net_5754)
	);

	bfr new_net_5756_bfr_before (
		.din(new_net_5756),
		.dout(new_net_5755)
	);

	bfr new_net_5757_bfr_before (
		.din(new_net_5757),
		.dout(new_net_5756)
	);

	bfr new_net_5758_bfr_before (
		.din(new_net_5758),
		.dout(new_net_5757)
	);

	bfr new_net_5759_bfr_before (
		.din(new_net_5759),
		.dout(new_net_5758)
	);

	bfr new_net_5760_bfr_before (
		.din(new_net_5760),
		.dout(new_net_5759)
	);

	bfr new_net_5761_bfr_before (
		.din(new_net_5761),
		.dout(new_net_5760)
	);

	bfr new_net_5762_bfr_before (
		.din(new_net_5762),
		.dout(new_net_5761)
	);

	bfr new_net_5763_bfr_before (
		.din(new_net_5763),
		.dout(new_net_5762)
	);

	bfr new_net_5764_bfr_before (
		.din(new_net_5764),
		.dout(new_net_5763)
	);

	bfr new_net_5765_bfr_before (
		.din(new_net_5765),
		.dout(new_net_5764)
	);

	bfr new_net_5766_bfr_before (
		.din(new_net_5766),
		.dout(new_net_5765)
	);

	bfr new_net_5767_bfr_before (
		.din(new_net_5767),
		.dout(new_net_5766)
	);

	bfr new_net_5768_bfr_before (
		.din(new_net_5768),
		.dout(new_net_5767)
	);

	bfr new_net_5769_bfr_before (
		.din(new_net_5769),
		.dout(new_net_5768)
	);

	bfr new_net_5770_bfr_before (
		.din(new_net_5770),
		.dout(new_net_5769)
	);

	bfr new_net_5771_bfr_before (
		.din(new_net_5771),
		.dout(new_net_5770)
	);

	bfr new_net_5772_bfr_before (
		.din(new_net_5772),
		.dout(new_net_5771)
	);

	bfr new_net_5773_bfr_before (
		.din(new_net_5773),
		.dout(new_net_5772)
	);

	bfr new_net_5774_bfr_before (
		.din(new_net_5774),
		.dout(new_net_5773)
	);

	bfr new_net_5775_bfr_before (
		.din(new_net_5775),
		.dout(new_net_5774)
	);

	bfr new_net_5776_bfr_before (
		.din(new_net_5776),
		.dout(new_net_5775)
	);

	bfr new_net_5777_bfr_before (
		.din(new_net_5777),
		.dout(new_net_5776)
	);

	bfr new_net_5778_bfr_before (
		.din(new_net_5778),
		.dout(new_net_5777)
	);

	bfr new_net_5779_bfr_before (
		.din(new_net_5779),
		.dout(new_net_5778)
	);

	bfr new_net_5780_bfr_before (
		.din(new_net_5780),
		.dout(new_net_5779)
	);

	bfr new_net_5781_bfr_before (
		.din(new_net_5781),
		.dout(new_net_5780)
	);

	bfr new_net_5782_bfr_before (
		.din(new_net_5782),
		.dout(new_net_5781)
	);

	bfr new_net_5783_bfr_before (
		.din(new_net_5783),
		.dout(new_net_5782)
	);

	bfr new_net_5784_bfr_before (
		.din(new_net_5784),
		.dout(new_net_5783)
	);

	bfr new_net_5785_bfr_before (
		.din(new_net_5785),
		.dout(new_net_5784)
	);

	bfr new_net_5786_bfr_before (
		.din(new_net_5786),
		.dout(new_net_5785)
	);

	bfr new_net_5787_bfr_before (
		.din(new_net_5787),
		.dout(new_net_5786)
	);

	bfr new_net_5788_bfr_before (
		.din(new_net_5788),
		.dout(new_net_5787)
	);

	bfr new_net_5789_bfr_before (
		.din(new_net_5789),
		.dout(new_net_5788)
	);

	bfr new_net_5790_bfr_before (
		.din(new_net_5790),
		.dout(new_net_5789)
	);

	bfr new_net_5791_bfr_before (
		.din(new_net_5791),
		.dout(new_net_5790)
	);

	bfr new_net_5792_bfr_before (
		.din(new_net_5792),
		.dout(new_net_5791)
	);

	bfr new_net_5793_bfr_before (
		.din(new_net_5793),
		.dout(new_net_5792)
	);

	bfr new_net_5794_bfr_before (
		.din(new_net_5794),
		.dout(new_net_5793)
	);

	bfr new_net_5795_bfr_before (
		.din(new_net_5795),
		.dout(new_net_5794)
	);

	bfr new_net_5796_bfr_before (
		.din(new_net_5796),
		.dout(new_net_5795)
	);

	bfr new_net_5797_bfr_before (
		.din(new_net_5797),
		.dout(new_net_5796)
	);

	spl3L new_net_2031_v_fanout (
		.a(new_net_2031),
		.b(new_net_5797),
		.c(new_net_1768),
		.d(new_net_1767)
	);

	spl4L n_0872__v_fanout (
		.a(n_0872_),
		.b(new_net_309),
		.c(new_net_310),
		.d(new_net_308),
		.e(new_net_307)
	);

	spl2 n_0833__v_fanout (
		.a(n_0833_),
		.b(new_net_1615),
		.c(new_net_1614)
	);

	spl3L n_1127__v_fanout (
		.a(n_1127_),
		.b(new_net_1462),
		.c(new_net_1461),
		.d(new_net_1463)
	);

	spl2 new_net_2085_v_fanout (
		.a(new_net_2085),
		.b(new_net_1246),
		.c(new_net_1247)
	);

	spl4L n_0881__v_fanout (
		.a(n_0881_),
		.b(new_net_1301),
		.c(new_net_1300),
		.d(new_net_1299),
		.e(new_net_1298)
	);

	spl2 new_net_2093_v_fanout (
		.a(new_net_2093),
		.b(new_net_1412),
		.c(new_net_1411)
	);

	bfr new_net_5798_bfr_before (
		.din(new_net_5798),
		.dout(N813)
	);

	bfr new_net_5799_bfr_before (
		.din(new_net_5799),
		.dout(new_net_5798)
	);

	bfr new_net_5800_bfr_before (
		.din(new_net_5800),
		.dout(new_net_5799)
	);

	bfr new_net_5801_bfr_before (
		.din(new_net_5801),
		.dout(new_net_5800)
	);

	bfr new_net_5802_bfr_before (
		.din(new_net_5802),
		.dout(new_net_5801)
	);

	bfr new_net_5803_bfr_before (
		.din(new_net_5803),
		.dout(new_net_5802)
	);

	bfr new_net_5804_bfr_before (
		.din(new_net_5804),
		.dout(new_net_5803)
	);

	bfr new_net_5805_bfr_before (
		.din(new_net_5805),
		.dout(new_net_5804)
	);

	bfr new_net_5806_bfr_before (
		.din(new_net_5806),
		.dout(new_net_5805)
	);

	bfr new_net_5807_bfr_before (
		.din(new_net_5807),
		.dout(new_net_5806)
	);

	bfr new_net_5808_bfr_before (
		.din(new_net_5808),
		.dout(new_net_5807)
	);

	bfr new_net_5809_bfr_before (
		.din(new_net_5809),
		.dout(new_net_5808)
	);

	bfr new_net_5810_bfr_before (
		.din(new_net_5810),
		.dout(new_net_5809)
	);

	bfr new_net_5811_bfr_before (
		.din(new_net_5811),
		.dout(new_net_5810)
	);

	bfr new_net_5812_bfr_before (
		.din(new_net_5812),
		.dout(new_net_5811)
	);

	bfr new_net_5813_bfr_before (
		.din(new_net_5813),
		.dout(new_net_5812)
	);

	bfr new_net_5814_bfr_before (
		.din(new_net_5814),
		.dout(new_net_5813)
	);

	bfr new_net_5815_bfr_before (
		.din(new_net_5815),
		.dout(new_net_5814)
	);

	bfr new_net_5816_bfr_before (
		.din(new_net_5816),
		.dout(new_net_5815)
	);

	bfr new_net_5817_bfr_before (
		.din(new_net_5817),
		.dout(new_net_5816)
	);

	bfr new_net_5818_bfr_before (
		.din(new_net_5818),
		.dout(new_net_5817)
	);

	bfr new_net_5819_bfr_before (
		.din(new_net_5819),
		.dout(new_net_5818)
	);

	bfr new_net_5820_bfr_before (
		.din(new_net_5820),
		.dout(new_net_5819)
	);

	bfr new_net_5821_bfr_before (
		.din(new_net_5821),
		.dout(new_net_5820)
	);

	bfr new_net_5822_bfr_before (
		.din(new_net_5822),
		.dout(new_net_5821)
	);

	bfr new_net_5823_bfr_before (
		.din(new_net_5823),
		.dout(new_net_5822)
	);

	bfr new_net_5824_bfr_before (
		.din(new_net_5824),
		.dout(new_net_5823)
	);

	bfr new_net_5825_bfr_before (
		.din(new_net_5825),
		.dout(new_net_5824)
	);

	bfr new_net_5826_bfr_before (
		.din(new_net_5826),
		.dout(new_net_5825)
	);

	bfr new_net_5827_bfr_before (
		.din(new_net_5827),
		.dout(new_net_5826)
	);

	bfr new_net_5828_bfr_before (
		.din(new_net_5828),
		.dout(new_net_5827)
	);

	bfr new_net_5829_bfr_before (
		.din(new_net_5829),
		.dout(new_net_5828)
	);

	bfr new_net_5830_bfr_before (
		.din(new_net_5830),
		.dout(new_net_5829)
	);

	bfr new_net_5831_bfr_before (
		.din(new_net_5831),
		.dout(new_net_5830)
	);

	bfr new_net_5832_bfr_before (
		.din(new_net_5832),
		.dout(new_net_5831)
	);

	bfr new_net_5833_bfr_before (
		.din(new_net_5833),
		.dout(new_net_5832)
	);

	bfr new_net_5834_bfr_before (
		.din(new_net_5834),
		.dout(new_net_5833)
	);

	bfr new_net_5835_bfr_before (
		.din(new_net_5835),
		.dout(new_net_5834)
	);

	bfr new_net_5836_bfr_before (
		.din(new_net_5836),
		.dout(new_net_5835)
	);

	bfr new_net_5837_bfr_before (
		.din(new_net_5837),
		.dout(new_net_5836)
	);

	bfr new_net_5838_bfr_before (
		.din(new_net_5838),
		.dout(new_net_5837)
	);

	bfr new_net_5839_bfr_before (
		.din(new_net_5839),
		.dout(new_net_5838)
	);

	bfr new_net_5840_bfr_before (
		.din(new_net_5840),
		.dout(new_net_5839)
	);

	bfr new_net_5841_bfr_before (
		.din(new_net_5841),
		.dout(new_net_5840)
	);

	bfr new_net_5842_bfr_before (
		.din(new_net_5842),
		.dout(new_net_5841)
	);

	bfr new_net_5843_bfr_before (
		.din(new_net_5843),
		.dout(new_net_5842)
	);

	bfr new_net_5844_bfr_before (
		.din(new_net_5844),
		.dout(new_net_5843)
	);

	bfr new_net_5845_bfr_before (
		.din(new_net_5845),
		.dout(new_net_5844)
	);

	bfr new_net_5846_bfr_before (
		.din(new_net_5846),
		.dout(new_net_5845)
	);

	bfr new_net_5847_bfr_before (
		.din(new_net_5847),
		.dout(new_net_5846)
	);

	bfr new_net_5848_bfr_before (
		.din(new_net_5848),
		.dout(new_net_5847)
	);

	bfr new_net_5849_bfr_before (
		.din(new_net_5849),
		.dout(new_net_5848)
	);

	bfr new_net_5850_bfr_before (
		.din(new_net_5850),
		.dout(new_net_5849)
	);

	bfr new_net_5851_bfr_before (
		.din(new_net_5851),
		.dout(new_net_5850)
	);

	bfr new_net_5852_bfr_before (
		.din(new_net_5852),
		.dout(new_net_5851)
	);

	bfr new_net_5853_bfr_before (
		.din(new_net_5853),
		.dout(new_net_5852)
	);

	bfr new_net_5854_bfr_before (
		.din(new_net_5854),
		.dout(new_net_5853)
	);

	bfr new_net_5855_bfr_before (
		.din(new_net_5855),
		.dout(new_net_5854)
	);

	spl3L new_net_2045_v_fanout (
		.a(new_net_2045),
		.b(new_net_1561),
		.c(new_net_1562),
		.d(new_net_5855)
	);

	bfr new_net_5856_bfr_before (
		.din(new_net_5856),
		.dout(N543)
	);

	bfr new_net_5857_bfr_before (
		.din(new_net_5857),
		.dout(new_net_5856)
	);

	bfr new_net_5858_bfr_before (
		.din(new_net_5858),
		.dout(new_net_5857)
	);

	bfr new_net_5859_bfr_before (
		.din(new_net_5859),
		.dout(new_net_5858)
	);

	bfr new_net_5860_bfr_before (
		.din(new_net_5860),
		.dout(new_net_5859)
	);

	bfr new_net_5861_bfr_before (
		.din(new_net_5861),
		.dout(new_net_5860)
	);

	bfr new_net_5862_bfr_before (
		.din(new_net_5862),
		.dout(new_net_5861)
	);

	bfr new_net_5863_bfr_before (
		.din(new_net_5863),
		.dout(new_net_5862)
	);

	bfr new_net_5864_bfr_before (
		.din(new_net_5864),
		.dout(new_net_5863)
	);

	bfr new_net_5865_bfr_before (
		.din(new_net_5865),
		.dout(new_net_5864)
	);

	bfr new_net_5866_bfr_before (
		.din(new_net_5866),
		.dout(new_net_5865)
	);

	bfr new_net_5867_bfr_before (
		.din(new_net_5867),
		.dout(new_net_5866)
	);

	bfr new_net_5868_bfr_before (
		.din(new_net_5868),
		.dout(new_net_5867)
	);

	bfr new_net_5869_bfr_before (
		.din(new_net_5869),
		.dout(new_net_5868)
	);

	bfr new_net_5870_bfr_before (
		.din(new_net_5870),
		.dout(new_net_5869)
	);

	bfr new_net_5871_bfr_before (
		.din(new_net_5871),
		.dout(new_net_5870)
	);

	bfr new_net_5872_bfr_before (
		.din(new_net_5872),
		.dout(new_net_5871)
	);

	bfr new_net_5873_bfr_before (
		.din(new_net_5873),
		.dout(new_net_5872)
	);

	bfr new_net_5874_bfr_before (
		.din(new_net_5874),
		.dout(new_net_5873)
	);

	bfr new_net_5875_bfr_before (
		.din(new_net_5875),
		.dout(new_net_5874)
	);

	bfr new_net_5876_bfr_before (
		.din(new_net_5876),
		.dout(new_net_5875)
	);

	bfr new_net_5877_bfr_before (
		.din(new_net_5877),
		.dout(new_net_5876)
	);

	bfr new_net_5878_bfr_before (
		.din(new_net_5878),
		.dout(new_net_5877)
	);

	bfr new_net_5879_bfr_before (
		.din(new_net_5879),
		.dout(new_net_5878)
	);

	bfr new_net_5880_bfr_before (
		.din(new_net_5880),
		.dout(new_net_5879)
	);

	bfr new_net_5881_bfr_before (
		.din(new_net_5881),
		.dout(new_net_5880)
	);

	bfr new_net_5882_bfr_before (
		.din(new_net_5882),
		.dout(new_net_5881)
	);

	bfr new_net_5883_bfr_before (
		.din(new_net_5883),
		.dout(new_net_5882)
	);

	bfr new_net_5884_bfr_before (
		.din(new_net_5884),
		.dout(new_net_5883)
	);

	bfr new_net_5885_bfr_before (
		.din(new_net_5885),
		.dout(new_net_5884)
	);

	bfr new_net_5886_bfr_before (
		.din(new_net_5886),
		.dout(new_net_5885)
	);

	bfr new_net_5887_bfr_before (
		.din(new_net_5887),
		.dout(new_net_5886)
	);

	bfr new_net_5888_bfr_before (
		.din(new_net_5888),
		.dout(new_net_5887)
	);

	bfr new_net_5889_bfr_before (
		.din(new_net_5889),
		.dout(new_net_5888)
	);

	bfr new_net_5890_bfr_before (
		.din(new_net_5890),
		.dout(new_net_5889)
	);

	bfr new_net_5891_bfr_before (
		.din(new_net_5891),
		.dout(new_net_5890)
	);

	bfr new_net_5892_bfr_before (
		.din(new_net_5892),
		.dout(new_net_5891)
	);

	bfr new_net_5893_bfr_before (
		.din(new_net_5893),
		.dout(new_net_5892)
	);

	bfr new_net_5894_bfr_before (
		.din(new_net_5894),
		.dout(new_net_5893)
	);

	bfr new_net_5895_bfr_before (
		.din(new_net_5895),
		.dout(new_net_5894)
	);

	bfr new_net_5896_bfr_before (
		.din(new_net_5896),
		.dout(new_net_5895)
	);

	bfr new_net_5897_bfr_before (
		.din(new_net_5897),
		.dout(new_net_5896)
	);

	bfr new_net_5898_bfr_before (
		.din(new_net_5898),
		.dout(new_net_5897)
	);

	bfr new_net_5899_bfr_before (
		.din(new_net_5899),
		.dout(new_net_5898)
	);

	bfr new_net_5900_bfr_before (
		.din(new_net_5900),
		.dout(new_net_5899)
	);

	bfr new_net_5901_bfr_before (
		.din(new_net_5901),
		.dout(new_net_5900)
	);

	bfr new_net_5902_bfr_before (
		.din(new_net_5902),
		.dout(new_net_5901)
	);

	bfr new_net_5903_bfr_before (
		.din(new_net_5903),
		.dout(new_net_5902)
	);

	bfr new_net_5904_bfr_before (
		.din(new_net_5904),
		.dout(new_net_5903)
	);

	bfr new_net_5905_bfr_before (
		.din(new_net_5905),
		.dout(new_net_5904)
	);

	bfr new_net_5906_bfr_before (
		.din(new_net_5906),
		.dout(new_net_5905)
	);

	bfr new_net_5907_bfr_before (
		.din(new_net_5907),
		.dout(new_net_5906)
	);

	bfr new_net_5908_bfr_before (
		.din(new_net_5908),
		.dout(new_net_5907)
	);

	bfr new_net_5909_bfr_before (
		.din(new_net_5909),
		.dout(new_net_5908)
	);

	bfr new_net_5910_bfr_before (
		.din(new_net_5910),
		.dout(new_net_5909)
	);

	bfr new_net_5911_bfr_before (
		.din(new_net_5911),
		.dout(new_net_5910)
	);

	bfr new_net_5912_bfr_before (
		.din(new_net_5912),
		.dout(new_net_5911)
	);

	bfr new_net_5913_bfr_before (
		.din(new_net_5913),
		.dout(new_net_5912)
	);

	spl3L new_net_2039_v_fanout (
		.a(new_net_2039),
		.b(new_net_5913),
		.c(new_net_1386),
		.d(new_net_1388)
	);

	spl2 n_0951__v_fanout (
		.a(n_0951_),
		.b(new_net_1446),
		.c(new_net_1445)
	);

	bfr new_net_5914_bfr_before (
		.din(new_net_5914),
		.dout(N515)
	);

	bfr new_net_5915_bfr_before (
		.din(new_net_5915),
		.dout(new_net_5914)
	);

	bfr new_net_5916_bfr_before (
		.din(new_net_5916),
		.dout(new_net_5915)
	);

	bfr new_net_5917_bfr_before (
		.din(new_net_5917),
		.dout(new_net_5916)
	);

	bfr new_net_5918_bfr_before (
		.din(new_net_5918),
		.dout(new_net_5917)
	);

	bfr new_net_5919_bfr_before (
		.din(new_net_5919),
		.dout(new_net_5918)
	);

	bfr new_net_5920_bfr_before (
		.din(new_net_5920),
		.dout(new_net_5919)
	);

	bfr new_net_5921_bfr_before (
		.din(new_net_5921),
		.dout(new_net_5920)
	);

	bfr new_net_5922_bfr_before (
		.din(new_net_5922),
		.dout(new_net_5921)
	);

	bfr new_net_5923_bfr_before (
		.din(new_net_5923),
		.dout(new_net_5922)
	);

	bfr new_net_5924_bfr_before (
		.din(new_net_5924),
		.dout(new_net_5923)
	);

	bfr new_net_5925_bfr_before (
		.din(new_net_5925),
		.dout(new_net_5924)
	);

	bfr new_net_5926_bfr_before (
		.din(new_net_5926),
		.dout(new_net_5925)
	);

	bfr new_net_5927_bfr_before (
		.din(new_net_5927),
		.dout(new_net_5926)
	);

	bfr new_net_5928_bfr_before (
		.din(new_net_5928),
		.dout(new_net_5927)
	);

	bfr new_net_5929_bfr_before (
		.din(new_net_5929),
		.dout(new_net_5928)
	);

	bfr new_net_5930_bfr_before (
		.din(new_net_5930),
		.dout(new_net_5929)
	);

	bfr new_net_5931_bfr_before (
		.din(new_net_5931),
		.dout(new_net_5930)
	);

	bfr new_net_5932_bfr_before (
		.din(new_net_5932),
		.dout(new_net_5931)
	);

	bfr new_net_5933_bfr_before (
		.din(new_net_5933),
		.dout(new_net_5932)
	);

	bfr new_net_5934_bfr_before (
		.din(new_net_5934),
		.dout(new_net_5933)
	);

	bfr new_net_5935_bfr_before (
		.din(new_net_5935),
		.dout(new_net_5934)
	);

	bfr new_net_5936_bfr_before (
		.din(new_net_5936),
		.dout(new_net_5935)
	);

	bfr new_net_5937_bfr_before (
		.din(new_net_5937),
		.dout(new_net_5936)
	);

	bfr new_net_5938_bfr_before (
		.din(new_net_5938),
		.dout(new_net_5937)
	);

	bfr new_net_5939_bfr_before (
		.din(new_net_5939),
		.dout(new_net_5938)
	);

	bfr new_net_5940_bfr_before (
		.din(new_net_5940),
		.dout(new_net_5939)
	);

	bfr new_net_5941_bfr_before (
		.din(new_net_5941),
		.dout(new_net_5940)
	);

	bfr new_net_5942_bfr_before (
		.din(new_net_5942),
		.dout(new_net_5941)
	);

	bfr new_net_5943_bfr_before (
		.din(new_net_5943),
		.dout(new_net_5942)
	);

	bfr new_net_5944_bfr_before (
		.din(new_net_5944),
		.dout(new_net_5943)
	);

	bfr new_net_5945_bfr_before (
		.din(new_net_5945),
		.dout(new_net_5944)
	);

	bfr new_net_5946_bfr_before (
		.din(new_net_5946),
		.dout(new_net_5945)
	);

	bfr new_net_5947_bfr_before (
		.din(new_net_5947),
		.dout(new_net_5946)
	);

	bfr new_net_5948_bfr_before (
		.din(new_net_5948),
		.dout(new_net_5947)
	);

	bfr new_net_5949_bfr_before (
		.din(new_net_5949),
		.dout(new_net_5948)
	);

	bfr new_net_5950_bfr_before (
		.din(new_net_5950),
		.dout(new_net_5949)
	);

	bfr new_net_5951_bfr_before (
		.din(new_net_5951),
		.dout(new_net_5950)
	);

	bfr new_net_5952_bfr_before (
		.din(new_net_5952),
		.dout(new_net_5951)
	);

	bfr new_net_5953_bfr_before (
		.din(new_net_5953),
		.dout(new_net_5952)
	);

	bfr new_net_5954_bfr_before (
		.din(new_net_5954),
		.dout(new_net_5953)
	);

	bfr new_net_5955_bfr_before (
		.din(new_net_5955),
		.dout(new_net_5954)
	);

	bfr new_net_5956_bfr_before (
		.din(new_net_5956),
		.dout(new_net_5955)
	);

	bfr new_net_5957_bfr_before (
		.din(new_net_5957),
		.dout(new_net_5956)
	);

	bfr new_net_5958_bfr_before (
		.din(new_net_5958),
		.dout(new_net_5957)
	);

	bfr new_net_5959_bfr_before (
		.din(new_net_5959),
		.dout(new_net_5958)
	);

	bfr new_net_5960_bfr_before (
		.din(new_net_5960),
		.dout(new_net_5959)
	);

	bfr new_net_5961_bfr_before (
		.din(new_net_5961),
		.dout(new_net_5960)
	);

	bfr new_net_5962_bfr_before (
		.din(new_net_5962),
		.dout(new_net_5961)
	);

	bfr new_net_5963_bfr_before (
		.din(new_net_5963),
		.dout(new_net_5962)
	);

	bfr new_net_5964_bfr_before (
		.din(new_net_5964),
		.dout(new_net_5963)
	);

	bfr new_net_5965_bfr_before (
		.din(new_net_5965),
		.dout(new_net_5964)
	);

	bfr new_net_5966_bfr_before (
		.din(new_net_5966),
		.dout(new_net_5965)
	);

	bfr new_net_5967_bfr_before (
		.din(new_net_5967),
		.dout(new_net_5966)
	);

	bfr new_net_5968_bfr_before (
		.din(new_net_5968),
		.dout(new_net_5967)
	);

	bfr new_net_5969_bfr_before (
		.din(new_net_5969),
		.dout(new_net_5968)
	);

	bfr new_net_5970_bfr_before (
		.din(new_net_5970),
		.dout(new_net_5969)
	);

	bfr new_net_5971_bfr_before (
		.din(new_net_5971),
		.dout(new_net_5970)
	);

	spl3L new_net_2032_v_fanout (
		.a(new_net_2032),
		.b(new_net_5971),
		.c(new_net_1879),
		.d(new_net_1880)
	);

	spl2 new_net_2074_v_fanout (
		.a(new_net_2074),
		.b(new_net_1882),
		.c(new_net_1884)
	);

	spl2 new_net_2092_v_fanout (
		.a(new_net_2092),
		.b(new_net_1198),
		.c(new_net_1199)
	);

	spl3L n_0720__v_fanout (
		.a(n_0720_),
		.b(new_net_649),
		.c(new_net_647),
		.d(new_net_648)
	);

	bfr new_net_5972_bfr_before (
		.din(new_net_5972),
		.dout(N509)
	);

	bfr new_net_5973_bfr_before (
		.din(new_net_5973),
		.dout(new_net_5972)
	);

	bfr new_net_5974_bfr_before (
		.din(new_net_5974),
		.dout(new_net_5973)
	);

	bfr new_net_5975_bfr_before (
		.din(new_net_5975),
		.dout(new_net_5974)
	);

	bfr new_net_5976_bfr_before (
		.din(new_net_5976),
		.dout(new_net_5975)
	);

	bfr new_net_5977_bfr_before (
		.din(new_net_5977),
		.dout(new_net_5976)
	);

	bfr new_net_5978_bfr_before (
		.din(new_net_5978),
		.dout(new_net_5977)
	);

	bfr new_net_5979_bfr_before (
		.din(new_net_5979),
		.dout(new_net_5978)
	);

	bfr new_net_5980_bfr_before (
		.din(new_net_5980),
		.dout(new_net_5979)
	);

	bfr new_net_5981_bfr_before (
		.din(new_net_5981),
		.dout(new_net_5980)
	);

	bfr new_net_5982_bfr_before (
		.din(new_net_5982),
		.dout(new_net_5981)
	);

	bfr new_net_5983_bfr_before (
		.din(new_net_5983),
		.dout(new_net_5982)
	);

	bfr new_net_5984_bfr_before (
		.din(new_net_5984),
		.dout(new_net_5983)
	);

	bfr new_net_5985_bfr_before (
		.din(new_net_5985),
		.dout(new_net_5984)
	);

	bfr new_net_5986_bfr_before (
		.din(new_net_5986),
		.dout(new_net_5985)
	);

	bfr new_net_5987_bfr_before (
		.din(new_net_5987),
		.dout(new_net_5986)
	);

	bfr new_net_5988_bfr_before (
		.din(new_net_5988),
		.dout(new_net_5987)
	);

	bfr new_net_5989_bfr_before (
		.din(new_net_5989),
		.dout(new_net_5988)
	);

	bfr new_net_5990_bfr_before (
		.din(new_net_5990),
		.dout(new_net_5989)
	);

	bfr new_net_5991_bfr_before (
		.din(new_net_5991),
		.dout(new_net_5990)
	);

	bfr new_net_5992_bfr_before (
		.din(new_net_5992),
		.dout(new_net_5991)
	);

	bfr new_net_5993_bfr_before (
		.din(new_net_5993),
		.dout(new_net_5992)
	);

	bfr new_net_5994_bfr_before (
		.din(new_net_5994),
		.dout(new_net_5993)
	);

	bfr new_net_5995_bfr_before (
		.din(new_net_5995),
		.dout(new_net_5994)
	);

	bfr new_net_5996_bfr_before (
		.din(new_net_5996),
		.dout(new_net_5995)
	);

	bfr new_net_5997_bfr_before (
		.din(new_net_5997),
		.dout(new_net_5996)
	);

	bfr new_net_5998_bfr_before (
		.din(new_net_5998),
		.dout(new_net_5997)
	);

	bfr new_net_5999_bfr_before (
		.din(new_net_5999),
		.dout(new_net_5998)
	);

	bfr new_net_6000_bfr_before (
		.din(new_net_6000),
		.dout(new_net_5999)
	);

	bfr new_net_6001_bfr_before (
		.din(new_net_6001),
		.dout(new_net_6000)
	);

	bfr new_net_6002_bfr_before (
		.din(new_net_6002),
		.dout(new_net_6001)
	);

	bfr new_net_6003_bfr_before (
		.din(new_net_6003),
		.dout(new_net_6002)
	);

	bfr new_net_6004_bfr_before (
		.din(new_net_6004),
		.dout(new_net_6003)
	);

	bfr new_net_6005_bfr_before (
		.din(new_net_6005),
		.dout(new_net_6004)
	);

	bfr new_net_6006_bfr_before (
		.din(new_net_6006),
		.dout(new_net_6005)
	);

	bfr new_net_6007_bfr_before (
		.din(new_net_6007),
		.dout(new_net_6006)
	);

	bfr new_net_6008_bfr_before (
		.din(new_net_6008),
		.dout(new_net_6007)
	);

	bfr new_net_6009_bfr_before (
		.din(new_net_6009),
		.dout(new_net_6008)
	);

	bfr new_net_6010_bfr_before (
		.din(new_net_6010),
		.dout(new_net_6009)
	);

	bfr new_net_6011_bfr_before (
		.din(new_net_6011),
		.dout(new_net_6010)
	);

	bfr new_net_6012_bfr_before (
		.din(new_net_6012),
		.dout(new_net_6011)
	);

	bfr new_net_6013_bfr_before (
		.din(new_net_6013),
		.dout(new_net_6012)
	);

	bfr new_net_6014_bfr_before (
		.din(new_net_6014),
		.dout(new_net_6013)
	);

	bfr new_net_6015_bfr_before (
		.din(new_net_6015),
		.dout(new_net_6014)
	);

	bfr new_net_6016_bfr_before (
		.din(new_net_6016),
		.dout(new_net_6015)
	);

	bfr new_net_6017_bfr_before (
		.din(new_net_6017),
		.dout(new_net_6016)
	);

	bfr new_net_6018_bfr_before (
		.din(new_net_6018),
		.dout(new_net_6017)
	);

	bfr new_net_6019_bfr_before (
		.din(new_net_6019),
		.dout(new_net_6018)
	);

	bfr new_net_6020_bfr_before (
		.din(new_net_6020),
		.dout(new_net_6019)
	);

	bfr new_net_6021_bfr_before (
		.din(new_net_6021),
		.dout(new_net_6020)
	);

	bfr new_net_6022_bfr_before (
		.din(new_net_6022),
		.dout(new_net_6021)
	);

	bfr new_net_6023_bfr_before (
		.din(new_net_6023),
		.dout(new_net_6022)
	);

	bfr new_net_6024_bfr_before (
		.din(new_net_6024),
		.dout(new_net_6023)
	);

	bfr new_net_6025_bfr_before (
		.din(new_net_6025),
		.dout(new_net_6024)
	);

	bfr new_net_6026_bfr_before (
		.din(new_net_6026),
		.dout(new_net_6025)
	);

	bfr new_net_6027_bfr_before (
		.din(new_net_6027),
		.dout(new_net_6026)
	);

	bfr new_net_6028_bfr_before (
		.din(new_net_6028),
		.dout(new_net_6027)
	);

	bfr new_net_6029_bfr_before (
		.din(new_net_6029),
		.dout(new_net_6028)
	);

	spl3L new_net_2029_v_fanout (
		.a(new_net_2029),
		.b(new_net_6029),
		.c(new_net_1459),
		.d(new_net_1458)
	);

	spl3L n_1124__v_fanout (
		.a(n_1124_),
		.b(new_net_668),
		.c(new_net_666),
		.d(new_net_667)
	);

	spl2 new_net_2076_v_fanout (
		.a(new_net_2076),
		.b(new_net_423),
		.c(new_net_424)
	);

	spl2 new_net_2075_v_fanout (
		.a(new_net_2075),
		.b(new_net_1948),
		.c(new_net_1949)
	);

	spl4L n_1253__v_fanout (
		.a(n_1253_),
		.b(new_net_732),
		.c(new_net_731),
		.d(new_net_730),
		.e(new_net_729)
	);

	spl2 new_net_2086_v_fanout (
		.a(new_net_2086),
		.b(new_net_1149),
		.c(new_net_1148)
	);

	spl4L n_1180__v_fanout (
		.a(n_1180_),
		.b(new_net_1853),
		.c(new_net_1854),
		.d(new_net_1852),
		.e(new_net_1851)
	);

	spl4L n_1153__v_fanout (
		.a(n_1153_),
		.b(new_net_823),
		.c(new_net_824),
		.d(new_net_825),
		.e(new_net_822)
	);

	spl3L n_1213__v_fanout (
		.a(n_1213_),
		.b(new_net_1043),
		.c(new_net_1041),
		.d(new_net_1042)
	);

	bfr new_net_6030_bfr_before (
		.din(new_net_6030),
		.dout(N539)
	);

	bfr new_net_6031_bfr_before (
		.din(new_net_6031),
		.dout(new_net_6030)
	);

	bfr new_net_6032_bfr_before (
		.din(new_net_6032),
		.dout(new_net_6031)
	);

	bfr new_net_6033_bfr_before (
		.din(new_net_6033),
		.dout(new_net_6032)
	);

	bfr new_net_6034_bfr_before (
		.din(new_net_6034),
		.dout(new_net_6033)
	);

	bfr new_net_6035_bfr_before (
		.din(new_net_6035),
		.dout(new_net_6034)
	);

	bfr new_net_6036_bfr_before (
		.din(new_net_6036),
		.dout(new_net_6035)
	);

	bfr new_net_6037_bfr_before (
		.din(new_net_6037),
		.dout(new_net_6036)
	);

	bfr new_net_6038_bfr_before (
		.din(new_net_6038),
		.dout(new_net_6037)
	);

	bfr new_net_6039_bfr_before (
		.din(new_net_6039),
		.dout(new_net_6038)
	);

	bfr new_net_6040_bfr_before (
		.din(new_net_6040),
		.dout(new_net_6039)
	);

	bfr new_net_6041_bfr_before (
		.din(new_net_6041),
		.dout(new_net_6040)
	);

	bfr new_net_6042_bfr_before (
		.din(new_net_6042),
		.dout(new_net_6041)
	);

	bfr new_net_6043_bfr_before (
		.din(new_net_6043),
		.dout(new_net_6042)
	);

	bfr new_net_6044_bfr_before (
		.din(new_net_6044),
		.dout(new_net_6043)
	);

	bfr new_net_6045_bfr_before (
		.din(new_net_6045),
		.dout(new_net_6044)
	);

	bfr new_net_6046_bfr_before (
		.din(new_net_6046),
		.dout(new_net_6045)
	);

	bfr new_net_6047_bfr_before (
		.din(new_net_6047),
		.dout(new_net_6046)
	);

	bfr new_net_6048_bfr_before (
		.din(new_net_6048),
		.dout(new_net_6047)
	);

	bfr new_net_6049_bfr_before (
		.din(new_net_6049),
		.dout(new_net_6048)
	);

	bfr new_net_6050_bfr_before (
		.din(new_net_6050),
		.dout(new_net_6049)
	);

	bfr new_net_6051_bfr_before (
		.din(new_net_6051),
		.dout(new_net_6050)
	);

	bfr new_net_6052_bfr_before (
		.din(new_net_6052),
		.dout(new_net_6051)
	);

	bfr new_net_6053_bfr_before (
		.din(new_net_6053),
		.dout(new_net_6052)
	);

	bfr new_net_6054_bfr_before (
		.din(new_net_6054),
		.dout(new_net_6053)
	);

	bfr new_net_6055_bfr_before (
		.din(new_net_6055),
		.dout(new_net_6054)
	);

	bfr new_net_6056_bfr_before (
		.din(new_net_6056),
		.dout(new_net_6055)
	);

	bfr new_net_6057_bfr_before (
		.din(new_net_6057),
		.dout(new_net_6056)
	);

	bfr new_net_6058_bfr_before (
		.din(new_net_6058),
		.dout(new_net_6057)
	);

	bfr new_net_6059_bfr_before (
		.din(new_net_6059),
		.dout(new_net_6058)
	);

	bfr new_net_6060_bfr_before (
		.din(new_net_6060),
		.dout(new_net_6059)
	);

	bfr new_net_6061_bfr_before (
		.din(new_net_6061),
		.dout(new_net_6060)
	);

	bfr new_net_6062_bfr_before (
		.din(new_net_6062),
		.dout(new_net_6061)
	);

	bfr new_net_6063_bfr_before (
		.din(new_net_6063),
		.dout(new_net_6062)
	);

	bfr new_net_6064_bfr_before (
		.din(new_net_6064),
		.dout(new_net_6063)
	);

	bfr new_net_6065_bfr_before (
		.din(new_net_6065),
		.dout(new_net_6064)
	);

	bfr new_net_6066_bfr_before (
		.din(new_net_6066),
		.dout(new_net_6065)
	);

	bfr new_net_6067_bfr_before (
		.din(new_net_6067),
		.dout(new_net_6066)
	);

	bfr new_net_6068_bfr_before (
		.din(new_net_6068),
		.dout(new_net_6067)
	);

	bfr new_net_6069_bfr_before (
		.din(new_net_6069),
		.dout(new_net_6068)
	);

	bfr new_net_6070_bfr_before (
		.din(new_net_6070),
		.dout(new_net_6069)
	);

	bfr new_net_6071_bfr_before (
		.din(new_net_6071),
		.dout(new_net_6070)
	);

	bfr new_net_6072_bfr_before (
		.din(new_net_6072),
		.dout(new_net_6071)
	);

	bfr new_net_6073_bfr_before (
		.din(new_net_6073),
		.dout(new_net_6072)
	);

	bfr new_net_6074_bfr_before (
		.din(new_net_6074),
		.dout(new_net_6073)
	);

	bfr new_net_6075_bfr_before (
		.din(new_net_6075),
		.dout(new_net_6074)
	);

	bfr new_net_6076_bfr_before (
		.din(new_net_6076),
		.dout(new_net_6075)
	);

	bfr new_net_6077_bfr_before (
		.din(new_net_6077),
		.dout(new_net_6076)
	);

	bfr new_net_6078_bfr_before (
		.din(new_net_6078),
		.dout(new_net_6077)
	);

	bfr new_net_6079_bfr_before (
		.din(new_net_6079),
		.dout(new_net_6078)
	);

	bfr new_net_6080_bfr_before (
		.din(new_net_6080),
		.dout(new_net_6079)
	);

	bfr new_net_6081_bfr_before (
		.din(new_net_6081),
		.dout(new_net_6080)
	);

	bfr new_net_6082_bfr_before (
		.din(new_net_6082),
		.dout(new_net_6081)
	);

	bfr new_net_6083_bfr_before (
		.din(new_net_6083),
		.dout(new_net_6082)
	);

	bfr new_net_6084_bfr_before (
		.din(new_net_6084),
		.dout(new_net_6083)
	);

	bfr new_net_6085_bfr_before (
		.din(new_net_6085),
		.dout(new_net_6084)
	);

	bfr new_net_6086_bfr_before (
		.din(new_net_6086),
		.dout(new_net_6085)
	);

	bfr new_net_6087_bfr_before (
		.din(new_net_6087),
		.dout(new_net_6086)
	);

	spl3L new_net_2037_v_fanout (
		.a(new_net_2037),
		.b(new_net_1330),
		.c(new_net_1329),
		.d(new_net_6087)
	);

	spl3L n_0730__v_fanout (
		.a(n_0730_),
		.b(new_net_1838),
		.c(new_net_1836),
		.d(new_net_1837)
	);

	spl4L n_1226__v_fanout (
		.a(n_1226_),
		.b(new_net_623),
		.c(new_net_624),
		.d(new_net_625),
		.e(new_net_622)
	);

	spl4L n_0683__v_fanout (
		.a(n_0683_),
		.b(new_net_1120),
		.c(new_net_1121),
		.d(new_net_1119),
		.e(new_net_1118)
	);

	spl4L n_0689__v_fanout (
		.a(n_0689_),
		.b(new_net_943),
		.c(new_net_944),
		.d(new_net_945),
		.e(new_net_942)
	);

	spl4L n_1165__v_fanout (
		.a(n_1165_),
		.b(new_net_88),
		.c(new_net_89),
		.d(new_net_90),
		.e(new_net_87)
	);

	spl2 new_net_2094_v_fanout (
		.a(new_net_2094),
		.b(new_net_1493),
		.c(new_net_1494)
	);

	spl2 new_net_2083_v_fanout (
		.a(new_net_2083),
		.b(new_net_1930),
		.c(new_net_1932)
	);

	bfr new_net_6088_bfr_before (
		.din(new_net_6088),
		.dout(N484)
	);

	bfr new_net_6089_bfr_before (
		.din(new_net_6089),
		.dout(new_net_6088)
	);

	bfr new_net_6090_bfr_before (
		.din(new_net_6090),
		.dout(new_net_6089)
	);

	bfr new_net_6091_bfr_before (
		.din(new_net_6091),
		.dout(new_net_6090)
	);

	bfr new_net_6092_bfr_before (
		.din(new_net_6092),
		.dout(new_net_6091)
	);

	bfr new_net_6093_bfr_before (
		.din(new_net_6093),
		.dout(new_net_6092)
	);

	bfr new_net_6094_bfr_before (
		.din(new_net_6094),
		.dout(new_net_6093)
	);

	bfr new_net_6095_bfr_before (
		.din(new_net_6095),
		.dout(new_net_6094)
	);

	bfr new_net_6096_bfr_before (
		.din(new_net_6096),
		.dout(new_net_6095)
	);

	bfr new_net_6097_bfr_before (
		.din(new_net_6097),
		.dout(new_net_6096)
	);

	bfr new_net_6098_bfr_before (
		.din(new_net_6098),
		.dout(new_net_6097)
	);

	bfr new_net_6099_bfr_before (
		.din(new_net_6099),
		.dout(new_net_6098)
	);

	bfr new_net_6100_bfr_before (
		.din(new_net_6100),
		.dout(new_net_6099)
	);

	bfr new_net_6101_bfr_before (
		.din(new_net_6101),
		.dout(new_net_6100)
	);

	bfr new_net_6102_bfr_before (
		.din(new_net_6102),
		.dout(new_net_6101)
	);

	bfr new_net_6103_bfr_before (
		.din(new_net_6103),
		.dout(new_net_6102)
	);

	bfr new_net_6104_bfr_before (
		.din(new_net_6104),
		.dout(new_net_6103)
	);

	bfr new_net_6105_bfr_before (
		.din(new_net_6105),
		.dout(new_net_6104)
	);

	bfr new_net_6106_bfr_before (
		.din(new_net_6106),
		.dout(new_net_6105)
	);

	bfr new_net_6107_bfr_before (
		.din(new_net_6107),
		.dout(new_net_6106)
	);

	bfr new_net_6108_bfr_before (
		.din(new_net_6108),
		.dout(new_net_6107)
	);

	bfr new_net_6109_bfr_before (
		.din(new_net_6109),
		.dout(new_net_6108)
	);

	bfr new_net_6110_bfr_before (
		.din(new_net_6110),
		.dout(new_net_6109)
	);

	bfr new_net_6111_bfr_before (
		.din(new_net_6111),
		.dout(new_net_6110)
	);

	bfr new_net_6112_bfr_before (
		.din(new_net_6112),
		.dout(new_net_6111)
	);

	bfr new_net_6113_bfr_before (
		.din(new_net_6113),
		.dout(new_net_6112)
	);

	bfr new_net_6114_bfr_before (
		.din(new_net_6114),
		.dout(new_net_6113)
	);

	bfr new_net_6115_bfr_before (
		.din(new_net_6115),
		.dout(new_net_6114)
	);

	bfr new_net_6116_bfr_before (
		.din(new_net_6116),
		.dout(new_net_6115)
	);

	bfr new_net_6117_bfr_before (
		.din(new_net_6117),
		.dout(new_net_6116)
	);

	bfr new_net_6118_bfr_before (
		.din(new_net_6118),
		.dout(new_net_6117)
	);

	bfr new_net_6119_bfr_before (
		.din(new_net_6119),
		.dout(new_net_6118)
	);

	bfr new_net_6120_bfr_before (
		.din(new_net_6120),
		.dout(new_net_6119)
	);

	bfr new_net_6121_bfr_before (
		.din(new_net_6121),
		.dout(new_net_6120)
	);

	bfr new_net_6122_bfr_before (
		.din(new_net_6122),
		.dout(new_net_6121)
	);

	bfr new_net_6123_bfr_before (
		.din(new_net_6123),
		.dout(new_net_6122)
	);

	bfr new_net_6124_bfr_before (
		.din(new_net_6124),
		.dout(new_net_6123)
	);

	bfr new_net_6125_bfr_before (
		.din(new_net_6125),
		.dout(new_net_6124)
	);

	bfr new_net_6126_bfr_before (
		.din(new_net_6126),
		.dout(new_net_6125)
	);

	bfr new_net_6127_bfr_before (
		.din(new_net_6127),
		.dout(new_net_6126)
	);

	bfr new_net_6128_bfr_before (
		.din(new_net_6128),
		.dout(new_net_6127)
	);

	bfr new_net_6129_bfr_before (
		.din(new_net_6129),
		.dout(new_net_6128)
	);

	bfr new_net_6130_bfr_before (
		.din(new_net_6130),
		.dout(new_net_6129)
	);

	bfr new_net_6131_bfr_before (
		.din(new_net_6131),
		.dout(new_net_6130)
	);

	bfr new_net_6132_bfr_before (
		.din(new_net_6132),
		.dout(new_net_6131)
	);

	bfr new_net_6133_bfr_before (
		.din(new_net_6133),
		.dout(new_net_6132)
	);

	bfr new_net_6134_bfr_before (
		.din(new_net_6134),
		.dout(new_net_6133)
	);

	bfr new_net_6135_bfr_before (
		.din(new_net_6135),
		.dout(new_net_6134)
	);

	bfr new_net_6136_bfr_before (
		.din(new_net_6136),
		.dout(new_net_6135)
	);

	bfr new_net_6137_bfr_before (
		.din(new_net_6137),
		.dout(new_net_6136)
	);

	bfr new_net_6138_bfr_before (
		.din(new_net_6138),
		.dout(new_net_6137)
	);

	bfr new_net_6139_bfr_before (
		.din(new_net_6139),
		.dout(new_net_6138)
	);

	bfr new_net_6140_bfr_before (
		.din(new_net_6140),
		.dout(new_net_6139)
	);

	bfr new_net_6141_bfr_before (
		.din(new_net_6141),
		.dout(new_net_6140)
	);

	bfr new_net_6142_bfr_before (
		.din(new_net_6142),
		.dout(new_net_6141)
	);

	bfr new_net_6143_bfr_before (
		.din(new_net_6143),
		.dout(new_net_6142)
	);

	bfr new_net_6144_bfr_before (
		.din(new_net_6144),
		.dout(new_net_6143)
	);

	bfr new_net_6145_bfr_before (
		.din(new_net_6145),
		.dout(new_net_6144)
	);

	spl3L new_net_2023_v_fanout (
		.a(new_net_2023),
		.b(new_net_6145),
		.c(new_net_1807),
		.d(new_net_1806)
	);

	spl2 new_net_2077_v_fanout (
		.a(new_net_2077),
		.b(new_net_1887),
		.c(new_net_1888)
	);

	spl4L n_1158__v_fanout (
		.a(n_1158_),
		.b(new_net_1321),
		.c(new_net_1322),
		.d(new_net_1323),
		.e(new_net_1320)
	);

	bfr new_net_6146_bfr_before (
		.din(new_net_6146),
		.dout(N565)
	);

	bfr new_net_6147_bfr_before (
		.din(new_net_6147),
		.dout(new_net_6146)
	);

	bfr new_net_6148_bfr_before (
		.din(new_net_6148),
		.dout(new_net_6147)
	);

	bfr new_net_6149_bfr_before (
		.din(new_net_6149),
		.dout(new_net_6148)
	);

	bfr new_net_6150_bfr_before (
		.din(new_net_6150),
		.dout(new_net_6149)
	);

	bfr new_net_6151_bfr_before (
		.din(new_net_6151),
		.dout(new_net_6150)
	);

	bfr new_net_6152_bfr_before (
		.din(new_net_6152),
		.dout(new_net_6151)
	);

	bfr new_net_6153_bfr_before (
		.din(new_net_6153),
		.dout(new_net_6152)
	);

	bfr new_net_6154_bfr_before (
		.din(new_net_6154),
		.dout(new_net_6153)
	);

	bfr new_net_6155_bfr_before (
		.din(new_net_6155),
		.dout(new_net_6154)
	);

	bfr new_net_6156_bfr_before (
		.din(new_net_6156),
		.dout(new_net_6155)
	);

	bfr new_net_6157_bfr_before (
		.din(new_net_6157),
		.dout(new_net_6156)
	);

	bfr new_net_6158_bfr_before (
		.din(new_net_6158),
		.dout(new_net_6157)
	);

	bfr new_net_6159_bfr_before (
		.din(new_net_6159),
		.dout(new_net_6158)
	);

	bfr new_net_6160_bfr_before (
		.din(new_net_6160),
		.dout(new_net_6159)
	);

	bfr new_net_6161_bfr_before (
		.din(new_net_6161),
		.dout(new_net_6160)
	);

	bfr new_net_6162_bfr_before (
		.din(new_net_6162),
		.dout(new_net_6161)
	);

	bfr new_net_6163_bfr_before (
		.din(new_net_6163),
		.dout(new_net_6162)
	);

	bfr new_net_6164_bfr_before (
		.din(new_net_6164),
		.dout(new_net_6163)
	);

	bfr new_net_6165_bfr_before (
		.din(new_net_6165),
		.dout(new_net_6164)
	);

	bfr new_net_6166_bfr_before (
		.din(new_net_6166),
		.dout(new_net_6165)
	);

	bfr new_net_6167_bfr_before (
		.din(new_net_6167),
		.dout(new_net_6166)
	);

	bfr new_net_6168_bfr_before (
		.din(new_net_6168),
		.dout(new_net_6167)
	);

	bfr new_net_6169_bfr_before (
		.din(new_net_6169),
		.dout(new_net_6168)
	);

	bfr new_net_6170_bfr_before (
		.din(new_net_6170),
		.dout(new_net_6169)
	);

	bfr new_net_6171_bfr_before (
		.din(new_net_6171),
		.dout(new_net_6170)
	);

	bfr new_net_6172_bfr_before (
		.din(new_net_6172),
		.dout(new_net_6171)
	);

	bfr new_net_6173_bfr_before (
		.din(new_net_6173),
		.dout(new_net_6172)
	);

	bfr new_net_6174_bfr_before (
		.din(new_net_6174),
		.dout(new_net_6173)
	);

	bfr new_net_6175_bfr_before (
		.din(new_net_6175),
		.dout(new_net_6174)
	);

	bfr new_net_6176_bfr_before (
		.din(new_net_6176),
		.dout(new_net_6175)
	);

	bfr new_net_6177_bfr_before (
		.din(new_net_6177),
		.dout(new_net_6176)
	);

	bfr new_net_6178_bfr_before (
		.din(new_net_6178),
		.dout(new_net_6177)
	);

	bfr new_net_6179_bfr_before (
		.din(new_net_6179),
		.dout(new_net_6178)
	);

	bfr new_net_6180_bfr_before (
		.din(new_net_6180),
		.dout(new_net_6179)
	);

	bfr new_net_6181_bfr_before (
		.din(new_net_6181),
		.dout(new_net_6180)
	);

	bfr new_net_6182_bfr_before (
		.din(new_net_6182),
		.dout(new_net_6181)
	);

	bfr new_net_6183_bfr_before (
		.din(new_net_6183),
		.dout(new_net_6182)
	);

	bfr new_net_6184_bfr_before (
		.din(new_net_6184),
		.dout(new_net_6183)
	);

	bfr new_net_6185_bfr_before (
		.din(new_net_6185),
		.dout(new_net_6184)
	);

	bfr new_net_6186_bfr_before (
		.din(new_net_6186),
		.dout(new_net_6185)
	);

	bfr new_net_6187_bfr_before (
		.din(new_net_6187),
		.dout(new_net_6186)
	);

	bfr new_net_6188_bfr_before (
		.din(new_net_6188),
		.dout(new_net_6187)
	);

	bfr new_net_6189_bfr_before (
		.din(new_net_6189),
		.dout(new_net_6188)
	);

	bfr new_net_6190_bfr_before (
		.din(new_net_6190),
		.dout(new_net_6189)
	);

	bfr new_net_6191_bfr_before (
		.din(new_net_6191),
		.dout(new_net_6190)
	);

	bfr new_net_6192_bfr_before (
		.din(new_net_6192),
		.dout(new_net_6191)
	);

	bfr new_net_6193_bfr_before (
		.din(new_net_6193),
		.dout(new_net_6192)
	);

	bfr new_net_6194_bfr_before (
		.din(new_net_6194),
		.dout(new_net_6193)
	);

	bfr new_net_6195_bfr_before (
		.din(new_net_6195),
		.dout(new_net_6194)
	);

	bfr new_net_6196_bfr_before (
		.din(new_net_6196),
		.dout(new_net_6195)
	);

	bfr new_net_6197_bfr_before (
		.din(new_net_6197),
		.dout(new_net_6196)
	);

	bfr new_net_6198_bfr_before (
		.din(new_net_6198),
		.dout(new_net_6197)
	);

	bfr new_net_6199_bfr_before (
		.din(new_net_6199),
		.dout(new_net_6198)
	);

	bfr new_net_6200_bfr_before (
		.din(new_net_6200),
		.dout(new_net_6199)
	);

	bfr new_net_6201_bfr_before (
		.din(new_net_6201),
		.dout(new_net_6200)
	);

	bfr new_net_6202_bfr_before (
		.din(new_net_6202),
		.dout(new_net_6201)
	);

	bfr new_net_6203_bfr_before (
		.din(new_net_6203),
		.dout(new_net_6202)
	);

	spl3L new_net_2049_v_fanout (
		.a(new_net_2049),
		.b(new_net_1660),
		.c(new_net_1662),
		.d(new_net_6203)
	);

	spl2 n_1246__v_fanout (
		.a(n_1246_),
		.b(new_net_1127),
		.c(new_net_1126)
	);

	spl3L n_1018__v_fanout (
		.a(n_1018_),
		.b(new_net_1245),
		.c(new_net_1244),
		.d(new_net_2085)
	);

	spl3L n_1030__v_fanout (
		.a(n_1030_),
		.b(new_net_2087),
		.c(new_net_748),
		.d(new_net_749)
	);

	bfr new_net_6204_bfr_after (
		.din(n_0665_),
		.dout(new_net_6204)
	);

	bfr new_net_6205_bfr_before (
		.din(new_net_6205),
		.dout(new_net_2069)
	);

	spl2 n_0665__v_fanout (
		.a(new_net_6204),
		.b(new_net_6205),
		.c(new_net_1611)
	);

	spl3L n_1066__v_fanout (
		.a(n_1066_),
		.b(new_net_2092),
		.c(new_net_1196),
		.d(new_net_1197)
	);

	spl3L n_0915__v_fanout (
		.a(n_0915_),
		.b(new_net_1584),
		.c(new_net_1582),
		.d(new_net_2071)
	);

	spl4L n_1069__v_fanout (
		.a(n_1069_),
		.b(new_net_540),
		.c(new_net_541),
		.d(new_net_539),
		.e(new_net_538)
	);

	bfr new_net_6206_bfr_after (
		.din(n_0987_),
		.dout(new_net_6206)
	);

	bfr new_net_6207_bfr_before (
		.din(new_net_6207),
		.dout(new_net_2080)
	);

	spl3L n_0987__v_fanout (
		.a(new_net_6206),
		.b(new_net_1393),
		.c(new_net_6207),
		.d(new_net_1394)
	);

	spl3L n_1033__v_fanout (
		.a(n_1033_),
		.b(new_net_1091),
		.c(new_net_1089),
		.d(new_net_2088)
	);

	spl3L n_0972__v_fanout (
		.a(n_0972_),
		.b(new_net_2077),
		.c(new_net_1885),
		.d(new_net_1886)
	);

	spl3L n_1075__v_fanout (
		.a(n_1075_),
		.b(new_net_2093),
		.c(new_net_1409),
		.d(new_net_1410)
	);

	spl3L n_1012__v_fanout (
		.a(n_1012_),
		.b(new_net_977),
		.c(new_net_974),
		.d(new_net_2084)
	);

	bfr new_net_6208_bfr_after (
		.din(n_0954_),
		.dout(new_net_6208)
	);

	spl2 n_0954__v_fanout (
		.a(new_net_6208),
		.b(new_net_1289),
		.c(new_net_1288)
	);

	spl3L n_1054__v_fanout (
		.a(n_1054_),
		.b(new_net_1491),
		.c(new_net_1488),
		.d(new_net_2091)
	);

	spl3L n_0960__v_fanout (
		.a(n_0960_),
		.b(new_net_2075),
		.c(new_net_1947),
		.d(new_net_1950)
	);

	spl3L n_0990__v_fanout (
		.a(n_0990_),
		.b(new_net_2081),
		.c(new_net_488),
		.d(new_net_491)
	);

	spl3L n_1021__v_fanout (
		.a(n_1021_),
		.b(new_net_2086),
		.c(new_net_1147),
		.d(new_net_1150)
	);

	spl3L n_0930__v_fanout (
		.a(n_0930_),
		.b(new_net_2074),
		.c(new_net_1881),
		.d(new_net_1883)
	);

	spl2 n_1051__v_fanout (
		.a(n_1051_),
		.b(new_net_1163),
		.c(new_net_1162)
	);

	spl3L n_1105__v_fanout (
		.a(n_1105_),
		.b(new_net_2098),
		.c(new_net_63),
		.d(new_net_65)
	);

	bfr new_net_6209_bfr_after (
		.din(n_1096_),
		.dout(new_net_6209)
	);

	bfr new_net_6210_bfr_before (
		.din(new_net_6210),
		.dout(new_net_2096)
	);

	spl3L n_1096__v_fanout (
		.a(new_net_6209),
		.b(new_net_1827),
		.c(new_net_6210),
		.d(new_net_1826)
	);

	spl3L n_0752__v_fanout (
		.a(n_0752_),
		.b(new_net_796),
		.c(new_net_2070),
		.d(new_net_794)
	);

	bfr new_net_6211_bfr_after (
		.din(n_1111_),
		.dout(new_net_6211)
	);

	bfr new_net_6212_bfr_before (
		.din(new_net_6212),
		.dout(new_net_2099)
	);

	spl3L n_1111__v_fanout (
		.a(new_net_6211),
		.b(new_net_321),
		.c(new_net_6212),
		.d(new_net_320)
	);

	spl3L n_1228__v_fanout (
		.a(n_1228_),
		.b(new_net_1016),
		.c(new_net_2100),
		.d(new_net_1015)
	);

	spl3L n_0918__v_fanout (
		.a(n_0918_),
		.b(new_net_2072),
		.c(new_net_1797),
		.d(new_net_1799)
	);

	spl3L n_1009__v_fanout (
		.a(n_1009_),
		.b(new_net_2083),
		.c(new_net_1929),
		.d(new_net_1931)
	);

	spl3L n_1102__v_fanout (
		.a(n_1102_),
		.b(new_net_2097),
		.c(new_net_637),
		.d(new_net_638)
	);

	spl4L n_0909__v_fanout (
		.a(n_0909_),
		.b(new_net_1442),
		.c(new_net_1440),
		.d(new_net_1441),
		.e(new_net_1439)
	);

	bfr new_net_6213_bfr_after (
		.din(n_0169_),
		.dout(new_net_6213)
	);

	bfr new_net_6214_bfr_after (
		.din(new_net_6213),
		.dout(new_net_6214)
	);

	bfr new_net_6215_bfr_after (
		.din(new_net_6214),
		.dout(new_net_6215)
	);

	bfr new_net_6216_bfr_after (
		.din(new_net_6215),
		.dout(new_net_6216)
	);

	bfr new_net_6217_bfr_after (
		.din(new_net_6216),
		.dout(new_net_6217)
	);

	bfr new_net_6218_bfr_after (
		.din(new_net_6217),
		.dout(new_net_6218)
	);

	bfr new_net_6219_bfr_after (
		.din(new_net_6218),
		.dout(new_net_6219)
	);

	bfr new_net_6220_bfr_after (
		.din(new_net_6219),
		.dout(new_net_6220)
	);

	bfr new_net_6221_bfr_after (
		.din(new_net_6220),
		.dout(new_net_6221)
	);

	bfr new_net_6222_bfr_after (
		.din(new_net_6221),
		.dout(new_net_6222)
	);

	bfr new_net_6223_bfr_after (
		.din(new_net_6222),
		.dout(new_net_6223)
	);

	bfr new_net_6224_bfr_after (
		.din(new_net_6223),
		.dout(new_net_6224)
	);

	bfr new_net_6225_bfr_after (
		.din(new_net_6224),
		.dout(new_net_6225)
	);

	bfr new_net_6226_bfr_after (
		.din(new_net_6225),
		.dout(new_net_6226)
	);

	bfr new_net_6227_bfr_after (
		.din(new_net_6226),
		.dout(new_net_6227)
	);

	bfr new_net_6228_bfr_after (
		.din(new_net_6227),
		.dout(new_net_6228)
	);

	bfr new_net_6229_bfr_after (
		.din(new_net_6228),
		.dout(new_net_6229)
	);

	bfr new_net_6230_bfr_after (
		.din(new_net_6229),
		.dout(new_net_6230)
	);

	bfr new_net_6231_bfr_after (
		.din(new_net_6230),
		.dout(new_net_6231)
	);

	bfr new_net_6232_bfr_after (
		.din(new_net_6231),
		.dout(new_net_6232)
	);

	bfr new_net_6233_bfr_after (
		.din(new_net_6232),
		.dout(new_net_6233)
	);

	bfr new_net_6234_bfr_after (
		.din(new_net_6233),
		.dout(new_net_6234)
	);

	bfr new_net_6235_bfr_after (
		.din(new_net_6234),
		.dout(new_net_6235)
	);

	bfr new_net_6236_bfr_after (
		.din(new_net_6235),
		.dout(new_net_6236)
	);

	bfr new_net_6237_bfr_after (
		.din(new_net_6236),
		.dout(new_net_6237)
	);

	bfr new_net_6238_bfr_after (
		.din(new_net_6237),
		.dout(new_net_6238)
	);

	bfr new_net_6239_bfr_after (
		.din(new_net_6238),
		.dout(new_net_6239)
	);

	bfr new_net_6240_bfr_after (
		.din(new_net_6239),
		.dout(new_net_6240)
	);

	bfr new_net_6241_bfr_after (
		.din(new_net_6240),
		.dout(new_net_6241)
	);

	bfr new_net_6242_bfr_after (
		.din(new_net_6241),
		.dout(new_net_6242)
	);

	bfr new_net_6243_bfr_after (
		.din(new_net_6242),
		.dout(new_net_6243)
	);

	bfr new_net_6244_bfr_after (
		.din(new_net_6243),
		.dout(new_net_6244)
	);

	bfr new_net_6245_bfr_after (
		.din(new_net_6244),
		.dout(new_net_6245)
	);

	bfr new_net_6246_bfr_after (
		.din(new_net_6245),
		.dout(new_net_6246)
	);

	bfr new_net_6247_bfr_after (
		.din(new_net_6246),
		.dout(new_net_6247)
	);

	bfr new_net_6248_bfr_after (
		.din(new_net_6247),
		.dout(new_net_6248)
	);

	bfr new_net_6249_bfr_after (
		.din(new_net_6248),
		.dout(new_net_6249)
	);

	bfr new_net_6250_bfr_after (
		.din(new_net_6249),
		.dout(new_net_6250)
	);

	bfr new_net_6251_bfr_after (
		.din(new_net_6250),
		.dout(new_net_6251)
	);

	bfr new_net_6252_bfr_after (
		.din(new_net_6251),
		.dout(new_net_6252)
	);

	bfr new_net_6253_bfr_after (
		.din(new_net_6252),
		.dout(new_net_6253)
	);

	bfr new_net_6254_bfr_after (
		.din(new_net_6253),
		.dout(new_net_6254)
	);

	bfr new_net_6255_bfr_after (
		.din(new_net_6254),
		.dout(new_net_6255)
	);

	bfr new_net_6256_bfr_after (
		.din(new_net_6255),
		.dout(new_net_6256)
	);

	bfr new_net_6257_bfr_after (
		.din(new_net_6256),
		.dout(new_net_6257)
	);

	bfr new_net_6258_bfr_after (
		.din(new_net_6257),
		.dout(new_net_6258)
	);

	bfr new_net_6259_bfr_after (
		.din(new_net_6258),
		.dout(new_net_6259)
	);

	bfr new_net_6260_bfr_after (
		.din(new_net_6259),
		.dout(new_net_6260)
	);

	bfr new_net_6261_bfr_after (
		.din(new_net_6260),
		.dout(new_net_6261)
	);

	bfr new_net_6262_bfr_after (
		.din(new_net_6261),
		.dout(new_net_6262)
	);

	bfr new_net_6263_bfr_after (
		.din(new_net_6262),
		.dout(new_net_6263)
	);

	bfr new_net_6264_bfr_after (
		.din(new_net_6263),
		.dout(new_net_6264)
	);

	bfr new_net_6265_bfr_after (
		.din(new_net_6264),
		.dout(new_net_6265)
	);

	spl2 n_0169__v_fanout (
		.a(new_net_6265),
		.b(new_net_1115),
		.c(new_net_1114)
	);

	spl2 n_0906__v_fanout (
		.a(n_0906_),
		.b(new_net_554),
		.c(new_net_553)
	);

	spl3L n_0927__v_fanout (
		.a(n_0927_),
		.b(new_net_998),
		.c(new_net_996),
		.d(new_net_2073)
	);

	spl3L n_1045__v_fanout (
		.a(n_1045_),
		.b(new_net_2090),
		.c(new_net_524),
		.d(new_net_527)
	);

	spl2 new_net_2064_v_fanout (
		.a(new_net_2064),
		.b(new_net_382),
		.c(new_net_373)
	);

	spl3L n_0963__v_fanout (
		.a(n_0963_),
		.b(new_net_425),
		.c(new_net_422),
		.d(new_net_2076)
	);

	bfr new_net_6266_bfr_after (
		.din(n_0981_),
		.dout(new_net_6266)
	);

	bfr new_net_6267_bfr_before (
		.din(new_net_6267),
		.dout(new_net_2079)
	);

	spl3L n_0981__v_fanout (
		.a(new_net_6266),
		.b(new_net_767),
		.c(new_net_6267),
		.d(new_net_765)
	);

	spl2 n_1087__v_fanout (
		.a(n_1087_),
		.b(new_net_1649),
		.c(new_net_1648)
	);

	spl3L n_0788__v_fanout (
		.a(n_0788_),
		.b(new_net_1019),
		.c(new_net_1017),
		.d(new_net_1018)
	);

	spl3L n_1090__v_fanout (
		.a(n_1090_),
		.b(new_net_983),
		.c(new_net_980),
		.d(new_net_2095)
	);

	spl3L n_1042__v_fanout (
		.a(n_1042_),
		.b(new_net_2089),
		.c(new_net_1601),
		.d(new_net_1602)
	);

	spl3L n_1078__v_fanout (
		.a(n_1078_),
		.b(new_net_2094),
		.c(new_net_1492),
		.d(new_net_1495)
	);

	bfr new_net_6268_bfr_before (
		.din(new_net_6268),
		.dout(N511)
	);

	bfr new_net_6269_bfr_before (
		.din(new_net_6269),
		.dout(new_net_6268)
	);

	bfr new_net_6270_bfr_before (
		.din(new_net_6270),
		.dout(new_net_6269)
	);

	bfr new_net_6271_bfr_before (
		.din(new_net_6271),
		.dout(new_net_6270)
	);

	bfr new_net_6272_bfr_before (
		.din(new_net_6272),
		.dout(new_net_6271)
	);

	bfr new_net_6273_bfr_before (
		.din(new_net_6273),
		.dout(new_net_6272)
	);

	bfr new_net_6274_bfr_before (
		.din(new_net_6274),
		.dout(new_net_6273)
	);

	bfr new_net_6275_bfr_before (
		.din(new_net_6275),
		.dout(new_net_6274)
	);

	bfr new_net_6276_bfr_before (
		.din(new_net_6276),
		.dout(new_net_6275)
	);

	bfr new_net_6277_bfr_before (
		.din(new_net_6277),
		.dout(new_net_6276)
	);

	bfr new_net_6278_bfr_before (
		.din(new_net_6278),
		.dout(new_net_6277)
	);

	bfr new_net_6279_bfr_before (
		.din(new_net_6279),
		.dout(new_net_6278)
	);

	bfr new_net_6280_bfr_before (
		.din(new_net_6280),
		.dout(new_net_6279)
	);

	bfr new_net_6281_bfr_before (
		.din(new_net_6281),
		.dout(new_net_6280)
	);

	bfr new_net_6282_bfr_before (
		.din(new_net_6282),
		.dout(new_net_6281)
	);

	bfr new_net_6283_bfr_before (
		.din(new_net_6283),
		.dout(new_net_6282)
	);

	bfr new_net_6284_bfr_before (
		.din(new_net_6284),
		.dout(new_net_6283)
	);

	bfr new_net_6285_bfr_before (
		.din(new_net_6285),
		.dout(new_net_6284)
	);

	bfr new_net_6286_bfr_before (
		.din(new_net_6286),
		.dout(new_net_6285)
	);

	bfr new_net_6287_bfr_before (
		.din(new_net_6287),
		.dout(new_net_6286)
	);

	bfr new_net_6288_bfr_before (
		.din(new_net_6288),
		.dout(new_net_6287)
	);

	bfr new_net_6289_bfr_before (
		.din(new_net_6289),
		.dout(new_net_6288)
	);

	bfr new_net_6290_bfr_before (
		.din(new_net_6290),
		.dout(new_net_6289)
	);

	bfr new_net_6291_bfr_before (
		.din(new_net_6291),
		.dout(new_net_6290)
	);

	bfr new_net_6292_bfr_before (
		.din(new_net_6292),
		.dout(new_net_6291)
	);

	bfr new_net_6293_bfr_before (
		.din(new_net_6293),
		.dout(new_net_6292)
	);

	bfr new_net_6294_bfr_before (
		.din(new_net_6294),
		.dout(new_net_6293)
	);

	bfr new_net_6295_bfr_before (
		.din(new_net_6295),
		.dout(new_net_6294)
	);

	bfr new_net_6296_bfr_before (
		.din(new_net_6296),
		.dout(new_net_6295)
	);

	bfr new_net_6297_bfr_before (
		.din(new_net_6297),
		.dout(new_net_6296)
	);

	bfr new_net_6298_bfr_before (
		.din(new_net_6298),
		.dout(new_net_6297)
	);

	bfr new_net_6299_bfr_before (
		.din(new_net_6299),
		.dout(new_net_6298)
	);

	bfr new_net_6300_bfr_before (
		.din(new_net_6300),
		.dout(new_net_6299)
	);

	bfr new_net_6301_bfr_before (
		.din(new_net_6301),
		.dout(new_net_6300)
	);

	bfr new_net_6302_bfr_before (
		.din(new_net_6302),
		.dout(new_net_6301)
	);

	bfr new_net_6303_bfr_before (
		.din(new_net_6303),
		.dout(new_net_6302)
	);

	bfr new_net_6304_bfr_before (
		.din(new_net_6304),
		.dout(new_net_6303)
	);

	bfr new_net_6305_bfr_before (
		.din(new_net_6305),
		.dout(new_net_6304)
	);

	bfr new_net_6306_bfr_before (
		.din(new_net_6306),
		.dout(new_net_6305)
	);

	bfr new_net_6307_bfr_before (
		.din(new_net_6307),
		.dout(new_net_6306)
	);

	bfr new_net_6308_bfr_before (
		.din(new_net_6308),
		.dout(new_net_6307)
	);

	bfr new_net_6309_bfr_before (
		.din(new_net_6309),
		.dout(new_net_6308)
	);

	bfr new_net_6310_bfr_before (
		.din(new_net_6310),
		.dout(new_net_6309)
	);

	bfr new_net_6311_bfr_before (
		.din(new_net_6311),
		.dout(new_net_6310)
	);

	bfr new_net_6312_bfr_before (
		.din(new_net_6312),
		.dout(new_net_6311)
	);

	bfr new_net_6313_bfr_before (
		.din(new_net_6313),
		.dout(new_net_6312)
	);

	bfr new_net_6314_bfr_before (
		.din(new_net_6314),
		.dout(new_net_6313)
	);

	bfr new_net_6315_bfr_before (
		.din(new_net_6315),
		.dout(new_net_6314)
	);

	bfr new_net_6316_bfr_before (
		.din(new_net_6316),
		.dout(new_net_6315)
	);

	bfr new_net_6317_bfr_before (
		.din(new_net_6317),
		.dout(new_net_6316)
	);

	bfr new_net_6318_bfr_before (
		.din(new_net_6318),
		.dout(new_net_6317)
	);

	bfr new_net_6319_bfr_before (
		.din(new_net_6319),
		.dout(new_net_6318)
	);

	bfr new_net_6320_bfr_before (
		.din(new_net_6320),
		.dout(new_net_6319)
	);

	bfr new_net_6321_bfr_before (
		.din(new_net_6321),
		.dout(new_net_6320)
	);

	bfr new_net_6322_bfr_before (
		.din(new_net_6322),
		.dout(new_net_6321)
	);

	bfr new_net_6323_bfr_before (
		.din(new_net_6323),
		.dout(new_net_6322)
	);

	bfr new_net_6324_bfr_before (
		.din(new_net_6324),
		.dout(new_net_6323)
	);

	bfr new_net_6325_bfr_before (
		.din(new_net_6325),
		.dout(new_net_6324)
	);

	bfr new_net_6326_bfr_before (
		.din(new_net_6326),
		.dout(new_net_6325)
	);

	spl3L new_net_2030_v_fanout (
		.a(new_net_2030),
		.b(new_net_1578),
		.c(new_net_1576),
		.d(new_net_6326)
	);

	spl3L n_0975__v_fanout (
		.a(n_0975_),
		.b(new_net_2078),
		.c(new_net_1925),
		.d(new_net_1928)
	);

	spl3L n_0993__v_fanout (
		.a(n_0993_),
		.b(new_net_44),
		.c(new_net_41),
		.d(new_net_2082)
	);

	spl2 n_0856__v_fanout (
		.a(n_0856_),
		.b(new_net_434),
		.c(new_net_433)
	);

	spl2 n_0850__v_fanout (
		.a(n_0850_),
		.b(new_net_1620),
		.c(new_net_1619)
	);

	spl4L n_0662__v_fanout (
		.a(n_0662_),
		.b(new_net_643),
		.c(new_net_644),
		.d(new_net_642),
		.e(new_net_641)
	);

	bfr new_net_6327_bfr_before (
		.din(new_net_6327),
		.dout(new_net_1508)
	);

	bfr new_net_6328_bfr_before (
		.din(new_net_6328),
		.dout(new_net_6327)
	);

	spl2 n_1205__v_fanout (
		.a(n_1205_),
		.b(new_net_6328),
		.c(new_net_1507)
	);

	spl2 n_0877__v_fanout (
		.a(n_0877_),
		.b(new_net_775),
		.c(new_net_774)
	);

	bfr new_net_6329_bfr_before (
		.din(new_net_6329),
		.dout(N537)
	);

	bfr new_net_6330_bfr_before (
		.din(new_net_6330),
		.dout(new_net_6329)
	);

	bfr new_net_6331_bfr_before (
		.din(new_net_6331),
		.dout(new_net_6330)
	);

	bfr new_net_6332_bfr_before (
		.din(new_net_6332),
		.dout(new_net_6331)
	);

	bfr new_net_6333_bfr_before (
		.din(new_net_6333),
		.dout(new_net_6332)
	);

	bfr new_net_6334_bfr_before (
		.din(new_net_6334),
		.dout(new_net_6333)
	);

	bfr new_net_6335_bfr_before (
		.din(new_net_6335),
		.dout(new_net_6334)
	);

	bfr new_net_6336_bfr_before (
		.din(new_net_6336),
		.dout(new_net_6335)
	);

	bfr new_net_6337_bfr_before (
		.din(new_net_6337),
		.dout(new_net_6336)
	);

	bfr new_net_6338_bfr_before (
		.din(new_net_6338),
		.dout(new_net_6337)
	);

	bfr new_net_6339_bfr_before (
		.din(new_net_6339),
		.dout(new_net_6338)
	);

	bfr new_net_6340_bfr_before (
		.din(new_net_6340),
		.dout(new_net_6339)
	);

	bfr new_net_6341_bfr_before (
		.din(new_net_6341),
		.dout(new_net_6340)
	);

	bfr new_net_6342_bfr_before (
		.din(new_net_6342),
		.dout(new_net_6341)
	);

	bfr new_net_6343_bfr_before (
		.din(new_net_6343),
		.dout(new_net_6342)
	);

	bfr new_net_6344_bfr_before (
		.din(new_net_6344),
		.dout(new_net_6343)
	);

	bfr new_net_6345_bfr_before (
		.din(new_net_6345),
		.dout(new_net_6344)
	);

	bfr new_net_6346_bfr_before (
		.din(new_net_6346),
		.dout(new_net_6345)
	);

	bfr new_net_6347_bfr_before (
		.din(new_net_6347),
		.dout(new_net_6346)
	);

	bfr new_net_6348_bfr_before (
		.din(new_net_6348),
		.dout(new_net_6347)
	);

	bfr new_net_6349_bfr_before (
		.din(new_net_6349),
		.dout(new_net_6348)
	);

	bfr new_net_6350_bfr_before (
		.din(new_net_6350),
		.dout(new_net_6349)
	);

	bfr new_net_6351_bfr_before (
		.din(new_net_6351),
		.dout(new_net_6350)
	);

	bfr new_net_6352_bfr_before (
		.din(new_net_6352),
		.dout(new_net_6351)
	);

	bfr new_net_6353_bfr_before (
		.din(new_net_6353),
		.dout(new_net_6352)
	);

	bfr new_net_6354_bfr_before (
		.din(new_net_6354),
		.dout(new_net_6353)
	);

	bfr new_net_6355_bfr_before (
		.din(new_net_6355),
		.dout(new_net_6354)
	);

	bfr new_net_6356_bfr_before (
		.din(new_net_6356),
		.dout(new_net_6355)
	);

	bfr new_net_6357_bfr_before (
		.din(new_net_6357),
		.dout(new_net_6356)
	);

	bfr new_net_6358_bfr_before (
		.din(new_net_6358),
		.dout(new_net_6357)
	);

	bfr new_net_6359_bfr_before (
		.din(new_net_6359),
		.dout(new_net_6358)
	);

	bfr new_net_6360_bfr_before (
		.din(new_net_6360),
		.dout(new_net_6359)
	);

	bfr new_net_6361_bfr_before (
		.din(new_net_6361),
		.dout(new_net_6360)
	);

	bfr new_net_6362_bfr_before (
		.din(new_net_6362),
		.dout(new_net_6361)
	);

	bfr new_net_6363_bfr_before (
		.din(new_net_6363),
		.dout(new_net_6362)
	);

	bfr new_net_6364_bfr_before (
		.din(new_net_6364),
		.dout(new_net_6363)
	);

	bfr new_net_6365_bfr_before (
		.din(new_net_6365),
		.dout(new_net_6364)
	);

	bfr new_net_6366_bfr_before (
		.din(new_net_6366),
		.dout(new_net_6365)
	);

	bfr new_net_6367_bfr_before (
		.din(new_net_6367),
		.dout(new_net_6366)
	);

	bfr new_net_6368_bfr_before (
		.din(new_net_6368),
		.dout(new_net_6367)
	);

	bfr new_net_6369_bfr_before (
		.din(new_net_6369),
		.dout(new_net_6368)
	);

	bfr new_net_6370_bfr_before (
		.din(new_net_6370),
		.dout(new_net_6369)
	);

	bfr new_net_6371_bfr_before (
		.din(new_net_6371),
		.dout(new_net_6370)
	);

	bfr new_net_6372_bfr_before (
		.din(new_net_6372),
		.dout(new_net_6371)
	);

	bfr new_net_6373_bfr_before (
		.din(new_net_6373),
		.dout(new_net_6372)
	);

	bfr new_net_6374_bfr_before (
		.din(new_net_6374),
		.dout(new_net_6373)
	);

	bfr new_net_6375_bfr_before (
		.din(new_net_6375),
		.dout(new_net_6374)
	);

	bfr new_net_6376_bfr_before (
		.din(new_net_6376),
		.dout(new_net_6375)
	);

	bfr new_net_6377_bfr_before (
		.din(new_net_6377),
		.dout(new_net_6376)
	);

	bfr new_net_6378_bfr_before (
		.din(new_net_6378),
		.dout(new_net_6377)
	);

	bfr new_net_6379_bfr_before (
		.din(new_net_6379),
		.dout(new_net_6378)
	);

	bfr new_net_6380_bfr_before (
		.din(new_net_6380),
		.dout(new_net_6379)
	);

	bfr new_net_6381_bfr_before (
		.din(new_net_6381),
		.dout(new_net_6380)
	);

	bfr new_net_6382_bfr_before (
		.din(new_net_6382),
		.dout(new_net_6381)
	);

	bfr new_net_6383_bfr_before (
		.din(new_net_6383),
		.dout(new_net_6382)
	);

	bfr new_net_6384_bfr_before (
		.din(new_net_6384),
		.dout(new_net_6383)
	);

	bfr new_net_6385_bfr_before (
		.din(new_net_6385),
		.dout(new_net_6384)
	);

	bfr new_net_6386_bfr_before (
		.din(new_net_6386),
		.dout(new_net_6385)
	);

	bfr new_net_6387_bfr_before (
		.din(new_net_6387),
		.dout(new_net_6386)
	);

	bfr new_net_6388_bfr_before (
		.din(new_net_6388),
		.dout(new_net_6387)
	);

	spl2 new_net_2036_v_fanout (
		.a(new_net_2036),
		.b(new_net_6388),
		.c(new_net_511)
	);

	bfr new_net_6389_bfr_before (
		.din(new_net_6389),
		.dout(new_net_79)
	);

	bfr new_net_6390_bfr_before (
		.din(new_net_6390),
		.dout(new_net_6389)
	);

	spl2 n_0728__v_fanout (
		.a(n_0728_),
		.b(new_net_80),
		.c(new_net_6390)
	);

	spl2 n_0733__v_fanout (
		.a(n_0733_),
		.b(new_net_339),
		.c(new_net_338)
	);

	spl2 n_0859__v_fanout (
		.a(n_0859_),
		.b(new_net_328),
		.c(new_net_327)
	);

	spl2 n_0832__v_fanout (
		.a(n_0832_),
		.b(new_net_1317),
		.c(new_net_1316)
	);

	spl2 n_0847__v_fanout (
		.a(n_0847_),
		.b(new_net_1920),
		.c(new_net_1919)
	);

	spl2 n_0880__v_fanout (
		.a(n_0880_),
		.b(new_net_842),
		.c(new_net_841)
	);

	spl2 n_0748__v_fanout (
		.a(n_0748_),
		.b(new_net_716),
		.c(new_net_715)
	);

	spl2 n_0889__v_fanout (
		.a(n_0889_),
		.b(new_net_1027),
		.c(new_net_1026)
	);

	spl2 n_0756__v_fanout (
		.a(n_0756_),
		.b(new_net_872),
		.c(new_net_871)
	);

	spl2 n_0769__v_fanout (
		.a(n_0769_),
		.b(new_net_808),
		.c(new_net_807)
	);

	spl2 n_0759__v_fanout (
		.a(n_0759_),
		.b(new_net_939),
		.c(new_net_938)
	);

	bfr new_net_6391_bfr_before (
		.din(new_net_6391),
		.dout(new_net_1443)
	);

	bfr new_net_6392_bfr_before (
		.din(new_net_6392),
		.dout(new_net_6391)
	);

	spl2 n_0783__v_fanout (
		.a(n_0783_),
		.b(new_net_1444),
		.c(new_net_6392)
	);

	bfr new_net_6393_bfr_before (
		.din(new_net_6393),
		.dout(new_net_346)
	);

	bfr new_net_6394_bfr_before (
		.din(new_net_6394),
		.dout(new_net_6393)
	);

	spl2 n_1207__v_fanout (
		.a(n_1207_),
		.b(new_net_347),
		.c(new_net_6394)
	);

	spl4L new_net_2063_v_fanout (
		.a(new_net_2063),
		.b(new_net_386),
		.c(new_net_389),
		.d(new_net_2064),
		.e(new_net_380)
	);

	bfr new_net_6395_bfr_before (
		.din(new_net_6395),
		.dout(new_net_1142)
	);

	bfr new_net_6396_bfr_before (
		.din(new_net_6396),
		.dout(new_net_6395)
	);

	spl2 n_1214__v_fanout (
		.a(n_1214_),
		.b(new_net_1143),
		.c(new_net_6396)
	);

	spl4L new_net_2060_v_fanout (
		.a(new_net_2060),
		.b(new_net_383),
		.c(new_net_388),
		.d(new_net_381),
		.e(new_net_379)
	);

	bfr new_net_6397_bfr_before (
		.din(new_net_6397),
		.dout(new_net_1191)
	);

	bfr new_net_6398_bfr_before (
		.din(new_net_6398),
		.dout(new_net_6397)
	);

	spl2 n_0773__v_fanout (
		.a(n_0773_),
		.b(new_net_1192),
		.c(new_net_6398)
	);

	spl4L new_net_2062_v_fanout (
		.a(new_net_2062),
		.b(new_net_378),
		.c(new_net_384),
		.d(new_net_376),
		.e(new_net_372)
	);

	spl3L new_net_2058_v_fanout (
		.a(new_net_2058),
		.b(new_net_375),
		.c(new_net_371),
		.d(new_net_377)
	);

	spl2 n_0736__v_fanout (
		.a(n_0736_),
		.b(new_net_722),
		.c(new_net_721)
	);

	spl2 n_0688__v_fanout (
		.a(n_0688_),
		.b(new_net_846),
		.c(new_net_845)
	);

	bfr new_net_6399_bfr_before (
		.din(new_net_6399),
		.dout(new_net_684)
	);

	bfr new_net_6400_bfr_before (
		.din(new_net_6400),
		.dout(new_net_6399)
	);

	spl2 n_1125__v_fanout (
		.a(n_1125_),
		.b(new_net_685),
		.c(new_net_6400)
	);

	spl2 n_0950__v_fanout (
		.a(n_0950_),
		.b(new_net_1429),
		.c(new_net_1428)
	);

	bfr new_net_6401_bfr_before (
		.din(new_net_6401),
		.dout(new_net_1921)
	);

	bfr new_net_6402_bfr_before (
		.din(new_net_6402),
		.dout(new_net_6401)
	);

	spl2 n_0721__v_fanout (
		.a(n_0721_),
		.b(new_net_1922),
		.c(new_net_6402)
	);

	spl2 n_0886__v_fanout (
		.a(n_0886_),
		.b(new_net_973),
		.c(new_net_972)
	);

	bfr new_net_6403_bfr_before (
		.din(new_net_6403),
		.dout(new_net_518)
	);

	bfr new_net_6404_bfr_before (
		.din(new_net_6404),
		.dout(new_net_6403)
	);

	spl2 n_0719__v_fanout (
		.a(n_0719_),
		.b(new_net_6404),
		.c(new_net_517)
	);

	bfr new_net_6405_bfr_before (
		.din(new_net_6405),
		.dout(new_net_660)
	);

	bfr new_net_6406_bfr_before (
		.din(new_net_6406),
		.dout(new_net_6405)
	);

	spl2 n_1123__v_fanout (
		.a(n_1123_),
		.b(new_net_6406),
		.c(new_net_659)
	);

	spl2 n_0811__v_fanout (
		.a(n_0811_),
		.b(new_net_1159),
		.c(new_net_1158)
	);

	bfr new_net_6407_bfr_before (
		.din(new_net_6407),
		.dout(new_net_857)
	);

	bfr new_net_6408_bfr_before (
		.din(new_net_6408),
		.dout(new_net_6407)
	);

	spl2 n_1133__v_fanout (
		.a(n_1133_),
		.b(new_net_6408),
		.c(new_net_856)
	);

	spl2 n_0672__v_fanout (
		.a(n_0672_),
		.b(new_net_1752),
		.c(new_net_1751)
	);

	bfr new_net_6409_bfr_before (
		.din(new_net_6409),
		.dout(new_net_48)
	);

	bfr new_net_6410_bfr_before (
		.din(new_net_6410),
		.dout(new_net_6409)
	);

	spl2 n_0726__v_fanout (
		.a(n_0726_),
		.b(new_net_6410),
		.c(new_net_47)
	);

	spl2 n_0803__v_fanout (
		.a(n_0803_),
		.b(new_net_1844),
		.c(new_net_1843)
	);

	bfr new_net_6411_bfr_before (
		.din(new_net_6411),
		.dout(new_net_937)
	);

	bfr new_net_6412_bfr_before (
		.din(new_net_6412),
		.dout(new_net_6411)
	);

	spl2 n_1212__v_fanout (
		.a(n_1212_),
		.b(new_net_6412),
		.c(new_net_936)
	);

	bfr new_net_6413_bfr_before (
		.din(new_net_6413),
		.dout(new_net_515)
	);

	bfr new_net_6414_bfr_before (
		.din(new_net_6414),
		.dout(new_net_6413)
	);

	spl2 n_1135__v_fanout (
		.a(n_1135_),
		.b(new_net_516),
		.c(new_net_6414)
	);

	spl2 n_0678__v_fanout (
		.a(n_0678_),
		.b(new_net_1890),
		.c(new_net_1889)
	);

	spl2 n_0823__v_fanout (
		.a(n_0823_),
		.b(new_net_1414),
		.c(new_net_1413)
	);

	bfr new_net_6415_bfr_before (
		.din(new_net_6415),
		.dout(new_net_1406)
	);

	bfr new_net_6416_bfr_before (
		.din(new_net_6416),
		.dout(new_net_6415)
	);

	spl2 n_0781__v_fanout (
		.a(n_0781_),
		.b(new_net_6416),
		.c(new_net_1405)
	);

	spl4L new_net_2061_v_fanout (
		.a(new_net_2061),
		.b(new_net_392),
		.c(new_net_370),
		.d(new_net_374),
		.e(new_net_390)
	);

	spl2 n_0826__v_fanout (
		.a(n_0826_),
		.b(new_net_711),
		.c(new_net_710)
	);

	spl2 new_net_2020_v_fanout (
		.a(new_net_2020),
		.b(new_net_121),
		.c(new_net_159)
	);

	spl2 n_0871__v_fanout (
		.a(n_0871_),
		.b(new_net_68),
		.c(new_net_67)
	);

	spl2 n_0682__v_fanout (
		.a(n_0682_),
		.b(new_net_1105),
		.c(new_net_1104)
	);

	spl2 n_0868__v_fanout (
		.a(n_0868_),
		.b(new_net_1727),
		.c(new_net_1726)
	);

	bfr new_net_6417_bfr_before (
		.din(new_net_6417),
		.dout(new_net_1012)
	);

	bfr new_net_6418_bfr_before (
		.din(new_net_6418),
		.dout(new_net_6417)
	);

	spl2 n_0771__v_fanout (
		.a(n_0771_),
		.b(new_net_6418),
		.c(new_net_1011)
	);

	bfr new_net_6419_bfr_after (
		.din(n_0180_),
		.dout(new_net_6419)
	);

	bfr new_net_6420_bfr_after (
		.din(new_net_6419),
		.dout(new_net_6420)
	);

	bfr new_net_6421_bfr_after (
		.din(new_net_6420),
		.dout(new_net_6421)
	);

	bfr new_net_6422_bfr_after (
		.din(new_net_6421),
		.dout(new_net_6422)
	);

	bfr new_net_6423_bfr_after (
		.din(new_net_6422),
		.dout(new_net_6423)
	);

	bfr new_net_6424_bfr_after (
		.din(new_net_6423),
		.dout(new_net_6424)
	);

	bfr new_net_6425_bfr_after (
		.din(new_net_6424),
		.dout(new_net_6425)
	);

	bfr new_net_6426_bfr_after (
		.din(new_net_6425),
		.dout(new_net_6426)
	);

	bfr new_net_6427_bfr_after (
		.din(new_net_6426),
		.dout(new_net_6427)
	);

	bfr new_net_6428_bfr_after (
		.din(new_net_6427),
		.dout(new_net_6428)
	);

	bfr new_net_6429_bfr_after (
		.din(new_net_6428),
		.dout(new_net_6429)
	);

	bfr new_net_6430_bfr_after (
		.din(new_net_6429),
		.dout(new_net_6430)
	);

	bfr new_net_6431_bfr_after (
		.din(new_net_6430),
		.dout(new_net_6431)
	);

	bfr new_net_6432_bfr_after (
		.din(new_net_6431),
		.dout(new_net_6432)
	);

	bfr new_net_6433_bfr_after (
		.din(new_net_6432),
		.dout(new_net_6433)
	);

	bfr new_net_6434_bfr_after (
		.din(new_net_6433),
		.dout(new_net_6434)
	);

	bfr new_net_6435_bfr_after (
		.din(new_net_6434),
		.dout(new_net_6435)
	);

	bfr new_net_6436_bfr_after (
		.din(new_net_6435),
		.dout(new_net_6436)
	);

	bfr new_net_6437_bfr_after (
		.din(new_net_6436),
		.dout(new_net_6437)
	);

	bfr new_net_6438_bfr_after (
		.din(new_net_6437),
		.dout(new_net_6438)
	);

	bfr new_net_6439_bfr_after (
		.din(new_net_6438),
		.dout(new_net_6439)
	);

	bfr new_net_6440_bfr_after (
		.din(new_net_6439),
		.dout(new_net_6440)
	);

	bfr new_net_6441_bfr_after (
		.din(new_net_6440),
		.dout(new_net_6441)
	);

	bfr new_net_6442_bfr_after (
		.din(new_net_6441),
		.dout(new_net_6442)
	);

	bfr new_net_6443_bfr_after (
		.din(new_net_6442),
		.dout(new_net_6443)
	);

	spl2 n_0180__v_fanout (
		.a(new_net_6443),
		.b(new_net_1135),
		.c(new_net_1134)
	);

	bfr new_net_6444_bfr_before (
		.din(new_net_6444),
		.dout(N945)
	);

	bfr new_net_6445_bfr_before (
		.din(new_net_6445),
		.dout(new_net_6444)
	);

	bfr new_net_6446_bfr_before (
		.din(new_net_6446),
		.dout(new_net_6445)
	);

	bfr new_net_6447_bfr_before (
		.din(new_net_6447),
		.dout(new_net_6446)
	);

	bfr new_net_6448_bfr_before (
		.din(new_net_6448),
		.dout(new_net_6447)
	);

	bfr new_net_6449_bfr_before (
		.din(new_net_6449),
		.dout(new_net_6448)
	);

	bfr new_net_6450_bfr_before (
		.din(new_net_6450),
		.dout(new_net_6449)
	);

	bfr new_net_6451_bfr_before (
		.din(new_net_6451),
		.dout(new_net_6450)
	);

	bfr new_net_6452_bfr_before (
		.din(new_net_6452),
		.dout(new_net_6451)
	);

	bfr new_net_6453_bfr_before (
		.din(new_net_6453),
		.dout(new_net_6452)
	);

	bfr new_net_6454_bfr_before (
		.din(new_net_6454),
		.dout(new_net_6453)
	);

	bfr new_net_6455_bfr_before (
		.din(new_net_6455),
		.dout(new_net_6454)
	);

	bfr new_net_6456_bfr_before (
		.din(new_net_6456),
		.dout(new_net_6455)
	);

	bfr new_net_6457_bfr_before (
		.din(new_net_6457),
		.dout(new_net_6456)
	);

	bfr new_net_6458_bfr_before (
		.din(new_net_6458),
		.dout(new_net_6457)
	);

	bfr new_net_6459_bfr_before (
		.din(new_net_6459),
		.dout(new_net_6458)
	);

	bfr new_net_6460_bfr_before (
		.din(new_net_6460),
		.dout(new_net_6459)
	);

	bfr new_net_6461_bfr_before (
		.din(new_net_6461),
		.dout(new_net_6460)
	);

	bfr new_net_6462_bfr_before (
		.din(new_net_6462),
		.dout(new_net_6461)
	);

	bfr new_net_6463_bfr_before (
		.din(new_net_6463),
		.dout(new_net_6462)
	);

	bfr new_net_6464_bfr_before (
		.din(new_net_6464),
		.dout(new_net_6463)
	);

	bfr new_net_6465_bfr_before (
		.din(new_net_6465),
		.dout(new_net_6464)
	);

	bfr new_net_6466_bfr_before (
		.din(new_net_6466),
		.dout(new_net_6465)
	);

	bfr new_net_6467_bfr_before (
		.din(new_net_6467),
		.dout(new_net_6466)
	);

	bfr new_net_6468_bfr_before (
		.din(new_net_6468),
		.dout(new_net_6467)
	);

	bfr new_net_6469_bfr_before (
		.din(new_net_6469),
		.dout(new_net_6468)
	);

	bfr new_net_6470_bfr_before (
		.din(new_net_6470),
		.dout(new_net_6469)
	);

	bfr new_net_6471_bfr_before (
		.din(new_net_6471),
		.dout(new_net_6470)
	);

	bfr new_net_6472_bfr_before (
		.din(new_net_6472),
		.dout(new_net_6471)
	);

	bfr new_net_6473_bfr_before (
		.din(new_net_6473),
		.dout(new_net_6472)
	);

	bfr new_net_6474_bfr_before (
		.din(new_net_6474),
		.dout(new_net_6473)
	);

	bfr new_net_6475_bfr_before (
		.din(new_net_6475),
		.dout(new_net_6474)
	);

	bfr new_net_6476_bfr_before (
		.din(new_net_6476),
		.dout(new_net_6475)
	);

	bfr new_net_6477_bfr_before (
		.din(new_net_6477),
		.dout(new_net_6476)
	);

	bfr new_net_6478_bfr_before (
		.din(new_net_6478),
		.dout(new_net_6477)
	);

	bfr new_net_6479_bfr_before (
		.din(new_net_6479),
		.dout(new_net_6478)
	);

	bfr new_net_6480_bfr_before (
		.din(new_net_6480),
		.dout(new_net_6479)
	);

	bfr new_net_6481_bfr_before (
		.din(new_net_6481),
		.dout(new_net_6480)
	);

	bfr new_net_6482_bfr_before (
		.din(new_net_6482),
		.dout(new_net_6481)
	);

	bfr new_net_6483_bfr_before (
		.din(new_net_6483),
		.dout(new_net_6482)
	);

	bfr new_net_6484_bfr_before (
		.din(new_net_6484),
		.dout(new_net_6483)
	);

	bfr new_net_6485_bfr_before (
		.din(new_net_6485),
		.dout(new_net_6484)
	);

	bfr new_net_6486_bfr_before (
		.din(new_net_6486),
		.dout(new_net_6485)
	);

	bfr new_net_6487_bfr_before (
		.din(new_net_6487),
		.dout(new_net_6486)
	);

	bfr new_net_6488_bfr_before (
		.din(new_net_6488),
		.dout(new_net_6487)
	);

	bfr new_net_6489_bfr_before (
		.din(new_net_6489),
		.dout(new_net_6488)
	);

	bfr new_net_6490_bfr_before (
		.din(new_net_6490),
		.dout(new_net_6489)
	);

	bfr new_net_6491_bfr_before (
		.din(new_net_6491),
		.dout(new_net_6490)
	);

	bfr new_net_6492_bfr_before (
		.din(new_net_6492),
		.dout(new_net_6491)
	);

	bfr new_net_6493_bfr_before (
		.din(new_net_6493),
		.dout(new_net_6492)
	);

	bfr new_net_6494_bfr_before (
		.din(new_net_6494),
		.dout(new_net_6493)
	);

	bfr new_net_6495_bfr_before (
		.din(new_net_6495),
		.dout(new_net_6494)
	);

	bfr new_net_6496_bfr_before (
		.din(new_net_6496),
		.dout(new_net_6495)
	);

	bfr new_net_6497_bfr_before (
		.din(new_net_6497),
		.dout(new_net_6496)
	);

	bfr new_net_6498_bfr_before (
		.din(new_net_6498),
		.dout(new_net_6497)
	);

	bfr new_net_6499_bfr_before (
		.din(new_net_6499),
		.dout(new_net_6498)
	);

	bfr new_net_6500_bfr_before (
		.din(new_net_6500),
		.dout(new_net_6499)
	);

	bfr new_net_6501_bfr_before (
		.din(new_net_6501),
		.dout(new_net_6500)
	);

	spl3L new_net_1962_v_fanout (
		.a(new_net_1962),
		.b(new_net_1725),
		.c(new_net_1724),
		.d(new_net_6501)
	);

	bfr new_net_6502_bfr_after (
		.din(n_0163_),
		.dout(new_net_6502)
	);

	bfr new_net_6503_bfr_after (
		.din(new_net_6502),
		.dout(new_net_6503)
	);

	bfr new_net_6504_bfr_after (
		.din(new_net_6503),
		.dout(new_net_6504)
	);

	bfr new_net_6505_bfr_after (
		.din(new_net_6504),
		.dout(new_net_6505)
	);

	bfr new_net_6506_bfr_after (
		.din(new_net_6505),
		.dout(new_net_6506)
	);

	bfr new_net_6507_bfr_after (
		.din(new_net_6506),
		.dout(new_net_6507)
	);

	bfr new_net_6508_bfr_after (
		.din(new_net_6507),
		.dout(new_net_6508)
	);

	bfr new_net_6509_bfr_after (
		.din(new_net_6508),
		.dout(new_net_6509)
	);

	bfr new_net_6510_bfr_after (
		.din(new_net_6509),
		.dout(new_net_6510)
	);

	bfr new_net_6511_bfr_after (
		.din(new_net_6510),
		.dout(new_net_6511)
	);

	bfr new_net_6512_bfr_after (
		.din(new_net_6511),
		.dout(new_net_6512)
	);

	bfr new_net_6513_bfr_after (
		.din(new_net_6512),
		.dout(new_net_6513)
	);

	bfr new_net_6514_bfr_after (
		.din(new_net_6513),
		.dout(new_net_6514)
	);

	bfr new_net_6515_bfr_after (
		.din(new_net_6514),
		.dout(new_net_6515)
	);

	bfr new_net_6516_bfr_after (
		.din(new_net_6515),
		.dout(new_net_6516)
	);

	bfr new_net_6517_bfr_after (
		.din(new_net_6516),
		.dout(new_net_6517)
	);

	bfr new_net_6518_bfr_after (
		.din(new_net_6517),
		.dout(new_net_6518)
	);

	bfr new_net_6519_bfr_after (
		.din(new_net_6518),
		.dout(new_net_6519)
	);

	bfr new_net_6520_bfr_after (
		.din(new_net_6519),
		.dout(new_net_6520)
	);

	bfr new_net_6521_bfr_after (
		.din(new_net_6520),
		.dout(new_net_6521)
	);

	bfr new_net_6522_bfr_after (
		.din(new_net_6521),
		.dout(new_net_6522)
	);

	bfr new_net_6523_bfr_after (
		.din(new_net_6522),
		.dout(new_net_6523)
	);

	bfr new_net_6524_bfr_after (
		.din(new_net_6523),
		.dout(new_net_6524)
	);

	bfr new_net_6525_bfr_after (
		.din(new_net_6524),
		.dout(new_net_6525)
	);

	bfr new_net_6526_bfr_after (
		.din(new_net_6525),
		.dout(new_net_6526)
	);

	bfr new_net_6527_bfr_after (
		.din(new_net_6526),
		.dout(new_net_6527)
	);

	bfr new_net_6528_bfr_after (
		.din(new_net_6527),
		.dout(new_net_6528)
	);

	bfr new_net_6529_bfr_after (
		.din(new_net_6528),
		.dout(new_net_6529)
	);

	bfr new_net_6530_bfr_after (
		.din(new_net_6529),
		.dout(new_net_6530)
	);

	bfr new_net_6531_bfr_after (
		.din(new_net_6530),
		.dout(new_net_6531)
	);

	bfr new_net_6532_bfr_after (
		.din(new_net_6531),
		.dout(new_net_6532)
	);

	bfr new_net_6533_bfr_after (
		.din(new_net_6532),
		.dout(new_net_6533)
	);

	bfr new_net_6534_bfr_after (
		.din(new_net_6533),
		.dout(new_net_6534)
	);

	bfr new_net_6535_bfr_after (
		.din(new_net_6534),
		.dout(new_net_6535)
	);

	bfr new_net_6536_bfr_after (
		.din(new_net_6535),
		.dout(new_net_6536)
	);

	bfr new_net_6537_bfr_after (
		.din(new_net_6536),
		.dout(new_net_6537)
	);

	bfr new_net_6538_bfr_after (
		.din(new_net_6537),
		.dout(new_net_6538)
	);

	bfr new_net_6539_bfr_after (
		.din(new_net_6538),
		.dout(new_net_6539)
	);

	bfr new_net_6540_bfr_after (
		.din(new_net_6539),
		.dout(new_net_6540)
	);

	bfr new_net_6541_bfr_after (
		.din(new_net_6540),
		.dout(new_net_6541)
	);

	bfr new_net_6542_bfr_after (
		.din(new_net_6541),
		.dout(new_net_6542)
	);

	bfr new_net_6543_bfr_after (
		.din(new_net_6542),
		.dout(new_net_6543)
	);

	bfr new_net_6544_bfr_after (
		.din(new_net_6543),
		.dout(new_net_6544)
	);

	bfr new_net_6545_bfr_after (
		.din(new_net_6544),
		.dout(new_net_6545)
	);

	bfr new_net_6546_bfr_after (
		.din(new_net_6545),
		.dout(new_net_6546)
	);

	bfr new_net_6547_bfr_after (
		.din(new_net_6546),
		.dout(new_net_6547)
	);

	bfr new_net_6548_bfr_after (
		.din(new_net_6547),
		.dout(new_net_6548)
	);

	bfr new_net_6549_bfr_after (
		.din(new_net_6548),
		.dout(new_net_6549)
	);

	bfr new_net_6550_bfr_after (
		.din(new_net_6549),
		.dout(new_net_6550)
	);

	bfr new_net_6551_bfr_after (
		.din(new_net_6550),
		.dout(new_net_6551)
	);

	bfr new_net_6552_bfr_after (
		.din(new_net_6551),
		.dout(new_net_6552)
	);

	bfr new_net_6553_bfr_after (
		.din(new_net_6552),
		.dout(new_net_6553)
	);

	bfr new_net_6554_bfr_after (
		.din(new_net_6553),
		.dout(new_net_6554)
	);

	bfr new_net_6555_bfr_after (
		.din(new_net_6554),
		.dout(new_net_6555)
	);

	bfr new_net_6556_bfr_after (
		.din(new_net_6555),
		.dout(new_net_6556)
	);

	bfr new_net_6557_bfr_after (
		.din(new_net_6556),
		.dout(new_net_6557)
	);

	bfr new_net_6558_bfr_after (
		.din(new_net_6557),
		.dout(new_net_6558)
	);

	bfr new_net_6559_bfr_after (
		.din(new_net_6558),
		.dout(new_net_6559)
	);

	bfr new_net_6560_bfr_after (
		.din(new_net_6559),
		.dout(new_net_6560)
	);

	spl4L n_0163__v_fanout (
		.a(new_net_6560),
		.b(new_net_454),
		.c(new_net_455),
		.d(new_net_453),
		.e(new_net_452)
	);

	spl2 new_net_2035_v_fanout (
		.a(new_net_2035),
		.b(new_net_2036),
		.c(new_net_512)
	);

	spl4L new_net_2057_v_fanout (
		.a(new_net_2057),
		.b(new_net_391),
		.c(new_net_387),
		.d(new_net_2058),
		.e(new_net_385)
	);

	spl4L new_net_2059_v_fanout (
		.a(new_net_2059),
		.b(new_net_2062),
		.c(new_net_2061),
		.d(new_net_2063),
		.e(new_net_2060)
	);

	bfr new_net_6561_bfr_before (
		.din(new_net_6561),
		.dout(new_net_2067)
	);

	bfr new_net_6562_bfr_before (
		.din(new_net_6562),
		.dout(new_net_6561)
	);

	bfr new_net_6563_bfr_before (
		.din(new_net_6563),
		.dout(new_net_6562)
	);

	bfr new_net_6564_bfr_before (
		.din(new_net_6564),
		.dout(new_net_6563)
	);

	bfr new_net_6565_bfr_before (
		.din(new_net_6565),
		.dout(new_net_6564)
	);

	bfr new_net_6566_bfr_before (
		.din(new_net_6566),
		.dout(new_net_6565)
	);

	bfr new_net_6567_bfr_before (
		.din(new_net_6567),
		.dout(new_net_6566)
	);

	bfr new_net_6568_bfr_before (
		.din(new_net_6568),
		.dout(new_net_6567)
	);

	bfr new_net_6569_bfr_before (
		.din(new_net_6569),
		.dout(new_net_6568)
	);

	bfr new_net_6570_bfr_before (
		.din(new_net_6570),
		.dout(new_net_6569)
	);

	bfr new_net_6571_bfr_before (
		.din(new_net_6571),
		.dout(new_net_6570)
	);

	bfr new_net_6572_bfr_before (
		.din(new_net_6572),
		.dout(new_net_6571)
	);

	bfr new_net_6573_bfr_before (
		.din(new_net_6573),
		.dout(new_net_6572)
	);

	bfr new_net_6574_bfr_before (
		.din(new_net_6574),
		.dout(new_net_6573)
	);

	bfr new_net_6575_bfr_before (
		.din(new_net_6575),
		.dout(new_net_6574)
	);

	bfr new_net_6576_bfr_before (
		.din(new_net_6576),
		.dout(new_net_6575)
	);

	bfr new_net_6577_bfr_before (
		.din(new_net_6577),
		.dout(new_net_6576)
	);

	bfr new_net_6578_bfr_before (
		.din(new_net_6578),
		.dout(new_net_6577)
	);

	bfr new_net_6579_bfr_before (
		.din(new_net_6579),
		.dout(new_net_6578)
	);

	bfr new_net_6580_bfr_before (
		.din(new_net_6580),
		.dout(new_net_6579)
	);

	bfr new_net_6581_bfr_before (
		.din(new_net_6581),
		.dout(new_net_6580)
	);

	bfr new_net_6582_bfr_before (
		.din(new_net_6582),
		.dout(new_net_6581)
	);

	bfr new_net_6583_bfr_before (
		.din(new_net_6583),
		.dout(new_net_6582)
	);

	bfr new_net_6584_bfr_before (
		.din(new_net_6584),
		.dout(new_net_6583)
	);

	bfr new_net_6585_bfr_before (
		.din(new_net_6585),
		.dout(new_net_6584)
	);

	bfr new_net_6586_bfr_before (
		.din(new_net_6586),
		.dout(new_net_6585)
	);

	bfr new_net_6587_bfr_before (
		.din(new_net_6587),
		.dout(new_net_6586)
	);

	bfr new_net_6588_bfr_before (
		.din(new_net_6588),
		.dout(new_net_6587)
	);

	bfr new_net_6589_bfr_before (
		.din(new_net_6589),
		.dout(new_net_6588)
	);

	bfr new_net_6590_bfr_before (
		.din(new_net_6590),
		.dout(new_net_6589)
	);

	bfr new_net_6591_bfr_before (
		.din(new_net_6591),
		.dout(new_net_6590)
	);

	bfr new_net_6592_bfr_before (
		.din(new_net_6592),
		.dout(new_net_6591)
	);

	bfr new_net_6593_bfr_before (
		.din(new_net_6593),
		.dout(new_net_6592)
	);

	bfr new_net_6594_bfr_before (
		.din(new_net_6594),
		.dout(new_net_6593)
	);

	bfr new_net_6595_bfr_before (
		.din(new_net_6595),
		.dout(new_net_6594)
	);

	bfr new_net_6596_bfr_before (
		.din(new_net_6596),
		.dout(new_net_6595)
	);

	bfr new_net_6597_bfr_before (
		.din(new_net_6597),
		.dout(new_net_6596)
	);

	bfr new_net_6598_bfr_before (
		.din(new_net_6598),
		.dout(new_net_6597)
	);

	bfr new_net_6599_bfr_before (
		.din(new_net_6599),
		.dout(new_net_6598)
	);

	bfr new_net_6600_bfr_before (
		.din(new_net_6600),
		.dout(new_net_6599)
	);

	bfr new_net_6601_bfr_before (
		.din(new_net_6601),
		.dout(new_net_6600)
	);

	bfr new_net_6602_bfr_before (
		.din(new_net_6602),
		.dout(new_net_6601)
	);

	bfr new_net_6603_bfr_before (
		.din(new_net_6603),
		.dout(new_net_6602)
	);

	bfr new_net_6604_bfr_before (
		.din(new_net_6604),
		.dout(new_net_6603)
	);

	bfr new_net_6605_bfr_before (
		.din(new_net_6605),
		.dout(new_net_6604)
	);

	bfr new_net_6606_bfr_before (
		.din(new_net_6606),
		.dout(new_net_6605)
	);

	bfr new_net_6607_bfr_before (
		.din(new_net_6607),
		.dout(new_net_6606)
	);

	bfr new_net_6608_bfr_before (
		.din(new_net_6608),
		.dout(new_net_6607)
	);

	bfr new_net_6609_bfr_before (
		.din(new_net_6609),
		.dout(new_net_6608)
	);

	bfr new_net_6610_bfr_before (
		.din(new_net_6610),
		.dout(new_net_6609)
	);

	bfr new_net_6611_bfr_before (
		.din(new_net_6611),
		.dout(new_net_6610)
	);

	bfr new_net_6612_bfr_before (
		.din(new_net_6612),
		.dout(new_net_6611)
	);

	bfr new_net_6613_bfr_before (
		.din(new_net_6613),
		.dout(new_net_6612)
	);

	bfr new_net_6614_bfr_before (
		.din(new_net_6614),
		.dout(new_net_6613)
	);

	spl2 n_0167__v_fanout (
		.a(n_0167_),
		.b(new_net_6614),
		.c(new_net_893)
	);

	spl2 new_net_2019_v_fanout (
		.a(new_net_2019),
		.b(new_net_2020),
		.c(new_net_151)
	);

	bfr new_net_6615_bfr_after (
		.din(n_0379_),
		.dout(new_net_6615)
	);

	bfr new_net_6616_bfr_after (
		.din(new_net_6615),
		.dout(new_net_6616)
	);

	bfr new_net_6617_bfr_after (
		.din(new_net_6616),
		.dout(new_net_6617)
	);

	bfr new_net_6618_bfr_after (
		.din(new_net_6617),
		.dout(new_net_6618)
	);

	bfr new_net_6619_bfr_after (
		.din(new_net_6618),
		.dout(new_net_6619)
	);

	bfr new_net_6620_bfr_after (
		.din(new_net_6619),
		.dout(new_net_6620)
	);

	bfr new_net_6621_bfr_after (
		.din(new_net_6620),
		.dout(new_net_6621)
	);

	bfr new_net_6622_bfr_after (
		.din(new_net_6621),
		.dout(new_net_6622)
	);

	bfr new_net_6623_bfr_after (
		.din(new_net_6622),
		.dout(new_net_6623)
	);

	bfr new_net_6624_bfr_after (
		.din(new_net_6623),
		.dout(new_net_6624)
	);

	bfr new_net_6625_bfr_before (
		.din(new_net_6625),
		.dout(new_net_876)
	);

	bfr new_net_6626_bfr_before (
		.din(new_net_6626),
		.dout(new_net_6625)
	);

	bfr new_net_6627_bfr_before (
		.din(new_net_6627),
		.dout(new_net_6626)
	);

	bfr new_net_6628_bfr_before (
		.din(new_net_6628),
		.dout(new_net_6627)
	);

	bfr new_net_6629_bfr_before (
		.din(new_net_6629),
		.dout(new_net_6628)
	);

	bfr new_net_6630_bfr_before (
		.din(new_net_6630),
		.dout(new_net_6629)
	);

	bfr new_net_6631_bfr_before (
		.din(new_net_6631),
		.dout(new_net_6630)
	);

	bfr new_net_6632_bfr_before (
		.din(new_net_6632),
		.dout(new_net_6631)
	);

	bfr new_net_6633_bfr_before (
		.din(new_net_6633),
		.dout(new_net_6632)
	);

	bfr new_net_6634_bfr_before (
		.din(new_net_6634),
		.dout(new_net_6633)
	);

	bfr new_net_6635_bfr_before (
		.din(new_net_6635),
		.dout(new_net_6634)
	);

	bfr new_net_6636_bfr_before (
		.din(new_net_6636),
		.dout(new_net_6635)
	);

	bfr new_net_6637_bfr_before (
		.din(new_net_6637),
		.dout(new_net_6636)
	);

	bfr new_net_6638_bfr_before (
		.din(new_net_6638),
		.dout(new_net_6637)
	);

	bfr new_net_6639_bfr_before (
		.din(new_net_6639),
		.dout(new_net_6638)
	);

	bfr new_net_6640_bfr_before (
		.din(new_net_6640),
		.dout(new_net_6639)
	);

	bfr new_net_6641_bfr_before (
		.din(new_net_6641),
		.dout(new_net_6640)
	);

	bfr new_net_6642_bfr_before (
		.din(new_net_6642),
		.dout(new_net_6641)
	);

	bfr new_net_6643_bfr_before (
		.din(new_net_6643),
		.dout(new_net_6642)
	);

	bfr new_net_6644_bfr_before (
		.din(new_net_6644),
		.dout(new_net_6643)
	);

	bfr new_net_6645_bfr_before (
		.din(new_net_6645),
		.dout(new_net_6644)
	);

	bfr new_net_6646_bfr_before (
		.din(new_net_6646),
		.dout(new_net_6645)
	);

	bfr new_net_6647_bfr_before (
		.din(new_net_6647),
		.dout(new_net_6646)
	);

	bfr new_net_6648_bfr_before (
		.din(new_net_6648),
		.dout(new_net_6647)
	);

	bfr new_net_6649_bfr_before (
		.din(new_net_6649),
		.dout(new_net_6648)
	);

	bfr new_net_6650_bfr_before (
		.din(new_net_6650),
		.dout(new_net_6649)
	);

	bfr new_net_6651_bfr_before (
		.din(new_net_6651),
		.dout(new_net_6650)
	);

	bfr new_net_6652_bfr_before (
		.din(new_net_6652),
		.dout(new_net_6651)
	);

	bfr new_net_6653_bfr_before (
		.din(new_net_6653),
		.dout(new_net_6652)
	);

	bfr new_net_6654_bfr_before (
		.din(new_net_6654),
		.dout(new_net_6653)
	);

	bfr new_net_6655_bfr_before (
		.din(new_net_6655),
		.dout(new_net_6654)
	);

	bfr new_net_6656_bfr_before (
		.din(new_net_6656),
		.dout(new_net_6655)
	);

	bfr new_net_6657_bfr_before (
		.din(new_net_6657),
		.dout(new_net_6656)
	);

	bfr new_net_6658_bfr_before (
		.din(new_net_6658),
		.dout(new_net_6657)
	);

	bfr new_net_6659_bfr_before (
		.din(new_net_6659),
		.dout(new_net_6658)
	);

	bfr new_net_6660_bfr_before (
		.din(new_net_6660),
		.dout(new_net_6659)
	);

	bfr new_net_6661_bfr_before (
		.din(new_net_6661),
		.dout(new_net_6660)
	);

	bfr new_net_6662_bfr_before (
		.din(new_net_6662),
		.dout(new_net_6661)
	);

	bfr new_net_6663_bfr_before (
		.din(new_net_6663),
		.dout(new_net_6662)
	);

	bfr new_net_6664_bfr_before (
		.din(new_net_6664),
		.dout(new_net_6663)
	);

	bfr new_net_6665_bfr_before (
		.din(new_net_6665),
		.dout(new_net_6664)
	);

	bfr new_net_6666_bfr_before (
		.din(new_net_6666),
		.dout(new_net_6665)
	);

	bfr new_net_6667_bfr_before (
		.din(new_net_6667),
		.dout(new_net_6666)
	);

	bfr new_net_6668_bfr_before (
		.din(new_net_6668),
		.dout(new_net_6667)
	);

	bfr new_net_6669_bfr_before (
		.din(new_net_6669),
		.dout(new_net_6668)
	);

	bfr new_net_6670_bfr_before (
		.din(new_net_6670),
		.dout(new_net_6669)
	);

	bfr new_net_6671_bfr_before (
		.din(new_net_6671),
		.dout(new_net_6670)
	);

	bfr new_net_6672_bfr_before (
		.din(new_net_6672),
		.dout(new_net_6671)
	);

	spl3L n_0379__v_fanout (
		.a(new_net_6624),
		.b(new_net_877),
		.c(new_net_6672),
		.d(new_net_878)
	);

	bfr new_net_6673_bfr_before (
		.din(new_net_6673),
		.dout(new_net_2068)
	);

	bfr new_net_6674_bfr_before (
		.din(new_net_6674),
		.dout(new_net_6673)
	);

	bfr new_net_6675_bfr_before (
		.din(new_net_6675),
		.dout(new_net_6674)
	);

	bfr new_net_6676_bfr_before (
		.din(new_net_6676),
		.dout(new_net_6675)
	);

	bfr new_net_6677_bfr_before (
		.din(new_net_6677),
		.dout(new_net_6676)
	);

	bfr new_net_6678_bfr_before (
		.din(new_net_6678),
		.dout(new_net_6677)
	);

	bfr new_net_6679_bfr_before (
		.din(new_net_6679),
		.dout(new_net_6678)
	);

	bfr new_net_6680_bfr_before (
		.din(new_net_6680),
		.dout(new_net_6679)
	);

	bfr new_net_6681_bfr_before (
		.din(new_net_6681),
		.dout(new_net_6680)
	);

	bfr new_net_6682_bfr_before (
		.din(new_net_6682),
		.dout(new_net_6681)
	);

	bfr new_net_6683_bfr_before (
		.din(new_net_6683),
		.dout(new_net_6682)
	);

	bfr new_net_6684_bfr_before (
		.din(new_net_6684),
		.dout(new_net_6683)
	);

	bfr new_net_6685_bfr_before (
		.din(new_net_6685),
		.dout(new_net_6684)
	);

	bfr new_net_6686_bfr_before (
		.din(new_net_6686),
		.dout(new_net_6685)
	);

	bfr new_net_6687_bfr_before (
		.din(new_net_6687),
		.dout(new_net_6686)
	);

	bfr new_net_6688_bfr_before (
		.din(new_net_6688),
		.dout(new_net_6687)
	);

	bfr new_net_6689_bfr_before (
		.din(new_net_6689),
		.dout(new_net_6688)
	);

	bfr new_net_6690_bfr_before (
		.din(new_net_6690),
		.dout(new_net_6689)
	);

	bfr new_net_6691_bfr_before (
		.din(new_net_6691),
		.dout(new_net_6690)
	);

	bfr new_net_6692_bfr_before (
		.din(new_net_6692),
		.dout(new_net_6691)
	);

	bfr new_net_6693_bfr_before (
		.din(new_net_6693),
		.dout(new_net_6692)
	);

	bfr new_net_6694_bfr_before (
		.din(new_net_6694),
		.dout(new_net_6693)
	);

	bfr new_net_6695_bfr_before (
		.din(new_net_6695),
		.dout(new_net_6694)
	);

	bfr new_net_6696_bfr_before (
		.din(new_net_6696),
		.dout(new_net_6695)
	);

	bfr new_net_6697_bfr_before (
		.din(new_net_6697),
		.dout(new_net_6696)
	);

	bfr new_net_6698_bfr_before (
		.din(new_net_6698),
		.dout(new_net_6697)
	);

	bfr new_net_6699_bfr_before (
		.din(new_net_6699),
		.dout(new_net_6698)
	);

	bfr new_net_6700_bfr_before (
		.din(new_net_6700),
		.dout(new_net_6699)
	);

	bfr new_net_6701_bfr_before (
		.din(new_net_6701),
		.dout(new_net_6700)
	);

	bfr new_net_6702_bfr_before (
		.din(new_net_6702),
		.dout(new_net_6701)
	);

	bfr new_net_6703_bfr_before (
		.din(new_net_6703),
		.dout(new_net_6702)
	);

	bfr new_net_6704_bfr_before (
		.din(new_net_6704),
		.dout(new_net_6703)
	);

	bfr new_net_6705_bfr_before (
		.din(new_net_6705),
		.dout(new_net_6704)
	);

	bfr new_net_6706_bfr_before (
		.din(new_net_6706),
		.dout(new_net_6705)
	);

	bfr new_net_6707_bfr_before (
		.din(new_net_6707),
		.dout(new_net_6706)
	);

	bfr new_net_6708_bfr_before (
		.din(new_net_6708),
		.dout(new_net_6707)
	);

	bfr new_net_6709_bfr_before (
		.din(new_net_6709),
		.dout(new_net_6708)
	);

	bfr new_net_6710_bfr_before (
		.din(new_net_6710),
		.dout(new_net_6709)
	);

	bfr new_net_6711_bfr_before (
		.din(new_net_6711),
		.dout(new_net_6710)
	);

	bfr new_net_6712_bfr_before (
		.din(new_net_6712),
		.dout(new_net_6711)
	);

	bfr new_net_6713_bfr_before (
		.din(new_net_6713),
		.dout(new_net_6712)
	);

	bfr new_net_6714_bfr_before (
		.din(new_net_6714),
		.dout(new_net_6713)
	);

	bfr new_net_6715_bfr_before (
		.din(new_net_6715),
		.dout(new_net_6714)
	);

	bfr new_net_6716_bfr_before (
		.din(new_net_6716),
		.dout(new_net_6715)
	);

	bfr new_net_6717_bfr_before (
		.din(new_net_6717),
		.dout(new_net_6716)
	);

	bfr new_net_6718_bfr_before (
		.din(new_net_6718),
		.dout(new_net_6717)
	);

	bfr new_net_6719_bfr_before (
		.din(new_net_6719),
		.dout(new_net_6718)
	);

	bfr new_net_6720_bfr_before (
		.din(new_net_6720),
		.dout(new_net_6719)
	);

	bfr new_net_6721_bfr_before (
		.din(new_net_6721),
		.dout(new_net_6720)
	);

	bfr new_net_6722_bfr_before (
		.din(new_net_6722),
		.dout(new_net_6721)
	);

	bfr new_net_6723_bfr_before (
		.din(new_net_6723),
		.dout(new_net_6722)
	);

	bfr new_net_6724_bfr_before (
		.din(new_net_6724),
		.dout(new_net_6723)
	);

	bfr new_net_6725_bfr_before (
		.din(new_net_6725),
		.dout(new_net_6724)
	);

	bfr new_net_6726_bfr_before (
		.din(new_net_6726),
		.dout(new_net_6725)
	);

	spl2 n_0168__v_fanout (
		.a(n_0168_),
		.b(new_net_6726),
		.c(new_net_1006)
	);

	spl4L new_net_2016_v_fanout (
		.a(new_net_2016),
		.b(new_net_287),
		.c(new_net_245),
		.d(new_net_254),
		.e(new_net_182)
	);

	spl4L new_net_1980_v_fanout (
		.a(new_net_1980),
		.b(new_net_128),
		.c(new_net_211),
		.d(new_net_120),
		.e(new_net_283)
	);

	spl4L new_net_1992_v_fanout (
		.a(new_net_1992),
		.b(new_net_230),
		.c(new_net_199),
		.d(new_net_209),
		.e(new_net_281)
	);

	spl4L new_net_1985_v_fanout (
		.a(new_net_1985),
		.b(new_net_240),
		.c(new_net_282),
		.d(new_net_219),
		.e(new_net_250)
	);

	bfr new_net_6727_bfr_before (
		.din(new_net_6727),
		.dout(N545)
	);

	bfr new_net_6728_bfr_before (
		.din(new_net_6728),
		.dout(new_net_6727)
	);

	bfr new_net_6729_bfr_before (
		.din(new_net_6729),
		.dout(new_net_6728)
	);

	bfr new_net_6730_bfr_before (
		.din(new_net_6730),
		.dout(new_net_6729)
	);

	bfr new_net_6731_bfr_before (
		.din(new_net_6731),
		.dout(new_net_6730)
	);

	bfr new_net_6732_bfr_before (
		.din(new_net_6732),
		.dout(new_net_6731)
	);

	bfr new_net_6733_bfr_before (
		.din(new_net_6733),
		.dout(new_net_6732)
	);

	bfr new_net_6734_bfr_before (
		.din(new_net_6734),
		.dout(new_net_6733)
	);

	bfr new_net_6735_bfr_before (
		.din(new_net_6735),
		.dout(new_net_6734)
	);

	bfr new_net_6736_bfr_before (
		.din(new_net_6736),
		.dout(new_net_6735)
	);

	bfr new_net_6737_bfr_before (
		.din(new_net_6737),
		.dout(new_net_6736)
	);

	bfr new_net_6738_bfr_before (
		.din(new_net_6738),
		.dout(new_net_6737)
	);

	bfr new_net_6739_bfr_before (
		.din(new_net_6739),
		.dout(new_net_6738)
	);

	bfr new_net_6740_bfr_before (
		.din(new_net_6740),
		.dout(new_net_6739)
	);

	bfr new_net_6741_bfr_before (
		.din(new_net_6741),
		.dout(new_net_6740)
	);

	bfr new_net_6742_bfr_before (
		.din(new_net_6742),
		.dout(new_net_6741)
	);

	bfr new_net_6743_bfr_before (
		.din(new_net_6743),
		.dout(new_net_6742)
	);

	bfr new_net_6744_bfr_before (
		.din(new_net_6744),
		.dout(new_net_6743)
	);

	bfr new_net_6745_bfr_before (
		.din(new_net_6745),
		.dout(new_net_6744)
	);

	bfr new_net_6746_bfr_before (
		.din(new_net_6746),
		.dout(new_net_6745)
	);

	bfr new_net_6747_bfr_before (
		.din(new_net_6747),
		.dout(new_net_6746)
	);

	bfr new_net_6748_bfr_before (
		.din(new_net_6748),
		.dout(new_net_6747)
	);

	bfr new_net_6749_bfr_before (
		.din(new_net_6749),
		.dout(new_net_6748)
	);

	bfr new_net_6750_bfr_before (
		.din(new_net_6750),
		.dout(new_net_6749)
	);

	bfr new_net_6751_bfr_before (
		.din(new_net_6751),
		.dout(new_net_6750)
	);

	bfr new_net_6752_bfr_before (
		.din(new_net_6752),
		.dout(new_net_6751)
	);

	bfr new_net_6753_bfr_before (
		.din(new_net_6753),
		.dout(new_net_6752)
	);

	bfr new_net_6754_bfr_before (
		.din(new_net_6754),
		.dout(new_net_6753)
	);

	bfr new_net_6755_bfr_before (
		.din(new_net_6755),
		.dout(new_net_6754)
	);

	bfr new_net_6756_bfr_before (
		.din(new_net_6756),
		.dout(new_net_6755)
	);

	bfr new_net_6757_bfr_before (
		.din(new_net_6757),
		.dout(new_net_6756)
	);

	bfr new_net_6758_bfr_before (
		.din(new_net_6758),
		.dout(new_net_6757)
	);

	bfr new_net_6759_bfr_before (
		.din(new_net_6759),
		.dout(new_net_6758)
	);

	bfr new_net_6760_bfr_before (
		.din(new_net_6760),
		.dout(new_net_6759)
	);

	bfr new_net_6761_bfr_before (
		.din(new_net_6761),
		.dout(new_net_6760)
	);

	bfr new_net_6762_bfr_before (
		.din(new_net_6762),
		.dout(new_net_6761)
	);

	bfr new_net_6763_bfr_before (
		.din(new_net_6763),
		.dout(new_net_6762)
	);

	bfr new_net_6764_bfr_before (
		.din(new_net_6764),
		.dout(new_net_6763)
	);

	bfr new_net_6765_bfr_before (
		.din(new_net_6765),
		.dout(new_net_6764)
	);

	bfr new_net_6766_bfr_before (
		.din(new_net_6766),
		.dout(new_net_6765)
	);

	bfr new_net_6767_bfr_before (
		.din(new_net_6767),
		.dout(new_net_6766)
	);

	bfr new_net_6768_bfr_before (
		.din(new_net_6768),
		.dout(new_net_6767)
	);

	bfr new_net_6769_bfr_before (
		.din(new_net_6769),
		.dout(new_net_6768)
	);

	bfr new_net_6770_bfr_before (
		.din(new_net_6770),
		.dout(new_net_6769)
	);

	bfr new_net_6771_bfr_before (
		.din(new_net_6771),
		.dout(new_net_6770)
	);

	bfr new_net_6772_bfr_before (
		.din(new_net_6772),
		.dout(new_net_6771)
	);

	bfr new_net_6773_bfr_before (
		.din(new_net_6773),
		.dout(new_net_6772)
	);

	bfr new_net_6774_bfr_before (
		.din(new_net_6774),
		.dout(new_net_6773)
	);

	bfr new_net_6775_bfr_before (
		.din(new_net_6775),
		.dout(new_net_6774)
	);

	bfr new_net_6776_bfr_before (
		.din(new_net_6776),
		.dout(new_net_6775)
	);

	bfr new_net_6777_bfr_before (
		.din(new_net_6777),
		.dout(new_net_6776)
	);

	bfr new_net_6778_bfr_before (
		.din(new_net_6778),
		.dout(new_net_6777)
	);

	bfr new_net_6779_bfr_before (
		.din(new_net_6779),
		.dout(new_net_6778)
	);

	bfr new_net_6780_bfr_before (
		.din(new_net_6780),
		.dout(new_net_6779)
	);

	bfr new_net_6781_bfr_before (
		.din(new_net_6781),
		.dout(new_net_6780)
	);

	bfr new_net_6782_bfr_before (
		.din(new_net_6782),
		.dout(new_net_6781)
	);

	bfr new_net_6783_bfr_before (
		.din(new_net_6783),
		.dout(new_net_6782)
	);

	bfr new_net_6784_bfr_before (
		.din(new_net_6784),
		.dout(new_net_6783)
	);

	bfr new_net_6785_bfr_before (
		.din(new_net_6785),
		.dout(new_net_6784)
	);

	bfr new_net_6786_bfr_before (
		.din(new_net_6786),
		.dout(new_net_6785)
	);

	bfr new_net_6787_bfr_before (
		.din(new_net_6787),
		.dout(new_net_6786)
	);

	bfr new_net_6788_bfr_before (
		.din(new_net_6788),
		.dout(new_net_6787)
	);

	spl2 new_net_2040_v_fanout (
		.a(new_net_2040),
		.b(new_net_6788),
		.c(new_net_1080)
	);

	spl4L new_net_2008_v_fanout (
		.a(new_net_2008),
		.b(new_net_195),
		.c(new_net_174),
		.d(new_net_208),
		.e(new_net_153)
	);

	spl4L new_net_1982_v_fanout (
		.a(new_net_1982),
		.b(new_net_157),
		.c(new_net_191),
		.d(new_net_170),
		.e(new_net_149)
	);

	spl4L new_net_1984_v_fanout (
		.a(new_net_1984),
		.b(new_net_223),
		.c(new_net_265),
		.d(new_net_259),
		.e(new_net_202)
	);

	bfr new_net_6789_bfr_before (
		.din(new_net_6789),
		.dout(N561)
	);

	bfr new_net_6790_bfr_before (
		.din(new_net_6790),
		.dout(new_net_6789)
	);

	bfr new_net_6791_bfr_before (
		.din(new_net_6791),
		.dout(new_net_6790)
	);

	bfr new_net_6792_bfr_before (
		.din(new_net_6792),
		.dout(new_net_6791)
	);

	bfr new_net_6793_bfr_before (
		.din(new_net_6793),
		.dout(new_net_6792)
	);

	bfr new_net_6794_bfr_before (
		.din(new_net_6794),
		.dout(new_net_6793)
	);

	bfr new_net_6795_bfr_before (
		.din(new_net_6795),
		.dout(new_net_6794)
	);

	bfr new_net_6796_bfr_before (
		.din(new_net_6796),
		.dout(new_net_6795)
	);

	bfr new_net_6797_bfr_before (
		.din(new_net_6797),
		.dout(new_net_6796)
	);

	bfr new_net_6798_bfr_before (
		.din(new_net_6798),
		.dout(new_net_6797)
	);

	bfr new_net_6799_bfr_before (
		.din(new_net_6799),
		.dout(new_net_6798)
	);

	bfr new_net_6800_bfr_before (
		.din(new_net_6800),
		.dout(new_net_6799)
	);

	bfr new_net_6801_bfr_before (
		.din(new_net_6801),
		.dout(new_net_6800)
	);

	bfr new_net_6802_bfr_before (
		.din(new_net_6802),
		.dout(new_net_6801)
	);

	bfr new_net_6803_bfr_before (
		.din(new_net_6803),
		.dout(new_net_6802)
	);

	bfr new_net_6804_bfr_before (
		.din(new_net_6804),
		.dout(new_net_6803)
	);

	bfr new_net_6805_bfr_before (
		.din(new_net_6805),
		.dout(new_net_6804)
	);

	bfr new_net_6806_bfr_before (
		.din(new_net_6806),
		.dout(new_net_6805)
	);

	bfr new_net_6807_bfr_before (
		.din(new_net_6807),
		.dout(new_net_6806)
	);

	bfr new_net_6808_bfr_before (
		.din(new_net_6808),
		.dout(new_net_6807)
	);

	bfr new_net_6809_bfr_before (
		.din(new_net_6809),
		.dout(new_net_6808)
	);

	bfr new_net_6810_bfr_before (
		.din(new_net_6810),
		.dout(new_net_6809)
	);

	bfr new_net_6811_bfr_before (
		.din(new_net_6811),
		.dout(new_net_6810)
	);

	bfr new_net_6812_bfr_before (
		.din(new_net_6812),
		.dout(new_net_6811)
	);

	bfr new_net_6813_bfr_before (
		.din(new_net_6813),
		.dout(new_net_6812)
	);

	bfr new_net_6814_bfr_before (
		.din(new_net_6814),
		.dout(new_net_6813)
	);

	bfr new_net_6815_bfr_before (
		.din(new_net_6815),
		.dout(new_net_6814)
	);

	bfr new_net_6816_bfr_before (
		.din(new_net_6816),
		.dout(new_net_6815)
	);

	bfr new_net_6817_bfr_before (
		.din(new_net_6817),
		.dout(new_net_6816)
	);

	bfr new_net_6818_bfr_before (
		.din(new_net_6818),
		.dout(new_net_6817)
	);

	bfr new_net_6819_bfr_before (
		.din(new_net_6819),
		.dout(new_net_6818)
	);

	bfr new_net_6820_bfr_before (
		.din(new_net_6820),
		.dout(new_net_6819)
	);

	bfr new_net_6821_bfr_before (
		.din(new_net_6821),
		.dout(new_net_6820)
	);

	bfr new_net_6822_bfr_before (
		.din(new_net_6822),
		.dout(new_net_6821)
	);

	bfr new_net_6823_bfr_before (
		.din(new_net_6823),
		.dout(new_net_6822)
	);

	bfr new_net_6824_bfr_before (
		.din(new_net_6824),
		.dout(new_net_6823)
	);

	bfr new_net_6825_bfr_before (
		.din(new_net_6825),
		.dout(new_net_6824)
	);

	bfr new_net_6826_bfr_before (
		.din(new_net_6826),
		.dout(new_net_6825)
	);

	bfr new_net_6827_bfr_before (
		.din(new_net_6827),
		.dout(new_net_6826)
	);

	bfr new_net_6828_bfr_before (
		.din(new_net_6828),
		.dout(new_net_6827)
	);

	bfr new_net_6829_bfr_before (
		.din(new_net_6829),
		.dout(new_net_6828)
	);

	bfr new_net_6830_bfr_before (
		.din(new_net_6830),
		.dout(new_net_6829)
	);

	bfr new_net_6831_bfr_before (
		.din(new_net_6831),
		.dout(new_net_6830)
	);

	bfr new_net_6832_bfr_before (
		.din(new_net_6832),
		.dout(new_net_6831)
	);

	bfr new_net_6833_bfr_before (
		.din(new_net_6833),
		.dout(new_net_6832)
	);

	bfr new_net_6834_bfr_before (
		.din(new_net_6834),
		.dout(new_net_6833)
	);

	bfr new_net_6835_bfr_before (
		.din(new_net_6835),
		.dout(new_net_6834)
	);

	bfr new_net_6836_bfr_before (
		.din(new_net_6836),
		.dout(new_net_6835)
	);

	bfr new_net_6837_bfr_before (
		.din(new_net_6837),
		.dout(new_net_6836)
	);

	bfr new_net_6838_bfr_before (
		.din(new_net_6838),
		.dout(new_net_6837)
	);

	bfr new_net_6839_bfr_before (
		.din(new_net_6839),
		.dout(new_net_6838)
	);

	bfr new_net_6840_bfr_before (
		.din(new_net_6840),
		.dout(new_net_6839)
	);

	bfr new_net_6841_bfr_before (
		.din(new_net_6841),
		.dout(new_net_6840)
	);

	bfr new_net_6842_bfr_before (
		.din(new_net_6842),
		.dout(new_net_6841)
	);

	bfr new_net_6843_bfr_before (
		.din(new_net_6843),
		.dout(new_net_6842)
	);

	bfr new_net_6844_bfr_before (
		.din(new_net_6844),
		.dout(new_net_6843)
	);

	bfr new_net_6845_bfr_before (
		.din(new_net_6845),
		.dout(new_net_6844)
	);

	bfr new_net_6846_bfr_before (
		.din(new_net_6846),
		.dout(new_net_6845)
	);

	bfr new_net_6847_bfr_before (
		.din(new_net_6847),
		.dout(new_net_6846)
	);

	bfr new_net_6848_bfr_before (
		.din(new_net_6848),
		.dout(new_net_6847)
	);

	bfr new_net_6849_bfr_before (
		.din(new_net_6849),
		.dout(new_net_6848)
	);

	bfr new_net_6850_bfr_before (
		.din(new_net_6850),
		.dout(new_net_6849)
	);

	spl2 new_net_2047_v_fanout (
		.a(new_net_2047),
		.b(new_net_6850),
		.c(new_net_1895)
	);

	spl4L new_net_1981_v_fanout (
		.a(new_net_1981),
		.b(new_net_183),
		.c(new_net_162),
		.d(new_net_141),
		.e(new_net_136)
	);

	spl4L new_net_1976_v_fanout (
		.a(new_net_1976),
		.b(new_net_184),
		.c(new_net_266),
		.d(new_net_224),
		.e(new_net_203)
	);

	spl4L new_net_1971_v_fanout (
		.a(new_net_1971),
		.b(new_net_154),
		.c(new_net_284),
		.d(new_net_175),
		.e(new_net_242)
	);

	bfr new_net_6851_bfr_before (
		.din(new_net_6851),
		.dout(N571)
	);

	bfr new_net_6852_bfr_before (
		.din(new_net_6852),
		.dout(new_net_6851)
	);

	bfr new_net_6853_bfr_before (
		.din(new_net_6853),
		.dout(new_net_6852)
	);

	bfr new_net_6854_bfr_before (
		.din(new_net_6854),
		.dout(new_net_6853)
	);

	bfr new_net_6855_bfr_before (
		.din(new_net_6855),
		.dout(new_net_6854)
	);

	bfr new_net_6856_bfr_before (
		.din(new_net_6856),
		.dout(new_net_6855)
	);

	bfr new_net_6857_bfr_before (
		.din(new_net_6857),
		.dout(new_net_6856)
	);

	bfr new_net_6858_bfr_before (
		.din(new_net_6858),
		.dout(new_net_6857)
	);

	bfr new_net_6859_bfr_before (
		.din(new_net_6859),
		.dout(new_net_6858)
	);

	bfr new_net_6860_bfr_before (
		.din(new_net_6860),
		.dout(new_net_6859)
	);

	bfr new_net_6861_bfr_before (
		.din(new_net_6861),
		.dout(new_net_6860)
	);

	bfr new_net_6862_bfr_before (
		.din(new_net_6862),
		.dout(new_net_6861)
	);

	bfr new_net_6863_bfr_before (
		.din(new_net_6863),
		.dout(new_net_6862)
	);

	bfr new_net_6864_bfr_before (
		.din(new_net_6864),
		.dout(new_net_6863)
	);

	bfr new_net_6865_bfr_before (
		.din(new_net_6865),
		.dout(new_net_6864)
	);

	bfr new_net_6866_bfr_before (
		.din(new_net_6866),
		.dout(new_net_6865)
	);

	bfr new_net_6867_bfr_before (
		.din(new_net_6867),
		.dout(new_net_6866)
	);

	bfr new_net_6868_bfr_before (
		.din(new_net_6868),
		.dout(new_net_6867)
	);

	bfr new_net_6869_bfr_before (
		.din(new_net_6869),
		.dout(new_net_6868)
	);

	bfr new_net_6870_bfr_before (
		.din(new_net_6870),
		.dout(new_net_6869)
	);

	bfr new_net_6871_bfr_before (
		.din(new_net_6871),
		.dout(new_net_6870)
	);

	bfr new_net_6872_bfr_before (
		.din(new_net_6872),
		.dout(new_net_6871)
	);

	bfr new_net_6873_bfr_before (
		.din(new_net_6873),
		.dout(new_net_6872)
	);

	bfr new_net_6874_bfr_before (
		.din(new_net_6874),
		.dout(new_net_6873)
	);

	bfr new_net_6875_bfr_before (
		.din(new_net_6875),
		.dout(new_net_6874)
	);

	bfr new_net_6876_bfr_before (
		.din(new_net_6876),
		.dout(new_net_6875)
	);

	bfr new_net_6877_bfr_before (
		.din(new_net_6877),
		.dout(new_net_6876)
	);

	bfr new_net_6878_bfr_before (
		.din(new_net_6878),
		.dout(new_net_6877)
	);

	bfr new_net_6879_bfr_before (
		.din(new_net_6879),
		.dout(new_net_6878)
	);

	bfr new_net_6880_bfr_before (
		.din(new_net_6880),
		.dout(new_net_6879)
	);

	bfr new_net_6881_bfr_before (
		.din(new_net_6881),
		.dout(new_net_6880)
	);

	bfr new_net_6882_bfr_before (
		.din(new_net_6882),
		.dout(new_net_6881)
	);

	bfr new_net_6883_bfr_before (
		.din(new_net_6883),
		.dout(new_net_6882)
	);

	bfr new_net_6884_bfr_before (
		.din(new_net_6884),
		.dout(new_net_6883)
	);

	bfr new_net_6885_bfr_before (
		.din(new_net_6885),
		.dout(new_net_6884)
	);

	bfr new_net_6886_bfr_before (
		.din(new_net_6886),
		.dout(new_net_6885)
	);

	bfr new_net_6887_bfr_before (
		.din(new_net_6887),
		.dout(new_net_6886)
	);

	bfr new_net_6888_bfr_before (
		.din(new_net_6888),
		.dout(new_net_6887)
	);

	bfr new_net_6889_bfr_before (
		.din(new_net_6889),
		.dout(new_net_6888)
	);

	bfr new_net_6890_bfr_before (
		.din(new_net_6890),
		.dout(new_net_6889)
	);

	bfr new_net_6891_bfr_before (
		.din(new_net_6891),
		.dout(new_net_6890)
	);

	bfr new_net_6892_bfr_before (
		.din(new_net_6892),
		.dout(new_net_6891)
	);

	bfr new_net_6893_bfr_before (
		.din(new_net_6893),
		.dout(new_net_6892)
	);

	bfr new_net_6894_bfr_before (
		.din(new_net_6894),
		.dout(new_net_6893)
	);

	bfr new_net_6895_bfr_before (
		.din(new_net_6895),
		.dout(new_net_6894)
	);

	bfr new_net_6896_bfr_before (
		.din(new_net_6896),
		.dout(new_net_6895)
	);

	bfr new_net_6897_bfr_before (
		.din(new_net_6897),
		.dout(new_net_6896)
	);

	bfr new_net_6898_bfr_before (
		.din(new_net_6898),
		.dout(new_net_6897)
	);

	bfr new_net_6899_bfr_before (
		.din(new_net_6899),
		.dout(new_net_6898)
	);

	bfr new_net_6900_bfr_before (
		.din(new_net_6900),
		.dout(new_net_6899)
	);

	bfr new_net_6901_bfr_before (
		.din(new_net_6901),
		.dout(new_net_6900)
	);

	bfr new_net_6902_bfr_before (
		.din(new_net_6902),
		.dout(new_net_6901)
	);

	bfr new_net_6903_bfr_before (
		.din(new_net_6903),
		.dout(new_net_6902)
	);

	bfr new_net_6904_bfr_before (
		.din(new_net_6904),
		.dout(new_net_6903)
	);

	bfr new_net_6905_bfr_before (
		.din(new_net_6905),
		.dout(new_net_6904)
	);

	bfr new_net_6906_bfr_before (
		.din(new_net_6906),
		.dout(new_net_6905)
	);

	bfr new_net_6907_bfr_before (
		.din(new_net_6907),
		.dout(new_net_6906)
	);

	bfr new_net_6908_bfr_before (
		.din(new_net_6908),
		.dout(new_net_6907)
	);

	bfr new_net_6909_bfr_before (
		.din(new_net_6909),
		.dout(new_net_6908)
	);

	bfr new_net_6910_bfr_before (
		.din(new_net_6910),
		.dout(new_net_6909)
	);

	bfr new_net_6911_bfr_before (
		.din(new_net_6911),
		.dout(new_net_6910)
	);

	bfr new_net_6912_bfr_before (
		.din(new_net_6912),
		.dout(new_net_6911)
	);

	spl2 new_net_2052_v_fanout (
		.a(new_net_2052),
		.b(new_net_6912),
		.c(new_net_1719)
	);

	spl4L new_net_2005_v_fanout (
		.a(new_net_2005),
		.b(new_net_228),
		.c(new_net_270),
		.d(new_net_197),
		.e(new_net_279)
	);

	spl4L new_net_1995_v_fanout (
		.a(new_net_1995),
		.b(new_net_168),
		.c(new_net_147),
		.d(new_net_181),
		.e(new_net_160)
	);

	spl4L new_net_2011_v_fanout (
		.a(new_net_2011),
		.b(new_net_227),
		.c(new_net_278),
		.d(new_net_236),
		.e(new_net_215)
	);

	spl4L new_net_2007_v_fanout (
		.a(new_net_2007),
		.b(new_net_166),
		.c(new_net_187),
		.d(new_net_145),
		.e(new_net_132)
	);

	spl4L new_net_2013_v_fanout (
		.a(new_net_2013),
		.b(new_net_119),
		.c(new_net_177),
		.d(new_net_190),
		.e(new_net_156)
	);

	bfr new_net_6913_bfr_before (
		.din(new_net_6913),
		.dout(N569)
	);

	bfr new_net_6914_bfr_before (
		.din(new_net_6914),
		.dout(new_net_6913)
	);

	bfr new_net_6915_bfr_before (
		.din(new_net_6915),
		.dout(new_net_6914)
	);

	bfr new_net_6916_bfr_before (
		.din(new_net_6916),
		.dout(new_net_6915)
	);

	bfr new_net_6917_bfr_before (
		.din(new_net_6917),
		.dout(new_net_6916)
	);

	bfr new_net_6918_bfr_before (
		.din(new_net_6918),
		.dout(new_net_6917)
	);

	bfr new_net_6919_bfr_before (
		.din(new_net_6919),
		.dout(new_net_6918)
	);

	bfr new_net_6920_bfr_before (
		.din(new_net_6920),
		.dout(new_net_6919)
	);

	bfr new_net_6921_bfr_before (
		.din(new_net_6921),
		.dout(new_net_6920)
	);

	bfr new_net_6922_bfr_before (
		.din(new_net_6922),
		.dout(new_net_6921)
	);

	bfr new_net_6923_bfr_before (
		.din(new_net_6923),
		.dout(new_net_6922)
	);

	bfr new_net_6924_bfr_before (
		.din(new_net_6924),
		.dout(new_net_6923)
	);

	bfr new_net_6925_bfr_before (
		.din(new_net_6925),
		.dout(new_net_6924)
	);

	bfr new_net_6926_bfr_before (
		.din(new_net_6926),
		.dout(new_net_6925)
	);

	bfr new_net_6927_bfr_before (
		.din(new_net_6927),
		.dout(new_net_6926)
	);

	bfr new_net_6928_bfr_before (
		.din(new_net_6928),
		.dout(new_net_6927)
	);

	bfr new_net_6929_bfr_before (
		.din(new_net_6929),
		.dout(new_net_6928)
	);

	bfr new_net_6930_bfr_before (
		.din(new_net_6930),
		.dout(new_net_6929)
	);

	bfr new_net_6931_bfr_before (
		.din(new_net_6931),
		.dout(new_net_6930)
	);

	bfr new_net_6932_bfr_before (
		.din(new_net_6932),
		.dout(new_net_6931)
	);

	bfr new_net_6933_bfr_before (
		.din(new_net_6933),
		.dout(new_net_6932)
	);

	bfr new_net_6934_bfr_before (
		.din(new_net_6934),
		.dout(new_net_6933)
	);

	bfr new_net_6935_bfr_before (
		.din(new_net_6935),
		.dout(new_net_6934)
	);

	bfr new_net_6936_bfr_before (
		.din(new_net_6936),
		.dout(new_net_6935)
	);

	bfr new_net_6937_bfr_before (
		.din(new_net_6937),
		.dout(new_net_6936)
	);

	bfr new_net_6938_bfr_before (
		.din(new_net_6938),
		.dout(new_net_6937)
	);

	bfr new_net_6939_bfr_before (
		.din(new_net_6939),
		.dout(new_net_6938)
	);

	bfr new_net_6940_bfr_before (
		.din(new_net_6940),
		.dout(new_net_6939)
	);

	bfr new_net_6941_bfr_before (
		.din(new_net_6941),
		.dout(new_net_6940)
	);

	bfr new_net_6942_bfr_before (
		.din(new_net_6942),
		.dout(new_net_6941)
	);

	bfr new_net_6943_bfr_before (
		.din(new_net_6943),
		.dout(new_net_6942)
	);

	bfr new_net_6944_bfr_before (
		.din(new_net_6944),
		.dout(new_net_6943)
	);

	bfr new_net_6945_bfr_before (
		.din(new_net_6945),
		.dout(new_net_6944)
	);

	bfr new_net_6946_bfr_before (
		.din(new_net_6946),
		.dout(new_net_6945)
	);

	bfr new_net_6947_bfr_before (
		.din(new_net_6947),
		.dout(new_net_6946)
	);

	bfr new_net_6948_bfr_before (
		.din(new_net_6948),
		.dout(new_net_6947)
	);

	bfr new_net_6949_bfr_before (
		.din(new_net_6949),
		.dout(new_net_6948)
	);

	bfr new_net_6950_bfr_before (
		.din(new_net_6950),
		.dout(new_net_6949)
	);

	bfr new_net_6951_bfr_before (
		.din(new_net_6951),
		.dout(new_net_6950)
	);

	bfr new_net_6952_bfr_before (
		.din(new_net_6952),
		.dout(new_net_6951)
	);

	bfr new_net_6953_bfr_before (
		.din(new_net_6953),
		.dout(new_net_6952)
	);

	bfr new_net_6954_bfr_before (
		.din(new_net_6954),
		.dout(new_net_6953)
	);

	bfr new_net_6955_bfr_before (
		.din(new_net_6955),
		.dout(new_net_6954)
	);

	bfr new_net_6956_bfr_before (
		.din(new_net_6956),
		.dout(new_net_6955)
	);

	bfr new_net_6957_bfr_before (
		.din(new_net_6957),
		.dout(new_net_6956)
	);

	bfr new_net_6958_bfr_before (
		.din(new_net_6958),
		.dout(new_net_6957)
	);

	bfr new_net_6959_bfr_before (
		.din(new_net_6959),
		.dout(new_net_6958)
	);

	bfr new_net_6960_bfr_before (
		.din(new_net_6960),
		.dout(new_net_6959)
	);

	bfr new_net_6961_bfr_before (
		.din(new_net_6961),
		.dout(new_net_6960)
	);

	bfr new_net_6962_bfr_before (
		.din(new_net_6962),
		.dout(new_net_6961)
	);

	bfr new_net_6963_bfr_before (
		.din(new_net_6963),
		.dout(new_net_6962)
	);

	bfr new_net_6964_bfr_before (
		.din(new_net_6964),
		.dout(new_net_6963)
	);

	bfr new_net_6965_bfr_before (
		.din(new_net_6965),
		.dout(new_net_6964)
	);

	bfr new_net_6966_bfr_before (
		.din(new_net_6966),
		.dout(new_net_6965)
	);

	bfr new_net_6967_bfr_before (
		.din(new_net_6967),
		.dout(new_net_6966)
	);

	bfr new_net_6968_bfr_before (
		.din(new_net_6968),
		.dout(new_net_6967)
	);

	bfr new_net_6969_bfr_before (
		.din(new_net_6969),
		.dout(new_net_6968)
	);

	bfr new_net_6970_bfr_before (
		.din(new_net_6970),
		.dout(new_net_6969)
	);

	bfr new_net_6971_bfr_before (
		.din(new_net_6971),
		.dout(new_net_6970)
	);

	bfr new_net_6972_bfr_before (
		.din(new_net_6972),
		.dout(new_net_6971)
	);

	bfr new_net_6973_bfr_before (
		.din(new_net_6973),
		.dout(new_net_6972)
	);

	bfr new_net_6974_bfr_before (
		.din(new_net_6974),
		.dout(new_net_6973)
	);

	spl2 new_net_2051_v_fanout (
		.a(new_net_2051),
		.b(new_net_6974),
		.c(new_net_650)
	);

	spl4L new_net_1968_v_fanout (
		.a(new_net_1968),
		.b(new_net_213),
		.c(new_net_234),
		.d(new_net_244),
		.e(new_net_214)
	);

	spl4L new_net_1990_v_fanout (
		.a(new_net_1990),
		.b(new_net_222),
		.c(new_net_264),
		.d(new_net_207),
		.e(new_net_201)
	);

	spl4L new_net_1986_v_fanout (
		.a(new_net_1986),
		.b(new_net_200),
		.c(new_net_273),
		.d(new_net_231),
		.e(new_net_210)
	);

	spl4L new_net_1991_v_fanout (
		.a(new_net_1991),
		.b(new_net_218),
		.c(new_net_239),
		.d(new_net_249),
		.e(new_net_258)
	);

	bfr new_net_6975_bfr_before (
		.din(new_net_6975),
		.dout(N707)
	);

	bfr new_net_6976_bfr_before (
		.din(new_net_6976),
		.dout(new_net_6975)
	);

	bfr new_net_6977_bfr_before (
		.din(new_net_6977),
		.dout(new_net_6976)
	);

	bfr new_net_6978_bfr_before (
		.din(new_net_6978),
		.dout(new_net_6977)
	);

	bfr new_net_6979_bfr_before (
		.din(new_net_6979),
		.dout(new_net_6978)
	);

	bfr new_net_6980_bfr_before (
		.din(new_net_6980),
		.dout(new_net_6979)
	);

	bfr new_net_6981_bfr_before (
		.din(new_net_6981),
		.dout(new_net_6980)
	);

	bfr new_net_6982_bfr_before (
		.din(new_net_6982),
		.dout(new_net_6981)
	);

	bfr new_net_6983_bfr_before (
		.din(new_net_6983),
		.dout(new_net_6982)
	);

	bfr new_net_6984_bfr_before (
		.din(new_net_6984),
		.dout(new_net_6983)
	);

	bfr new_net_6985_bfr_before (
		.din(new_net_6985),
		.dout(new_net_6984)
	);

	bfr new_net_6986_bfr_before (
		.din(new_net_6986),
		.dout(new_net_6985)
	);

	bfr new_net_6987_bfr_before (
		.din(new_net_6987),
		.dout(new_net_6986)
	);

	bfr new_net_6988_bfr_before (
		.din(new_net_6988),
		.dout(new_net_6987)
	);

	bfr new_net_6989_bfr_before (
		.din(new_net_6989),
		.dout(new_net_6988)
	);

	bfr new_net_6990_bfr_before (
		.din(new_net_6990),
		.dout(new_net_6989)
	);

	bfr new_net_6991_bfr_before (
		.din(new_net_6991),
		.dout(new_net_6990)
	);

	bfr new_net_6992_bfr_before (
		.din(new_net_6992),
		.dout(new_net_6991)
	);

	bfr new_net_6993_bfr_before (
		.din(new_net_6993),
		.dout(new_net_6992)
	);

	bfr new_net_6994_bfr_before (
		.din(new_net_6994),
		.dout(new_net_6993)
	);

	bfr new_net_6995_bfr_before (
		.din(new_net_6995),
		.dout(new_net_6994)
	);

	bfr new_net_6996_bfr_before (
		.din(new_net_6996),
		.dout(new_net_6995)
	);

	bfr new_net_6997_bfr_before (
		.din(new_net_6997),
		.dout(new_net_6996)
	);

	bfr new_net_6998_bfr_before (
		.din(new_net_6998),
		.dout(new_net_6997)
	);

	bfr new_net_6999_bfr_before (
		.din(new_net_6999),
		.dout(new_net_6998)
	);

	bfr new_net_7000_bfr_before (
		.din(new_net_7000),
		.dout(new_net_6999)
	);

	bfr new_net_7001_bfr_before (
		.din(new_net_7001),
		.dout(new_net_7000)
	);

	bfr new_net_7002_bfr_before (
		.din(new_net_7002),
		.dout(new_net_7001)
	);

	bfr new_net_7003_bfr_before (
		.din(new_net_7003),
		.dout(new_net_7002)
	);

	bfr new_net_7004_bfr_before (
		.din(new_net_7004),
		.dout(new_net_7003)
	);

	bfr new_net_7005_bfr_before (
		.din(new_net_7005),
		.dout(new_net_7004)
	);

	bfr new_net_7006_bfr_before (
		.din(new_net_7006),
		.dout(new_net_7005)
	);

	bfr new_net_7007_bfr_before (
		.din(new_net_7007),
		.dout(new_net_7006)
	);

	bfr new_net_7008_bfr_before (
		.din(new_net_7008),
		.dout(new_net_7007)
	);

	bfr new_net_7009_bfr_before (
		.din(new_net_7009),
		.dout(new_net_7008)
	);

	bfr new_net_7010_bfr_before (
		.din(new_net_7010),
		.dout(new_net_7009)
	);

	bfr new_net_7011_bfr_before (
		.din(new_net_7011),
		.dout(new_net_7010)
	);

	bfr new_net_7012_bfr_before (
		.din(new_net_7012),
		.dout(new_net_7011)
	);

	bfr new_net_7013_bfr_before (
		.din(new_net_7013),
		.dout(new_net_7012)
	);

	bfr new_net_7014_bfr_before (
		.din(new_net_7014),
		.dout(new_net_7013)
	);

	bfr new_net_7015_bfr_before (
		.din(new_net_7015),
		.dout(new_net_7014)
	);

	bfr new_net_7016_bfr_before (
		.din(new_net_7016),
		.dout(new_net_7015)
	);

	bfr new_net_7017_bfr_before (
		.din(new_net_7017),
		.dout(new_net_7016)
	);

	bfr new_net_7018_bfr_before (
		.din(new_net_7018),
		.dout(new_net_7017)
	);

	bfr new_net_7019_bfr_before (
		.din(new_net_7019),
		.dout(new_net_7018)
	);

	bfr new_net_7020_bfr_before (
		.din(new_net_7020),
		.dout(new_net_7019)
	);

	bfr new_net_7021_bfr_before (
		.din(new_net_7021),
		.dout(new_net_7020)
	);

	bfr new_net_7022_bfr_before (
		.din(new_net_7022),
		.dout(new_net_7021)
	);

	bfr new_net_7023_bfr_before (
		.din(new_net_7023),
		.dout(new_net_7022)
	);

	bfr new_net_7024_bfr_before (
		.din(new_net_7024),
		.dout(new_net_7023)
	);

	bfr new_net_7025_bfr_before (
		.din(new_net_7025),
		.dout(new_net_7024)
	);

	bfr new_net_7026_bfr_before (
		.din(new_net_7026),
		.dout(new_net_7025)
	);

	bfr new_net_7027_bfr_before (
		.din(new_net_7027),
		.dout(new_net_7026)
	);

	bfr new_net_7028_bfr_before (
		.din(new_net_7028),
		.dout(new_net_7027)
	);

	bfr new_net_7029_bfr_before (
		.din(new_net_7029),
		.dout(new_net_7028)
	);

	bfr new_net_7030_bfr_before (
		.din(new_net_7030),
		.dout(new_net_7029)
	);

	bfr new_net_7031_bfr_before (
		.din(new_net_7031),
		.dout(new_net_7030)
	);

	bfr new_net_7032_bfr_before (
		.din(new_net_7032),
		.dout(new_net_7031)
	);

	bfr new_net_7033_bfr_before (
		.din(new_net_7033),
		.dout(new_net_7032)
	);

	bfr new_net_7034_bfr_before (
		.din(new_net_7034),
		.dout(new_net_7033)
	);

	bfr new_net_7035_bfr_before (
		.din(new_net_7035),
		.dout(new_net_7034)
	);

	bfr new_net_7036_bfr_before (
		.din(new_net_7036),
		.dout(new_net_7035)
	);

	spl2 new_net_2026_v_fanout (
		.a(new_net_2026),
		.b(new_net_7036),
		.c(new_net_1144)
	);

	spl4L new_net_1970_v_fanout (
		.a(new_net_1970),
		.b(new_net_221),
		.c(new_net_261),
		.d(new_net_252),
		.e(new_net_267)
	);

	spl4L new_net_1997_v_fanout (
		.a(new_net_1997),
		.b(new_net_217),
		.c(new_net_238),
		.d(new_net_280),
		.e(new_net_248)
	);

	spl4L new_net_1969_v_fanout (
		.a(new_net_1969),
		.b(new_net_204),
		.c(new_net_225),
		.d(new_net_286),
		.e(new_net_276)
	);

	bfr new_net_7037_bfr_before (
		.din(new_net_7037),
		.dout(N547)
	);

	bfr new_net_7038_bfr_before (
		.din(new_net_7038),
		.dout(new_net_7037)
	);

	bfr new_net_7039_bfr_before (
		.din(new_net_7039),
		.dout(new_net_7038)
	);

	bfr new_net_7040_bfr_before (
		.din(new_net_7040),
		.dout(new_net_7039)
	);

	bfr new_net_7041_bfr_before (
		.din(new_net_7041),
		.dout(new_net_7040)
	);

	bfr new_net_7042_bfr_before (
		.din(new_net_7042),
		.dout(new_net_7041)
	);

	bfr new_net_7043_bfr_before (
		.din(new_net_7043),
		.dout(new_net_7042)
	);

	bfr new_net_7044_bfr_before (
		.din(new_net_7044),
		.dout(new_net_7043)
	);

	bfr new_net_7045_bfr_before (
		.din(new_net_7045),
		.dout(new_net_7044)
	);

	bfr new_net_7046_bfr_before (
		.din(new_net_7046),
		.dout(new_net_7045)
	);

	bfr new_net_7047_bfr_before (
		.din(new_net_7047),
		.dout(new_net_7046)
	);

	bfr new_net_7048_bfr_before (
		.din(new_net_7048),
		.dout(new_net_7047)
	);

	bfr new_net_7049_bfr_before (
		.din(new_net_7049),
		.dout(new_net_7048)
	);

	bfr new_net_7050_bfr_before (
		.din(new_net_7050),
		.dout(new_net_7049)
	);

	bfr new_net_7051_bfr_before (
		.din(new_net_7051),
		.dout(new_net_7050)
	);

	bfr new_net_7052_bfr_before (
		.din(new_net_7052),
		.dout(new_net_7051)
	);

	bfr new_net_7053_bfr_before (
		.din(new_net_7053),
		.dout(new_net_7052)
	);

	bfr new_net_7054_bfr_before (
		.din(new_net_7054),
		.dout(new_net_7053)
	);

	bfr new_net_7055_bfr_before (
		.din(new_net_7055),
		.dout(new_net_7054)
	);

	bfr new_net_7056_bfr_before (
		.din(new_net_7056),
		.dout(new_net_7055)
	);

	bfr new_net_7057_bfr_before (
		.din(new_net_7057),
		.dout(new_net_7056)
	);

	bfr new_net_7058_bfr_before (
		.din(new_net_7058),
		.dout(new_net_7057)
	);

	bfr new_net_7059_bfr_before (
		.din(new_net_7059),
		.dout(new_net_7058)
	);

	bfr new_net_7060_bfr_before (
		.din(new_net_7060),
		.dout(new_net_7059)
	);

	bfr new_net_7061_bfr_before (
		.din(new_net_7061),
		.dout(new_net_7060)
	);

	bfr new_net_7062_bfr_before (
		.din(new_net_7062),
		.dout(new_net_7061)
	);

	bfr new_net_7063_bfr_before (
		.din(new_net_7063),
		.dout(new_net_7062)
	);

	bfr new_net_7064_bfr_before (
		.din(new_net_7064),
		.dout(new_net_7063)
	);

	bfr new_net_7065_bfr_before (
		.din(new_net_7065),
		.dout(new_net_7064)
	);

	bfr new_net_7066_bfr_before (
		.din(new_net_7066),
		.dout(new_net_7065)
	);

	bfr new_net_7067_bfr_before (
		.din(new_net_7067),
		.dout(new_net_7066)
	);

	bfr new_net_7068_bfr_before (
		.din(new_net_7068),
		.dout(new_net_7067)
	);

	bfr new_net_7069_bfr_before (
		.din(new_net_7069),
		.dout(new_net_7068)
	);

	bfr new_net_7070_bfr_before (
		.din(new_net_7070),
		.dout(new_net_7069)
	);

	bfr new_net_7071_bfr_before (
		.din(new_net_7071),
		.dout(new_net_7070)
	);

	bfr new_net_7072_bfr_before (
		.din(new_net_7072),
		.dout(new_net_7071)
	);

	bfr new_net_7073_bfr_before (
		.din(new_net_7073),
		.dout(new_net_7072)
	);

	bfr new_net_7074_bfr_before (
		.din(new_net_7074),
		.dout(new_net_7073)
	);

	bfr new_net_7075_bfr_before (
		.din(new_net_7075),
		.dout(new_net_7074)
	);

	bfr new_net_7076_bfr_before (
		.din(new_net_7076),
		.dout(new_net_7075)
	);

	bfr new_net_7077_bfr_before (
		.din(new_net_7077),
		.dout(new_net_7076)
	);

	bfr new_net_7078_bfr_before (
		.din(new_net_7078),
		.dout(new_net_7077)
	);

	bfr new_net_7079_bfr_before (
		.din(new_net_7079),
		.dout(new_net_7078)
	);

	bfr new_net_7080_bfr_before (
		.din(new_net_7080),
		.dout(new_net_7079)
	);

	bfr new_net_7081_bfr_before (
		.din(new_net_7081),
		.dout(new_net_7080)
	);

	bfr new_net_7082_bfr_before (
		.din(new_net_7082),
		.dout(new_net_7081)
	);

	bfr new_net_7083_bfr_before (
		.din(new_net_7083),
		.dout(new_net_7082)
	);

	bfr new_net_7084_bfr_before (
		.din(new_net_7084),
		.dout(new_net_7083)
	);

	bfr new_net_7085_bfr_before (
		.din(new_net_7085),
		.dout(new_net_7084)
	);

	bfr new_net_7086_bfr_before (
		.din(new_net_7086),
		.dout(new_net_7085)
	);

	bfr new_net_7087_bfr_before (
		.din(new_net_7087),
		.dout(new_net_7086)
	);

	bfr new_net_7088_bfr_before (
		.din(new_net_7088),
		.dout(new_net_7087)
	);

	bfr new_net_7089_bfr_before (
		.din(new_net_7089),
		.dout(new_net_7088)
	);

	bfr new_net_7090_bfr_before (
		.din(new_net_7090),
		.dout(new_net_7089)
	);

	bfr new_net_7091_bfr_before (
		.din(new_net_7091),
		.dout(new_net_7090)
	);

	bfr new_net_7092_bfr_before (
		.din(new_net_7092),
		.dout(new_net_7091)
	);

	bfr new_net_7093_bfr_before (
		.din(new_net_7093),
		.dout(new_net_7092)
	);

	bfr new_net_7094_bfr_before (
		.din(new_net_7094),
		.dout(new_net_7093)
	);

	bfr new_net_7095_bfr_before (
		.din(new_net_7095),
		.dout(new_net_7094)
	);

	bfr new_net_7096_bfr_before (
		.din(new_net_7096),
		.dout(new_net_7095)
	);

	bfr new_net_7097_bfr_before (
		.din(new_net_7097),
		.dout(new_net_7096)
	);

	bfr new_net_7098_bfr_before (
		.din(new_net_7098),
		.dout(new_net_7097)
	);

	spl2 new_net_2041_v_fanout (
		.a(new_net_2041),
		.b(new_net_7098),
		.c(new_net_1432)
	);

	spl4L new_net_2010_v_fanout (
		.a(new_net_2010),
		.b(new_net_288),
		.c(new_net_255),
		.d(new_net_246),
		.e(new_net_216)
	);

	spl4L new_net_1974_v_fanout (
		.a(new_net_1974),
		.b(new_net_188),
		.c(new_net_167),
		.d(new_net_212),
		.e(new_net_146)
	);

	spl4L new_net_2015_v_fanout (
		.a(new_net_2015),
		.b(new_net_135),
		.c(new_net_140),
		.d(new_net_161),
		.e(new_net_127)
	);

	spl4L new_net_2018_v_fanout (
		.a(new_net_2018),
		.b(new_net_268),
		.c(new_net_2019),
		.d(new_net_253),
		.e(new_net_262)
	);

	bfr new_net_7099_bfr_before (
		.din(new_net_7099),
		.dout(N553)
	);

	bfr new_net_7100_bfr_before (
		.din(new_net_7100),
		.dout(new_net_7099)
	);

	bfr new_net_7101_bfr_before (
		.din(new_net_7101),
		.dout(new_net_7100)
	);

	bfr new_net_7102_bfr_before (
		.din(new_net_7102),
		.dout(new_net_7101)
	);

	bfr new_net_7103_bfr_before (
		.din(new_net_7103),
		.dout(new_net_7102)
	);

	bfr new_net_7104_bfr_before (
		.din(new_net_7104),
		.dout(new_net_7103)
	);

	bfr new_net_7105_bfr_before (
		.din(new_net_7105),
		.dout(new_net_7104)
	);

	bfr new_net_7106_bfr_before (
		.din(new_net_7106),
		.dout(new_net_7105)
	);

	bfr new_net_7107_bfr_before (
		.din(new_net_7107),
		.dout(new_net_7106)
	);

	bfr new_net_7108_bfr_before (
		.din(new_net_7108),
		.dout(new_net_7107)
	);

	bfr new_net_7109_bfr_before (
		.din(new_net_7109),
		.dout(new_net_7108)
	);

	bfr new_net_7110_bfr_before (
		.din(new_net_7110),
		.dout(new_net_7109)
	);

	bfr new_net_7111_bfr_before (
		.din(new_net_7111),
		.dout(new_net_7110)
	);

	bfr new_net_7112_bfr_before (
		.din(new_net_7112),
		.dout(new_net_7111)
	);

	bfr new_net_7113_bfr_before (
		.din(new_net_7113),
		.dout(new_net_7112)
	);

	bfr new_net_7114_bfr_before (
		.din(new_net_7114),
		.dout(new_net_7113)
	);

	bfr new_net_7115_bfr_before (
		.din(new_net_7115),
		.dout(new_net_7114)
	);

	bfr new_net_7116_bfr_before (
		.din(new_net_7116),
		.dout(new_net_7115)
	);

	bfr new_net_7117_bfr_before (
		.din(new_net_7117),
		.dout(new_net_7116)
	);

	bfr new_net_7118_bfr_before (
		.din(new_net_7118),
		.dout(new_net_7117)
	);

	bfr new_net_7119_bfr_before (
		.din(new_net_7119),
		.dout(new_net_7118)
	);

	bfr new_net_7120_bfr_before (
		.din(new_net_7120),
		.dout(new_net_7119)
	);

	bfr new_net_7121_bfr_before (
		.din(new_net_7121),
		.dout(new_net_7120)
	);

	bfr new_net_7122_bfr_before (
		.din(new_net_7122),
		.dout(new_net_7121)
	);

	bfr new_net_7123_bfr_before (
		.din(new_net_7123),
		.dout(new_net_7122)
	);

	bfr new_net_7124_bfr_before (
		.din(new_net_7124),
		.dout(new_net_7123)
	);

	bfr new_net_7125_bfr_before (
		.din(new_net_7125),
		.dout(new_net_7124)
	);

	bfr new_net_7126_bfr_before (
		.din(new_net_7126),
		.dout(new_net_7125)
	);

	bfr new_net_7127_bfr_before (
		.din(new_net_7127),
		.dout(new_net_7126)
	);

	bfr new_net_7128_bfr_before (
		.din(new_net_7128),
		.dout(new_net_7127)
	);

	bfr new_net_7129_bfr_before (
		.din(new_net_7129),
		.dout(new_net_7128)
	);

	bfr new_net_7130_bfr_before (
		.din(new_net_7130),
		.dout(new_net_7129)
	);

	bfr new_net_7131_bfr_before (
		.din(new_net_7131),
		.dout(new_net_7130)
	);

	bfr new_net_7132_bfr_before (
		.din(new_net_7132),
		.dout(new_net_7131)
	);

	bfr new_net_7133_bfr_before (
		.din(new_net_7133),
		.dout(new_net_7132)
	);

	bfr new_net_7134_bfr_before (
		.din(new_net_7134),
		.dout(new_net_7133)
	);

	bfr new_net_7135_bfr_before (
		.din(new_net_7135),
		.dout(new_net_7134)
	);

	bfr new_net_7136_bfr_before (
		.din(new_net_7136),
		.dout(new_net_7135)
	);

	bfr new_net_7137_bfr_before (
		.din(new_net_7137),
		.dout(new_net_7136)
	);

	bfr new_net_7138_bfr_before (
		.din(new_net_7138),
		.dout(new_net_7137)
	);

	bfr new_net_7139_bfr_before (
		.din(new_net_7139),
		.dout(new_net_7138)
	);

	bfr new_net_7140_bfr_before (
		.din(new_net_7140),
		.dout(new_net_7139)
	);

	bfr new_net_7141_bfr_before (
		.din(new_net_7141),
		.dout(new_net_7140)
	);

	bfr new_net_7142_bfr_before (
		.din(new_net_7142),
		.dout(new_net_7141)
	);

	bfr new_net_7143_bfr_before (
		.din(new_net_7143),
		.dout(new_net_7142)
	);

	bfr new_net_7144_bfr_before (
		.din(new_net_7144),
		.dout(new_net_7143)
	);

	bfr new_net_7145_bfr_before (
		.din(new_net_7145),
		.dout(new_net_7144)
	);

	bfr new_net_7146_bfr_before (
		.din(new_net_7146),
		.dout(new_net_7145)
	);

	bfr new_net_7147_bfr_before (
		.din(new_net_7147),
		.dout(new_net_7146)
	);

	bfr new_net_7148_bfr_before (
		.din(new_net_7148),
		.dout(new_net_7147)
	);

	bfr new_net_7149_bfr_before (
		.din(new_net_7149),
		.dout(new_net_7148)
	);

	bfr new_net_7150_bfr_before (
		.din(new_net_7150),
		.dout(new_net_7149)
	);

	bfr new_net_7151_bfr_before (
		.din(new_net_7151),
		.dout(new_net_7150)
	);

	bfr new_net_7152_bfr_before (
		.din(new_net_7152),
		.dout(new_net_7151)
	);

	bfr new_net_7153_bfr_before (
		.din(new_net_7153),
		.dout(new_net_7152)
	);

	bfr new_net_7154_bfr_before (
		.din(new_net_7154),
		.dout(new_net_7153)
	);

	bfr new_net_7155_bfr_before (
		.din(new_net_7155),
		.dout(new_net_7154)
	);

	bfr new_net_7156_bfr_before (
		.din(new_net_7156),
		.dout(new_net_7155)
	);

	bfr new_net_7157_bfr_before (
		.din(new_net_7157),
		.dout(new_net_7156)
	);

	bfr new_net_7158_bfr_before (
		.din(new_net_7158),
		.dout(new_net_7157)
	);

	bfr new_net_7159_bfr_before (
		.din(new_net_7159),
		.dout(new_net_7158)
	);

	bfr new_net_7160_bfr_before (
		.din(new_net_7160),
		.dout(new_net_7159)
	);

	spl2 new_net_2044_v_fanout (
		.a(new_net_2044),
		.b(new_net_7160),
		.c(new_net_1479)
	);

	bfr new_net_7161_bfr_before (
		.din(new_net_7161),
		.dout(N507)
	);

	bfr new_net_7162_bfr_before (
		.din(new_net_7162),
		.dout(new_net_7161)
	);

	bfr new_net_7163_bfr_before (
		.din(new_net_7163),
		.dout(new_net_7162)
	);

	bfr new_net_7164_bfr_before (
		.din(new_net_7164),
		.dout(new_net_7163)
	);

	bfr new_net_7165_bfr_before (
		.din(new_net_7165),
		.dout(new_net_7164)
	);

	bfr new_net_7166_bfr_before (
		.din(new_net_7166),
		.dout(new_net_7165)
	);

	bfr new_net_7167_bfr_before (
		.din(new_net_7167),
		.dout(new_net_7166)
	);

	bfr new_net_7168_bfr_before (
		.din(new_net_7168),
		.dout(new_net_7167)
	);

	bfr new_net_7169_bfr_before (
		.din(new_net_7169),
		.dout(new_net_7168)
	);

	bfr new_net_7170_bfr_before (
		.din(new_net_7170),
		.dout(new_net_7169)
	);

	bfr new_net_7171_bfr_before (
		.din(new_net_7171),
		.dout(new_net_7170)
	);

	bfr new_net_7172_bfr_before (
		.din(new_net_7172),
		.dout(new_net_7171)
	);

	bfr new_net_7173_bfr_before (
		.din(new_net_7173),
		.dout(new_net_7172)
	);

	bfr new_net_7174_bfr_before (
		.din(new_net_7174),
		.dout(new_net_7173)
	);

	bfr new_net_7175_bfr_before (
		.din(new_net_7175),
		.dout(new_net_7174)
	);

	bfr new_net_7176_bfr_before (
		.din(new_net_7176),
		.dout(new_net_7175)
	);

	bfr new_net_7177_bfr_before (
		.din(new_net_7177),
		.dout(new_net_7176)
	);

	bfr new_net_7178_bfr_before (
		.din(new_net_7178),
		.dout(new_net_7177)
	);

	bfr new_net_7179_bfr_before (
		.din(new_net_7179),
		.dout(new_net_7178)
	);

	bfr new_net_7180_bfr_before (
		.din(new_net_7180),
		.dout(new_net_7179)
	);

	bfr new_net_7181_bfr_before (
		.din(new_net_7181),
		.dout(new_net_7180)
	);

	bfr new_net_7182_bfr_before (
		.din(new_net_7182),
		.dout(new_net_7181)
	);

	bfr new_net_7183_bfr_before (
		.din(new_net_7183),
		.dout(new_net_7182)
	);

	bfr new_net_7184_bfr_before (
		.din(new_net_7184),
		.dout(new_net_7183)
	);

	bfr new_net_7185_bfr_before (
		.din(new_net_7185),
		.dout(new_net_7184)
	);

	bfr new_net_7186_bfr_before (
		.din(new_net_7186),
		.dout(new_net_7185)
	);

	bfr new_net_7187_bfr_before (
		.din(new_net_7187),
		.dout(new_net_7186)
	);

	bfr new_net_7188_bfr_before (
		.din(new_net_7188),
		.dout(new_net_7187)
	);

	bfr new_net_7189_bfr_before (
		.din(new_net_7189),
		.dout(new_net_7188)
	);

	bfr new_net_7190_bfr_before (
		.din(new_net_7190),
		.dout(new_net_7189)
	);

	bfr new_net_7191_bfr_before (
		.din(new_net_7191),
		.dout(new_net_7190)
	);

	bfr new_net_7192_bfr_before (
		.din(new_net_7192),
		.dout(new_net_7191)
	);

	bfr new_net_7193_bfr_before (
		.din(new_net_7193),
		.dout(new_net_7192)
	);

	bfr new_net_7194_bfr_before (
		.din(new_net_7194),
		.dout(new_net_7193)
	);

	bfr new_net_7195_bfr_before (
		.din(new_net_7195),
		.dout(new_net_7194)
	);

	bfr new_net_7196_bfr_before (
		.din(new_net_7196),
		.dout(new_net_7195)
	);

	bfr new_net_7197_bfr_before (
		.din(new_net_7197),
		.dout(new_net_7196)
	);

	bfr new_net_7198_bfr_before (
		.din(new_net_7198),
		.dout(new_net_7197)
	);

	bfr new_net_7199_bfr_before (
		.din(new_net_7199),
		.dout(new_net_7198)
	);

	bfr new_net_7200_bfr_before (
		.din(new_net_7200),
		.dout(new_net_7199)
	);

	bfr new_net_7201_bfr_before (
		.din(new_net_7201),
		.dout(new_net_7200)
	);

	bfr new_net_7202_bfr_before (
		.din(new_net_7202),
		.dout(new_net_7201)
	);

	bfr new_net_7203_bfr_before (
		.din(new_net_7203),
		.dout(new_net_7202)
	);

	bfr new_net_7204_bfr_before (
		.din(new_net_7204),
		.dout(new_net_7203)
	);

	bfr new_net_7205_bfr_before (
		.din(new_net_7205),
		.dout(new_net_7204)
	);

	bfr new_net_7206_bfr_before (
		.din(new_net_7206),
		.dout(new_net_7205)
	);

	bfr new_net_7207_bfr_before (
		.din(new_net_7207),
		.dout(new_net_7206)
	);

	bfr new_net_7208_bfr_before (
		.din(new_net_7208),
		.dout(new_net_7207)
	);

	bfr new_net_7209_bfr_before (
		.din(new_net_7209),
		.dout(new_net_7208)
	);

	bfr new_net_7210_bfr_before (
		.din(new_net_7210),
		.dout(new_net_7209)
	);

	bfr new_net_7211_bfr_before (
		.din(new_net_7211),
		.dout(new_net_7210)
	);

	bfr new_net_7212_bfr_before (
		.din(new_net_7212),
		.dout(new_net_7211)
	);

	bfr new_net_7213_bfr_before (
		.din(new_net_7213),
		.dout(new_net_7212)
	);

	bfr new_net_7214_bfr_before (
		.din(new_net_7214),
		.dout(new_net_7213)
	);

	bfr new_net_7215_bfr_before (
		.din(new_net_7215),
		.dout(new_net_7214)
	);

	bfr new_net_7216_bfr_before (
		.din(new_net_7216),
		.dout(new_net_7215)
	);

	bfr new_net_7217_bfr_before (
		.din(new_net_7217),
		.dout(new_net_7216)
	);

	bfr new_net_7218_bfr_before (
		.din(new_net_7218),
		.dout(new_net_7217)
	);

	bfr new_net_7219_bfr_before (
		.din(new_net_7219),
		.dout(new_net_7218)
	);

	bfr new_net_7220_bfr_before (
		.din(new_net_7220),
		.dout(new_net_7219)
	);

	bfr new_net_7221_bfr_before (
		.din(new_net_7221),
		.dout(new_net_7220)
	);

	bfr new_net_7222_bfr_before (
		.din(new_net_7222),
		.dout(new_net_7221)
	);

	spl2 new_net_2028_v_fanout (
		.a(new_net_2028),
		.b(new_net_7222),
		.c(new_net_1340)
	);

	spl4L new_net_2003_v_fanout (
		.a(new_net_2003),
		.b(new_net_247),
		.c(new_net_237),
		.d(new_net_256),
		.e(new_net_232)
	);

	spl4L new_net_2017_v_fanout (
		.a(new_net_2017),
		.b(new_net_205),
		.c(new_net_226),
		.d(new_net_277),
		.e(new_net_235)
	);

	spl4L new_net_2002_v_fanout (
		.a(new_net_2002),
		.b(new_net_142),
		.c(new_net_137),
		.d(new_net_163),
		.e(new_net_129)
	);

	bfr new_net_7223_bfr_before (
		.din(new_net_7223),
		.dout(N567)
	);

	bfr new_net_7224_bfr_before (
		.din(new_net_7224),
		.dout(new_net_7223)
	);

	bfr new_net_7225_bfr_before (
		.din(new_net_7225),
		.dout(new_net_7224)
	);

	bfr new_net_7226_bfr_before (
		.din(new_net_7226),
		.dout(new_net_7225)
	);

	bfr new_net_7227_bfr_before (
		.din(new_net_7227),
		.dout(new_net_7226)
	);

	bfr new_net_7228_bfr_before (
		.din(new_net_7228),
		.dout(new_net_7227)
	);

	bfr new_net_7229_bfr_before (
		.din(new_net_7229),
		.dout(new_net_7228)
	);

	bfr new_net_7230_bfr_before (
		.din(new_net_7230),
		.dout(new_net_7229)
	);

	bfr new_net_7231_bfr_before (
		.din(new_net_7231),
		.dout(new_net_7230)
	);

	bfr new_net_7232_bfr_before (
		.din(new_net_7232),
		.dout(new_net_7231)
	);

	bfr new_net_7233_bfr_before (
		.din(new_net_7233),
		.dout(new_net_7232)
	);

	bfr new_net_7234_bfr_before (
		.din(new_net_7234),
		.dout(new_net_7233)
	);

	bfr new_net_7235_bfr_before (
		.din(new_net_7235),
		.dout(new_net_7234)
	);

	bfr new_net_7236_bfr_before (
		.din(new_net_7236),
		.dout(new_net_7235)
	);

	bfr new_net_7237_bfr_before (
		.din(new_net_7237),
		.dout(new_net_7236)
	);

	bfr new_net_7238_bfr_before (
		.din(new_net_7238),
		.dout(new_net_7237)
	);

	bfr new_net_7239_bfr_before (
		.din(new_net_7239),
		.dout(new_net_7238)
	);

	bfr new_net_7240_bfr_before (
		.din(new_net_7240),
		.dout(new_net_7239)
	);

	bfr new_net_7241_bfr_before (
		.din(new_net_7241),
		.dout(new_net_7240)
	);

	bfr new_net_7242_bfr_before (
		.din(new_net_7242),
		.dout(new_net_7241)
	);

	bfr new_net_7243_bfr_before (
		.din(new_net_7243),
		.dout(new_net_7242)
	);

	bfr new_net_7244_bfr_before (
		.din(new_net_7244),
		.dout(new_net_7243)
	);

	bfr new_net_7245_bfr_before (
		.din(new_net_7245),
		.dout(new_net_7244)
	);

	bfr new_net_7246_bfr_before (
		.din(new_net_7246),
		.dout(new_net_7245)
	);

	bfr new_net_7247_bfr_before (
		.din(new_net_7247),
		.dout(new_net_7246)
	);

	bfr new_net_7248_bfr_before (
		.din(new_net_7248),
		.dout(new_net_7247)
	);

	bfr new_net_7249_bfr_before (
		.din(new_net_7249),
		.dout(new_net_7248)
	);

	bfr new_net_7250_bfr_before (
		.din(new_net_7250),
		.dout(new_net_7249)
	);

	bfr new_net_7251_bfr_before (
		.din(new_net_7251),
		.dout(new_net_7250)
	);

	bfr new_net_7252_bfr_before (
		.din(new_net_7252),
		.dout(new_net_7251)
	);

	bfr new_net_7253_bfr_before (
		.din(new_net_7253),
		.dout(new_net_7252)
	);

	bfr new_net_7254_bfr_before (
		.din(new_net_7254),
		.dout(new_net_7253)
	);

	bfr new_net_7255_bfr_before (
		.din(new_net_7255),
		.dout(new_net_7254)
	);

	bfr new_net_7256_bfr_before (
		.din(new_net_7256),
		.dout(new_net_7255)
	);

	bfr new_net_7257_bfr_before (
		.din(new_net_7257),
		.dout(new_net_7256)
	);

	bfr new_net_7258_bfr_before (
		.din(new_net_7258),
		.dout(new_net_7257)
	);

	bfr new_net_7259_bfr_before (
		.din(new_net_7259),
		.dout(new_net_7258)
	);

	bfr new_net_7260_bfr_before (
		.din(new_net_7260),
		.dout(new_net_7259)
	);

	bfr new_net_7261_bfr_before (
		.din(new_net_7261),
		.dout(new_net_7260)
	);

	bfr new_net_7262_bfr_before (
		.din(new_net_7262),
		.dout(new_net_7261)
	);

	bfr new_net_7263_bfr_before (
		.din(new_net_7263),
		.dout(new_net_7262)
	);

	bfr new_net_7264_bfr_before (
		.din(new_net_7264),
		.dout(new_net_7263)
	);

	bfr new_net_7265_bfr_before (
		.din(new_net_7265),
		.dout(new_net_7264)
	);

	bfr new_net_7266_bfr_before (
		.din(new_net_7266),
		.dout(new_net_7265)
	);

	bfr new_net_7267_bfr_before (
		.din(new_net_7267),
		.dout(new_net_7266)
	);

	bfr new_net_7268_bfr_before (
		.din(new_net_7268),
		.dout(new_net_7267)
	);

	bfr new_net_7269_bfr_before (
		.din(new_net_7269),
		.dout(new_net_7268)
	);

	bfr new_net_7270_bfr_before (
		.din(new_net_7270),
		.dout(new_net_7269)
	);

	bfr new_net_7271_bfr_before (
		.din(new_net_7271),
		.dout(new_net_7270)
	);

	bfr new_net_7272_bfr_before (
		.din(new_net_7272),
		.dout(new_net_7271)
	);

	bfr new_net_7273_bfr_before (
		.din(new_net_7273),
		.dout(new_net_7272)
	);

	bfr new_net_7274_bfr_before (
		.din(new_net_7274),
		.dout(new_net_7273)
	);

	bfr new_net_7275_bfr_before (
		.din(new_net_7275),
		.dout(new_net_7274)
	);

	bfr new_net_7276_bfr_before (
		.din(new_net_7276),
		.dout(new_net_7275)
	);

	bfr new_net_7277_bfr_before (
		.din(new_net_7277),
		.dout(new_net_7276)
	);

	bfr new_net_7278_bfr_before (
		.din(new_net_7278),
		.dout(new_net_7277)
	);

	bfr new_net_7279_bfr_before (
		.din(new_net_7279),
		.dout(new_net_7278)
	);

	bfr new_net_7280_bfr_before (
		.din(new_net_7280),
		.dout(new_net_7279)
	);

	bfr new_net_7281_bfr_before (
		.din(new_net_7281),
		.dout(new_net_7280)
	);

	bfr new_net_7282_bfr_before (
		.din(new_net_7282),
		.dout(new_net_7281)
	);

	bfr new_net_7283_bfr_before (
		.din(new_net_7283),
		.dout(new_net_7282)
	);

	bfr new_net_7284_bfr_before (
		.din(new_net_7284),
		.dout(new_net_7283)
	);

	spl2 new_net_2050_v_fanout (
		.a(new_net_2050),
		.b(new_net_7284),
		.c(new_net_519)
	);

	spl4L new_net_1996_v_fanout (
		.a(new_net_1996),
		.b(new_net_155),
		.c(new_net_257),
		.d(new_net_176),
		.e(new_net_189)
	);

	bfr new_net_7285_bfr_before (
		.din(new_net_7285),
		.dout(N573)
	);

	bfr new_net_7286_bfr_before (
		.din(new_net_7286),
		.dout(new_net_7285)
	);

	bfr new_net_7287_bfr_before (
		.din(new_net_7287),
		.dout(new_net_7286)
	);

	bfr new_net_7288_bfr_before (
		.din(new_net_7288),
		.dout(new_net_7287)
	);

	bfr new_net_7289_bfr_before (
		.din(new_net_7289),
		.dout(new_net_7288)
	);

	bfr new_net_7290_bfr_before (
		.din(new_net_7290),
		.dout(new_net_7289)
	);

	bfr new_net_7291_bfr_before (
		.din(new_net_7291),
		.dout(new_net_7290)
	);

	bfr new_net_7292_bfr_before (
		.din(new_net_7292),
		.dout(new_net_7291)
	);

	bfr new_net_7293_bfr_before (
		.din(new_net_7293),
		.dout(new_net_7292)
	);

	bfr new_net_7294_bfr_before (
		.din(new_net_7294),
		.dout(new_net_7293)
	);

	bfr new_net_7295_bfr_before (
		.din(new_net_7295),
		.dout(new_net_7294)
	);

	bfr new_net_7296_bfr_before (
		.din(new_net_7296),
		.dout(new_net_7295)
	);

	bfr new_net_7297_bfr_before (
		.din(new_net_7297),
		.dout(new_net_7296)
	);

	bfr new_net_7298_bfr_before (
		.din(new_net_7298),
		.dout(new_net_7297)
	);

	bfr new_net_7299_bfr_before (
		.din(new_net_7299),
		.dout(new_net_7298)
	);

	bfr new_net_7300_bfr_before (
		.din(new_net_7300),
		.dout(new_net_7299)
	);

	bfr new_net_7301_bfr_before (
		.din(new_net_7301),
		.dout(new_net_7300)
	);

	bfr new_net_7302_bfr_before (
		.din(new_net_7302),
		.dout(new_net_7301)
	);

	bfr new_net_7303_bfr_before (
		.din(new_net_7303),
		.dout(new_net_7302)
	);

	bfr new_net_7304_bfr_before (
		.din(new_net_7304),
		.dout(new_net_7303)
	);

	bfr new_net_7305_bfr_before (
		.din(new_net_7305),
		.dout(new_net_7304)
	);

	bfr new_net_7306_bfr_before (
		.din(new_net_7306),
		.dout(new_net_7305)
	);

	bfr new_net_7307_bfr_before (
		.din(new_net_7307),
		.dout(new_net_7306)
	);

	bfr new_net_7308_bfr_before (
		.din(new_net_7308),
		.dout(new_net_7307)
	);

	bfr new_net_7309_bfr_before (
		.din(new_net_7309),
		.dout(new_net_7308)
	);

	bfr new_net_7310_bfr_before (
		.din(new_net_7310),
		.dout(new_net_7309)
	);

	bfr new_net_7311_bfr_before (
		.din(new_net_7311),
		.dout(new_net_7310)
	);

	bfr new_net_7312_bfr_before (
		.din(new_net_7312),
		.dout(new_net_7311)
	);

	bfr new_net_7313_bfr_before (
		.din(new_net_7313),
		.dout(new_net_7312)
	);

	bfr new_net_7314_bfr_before (
		.din(new_net_7314),
		.dout(new_net_7313)
	);

	bfr new_net_7315_bfr_before (
		.din(new_net_7315),
		.dout(new_net_7314)
	);

	bfr new_net_7316_bfr_before (
		.din(new_net_7316),
		.dout(new_net_7315)
	);

	bfr new_net_7317_bfr_before (
		.din(new_net_7317),
		.dout(new_net_7316)
	);

	bfr new_net_7318_bfr_before (
		.din(new_net_7318),
		.dout(new_net_7317)
	);

	bfr new_net_7319_bfr_before (
		.din(new_net_7319),
		.dout(new_net_7318)
	);

	bfr new_net_7320_bfr_before (
		.din(new_net_7320),
		.dout(new_net_7319)
	);

	bfr new_net_7321_bfr_before (
		.din(new_net_7321),
		.dout(new_net_7320)
	);

	bfr new_net_7322_bfr_before (
		.din(new_net_7322),
		.dout(new_net_7321)
	);

	bfr new_net_7323_bfr_before (
		.din(new_net_7323),
		.dout(new_net_7322)
	);

	bfr new_net_7324_bfr_before (
		.din(new_net_7324),
		.dout(new_net_7323)
	);

	bfr new_net_7325_bfr_before (
		.din(new_net_7325),
		.dout(new_net_7324)
	);

	bfr new_net_7326_bfr_before (
		.din(new_net_7326),
		.dout(new_net_7325)
	);

	bfr new_net_7327_bfr_before (
		.din(new_net_7327),
		.dout(new_net_7326)
	);

	bfr new_net_7328_bfr_before (
		.din(new_net_7328),
		.dout(new_net_7327)
	);

	bfr new_net_7329_bfr_before (
		.din(new_net_7329),
		.dout(new_net_7328)
	);

	bfr new_net_7330_bfr_before (
		.din(new_net_7330),
		.dout(new_net_7329)
	);

	bfr new_net_7331_bfr_before (
		.din(new_net_7331),
		.dout(new_net_7330)
	);

	bfr new_net_7332_bfr_before (
		.din(new_net_7332),
		.dout(new_net_7331)
	);

	bfr new_net_7333_bfr_before (
		.din(new_net_7333),
		.dout(new_net_7332)
	);

	bfr new_net_7334_bfr_before (
		.din(new_net_7334),
		.dout(new_net_7333)
	);

	bfr new_net_7335_bfr_before (
		.din(new_net_7335),
		.dout(new_net_7334)
	);

	bfr new_net_7336_bfr_before (
		.din(new_net_7336),
		.dout(new_net_7335)
	);

	bfr new_net_7337_bfr_before (
		.din(new_net_7337),
		.dout(new_net_7336)
	);

	bfr new_net_7338_bfr_before (
		.din(new_net_7338),
		.dout(new_net_7337)
	);

	bfr new_net_7339_bfr_before (
		.din(new_net_7339),
		.dout(new_net_7338)
	);

	bfr new_net_7340_bfr_before (
		.din(new_net_7340),
		.dout(new_net_7339)
	);

	bfr new_net_7341_bfr_before (
		.din(new_net_7341),
		.dout(new_net_7340)
	);

	bfr new_net_7342_bfr_before (
		.din(new_net_7342),
		.dout(new_net_7341)
	);

	bfr new_net_7343_bfr_before (
		.din(new_net_7343),
		.dout(new_net_7342)
	);

	bfr new_net_7344_bfr_before (
		.din(new_net_7344),
		.dout(new_net_7343)
	);

	bfr new_net_7345_bfr_before (
		.din(new_net_7345),
		.dout(new_net_7344)
	);

	bfr new_net_7346_bfr_before (
		.din(new_net_7346),
		.dout(new_net_7345)
	);

	spl2 new_net_2053_v_fanout (
		.a(new_net_2053),
		.b(new_net_7346),
		.c(new_net_849)
	);

	spl4L new_net_1965_v_fanout (
		.a(new_net_1965),
		.b(new_net_164),
		.c(new_net_143),
		.d(new_net_130),
		.e(new_net_122)
	);

	spl2 new_net_2056_v_fanout (
		.a(new_net_2056),
		.b(new_net_1084),
		.c(new_net_1086)
	);

	spl4L new_net_2000_v_fanout (
		.a(new_net_2000),
		.b(new_net_271),
		.c(new_net_198),
		.d(new_net_150),
		.e(new_net_229)
	);

	spl4L new_net_1973_v_fanout (
		.a(new_net_1973),
		.b(new_net_133),
		.c(new_net_138),
		.d(new_net_180),
		.e(new_net_125)
	);

	spl4L new_net_1975_v_fanout (
		.a(new_net_1975),
		.b(new_net_243),
		.c(new_net_285),
		.d(new_net_275),
		.e(new_net_233)
	);

	spl4L new_net_1987_v_fanout (
		.a(new_net_1987),
		.b(new_net_194),
		.c(new_net_123),
		.d(new_net_173),
		.e(new_net_152)
	);

	spl4L new_net_1966_v_fanout (
		.a(new_net_1966),
		.b(new_net_206),
		.c(new_net_193),
		.d(new_net_172),
		.e(new_net_185)
	);

	spl4L new_net_1994_v_fanout (
		.a(new_net_1994),
		.b(new_net_126),
		.c(new_net_134),
		.d(new_net_139),
		.e(new_net_272)
	);

	bfr new_net_7347_bfr_after (
		.din(new_net_12),
		.dout(new_net_7347)
	);

	bfr new_net_7348_bfr_after (
		.din(new_net_7347),
		.dout(new_net_7348)
	);

	bfr new_net_7349_bfr_after (
		.din(new_net_7348),
		.dout(new_net_7349)
	);

	bfr new_net_7350_bfr_after (
		.din(new_net_7349),
		.dout(new_net_7350)
	);

	bfr new_net_7351_bfr_after (
		.din(new_net_7350),
		.dout(new_net_7351)
	);

	bfr new_net_7352_bfr_after (
		.din(new_net_7351),
		.dout(new_net_7352)
	);

	bfr new_net_7353_bfr_after (
		.din(new_net_7352),
		.dout(new_net_7353)
	);

	bfr new_net_7354_bfr_after (
		.din(new_net_7353),
		.dout(new_net_7354)
	);

	bfr new_net_7355_bfr_after (
		.din(new_net_7354),
		.dout(new_net_7355)
	);

	bfr new_net_7356_bfr_after (
		.din(new_net_7355),
		.dout(new_net_7356)
	);

	bfr new_net_7357_bfr_after (
		.din(new_net_7356),
		.dout(new_net_7357)
	);

	bfr new_net_7358_bfr_after (
		.din(new_net_7357),
		.dout(new_net_7358)
	);

	bfr new_net_7359_bfr_after (
		.din(new_net_7358),
		.dout(new_net_7359)
	);

	bfr new_net_7360_bfr_after (
		.din(new_net_7359),
		.dout(new_net_7360)
	);

	bfr new_net_7361_bfr_after (
		.din(new_net_7360),
		.dout(new_net_7361)
	);

	bfr new_net_7362_bfr_after (
		.din(new_net_7361),
		.dout(new_net_7362)
	);

	bfr new_net_7363_bfr_after (
		.din(new_net_7362),
		.dout(new_net_7363)
	);

	bfr new_net_7364_bfr_after (
		.din(new_net_7363),
		.dout(new_net_7364)
	);

	bfr new_net_7365_bfr_after (
		.din(new_net_7364),
		.dout(new_net_7365)
	);

	bfr new_net_7366_bfr_after (
		.din(new_net_7365),
		.dout(new_net_7366)
	);

	bfr new_net_7367_bfr_after (
		.din(new_net_7366),
		.dout(new_net_7367)
	);

	bfr new_net_7368_bfr_after (
		.din(new_net_7367),
		.dout(new_net_7368)
	);

	bfr new_net_7369_bfr_after (
		.din(new_net_7368),
		.dout(new_net_7369)
	);

	bfr new_net_7370_bfr_after (
		.din(new_net_7369),
		.dout(new_net_7370)
	);

	bfr new_net_7371_bfr_after (
		.din(new_net_7370),
		.dout(new_net_7371)
	);

	bfr new_net_7372_bfr_after (
		.din(new_net_7371),
		.dout(new_net_7372)
	);

	bfr new_net_7373_bfr_after (
		.din(new_net_7372),
		.dout(new_net_7373)
	);

	bfr new_net_7374_bfr_after (
		.din(new_net_7373),
		.dout(new_net_7374)
	);

	bfr new_net_7375_bfr_after (
		.din(new_net_7374),
		.dout(new_net_7375)
	);

	bfr new_net_7376_bfr_after (
		.din(new_net_7375),
		.dout(new_net_7376)
	);

	bfr new_net_7377_bfr_after (
		.din(new_net_7376),
		.dout(new_net_7377)
	);

	bfr new_net_7378_bfr_after (
		.din(new_net_7377),
		.dout(new_net_7378)
	);

	bfr new_net_7379_bfr_after (
		.din(new_net_7378),
		.dout(new_net_7379)
	);

	bfr new_net_7380_bfr_after (
		.din(new_net_7379),
		.dout(new_net_7380)
	);

	bfr new_net_7381_bfr_after (
		.din(new_net_7380),
		.dout(new_net_7381)
	);

	bfr new_net_7382_bfr_after (
		.din(new_net_7381),
		.dout(new_net_7382)
	);

	bfr new_net_7383_bfr_after (
		.din(new_net_7382),
		.dout(new_net_7383)
	);

	bfr new_net_7384_bfr_after (
		.din(new_net_7383),
		.dout(new_net_7384)
	);

	bfr new_net_7385_bfr_after (
		.din(new_net_7384),
		.dout(new_net_7385)
	);

	bfr new_net_7386_bfr_after (
		.din(new_net_7385),
		.dout(new_net_7386)
	);

	bfr new_net_7387_bfr_after (
		.din(new_net_7386),
		.dout(new_net_7387)
	);

	bfr new_net_7388_bfr_after (
		.din(new_net_7387),
		.dout(new_net_7388)
	);

	bfr new_net_7389_bfr_after (
		.din(new_net_7388),
		.dout(new_net_7389)
	);

	bfr new_net_7390_bfr_after (
		.din(new_net_7389),
		.dout(new_net_7390)
	);

	bfr new_net_7391_bfr_after (
		.din(new_net_7390),
		.dout(new_net_7391)
	);

	bfr new_net_7392_bfr_after (
		.din(new_net_7391),
		.dout(new_net_7392)
	);

	bfr new_net_7393_bfr_after (
		.din(new_net_7392),
		.dout(new_net_7393)
	);

	bfr new_net_7394_bfr_after (
		.din(new_net_7393),
		.dout(new_net_7394)
	);

	bfr new_net_7395_bfr_after (
		.din(new_net_7394),
		.dout(new_net_7395)
	);

	bfr new_net_7396_bfr_after (
		.din(new_net_7395),
		.dout(new_net_7396)
	);

	bfr new_net_7397_bfr_after (
		.din(new_net_7396),
		.dout(new_net_7397)
	);

	bfr new_net_7398_bfr_after (
		.din(new_net_7397),
		.dout(new_net_7398)
	);

	bfr new_net_7399_bfr_after (
		.din(new_net_7398),
		.dout(new_net_7399)
	);

	bfr new_net_7400_bfr_after (
		.din(new_net_7399),
		.dout(new_net_7400)
	);

	bfr new_net_7401_bfr_after (
		.din(new_net_7400),
		.dout(new_net_7401)
	);

	bfr new_net_7402_bfr_after (
		.din(new_net_7401),
		.dout(new_net_7402)
	);

	bfr new_net_7403_bfr_after (
		.din(new_net_7402),
		.dout(new_net_7403)
	);

	bfr new_net_7404_bfr_after (
		.din(new_net_7403),
		.dout(new_net_7404)
	);

	bfr new_net_7405_bfr_after (
		.din(new_net_7404),
		.dout(new_net_7405)
	);

	bfr new_net_7406_bfr_after (
		.din(new_net_7405),
		.dout(new_net_7406)
	);

	bfr new_net_7407_bfr_after (
		.din(new_net_7406),
		.dout(new_net_7407)
	);

	bfr new_net_7408_bfr_after (
		.din(new_net_7407),
		.dout(new_net_7408)
	);

	spl2 new_net_12_v_fanout (
		.a(new_net_7408),
		.b(N1489),
		.c(N1113)
	);

	spl4L new_net_2001_v_fanout (
		.a(new_net_2001),
		.b(new_net_179),
		.c(new_net_158),
		.d(new_net_192),
		.e(new_net_171)
	);

	spl4L new_net_1979_v_fanout (
		.a(new_net_1979),
		.b(new_net_220),
		.c(new_net_241),
		.d(new_net_251),
		.e(new_net_260)
	);

	spl4L new_net_2006_v_fanout (
		.a(new_net_2006),
		.b(new_net_124),
		.c(new_net_148),
		.d(new_net_178),
		.e(new_net_274)
	);

	bfr new_net_7409_bfr_before (
		.din(new_net_7409),
		.dout(N551)
	);

	bfr new_net_7410_bfr_before (
		.din(new_net_7410),
		.dout(new_net_7409)
	);

	bfr new_net_7411_bfr_before (
		.din(new_net_7411),
		.dout(new_net_7410)
	);

	bfr new_net_7412_bfr_before (
		.din(new_net_7412),
		.dout(new_net_7411)
	);

	bfr new_net_7413_bfr_before (
		.din(new_net_7413),
		.dout(new_net_7412)
	);

	bfr new_net_7414_bfr_before (
		.din(new_net_7414),
		.dout(new_net_7413)
	);

	bfr new_net_7415_bfr_before (
		.din(new_net_7415),
		.dout(new_net_7414)
	);

	bfr new_net_7416_bfr_before (
		.din(new_net_7416),
		.dout(new_net_7415)
	);

	bfr new_net_7417_bfr_before (
		.din(new_net_7417),
		.dout(new_net_7416)
	);

	bfr new_net_7418_bfr_before (
		.din(new_net_7418),
		.dout(new_net_7417)
	);

	bfr new_net_7419_bfr_before (
		.din(new_net_7419),
		.dout(new_net_7418)
	);

	bfr new_net_7420_bfr_before (
		.din(new_net_7420),
		.dout(new_net_7419)
	);

	bfr new_net_7421_bfr_before (
		.din(new_net_7421),
		.dout(new_net_7420)
	);

	bfr new_net_7422_bfr_before (
		.din(new_net_7422),
		.dout(new_net_7421)
	);

	bfr new_net_7423_bfr_before (
		.din(new_net_7423),
		.dout(new_net_7422)
	);

	bfr new_net_7424_bfr_before (
		.din(new_net_7424),
		.dout(new_net_7423)
	);

	bfr new_net_7425_bfr_before (
		.din(new_net_7425),
		.dout(new_net_7424)
	);

	bfr new_net_7426_bfr_before (
		.din(new_net_7426),
		.dout(new_net_7425)
	);

	bfr new_net_7427_bfr_before (
		.din(new_net_7427),
		.dout(new_net_7426)
	);

	bfr new_net_7428_bfr_before (
		.din(new_net_7428),
		.dout(new_net_7427)
	);

	bfr new_net_7429_bfr_before (
		.din(new_net_7429),
		.dout(new_net_7428)
	);

	bfr new_net_7430_bfr_before (
		.din(new_net_7430),
		.dout(new_net_7429)
	);

	bfr new_net_7431_bfr_before (
		.din(new_net_7431),
		.dout(new_net_7430)
	);

	bfr new_net_7432_bfr_before (
		.din(new_net_7432),
		.dout(new_net_7431)
	);

	bfr new_net_7433_bfr_before (
		.din(new_net_7433),
		.dout(new_net_7432)
	);

	bfr new_net_7434_bfr_before (
		.din(new_net_7434),
		.dout(new_net_7433)
	);

	bfr new_net_7435_bfr_before (
		.din(new_net_7435),
		.dout(new_net_7434)
	);

	bfr new_net_7436_bfr_before (
		.din(new_net_7436),
		.dout(new_net_7435)
	);

	bfr new_net_7437_bfr_before (
		.din(new_net_7437),
		.dout(new_net_7436)
	);

	bfr new_net_7438_bfr_before (
		.din(new_net_7438),
		.dout(new_net_7437)
	);

	bfr new_net_7439_bfr_before (
		.din(new_net_7439),
		.dout(new_net_7438)
	);

	bfr new_net_7440_bfr_before (
		.din(new_net_7440),
		.dout(new_net_7439)
	);

	bfr new_net_7441_bfr_before (
		.din(new_net_7441),
		.dout(new_net_7440)
	);

	bfr new_net_7442_bfr_before (
		.din(new_net_7442),
		.dout(new_net_7441)
	);

	bfr new_net_7443_bfr_before (
		.din(new_net_7443),
		.dout(new_net_7442)
	);

	bfr new_net_7444_bfr_before (
		.din(new_net_7444),
		.dout(new_net_7443)
	);

	bfr new_net_7445_bfr_before (
		.din(new_net_7445),
		.dout(new_net_7444)
	);

	bfr new_net_7446_bfr_before (
		.din(new_net_7446),
		.dout(new_net_7445)
	);

	bfr new_net_7447_bfr_before (
		.din(new_net_7447),
		.dout(new_net_7446)
	);

	bfr new_net_7448_bfr_before (
		.din(new_net_7448),
		.dout(new_net_7447)
	);

	bfr new_net_7449_bfr_before (
		.din(new_net_7449),
		.dout(new_net_7448)
	);

	bfr new_net_7450_bfr_before (
		.din(new_net_7450),
		.dout(new_net_7449)
	);

	bfr new_net_7451_bfr_before (
		.din(new_net_7451),
		.dout(new_net_7450)
	);

	bfr new_net_7452_bfr_before (
		.din(new_net_7452),
		.dout(new_net_7451)
	);

	bfr new_net_7453_bfr_before (
		.din(new_net_7453),
		.dout(new_net_7452)
	);

	bfr new_net_7454_bfr_before (
		.din(new_net_7454),
		.dout(new_net_7453)
	);

	bfr new_net_7455_bfr_before (
		.din(new_net_7455),
		.dout(new_net_7454)
	);

	bfr new_net_7456_bfr_before (
		.din(new_net_7456),
		.dout(new_net_7455)
	);

	bfr new_net_7457_bfr_before (
		.din(new_net_7457),
		.dout(new_net_7456)
	);

	bfr new_net_7458_bfr_before (
		.din(new_net_7458),
		.dout(new_net_7457)
	);

	bfr new_net_7459_bfr_before (
		.din(new_net_7459),
		.dout(new_net_7458)
	);

	bfr new_net_7460_bfr_before (
		.din(new_net_7460),
		.dout(new_net_7459)
	);

	bfr new_net_7461_bfr_before (
		.din(new_net_7461),
		.dout(new_net_7460)
	);

	bfr new_net_7462_bfr_before (
		.din(new_net_7462),
		.dout(new_net_7461)
	);

	bfr new_net_7463_bfr_before (
		.din(new_net_7463),
		.dout(new_net_7462)
	);

	bfr new_net_7464_bfr_before (
		.din(new_net_7464),
		.dout(new_net_7463)
	);

	bfr new_net_7465_bfr_before (
		.din(new_net_7465),
		.dout(new_net_7464)
	);

	bfr new_net_7466_bfr_before (
		.din(new_net_7466),
		.dout(new_net_7465)
	);

	bfr new_net_7467_bfr_before (
		.din(new_net_7467),
		.dout(new_net_7466)
	);

	bfr new_net_7468_bfr_before (
		.din(new_net_7468),
		.dout(new_net_7467)
	);

	bfr new_net_7469_bfr_before (
		.din(new_net_7469),
		.dout(new_net_7468)
	);

	bfr new_net_7470_bfr_before (
		.din(new_net_7470),
		.dout(new_net_7469)
	);

	spl2 new_net_2043_v_fanout (
		.a(new_net_2043),
		.b(new_net_7470),
		.c(new_net_1349)
	);

	spl4L new_net_1989_v_fanout (
		.a(new_net_1989),
		.b(new_net_144),
		.c(new_net_186),
		.d(new_net_165),
		.e(new_net_131)
	);

	spl4L new_net_2012_v_fanout (
		.a(new_net_2012),
		.b(new_net_196),
		.c(new_net_263),
		.d(new_net_169),
		.e(new_net_269)
	);

	bfr new_net_7471_bfr_before (
		.din(new_net_7471),
		.dout(N559)
	);

	bfr new_net_7472_bfr_before (
		.din(new_net_7472),
		.dout(new_net_7471)
	);

	bfr new_net_7473_bfr_before (
		.din(new_net_7473),
		.dout(new_net_7472)
	);

	bfr new_net_7474_bfr_before (
		.din(new_net_7474),
		.dout(new_net_7473)
	);

	bfr new_net_7475_bfr_before (
		.din(new_net_7475),
		.dout(new_net_7474)
	);

	bfr new_net_7476_bfr_before (
		.din(new_net_7476),
		.dout(new_net_7475)
	);

	bfr new_net_7477_bfr_before (
		.din(new_net_7477),
		.dout(new_net_7476)
	);

	bfr new_net_7478_bfr_before (
		.din(new_net_7478),
		.dout(new_net_7477)
	);

	bfr new_net_7479_bfr_before (
		.din(new_net_7479),
		.dout(new_net_7478)
	);

	bfr new_net_7480_bfr_before (
		.din(new_net_7480),
		.dout(new_net_7479)
	);

	bfr new_net_7481_bfr_before (
		.din(new_net_7481),
		.dout(new_net_7480)
	);

	bfr new_net_7482_bfr_before (
		.din(new_net_7482),
		.dout(new_net_7481)
	);

	bfr new_net_7483_bfr_before (
		.din(new_net_7483),
		.dout(new_net_7482)
	);

	bfr new_net_7484_bfr_before (
		.din(new_net_7484),
		.dout(new_net_7483)
	);

	bfr new_net_7485_bfr_before (
		.din(new_net_7485),
		.dout(new_net_7484)
	);

	bfr new_net_7486_bfr_before (
		.din(new_net_7486),
		.dout(new_net_7485)
	);

	bfr new_net_7487_bfr_before (
		.din(new_net_7487),
		.dout(new_net_7486)
	);

	bfr new_net_7488_bfr_before (
		.din(new_net_7488),
		.dout(new_net_7487)
	);

	bfr new_net_7489_bfr_before (
		.din(new_net_7489),
		.dout(new_net_7488)
	);

	bfr new_net_7490_bfr_before (
		.din(new_net_7490),
		.dout(new_net_7489)
	);

	bfr new_net_7491_bfr_before (
		.din(new_net_7491),
		.dout(new_net_7490)
	);

	bfr new_net_7492_bfr_before (
		.din(new_net_7492),
		.dout(new_net_7491)
	);

	bfr new_net_7493_bfr_before (
		.din(new_net_7493),
		.dout(new_net_7492)
	);

	bfr new_net_7494_bfr_before (
		.din(new_net_7494),
		.dout(new_net_7493)
	);

	bfr new_net_7495_bfr_before (
		.din(new_net_7495),
		.dout(new_net_7494)
	);

	bfr new_net_7496_bfr_before (
		.din(new_net_7496),
		.dout(new_net_7495)
	);

	bfr new_net_7497_bfr_before (
		.din(new_net_7497),
		.dout(new_net_7496)
	);

	bfr new_net_7498_bfr_before (
		.din(new_net_7498),
		.dout(new_net_7497)
	);

	bfr new_net_7499_bfr_before (
		.din(new_net_7499),
		.dout(new_net_7498)
	);

	bfr new_net_7500_bfr_before (
		.din(new_net_7500),
		.dout(new_net_7499)
	);

	bfr new_net_7501_bfr_before (
		.din(new_net_7501),
		.dout(new_net_7500)
	);

	bfr new_net_7502_bfr_before (
		.din(new_net_7502),
		.dout(new_net_7501)
	);

	bfr new_net_7503_bfr_before (
		.din(new_net_7503),
		.dout(new_net_7502)
	);

	bfr new_net_7504_bfr_before (
		.din(new_net_7504),
		.dout(new_net_7503)
	);

	bfr new_net_7505_bfr_before (
		.din(new_net_7505),
		.dout(new_net_7504)
	);

	bfr new_net_7506_bfr_before (
		.din(new_net_7506),
		.dout(new_net_7505)
	);

	bfr new_net_7507_bfr_before (
		.din(new_net_7507),
		.dout(new_net_7506)
	);

	bfr new_net_7508_bfr_before (
		.din(new_net_7508),
		.dout(new_net_7507)
	);

	bfr new_net_7509_bfr_before (
		.din(new_net_7509),
		.dout(new_net_7508)
	);

	bfr new_net_7510_bfr_before (
		.din(new_net_7510),
		.dout(new_net_7509)
	);

	bfr new_net_7511_bfr_before (
		.din(new_net_7511),
		.dout(new_net_7510)
	);

	bfr new_net_7512_bfr_before (
		.din(new_net_7512),
		.dout(new_net_7511)
	);

	bfr new_net_7513_bfr_before (
		.din(new_net_7513),
		.dout(new_net_7512)
	);

	bfr new_net_7514_bfr_before (
		.din(new_net_7514),
		.dout(new_net_7513)
	);

	bfr new_net_7515_bfr_before (
		.din(new_net_7515),
		.dout(new_net_7514)
	);

	bfr new_net_7516_bfr_before (
		.din(new_net_7516),
		.dout(new_net_7515)
	);

	bfr new_net_7517_bfr_before (
		.din(new_net_7517),
		.dout(new_net_7516)
	);

	bfr new_net_7518_bfr_before (
		.din(new_net_7518),
		.dout(new_net_7517)
	);

	bfr new_net_7519_bfr_before (
		.din(new_net_7519),
		.dout(new_net_7518)
	);

	bfr new_net_7520_bfr_before (
		.din(new_net_7520),
		.dout(new_net_7519)
	);

	bfr new_net_7521_bfr_before (
		.din(new_net_7521),
		.dout(new_net_7520)
	);

	bfr new_net_7522_bfr_before (
		.din(new_net_7522),
		.dout(new_net_7521)
	);

	bfr new_net_7523_bfr_before (
		.din(new_net_7523),
		.dout(new_net_7522)
	);

	bfr new_net_7524_bfr_before (
		.din(new_net_7524),
		.dout(new_net_7523)
	);

	bfr new_net_7525_bfr_before (
		.din(new_net_7525),
		.dout(new_net_7524)
	);

	bfr new_net_7526_bfr_before (
		.din(new_net_7526),
		.dout(new_net_7525)
	);

	bfr new_net_7527_bfr_before (
		.din(new_net_7527),
		.dout(new_net_7526)
	);

	bfr new_net_7528_bfr_before (
		.din(new_net_7528),
		.dout(new_net_7527)
	);

	bfr new_net_7529_bfr_before (
		.din(new_net_7529),
		.dout(new_net_7528)
	);

	bfr new_net_7530_bfr_before (
		.din(new_net_7530),
		.dout(new_net_7529)
	);

	bfr new_net_7531_bfr_before (
		.din(new_net_7531),
		.dout(new_net_7530)
	);

	bfr new_net_7532_bfr_before (
		.din(new_net_7532),
		.dout(new_net_7531)
	);

	spl2 new_net_2046_v_fanout (
		.a(new_net_2046),
		.b(new_net_7532),
		.c(new_net_1579)
	);

	bfr new_net_7533_bfr_before (
		.din(new_net_7533),
		.dout(new_net_1169)
	);

	bfr new_net_7534_bfr_before (
		.din(new_net_7534),
		.dout(new_net_7533)
	);

	bfr new_net_7535_bfr_before (
		.din(new_net_7535),
		.dout(new_net_7534)
	);

	bfr new_net_7536_bfr_before (
		.din(new_net_7536),
		.dout(new_net_7535)
	);

	spl2 n_0938__v_fanout (
		.a(n_0938_),
		.b(new_net_1170),
		.c(new_net_7536)
	);

	spl4L new_net_1988_v_fanout (
		.a(new_net_1988),
		.b(new_net_1990),
		.c(new_net_1989),
		.d(new_net_1991),
		.e(new_net_1992)
	);

	bfr new_net_7537_bfr_after (
		.din(n_0668_),
		.dout(new_net_7537)
	);

	bfr new_net_7538_bfr_after (
		.din(new_net_7537),
		.dout(new_net_7538)
	);

	bfr new_net_7539_bfr_after (
		.din(new_net_7538),
		.dout(new_net_7539)
	);

	bfr new_net_7540_bfr_after (
		.din(new_net_7539),
		.dout(new_net_7540)
	);

	bfr new_net_7541_bfr_after (
		.din(new_net_7540),
		.dout(new_net_7541)
	);

	bfr new_net_7542_bfr_after (
		.din(new_net_7541),
		.dout(new_net_7542)
	);

	bfr new_net_7543_bfr_after (
		.din(new_net_7542),
		.dout(new_net_7543)
	);

	bfr new_net_7544_bfr_before (
		.din(new_net_7544),
		.dout(new_net_2065)
	);

	bfr new_net_7545_bfr_before (
		.din(new_net_7545),
		.dout(new_net_7544)
	);

	bfr new_net_7546_bfr_before (
		.din(new_net_7546),
		.dout(new_net_7545)
	);

	bfr new_net_7547_bfr_before (
		.din(new_net_7547),
		.dout(new_net_7546)
	);

	bfr new_net_7548_bfr_before (
		.din(new_net_7548),
		.dout(new_net_7547)
	);

	bfr new_net_7549_bfr_before (
		.din(new_net_7549),
		.dout(new_net_7548)
	);

	bfr new_net_7550_bfr_before (
		.din(new_net_7550),
		.dout(new_net_7549)
	);

	bfr new_net_7551_bfr_before (
		.din(new_net_7551),
		.dout(new_net_7550)
	);

	bfr new_net_7552_bfr_before (
		.din(new_net_7552),
		.dout(new_net_7551)
	);

	bfr new_net_7553_bfr_before (
		.din(new_net_7553),
		.dout(new_net_7552)
	);

	bfr new_net_7554_bfr_before (
		.din(new_net_7554),
		.dout(new_net_7553)
	);

	spl2 n_0668__v_fanout (
		.a(new_net_7543),
		.b(new_net_7554),
		.c(new_net_1676)
	);

	bfr new_net_7555_bfr_after (
		.din(n_0670_),
		.dout(new_net_7555)
	);

	bfr new_net_7556_bfr_after (
		.din(new_net_7555),
		.dout(new_net_7556)
	);

	bfr new_net_7557_bfr_after (
		.din(new_net_7556),
		.dout(new_net_7557)
	);

	bfr new_net_7558_bfr_after (
		.din(new_net_7557),
		.dout(new_net_7558)
	);

	bfr new_net_7559_bfr_after (
		.din(new_net_7558),
		.dout(new_net_7559)
	);

	spl2 n_0670__v_fanout (
		.a(new_net_7559),
		.b(new_net_1453),
		.c(new_net_1452)
	);

	bfr new_net_7560_bfr_after (
		.din(n_1321_),
		.dout(new_net_7560)
	);

	bfr new_net_7561_bfr_after (
		.din(new_net_7560),
		.dout(new_net_7561)
	);

	bfr new_net_7562_bfr_after (
		.din(new_net_7561),
		.dout(new_net_7562)
	);

	bfr new_net_7563_bfr_after (
		.din(new_net_7562),
		.dout(new_net_7563)
	);

	bfr new_net_7564_bfr_after (
		.din(new_net_7563),
		.dout(new_net_7564)
	);

	spl2 n_1321__v_fanout (
		.a(new_net_7564),
		.b(new_net_1297),
		.c(new_net_1296)
	);

	bfr new_net_7565_bfr_before (
		.din(new_net_7565),
		.dout(N884)
	);

	bfr new_net_7566_bfr_before (
		.din(new_net_7566),
		.dout(new_net_7565)
	);

	bfr new_net_7567_bfr_before (
		.din(new_net_7567),
		.dout(new_net_7566)
	);

	bfr new_net_7568_bfr_before (
		.din(new_net_7568),
		.dout(new_net_7567)
	);

	bfr new_net_7569_bfr_before (
		.din(new_net_7569),
		.dout(new_net_7568)
	);

	bfr new_net_7570_bfr_before (
		.din(new_net_7570),
		.dout(new_net_7569)
	);

	bfr new_net_7571_bfr_before (
		.din(new_net_7571),
		.dout(new_net_7570)
	);

	bfr new_net_7572_bfr_before (
		.din(new_net_7572),
		.dout(new_net_7571)
	);

	bfr new_net_7573_bfr_before (
		.din(new_net_7573),
		.dout(new_net_7572)
	);

	bfr new_net_7574_bfr_before (
		.din(new_net_7574),
		.dout(new_net_7573)
	);

	bfr new_net_7575_bfr_before (
		.din(new_net_7575),
		.dout(new_net_7574)
	);

	bfr new_net_7576_bfr_before (
		.din(new_net_7576),
		.dout(new_net_7575)
	);

	bfr new_net_7577_bfr_before (
		.din(new_net_7577),
		.dout(new_net_7576)
	);

	bfr new_net_7578_bfr_before (
		.din(new_net_7578),
		.dout(new_net_7577)
	);

	bfr new_net_7579_bfr_before (
		.din(new_net_7579),
		.dout(new_net_7578)
	);

	bfr new_net_7580_bfr_before (
		.din(new_net_7580),
		.dout(new_net_7579)
	);

	bfr new_net_7581_bfr_before (
		.din(new_net_7581),
		.dout(new_net_7580)
	);

	bfr new_net_7582_bfr_before (
		.din(new_net_7582),
		.dout(new_net_7581)
	);

	bfr new_net_7583_bfr_before (
		.din(new_net_7583),
		.dout(new_net_7582)
	);

	bfr new_net_7584_bfr_before (
		.din(new_net_7584),
		.dout(new_net_7583)
	);

	bfr new_net_7585_bfr_before (
		.din(new_net_7585),
		.dout(new_net_7584)
	);

	bfr new_net_7586_bfr_before (
		.din(new_net_7586),
		.dout(new_net_7585)
	);

	bfr new_net_7587_bfr_before (
		.din(new_net_7587),
		.dout(new_net_7586)
	);

	bfr new_net_7588_bfr_before (
		.din(new_net_7588),
		.dout(new_net_7587)
	);

	bfr new_net_7589_bfr_before (
		.din(new_net_7589),
		.dout(new_net_7588)
	);

	bfr new_net_7590_bfr_before (
		.din(new_net_7590),
		.dout(new_net_7589)
	);

	bfr new_net_7591_bfr_before (
		.din(new_net_7591),
		.dout(new_net_7590)
	);

	bfr new_net_7592_bfr_before (
		.din(new_net_7592),
		.dout(new_net_7591)
	);

	bfr new_net_7593_bfr_before (
		.din(new_net_7593),
		.dout(new_net_7592)
	);

	bfr new_net_7594_bfr_before (
		.din(new_net_7594),
		.dout(new_net_7593)
	);

	bfr new_net_7595_bfr_before (
		.din(new_net_7595),
		.dout(new_net_7594)
	);

	bfr new_net_7596_bfr_before (
		.din(new_net_7596),
		.dout(new_net_7595)
	);

	bfr new_net_7597_bfr_before (
		.din(new_net_7597),
		.dout(new_net_7596)
	);

	bfr new_net_7598_bfr_before (
		.din(new_net_7598),
		.dout(new_net_7597)
	);

	bfr new_net_7599_bfr_before (
		.din(new_net_7599),
		.dout(new_net_7598)
	);

	bfr new_net_7600_bfr_before (
		.din(new_net_7600),
		.dout(new_net_7599)
	);

	bfr new_net_7601_bfr_before (
		.din(new_net_7601),
		.dout(new_net_7600)
	);

	bfr new_net_7602_bfr_before (
		.din(new_net_7602),
		.dout(new_net_7601)
	);

	bfr new_net_7603_bfr_before (
		.din(new_net_7603),
		.dout(new_net_7602)
	);

	bfr new_net_7604_bfr_before (
		.din(new_net_7604),
		.dout(new_net_7603)
	);

	bfr new_net_7605_bfr_before (
		.din(new_net_7605),
		.dout(new_net_7604)
	);

	bfr new_net_7606_bfr_before (
		.din(new_net_7606),
		.dout(new_net_7605)
	);

	bfr new_net_7607_bfr_before (
		.din(new_net_7607),
		.dout(new_net_7606)
	);

	bfr new_net_7608_bfr_before (
		.din(new_net_7608),
		.dout(new_net_7607)
	);

	bfr new_net_7609_bfr_before (
		.din(new_net_7609),
		.dout(new_net_7608)
	);

	bfr new_net_7610_bfr_before (
		.din(new_net_7610),
		.dout(new_net_7609)
	);

	bfr new_net_7611_bfr_before (
		.din(new_net_7611),
		.dout(new_net_7610)
	);

	bfr new_net_7612_bfr_before (
		.din(new_net_7612),
		.dout(new_net_7611)
	);

	bfr new_net_7613_bfr_before (
		.din(new_net_7613),
		.dout(new_net_7612)
	);

	bfr new_net_7614_bfr_before (
		.din(new_net_7614),
		.dout(new_net_7613)
	);

	bfr new_net_7615_bfr_before (
		.din(new_net_7615),
		.dout(new_net_7614)
	);

	bfr new_net_7616_bfr_before (
		.din(new_net_7616),
		.dout(new_net_7615)
	);

	bfr new_net_7617_bfr_before (
		.din(new_net_7617),
		.dout(new_net_7616)
	);

	bfr new_net_7618_bfr_before (
		.din(new_net_7618),
		.dout(new_net_7617)
	);

	bfr new_net_7619_bfr_before (
		.din(new_net_7619),
		.dout(new_net_7618)
	);

	bfr new_net_7620_bfr_before (
		.din(new_net_7620),
		.dout(new_net_7619)
	);

	bfr new_net_7621_bfr_before (
		.din(new_net_7621),
		.dout(new_net_7620)
	);

	bfr new_net_7622_bfr_before (
		.din(new_net_7622),
		.dout(new_net_7621)
	);

	bfr new_net_7623_bfr_before (
		.din(new_net_7623),
		.dout(new_net_7622)
	);

	bfr new_net_7624_bfr_before (
		.din(new_net_7624),
		.dout(new_net_7623)
	);

	bfr new_net_7625_bfr_before (
		.din(new_net_7625),
		.dout(new_net_7624)
	);

	bfr new_net_7626_bfr_before (
		.din(new_net_7626),
		.dout(new_net_7625)
	);

	bfr new_net_7627_bfr_before (
		.din(new_net_7627),
		.dout(new_net_7626)
	);

	spl2 new_net_3_v_fanout (
		.a(new_net_3),
		.b(new_net_53),
		.c(new_net_7627)
	);

	bfr new_net_7628_bfr_after (
		.din(n_1341_),
		.dout(new_net_7628)
	);

	bfr new_net_7629_bfr_after (
		.din(new_net_7628),
		.dout(new_net_7629)
	);

	bfr new_net_7630_bfr_after (
		.din(new_net_7629),
		.dout(new_net_7630)
	);

	bfr new_net_7631_bfr_after (
		.din(new_net_7630),
		.dout(new_net_7631)
	);

	bfr new_net_7632_bfr_after (
		.din(new_net_7631),
		.dout(new_net_7632)
	);

	spl2 n_1341__v_fanout (
		.a(new_net_7632),
		.b(new_net_1697),
		.c(new_net_1696)
	);

	bfr new_net_7633_bfr_after (
		.din(n_0048_),
		.dout(new_net_7633)
	);

	bfr new_net_7634_bfr_after (
		.din(new_net_7633),
		.dout(new_net_7634)
	);

	bfr new_net_7635_bfr_after (
		.din(new_net_7634),
		.dout(new_net_7635)
	);

	bfr new_net_7636_bfr_after (
		.din(new_net_7635),
		.dout(new_net_7636)
	);

	bfr new_net_7637_bfr_after (
		.din(new_net_7636),
		.dout(new_net_7637)
	);

	spl2 n_0048__v_fanout (
		.a(new_net_7637),
		.b(new_net_1001),
		.c(new_net_1000)
	);

	bfr new_net_7638_bfr_before (
		.din(new_net_7638),
		.dout(N883)
	);

	bfr new_net_7639_bfr_before (
		.din(new_net_7639),
		.dout(new_net_7638)
	);

	bfr new_net_7640_bfr_before (
		.din(new_net_7640),
		.dout(new_net_7639)
	);

	bfr new_net_7641_bfr_before (
		.din(new_net_7641),
		.dout(new_net_7640)
	);

	bfr new_net_7642_bfr_before (
		.din(new_net_7642),
		.dout(new_net_7641)
	);

	bfr new_net_7643_bfr_before (
		.din(new_net_7643),
		.dout(new_net_7642)
	);

	bfr new_net_7644_bfr_before (
		.din(new_net_7644),
		.dout(new_net_7643)
	);

	bfr new_net_7645_bfr_before (
		.din(new_net_7645),
		.dout(new_net_7644)
	);

	bfr new_net_7646_bfr_before (
		.din(new_net_7646),
		.dout(new_net_7645)
	);

	bfr new_net_7647_bfr_before (
		.din(new_net_7647),
		.dout(new_net_7646)
	);

	bfr new_net_7648_bfr_before (
		.din(new_net_7648),
		.dout(new_net_7647)
	);

	bfr new_net_7649_bfr_before (
		.din(new_net_7649),
		.dout(new_net_7648)
	);

	bfr new_net_7650_bfr_before (
		.din(new_net_7650),
		.dout(new_net_7649)
	);

	bfr new_net_7651_bfr_before (
		.din(new_net_7651),
		.dout(new_net_7650)
	);

	bfr new_net_7652_bfr_before (
		.din(new_net_7652),
		.dout(new_net_7651)
	);

	bfr new_net_7653_bfr_before (
		.din(new_net_7653),
		.dout(new_net_7652)
	);

	bfr new_net_7654_bfr_before (
		.din(new_net_7654),
		.dout(new_net_7653)
	);

	bfr new_net_7655_bfr_before (
		.din(new_net_7655),
		.dout(new_net_7654)
	);

	bfr new_net_7656_bfr_before (
		.din(new_net_7656),
		.dout(new_net_7655)
	);

	bfr new_net_7657_bfr_before (
		.din(new_net_7657),
		.dout(new_net_7656)
	);

	bfr new_net_7658_bfr_before (
		.din(new_net_7658),
		.dout(new_net_7657)
	);

	bfr new_net_7659_bfr_before (
		.din(new_net_7659),
		.dout(new_net_7658)
	);

	bfr new_net_7660_bfr_before (
		.din(new_net_7660),
		.dout(new_net_7659)
	);

	bfr new_net_7661_bfr_before (
		.din(new_net_7661),
		.dout(new_net_7660)
	);

	bfr new_net_7662_bfr_before (
		.din(new_net_7662),
		.dout(new_net_7661)
	);

	bfr new_net_7663_bfr_before (
		.din(new_net_7663),
		.dout(new_net_7662)
	);

	bfr new_net_7664_bfr_before (
		.din(new_net_7664),
		.dout(new_net_7663)
	);

	bfr new_net_7665_bfr_before (
		.din(new_net_7665),
		.dout(new_net_7664)
	);

	bfr new_net_7666_bfr_before (
		.din(new_net_7666),
		.dout(new_net_7665)
	);

	bfr new_net_7667_bfr_before (
		.din(new_net_7667),
		.dout(new_net_7666)
	);

	bfr new_net_7668_bfr_before (
		.din(new_net_7668),
		.dout(new_net_7667)
	);

	bfr new_net_7669_bfr_before (
		.din(new_net_7669),
		.dout(new_net_7668)
	);

	bfr new_net_7670_bfr_before (
		.din(new_net_7670),
		.dout(new_net_7669)
	);

	bfr new_net_7671_bfr_before (
		.din(new_net_7671),
		.dout(new_net_7670)
	);

	bfr new_net_7672_bfr_before (
		.din(new_net_7672),
		.dout(new_net_7671)
	);

	bfr new_net_7673_bfr_before (
		.din(new_net_7673),
		.dout(new_net_7672)
	);

	bfr new_net_7674_bfr_before (
		.din(new_net_7674),
		.dout(new_net_7673)
	);

	bfr new_net_7675_bfr_before (
		.din(new_net_7675),
		.dout(new_net_7674)
	);

	bfr new_net_7676_bfr_before (
		.din(new_net_7676),
		.dout(new_net_7675)
	);

	bfr new_net_7677_bfr_before (
		.din(new_net_7677),
		.dout(new_net_7676)
	);

	bfr new_net_7678_bfr_before (
		.din(new_net_7678),
		.dout(new_net_7677)
	);

	bfr new_net_7679_bfr_before (
		.din(new_net_7679),
		.dout(new_net_7678)
	);

	bfr new_net_7680_bfr_before (
		.din(new_net_7680),
		.dout(new_net_7679)
	);

	bfr new_net_7681_bfr_before (
		.din(new_net_7681),
		.dout(new_net_7680)
	);

	bfr new_net_7682_bfr_before (
		.din(new_net_7682),
		.dout(new_net_7681)
	);

	bfr new_net_7683_bfr_before (
		.din(new_net_7683),
		.dout(new_net_7682)
	);

	bfr new_net_7684_bfr_before (
		.din(new_net_7684),
		.dout(new_net_7683)
	);

	bfr new_net_7685_bfr_before (
		.din(new_net_7685),
		.dout(new_net_7684)
	);

	bfr new_net_7686_bfr_before (
		.din(new_net_7686),
		.dout(new_net_7685)
	);

	bfr new_net_7687_bfr_before (
		.din(new_net_7687),
		.dout(new_net_7686)
	);

	bfr new_net_7688_bfr_before (
		.din(new_net_7688),
		.dout(new_net_7687)
	);

	bfr new_net_7689_bfr_before (
		.din(new_net_7689),
		.dout(new_net_7688)
	);

	bfr new_net_7690_bfr_before (
		.din(new_net_7690),
		.dout(new_net_7689)
	);

	bfr new_net_7691_bfr_before (
		.din(new_net_7691),
		.dout(new_net_7690)
	);

	bfr new_net_7692_bfr_before (
		.din(new_net_7692),
		.dout(new_net_7691)
	);

	bfr new_net_7693_bfr_before (
		.din(new_net_7693),
		.dout(new_net_7692)
	);

	bfr new_net_7694_bfr_before (
		.din(new_net_7694),
		.dout(new_net_7693)
	);

	bfr new_net_7695_bfr_before (
		.din(new_net_7695),
		.dout(new_net_7694)
	);

	bfr new_net_7696_bfr_before (
		.din(new_net_7696),
		.dout(new_net_7695)
	);

	bfr new_net_7697_bfr_before (
		.din(new_net_7697),
		.dout(new_net_7696)
	);

	bfr new_net_7698_bfr_before (
		.din(new_net_7698),
		.dout(new_net_7697)
	);

	bfr new_net_7699_bfr_before (
		.din(new_net_7699),
		.dout(new_net_7698)
	);

	bfr new_net_7700_bfr_before (
		.din(new_net_7700),
		.dout(new_net_7699)
	);

	spl2 new_net_0_v_fanout (
		.a(new_net_0),
		.b(new_net_1687),
		.c(new_net_7700)
	);

	spl4L new_net_1983_v_fanout (
		.a(new_net_1983),
		.b(new_net_1985),
		.c(new_net_1987),
		.d(new_net_1986),
		.e(new_net_1984)
	);

	spl4L new_net_1972_v_fanout (
		.a(new_net_1972),
		.b(new_net_1973),
		.c(new_net_1974),
		.d(new_net_1976),
		.e(new_net_1975)
	);

	spl4L new_net_1993_v_fanout (
		.a(new_net_1993),
		.b(new_net_1994),
		.c(new_net_1997),
		.d(new_net_1995),
		.e(new_net_1996)
	);

	bfr new_net_7701_bfr_after (
		.din(n_1293_),
		.dout(new_net_7701)
	);

	bfr new_net_7702_bfr_after (
		.din(new_net_7701),
		.dout(new_net_7702)
	);

	bfr new_net_7703_bfr_after (
		.din(new_net_7702),
		.dout(new_net_7703)
	);

	bfr new_net_7704_bfr_after (
		.din(new_net_7703),
		.dout(new_net_7704)
	);

	bfr new_net_7705_bfr_after (
		.din(new_net_7704),
		.dout(new_net_7705)
	);

	spl2 n_1293__v_fanout (
		.a(new_net_7705),
		.b(new_net_886),
		.c(new_net_885)
	);

	spl4L new_net_1978_v_fanout (
		.a(new_net_1978),
		.b(new_net_1981),
		.c(new_net_1980),
		.d(new_net_1982),
		.e(new_net_1979)
	);

	bfr new_net_7706_bfr_before (
		.din(new_net_7706),
		.dout(N882)
	);

	bfr new_net_7707_bfr_before (
		.din(new_net_7707),
		.dout(new_net_7706)
	);

	bfr new_net_7708_bfr_before (
		.din(new_net_7708),
		.dout(new_net_7707)
	);

	bfr new_net_7709_bfr_before (
		.din(new_net_7709),
		.dout(new_net_7708)
	);

	bfr new_net_7710_bfr_before (
		.din(new_net_7710),
		.dout(new_net_7709)
	);

	bfr new_net_7711_bfr_before (
		.din(new_net_7711),
		.dout(new_net_7710)
	);

	bfr new_net_7712_bfr_before (
		.din(new_net_7712),
		.dout(new_net_7711)
	);

	bfr new_net_7713_bfr_before (
		.din(new_net_7713),
		.dout(new_net_7712)
	);

	bfr new_net_7714_bfr_before (
		.din(new_net_7714),
		.dout(new_net_7713)
	);

	bfr new_net_7715_bfr_before (
		.din(new_net_7715),
		.dout(new_net_7714)
	);

	bfr new_net_7716_bfr_before (
		.din(new_net_7716),
		.dout(new_net_7715)
	);

	bfr new_net_7717_bfr_before (
		.din(new_net_7717),
		.dout(new_net_7716)
	);

	bfr new_net_7718_bfr_before (
		.din(new_net_7718),
		.dout(new_net_7717)
	);

	bfr new_net_7719_bfr_before (
		.din(new_net_7719),
		.dout(new_net_7718)
	);

	bfr new_net_7720_bfr_before (
		.din(new_net_7720),
		.dout(new_net_7719)
	);

	bfr new_net_7721_bfr_before (
		.din(new_net_7721),
		.dout(new_net_7720)
	);

	bfr new_net_7722_bfr_before (
		.din(new_net_7722),
		.dout(new_net_7721)
	);

	bfr new_net_7723_bfr_before (
		.din(new_net_7723),
		.dout(new_net_7722)
	);

	bfr new_net_7724_bfr_before (
		.din(new_net_7724),
		.dout(new_net_7723)
	);

	bfr new_net_7725_bfr_before (
		.din(new_net_7725),
		.dout(new_net_7724)
	);

	bfr new_net_7726_bfr_before (
		.din(new_net_7726),
		.dout(new_net_7725)
	);

	bfr new_net_7727_bfr_before (
		.din(new_net_7727),
		.dout(new_net_7726)
	);

	bfr new_net_7728_bfr_before (
		.din(new_net_7728),
		.dout(new_net_7727)
	);

	bfr new_net_7729_bfr_before (
		.din(new_net_7729),
		.dout(new_net_7728)
	);

	bfr new_net_7730_bfr_before (
		.din(new_net_7730),
		.dout(new_net_7729)
	);

	bfr new_net_7731_bfr_before (
		.din(new_net_7731),
		.dout(new_net_7730)
	);

	bfr new_net_7732_bfr_before (
		.din(new_net_7732),
		.dout(new_net_7731)
	);

	bfr new_net_7733_bfr_before (
		.din(new_net_7733),
		.dout(new_net_7732)
	);

	bfr new_net_7734_bfr_before (
		.din(new_net_7734),
		.dout(new_net_7733)
	);

	bfr new_net_7735_bfr_before (
		.din(new_net_7735),
		.dout(new_net_7734)
	);

	bfr new_net_7736_bfr_before (
		.din(new_net_7736),
		.dout(new_net_7735)
	);

	bfr new_net_7737_bfr_before (
		.din(new_net_7737),
		.dout(new_net_7736)
	);

	bfr new_net_7738_bfr_before (
		.din(new_net_7738),
		.dout(new_net_7737)
	);

	bfr new_net_7739_bfr_before (
		.din(new_net_7739),
		.dout(new_net_7738)
	);

	bfr new_net_7740_bfr_before (
		.din(new_net_7740),
		.dout(new_net_7739)
	);

	bfr new_net_7741_bfr_before (
		.din(new_net_7741),
		.dout(new_net_7740)
	);

	bfr new_net_7742_bfr_before (
		.din(new_net_7742),
		.dout(new_net_7741)
	);

	bfr new_net_7743_bfr_before (
		.din(new_net_7743),
		.dout(new_net_7742)
	);

	bfr new_net_7744_bfr_before (
		.din(new_net_7744),
		.dout(new_net_7743)
	);

	bfr new_net_7745_bfr_before (
		.din(new_net_7745),
		.dout(new_net_7744)
	);

	bfr new_net_7746_bfr_before (
		.din(new_net_7746),
		.dout(new_net_7745)
	);

	bfr new_net_7747_bfr_before (
		.din(new_net_7747),
		.dout(new_net_7746)
	);

	bfr new_net_7748_bfr_before (
		.din(new_net_7748),
		.dout(new_net_7747)
	);

	bfr new_net_7749_bfr_before (
		.din(new_net_7749),
		.dout(new_net_7748)
	);

	bfr new_net_7750_bfr_before (
		.din(new_net_7750),
		.dout(new_net_7749)
	);

	bfr new_net_7751_bfr_before (
		.din(new_net_7751),
		.dout(new_net_7750)
	);

	bfr new_net_7752_bfr_before (
		.din(new_net_7752),
		.dout(new_net_7751)
	);

	bfr new_net_7753_bfr_before (
		.din(new_net_7753),
		.dout(new_net_7752)
	);

	bfr new_net_7754_bfr_before (
		.din(new_net_7754),
		.dout(new_net_7753)
	);

	bfr new_net_7755_bfr_before (
		.din(new_net_7755),
		.dout(new_net_7754)
	);

	bfr new_net_7756_bfr_before (
		.din(new_net_7756),
		.dout(new_net_7755)
	);

	bfr new_net_7757_bfr_before (
		.din(new_net_7757),
		.dout(new_net_7756)
	);

	bfr new_net_7758_bfr_before (
		.din(new_net_7758),
		.dout(new_net_7757)
	);

	bfr new_net_7759_bfr_before (
		.din(new_net_7759),
		.dout(new_net_7758)
	);

	bfr new_net_7760_bfr_before (
		.din(new_net_7760),
		.dout(new_net_7759)
	);

	bfr new_net_7761_bfr_before (
		.din(new_net_7761),
		.dout(new_net_7760)
	);

	bfr new_net_7762_bfr_before (
		.din(new_net_7762),
		.dout(new_net_7761)
	);

	bfr new_net_7763_bfr_before (
		.din(new_net_7763),
		.dout(new_net_7762)
	);

	bfr new_net_7764_bfr_before (
		.din(new_net_7764),
		.dout(new_net_7763)
	);

	bfr new_net_7765_bfr_before (
		.din(new_net_7765),
		.dout(new_net_7764)
	);

	bfr new_net_7766_bfr_before (
		.din(new_net_7766),
		.dout(new_net_7765)
	);

	bfr new_net_7767_bfr_before (
		.din(new_net_7767),
		.dout(new_net_7766)
	);

	bfr new_net_7768_bfr_before (
		.din(new_net_7768),
		.dout(new_net_7767)
	);

	spl2 new_net_1_v_fanout (
		.a(new_net_1),
		.b(new_net_1391),
		.c(new_net_7768)
	);

	bfr new_net_7769_bfr_after (
		.din(n_1297_),
		.dout(new_net_7769)
	);

	bfr new_net_7770_bfr_after (
		.din(new_net_7769),
		.dout(new_net_7770)
	);

	bfr new_net_7771_bfr_after (
		.din(new_net_7770),
		.dout(new_net_7771)
	);

	bfr new_net_7772_bfr_after (
		.din(new_net_7771),
		.dout(new_net_7772)
	);

	bfr new_net_7773_bfr_after (
		.din(new_net_7772),
		.dout(new_net_7773)
	);

	spl2 n_1297__v_fanout (
		.a(new_net_7773),
		.b(new_net_1295),
		.c(new_net_1294)
	);

	bfr new_net_7774_bfr_before (
		.din(new_net_7774),
		.dout(new_net_1176)
	);

	bfr new_net_7775_bfr_before (
		.din(new_net_7775),
		.dout(new_net_7774)
	);

	bfr new_net_7776_bfr_before (
		.din(new_net_7776),
		.dout(new_net_7775)
	);

	spl2 n_0939__v_fanout (
		.a(n_0939_),
		.b(new_net_1177),
		.c(new_net_7776)
	);

	bfr new_net_7777_bfr_after (
		.din(n_1331_),
		.dout(new_net_7777)
	);

	bfr new_net_7778_bfr_after (
		.din(new_net_7777),
		.dout(new_net_7778)
	);

	bfr new_net_7779_bfr_after (
		.din(new_net_7778),
		.dout(new_net_7779)
	);

	bfr new_net_7780_bfr_after (
		.din(new_net_7779),
		.dout(new_net_7780)
	);

	bfr new_net_7781_bfr_after (
		.din(new_net_7780),
		.dout(new_net_7781)
	);

	spl2 n_1331__v_fanout (
		.a(new_net_7781),
		.b(new_net_585),
		.c(new_net_584)
	);

	spl4L new_net_1999_v_fanout (
		.a(new_net_1999),
		.b(new_net_2002),
		.c(new_net_2001),
		.d(new_net_2003),
		.e(new_net_2000)
	);

	spl4L new_net_2014_v_fanout (
		.a(new_net_2014),
		.b(new_net_2016),
		.c(new_net_2018),
		.d(new_net_2017),
		.e(new_net_2015)
	);

	spl4L new_net_2009_v_fanout (
		.a(new_net_2009),
		.b(new_net_2013),
		.c(new_net_2012),
		.d(new_net_2010),
		.e(new_net_2011)
	);

	bfr new_net_7782_bfr_before (
		.din(new_net_7782),
		.dout(N885)
	);

	bfr new_net_7783_bfr_before (
		.din(new_net_7783),
		.dout(new_net_7782)
	);

	bfr new_net_7784_bfr_before (
		.din(new_net_7784),
		.dout(new_net_7783)
	);

	bfr new_net_7785_bfr_before (
		.din(new_net_7785),
		.dout(new_net_7784)
	);

	bfr new_net_7786_bfr_before (
		.din(new_net_7786),
		.dout(new_net_7785)
	);

	bfr new_net_7787_bfr_before (
		.din(new_net_7787),
		.dout(new_net_7786)
	);

	bfr new_net_7788_bfr_before (
		.din(new_net_7788),
		.dout(new_net_7787)
	);

	bfr new_net_7789_bfr_before (
		.din(new_net_7789),
		.dout(new_net_7788)
	);

	bfr new_net_7790_bfr_before (
		.din(new_net_7790),
		.dout(new_net_7789)
	);

	bfr new_net_7791_bfr_before (
		.din(new_net_7791),
		.dout(new_net_7790)
	);

	bfr new_net_7792_bfr_before (
		.din(new_net_7792),
		.dout(new_net_7791)
	);

	bfr new_net_7793_bfr_before (
		.din(new_net_7793),
		.dout(new_net_7792)
	);

	bfr new_net_7794_bfr_before (
		.din(new_net_7794),
		.dout(new_net_7793)
	);

	bfr new_net_7795_bfr_before (
		.din(new_net_7795),
		.dout(new_net_7794)
	);

	bfr new_net_7796_bfr_before (
		.din(new_net_7796),
		.dout(new_net_7795)
	);

	bfr new_net_7797_bfr_before (
		.din(new_net_7797),
		.dout(new_net_7796)
	);

	bfr new_net_7798_bfr_before (
		.din(new_net_7798),
		.dout(new_net_7797)
	);

	bfr new_net_7799_bfr_before (
		.din(new_net_7799),
		.dout(new_net_7798)
	);

	bfr new_net_7800_bfr_before (
		.din(new_net_7800),
		.dout(new_net_7799)
	);

	bfr new_net_7801_bfr_before (
		.din(new_net_7801),
		.dout(new_net_7800)
	);

	bfr new_net_7802_bfr_before (
		.din(new_net_7802),
		.dout(new_net_7801)
	);

	bfr new_net_7803_bfr_before (
		.din(new_net_7803),
		.dout(new_net_7802)
	);

	bfr new_net_7804_bfr_before (
		.din(new_net_7804),
		.dout(new_net_7803)
	);

	bfr new_net_7805_bfr_before (
		.din(new_net_7805),
		.dout(new_net_7804)
	);

	bfr new_net_7806_bfr_before (
		.din(new_net_7806),
		.dout(new_net_7805)
	);

	bfr new_net_7807_bfr_before (
		.din(new_net_7807),
		.dout(new_net_7806)
	);

	bfr new_net_7808_bfr_before (
		.din(new_net_7808),
		.dout(new_net_7807)
	);

	bfr new_net_7809_bfr_before (
		.din(new_net_7809),
		.dout(new_net_7808)
	);

	bfr new_net_7810_bfr_before (
		.din(new_net_7810),
		.dout(new_net_7809)
	);

	bfr new_net_7811_bfr_before (
		.din(new_net_7811),
		.dout(new_net_7810)
	);

	bfr new_net_7812_bfr_before (
		.din(new_net_7812),
		.dout(new_net_7811)
	);

	bfr new_net_7813_bfr_before (
		.din(new_net_7813),
		.dout(new_net_7812)
	);

	bfr new_net_7814_bfr_before (
		.din(new_net_7814),
		.dout(new_net_7813)
	);

	bfr new_net_7815_bfr_before (
		.din(new_net_7815),
		.dout(new_net_7814)
	);

	bfr new_net_7816_bfr_before (
		.din(new_net_7816),
		.dout(new_net_7815)
	);

	bfr new_net_7817_bfr_before (
		.din(new_net_7817),
		.dout(new_net_7816)
	);

	bfr new_net_7818_bfr_before (
		.din(new_net_7818),
		.dout(new_net_7817)
	);

	bfr new_net_7819_bfr_before (
		.din(new_net_7819),
		.dout(new_net_7818)
	);

	bfr new_net_7820_bfr_before (
		.din(new_net_7820),
		.dout(new_net_7819)
	);

	bfr new_net_7821_bfr_before (
		.din(new_net_7821),
		.dout(new_net_7820)
	);

	bfr new_net_7822_bfr_before (
		.din(new_net_7822),
		.dout(new_net_7821)
	);

	bfr new_net_7823_bfr_before (
		.din(new_net_7823),
		.dout(new_net_7822)
	);

	bfr new_net_7824_bfr_before (
		.din(new_net_7824),
		.dout(new_net_7823)
	);

	bfr new_net_7825_bfr_before (
		.din(new_net_7825),
		.dout(new_net_7824)
	);

	bfr new_net_7826_bfr_before (
		.din(new_net_7826),
		.dout(new_net_7825)
	);

	bfr new_net_7827_bfr_before (
		.din(new_net_7827),
		.dout(new_net_7826)
	);

	bfr new_net_7828_bfr_before (
		.din(new_net_7828),
		.dout(new_net_7827)
	);

	bfr new_net_7829_bfr_before (
		.din(new_net_7829),
		.dout(new_net_7828)
	);

	bfr new_net_7830_bfr_before (
		.din(new_net_7830),
		.dout(new_net_7829)
	);

	bfr new_net_7831_bfr_before (
		.din(new_net_7831),
		.dout(new_net_7830)
	);

	bfr new_net_7832_bfr_before (
		.din(new_net_7832),
		.dout(new_net_7831)
	);

	bfr new_net_7833_bfr_before (
		.din(new_net_7833),
		.dout(new_net_7832)
	);

	bfr new_net_7834_bfr_before (
		.din(new_net_7834),
		.dout(new_net_7833)
	);

	bfr new_net_7835_bfr_before (
		.din(new_net_7835),
		.dout(new_net_7834)
	);

	bfr new_net_7836_bfr_before (
		.din(new_net_7836),
		.dout(new_net_7835)
	);

	bfr new_net_7837_bfr_before (
		.din(new_net_7837),
		.dout(new_net_7836)
	);

	bfr new_net_7838_bfr_before (
		.din(new_net_7838),
		.dout(new_net_7837)
	);

	bfr new_net_7839_bfr_before (
		.din(new_net_7839),
		.dout(new_net_7838)
	);

	bfr new_net_7840_bfr_before (
		.din(new_net_7840),
		.dout(new_net_7839)
	);

	bfr new_net_7841_bfr_before (
		.din(new_net_7841),
		.dout(new_net_7840)
	);

	bfr new_net_7842_bfr_before (
		.din(new_net_7842),
		.dout(new_net_7841)
	);

	bfr new_net_7843_bfr_before (
		.din(new_net_7843),
		.dout(new_net_7842)
	);

	bfr new_net_7844_bfr_before (
		.din(new_net_7844),
		.dout(new_net_7843)
	);

	spl2 new_net_2_v_fanout (
		.a(new_net_2),
		.b(new_net_1934),
		.c(new_net_7844)
	);

	spl4L new_net_1967_v_fanout (
		.a(new_net_1967),
		.b(new_net_1969),
		.c(new_net_1971),
		.d(new_net_1970),
		.e(new_net_1968)
	);

	bfr new_net_7845_bfr_before (
		.din(new_net_7845),
		.dout(new_net_316)
	);

	bfr new_net_7846_bfr_before (
		.din(new_net_7846),
		.dout(new_net_7845)
	);

	bfr new_net_7847_bfr_before (
		.din(new_net_7847),
		.dout(new_net_7846)
	);

	bfr new_net_7848_bfr_before (
		.din(new_net_7848),
		.dout(new_net_7847)
	);

	bfr new_net_7849_bfr_before (
		.din(new_net_7849),
		.dout(new_net_7848)
	);

	bfr new_net_7850_bfr_before (
		.din(new_net_7850),
		.dout(new_net_7849)
	);

	bfr new_net_7851_bfr_before (
		.din(new_net_7851),
		.dout(new_net_7850)
	);

	bfr new_net_7852_bfr_before (
		.din(new_net_7852),
		.dout(new_net_7851)
	);

	bfr new_net_7853_bfr_before (
		.din(new_net_7853),
		.dout(new_net_7852)
	);

	bfr new_net_7854_bfr_before (
		.din(new_net_7854),
		.dout(new_net_7853)
	);

	bfr new_net_7855_bfr_before (
		.din(new_net_7855),
		.dout(new_net_7854)
	);

	bfr new_net_7856_bfr_before (
		.din(new_net_7856),
		.dout(new_net_7855)
	);

	bfr new_net_7857_bfr_before (
		.din(new_net_7857),
		.dout(new_net_7856)
	);

	bfr new_net_7858_bfr_before (
		.din(new_net_7858),
		.dout(new_net_7857)
	);

	bfr new_net_7859_bfr_before (
		.din(new_net_7859),
		.dout(new_net_7858)
	);

	bfr new_net_7860_bfr_before (
		.din(new_net_7860),
		.dout(new_net_7859)
	);

	bfr new_net_7861_bfr_before (
		.din(new_net_7861),
		.dout(new_net_7860)
	);

	bfr new_net_7862_bfr_before (
		.din(new_net_7862),
		.dout(new_net_7861)
	);

	bfr new_net_7863_bfr_before (
		.din(new_net_7863),
		.dout(new_net_7862)
	);

	bfr new_net_7864_bfr_before (
		.din(new_net_7864),
		.dout(new_net_7863)
	);

	bfr new_net_7865_bfr_before (
		.din(new_net_7865),
		.dout(new_net_7864)
	);

	bfr new_net_7866_bfr_before (
		.din(new_net_7866),
		.dout(new_net_7865)
	);

	bfr new_net_7867_bfr_before (
		.din(new_net_7867),
		.dout(new_net_7866)
	);

	bfr new_net_7868_bfr_before (
		.din(new_net_7868),
		.dout(new_net_7867)
	);

	bfr new_net_7869_bfr_before (
		.din(new_net_7869),
		.dout(new_net_7868)
	);

	bfr new_net_7870_bfr_before (
		.din(new_net_7870),
		.dout(new_net_7869)
	);

	bfr new_net_7871_bfr_before (
		.din(new_net_7871),
		.dout(new_net_7870)
	);

	bfr new_net_7872_bfr_before (
		.din(new_net_7872),
		.dout(new_net_7871)
	);

	bfr new_net_7873_bfr_before (
		.din(new_net_7873),
		.dout(new_net_7872)
	);

	bfr new_net_7874_bfr_before (
		.din(new_net_7874),
		.dout(new_net_7873)
	);

	bfr new_net_7875_bfr_before (
		.din(new_net_7875),
		.dout(new_net_7874)
	);

	bfr new_net_7876_bfr_before (
		.din(new_net_7876),
		.dout(new_net_7875)
	);

	bfr new_net_7877_bfr_before (
		.din(new_net_7877),
		.dout(new_net_7876)
	);

	bfr new_net_7878_bfr_before (
		.din(new_net_7878),
		.dout(new_net_7877)
	);

	bfr new_net_7879_bfr_before (
		.din(new_net_7879),
		.dout(new_net_7878)
	);

	bfr new_net_7880_bfr_before (
		.din(new_net_7880),
		.dout(new_net_7879)
	);

	bfr new_net_7881_bfr_before (
		.din(new_net_7881),
		.dout(new_net_7880)
	);

	bfr new_net_7882_bfr_before (
		.din(new_net_7882),
		.dout(new_net_7881)
	);

	bfr new_net_7883_bfr_before (
		.din(new_net_7883),
		.dout(new_net_7882)
	);

	bfr new_net_7884_bfr_before (
		.din(new_net_7884),
		.dout(new_net_7883)
	);

	bfr new_net_7885_bfr_before (
		.din(new_net_7885),
		.dout(new_net_7884)
	);

	bfr new_net_7886_bfr_before (
		.din(new_net_7886),
		.dout(new_net_7885)
	);

	bfr new_net_7887_bfr_before (
		.din(new_net_7887),
		.dout(new_net_7886)
	);

	bfr new_net_7888_bfr_before (
		.din(new_net_7888),
		.dout(new_net_7887)
	);

	bfr new_net_7889_bfr_before (
		.din(new_net_7889),
		.dout(new_net_7888)
	);

	bfr new_net_7890_bfr_before (
		.din(new_net_7890),
		.dout(new_net_7889)
	);

	bfr new_net_7891_bfr_before (
		.din(new_net_7891),
		.dout(new_net_7890)
	);

	bfr new_net_7892_bfr_before (
		.din(new_net_7892),
		.dout(new_net_7891)
	);

	bfr new_net_7893_bfr_before (
		.din(new_net_7893),
		.dout(new_net_7892)
	);

	bfr new_net_7894_bfr_before (
		.din(new_net_7894),
		.dout(new_net_7893)
	);

	bfr new_net_7895_bfr_before (
		.din(new_net_7895),
		.dout(new_net_7894)
	);

	bfr new_net_7896_bfr_before (
		.din(new_net_7896),
		.dout(new_net_7895)
	);

	bfr new_net_7897_bfr_before (
		.din(new_net_7897),
		.dout(new_net_7896)
	);

	bfr new_net_7898_bfr_before (
		.din(new_net_7898),
		.dout(new_net_7897)
	);

	bfr new_net_7899_bfr_before (
		.din(new_net_7899),
		.dout(new_net_7898)
	);

	bfr new_net_7900_bfr_before (
		.din(new_net_7900),
		.dout(new_net_7899)
	);

	bfr new_net_7901_bfr_before (
		.din(new_net_7901),
		.dout(new_net_7900)
	);

	bfr new_net_7902_bfr_before (
		.din(new_net_7902),
		.dout(new_net_7901)
	);

	bfr new_net_7903_bfr_before (
		.din(new_net_7903),
		.dout(new_net_7902)
	);

	bfr new_net_7904_bfr_before (
		.din(new_net_7904),
		.dout(new_net_7903)
	);

	spl4L n_0162__v_fanout (
		.a(n_0162_),
		.b(new_net_315),
		.c(new_net_7904),
		.d(new_net_314),
		.e(new_net_313)
	);

	bfr new_net_7905_bfr_after (
		.din(n_1304_),
		.dout(new_net_7905)
	);

	bfr new_net_7906_bfr_after (
		.din(new_net_7905),
		.dout(new_net_7906)
	);

	bfr new_net_7907_bfr_after (
		.din(new_net_7906),
		.dout(new_net_7907)
	);

	bfr new_net_7908_bfr_after (
		.din(new_net_7907),
		.dout(new_net_7908)
	);

	bfr new_net_7909_bfr_after (
		.din(new_net_7908),
		.dout(new_net_7909)
	);

	spl2 n_1304__v_fanout (
		.a(new_net_7909),
		.b(new_net_1786),
		.c(new_net_1785)
	);

	bfr new_net_7910_bfr_after (
		.din(n_1307_),
		.dout(new_net_7910)
	);

	bfr new_net_7911_bfr_after (
		.din(new_net_7910),
		.dout(new_net_7911)
	);

	bfr new_net_7912_bfr_after (
		.din(new_net_7911),
		.dout(new_net_7912)
	);

	bfr new_net_7913_bfr_after (
		.din(new_net_7912),
		.dout(new_net_7913)
	);

	bfr new_net_7914_bfr_after (
		.din(new_net_7913),
		.dout(new_net_7914)
	);

	spl2 n_1307__v_fanout (
		.a(new_net_7914),
		.b(new_net_583),
		.c(new_net_582)
	);

	bfr new_net_7915_bfr_after (
		.din(n_1300_),
		.dout(new_net_7915)
	);

	bfr new_net_7916_bfr_after (
		.din(new_net_7915),
		.dout(new_net_7916)
	);

	bfr new_net_7917_bfr_after (
		.din(new_net_7916),
		.dout(new_net_7917)
	);

	bfr new_net_7918_bfr_after (
		.din(new_net_7917),
		.dout(new_net_7918)
	);

	bfr new_net_7919_bfr_after (
		.din(new_net_7918),
		.dout(new_net_7919)
	);

	spl2 n_1300__v_fanout (
		.a(new_net_7919),
		.b(new_net_1625),
		.c(new_net_1624)
	);

	spl2 n_0166__v_fanout (
		.a(n_0166_),
		.b(new_net_806),
		.c(new_net_805)
	);

	spl4L new_net_2004_v_fanout (
		.a(new_net_2004),
		.b(new_net_2006),
		.c(new_net_2008),
		.d(new_net_2007),
		.e(new_net_2005)
	);

	spl2 new_net_1964_v_fanout (
		.a(new_net_1964),
		.b(new_net_1966),
		.c(new_net_1965)
	);

	bfr new_net_7920_bfr_before (
		.din(new_net_7920),
		.dout(N489)
	);

	bfr new_net_7921_bfr_before (
		.din(new_net_7921),
		.dout(new_net_7920)
	);

	bfr new_net_7922_bfr_before (
		.din(new_net_7922),
		.dout(new_net_7921)
	);

	bfr new_net_7923_bfr_before (
		.din(new_net_7923),
		.dout(new_net_7922)
	);

	bfr new_net_7924_bfr_before (
		.din(new_net_7924),
		.dout(new_net_7923)
	);

	bfr new_net_7925_bfr_before (
		.din(new_net_7925),
		.dout(new_net_7924)
	);

	bfr new_net_7926_bfr_before (
		.din(new_net_7926),
		.dout(new_net_7925)
	);

	bfr new_net_7927_bfr_before (
		.din(new_net_7927),
		.dout(new_net_7926)
	);

	bfr new_net_7928_bfr_before (
		.din(new_net_7928),
		.dout(new_net_7927)
	);

	bfr new_net_7929_bfr_before (
		.din(new_net_7929),
		.dout(new_net_7928)
	);

	bfr new_net_7930_bfr_before (
		.din(new_net_7930),
		.dout(new_net_7929)
	);

	bfr new_net_7931_bfr_before (
		.din(new_net_7931),
		.dout(new_net_7930)
	);

	bfr new_net_7932_bfr_before (
		.din(new_net_7932),
		.dout(new_net_7931)
	);

	bfr new_net_7933_bfr_before (
		.din(new_net_7933),
		.dout(new_net_7932)
	);

	bfr new_net_7934_bfr_before (
		.din(new_net_7934),
		.dout(new_net_7933)
	);

	bfr new_net_7935_bfr_before (
		.din(new_net_7935),
		.dout(new_net_7934)
	);

	bfr new_net_7936_bfr_before (
		.din(new_net_7936),
		.dout(new_net_7935)
	);

	bfr new_net_7937_bfr_before (
		.din(new_net_7937),
		.dout(new_net_7936)
	);

	bfr new_net_7938_bfr_before (
		.din(new_net_7938),
		.dout(new_net_7937)
	);

	bfr new_net_7939_bfr_before (
		.din(new_net_7939),
		.dout(new_net_7938)
	);

	bfr new_net_7940_bfr_before (
		.din(new_net_7940),
		.dout(new_net_7939)
	);

	bfr new_net_7941_bfr_before (
		.din(new_net_7941),
		.dout(new_net_7940)
	);

	bfr new_net_7942_bfr_before (
		.din(new_net_7942),
		.dout(new_net_7941)
	);

	bfr new_net_7943_bfr_before (
		.din(new_net_7943),
		.dout(new_net_7942)
	);

	bfr new_net_7944_bfr_before (
		.din(new_net_7944),
		.dout(new_net_7943)
	);

	bfr new_net_7945_bfr_before (
		.din(new_net_7945),
		.dout(new_net_7944)
	);

	bfr new_net_7946_bfr_before (
		.din(new_net_7946),
		.dout(new_net_7945)
	);

	bfr new_net_7947_bfr_before (
		.din(new_net_7947),
		.dout(new_net_7946)
	);

	bfr new_net_7948_bfr_before (
		.din(new_net_7948),
		.dout(new_net_7947)
	);

	bfr new_net_7949_bfr_before (
		.din(new_net_7949),
		.dout(new_net_7948)
	);

	bfr new_net_7950_bfr_before (
		.din(new_net_7950),
		.dout(new_net_7949)
	);

	bfr new_net_7951_bfr_before (
		.din(new_net_7951),
		.dout(new_net_7950)
	);

	bfr new_net_7952_bfr_before (
		.din(new_net_7952),
		.dout(new_net_7951)
	);

	bfr new_net_7953_bfr_before (
		.din(new_net_7953),
		.dout(new_net_7952)
	);

	bfr new_net_7954_bfr_before (
		.din(new_net_7954),
		.dout(new_net_7953)
	);

	bfr new_net_7955_bfr_before (
		.din(new_net_7955),
		.dout(new_net_7954)
	);

	bfr new_net_7956_bfr_before (
		.din(new_net_7956),
		.dout(new_net_7955)
	);

	bfr new_net_7957_bfr_before (
		.din(new_net_7957),
		.dout(new_net_7956)
	);

	bfr new_net_7958_bfr_before (
		.din(new_net_7958),
		.dout(new_net_7957)
	);

	bfr new_net_7959_bfr_before (
		.din(new_net_7959),
		.dout(new_net_7958)
	);

	bfr new_net_7960_bfr_before (
		.din(new_net_7960),
		.dout(new_net_7959)
	);

	bfr new_net_7961_bfr_before (
		.din(new_net_7961),
		.dout(new_net_7960)
	);

	bfr new_net_7962_bfr_before (
		.din(new_net_7962),
		.dout(new_net_7961)
	);

	bfr new_net_7963_bfr_before (
		.din(new_net_7963),
		.dout(new_net_7962)
	);

	bfr new_net_7964_bfr_before (
		.din(new_net_7964),
		.dout(new_net_7963)
	);

	bfr new_net_7965_bfr_before (
		.din(new_net_7965),
		.dout(new_net_7964)
	);

	bfr new_net_7966_bfr_before (
		.din(new_net_7966),
		.dout(new_net_7965)
	);

	bfr new_net_7967_bfr_before (
		.din(new_net_7967),
		.dout(new_net_7966)
	);

	bfr new_net_7968_bfr_before (
		.din(new_net_7968),
		.dout(new_net_7967)
	);

	bfr new_net_7969_bfr_before (
		.din(new_net_7969),
		.dout(new_net_7968)
	);

	bfr new_net_7970_bfr_before (
		.din(new_net_7970),
		.dout(new_net_7969)
	);

	bfr new_net_7971_bfr_before (
		.din(new_net_7971),
		.dout(new_net_7970)
	);

	bfr new_net_7972_bfr_before (
		.din(new_net_7972),
		.dout(new_net_7971)
	);

	bfr new_net_7973_bfr_before (
		.din(new_net_7973),
		.dout(new_net_7972)
	);

	bfr new_net_7974_bfr_before (
		.din(new_net_7974),
		.dout(new_net_7973)
	);

	bfr new_net_7975_bfr_before (
		.din(new_net_7975),
		.dout(new_net_7974)
	);

	bfr new_net_7976_bfr_before (
		.din(new_net_7976),
		.dout(new_net_7975)
	);

	bfr new_net_7977_bfr_before (
		.din(new_net_7977),
		.dout(new_net_7976)
	);

	bfr new_net_7978_bfr_before (
		.din(new_net_7978),
		.dout(new_net_7977)
	);

	bfr new_net_7979_bfr_before (
		.din(new_net_7979),
		.dout(new_net_7978)
	);

	bfr new_net_7980_bfr_before (
		.din(new_net_7980),
		.dout(new_net_7979)
	);

	bfr new_net_7981_bfr_before (
		.din(new_net_7981),
		.dout(new_net_7980)
	);

	bfr new_net_7982_bfr_before (
		.din(new_net_7982),
		.dout(new_net_7981)
	);

	spl2 new_net_2025_v_fanout (
		.a(new_net_2025),
		.b(new_net_7982),
		.c(new_net_1467)
	);

	bfr new_net_7983_bfr_after (
		.din(n_1350_),
		.dout(new_net_7983)
	);

	bfr new_net_7984_bfr_after (
		.din(new_net_7983),
		.dout(new_net_7984)
	);

	bfr new_net_7985_bfr_after (
		.din(new_net_7984),
		.dout(new_net_7985)
	);

	bfr new_net_7986_bfr_after (
		.din(new_net_7985),
		.dout(new_net_7986)
	);

	bfr new_net_7987_bfr_after (
		.din(new_net_7986),
		.dout(new_net_7987)
	);

	spl2 n_1350__v_fanout (
		.a(new_net_7987),
		.b(new_net_810),
		.c(new_net_809)
	);

	spl3L n_0161__v_fanout (
		.a(n_0161_),
		.b(new_net_1618),
		.c(new_net_1616),
		.d(new_net_1617)
	);

	bfr new_net_7988_bfr_after (
		.din(n_1344_),
		.dout(new_net_7988)
	);

	bfr new_net_7989_bfr_after (
		.din(new_net_7988),
		.dout(new_net_7989)
	);

	bfr new_net_7990_bfr_after (
		.din(new_net_7989),
		.dout(new_net_7990)
	);

	bfr new_net_7991_bfr_after (
		.din(new_net_7990),
		.dout(new_net_7991)
	);

	bfr new_net_7992_bfr_after (
		.din(new_net_7991),
		.dout(new_net_7992)
	);

	spl2 n_1344__v_fanout (
		.a(new_net_7992),
		.b(new_net_14),
		.c(new_net_13)
	);

	bfr new_net_7993_bfr_after (
		.din(new_net_10),
		.dout(new_net_7993)
	);

	bfr new_net_7994_bfr_after (
		.din(new_net_7993),
		.dout(new_net_7994)
	);

	bfr new_net_7995_bfr_after (
		.din(new_net_7994),
		.dout(new_net_7995)
	);

	bfr new_net_7996_bfr_after (
		.din(new_net_7995),
		.dout(new_net_7996)
	);

	bfr new_net_7997_bfr_after (
		.din(new_net_7996),
		.dout(new_net_7997)
	);

	bfr new_net_7998_bfr_after (
		.din(new_net_7997),
		.dout(new_net_7998)
	);

	bfr new_net_7999_bfr_after (
		.din(new_net_7998),
		.dout(new_net_7999)
	);

	bfr new_net_8000_bfr_after (
		.din(new_net_7999),
		.dout(new_net_8000)
	);

	bfr new_net_8001_bfr_after (
		.din(new_net_8000),
		.dout(new_net_8001)
	);

	bfr new_net_8002_bfr_after (
		.din(new_net_8001),
		.dout(new_net_8002)
	);

	bfr new_net_8003_bfr_after (
		.din(new_net_8002),
		.dout(new_net_8003)
	);

	bfr new_net_8004_bfr_after (
		.din(new_net_8003),
		.dout(new_net_8004)
	);

	bfr new_net_8005_bfr_after (
		.din(new_net_8004),
		.dout(new_net_8005)
	);

	bfr new_net_8006_bfr_after (
		.din(new_net_8005),
		.dout(new_net_8006)
	);

	bfr new_net_8007_bfr_after (
		.din(new_net_8006),
		.dout(new_net_8007)
	);

	bfr new_net_8008_bfr_after (
		.din(new_net_8007),
		.dout(new_net_8008)
	);

	bfr new_net_8009_bfr_after (
		.din(new_net_8008),
		.dout(new_net_8009)
	);

	bfr new_net_8010_bfr_after (
		.din(new_net_8009),
		.dout(new_net_8010)
	);

	bfr new_net_8011_bfr_after (
		.din(new_net_8010),
		.dout(new_net_8011)
	);

	bfr new_net_8012_bfr_after (
		.din(new_net_8011),
		.dout(new_net_8012)
	);

	bfr new_net_8013_bfr_after (
		.din(new_net_8012),
		.dout(new_net_8013)
	);

	bfr new_net_8014_bfr_after (
		.din(new_net_8013),
		.dout(new_net_8014)
	);

	bfr new_net_8015_bfr_after (
		.din(new_net_8014),
		.dout(new_net_8015)
	);

	bfr new_net_8016_bfr_after (
		.din(new_net_8015),
		.dout(new_net_8016)
	);

	bfr new_net_8017_bfr_after (
		.din(new_net_8016),
		.dout(new_net_8017)
	);

	bfr new_net_8018_bfr_after (
		.din(new_net_8017),
		.dout(new_net_8018)
	);

	bfr new_net_8019_bfr_after (
		.din(new_net_8018),
		.dout(new_net_8019)
	);

	bfr new_net_8020_bfr_after (
		.din(new_net_8019),
		.dout(new_net_8020)
	);

	bfr new_net_8021_bfr_after (
		.din(new_net_8020),
		.dout(new_net_8021)
	);

	bfr new_net_8022_bfr_after (
		.din(new_net_8021),
		.dout(new_net_8022)
	);

	bfr new_net_8023_bfr_after (
		.din(new_net_8022),
		.dout(new_net_8023)
	);

	bfr new_net_8024_bfr_after (
		.din(new_net_8023),
		.dout(new_net_8024)
	);

	bfr new_net_8025_bfr_after (
		.din(new_net_8024),
		.dout(new_net_8025)
	);

	bfr new_net_8026_bfr_after (
		.din(new_net_8025),
		.dout(new_net_8026)
	);

	bfr new_net_8027_bfr_after (
		.din(new_net_8026),
		.dout(new_net_8027)
	);

	bfr new_net_8028_bfr_after (
		.din(new_net_8027),
		.dout(new_net_8028)
	);

	bfr new_net_8029_bfr_after (
		.din(new_net_8028),
		.dout(new_net_8029)
	);

	bfr new_net_8030_bfr_after (
		.din(new_net_8029),
		.dout(new_net_8030)
	);

	bfr new_net_8031_bfr_after (
		.din(new_net_8030),
		.dout(new_net_8031)
	);

	bfr new_net_8032_bfr_after (
		.din(new_net_8031),
		.dout(new_net_8032)
	);

	bfr new_net_8033_bfr_after (
		.din(new_net_8032),
		.dout(new_net_8033)
	);

	bfr new_net_8034_bfr_after (
		.din(new_net_8033),
		.dout(new_net_8034)
	);

	bfr new_net_8035_bfr_after (
		.din(new_net_8034),
		.dout(new_net_8035)
	);

	bfr new_net_8036_bfr_after (
		.din(new_net_8035),
		.dout(new_net_8036)
	);

	bfr new_net_8037_bfr_after (
		.din(new_net_8036),
		.dout(new_net_8037)
	);

	bfr new_net_8038_bfr_after (
		.din(new_net_8037),
		.dout(new_net_8038)
	);

	bfr new_net_8039_bfr_after (
		.din(new_net_8038),
		.dout(new_net_8039)
	);

	bfr new_net_8040_bfr_after (
		.din(new_net_8039),
		.dout(new_net_8040)
	);

	bfr new_net_8041_bfr_after (
		.din(new_net_8040),
		.dout(new_net_8041)
	);

	bfr new_net_8042_bfr_after (
		.din(new_net_8041),
		.dout(new_net_8042)
	);

	bfr new_net_8043_bfr_after (
		.din(new_net_8042),
		.dout(new_net_8043)
	);

	bfr new_net_8044_bfr_after (
		.din(new_net_8043),
		.dout(new_net_8044)
	);

	bfr new_net_8045_bfr_after (
		.din(new_net_8044),
		.dout(new_net_8045)
	);

	bfr new_net_8046_bfr_after (
		.din(new_net_8045),
		.dout(new_net_8046)
	);

	bfr new_net_8047_bfr_after (
		.din(new_net_8046),
		.dout(new_net_8047)
	);

	bfr new_net_8048_bfr_after (
		.din(new_net_8047),
		.dout(new_net_8048)
	);

	bfr new_net_8049_bfr_after (
		.din(new_net_8048),
		.dout(new_net_8049)
	);

	bfr new_net_8050_bfr_after (
		.din(new_net_8049),
		.dout(new_net_8050)
	);

	bfr new_net_8051_bfr_after (
		.din(new_net_8050),
		.dout(new_net_8051)
	);

	bfr new_net_8052_bfr_after (
		.din(new_net_8051),
		.dout(new_net_8052)
	);

	bfr new_net_8053_bfr_after (
		.din(new_net_8052),
		.dout(new_net_8053)
	);

	bfr new_net_8054_bfr_after (
		.din(new_net_8053),
		.dout(new_net_8054)
	);

	bfr new_net_8055_bfr_after (
		.din(new_net_8054),
		.dout(new_net_8055)
	);

	spl2 new_net_10_v_fanout (
		.a(new_net_8055),
		.b(N1112),
		.c(N1110)
	);

	bfr new_net_8056_bfr_after (
		.din(n_0718_),
		.dout(new_net_8056)
	);

	bfr new_net_8057_bfr_after (
		.din(new_net_8056),
		.dout(new_net_8057)
	);

	spl2 n_0718__v_fanout (
		.a(new_net_8057),
		.b(new_net_2059),
		.c(new_net_2057)
	);

	bfr new_net_8058_bfr_after (
		.din(new_net_11),
		.dout(new_net_8058)
	);

	bfr new_net_8059_bfr_after (
		.din(new_net_8058),
		.dout(new_net_8059)
	);

	bfr new_net_8060_bfr_after (
		.din(new_net_8059),
		.dout(new_net_8060)
	);

	bfr new_net_8061_bfr_after (
		.din(new_net_8060),
		.dout(new_net_8061)
	);

	bfr new_net_8062_bfr_after (
		.din(new_net_8061),
		.dout(new_net_8062)
	);

	bfr new_net_8063_bfr_after (
		.din(new_net_8062),
		.dout(new_net_8063)
	);

	bfr new_net_8064_bfr_after (
		.din(new_net_8063),
		.dout(new_net_8064)
	);

	bfr new_net_8065_bfr_after (
		.din(new_net_8064),
		.dout(new_net_8065)
	);

	bfr new_net_8066_bfr_after (
		.din(new_net_8065),
		.dout(new_net_8066)
	);

	bfr new_net_8067_bfr_after (
		.din(new_net_8066),
		.dout(new_net_8067)
	);

	bfr new_net_8068_bfr_after (
		.din(new_net_8067),
		.dout(new_net_8068)
	);

	bfr new_net_8069_bfr_after (
		.din(new_net_8068),
		.dout(new_net_8069)
	);

	bfr new_net_8070_bfr_after (
		.din(new_net_8069),
		.dout(new_net_8070)
	);

	bfr new_net_8071_bfr_after (
		.din(new_net_8070),
		.dout(new_net_8071)
	);

	bfr new_net_8072_bfr_after (
		.din(new_net_8071),
		.dout(new_net_8072)
	);

	bfr new_net_8073_bfr_after (
		.din(new_net_8072),
		.dout(new_net_8073)
	);

	bfr new_net_8074_bfr_after (
		.din(new_net_8073),
		.dout(new_net_8074)
	);

	bfr new_net_8075_bfr_after (
		.din(new_net_8074),
		.dout(new_net_8075)
	);

	bfr new_net_8076_bfr_after (
		.din(new_net_8075),
		.dout(new_net_8076)
	);

	bfr new_net_8077_bfr_after (
		.din(new_net_8076),
		.dout(new_net_8077)
	);

	bfr new_net_8078_bfr_after (
		.din(new_net_8077),
		.dout(new_net_8078)
	);

	bfr new_net_8079_bfr_after (
		.din(new_net_8078),
		.dout(new_net_8079)
	);

	bfr new_net_8080_bfr_after (
		.din(new_net_8079),
		.dout(new_net_8080)
	);

	bfr new_net_8081_bfr_after (
		.din(new_net_8080),
		.dout(new_net_8081)
	);

	bfr new_net_8082_bfr_after (
		.din(new_net_8081),
		.dout(new_net_8082)
	);

	bfr new_net_8083_bfr_after (
		.din(new_net_8082),
		.dout(new_net_8083)
	);

	bfr new_net_8084_bfr_after (
		.din(new_net_8083),
		.dout(new_net_8084)
	);

	bfr new_net_8085_bfr_after (
		.din(new_net_8084),
		.dout(new_net_8085)
	);

	bfr new_net_8086_bfr_after (
		.din(new_net_8085),
		.dout(new_net_8086)
	);

	bfr new_net_8087_bfr_after (
		.din(new_net_8086),
		.dout(new_net_8087)
	);

	bfr new_net_8088_bfr_after (
		.din(new_net_8087),
		.dout(new_net_8088)
	);

	bfr new_net_8089_bfr_after (
		.din(new_net_8088),
		.dout(new_net_8089)
	);

	bfr new_net_8090_bfr_after (
		.din(new_net_8089),
		.dout(new_net_8090)
	);

	bfr new_net_8091_bfr_after (
		.din(new_net_8090),
		.dout(new_net_8091)
	);

	bfr new_net_8092_bfr_after (
		.din(new_net_8091),
		.dout(new_net_8092)
	);

	bfr new_net_8093_bfr_after (
		.din(new_net_8092),
		.dout(new_net_8093)
	);

	bfr new_net_8094_bfr_after (
		.din(new_net_8093),
		.dout(new_net_8094)
	);

	bfr new_net_8095_bfr_after (
		.din(new_net_8094),
		.dout(new_net_8095)
	);

	bfr new_net_8096_bfr_after (
		.din(new_net_8095),
		.dout(new_net_8096)
	);

	bfr new_net_8097_bfr_after (
		.din(new_net_8096),
		.dout(new_net_8097)
	);

	bfr new_net_8098_bfr_after (
		.din(new_net_8097),
		.dout(new_net_8098)
	);

	bfr new_net_8099_bfr_after (
		.din(new_net_8098),
		.dout(new_net_8099)
	);

	bfr new_net_8100_bfr_after (
		.din(new_net_8099),
		.dout(new_net_8100)
	);

	bfr new_net_8101_bfr_after (
		.din(new_net_8100),
		.dout(new_net_8101)
	);

	bfr new_net_8102_bfr_after (
		.din(new_net_8101),
		.dout(new_net_8102)
	);

	bfr new_net_8103_bfr_after (
		.din(new_net_8102),
		.dout(new_net_8103)
	);

	bfr new_net_8104_bfr_after (
		.din(new_net_8103),
		.dout(new_net_8104)
	);

	bfr new_net_8105_bfr_after (
		.din(new_net_8104),
		.dout(new_net_8105)
	);

	bfr new_net_8106_bfr_after (
		.din(new_net_8105),
		.dout(new_net_8106)
	);

	bfr new_net_8107_bfr_after (
		.din(new_net_8106),
		.dout(new_net_8107)
	);

	bfr new_net_8108_bfr_after (
		.din(new_net_8107),
		.dout(new_net_8108)
	);

	bfr new_net_8109_bfr_after (
		.din(new_net_8108),
		.dout(new_net_8109)
	);

	bfr new_net_8110_bfr_after (
		.din(new_net_8109),
		.dout(new_net_8110)
	);

	bfr new_net_8111_bfr_after (
		.din(new_net_8110),
		.dout(new_net_8111)
	);

	bfr new_net_8112_bfr_after (
		.din(new_net_8111),
		.dout(new_net_8112)
	);

	bfr new_net_8113_bfr_after (
		.din(new_net_8112),
		.dout(new_net_8113)
	);

	bfr new_net_8114_bfr_after (
		.din(new_net_8113),
		.dout(new_net_8114)
	);

	bfr new_net_8115_bfr_after (
		.din(new_net_8114),
		.dout(new_net_8115)
	);

	bfr new_net_8116_bfr_after (
		.din(new_net_8115),
		.dout(new_net_8116)
	);

	bfr new_net_8117_bfr_after (
		.din(new_net_8116),
		.dout(new_net_8117)
	);

	bfr new_net_8118_bfr_after (
		.din(new_net_8117),
		.dout(new_net_8118)
	);

	bfr new_net_8119_bfr_after (
		.din(new_net_8118),
		.dout(new_net_8119)
	);

	bfr new_net_8120_bfr_after (
		.din(new_net_8119),
		.dout(new_net_8120)
	);

	bfr new_net_8121_bfr_after (
		.din(new_net_8120),
		.dout(new_net_8121)
	);

	spl3L new_net_11_v_fanout (
		.a(new_net_8121),
		.b(N1114),
		.c(N1111),
		.d(N582)
	);

	spl4L new_net_1977_v_fanout (
		.a(new_net_1977),
		.b(new_net_1993),
		.c(new_net_1983),
		.d(new_net_1988),
		.e(new_net_1978)
	);

	spl3L new_net_1963_v_fanout (
		.a(new_net_1963),
		.b(new_net_1967),
		.c(new_net_1964),
		.d(new_net_1972)
	);

	spl4L new_net_1998_v_fanout (
		.a(new_net_1998),
		.b(new_net_2014),
		.c(new_net_2009),
		.d(new_net_2004),
		.e(new_net_1999)
	);

	bfr new_net_8122_bfr_after (
		.din(N289),
		.dout(new_net_8122)
	);

	bfr new_net_8123_bfr_after (
		.din(new_net_8122),
		.dout(new_net_8123)
	);

	bfr new_net_8124_bfr_after (
		.din(new_net_8123),
		.dout(new_net_8124)
	);

	bfr new_net_8125_bfr_before (
		.din(new_net_8125),
		.dout(new_net_2030)
	);

	bfr new_net_8126_bfr_before (
		.din(new_net_8126),
		.dout(new_net_8125)
	);

	spl2 N289_v_fanout (
		.a(new_net_8124),
		.b(new_net_8126),
		.c(new_net_1575)
	);

	bfr new_net_8127_bfr_before (
		.din(new_net_8127),
		.dout(new_net_2041)
	);

	bfr new_net_8128_bfr_before (
		.din(new_net_8128),
		.dout(new_net_8127)
	);

	spl2 N325_v_fanout (
		.a(N325),
		.b(new_net_1433),
		.c(new_net_8128)
	);

	bfr new_net_8129_bfr_after (
		.din(N296),
		.dout(new_net_8129)
	);

	bfr new_net_8130_bfr_after (
		.din(new_net_8129),
		.dout(new_net_8130)
	);

	bfr new_net_8131_bfr_after (
		.din(new_net_8130),
		.dout(new_net_8131)
	);

	bfr new_net_8132_bfr_before (
		.din(new_net_8132),
		.dout(new_net_2032)
	);

	bfr new_net_8133_bfr_before (
		.din(new_net_8133),
		.dout(new_net_8132)
	);

	bfr new_net_8134_bfr_before (
		.din(new_net_8134),
		.dout(new_net_8133)
	);

	spl2 N296_v_fanout (
		.a(new_net_8131),
		.b(new_net_8134),
		.c(new_net_1877)
	);

	bfr new_net_8135_bfr_after (
		.din(N307),
		.dout(new_net_8135)
	);

	bfr new_net_8136_bfr_after (
		.din(new_net_8135),
		.dout(new_net_8136)
	);

	bfr new_net_8137_bfr_after (
		.din(new_net_8136),
		.dout(new_net_8137)
	);

	bfr new_net_8138_bfr_before (
		.din(new_net_8138),
		.dout(N535)
	);

	bfr new_net_8139_bfr_before (
		.din(new_net_8139),
		.dout(new_net_8138)
	);

	bfr new_net_8140_bfr_before (
		.din(new_net_8140),
		.dout(new_net_8139)
	);

	bfr new_net_8141_bfr_before (
		.din(new_net_8141),
		.dout(new_net_8140)
	);

	bfr new_net_8142_bfr_before (
		.din(new_net_8142),
		.dout(new_net_8141)
	);

	bfr new_net_8143_bfr_before (
		.din(new_net_8143),
		.dout(new_net_8142)
	);

	bfr new_net_8144_bfr_before (
		.din(new_net_8144),
		.dout(new_net_8143)
	);

	bfr new_net_8145_bfr_before (
		.din(new_net_8145),
		.dout(new_net_8144)
	);

	bfr new_net_8146_bfr_before (
		.din(new_net_8146),
		.dout(new_net_8145)
	);

	bfr new_net_8147_bfr_before (
		.din(new_net_8147),
		.dout(new_net_8146)
	);

	bfr new_net_8148_bfr_before (
		.din(new_net_8148),
		.dout(new_net_8147)
	);

	bfr new_net_8149_bfr_before (
		.din(new_net_8149),
		.dout(new_net_8148)
	);

	bfr new_net_8150_bfr_before (
		.din(new_net_8150),
		.dout(new_net_8149)
	);

	bfr new_net_8151_bfr_before (
		.din(new_net_8151),
		.dout(new_net_8150)
	);

	bfr new_net_8152_bfr_before (
		.din(new_net_8152),
		.dout(new_net_8151)
	);

	bfr new_net_8153_bfr_before (
		.din(new_net_8153),
		.dout(new_net_8152)
	);

	bfr new_net_8154_bfr_before (
		.din(new_net_8154),
		.dout(new_net_8153)
	);

	bfr new_net_8155_bfr_before (
		.din(new_net_8155),
		.dout(new_net_8154)
	);

	bfr new_net_8156_bfr_before (
		.din(new_net_8156),
		.dout(new_net_8155)
	);

	bfr new_net_8157_bfr_before (
		.din(new_net_8157),
		.dout(new_net_8156)
	);

	bfr new_net_8158_bfr_before (
		.din(new_net_8158),
		.dout(new_net_8157)
	);

	bfr new_net_8159_bfr_before (
		.din(new_net_8159),
		.dout(new_net_8158)
	);

	bfr new_net_8160_bfr_before (
		.din(new_net_8160),
		.dout(new_net_8159)
	);

	bfr new_net_8161_bfr_before (
		.din(new_net_8161),
		.dout(new_net_8160)
	);

	bfr new_net_8162_bfr_before (
		.din(new_net_8162),
		.dout(new_net_8161)
	);

	bfr new_net_8163_bfr_before (
		.din(new_net_8163),
		.dout(new_net_8162)
	);

	bfr new_net_8164_bfr_before (
		.din(new_net_8164),
		.dout(new_net_8163)
	);

	bfr new_net_8165_bfr_before (
		.din(new_net_8165),
		.dout(new_net_8164)
	);

	bfr new_net_8166_bfr_before (
		.din(new_net_8166),
		.dout(new_net_8165)
	);

	bfr new_net_8167_bfr_before (
		.din(new_net_8167),
		.dout(new_net_8166)
	);

	bfr new_net_8168_bfr_before (
		.din(new_net_8168),
		.dout(new_net_8167)
	);

	bfr new_net_8169_bfr_before (
		.din(new_net_8169),
		.dout(new_net_8168)
	);

	bfr new_net_8170_bfr_before (
		.din(new_net_8170),
		.dout(new_net_8169)
	);

	bfr new_net_8171_bfr_before (
		.din(new_net_8171),
		.dout(new_net_8170)
	);

	bfr new_net_8172_bfr_before (
		.din(new_net_8172),
		.dout(new_net_8171)
	);

	bfr new_net_8173_bfr_before (
		.din(new_net_8173),
		.dout(new_net_8172)
	);

	bfr new_net_8174_bfr_before (
		.din(new_net_8174),
		.dout(new_net_8173)
	);

	bfr new_net_8175_bfr_before (
		.din(new_net_8175),
		.dout(new_net_8174)
	);

	bfr new_net_8176_bfr_before (
		.din(new_net_8176),
		.dout(new_net_8175)
	);

	bfr new_net_8177_bfr_before (
		.din(new_net_8177),
		.dout(new_net_8176)
	);

	bfr new_net_8178_bfr_before (
		.din(new_net_8178),
		.dout(new_net_8177)
	);

	bfr new_net_8179_bfr_before (
		.din(new_net_8179),
		.dout(new_net_8178)
	);

	bfr new_net_8180_bfr_before (
		.din(new_net_8180),
		.dout(new_net_8179)
	);

	bfr new_net_8181_bfr_before (
		.din(new_net_8181),
		.dout(new_net_8180)
	);

	bfr new_net_8182_bfr_before (
		.din(new_net_8182),
		.dout(new_net_8181)
	);

	bfr new_net_8183_bfr_before (
		.din(new_net_8183),
		.dout(new_net_8182)
	);

	bfr new_net_8184_bfr_before (
		.din(new_net_8184),
		.dout(new_net_8183)
	);

	bfr new_net_8185_bfr_before (
		.din(new_net_8185),
		.dout(new_net_8184)
	);

	bfr new_net_8186_bfr_before (
		.din(new_net_8186),
		.dout(new_net_8185)
	);

	bfr new_net_8187_bfr_before (
		.din(new_net_8187),
		.dout(new_net_8186)
	);

	bfr new_net_8188_bfr_before (
		.din(new_net_8188),
		.dout(new_net_8187)
	);

	bfr new_net_8189_bfr_before (
		.din(new_net_8189),
		.dout(new_net_8188)
	);

	bfr new_net_8190_bfr_before (
		.din(new_net_8190),
		.dout(new_net_8189)
	);

	bfr new_net_8191_bfr_before (
		.din(new_net_8191),
		.dout(new_net_8190)
	);

	bfr new_net_8192_bfr_before (
		.din(new_net_8192),
		.dout(new_net_8191)
	);

	bfr new_net_8193_bfr_before (
		.din(new_net_8193),
		.dout(new_net_8192)
	);

	bfr new_net_8194_bfr_before (
		.din(new_net_8194),
		.dout(new_net_8193)
	);

	bfr new_net_8195_bfr_before (
		.din(new_net_8195),
		.dout(new_net_8194)
	);

	bfr new_net_8196_bfr_before (
		.din(new_net_8196),
		.dout(new_net_8195)
	);

	bfr new_net_8197_bfr_before (
		.din(new_net_8197),
		.dout(new_net_8196)
	);

	bfr new_net_8198_bfr_before (
		.din(new_net_8198),
		.dout(new_net_8197)
	);

	bfr new_net_8199_bfr_before (
		.din(new_net_8199),
		.dout(new_net_8198)
	);

	spl2 N307_v_fanout (
		.a(new_net_8137),
		.b(new_net_8199),
		.c(new_net_363)
	);

	bfr new_net_8200_bfr_before (
		.din(new_net_8200),
		.dout(new_net_2026)
	);

	bfr new_net_8201_bfr_before (
		.din(new_net_8201),
		.dout(new_net_8200)
	);

	spl2 N277_v_fanout (
		.a(N277),
		.b(new_net_1146),
		.c(new_net_8201)
	);

	bfr new_net_8202_bfr_before (
		.din(new_net_8202),
		.dout(new_net_2043)
	);

	bfr new_net_8203_bfr_before (
		.din(new_net_8203),
		.dout(new_net_8202)
	);

	spl2 N331_v_fanout (
		.a(N331),
		.b(new_net_1350),
		.c(new_net_8203)
	);

	bfr new_net_8204_bfr_after (
		.din(N328),
		.dout(new_net_8204)
	);

	bfr new_net_8205_bfr_after (
		.din(new_net_8204),
		.dout(new_net_8205)
	);

	bfr new_net_8206_bfr_after (
		.din(new_net_8205),
		.dout(new_net_8206)
	);

	bfr new_net_8207_bfr_before (
		.din(new_net_8207),
		.dout(new_net_2042)
	);

	bfr new_net_8208_bfr_before (
		.din(new_net_8208),
		.dout(new_net_8207)
	);

	bfr new_net_8209_bfr_before (
		.din(new_net_8209),
		.dout(new_net_8208)
	);

	spl2 N328_v_fanout (
		.a(new_net_8206),
		.b(new_net_8209),
		.c(new_net_1225)
	);

	bfr new_net_8210_bfr_after (
		.din(N303),
		.dout(new_net_8210)
	);

	bfr new_net_8211_bfr_after (
		.din(new_net_8210),
		.dout(new_net_8211)
	);

	bfr new_net_8212_bfr_after (
		.din(new_net_8211),
		.dout(new_net_8212)
	);

	bfr new_net_8213_bfr_before (
		.din(new_net_8213),
		.dout(new_net_2034)
	);

	bfr new_net_8214_bfr_before (
		.din(new_net_8214),
		.dout(new_net_8213)
	);

	bfr new_net_8215_bfr_before (
		.din(new_net_8215),
		.dout(new_net_8214)
	);

	spl2 N303_v_fanout (
		.a(new_net_8212),
		.b(new_net_8215),
		.c(new_net_1266)
	);

	spl2 N164_v_fanout (
		.a(N164),
		.b(new_net_552),
		.c(new_net_551)
	);

	spl3L N5_v_fanout (
		.a(N5),
		.b(new_net_828),
		.c(new_net_826),
		.d(new_net_827)
	);

	bfr new_net_8216_bfr_before (
		.din(new_net_8216),
		.dout(new_net_2051)
	);

	bfr new_net_8217_bfr_before (
		.din(new_net_8217),
		.dout(new_net_8216)
	);

	spl2 N358_v_fanout (
		.a(N358),
		.b(new_net_652),
		.c(new_net_8217)
	);

	bfr new_net_8218_bfr_after (
		.din(N340),
		.dout(new_net_8218)
	);

	bfr new_net_8219_bfr_after (
		.din(new_net_8218),
		.dout(new_net_8219)
	);

	bfr new_net_8220_bfr_after (
		.din(new_net_8219),
		.dout(new_net_8220)
	);

	bfr new_net_8221_bfr_before (
		.din(new_net_8221),
		.dout(new_net_2045)
	);

	bfr new_net_8222_bfr_before (
		.din(new_net_8222),
		.dout(new_net_8221)
	);

	bfr new_net_8223_bfr_before (
		.din(new_net_8223),
		.dout(new_net_8222)
	);

	spl2 N340_v_fanout (
		.a(new_net_8220),
		.b(new_net_8223),
		.c(new_net_1560)
	);

	bfr new_net_8224_bfr_after (
		.din(N257),
		.dout(new_net_8224)
	);

	bfr new_net_8225_bfr_after (
		.din(new_net_8224),
		.dout(new_net_8225)
	);

	bfr new_net_8226_bfr_after (
		.din(new_net_8225),
		.dout(new_net_8226)
	);

	bfr new_net_8227_bfr_before (
		.din(new_net_8227),
		.dout(new_net_2023)
	);

	bfr new_net_8228_bfr_before (
		.din(new_net_8228),
		.dout(new_net_8227)
	);

	bfr new_net_8229_bfr_before (
		.din(new_net_8229),
		.dout(new_net_8228)
	);

	spl2 N257_v_fanout (
		.a(new_net_8226),
		.b(new_net_8229),
		.c(new_net_1805)
	);

	bfr new_net_8230_bfr_after (
		.din(N106),
		.dout(new_net_8230)
	);

	bfr new_net_8231_bfr_after (
		.din(new_net_8230),
		.dout(new_net_8231)
	);

	bfr new_net_8232_bfr_after (
		.din(new_net_8231),
		.dout(new_net_8232)
	);

	bfr new_net_8233_bfr_before (
		.din(new_net_8233),
		.dout(new_net_1962)
	);

	bfr new_net_8234_bfr_before (
		.din(new_net_8234),
		.dout(new_net_8233)
	);

	bfr new_net_8235_bfr_before (
		.din(new_net_8235),
		.dout(new_net_8234)
	);

	spl2 N106_v_fanout (
		.a(new_net_8232),
		.b(new_net_8235),
		.c(new_net_1722)
	);

	bfr new_net_8236_bfr_after (
		.din(N352),
		.dout(new_net_8236)
	);

	bfr new_net_8237_bfr_after (
		.din(new_net_8236),
		.dout(new_net_8237)
	);

	bfr new_net_8238_bfr_after (
		.din(new_net_8237),
		.dout(new_net_8238)
	);

	bfr new_net_8239_bfr_before (
		.din(new_net_8239),
		.dout(new_net_2049)
	);

	bfr new_net_8240_bfr_before (
		.din(new_net_8240),
		.dout(new_net_8239)
	);

	bfr new_net_8241_bfr_before (
		.din(new_net_8241),
		.dout(new_net_8240)
	);

	spl2 N352_v_fanout (
		.a(new_net_8238),
		.b(new_net_8241),
		.c(new_net_1659)
	);

	bfr new_net_8242_bfr_before (
		.din(new_net_8242),
		.dout(new_net_2050)
	);

	bfr new_net_8243_bfr_before (
		.din(new_net_8243),
		.dout(new_net_8242)
	);

	spl2 N355_v_fanout (
		.a(N355),
		.b(new_net_520),
		.c(new_net_8243)
	);

	spl2 N212_v_fanout (
		.a(N212),
		.b(new_net_1058),
		.c(new_net_1057)
	);

	bfr new_net_8244_bfr_after (
		.din(N260),
		.dout(new_net_8244)
	);

	bfr new_net_8245_bfr_after (
		.din(new_net_8244),
		.dout(new_net_8245)
	);

	bfr new_net_8246_bfr_after (
		.din(new_net_8245),
		.dout(new_net_8246)
	);

	bfr new_net_8247_bfr_before (
		.din(new_net_8247),
		.dout(new_net_2024)
	);

	bfr new_net_8248_bfr_before (
		.din(new_net_8248),
		.dout(new_net_8247)
	);

	bfr new_net_8249_bfr_before (
		.din(new_net_8249),
		.dout(new_net_8248)
	);

	spl2 N260_v_fanout (
		.a(new_net_8246),
		.b(new_net_8249),
		.c(new_net_1343)
	);

	bfr new_net_8250_bfr_after (
		.din(N319),
		.dout(new_net_8250)
	);

	bfr new_net_8251_bfr_after (
		.din(new_net_8250),
		.dout(new_net_8251)
	);

	bfr new_net_8252_bfr_after (
		.din(new_net_8251),
		.dout(new_net_8252)
	);

	bfr new_net_8253_bfr_before (
		.din(new_net_8253),
		.dout(new_net_2039)
	);

	bfr new_net_8254_bfr_before (
		.din(new_net_8254),
		.dout(new_net_8253)
	);

	bfr new_net_8255_bfr_before (
		.din(new_net_8255),
		.dout(new_net_8254)
	);

	spl2 N319_v_fanout (
		.a(new_net_8252),
		.b(new_net_1389),
		.c(new_net_8255)
	);

	spl2 N165_v_fanout (
		.a(N165),
		.b(new_net_1776),
		.c(new_net_1775)
	);

	bfr new_net_8256_bfr_before (
		.din(new_net_8256),
		.dout(new_net_2040)
	);

	bfr new_net_8257_bfr_before (
		.din(new_net_8257),
		.dout(new_net_8256)
	);

	spl2 N322_v_fanout (
		.a(N322),
		.b(new_net_8257),
		.c(new_net_1078)
	);

	bfr new_net_8258_bfr_after (
		.din(N349),
		.dout(new_net_8258)
	);

	bfr new_net_8259_bfr_after (
		.din(new_net_8258),
		.dout(new_net_8259)
	);

	bfr new_net_8260_bfr_after (
		.din(new_net_8259),
		.dout(new_net_8260)
	);

	bfr new_net_8261_bfr_before (
		.din(new_net_8261),
		.dout(new_net_2048)
	);

	bfr new_net_8262_bfr_before (
		.din(new_net_8262),
		.dout(new_net_8261)
	);

	bfr new_net_8263_bfr_before (
		.din(new_net_8263),
		.dout(new_net_8262)
	);

	spl2 N349_v_fanout (
		.a(new_net_8260),
		.b(new_net_8263),
		.c(new_net_1607)
	);

	bfr new_net_8264_bfr_after (
		.din(N41),
		.dout(new_net_8264)
	);

	bfr new_net_8265_bfr_after (
		.din(new_net_8264),
		.dout(new_net_8265)
	);

	bfr new_net_8266_bfr_after (
		.din(new_net_8265),
		.dout(new_net_8266)
	);

	spl2 N41_v_fanout (
		.a(new_net_8266),
		.b(new_net_1487),
		.c(new_net_1486)
	);

	bfr new_net_8267_bfr_after (
		.din(N310),
		.dout(new_net_8267)
	);

	bfr new_net_8268_bfr_after (
		.din(new_net_8267),
		.dout(new_net_8268)
	);

	bfr new_net_8269_bfr_after (
		.din(new_net_8268),
		.dout(new_net_8269)
	);

	spl2 N310_v_fanout (
		.a(new_net_8269),
		.b(new_net_513),
		.c(new_net_2035)
	);

	bfr new_net_8270_bfr_before (
		.din(new_net_8270),
		.dout(N492)
	);

	bfr new_net_8271_bfr_before (
		.din(new_net_8271),
		.dout(new_net_8270)
	);

	bfr new_net_8272_bfr_before (
		.din(new_net_8272),
		.dout(new_net_8271)
	);

	bfr new_net_8273_bfr_before (
		.din(new_net_8273),
		.dout(new_net_8272)
	);

	bfr new_net_8274_bfr_before (
		.din(new_net_8274),
		.dout(new_net_8273)
	);

	bfr new_net_8275_bfr_before (
		.din(new_net_8275),
		.dout(new_net_8274)
	);

	bfr new_net_8276_bfr_before (
		.din(new_net_8276),
		.dout(new_net_8275)
	);

	bfr new_net_8277_bfr_before (
		.din(new_net_8277),
		.dout(new_net_8276)
	);

	bfr new_net_8278_bfr_before (
		.din(new_net_8278),
		.dout(new_net_8277)
	);

	bfr new_net_8279_bfr_before (
		.din(new_net_8279),
		.dout(new_net_8278)
	);

	bfr new_net_8280_bfr_before (
		.din(new_net_8280),
		.dout(new_net_8279)
	);

	bfr new_net_8281_bfr_before (
		.din(new_net_8281),
		.dout(new_net_8280)
	);

	bfr new_net_8282_bfr_before (
		.din(new_net_8282),
		.dout(new_net_8281)
	);

	bfr new_net_8283_bfr_before (
		.din(new_net_8283),
		.dout(new_net_8282)
	);

	bfr new_net_8284_bfr_before (
		.din(new_net_8284),
		.dout(new_net_8283)
	);

	bfr new_net_8285_bfr_before (
		.din(new_net_8285),
		.dout(new_net_8284)
	);

	bfr new_net_8286_bfr_before (
		.din(new_net_8286),
		.dout(new_net_8285)
	);

	bfr new_net_8287_bfr_before (
		.din(new_net_8287),
		.dout(new_net_8286)
	);

	bfr new_net_8288_bfr_before (
		.din(new_net_8288),
		.dout(new_net_8287)
	);

	bfr new_net_8289_bfr_before (
		.din(new_net_8289),
		.dout(new_net_8288)
	);

	bfr new_net_8290_bfr_before (
		.din(new_net_8290),
		.dout(new_net_8289)
	);

	bfr new_net_8291_bfr_before (
		.din(new_net_8291),
		.dout(new_net_8290)
	);

	bfr new_net_8292_bfr_before (
		.din(new_net_8292),
		.dout(new_net_8291)
	);

	bfr new_net_8293_bfr_before (
		.din(new_net_8293),
		.dout(new_net_8292)
	);

	bfr new_net_8294_bfr_before (
		.din(new_net_8294),
		.dout(new_net_8293)
	);

	bfr new_net_8295_bfr_before (
		.din(new_net_8295),
		.dout(new_net_8294)
	);

	bfr new_net_8296_bfr_before (
		.din(new_net_8296),
		.dout(new_net_8295)
	);

	bfr new_net_8297_bfr_before (
		.din(new_net_8297),
		.dout(new_net_8296)
	);

	bfr new_net_8298_bfr_before (
		.din(new_net_8298),
		.dout(new_net_8297)
	);

	bfr new_net_8299_bfr_before (
		.din(new_net_8299),
		.dout(new_net_8298)
	);

	bfr new_net_8300_bfr_before (
		.din(new_net_8300),
		.dout(new_net_8299)
	);

	bfr new_net_8301_bfr_before (
		.din(new_net_8301),
		.dout(new_net_8300)
	);

	bfr new_net_8302_bfr_before (
		.din(new_net_8302),
		.dout(new_net_8301)
	);

	bfr new_net_8303_bfr_before (
		.din(new_net_8303),
		.dout(new_net_8302)
	);

	bfr new_net_8304_bfr_before (
		.din(new_net_8304),
		.dout(new_net_8303)
	);

	bfr new_net_8305_bfr_before (
		.din(new_net_8305),
		.dout(new_net_8304)
	);

	bfr new_net_8306_bfr_before (
		.din(new_net_8306),
		.dout(new_net_8305)
	);

	bfr new_net_8307_bfr_before (
		.din(new_net_8307),
		.dout(new_net_8306)
	);

	bfr new_net_8308_bfr_before (
		.din(new_net_8308),
		.dout(new_net_8307)
	);

	bfr new_net_8309_bfr_before (
		.din(new_net_8309),
		.dout(new_net_8308)
	);

	bfr new_net_8310_bfr_before (
		.din(new_net_8310),
		.dout(new_net_8309)
	);

	bfr new_net_8311_bfr_before (
		.din(new_net_8311),
		.dout(new_net_8310)
	);

	bfr new_net_8312_bfr_before (
		.din(new_net_8312),
		.dout(new_net_8311)
	);

	bfr new_net_8313_bfr_before (
		.din(new_net_8313),
		.dout(new_net_8312)
	);

	bfr new_net_8314_bfr_before (
		.din(new_net_8314),
		.dout(new_net_8313)
	);

	bfr new_net_8315_bfr_before (
		.din(new_net_8315),
		.dout(new_net_8314)
	);

	bfr new_net_8316_bfr_before (
		.din(new_net_8316),
		.dout(new_net_8315)
	);

	bfr new_net_8317_bfr_before (
		.din(new_net_8317),
		.dout(new_net_8316)
	);

	bfr new_net_8318_bfr_before (
		.din(new_net_8318),
		.dout(new_net_8317)
	);

	bfr new_net_8319_bfr_before (
		.din(new_net_8319),
		.dout(new_net_8318)
	);

	bfr new_net_8320_bfr_before (
		.din(new_net_8320),
		.dout(new_net_8319)
	);

	bfr new_net_8321_bfr_before (
		.din(new_net_8321),
		.dout(new_net_8320)
	);

	bfr new_net_8322_bfr_before (
		.din(new_net_8322),
		.dout(new_net_8321)
	);

	bfr new_net_8323_bfr_before (
		.din(new_net_8323),
		.dout(new_net_8322)
	);

	bfr new_net_8324_bfr_before (
		.din(new_net_8324),
		.dout(new_net_8323)
	);

	bfr new_net_8325_bfr_before (
		.din(new_net_8325),
		.dout(new_net_8324)
	);

	bfr new_net_8326_bfr_before (
		.din(new_net_8326),
		.dout(new_net_8325)
	);

	bfr new_net_8327_bfr_before (
		.din(new_net_8327),
		.dout(new_net_8326)
	);

	bfr new_net_8328_bfr_before (
		.din(new_net_8328),
		.dout(new_net_8327)
	);

	bfr new_net_8329_bfr_before (
		.din(new_net_8329),
		.dout(new_net_8328)
	);

	bfr new_net_8330_bfr_before (
		.din(new_net_8330),
		.dout(new_net_8329)
	);

	bfr new_net_8331_bfr_before (
		.din(new_net_8331),
		.dout(new_net_8330)
	);

	bfr new_net_8332_bfr_before (
		.din(new_net_8332),
		.dout(new_net_8331)
	);

	bfr new_net_8333_bfr_before (
		.din(new_net_8333),
		.dout(new_net_8332)
	);

	bfr new_net_8334_bfr_before (
		.din(new_net_8334),
		.dout(new_net_8333)
	);

	spl4L N267_v_fanout (
		.a(N267),
		.b(new_net_1917),
		.c(new_net_8334),
		.d(new_net_1918),
		.e(new_net_1915)
	);

	spl2 N211_v_fanout (
		.a(N211),
		.b(new_net_1033),
		.c(new_net_1032)
	);

	bfr new_net_8335_bfr_after (
		.din(N313),
		.dout(new_net_8335)
	);

	bfr new_net_8336_bfr_after (
		.din(new_net_8335),
		.dout(new_net_8336)
	);

	bfr new_net_8337_bfr_after (
		.din(new_net_8336),
		.dout(new_net_8337)
	);

	bfr new_net_8338_bfr_before (
		.din(new_net_8338),
		.dout(new_net_2037)
	);

	bfr new_net_8339_bfr_before (
		.din(new_net_8339),
		.dout(new_net_8338)
	);

	bfr new_net_8340_bfr_before (
		.din(new_net_8340),
		.dout(new_net_8339)
	);

	spl2 N313_v_fanout (
		.a(new_net_8337),
		.b(new_net_1332),
		.c(new_net_8340)
	);

	bfr new_net_8341_bfr_before (
		.din(new_net_8341),
		.dout(new_net_2053)
	);

	bfr new_net_8342_bfr_before (
		.din(new_net_8342),
		.dout(new_net_8341)
	);

	spl2 N364_v_fanout (
		.a(N364),
		.b(new_net_850),
		.c(new_net_8342)
	);

	bfr new_net_8343_bfr_after (
		.din(N299),
		.dout(new_net_8343)
	);

	bfr new_net_8344_bfr_after (
		.din(new_net_8343),
		.dout(new_net_8344)
	);

	bfr new_net_8345_bfr_after (
		.din(new_net_8344),
		.dout(new_net_8345)
	);

	bfr new_net_8346_bfr_before (
		.din(new_net_8346),
		.dout(new_net_2033)
	);

	bfr new_net_8347_bfr_before (
		.din(new_net_8347),
		.dout(new_net_8346)
	);

	bfr new_net_8348_bfr_before (
		.din(new_net_8348),
		.dout(new_net_8347)
	);

	spl2 N299_v_fanout (
		.a(new_net_8345),
		.b(new_net_8348),
		.c(new_net_1233)
	);

	bfr new_net_8349_bfr_after (
		.din(N254),
		.dout(new_net_8349)
	);

	bfr new_net_8350_bfr_after (
		.din(new_net_8349),
		.dout(new_net_8350)
	);

	bfr new_net_8351_bfr_after (
		.din(new_net_8350),
		.dout(new_net_8351)
	);

	bfr new_net_8352_bfr_before (
		.din(new_net_8352),
		.dout(new_net_2022)
	);

	bfr new_net_8353_bfr_before (
		.din(new_net_8353),
		.dout(new_net_8352)
	);

	bfr new_net_8354_bfr_before (
		.din(new_net_8354),
		.dout(new_net_8353)
	);

	spl2 N254_v_fanout (
		.a(new_net_8351),
		.b(new_net_8354),
		.c(new_net_1069)
	);

	bfr new_net_8355_bfr_before (
		.din(new_net_8355),
		.dout(new_net_1431)
	);

	bfr new_net_8356_bfr_before (
		.din(new_net_8356),
		.dout(new_net_8355)
	);

	bfr new_net_8357_bfr_before (
		.din(new_net_8357),
		.dout(new_net_8356)
	);

	bfr new_net_8358_bfr_before (
		.din(new_net_8358),
		.dout(new_net_8357)
	);

	bfr new_net_8359_bfr_before (
		.din(new_net_8359),
		.dout(new_net_8358)
	);

	spl2 N89_v_fanout (
		.a(N89),
		.b(new_net_8359),
		.c(new_net_1430)
	);

	bfr new_net_8360_bfr_before (
		.din(new_net_8360),
		.dout(new_net_2047)
	);

	bfr new_net_8361_bfr_before (
		.din(new_net_8361),
		.dout(new_net_8360)
	);

	spl2 N346_v_fanout (
		.a(N346),
		.b(new_net_1896),
		.c(new_net_8361)
	);

	bfr new_net_8362_bfr_before (
		.din(new_net_8362),
		.dout(new_net_2054)
	);

	bfr new_net_8363_bfr_before (
		.din(new_net_8363),
		.dout(new_net_8362)
	);

	bfr new_net_8364_bfr_before (
		.din(new_net_8364),
		.dout(new_net_8363)
	);

	bfr new_net_8365_bfr_before (
		.din(new_net_8365),
		.dout(new_net_8364)
	);

	bfr new_net_8366_bfr_before (
		.din(new_net_8366),
		.dout(new_net_8365)
	);

	bfr new_net_8367_bfr_before (
		.din(new_net_8367),
		.dout(new_net_8366)
	);

	bfr new_net_8368_bfr_before (
		.din(new_net_8368),
		.dout(new_net_8367)
	);

	bfr new_net_8369_bfr_before (
		.din(new_net_8369),
		.dout(new_net_8368)
	);

	spl2 N367_v_fanout (
		.a(N367),
		.b(new_net_962),
		.c(new_net_8369)
	);

	bfr new_net_8370_bfr_before (
		.din(new_net_8370),
		.dout(new_net_2046)
	);

	bfr new_net_8371_bfr_before (
		.din(new_net_8371),
		.dout(new_net_8370)
	);

	spl2 N343_v_fanout (
		.a(N343),
		.b(new_net_1580),
		.c(new_net_8371)
	);

	bfr new_net_8372_bfr_before (
		.din(new_net_8372),
		.dout(new_net_2025)
	);

	spl4L N263_v_fanout (
		.a(N263),
		.b(new_net_8372),
		.c(new_net_1468),
		.d(new_net_1466),
		.e(new_net_1464)
	);

	bfr new_net_8373_bfr_before (
		.din(new_net_8373),
		.dout(new_net_2044)
	);

	bfr new_net_8374_bfr_before (
		.din(new_net_8374),
		.dout(new_net_8373)
	);

	spl2 N334_v_fanout (
		.a(N334),
		.b(new_net_1480),
		.c(new_net_8374)
	);

	bfr new_net_8375_bfr_after (
		.din(N286),
		.dout(new_net_8375)
	);

	bfr new_net_8376_bfr_after (
		.din(new_net_8375),
		.dout(new_net_8376)
	);

	bfr new_net_8377_bfr_after (
		.din(new_net_8376),
		.dout(new_net_8377)
	);

	bfr new_net_8378_bfr_before (
		.din(new_net_8378),
		.dout(new_net_2029)
	);

	bfr new_net_8379_bfr_before (
		.din(new_net_8379),
		.dout(new_net_8378)
	);

	bfr new_net_8380_bfr_before (
		.din(new_net_8380),
		.dout(new_net_8379)
	);

	spl2 N286_v_fanout (
		.a(new_net_8377),
		.b(new_net_8380),
		.c(new_net_1457)
	);

	bfr new_net_8381_bfr_after (
		.din(N251),
		.dout(new_net_8381)
	);

	bfr new_net_8382_bfr_after (
		.din(new_net_8381),
		.dout(new_net_8382)
	);

	bfr new_net_8383_bfr_after (
		.din(new_net_8382),
		.dout(new_net_8383)
	);

	bfr new_net_8384_bfr_before (
		.din(new_net_8384),
		.dout(new_net_2021)
	);

	bfr new_net_8385_bfr_before (
		.din(new_net_8385),
		.dout(new_net_8384)
	);

	bfr new_net_8386_bfr_before (
		.din(new_net_8386),
		.dout(new_net_8385)
	);

	spl2 N251_v_fanout (
		.a(new_net_8383),
		.b(new_net_8386),
		.c(new_net_946)
	);

	bfr new_net_8387_bfr_after (
		.din(N293),
		.dout(new_net_8387)
	);

	bfr new_net_8388_bfr_after (
		.din(new_net_8387),
		.dout(new_net_8388)
	);

	bfr new_net_8389_bfr_after (
		.din(new_net_8388),
		.dout(new_net_8389)
	);

	bfr new_net_8390_bfr_before (
		.din(new_net_8390),
		.dout(new_net_2031)
	);

	bfr new_net_8391_bfr_before (
		.din(new_net_8391),
		.dout(new_net_8390)
	);

	bfr new_net_8392_bfr_before (
		.din(new_net_8392),
		.dout(new_net_8391)
	);

	spl2 N293_v_fanout (
		.a(new_net_8389),
		.b(new_net_8392),
		.c(new_net_1765)
	);

	bfr new_net_8393_bfr_after (
		.din(N337),
		.dout(new_net_8393)
	);

	bfr new_net_8394_bfr_after (
		.din(new_net_8393),
		.dout(new_net_8394)
	);

	bfr new_net_8395_bfr_after (
		.din(new_net_8394),
		.dout(new_net_8395)
	);

	bfr new_net_8396_bfr_before (
		.din(new_net_8396),
		.dout(N556)
	);

	bfr new_net_8397_bfr_before (
		.din(new_net_8397),
		.dout(new_net_8396)
	);

	bfr new_net_8398_bfr_before (
		.din(new_net_8398),
		.dout(new_net_8397)
	);

	bfr new_net_8399_bfr_before (
		.din(new_net_8399),
		.dout(new_net_8398)
	);

	bfr new_net_8400_bfr_before (
		.din(new_net_8400),
		.dout(new_net_8399)
	);

	bfr new_net_8401_bfr_before (
		.din(new_net_8401),
		.dout(new_net_8400)
	);

	bfr new_net_8402_bfr_before (
		.din(new_net_8402),
		.dout(new_net_8401)
	);

	bfr new_net_8403_bfr_before (
		.din(new_net_8403),
		.dout(new_net_8402)
	);

	bfr new_net_8404_bfr_before (
		.din(new_net_8404),
		.dout(new_net_8403)
	);

	bfr new_net_8405_bfr_before (
		.din(new_net_8405),
		.dout(new_net_8404)
	);

	bfr new_net_8406_bfr_before (
		.din(new_net_8406),
		.dout(new_net_8405)
	);

	bfr new_net_8407_bfr_before (
		.din(new_net_8407),
		.dout(new_net_8406)
	);

	bfr new_net_8408_bfr_before (
		.din(new_net_8408),
		.dout(new_net_8407)
	);

	bfr new_net_8409_bfr_before (
		.din(new_net_8409),
		.dout(new_net_8408)
	);

	bfr new_net_8410_bfr_before (
		.din(new_net_8410),
		.dout(new_net_8409)
	);

	bfr new_net_8411_bfr_before (
		.din(new_net_8411),
		.dout(new_net_8410)
	);

	bfr new_net_8412_bfr_before (
		.din(new_net_8412),
		.dout(new_net_8411)
	);

	bfr new_net_8413_bfr_before (
		.din(new_net_8413),
		.dout(new_net_8412)
	);

	bfr new_net_8414_bfr_before (
		.din(new_net_8414),
		.dout(new_net_8413)
	);

	bfr new_net_8415_bfr_before (
		.din(new_net_8415),
		.dout(new_net_8414)
	);

	bfr new_net_8416_bfr_before (
		.din(new_net_8416),
		.dout(new_net_8415)
	);

	bfr new_net_8417_bfr_before (
		.din(new_net_8417),
		.dout(new_net_8416)
	);

	bfr new_net_8418_bfr_before (
		.din(new_net_8418),
		.dout(new_net_8417)
	);

	bfr new_net_8419_bfr_before (
		.din(new_net_8419),
		.dout(new_net_8418)
	);

	bfr new_net_8420_bfr_before (
		.din(new_net_8420),
		.dout(new_net_8419)
	);

	bfr new_net_8421_bfr_before (
		.din(new_net_8421),
		.dout(new_net_8420)
	);

	bfr new_net_8422_bfr_before (
		.din(new_net_8422),
		.dout(new_net_8421)
	);

	bfr new_net_8423_bfr_before (
		.din(new_net_8423),
		.dout(new_net_8422)
	);

	bfr new_net_8424_bfr_before (
		.din(new_net_8424),
		.dout(new_net_8423)
	);

	bfr new_net_8425_bfr_before (
		.din(new_net_8425),
		.dout(new_net_8424)
	);

	bfr new_net_8426_bfr_before (
		.din(new_net_8426),
		.dout(new_net_8425)
	);

	bfr new_net_8427_bfr_before (
		.din(new_net_8427),
		.dout(new_net_8426)
	);

	bfr new_net_8428_bfr_before (
		.din(new_net_8428),
		.dout(new_net_8427)
	);

	bfr new_net_8429_bfr_before (
		.din(new_net_8429),
		.dout(new_net_8428)
	);

	bfr new_net_8430_bfr_before (
		.din(new_net_8430),
		.dout(new_net_8429)
	);

	bfr new_net_8431_bfr_before (
		.din(new_net_8431),
		.dout(new_net_8430)
	);

	bfr new_net_8432_bfr_before (
		.din(new_net_8432),
		.dout(new_net_8431)
	);

	bfr new_net_8433_bfr_before (
		.din(new_net_8433),
		.dout(new_net_8432)
	);

	bfr new_net_8434_bfr_before (
		.din(new_net_8434),
		.dout(new_net_8433)
	);

	bfr new_net_8435_bfr_before (
		.din(new_net_8435),
		.dout(new_net_8434)
	);

	bfr new_net_8436_bfr_before (
		.din(new_net_8436),
		.dout(new_net_8435)
	);

	bfr new_net_8437_bfr_before (
		.din(new_net_8437),
		.dout(new_net_8436)
	);

	bfr new_net_8438_bfr_before (
		.din(new_net_8438),
		.dout(new_net_8437)
	);

	bfr new_net_8439_bfr_before (
		.din(new_net_8439),
		.dout(new_net_8438)
	);

	bfr new_net_8440_bfr_before (
		.din(new_net_8440),
		.dout(new_net_8439)
	);

	bfr new_net_8441_bfr_before (
		.din(new_net_8441),
		.dout(new_net_8440)
	);

	bfr new_net_8442_bfr_before (
		.din(new_net_8442),
		.dout(new_net_8441)
	);

	bfr new_net_8443_bfr_before (
		.din(new_net_8443),
		.dout(new_net_8442)
	);

	bfr new_net_8444_bfr_before (
		.din(new_net_8444),
		.dout(new_net_8443)
	);

	bfr new_net_8445_bfr_before (
		.din(new_net_8445),
		.dout(new_net_8444)
	);

	bfr new_net_8446_bfr_before (
		.din(new_net_8446),
		.dout(new_net_8445)
	);

	bfr new_net_8447_bfr_before (
		.din(new_net_8447),
		.dout(new_net_8446)
	);

	bfr new_net_8448_bfr_before (
		.din(new_net_8448),
		.dout(new_net_8447)
	);

	bfr new_net_8449_bfr_before (
		.din(new_net_8449),
		.dout(new_net_8448)
	);

	bfr new_net_8450_bfr_before (
		.din(new_net_8450),
		.dout(new_net_8449)
	);

	bfr new_net_8451_bfr_before (
		.din(new_net_8451),
		.dout(new_net_8450)
	);

	bfr new_net_8452_bfr_before (
		.din(new_net_8452),
		.dout(new_net_8451)
	);

	bfr new_net_8453_bfr_before (
		.din(new_net_8453),
		.dout(new_net_8452)
	);

	bfr new_net_8454_bfr_before (
		.din(new_net_8454),
		.dout(new_net_8453)
	);

	bfr new_net_8455_bfr_before (
		.din(new_net_8455),
		.dout(new_net_8454)
	);

	bfr new_net_8456_bfr_before (
		.din(new_net_8456),
		.dout(new_net_8455)
	);

	bfr new_net_8457_bfr_before (
		.din(new_net_8457),
		.dout(new_net_8456)
	);

	spl2 N337_v_fanout (
		.a(new_net_8395),
		.b(new_net_8457),
		.c(new_net_1590)
	);

	bfr new_net_8458_bfr_before (
		.din(new_net_8458),
		.dout(new_net_1790)
	);

	bfr new_net_8459_bfr_before (
		.din(new_net_8459),
		.dout(new_net_8458)
	);

	spl4L N382_v_fanout (
		.a(N382),
		.b(new_net_1789),
		.c(new_net_1788),
		.d(new_net_8459),
		.e(new_net_1787)
	);

	bfr new_net_8460_bfr_before (
		.din(new_net_8460),
		.dout(new_net_2052)
	);

	bfr new_net_8461_bfr_before (
		.din(new_net_8461),
		.dout(new_net_8460)
	);

	spl2 N361_v_fanout (
		.a(N361),
		.b(new_net_1720),
		.c(new_net_8461)
	);

	spl3L N18_v_fanout (
		.a(N18),
		.b(new_net_1977),
		.c(new_net_1963),
		.d(new_net_1998)
	);

	bfr new_net_8462_bfr_before (
		.din(new_net_8462),
		.dout(new_net_1257)
	);

	bfr new_net_8463_bfr_before (
		.din(new_net_8463),
		.dout(new_net_8462)
	);

	bfr new_net_8464_bfr_before (
		.din(new_net_8464),
		.dout(new_net_8463)
	);

	spl2 N70_v_fanout (
		.a(N70),
		.b(new_net_1258),
		.c(new_net_8464)
	);

	bfr new_net_8465_bfr_before (
		.din(new_net_8465),
		.dout(new_net_2028)
	);

	bfr new_net_8466_bfr_before (
		.din(new_net_8466),
		.dout(new_net_8465)
	);

	spl2 N283_v_fanout (
		.a(N283),
		.b(new_net_1341),
		.c(new_net_8466)
	);

	bfr new_net_8467_bfr_before (
		.din(new_net_8467),
		.dout(new_net_1961)
	);

	bfr new_net_8468_bfr_before (
		.din(new_net_8468),
		.dout(new_net_8467)
	);

	bfr new_net_8469_bfr_before (
		.din(new_net_8469),
		.dout(new_net_8468)
	);

	bfr new_net_8470_bfr_before (
		.din(new_net_8470),
		.dout(new_net_8469)
	);

	bfr new_net_8471_bfr_before (
		.din(new_net_8471),
		.dout(new_net_8470)
	);

	bfr new_net_8472_bfr_before (
		.din(new_net_8472),
		.dout(new_net_8471)
	);

	bfr new_net_8473_bfr_before (
		.din(new_net_8473),
		.dout(new_net_8472)
	);

	bfr new_net_8474_bfr_before (
		.din(new_net_8474),
		.dout(new_net_8473)
	);

	bfr new_net_8475_bfr_before (
		.din(new_net_8475),
		.dout(new_net_8474)
	);

	bfr new_net_8476_bfr_before (
		.din(new_net_8476),
		.dout(new_net_8475)
	);

	bfr new_net_8477_bfr_before (
		.din(new_net_8477),
		.dout(new_net_8476)
	);

	bfr new_net_8478_bfr_before (
		.din(new_net_8478),
		.dout(new_net_8477)
	);

	bfr new_net_8479_bfr_before (
		.din(new_net_8479),
		.dout(new_net_8478)
	);

	bfr new_net_8480_bfr_before (
		.din(new_net_8480),
		.dout(new_net_8479)
	);

	bfr new_net_8481_bfr_before (
		.din(new_net_8481),
		.dout(new_net_8480)
	);

	bfr new_net_8482_bfr_before (
		.din(new_net_8482),
		.dout(new_net_8481)
	);

	bfr new_net_8483_bfr_before (
		.din(new_net_8483),
		.dout(new_net_8482)
	);

	bfr new_net_8484_bfr_before (
		.din(new_net_8484),
		.dout(new_net_8483)
	);

	bfr new_net_8485_bfr_before (
		.din(new_net_8485),
		.dout(new_net_8484)
	);

	bfr new_net_8486_bfr_before (
		.din(new_net_8486),
		.dout(new_net_8485)
	);

	bfr new_net_8487_bfr_before (
		.din(new_net_8487),
		.dout(new_net_8486)
	);

	bfr new_net_8488_bfr_before (
		.din(new_net_8488),
		.dout(new_net_8487)
	);

	bfr new_net_8489_bfr_before (
		.din(new_net_8489),
		.dout(new_net_8488)
	);

	bfr new_net_8490_bfr_before (
		.din(new_net_8490),
		.dout(new_net_8489)
	);

	bfr new_net_8491_bfr_before (
		.din(new_net_8491),
		.dout(new_net_8490)
	);

	bfr new_net_8492_bfr_before (
		.din(new_net_8492),
		.dout(new_net_8491)
	);

	bfr new_net_8493_bfr_before (
		.din(new_net_8493),
		.dout(new_net_8492)
	);

	bfr new_net_8494_bfr_before (
		.din(new_net_8494),
		.dout(new_net_8493)
	);

	bfr new_net_8495_bfr_before (
		.din(new_net_8495),
		.dout(new_net_8494)
	);

	bfr new_net_8496_bfr_before (
		.din(new_net_8496),
		.dout(new_net_8495)
	);

	bfr new_net_8497_bfr_before (
		.din(new_net_8497),
		.dout(new_net_8496)
	);

	bfr new_net_8498_bfr_before (
		.din(new_net_8498),
		.dout(new_net_8497)
	);

	bfr new_net_8499_bfr_before (
		.din(new_net_8499),
		.dout(new_net_8498)
	);

	bfr new_net_8500_bfr_before (
		.din(new_net_8500),
		.dout(new_net_8499)
	);

	bfr new_net_8501_bfr_before (
		.din(new_net_8501),
		.dout(new_net_8500)
	);

	bfr new_net_8502_bfr_before (
		.din(new_net_8502),
		.dout(new_net_8501)
	);

	bfr new_net_8503_bfr_before (
		.din(new_net_8503),
		.dout(new_net_8502)
	);

	bfr new_net_8504_bfr_before (
		.din(new_net_8504),
		.dout(new_net_8503)
	);

	bfr new_net_8505_bfr_before (
		.din(new_net_8505),
		.dout(new_net_8504)
	);

	bfr new_net_8506_bfr_before (
		.din(new_net_8506),
		.dout(new_net_8505)
	);

	bfr new_net_8507_bfr_before (
		.din(new_net_8507),
		.dout(new_net_8506)
	);

	bfr new_net_8508_bfr_before (
		.din(new_net_8508),
		.dout(new_net_8507)
	);

	bfr new_net_8509_bfr_before (
		.din(new_net_8509),
		.dout(new_net_8508)
	);

	bfr new_net_8510_bfr_before (
		.din(new_net_8510),
		.dout(new_net_8509)
	);

	bfr new_net_8511_bfr_before (
		.din(new_net_8511),
		.dout(new_net_8510)
	);

	bfr new_net_8512_bfr_before (
		.din(new_net_8512),
		.dout(new_net_8511)
	);

	bfr new_net_8513_bfr_before (
		.din(new_net_8513),
		.dout(new_net_8512)
	);

	bfr new_net_8514_bfr_before (
		.din(new_net_8514),
		.dout(new_net_8513)
	);

	bfr new_net_8515_bfr_before (
		.din(new_net_8515),
		.dout(new_net_8514)
	);

	bfr new_net_8516_bfr_before (
		.din(new_net_8516),
		.dout(new_net_8515)
	);

	bfr new_net_8517_bfr_before (
		.din(new_net_8517),
		.dout(new_net_8516)
	);

	bfr new_net_8518_bfr_before (
		.din(new_net_8518),
		.dout(new_net_8517)
	);

	bfr new_net_8519_bfr_before (
		.din(new_net_8519),
		.dout(new_net_8518)
	);

	bfr new_net_8520_bfr_before (
		.din(new_net_8520),
		.dout(new_net_8519)
	);

	bfr new_net_8521_bfr_before (
		.din(new_net_8521),
		.dout(new_net_8520)
	);

	bfr new_net_8522_bfr_before (
		.din(new_net_8522),
		.dout(new_net_8521)
	);

	bfr new_net_8523_bfr_before (
		.din(new_net_8523),
		.dout(new_net_8522)
	);

	bfr new_net_8524_bfr_before (
		.din(new_net_8524),
		.dout(new_net_8523)
	);

	bfr new_net_8525_bfr_before (
		.din(new_net_8525),
		.dout(new_net_8524)
	);

	bfr new_net_8526_bfr_before (
		.din(new_net_8526),
		.dout(new_net_8525)
	);

	bfr new_net_8527_bfr_before (
		.din(new_net_8527),
		.dout(new_net_8526)
	);

	bfr new_net_8528_bfr_before (
		.din(new_net_8528),
		.dout(new_net_8527)
	);

	bfr new_net_8529_bfr_before (
		.din(new_net_8529),
		.dout(new_net_8528)
	);

	bfr new_net_8530_bfr_before (
		.din(new_net_8530),
		.dout(new_net_8529)
	);

	spl2 N1_v_fanout (
		.a(N1),
		.b(new_net_8530),
		.c(new_net_573)
	);

	bfr new_net_8531_bfr_after (
		.din(N274),
		.dout(new_net_8531)
	);

	bfr new_net_8532_bfr_after (
		.din(new_net_8531),
		.dout(new_net_8532)
	);

	bfr new_net_8533_bfr_after (
		.din(new_net_8532),
		.dout(new_net_8533)
	);

	bfr new_net_8534_bfr_before (
		.din(new_net_8534),
		.dout(N501)
	);

	bfr new_net_8535_bfr_before (
		.din(new_net_8535),
		.dout(new_net_8534)
	);

	bfr new_net_8536_bfr_before (
		.din(new_net_8536),
		.dout(new_net_8535)
	);

	bfr new_net_8537_bfr_before (
		.din(new_net_8537),
		.dout(new_net_8536)
	);

	bfr new_net_8538_bfr_before (
		.din(new_net_8538),
		.dout(new_net_8537)
	);

	bfr new_net_8539_bfr_before (
		.din(new_net_8539),
		.dout(new_net_8538)
	);

	bfr new_net_8540_bfr_before (
		.din(new_net_8540),
		.dout(new_net_8539)
	);

	bfr new_net_8541_bfr_before (
		.din(new_net_8541),
		.dout(new_net_8540)
	);

	bfr new_net_8542_bfr_before (
		.din(new_net_8542),
		.dout(new_net_8541)
	);

	bfr new_net_8543_bfr_before (
		.din(new_net_8543),
		.dout(new_net_8542)
	);

	bfr new_net_8544_bfr_before (
		.din(new_net_8544),
		.dout(new_net_8543)
	);

	bfr new_net_8545_bfr_before (
		.din(new_net_8545),
		.dout(new_net_8544)
	);

	bfr new_net_8546_bfr_before (
		.din(new_net_8546),
		.dout(new_net_8545)
	);

	bfr new_net_8547_bfr_before (
		.din(new_net_8547),
		.dout(new_net_8546)
	);

	bfr new_net_8548_bfr_before (
		.din(new_net_8548),
		.dout(new_net_8547)
	);

	bfr new_net_8549_bfr_before (
		.din(new_net_8549),
		.dout(new_net_8548)
	);

	bfr new_net_8550_bfr_before (
		.din(new_net_8550),
		.dout(new_net_8549)
	);

	bfr new_net_8551_bfr_before (
		.din(new_net_8551),
		.dout(new_net_8550)
	);

	bfr new_net_8552_bfr_before (
		.din(new_net_8552),
		.dout(new_net_8551)
	);

	bfr new_net_8553_bfr_before (
		.din(new_net_8553),
		.dout(new_net_8552)
	);

	bfr new_net_8554_bfr_before (
		.din(new_net_8554),
		.dout(new_net_8553)
	);

	bfr new_net_8555_bfr_before (
		.din(new_net_8555),
		.dout(new_net_8554)
	);

	bfr new_net_8556_bfr_before (
		.din(new_net_8556),
		.dout(new_net_8555)
	);

	bfr new_net_8557_bfr_before (
		.din(new_net_8557),
		.dout(new_net_8556)
	);

	bfr new_net_8558_bfr_before (
		.din(new_net_8558),
		.dout(new_net_8557)
	);

	bfr new_net_8559_bfr_before (
		.din(new_net_8559),
		.dout(new_net_8558)
	);

	bfr new_net_8560_bfr_before (
		.din(new_net_8560),
		.dout(new_net_8559)
	);

	bfr new_net_8561_bfr_before (
		.din(new_net_8561),
		.dout(new_net_8560)
	);

	bfr new_net_8562_bfr_before (
		.din(new_net_8562),
		.dout(new_net_8561)
	);

	bfr new_net_8563_bfr_before (
		.din(new_net_8563),
		.dout(new_net_8562)
	);

	bfr new_net_8564_bfr_before (
		.din(new_net_8564),
		.dout(new_net_8563)
	);

	bfr new_net_8565_bfr_before (
		.din(new_net_8565),
		.dout(new_net_8564)
	);

	bfr new_net_8566_bfr_before (
		.din(new_net_8566),
		.dout(new_net_8565)
	);

	bfr new_net_8567_bfr_before (
		.din(new_net_8567),
		.dout(new_net_8566)
	);

	bfr new_net_8568_bfr_before (
		.din(new_net_8568),
		.dout(new_net_8567)
	);

	bfr new_net_8569_bfr_before (
		.din(new_net_8569),
		.dout(new_net_8568)
	);

	bfr new_net_8570_bfr_before (
		.din(new_net_8570),
		.dout(new_net_8569)
	);

	bfr new_net_8571_bfr_before (
		.din(new_net_8571),
		.dout(new_net_8570)
	);

	bfr new_net_8572_bfr_before (
		.din(new_net_8572),
		.dout(new_net_8571)
	);

	bfr new_net_8573_bfr_before (
		.din(new_net_8573),
		.dout(new_net_8572)
	);

	bfr new_net_8574_bfr_before (
		.din(new_net_8574),
		.dout(new_net_8573)
	);

	bfr new_net_8575_bfr_before (
		.din(new_net_8575),
		.dout(new_net_8574)
	);

	bfr new_net_8576_bfr_before (
		.din(new_net_8576),
		.dout(new_net_8575)
	);

	bfr new_net_8577_bfr_before (
		.din(new_net_8577),
		.dout(new_net_8576)
	);

	bfr new_net_8578_bfr_before (
		.din(new_net_8578),
		.dout(new_net_8577)
	);

	bfr new_net_8579_bfr_before (
		.din(new_net_8579),
		.dout(new_net_8578)
	);

	bfr new_net_8580_bfr_before (
		.din(new_net_8580),
		.dout(new_net_8579)
	);

	bfr new_net_8581_bfr_before (
		.din(new_net_8581),
		.dout(new_net_8580)
	);

	bfr new_net_8582_bfr_before (
		.din(new_net_8582),
		.dout(new_net_8581)
	);

	bfr new_net_8583_bfr_before (
		.din(new_net_8583),
		.dout(new_net_8582)
	);

	bfr new_net_8584_bfr_before (
		.din(new_net_8584),
		.dout(new_net_8583)
	);

	bfr new_net_8585_bfr_before (
		.din(new_net_8585),
		.dout(new_net_8584)
	);

	bfr new_net_8586_bfr_before (
		.din(new_net_8586),
		.dout(new_net_8585)
	);

	bfr new_net_8587_bfr_before (
		.din(new_net_8587),
		.dout(new_net_8586)
	);

	bfr new_net_8588_bfr_before (
		.din(new_net_8588),
		.dout(new_net_8587)
	);

	bfr new_net_8589_bfr_before (
		.din(new_net_8589),
		.dout(new_net_8588)
	);

	bfr new_net_8590_bfr_before (
		.din(new_net_8590),
		.dout(new_net_8589)
	);

	bfr new_net_8591_bfr_before (
		.din(new_net_8591),
		.dout(new_net_8590)
	);

	bfr new_net_8592_bfr_before (
		.din(new_net_8592),
		.dout(new_net_8591)
	);

	bfr new_net_8593_bfr_before (
		.din(new_net_8593),
		.dout(new_net_8592)
	);

	bfr new_net_8594_bfr_before (
		.din(new_net_8594),
		.dout(new_net_8593)
	);

	bfr new_net_8595_bfr_before (
		.din(new_net_8595),
		.dout(new_net_8594)
	);

	spl2 N274_v_fanout (
		.a(new_net_8533),
		.b(new_net_8595),
		.c(new_net_1067)
	);

	bfr new_net_8596_bfr_after (
		.din(N248),
		.dout(new_net_8596)
	);

	bfr new_net_8597_bfr_after (
		.din(new_net_8596),
		.dout(new_net_8597)
	);

	bfr new_net_8598_bfr_after (
		.din(new_net_8597),
		.dout(new_net_8598)
	);

	bfr new_net_8599_bfr_before (
		.din(new_net_8599),
		.dout(N478)
	);

	bfr new_net_8600_bfr_before (
		.din(new_net_8600),
		.dout(new_net_8599)
	);

	bfr new_net_8601_bfr_before (
		.din(new_net_8601),
		.dout(new_net_8600)
	);

	bfr new_net_8602_bfr_before (
		.din(new_net_8602),
		.dout(new_net_8601)
	);

	bfr new_net_8603_bfr_before (
		.din(new_net_8603),
		.dout(new_net_8602)
	);

	bfr new_net_8604_bfr_before (
		.din(new_net_8604),
		.dout(new_net_8603)
	);

	bfr new_net_8605_bfr_before (
		.din(new_net_8605),
		.dout(new_net_8604)
	);

	bfr new_net_8606_bfr_before (
		.din(new_net_8606),
		.dout(new_net_8605)
	);

	bfr new_net_8607_bfr_before (
		.din(new_net_8607),
		.dout(new_net_8606)
	);

	bfr new_net_8608_bfr_before (
		.din(new_net_8608),
		.dout(new_net_8607)
	);

	bfr new_net_8609_bfr_before (
		.din(new_net_8609),
		.dout(new_net_8608)
	);

	bfr new_net_8610_bfr_before (
		.din(new_net_8610),
		.dout(new_net_8609)
	);

	bfr new_net_8611_bfr_before (
		.din(new_net_8611),
		.dout(new_net_8610)
	);

	bfr new_net_8612_bfr_before (
		.din(new_net_8612),
		.dout(new_net_8611)
	);

	bfr new_net_8613_bfr_before (
		.din(new_net_8613),
		.dout(new_net_8612)
	);

	bfr new_net_8614_bfr_before (
		.din(new_net_8614),
		.dout(new_net_8613)
	);

	bfr new_net_8615_bfr_before (
		.din(new_net_8615),
		.dout(new_net_8614)
	);

	bfr new_net_8616_bfr_before (
		.din(new_net_8616),
		.dout(new_net_8615)
	);

	bfr new_net_8617_bfr_before (
		.din(new_net_8617),
		.dout(new_net_8616)
	);

	bfr new_net_8618_bfr_before (
		.din(new_net_8618),
		.dout(new_net_8617)
	);

	bfr new_net_8619_bfr_before (
		.din(new_net_8619),
		.dout(new_net_8618)
	);

	bfr new_net_8620_bfr_before (
		.din(new_net_8620),
		.dout(new_net_8619)
	);

	bfr new_net_8621_bfr_before (
		.din(new_net_8621),
		.dout(new_net_8620)
	);

	bfr new_net_8622_bfr_before (
		.din(new_net_8622),
		.dout(new_net_8621)
	);

	bfr new_net_8623_bfr_before (
		.din(new_net_8623),
		.dout(new_net_8622)
	);

	bfr new_net_8624_bfr_before (
		.din(new_net_8624),
		.dout(new_net_8623)
	);

	bfr new_net_8625_bfr_before (
		.din(new_net_8625),
		.dout(new_net_8624)
	);

	bfr new_net_8626_bfr_before (
		.din(new_net_8626),
		.dout(new_net_8625)
	);

	bfr new_net_8627_bfr_before (
		.din(new_net_8627),
		.dout(new_net_8626)
	);

	bfr new_net_8628_bfr_before (
		.din(new_net_8628),
		.dout(new_net_8627)
	);

	bfr new_net_8629_bfr_before (
		.din(new_net_8629),
		.dout(new_net_8628)
	);

	bfr new_net_8630_bfr_before (
		.din(new_net_8630),
		.dout(new_net_8629)
	);

	bfr new_net_8631_bfr_before (
		.din(new_net_8631),
		.dout(new_net_8630)
	);

	bfr new_net_8632_bfr_before (
		.din(new_net_8632),
		.dout(new_net_8631)
	);

	bfr new_net_8633_bfr_before (
		.din(new_net_8633),
		.dout(new_net_8632)
	);

	bfr new_net_8634_bfr_before (
		.din(new_net_8634),
		.dout(new_net_8633)
	);

	bfr new_net_8635_bfr_before (
		.din(new_net_8635),
		.dout(new_net_8634)
	);

	bfr new_net_8636_bfr_before (
		.din(new_net_8636),
		.dout(new_net_8635)
	);

	bfr new_net_8637_bfr_before (
		.din(new_net_8637),
		.dout(new_net_8636)
	);

	bfr new_net_8638_bfr_before (
		.din(new_net_8638),
		.dout(new_net_8637)
	);

	bfr new_net_8639_bfr_before (
		.din(new_net_8639),
		.dout(new_net_8638)
	);

	bfr new_net_8640_bfr_before (
		.din(new_net_8640),
		.dout(new_net_8639)
	);

	bfr new_net_8641_bfr_before (
		.din(new_net_8641),
		.dout(new_net_8640)
	);

	bfr new_net_8642_bfr_before (
		.din(new_net_8642),
		.dout(new_net_8641)
	);

	bfr new_net_8643_bfr_before (
		.din(new_net_8643),
		.dout(new_net_8642)
	);

	bfr new_net_8644_bfr_before (
		.din(new_net_8644),
		.dout(new_net_8643)
	);

	bfr new_net_8645_bfr_before (
		.din(new_net_8645),
		.dout(new_net_8644)
	);

	bfr new_net_8646_bfr_before (
		.din(new_net_8646),
		.dout(new_net_8645)
	);

	bfr new_net_8647_bfr_before (
		.din(new_net_8647),
		.dout(new_net_8646)
	);

	bfr new_net_8648_bfr_before (
		.din(new_net_8648),
		.dout(new_net_8647)
	);

	bfr new_net_8649_bfr_before (
		.din(new_net_8649),
		.dout(new_net_8648)
	);

	bfr new_net_8650_bfr_before (
		.din(new_net_8650),
		.dout(new_net_8649)
	);

	bfr new_net_8651_bfr_before (
		.din(new_net_8651),
		.dout(new_net_8650)
	);

	bfr new_net_8652_bfr_before (
		.din(new_net_8652),
		.dout(new_net_8651)
	);

	bfr new_net_8653_bfr_before (
		.din(new_net_8653),
		.dout(new_net_8652)
	);

	bfr new_net_8654_bfr_before (
		.din(new_net_8654),
		.dout(new_net_8653)
	);

	bfr new_net_8655_bfr_before (
		.din(new_net_8655),
		.dout(new_net_8654)
	);

	bfr new_net_8656_bfr_before (
		.din(new_net_8656),
		.dout(new_net_8655)
	);

	bfr new_net_8657_bfr_before (
		.din(new_net_8657),
		.dout(new_net_8656)
	);

	bfr new_net_8658_bfr_before (
		.din(new_net_8658),
		.dout(new_net_8657)
	);

	bfr new_net_8659_bfr_before (
		.din(new_net_8659),
		.dout(new_net_8658)
	);

	bfr new_net_8660_bfr_before (
		.din(new_net_8660),
		.dout(new_net_8659)
	);

	spl2 N248_v_fanout (
		.a(new_net_8598),
		.b(new_net_8660),
		.c(new_net_847)
	);

	bfr new_net_8661_bfr_after (
		.din(N280),
		.dout(new_net_8661)
	);

	bfr new_net_8662_bfr_after (
		.din(new_net_8661),
		.dout(new_net_8662)
	);

	bfr new_net_8663_bfr_after (
		.din(new_net_8662),
		.dout(new_net_8663)
	);

	bfr new_net_8664_bfr_before (
		.din(new_net_8664),
		.dout(new_net_2027)
	);

	bfr new_net_8665_bfr_before (
		.din(new_net_8665),
		.dout(new_net_8664)
	);

	bfr new_net_8666_bfr_before (
		.din(new_net_8666),
		.dout(new_net_8665)
	);

	spl2 N280_v_fanout (
		.a(new_net_8663),
		.b(new_net_8666),
		.c(new_net_1122)
	);

	bfr new_net_8667_bfr_after (
		.din(N316),
		.dout(new_net_8667)
	);

	bfr new_net_8668_bfr_after (
		.din(new_net_8667),
		.dout(new_net_8668)
	);

	bfr new_net_8669_bfr_after (
		.din(new_net_8668),
		.dout(new_net_8669)
	);

	bfr new_net_8670_bfr_before (
		.din(new_net_8670),
		.dout(new_net_2038)
	);

	bfr new_net_8671_bfr_before (
		.din(new_net_8671),
		.dout(new_net_8670)
	);

	bfr new_net_8672_bfr_before (
		.din(new_net_8672),
		.dout(new_net_8671)
	);

	spl2 N316_v_fanout (
		.a(new_net_8669),
		.b(new_net_1357),
		.c(new_net_8672)
	);

	spl2 N245_v_fanout (
		.a(N245),
		.b(new_net_1731),
		.c(new_net_1730)
	);

	spl2 N271_v_fanout (
		.a(N271),
		.b(new_net_1675),
		.c(new_net_1674)
	);

	bfr new_net_8673_bfr_before (
		.din(new_net_8673),
		.dout(new_net_2056)
	);

	bfr new_net_8674_bfr_before (
		.din(new_net_8674),
		.dout(new_net_8673)
	);

	spl3L N38_v_fanout (
		.a(N38),
		.b(new_net_8674),
		.c(new_net_1083),
		.d(new_net_1085)
	);

	bfr new_net_8675_bfr_after (
		.din(N26),
		.dout(new_net_8675)
	);

	bfr new_net_8676_bfr_after (
		.din(new_net_8675),
		.dout(new_net_8676)
	);

	bfr new_net_8677_bfr_after (
		.din(new_net_8676),
		.dout(new_net_8677)
	);

	bfr new_net_2195_bfr_after (
		.din(new_net_8677),
		.dout(new_net_2195)
	);

	bfr new_net_8678_bfr_after (
		.din(n_0311_),
		.dout(new_net_8678)
	);

	bfr new_net_8679_bfr_after (
		.din(new_net_8678),
		.dout(new_net_8679)
	);

	bfr new_net_8680_bfr_after (
		.din(new_net_8679),
		.dout(new_net_8680)
	);

	bfr new_net_8681_bfr_after (
		.din(new_net_8680),
		.dout(new_net_8681)
	);

	bfr new_net_8682_bfr_after (
		.din(new_net_8681),
		.dout(new_net_8682)
	);

	bfr new_net_8683_bfr_after (
		.din(new_net_8682),
		.dout(new_net_8683)
	);

	bfr new_net_8684_bfr_after (
		.din(new_net_8683),
		.dout(new_net_8684)
	);

	bfr new_net_8685_bfr_after (
		.din(new_net_8684),
		.dout(new_net_8685)
	);

	bfr new_net_8686_bfr_after (
		.din(new_net_8685),
		.dout(new_net_8686)
	);

	bfr new_net_8687_bfr_after (
		.din(new_net_8686),
		.dout(new_net_8687)
	);

	bfr new_net_2438_bfr_after (
		.din(new_net_8687),
		.dout(new_net_2438)
	);

	bfr new_net_8688_bfr_after (
		.din(new_net_2556),
		.dout(new_net_8688)
	);

	bfr new_net_8689_bfr_after (
		.din(new_net_8688),
		.dout(new_net_8689)
	);

	bfr new_net_8690_bfr_after (
		.din(new_net_8689),
		.dout(new_net_8690)
	);

	bfr new_net_8691_bfr_after (
		.din(new_net_8690),
		.dout(new_net_8691)
	);

	bfr N10715_bfr_after (
		.din(new_net_8691),
		.dout(N10715)
	);

	bfr new_net_8692_bfr_after (
		.din(N222),
		.dout(new_net_8692)
	);

	bfr new_net_8693_bfr_after (
		.din(new_net_8692),
		.dout(new_net_8693)
	);

	bfr new_net_8694_bfr_after (
		.din(new_net_8693),
		.dout(new_net_8694)
	);

	bfr new_net_2270_bfr_after (
		.din(new_net_8694),
		.dout(new_net_2270)
	);

	bfr new_net_8695_bfr_after (
		.din(N194),
		.dout(new_net_8695)
	);

	bfr new_net_8696_bfr_after (
		.din(new_net_8695),
		.dout(new_net_8696)
	);

	bfr new_net_8697_bfr_after (
		.din(new_net_8696),
		.dout(new_net_8697)
	);

	bfr new_net_2333_bfr_after (
		.din(new_net_8697),
		.dout(new_net_2333)
	);

	bfr new_net_2228_bfr_after (
		.din(n_0768_),
		.dout(new_net_2228)
	);

	bfr new_net_8698_bfr_after (
		.din(N223),
		.dout(new_net_8698)
	);

	bfr new_net_8699_bfr_after (
		.din(new_net_8698),
		.dout(new_net_8699)
	);

	bfr new_net_8700_bfr_after (
		.din(new_net_8699),
		.dout(new_net_8700)
	);

	bfr new_net_2249_bfr_after (
		.din(new_net_8700),
		.dout(new_net_2249)
	);

	bfr new_net_2207_bfr_after (
		.din(n_0734_),
		.dout(new_net_2207)
	);

	bfr new_net_2354_bfr_after (
		.din(n_1232_),
		.dout(new_net_2354)
	);

	bfr new_net_8701_bfr_after (
		.din(n_0465_),
		.dout(new_net_8701)
	);

	bfr new_net_8702_bfr_after (
		.din(new_net_8701),
		.dout(new_net_8702)
	);

	bfr new_net_8703_bfr_after (
		.din(new_net_8702),
		.dout(new_net_8703)
	);

	bfr new_net_8704_bfr_after (
		.din(new_net_8703),
		.dout(new_net_8704)
	);

	bfr new_net_8705_bfr_after (
		.din(new_net_8704),
		.dout(new_net_8705)
	);

	bfr new_net_8706_bfr_after (
		.din(new_net_8705),
		.dout(new_net_8706)
	);

	bfr new_net_8707_bfr_after (
		.din(new_net_8706),
		.dout(new_net_8707)
	);

	bfr new_net_8708_bfr_after (
		.din(new_net_8707),
		.dout(new_net_8708)
	);

	bfr new_net_8709_bfr_after (
		.din(new_net_8708),
		.dout(new_net_8709)
	);

	bfr new_net_8710_bfr_after (
		.din(new_net_8709),
		.dout(new_net_8710)
	);

	bfr new_net_8711_bfr_after (
		.din(new_net_8710),
		.dout(new_net_8711)
	);

	bfr new_net_8712_bfr_after (
		.din(new_net_8711),
		.dout(new_net_8712)
	);

	bfr new_net_8713_bfr_after (
		.din(new_net_8712),
		.dout(new_net_8713)
	);

	bfr new_net_8714_bfr_after (
		.din(new_net_8713),
		.dout(new_net_8714)
	);

	bfr new_net_8715_bfr_after (
		.din(new_net_8714),
		.dout(new_net_8715)
	);

	bfr new_net_8716_bfr_after (
		.din(new_net_8715),
		.dout(new_net_8716)
	);

	bfr new_net_8717_bfr_after (
		.din(new_net_8716),
		.dout(new_net_8717)
	);

	bfr new_net_8718_bfr_after (
		.din(new_net_8717),
		.dout(new_net_8718)
	);

	bfr new_net_8719_bfr_after (
		.din(new_net_8718),
		.dout(new_net_8719)
	);

	bfr new_net_8720_bfr_after (
		.din(new_net_8719),
		.dout(new_net_8720)
	);

	bfr new_net_8721_bfr_after (
		.din(new_net_8720),
		.dout(new_net_8721)
	);

	bfr new_net_2459_bfr_after (
		.din(new_net_8721),
		.dout(new_net_2459)
	);

	bfr new_net_8722_bfr_after (
		.din(n_0610_),
		.dout(new_net_8722)
	);

	bfr new_net_2480_bfr_after (
		.din(new_net_8722),
		.dout(new_net_2480)
	);

	bfr new_net_8723_bfr_after (
		.din(N75),
		.dout(new_net_8723)
	);

	bfr new_net_8724_bfr_after (
		.din(new_net_8723),
		.dout(new_net_8724)
	);

	bfr new_net_8725_bfr_after (
		.din(new_net_8724),
		.dout(new_net_8725)
	);

	bfr new_net_2291_bfr_after (
		.din(new_net_8725),
		.dout(new_net_2291)
	);

	bfr new_net_8726_bfr_after (
		.din(N202),
		.dout(new_net_8726)
	);

	bfr new_net_8727_bfr_after (
		.din(new_net_8726),
		.dout(new_net_8727)
	);

	bfr new_net_8728_bfr_after (
		.din(new_net_8727),
		.dout(new_net_8728)
	);

	bfr new_net_2375_bfr_after (
		.din(new_net_8728),
		.dout(new_net_2375)
	);

	bfr new_net_8729_bfr_after (
		.din(new_net_2495),
		.dout(new_net_8729)
	);

	bfr new_net_8730_bfr_after (
		.din(new_net_8729),
		.dout(new_net_8730)
	);

	bfr new_net_8731_bfr_after (
		.din(new_net_8730),
		.dout(new_net_8731)
	);

	bfr new_net_8732_bfr_after (
		.din(new_net_8731),
		.dout(new_net_8732)
	);

	bfr new_net_8733_bfr_after (
		.din(new_net_8732),
		.dout(new_net_8733)
	);

	bfr new_net_8734_bfr_after (
		.din(new_net_8733),
		.dout(new_net_8734)
	);

	bfr new_net_8735_bfr_after (
		.din(new_net_8734),
		.dout(new_net_8735)
	);

	bfr new_net_8736_bfr_after (
		.din(new_net_8735),
		.dout(new_net_8736)
	);

	bfr new_net_8737_bfr_after (
		.din(new_net_8736),
		.dout(new_net_8737)
	);

	bfr new_net_8738_bfr_after (
		.din(new_net_8737),
		.dout(new_net_8738)
	);

	bfr new_net_8739_bfr_after (
		.din(new_net_8738),
		.dout(new_net_8739)
	);

	bfr new_net_8740_bfr_after (
		.din(new_net_8739),
		.dout(new_net_8740)
	);

	bfr new_net_8741_bfr_after (
		.din(new_net_8740),
		.dout(new_net_8741)
	);

	bfr new_net_8742_bfr_after (
		.din(new_net_8741),
		.dout(new_net_8742)
	);

	bfr new_net_8743_bfr_after (
		.din(new_net_8742),
		.dout(new_net_8743)
	);

	bfr new_net_8744_bfr_after (
		.din(new_net_8743),
		.dout(new_net_8744)
	);

	bfr N10714_bfr_after (
		.din(new_net_8744),
		.dout(N10714)
	);

	bfr new_net_8745_bfr_after (
		.din(N50),
		.dout(new_net_8745)
	);

	bfr new_net_8746_bfr_after (
		.din(new_net_8745),
		.dout(new_net_8746)
	);

	bfr new_net_8747_bfr_after (
		.din(new_net_8746),
		.dout(new_net_8747)
	);

	bfr new_net_2265_bfr_after (
		.din(new_net_8747),
		.dout(new_net_2265)
	);

	bfr new_net_8748_bfr_after (
		.din(N109),
		.dout(new_net_8748)
	);

	bfr new_net_8749_bfr_after (
		.din(new_net_8748),
		.dout(new_net_8749)
	);

	bfr new_net_8750_bfr_after (
		.din(new_net_8749),
		.dout(new_net_8750)
	);

	bfr new_net_2307_bfr_after (
		.din(new_net_8750),
		.dout(new_net_2307)
	);

	bfr new_net_2391_bfr_after (
		.din(N163),
		.dout(new_net_2391)
	);

	bfr new_net_8751_bfr_after (
		.din(n_0240_),
		.dout(new_net_8751)
	);

	bfr new_net_8752_bfr_after (
		.din(new_net_8751),
		.dout(new_net_8752)
	);

	bfr new_net_2412_bfr_after (
		.din(new_net_8752),
		.dout(new_net_2412)
	);

	bfr new_net_8753_bfr_after (
		.din(N153),
		.dout(new_net_8753)
	);

	bfr new_net_8754_bfr_after (
		.din(new_net_8753),
		.dout(new_net_8754)
	);

	bfr new_net_8755_bfr_after (
		.din(new_net_8754),
		.dout(new_net_8755)
	);

	bfr new_net_2202_bfr_after (
		.din(new_net_8755),
		.dout(new_net_2202)
	);

	bfr new_net_8756_bfr_after (
		.din(N213),
		.dout(new_net_8756)
	);

	bfr new_net_8757_bfr_after (
		.din(new_net_8756),
		.dout(new_net_8757)
	);

	bfr new_net_8758_bfr_after (
		.din(new_net_8757),
		.dout(new_net_8758)
	);

	bfr new_net_2223_bfr_after (
		.din(new_net_8758),
		.dout(new_net_2223)
	);

	bfr new_net_8759_bfr_after (
		.din(N44),
		.dout(new_net_8759)
	);

	bfr new_net_8760_bfr_after (
		.din(new_net_8759),
		.dout(new_net_8760)
	);

	bfr new_net_8761_bfr_after (
		.din(new_net_8760),
		.dout(new_net_8761)
	);

	bfr new_net_2244_bfr_after (
		.din(new_net_8761),
		.dout(new_net_2244)
	);

	bfr new_net_8762_bfr_after (
		.din(N76),
		.dout(new_net_8762)
	);

	bfr new_net_8763_bfr_after (
		.din(new_net_8762),
		.dout(new_net_8763)
	);

	bfr new_net_8764_bfr_after (
		.din(new_net_8763),
		.dout(new_net_8764)
	);

	bfr new_net_2286_bfr_after (
		.din(new_net_8764),
		.dout(new_net_2286)
	);

	bfr new_net_2328_bfr_after (
		.din(n_1159_),
		.dout(new_net_2328)
	);

	bfr new_net_8765_bfr_after (
		.din(N175),
		.dout(new_net_8765)
	);

	bfr new_net_8766_bfr_after (
		.din(new_net_8765),
		.dout(new_net_8766)
	);

	bfr new_net_8767_bfr_after (
		.din(new_net_8766),
		.dout(new_net_8767)
	);

	bfr new_net_2349_bfr_after (
		.din(new_net_8767),
		.dout(new_net_2349)
	);

	bfr new_net_8768_bfr_after (
		.din(new_net_2527),
		.dout(new_net_8768)
	);

	bfr new_net_8769_bfr_after (
		.din(new_net_8768),
		.dout(new_net_8769)
	);

	bfr new_net_8770_bfr_after (
		.din(new_net_8769),
		.dout(new_net_8770)
	);

	bfr new_net_8771_bfr_after (
		.din(new_net_8770),
		.dout(new_net_8771)
	);

	bfr new_net_8772_bfr_after (
		.din(new_net_8771),
		.dout(new_net_8772)
	);

	bfr new_net_8773_bfr_after (
		.din(new_net_8772),
		.dout(new_net_8773)
	);

	bfr new_net_8774_bfr_after (
		.din(new_net_8773),
		.dout(new_net_8774)
	);

	bfr new_net_8775_bfr_after (
		.din(new_net_8774),
		.dout(new_net_8775)
	);

	bfr new_net_8776_bfr_after (
		.din(new_net_8775),
		.dout(new_net_8776)
	);

	bfr new_net_8777_bfr_after (
		.din(new_net_8776),
		.dout(new_net_8777)
	);

	bfr new_net_8778_bfr_after (
		.din(new_net_8777),
		.dout(new_net_8778)
	);

	bfr new_net_8779_bfr_after (
		.din(new_net_8778),
		.dout(new_net_8779)
	);

	bfr new_net_8780_bfr_after (
		.din(new_net_8779),
		.dout(new_net_8780)
	);

	bfr N11333_bfr_after (
		.din(new_net_8780),
		.dout(N11333)
	);

	bfr new_net_2251_bfr_after (
		.din(n_0849_),
		.dout(new_net_2251)
	);

	bfr new_net_8781_bfr_after (
		.din(N113),
		.dout(new_net_8781)
	);

	bfr new_net_8782_bfr_after (
		.din(new_net_8781),
		.dout(new_net_8782)
	);

	bfr new_net_8783_bfr_after (
		.din(new_net_8782),
		.dout(new_net_8783)
	);

	bfr new_net_2277_bfr_after (
		.din(new_net_8783),
		.dout(new_net_2277)
	);

	bfr new_net_2340_bfr_after (
		.din(n_1186_),
		.dout(new_net_2340)
	);

	bfr new_net_8784_bfr_after (
		.din(N160),
		.dout(new_net_8784)
	);

	bfr new_net_8785_bfr_after (
		.din(new_net_8784),
		.dout(new_net_8785)
	);

	bfr new_net_8786_bfr_after (
		.din(new_net_8785),
		.dout(new_net_8786)
	);

	bfr new_net_2216_bfr_after (
		.din(new_net_8786),
		.dout(new_net_2216)
	);

	bfr new_net_2260_bfr_after (
		.din(n_0867_),
		.dout(new_net_2260)
	);

	bfr new_net_8787_bfr_after (
		.din(N60),
		.dout(new_net_8787)
	);

	bfr new_net_8788_bfr_after (
		.din(new_net_8787),
		.dout(new_net_8788)
	);

	bfr new_net_8789_bfr_after (
		.din(new_net_8788),
		.dout(new_net_8789)
	);

	bfr new_net_2302_bfr_after (
		.din(new_net_8789),
		.dout(new_net_2302)
	);

	bfr new_net_8790_bfr_after (
		.din(n_0068_),
		.dout(new_net_8790)
	);

	bfr new_net_8791_bfr_after (
		.din(new_net_8790),
		.dout(new_net_8791)
	);

	bfr new_net_8792_bfr_after (
		.din(new_net_8791),
		.dout(new_net_8792)
	);

	bfr new_net_8793_bfr_after (
		.din(new_net_8792),
		.dout(new_net_8793)
	);

	bfr new_net_8794_bfr_after (
		.din(new_net_8793),
		.dout(new_net_8794)
	);

	bfr new_net_8795_bfr_after (
		.din(new_net_8794),
		.dout(new_net_8795)
	);

	bfr new_net_8796_bfr_after (
		.din(new_net_8795),
		.dout(new_net_8796)
	);

	bfr new_net_8797_bfr_after (
		.din(new_net_8796),
		.dout(new_net_8797)
	);

	bfr new_net_8798_bfr_after (
		.din(new_net_8797),
		.dout(new_net_8798)
	);

	bfr new_net_8799_bfr_after (
		.din(new_net_8798),
		.dout(new_net_8799)
	);

	bfr new_net_8800_bfr_after (
		.din(new_net_8799),
		.dout(new_net_8800)
	);

	bfr new_net_8801_bfr_after (
		.din(new_net_8800),
		.dout(new_net_8801)
	);

	bfr new_net_8802_bfr_after (
		.din(new_net_8801),
		.dout(new_net_8802)
	);

	bfr new_net_8803_bfr_after (
		.din(new_net_8802),
		.dout(new_net_8803)
	);

	bfr new_net_8804_bfr_after (
		.din(new_net_8803),
		.dout(new_net_8804)
	);

	bfr new_net_8805_bfr_after (
		.din(new_net_8804),
		.dout(new_net_8805)
	);

	bfr new_net_8806_bfr_after (
		.din(new_net_8805),
		.dout(new_net_8806)
	);

	bfr new_net_8807_bfr_after (
		.din(new_net_8806),
		.dout(new_net_8807)
	);

	bfr new_net_2386_bfr_after (
		.din(new_net_8807),
		.dout(new_net_2386)
	);

	bfr new_net_2407_bfr_after (
		.din(n_0225_),
		.dout(new_net_2407)
	);

	bfr new_net_8808_bfr_after (
		.din(N87),
		.dout(new_net_8808)
	);

	bfr new_net_8809_bfr_after (
		.din(new_net_8808),
		.dout(new_net_8809)
	);

	bfr new_net_8810_bfr_after (
		.din(new_net_8809),
		.dout(new_net_8810)
	);

	bfr new_net_2281_bfr_after (
		.din(new_net_8810),
		.dout(new_net_2281)
	);

	bfr new_net_8811_bfr_after (
		.din(N195),
		.dout(new_net_8811)
	);

	bfr new_net_8812_bfr_after (
		.din(new_net_8811),
		.dout(new_net_8812)
	);

	bfr new_net_8813_bfr_after (
		.din(new_net_8812),
		.dout(new_net_8813)
	);

	bfr new_net_2323_bfr_after (
		.din(new_net_8813),
		.dout(new_net_2323)
	);

	bfr new_net_8814_bfr_after (
		.din(N171),
		.dout(new_net_8814)
	);

	bfr new_net_8815_bfr_after (
		.din(new_net_8814),
		.dout(new_net_8815)
	);

	bfr new_net_8816_bfr_after (
		.din(new_net_8815),
		.dout(new_net_8816)
	);

	bfr new_net_2344_bfr_after (
		.din(new_net_8816),
		.dout(new_net_2344)
	);

	bfr new_net_2239_bfr_after (
		.din(n_0822_),
		.dout(new_net_2239)
	);

	bfr new_net_2187_bfr_after (
		.din(n_0669_),
		.dout(new_net_2187)
	);

	bfr new_net_8817_bfr_after (
		.din(N238),
		.dout(new_net_8817)
	);

	bfr new_net_8818_bfr_after (
		.din(new_net_8817),
		.dout(new_net_8818)
	);

	bfr new_net_8819_bfr_after (
		.din(new_net_8818),
		.dout(new_net_8819)
	);

	bfr new_net_2197_bfr_after (
		.din(new_net_8819),
		.dout(new_net_2197)
	);

	bfr new_net_2370_bfr_after (
		.din(n_1272_),
		.dout(new_net_2370)
	);

	bfr new_net_2433_bfr_after (
		.din(n_0303_),
		.dout(new_net_2433)
	);

	bfr new_net_8820_bfr_after (
		.din(N47),
		.dout(new_net_8820)
	);

	bfr new_net_8821_bfr_after (
		.din(new_net_8820),
		.dout(new_net_8821)
	);

	bfr new_net_8822_bfr_after (
		.din(new_net_8821),
		.dout(new_net_8822)
	);

	bfr new_net_2250_bfr_after (
		.din(new_net_8822),
		.dout(new_net_2250)
	);

	bfr new_net_2463_bfr_after (
		.din(n_0499_),
		.dout(new_net_2463)
	);

	bfr new_net_2458_bfr_after (
		.din(n_0455_),
		.dout(new_net_2458)
	);

	bfr new_net_2254_bfr_after (
		.din(n_0855_),
		.dout(new_net_2254)
	);

	bfr new_net_2213_bfr_after (
		.din(n_0749_),
		.dout(new_net_2213)
	);

	bfr new_net_8823_bfr_after (
		.din(N61),
		.dout(new_net_8823)
	);

	bfr new_net_8824_bfr_after (
		.din(new_net_8823),
		.dout(new_net_8824)
	);

	bfr new_net_8825_bfr_after (
		.din(new_net_8824),
		.dout(new_net_8825)
	);

	bfr new_net_2297_bfr_after (
		.din(new_net_8825),
		.dout(new_net_2297)
	);

	bfr new_net_8826_bfr_after (
		.din(n_1357_),
		.dout(new_net_8826)
	);

	bfr new_net_8827_bfr_after (
		.din(new_net_8826),
		.dout(new_net_8827)
	);

	bfr new_net_8828_bfr_after (
		.din(new_net_8827),
		.dout(new_net_8828)
	);

	bfr new_net_8829_bfr_after (
		.din(new_net_8828),
		.dout(new_net_8829)
	);

	bfr new_net_8830_bfr_after (
		.din(new_net_8829),
		.dout(new_net_8830)
	);

	bfr new_net_8831_bfr_after (
		.din(new_net_8830),
		.dout(new_net_8831)
	);

	bfr new_net_8832_bfr_after (
		.din(new_net_8831),
		.dout(new_net_8832)
	);

	bfr new_net_2381_bfr_after (
		.din(new_net_8832),
		.dout(new_net_2381)
	);

	bfr new_net_2465_bfr_after (
		.din(n_0517_),
		.dout(new_net_2465)
	);

	bfr new_net_8833_bfr_after (
		.din(n_0630_),
		.dout(new_net_8833)
	);

	bfr new_net_8834_bfr_after (
		.din(new_net_8833),
		.dout(new_net_8834)
	);

	bfr new_net_2486_bfr_after (
		.din(new_net_8834),
		.dout(new_net_2486)
	);

	bfr new_net_8835_bfr_after (
		.din(N169),
		.dout(new_net_8835)
	);

	bfr new_net_8836_bfr_after (
		.din(new_net_8835),
		.dout(new_net_8836)
	);

	bfr new_net_8837_bfr_after (
		.din(new_net_8836),
		.dout(new_net_8837)
	);

	bfr new_net_2318_bfr_after (
		.din(new_net_8837),
		.dout(new_net_2318)
	);

	bfr new_net_8838_bfr_after (
		.din(n_0205_),
		.dout(new_net_8838)
	);

	bfr new_net_8839_bfr_after (
		.din(new_net_8838),
		.dout(new_net_8839)
	);

	bfr new_net_8840_bfr_after (
		.din(new_net_8839),
		.dout(new_net_8840)
	);

	bfr new_net_8841_bfr_after (
		.din(new_net_8840),
		.dout(new_net_8841)
	);

	bfr new_net_2402_bfr_after (
		.din(new_net_8841),
		.dout(new_net_2402)
	);

	bfr new_net_8842_bfr_after (
		.din(N231),
		.dout(new_net_8842)
	);

	bfr new_net_8843_bfr_after (
		.din(new_net_8842),
		.dout(new_net_8843)
	);

	bfr new_net_8844_bfr_after (
		.din(new_net_8843),
		.dout(new_net_8844)
	);

	bfr new_net_2234_bfr_after (
		.din(new_net_8844),
		.dout(new_net_2234)
	);

	bfr new_net_8845_bfr_after (
		.din(N225),
		.dout(new_net_8845)
	);

	bfr new_net_8846_bfr_after (
		.din(new_net_8845),
		.dout(new_net_8846)
	);

	bfr new_net_8847_bfr_after (
		.din(new_net_8846),
		.dout(new_net_8847)
	);

	bfr new_net_2255_bfr_after (
		.din(new_net_8847),
		.dout(new_net_2255)
	);

	bfr new_net_8848_bfr_after (
		.din(N23),
		.dout(new_net_8848)
	);

	bfr new_net_8849_bfr_after (
		.din(new_net_8848),
		.dout(new_net_8849)
	);

	bfr new_net_8850_bfr_after (
		.din(new_net_8849),
		.dout(new_net_8850)
	);

	bfr new_net_2192_bfr_after (
		.din(new_net_8850),
		.dout(new_net_2192)
	);

	bfr new_net_8851_bfr_after (
		.din(N144),
		.dout(new_net_8851)
	);

	bfr new_net_8852_bfr_after (
		.din(new_net_8851),
		.dout(new_net_8852)
	);

	bfr new_net_8853_bfr_after (
		.din(new_net_8852),
		.dout(new_net_8853)
	);

	bfr new_net_2218_bfr_after (
		.din(new_net_8853),
		.dout(new_net_2218)
	);

	bfr new_net_8854_bfr_after (
		.din(N114),
		.dout(new_net_8854)
	);

	bfr new_net_8855_bfr_after (
		.din(new_net_8854),
		.dout(new_net_8855)
	);

	bfr new_net_8856_bfr_after (
		.din(new_net_8855),
		.dout(new_net_8856)
	);

	bfr new_net_2276_bfr_after (
		.din(new_net_8856),
		.dout(new_net_2276)
	);

	bfr new_net_8857_bfr_after (
		.din(N187),
		.dout(new_net_8857)
	);

	bfr new_net_8858_bfr_after (
		.din(new_net_8857),
		.dout(new_net_8858)
	);

	bfr new_net_8859_bfr_after (
		.din(new_net_8858),
		.dout(new_net_8859)
	);

	bfr new_net_2339_bfr_after (
		.din(new_net_8859),
		.dout(new_net_2339)
	);

	bfr new_net_8860_bfr_after (
		.din(n_0628_),
		.dout(new_net_8860)
	);

	bfr new_net_2488_bfr_after (
		.din(new_net_8860),
		.dout(new_net_2488)
	);

	bfr new_net_8861_bfr_after (
		.din(new_net_2574),
		.dout(new_net_8861)
	);

	bfr new_net_8862_bfr_after (
		.din(new_net_8861),
		.dout(new_net_8862)
	);

	bfr new_net_8863_bfr_after (
		.din(new_net_8862),
		.dout(new_net_8863)
	);

	bfr new_net_8864_bfr_after (
		.din(new_net_8863),
		.dout(new_net_8864)
	);

	bfr new_net_8865_bfr_after (
		.din(new_net_8864),
		.dout(new_net_8865)
	);

	bfr new_net_8866_bfr_after (
		.din(new_net_8865),
		.dout(new_net_8866)
	);

	bfr new_net_8867_bfr_after (
		.din(new_net_8866),
		.dout(new_net_8867)
	);

	bfr new_net_8868_bfr_after (
		.din(new_net_8867),
		.dout(new_net_8868)
	);

	bfr new_net_8869_bfr_after (
		.din(new_net_8868),
		.dout(new_net_8869)
	);

	bfr new_net_8870_bfr_after (
		.din(new_net_8869),
		.dout(new_net_8870)
	);

	bfr new_net_8871_bfr_after (
		.din(new_net_8870),
		.dout(new_net_8871)
	);

	bfr new_net_8872_bfr_after (
		.din(new_net_8871),
		.dout(new_net_8872)
	);

	bfr new_net_8873_bfr_after (
		.din(new_net_8872),
		.dout(new_net_8873)
	);

	bfr new_net_8874_bfr_after (
		.din(new_net_8873),
		.dout(new_net_8874)
	);

	bfr new_net_8875_bfr_after (
		.din(new_net_8874),
		.dout(new_net_8875)
	);

	bfr new_net_8876_bfr_after (
		.din(new_net_8875),
		.dout(new_net_8876)
	);

	bfr new_net_8877_bfr_after (
		.din(new_net_8876),
		.dout(new_net_8877)
	);

	bfr new_net_8878_bfr_after (
		.din(new_net_8877),
		.dout(new_net_8878)
	);

	bfr new_net_8879_bfr_after (
		.din(new_net_8878),
		.dout(new_net_8879)
	);

	bfr new_net_8880_bfr_after (
		.din(new_net_8879),
		.dout(new_net_8880)
	);

	bfr new_net_8881_bfr_after (
		.din(new_net_8880),
		.dout(new_net_8881)
	);

	bfr new_net_8882_bfr_after (
		.din(new_net_8881),
		.dout(new_net_8882)
	);

	bfr new_net_8883_bfr_after (
		.din(new_net_8882),
		.dout(new_net_8883)
	);

	bfr new_net_8884_bfr_after (
		.din(new_net_8883),
		.dout(new_net_8884)
	);

	bfr N10907_bfr_after (
		.din(new_net_8884),
		.dout(N10907)
	);

	bfr new_net_8885_bfr_after (
		.din(N201),
		.dout(new_net_8885)
	);

	bfr new_net_8886_bfr_after (
		.din(new_net_8885),
		.dout(new_net_8886)
	);

	bfr new_net_8887_bfr_after (
		.din(new_net_8886),
		.dout(new_net_8887)
	);

	bfr new_net_2369_bfr_after (
		.din(new_net_8887),
		.dout(new_net_2369)
	);

	bfr new_net_2432_bfr_after (
		.din(n_0295_),
		.dout(new_net_2432)
	);

	bfr new_net_8888_bfr_after (
		.din(n_0283_),
		.dout(new_net_8888)
	);

	bfr new_net_8889_bfr_after (
		.din(new_net_8888),
		.dout(new_net_8889)
	);

	bfr new_net_8890_bfr_after (
		.din(new_net_8889),
		.dout(new_net_8890)
	);

	bfr new_net_8891_bfr_after (
		.din(new_net_8890),
		.dout(new_net_8891)
	);

	bfr new_net_8892_bfr_after (
		.din(new_net_8891),
		.dout(new_net_8892)
	);

	bfr new_net_8893_bfr_after (
		.din(new_net_8892),
		.dout(new_net_8893)
	);

	bfr new_net_2427_bfr_after (
		.din(new_net_8893),
		.dout(new_net_2427)
	);

	bfr new_net_8894_bfr_after (
		.din(new_net_2507),
		.dout(new_net_8894)
	);

	bfr new_net_8895_bfr_after (
		.din(new_net_8894),
		.dout(new_net_8895)
	);

	bfr new_net_8896_bfr_after (
		.din(new_net_8895),
		.dout(new_net_8896)
	);

	bfr new_net_8897_bfr_after (
		.din(new_net_8896),
		.dout(new_net_8897)
	);

	bfr new_net_8898_bfr_after (
		.din(new_net_8897),
		.dout(new_net_8898)
	);

	bfr new_net_8899_bfr_after (
		.din(new_net_8898),
		.dout(new_net_8899)
	);

	bfr new_net_8900_bfr_after (
		.din(new_net_8899),
		.dout(new_net_8900)
	);

	bfr new_net_8901_bfr_after (
		.din(new_net_8900),
		.dout(new_net_8901)
	);

	bfr new_net_8902_bfr_after (
		.din(new_net_8901),
		.dout(new_net_8902)
	);

	bfr new_net_8903_bfr_after (
		.din(new_net_8902),
		.dout(new_net_8903)
	);

	bfr new_net_8904_bfr_after (
		.din(new_net_8903),
		.dout(new_net_8904)
	);

	bfr new_net_8905_bfr_after (
		.din(new_net_8904),
		.dout(new_net_8905)
	);

	bfr new_net_8906_bfr_after (
		.din(new_net_8905),
		.dout(new_net_8906)
	);

	bfr new_net_8907_bfr_after (
		.din(new_net_8906),
		.dout(new_net_8907)
	);

	bfr new_net_8908_bfr_after (
		.din(new_net_8907),
		.dout(new_net_8908)
	);

	bfr new_net_8909_bfr_after (
		.din(new_net_8908),
		.dout(new_net_8909)
	);

	bfr new_net_8910_bfr_after (
		.din(new_net_8909),
		.dout(new_net_8910)
	);

	bfr new_net_8911_bfr_after (
		.din(new_net_8910),
		.dout(new_net_8911)
	);

	bfr new_net_8912_bfr_after (
		.din(new_net_8911),
		.dout(new_net_8912)
	);

	bfr new_net_8913_bfr_after (
		.din(new_net_8912),
		.dout(new_net_8913)
	);

	bfr new_net_8914_bfr_after (
		.din(new_net_8913),
		.dout(new_net_8914)
	);

	bfr new_net_8915_bfr_after (
		.din(new_net_8914),
		.dout(new_net_8915)
	);

	bfr new_net_8916_bfr_after (
		.din(new_net_8915),
		.dout(new_net_8916)
	);

	bfr new_net_8917_bfr_after (
		.din(new_net_8916),
		.dout(new_net_8917)
	);

	bfr new_net_8918_bfr_after (
		.din(new_net_8917),
		.dout(new_net_8918)
	);

	bfr new_net_8919_bfr_after (
		.din(new_net_8918),
		.dout(new_net_8919)
	);

	bfr new_net_8920_bfr_after (
		.din(new_net_8919),
		.dout(new_net_8920)
	);

	bfr new_net_8921_bfr_after (
		.din(new_net_8920),
		.dout(new_net_8921)
	);

	bfr new_net_8922_bfr_after (
		.din(new_net_8921),
		.dout(new_net_8922)
	);

	bfr new_net_8923_bfr_after (
		.din(new_net_8922),
		.dout(new_net_8923)
	);

	bfr new_net_8924_bfr_after (
		.din(new_net_8923),
		.dout(new_net_8924)
	);

	bfr new_net_8925_bfr_after (
		.din(new_net_8924),
		.dout(new_net_8925)
	);

	bfr new_net_8926_bfr_after (
		.din(new_net_8925),
		.dout(new_net_8926)
	);

	bfr new_net_8927_bfr_after (
		.din(new_net_8926),
		.dout(new_net_8927)
	);

	bfr new_net_8928_bfr_after (
		.din(new_net_8927),
		.dout(new_net_8928)
	);

	bfr new_net_8929_bfr_after (
		.din(new_net_8928),
		.dout(new_net_8929)
	);

	bfr new_net_8930_bfr_after (
		.din(new_net_8929),
		.dout(new_net_8930)
	);

	bfr new_net_8931_bfr_after (
		.din(new_net_8930),
		.dout(new_net_8931)
	);

	bfr new_net_8932_bfr_after (
		.din(new_net_8931),
		.dout(new_net_8932)
	);

	bfr new_net_8933_bfr_after (
		.din(new_net_8932),
		.dout(new_net_8933)
	);

	bfr new_net_8934_bfr_after (
		.din(new_net_8933),
		.dout(new_net_8934)
	);

	bfr new_net_8935_bfr_after (
		.din(new_net_8934),
		.dout(new_net_8935)
	);

	bfr new_net_8936_bfr_after (
		.din(new_net_8935),
		.dout(new_net_8936)
	);

	bfr new_net_8937_bfr_after (
		.din(new_net_8936),
		.dout(new_net_8937)
	);

	bfr new_net_8938_bfr_after (
		.din(new_net_8937),
		.dout(new_net_8938)
	);

	bfr new_net_8939_bfr_after (
		.din(new_net_8938),
		.dout(new_net_8939)
	);

	bfr new_net_8940_bfr_after (
		.din(new_net_8939),
		.dout(new_net_8940)
	);

	bfr new_net_8941_bfr_after (
		.din(new_net_8940),
		.dout(new_net_8941)
	);

	bfr new_net_8942_bfr_after (
		.din(new_net_8941),
		.dout(new_net_8942)
	);

	bfr N10112_bfr_after (
		.din(new_net_8942),
		.dout(N10112)
	);

	bfr new_net_8943_bfr_after (
		.din(N63),
		.dout(new_net_8943)
	);

	bfr new_net_8944_bfr_after (
		.din(new_net_8943),
		.dout(new_net_8944)
	);

	bfr new_net_8945_bfr_after (
		.din(new_net_8944),
		.dout(new_net_8945)
	);

	bfr new_net_2312_bfr_after (
		.din(new_net_8945),
		.dout(new_net_2312)
	);

	bfr new_net_8946_bfr_after (
		.din(N110),
		.dout(new_net_8946)
	);

	bfr new_net_8947_bfr_after (
		.din(new_net_8946),
		.dout(new_net_8947)
	);

	bfr new_net_8948_bfr_after (
		.din(new_net_8947),
		.dout(new_net_8948)
	);

	bfr new_net_2308_bfr_after (
		.din(new_net_8948),
		.dout(new_net_2308)
	);

	bfr new_net_8949_bfr_after (
		.din(new_net_2497),
		.dout(new_net_8949)
	);

	bfr new_net_8950_bfr_after (
		.din(new_net_8949),
		.dout(new_net_8950)
	);

	bfr new_net_8951_bfr_after (
		.din(new_net_8950),
		.dout(new_net_8951)
	);

	bfr new_net_8952_bfr_after (
		.din(new_net_8951),
		.dout(new_net_8952)
	);

	bfr new_net_8953_bfr_after (
		.din(new_net_8952),
		.dout(new_net_8953)
	);

	bfr N10716_bfr_after (
		.din(new_net_8953),
		.dout(N10716)
	);

	bfr new_net_8954_bfr_after (
		.din(new_net_2509),
		.dout(new_net_8954)
	);

	bfr new_net_8955_bfr_after (
		.din(new_net_8954),
		.dout(new_net_8955)
	);

	bfr new_net_8956_bfr_after (
		.din(new_net_8955),
		.dout(new_net_8956)
	);

	bfr new_net_8957_bfr_after (
		.din(new_net_8956),
		.dout(new_net_8957)
	);

	bfr new_net_8958_bfr_after (
		.din(new_net_8957),
		.dout(new_net_8958)
	);

	bfr new_net_8959_bfr_after (
		.din(new_net_8958),
		.dout(new_net_8959)
	);

	bfr new_net_8960_bfr_after (
		.din(new_net_8959),
		.dout(new_net_8960)
	);

	bfr new_net_8961_bfr_after (
		.din(new_net_8960),
		.dout(new_net_8961)
	);

	bfr new_net_8962_bfr_after (
		.din(new_net_8961),
		.dout(new_net_8962)
	);

	bfr new_net_8963_bfr_after (
		.din(new_net_8962),
		.dout(new_net_8963)
	);

	bfr new_net_8964_bfr_after (
		.din(new_net_8963),
		.dout(new_net_8964)
	);

	bfr new_net_8965_bfr_after (
		.din(new_net_8964),
		.dout(new_net_8965)
	);

	bfr new_net_8966_bfr_after (
		.din(new_net_8965),
		.dout(new_net_8966)
	);

	bfr new_net_8967_bfr_after (
		.din(new_net_8966),
		.dout(new_net_8967)
	);

	bfr new_net_8968_bfr_after (
		.din(new_net_8967),
		.dout(new_net_8968)
	);

	bfr new_net_8969_bfr_after (
		.din(new_net_8968),
		.dout(new_net_8969)
	);

	bfr new_net_8970_bfr_after (
		.din(new_net_8969),
		.dout(new_net_8970)
	);

	bfr new_net_8971_bfr_after (
		.din(new_net_8970),
		.dout(new_net_8971)
	);

	bfr new_net_8972_bfr_after (
		.din(new_net_8971),
		.dout(new_net_8972)
	);

	bfr new_net_8973_bfr_after (
		.din(new_net_8972),
		.dout(new_net_8973)
	);

	bfr new_net_8974_bfr_after (
		.din(new_net_8973),
		.dout(new_net_8974)
	);

	bfr new_net_8975_bfr_after (
		.din(new_net_8974),
		.dout(new_net_8975)
	);

	bfr new_net_8976_bfr_after (
		.din(new_net_8975),
		.dout(new_net_8976)
	);

	bfr new_net_8977_bfr_after (
		.din(new_net_8976),
		.dout(new_net_8977)
	);

	bfr N10905_bfr_after (
		.din(new_net_8977),
		.dout(N10905)
	);

	bfr new_net_8978_bfr_after (
		.din(new_net_2521),
		.dout(new_net_8978)
	);

	bfr new_net_8979_bfr_after (
		.din(new_net_8978),
		.dout(new_net_8979)
	);

	bfr new_net_8980_bfr_after (
		.din(new_net_8979),
		.dout(new_net_8980)
	);

	bfr new_net_8981_bfr_after (
		.din(new_net_8980),
		.dout(new_net_8981)
	);

	bfr new_net_8982_bfr_after (
		.din(new_net_8981),
		.dout(new_net_8982)
	);

	bfr new_net_8983_bfr_after (
		.din(new_net_8982),
		.dout(new_net_8983)
	);

	bfr new_net_8984_bfr_after (
		.din(new_net_8983),
		.dout(new_net_8984)
	);

	bfr new_net_8985_bfr_after (
		.din(new_net_8984),
		.dout(new_net_8985)
	);

	bfr new_net_8986_bfr_after (
		.din(new_net_8985),
		.dout(new_net_8986)
	);

	bfr new_net_8987_bfr_after (
		.din(new_net_8986),
		.dout(new_net_8987)
	);

	bfr new_net_8988_bfr_after (
		.din(new_net_8987),
		.dout(new_net_8988)
	);

	bfr new_net_8989_bfr_after (
		.din(new_net_8988),
		.dout(new_net_8989)
	);

	bfr new_net_8990_bfr_after (
		.din(new_net_8989),
		.dout(new_net_8990)
	);

	bfr N10761_bfr_after (
		.din(new_net_8990),
		.dout(N10761)
	);

	bfr new_net_8991_bfr_after (
		.din(new_net_2533),
		.dout(new_net_8991)
	);

	bfr new_net_8992_bfr_after (
		.din(new_net_8991),
		.dout(new_net_8992)
	);

	bfr new_net_8993_bfr_after (
		.din(new_net_8992),
		.dout(new_net_8993)
	);

	bfr new_net_8994_bfr_after (
		.din(new_net_8993),
		.dout(new_net_8994)
	);

	bfr new_net_8995_bfr_after (
		.din(new_net_8994),
		.dout(new_net_8995)
	);

	bfr new_net_8996_bfr_after (
		.din(new_net_8995),
		.dout(new_net_8996)
	);

	bfr new_net_8997_bfr_after (
		.din(new_net_8996),
		.dout(new_net_8997)
	);

	bfr new_net_8998_bfr_after (
		.din(new_net_8997),
		.dout(new_net_8998)
	);

	bfr new_net_8999_bfr_after (
		.din(new_net_8998),
		.dout(new_net_8999)
	);

	bfr new_net_9000_bfr_after (
		.din(new_net_8999),
		.dout(new_net_9000)
	);

	bfr new_net_9001_bfr_after (
		.din(new_net_9000),
		.dout(new_net_9001)
	);

	bfr new_net_9002_bfr_after (
		.din(new_net_9001),
		.dout(new_net_9002)
	);

	bfr new_net_9003_bfr_after (
		.din(new_net_9002),
		.dout(new_net_9003)
	);

	bfr new_net_9004_bfr_after (
		.din(new_net_9003),
		.dout(new_net_9004)
	);

	bfr new_net_9005_bfr_after (
		.din(new_net_9004),
		.dout(new_net_9005)
	);

	bfr new_net_9006_bfr_after (
		.din(new_net_9005),
		.dout(new_net_9006)
	);

	bfr new_net_9007_bfr_after (
		.din(new_net_9006),
		.dout(new_net_9007)
	);

	bfr new_net_9008_bfr_after (
		.din(new_net_9007),
		.dout(new_net_9008)
	);

	bfr new_net_9009_bfr_after (
		.din(new_net_9008),
		.dout(new_net_9009)
	);

	bfr new_net_9010_bfr_after (
		.din(new_net_9009),
		.dout(new_net_9010)
	);

	bfr new_net_9011_bfr_after (
		.din(new_net_9010),
		.dout(new_net_9011)
	);

	bfr new_net_9012_bfr_after (
		.din(new_net_9011),
		.dout(new_net_9012)
	);

	bfr new_net_9013_bfr_after (
		.din(new_net_9012),
		.dout(new_net_9013)
	);

	bfr new_net_9014_bfr_after (
		.din(new_net_9013),
		.dout(new_net_9014)
	);

	bfr new_net_9015_bfr_after (
		.din(new_net_9014),
		.dout(new_net_9015)
	);

	bfr new_net_9016_bfr_after (
		.din(new_net_9015),
		.dout(new_net_9016)
	);

	bfr new_net_9017_bfr_after (
		.din(new_net_9016),
		.dout(new_net_9017)
	);

	bfr new_net_9018_bfr_after (
		.din(new_net_9017),
		.dout(new_net_9018)
	);

	bfr new_net_9019_bfr_after (
		.din(new_net_9018),
		.dout(new_net_9019)
	);

	bfr new_net_9020_bfr_after (
		.din(new_net_9019),
		.dout(new_net_9020)
	);

	bfr new_net_9021_bfr_after (
		.din(new_net_9020),
		.dout(new_net_9021)
	);

	bfr new_net_9022_bfr_after (
		.din(new_net_9021),
		.dout(new_net_9022)
	);

	bfr new_net_9023_bfr_after (
		.din(new_net_9022),
		.dout(new_net_9023)
	);

	bfr new_net_9024_bfr_after (
		.din(new_net_9023),
		.dout(new_net_9024)
	);

	bfr N10628_bfr_after (
		.din(new_net_9024),
		.dout(N10628)
	);

	bfr new_net_9025_bfr_after (
		.din(new_net_2545),
		.dout(new_net_9025)
	);

	bfr new_net_9026_bfr_after (
		.din(new_net_9025),
		.dout(new_net_9026)
	);

	bfr new_net_9027_bfr_after (
		.din(new_net_9026),
		.dout(new_net_9027)
	);

	bfr new_net_9028_bfr_after (
		.din(new_net_9027),
		.dout(new_net_9028)
	);

	bfr new_net_9029_bfr_after (
		.din(new_net_9028),
		.dout(new_net_9029)
	);

	bfr new_net_9030_bfr_after (
		.din(new_net_9029),
		.dout(new_net_9030)
	);

	bfr new_net_9031_bfr_after (
		.din(new_net_9030),
		.dout(new_net_9031)
	);

	bfr new_net_9032_bfr_after (
		.din(new_net_9031),
		.dout(new_net_9032)
	);

	bfr N10641_bfr_after (
		.din(new_net_9032),
		.dout(N10641)
	);

	bfr new_net_9033_bfr_after (
		.din(n_0497_),
		.dout(new_net_9033)
	);

	bfr new_net_9034_bfr_after (
		.din(new_net_9033),
		.dout(new_net_9034)
	);

	bfr new_net_9035_bfr_after (
		.din(new_net_9034),
		.dout(new_net_9035)
	);

	bfr new_net_9036_bfr_after (
		.din(new_net_9035),
		.dout(new_net_9036)
	);

	bfr new_net_9037_bfr_after (
		.din(new_net_9036),
		.dout(new_net_9037)
	);

	bfr new_net_9038_bfr_after (
		.din(new_net_9037),
		.dout(new_net_9038)
	);

	bfr new_net_9039_bfr_after (
		.din(new_net_9038),
		.dout(new_net_9039)
	);

	bfr new_net_9040_bfr_after (
		.din(new_net_9039),
		.dout(new_net_9040)
	);

	bfr new_net_9041_bfr_after (
		.din(new_net_9040),
		.dout(new_net_9041)
	);

	bfr new_net_9042_bfr_after (
		.din(new_net_9041),
		.dout(new_net_9042)
	);

	bfr new_net_9043_bfr_after (
		.din(new_net_9042),
		.dout(new_net_9043)
	);

	bfr new_net_9044_bfr_after (
		.din(new_net_9043),
		.dout(new_net_9044)
	);

	bfr new_net_9045_bfr_after (
		.din(new_net_9044),
		.dout(new_net_9045)
	);

	bfr new_net_9046_bfr_after (
		.din(new_net_9045),
		.dout(new_net_9046)
	);

	bfr new_net_9047_bfr_after (
		.din(new_net_9046),
		.dout(new_net_9047)
	);

	bfr new_net_9048_bfr_after (
		.din(new_net_9047),
		.dout(new_net_9048)
	);

	bfr new_net_9049_bfr_after (
		.din(new_net_9048),
		.dout(new_net_9049)
	);

	bfr new_net_9050_bfr_after (
		.din(new_net_9049),
		.dout(new_net_9050)
	);

	bfr new_net_9051_bfr_after (
		.din(new_net_9050),
		.dout(new_net_9051)
	);

	bfr new_net_9052_bfr_after (
		.din(new_net_9051),
		.dout(new_net_9052)
	);

	bfr new_net_9053_bfr_after (
		.din(new_net_9052),
		.dout(new_net_9053)
	);

	bfr new_net_9054_bfr_after (
		.din(new_net_9053),
		.dout(new_net_9054)
	);

	bfr new_net_9055_bfr_after (
		.din(new_net_9054),
		.dout(new_net_9055)
	);

	bfr new_net_9056_bfr_after (
		.din(new_net_9055),
		.dout(new_net_9056)
	);

	bfr new_net_9057_bfr_after (
		.din(new_net_9056),
		.dout(new_net_9057)
	);

	bfr new_net_2462_bfr_after (
		.din(new_net_9057),
		.dout(new_net_2462)
	);

	bfr new_net_2457_bfr_after (
		.din(n_0450_),
		.dout(new_net_2457)
	);

	bfr new_net_9058_bfr_after (
		.din(n_0182_),
		.dout(new_net_9058)
	);

	bfr new_net_9059_bfr_after (
		.din(new_net_9058),
		.dout(new_net_9059)
	);

	bfr new_net_9060_bfr_after (
		.din(new_net_9059),
		.dout(new_net_9060)
	);

	bfr new_net_2400_bfr_after (
		.din(new_net_9060),
		.dout(new_net_2400)
	);

	bfr new_net_9061_bfr_after (
		.din(N179),
		.dout(new_net_9061)
	);

	bfr new_net_9062_bfr_after (
		.din(new_net_9061),
		.dout(new_net_9062)
	);

	bfr new_net_9063_bfr_after (
		.din(new_net_9062),
		.dout(new_net_9063)
	);

	bfr new_net_2355_bfr_after (
		.din(new_net_9063),
		.dout(new_net_2355)
	);

	bfr new_net_9064_bfr_after (
		.din(N147),
		.dout(new_net_9064)
	);

	bfr new_net_9065_bfr_after (
		.din(new_net_9064),
		.dout(new_net_9065)
	);

	bfr new_net_9066_bfr_after (
		.din(new_net_9065),
		.dout(new_net_9066)
	);

	bfr new_net_2208_bfr_after (
		.din(new_net_9066),
		.dout(new_net_2208)
	);

	bfr new_net_9067_bfr_after (
		.din(N73),
		.dout(new_net_9067)
	);

	bfr new_net_9068_bfr_after (
		.din(new_net_9067),
		.dout(new_net_9068)
	);

	bfr new_net_9069_bfr_after (
		.din(new_net_9068),
		.dout(new_net_9069)
	);

	bfr new_net_2292_bfr_after (
		.din(new_net_9069),
		.dout(new_net_2292)
	);

	bfr new_net_2376_bfr_after (
		.din(n_1281_),
		.dout(new_net_2376)
	);

	bfr new_net_2460_bfr_after (
		.din(n_0478_),
		.dout(new_net_2460)
	);

	bfr new_net_2481_bfr_after (
		.din(n_0609_),
		.dout(new_net_2481)
	);

	bfr new_net_9070_bfr_after (
		.din(N86),
		.dout(new_net_9070)
	);

	bfr new_net_9071_bfr_after (
		.din(new_net_9070),
		.dout(new_net_9071)
	);

	bfr new_net_9072_bfr_after (
		.din(new_net_9071),
		.dout(new_net_9072)
	);

	bfr new_net_2313_bfr_after (
		.din(new_net_9072),
		.dout(new_net_2313)
	);

	bfr new_net_2397_bfr_after (
		.din(n_0187_),
		.dout(new_net_2397)
	);

	bfr new_net_9073_bfr_after (
		.din(N35),
		.dout(new_net_9073)
	);

	bfr new_net_9074_bfr_after (
		.din(new_net_9073),
		.dout(new_net_9074)
	);

	bfr new_net_9075_bfr_after (
		.din(new_net_9074),
		.dout(new_net_9075)
	);

	bfr new_net_2271_bfr_after (
		.din(new_net_9075),
		.dout(new_net_2271)
	);

	bfr new_net_2334_bfr_after (
		.din(n_1177_),
		.dout(new_net_2334)
	);

	bfr N10759_bfr_after (
		.din(new_net_2519),
		.dout(N10759)
	);

	bfr new_net_9076_bfr_after (
		.din(N156),
		.dout(new_net_9076)
	);

	bfr new_net_9077_bfr_after (
		.din(new_net_9076),
		.dout(new_net_9077)
	);

	bfr new_net_9078_bfr_after (
		.din(new_net_9077),
		.dout(new_net_9078)
	);

	bfr new_net_2203_bfr_after (
		.din(new_net_9078),
		.dout(new_net_2203)
	);

	bfr new_net_9079_bfr_after (
		.din(N216),
		.dout(new_net_9079)
	);

	bfr new_net_9080_bfr_after (
		.din(new_net_9079),
		.dout(new_net_9080)
	);

	bfr new_net_9081_bfr_after (
		.din(new_net_9080),
		.dout(new_net_9081)
	);

	bfr new_net_2224_bfr_after (
		.din(new_net_9081),
		.dout(new_net_2224)
	);

	bfr new_net_2245_bfr_after (
		.din(n_0831_),
		.dout(new_net_2245)
	);

	bfr new_net_2266_bfr_after (
		.din(n_0876_),
		.dout(new_net_2266)
	);

	bfr new_net_9082_bfr_after (
		.din(N74),
		.dout(new_net_9082)
	);

	bfr new_net_9083_bfr_after (
		.din(new_net_9082),
		.dout(new_net_9083)
	);

	bfr new_net_9084_bfr_after (
		.din(new_net_9083),
		.dout(new_net_9084)
	);

	bfr new_net_2287_bfr_after (
		.din(new_net_9084),
		.dout(new_net_2287)
	);

	bfr new_net_9085_bfr_after (
		.din(N192),
		.dout(new_net_9085)
	);

	bfr new_net_9086_bfr_after (
		.din(new_net_9085),
		.dout(new_net_9086)
	);

	bfr new_net_9087_bfr_after (
		.din(new_net_9086),
		.dout(new_net_9087)
	);

	bfr new_net_2329_bfr_after (
		.din(new_net_9087),
		.dout(new_net_2329)
	);

	bfr new_net_9088_bfr_after (
		.din(N178),
		.dout(new_net_9088)
	);

	bfr new_net_9089_bfr_after (
		.din(new_net_9088),
		.dout(new_net_9089)
	);

	bfr new_net_9090_bfr_after (
		.din(new_net_9089),
		.dout(new_net_9090)
	);

	bfr new_net_2350_bfr_after (
		.din(new_net_9090),
		.dout(new_net_2350)
	);

	bfr new_net_9091_bfr_after (
		.din(N200),
		.dout(new_net_9091)
	);

	bfr new_net_9092_bfr_after (
		.din(new_net_9091),
		.dout(new_net_9092)
	);

	bfr new_net_9093_bfr_after (
		.din(new_net_9092),
		.dout(new_net_9093)
	);

	bfr new_net_2371_bfr_after (
		.din(new_net_9093),
		.dout(new_net_2371)
	);

	bfr new_net_2434_bfr_after (
		.din(n_0305_),
		.dout(new_net_2434)
	);

	bfr new_net_2455_bfr_after (
		.din(n_0435_),
		.dout(new_net_2455)
	);

	bfr new_net_9094_bfr_after (
		.din(new_net_2539),
		.dout(new_net_9094)
	);

	bfr new_net_9095_bfr_after (
		.din(new_net_9094),
		.dout(new_net_9095)
	);

	bfr new_net_9096_bfr_after (
		.din(new_net_9095),
		.dout(new_net_9096)
	);

	bfr new_net_9097_bfr_after (
		.din(new_net_9096),
		.dout(new_net_9097)
	);

	bfr new_net_9098_bfr_after (
		.din(new_net_9097),
		.dout(new_net_9098)
	);

	bfr new_net_9099_bfr_after (
		.din(new_net_9098),
		.dout(new_net_9099)
	);

	bfr new_net_9100_bfr_after (
		.din(new_net_9099),
		.dout(new_net_9100)
	);

	bfr new_net_9101_bfr_after (
		.din(new_net_9100),
		.dout(new_net_9101)
	);

	bfr new_net_9102_bfr_after (
		.din(new_net_9101),
		.dout(new_net_9102)
	);

	bfr new_net_9103_bfr_after (
		.din(new_net_9102),
		.dout(new_net_9103)
	);

	bfr new_net_9104_bfr_after (
		.din(new_net_9103),
		.dout(new_net_9104)
	);

	bfr new_net_9105_bfr_after (
		.din(new_net_9104),
		.dout(new_net_9105)
	);

	bfr new_net_9106_bfr_after (
		.din(new_net_9105),
		.dout(new_net_9106)
	);

	bfr new_net_9107_bfr_after (
		.din(new_net_9106),
		.dout(new_net_9107)
	);

	bfr new_net_9108_bfr_after (
		.din(new_net_9107),
		.dout(new_net_9108)
	);

	bfr new_net_9109_bfr_after (
		.din(new_net_9108),
		.dout(new_net_9109)
	);

	bfr new_net_9110_bfr_after (
		.din(new_net_9109),
		.dout(new_net_9110)
	);

	bfr new_net_9111_bfr_after (
		.din(new_net_9110),
		.dout(new_net_9111)
	);

	bfr new_net_9112_bfr_after (
		.din(new_net_9111),
		.dout(new_net_9112)
	);

	bfr new_net_9113_bfr_after (
		.din(new_net_9112),
		.dout(new_net_9113)
	);

	bfr new_net_9114_bfr_after (
		.din(new_net_9113),
		.dout(new_net_9114)
	);

	bfr new_net_9115_bfr_after (
		.din(new_net_9114),
		.dout(new_net_9115)
	);

	bfr new_net_9116_bfr_after (
		.din(new_net_9115),
		.dout(new_net_9116)
	);

	bfr new_net_9117_bfr_after (
		.din(new_net_9116),
		.dout(new_net_9117)
	);

	bfr N11340_bfr_after (
		.din(new_net_9117),
		.dout(N11340)
	);

	bfr new_net_9118_bfr_after (
		.din(N217),
		.dout(new_net_9118)
	);

	bfr new_net_9119_bfr_after (
		.din(new_net_9118),
		.dout(new_net_9119)
	);

	bfr new_net_9120_bfr_after (
		.din(new_net_9119),
		.dout(new_net_9120)
	);

	bfr new_net_2261_bfr_after (
		.din(new_net_9120),
		.dout(new_net_2261)
	);

	bfr new_net_9121_bfr_after (
		.din(N58),
		.dout(new_net_9121)
	);

	bfr new_net_9122_bfr_after (
		.din(new_net_9121),
		.dout(new_net_9122)
	);

	bfr new_net_9123_bfr_after (
		.din(new_net_9122),
		.dout(new_net_9123)
	);

	bfr new_net_2303_bfr_after (
		.din(new_net_9123),
		.dout(new_net_2303)
	);

	bfr new_net_2387_bfr_after (
		.din(n_0077_),
		.dout(new_net_2387)
	);

	bfr new_net_9124_bfr_after (
		.din(n_0224_),
		.dout(new_net_9124)
	);

	bfr new_net_2408_bfr_after (
		.din(new_net_9124),
		.dout(new_net_2408)
	);

	bfr new_net_9125_bfr_after (
		.din(n_0936_),
		.dout(new_net_9125)
	);

	bfr new_net_9126_bfr_after (
		.din(new_net_9125),
		.dout(new_net_9126)
	);

	bfr new_net_2282_bfr_after (
		.din(new_net_9126),
		.dout(new_net_2282)
	);

	bfr new_net_2324_bfr_after (
		.din(n_1152_),
		.dout(new_net_2324)
	);

	bfr new_net_2345_bfr_after (
		.din(n_1200_),
		.dout(new_net_2345)
	);

	bfr new_net_9127_bfr_after (
		.din(N159),
		.dout(new_net_9127)
	);

	bfr new_net_9128_bfr_after (
		.din(new_net_9127),
		.dout(new_net_9128)
	);

	bfr new_net_9129_bfr_after (
		.din(new_net_9128),
		.dout(new_net_9129)
	);

	bfr new_net_2219_bfr_after (
		.din(new_net_9129),
		.dout(new_net_2219)
	);

	bfr new_net_9130_bfr_after (
		.din(N233),
		.dout(new_net_9130)
	);

	bfr new_net_9131_bfr_after (
		.din(new_net_9130),
		.dout(new_net_9131)
	);

	bfr new_net_9132_bfr_after (
		.din(new_net_9131),
		.dout(new_net_9132)
	);

	bfr new_net_2240_bfr_after (
		.din(new_net_9132),
		.dout(new_net_2240)
	);

	bfr new_net_9133_bfr_after (
		.din(N29),
		.dout(new_net_9133)
	);

	bfr new_net_9134_bfr_after (
		.din(new_net_9133),
		.dout(new_net_9134)
	);

	bfr new_net_9135_bfr_after (
		.din(new_net_9134),
		.dout(new_net_9135)
	);

	bfr new_net_2198_bfr_after (
		.din(new_net_9135),
		.dout(new_net_2198)
	);

	bfr new_net_9136_bfr_after (
		.din(N158),
		.dout(new_net_9136)
	);

	bfr new_net_9137_bfr_after (
		.din(new_net_9136),
		.dout(new_net_9137)
	);

	bfr new_net_9138_bfr_after (
		.din(new_net_9137),
		.dout(new_net_9138)
	);

	bfr new_net_2212_bfr_after (
		.din(new_net_9138),
		.dout(new_net_2212)
	);

	bfr new_net_9139_bfr_after (
		.din(N62),
		.dout(new_net_9139)
	);

	bfr new_net_9140_bfr_after (
		.din(new_net_9139),
		.dout(new_net_9140)
	);

	bfr new_net_9141_bfr_after (
		.din(new_net_9140),
		.dout(new_net_9141)
	);

	bfr new_net_2298_bfr_after (
		.din(new_net_9141),
		.dout(new_net_2298)
	);

	bfr new_net_9142_bfr_after (
		.din(n_0014_),
		.dout(new_net_9142)
	);

	bfr new_net_9143_bfr_after (
		.din(new_net_9142),
		.dout(new_net_9143)
	);

	bfr new_net_9144_bfr_after (
		.din(new_net_9143),
		.dout(new_net_9144)
	);

	bfr new_net_9145_bfr_after (
		.din(new_net_9144),
		.dout(new_net_9145)
	);

	bfr new_net_9146_bfr_after (
		.din(new_net_9145),
		.dout(new_net_9146)
	);

	bfr new_net_9147_bfr_after (
		.din(new_net_9146),
		.dout(new_net_9147)
	);

	bfr new_net_9148_bfr_after (
		.din(new_net_9147),
		.dout(new_net_9148)
	);

	bfr new_net_9149_bfr_after (
		.din(new_net_9148),
		.dout(new_net_9149)
	);

	bfr new_net_9150_bfr_after (
		.din(new_net_9149),
		.dout(new_net_9150)
	);

	bfr new_net_2382_bfr_after (
		.din(new_net_9150),
		.dout(new_net_2382)
	);

	bfr new_net_9151_bfr_after (
		.din(n_0529_),
		.dout(new_net_9151)
	);

	bfr new_net_9152_bfr_after (
		.din(new_net_9151),
		.dout(new_net_9152)
	);

	bfr new_net_9153_bfr_after (
		.din(new_net_9152),
		.dout(new_net_9153)
	);

	bfr new_net_9154_bfr_after (
		.din(new_net_9153),
		.dout(new_net_9154)
	);

	bfr new_net_9155_bfr_after (
		.din(new_net_9154),
		.dout(new_net_9155)
	);

	bfr new_net_9156_bfr_after (
		.din(new_net_9155),
		.dout(new_net_9156)
	);

	bfr new_net_9157_bfr_after (
		.din(new_net_9156),
		.dout(new_net_9157)
	);

	bfr new_net_9158_bfr_after (
		.din(new_net_9157),
		.dout(new_net_9158)
	);

	bfr new_net_9159_bfr_after (
		.din(new_net_9158),
		.dout(new_net_9159)
	);

	bfr new_net_9160_bfr_after (
		.din(new_net_9159),
		.dout(new_net_9160)
	);

	bfr new_net_9161_bfr_after (
		.din(new_net_9160),
		.dout(new_net_9161)
	);

	bfr new_net_9162_bfr_after (
		.din(new_net_9161),
		.dout(new_net_9162)
	);

	bfr new_net_9163_bfr_after (
		.din(new_net_9162),
		.dout(new_net_9163)
	);

	bfr new_net_9164_bfr_after (
		.din(new_net_9163),
		.dout(new_net_9164)
	);

	bfr new_net_2466_bfr_after (
		.din(new_net_9164),
		.dout(new_net_2466)
	);

	bfr new_net_2487_bfr_after (
		.din(n_0640_),
		.dout(new_net_2487)
	);

	bfr new_net_9165_bfr_after (
		.din(N168),
		.dout(new_net_9165)
	);

	bfr new_net_9166_bfr_after (
		.din(new_net_9165),
		.dout(new_net_9166)
	);

	bfr new_net_9167_bfr_after (
		.din(new_net_9166),
		.dout(new_net_9167)
	);

	bfr new_net_2319_bfr_after (
		.din(new_net_9167),
		.dout(new_net_2319)
	);

	bfr new_net_2403_bfr_after (
		.din(n_0212_),
		.dout(new_net_2403)
	);

	bfr new_net_9168_bfr_after (
		.din(N157),
		.dout(new_net_9168)
	);

	bfr new_net_9169_bfr_after (
		.din(new_net_9168),
		.dout(new_net_9169)
	);

	bfr new_net_9170_bfr_after (
		.din(new_net_9169),
		.dout(new_net_9170)
	);

	bfr new_net_2214_bfr_after (
		.din(new_net_9170),
		.dout(new_net_2214)
	);

	bfr new_net_9171_bfr_after (
		.din(N100),
		.dout(new_net_9171)
	);

	bfr new_net_9172_bfr_after (
		.din(new_net_9171),
		.dout(new_net_9172)
	);

	bfr new_net_9173_bfr_after (
		.din(new_net_9172),
		.dout(new_net_9173)
	);

	bfr new_net_2235_bfr_after (
		.din(new_net_9173),
		.dout(new_net_2235)
	);

	bfr new_net_9174_bfr_after (
		.din(N94),
		.dout(new_net_9174)
	);

	bfr new_net_9175_bfr_after (
		.din(new_net_9174),
		.dout(new_net_9175)
	);

	bfr new_net_9176_bfr_after (
		.din(new_net_9175),
		.dout(new_net_9176)
	);

	bfr new_net_2256_bfr_after (
		.din(new_net_9176),
		.dout(new_net_2256)
	);

	bfr new_net_2193_bfr_after (
		.din(n_0677_),
		.dout(new_net_2193)
	);

	bfr new_net_2366_bfr_after (
		.din(n_1259_),
		.dout(new_net_2366)
	);

	bfr new_net_9177_bfr_after (
		.din(n_0288_),
		.dout(new_net_9177)
	);

	bfr new_net_2429_bfr_after (
		.din(new_net_9177),
		.dout(new_net_2429)
	);

	bfr new_net_2424_bfr_after (
		.din(n_0278_),
		.dout(new_net_2424)
	);

	bfr N10706_bfr_after (
		.din(new_net_2552),
		.dout(N10706)
	);

	bfr new_net_9178_bfr_after (
		.din(new_net_2564),
		.dout(new_net_9178)
	);

	bfr new_net_9179_bfr_after (
		.din(new_net_9178),
		.dout(new_net_9179)
	);

	bfr new_net_9180_bfr_after (
		.din(new_net_9179),
		.dout(new_net_9180)
	);

	bfr new_net_9181_bfr_after (
		.din(new_net_9180),
		.dout(new_net_9181)
	);

	bfr new_net_9182_bfr_after (
		.din(new_net_9181),
		.dout(new_net_9182)
	);

	bfr new_net_9183_bfr_after (
		.din(new_net_9182),
		.dout(new_net_9183)
	);

	bfr new_net_9184_bfr_after (
		.din(new_net_9183),
		.dout(new_net_9184)
	);

	bfr new_net_9185_bfr_after (
		.din(new_net_9184),
		.dout(new_net_9185)
	);

	bfr new_net_9186_bfr_after (
		.din(new_net_9185),
		.dout(new_net_9186)
	);

	bfr new_net_9187_bfr_after (
		.din(new_net_9186),
		.dout(new_net_9187)
	);

	bfr new_net_9188_bfr_after (
		.din(new_net_9187),
		.dout(new_net_9188)
	);

	bfr new_net_9189_bfr_after (
		.din(new_net_9188),
		.dout(new_net_9189)
	);

	bfr new_net_9190_bfr_after (
		.din(new_net_9189),
		.dout(new_net_9190)
	);

	bfr new_net_9191_bfr_after (
		.din(new_net_9190),
		.dout(new_net_9191)
	);

	bfr new_net_9192_bfr_after (
		.din(new_net_9191),
		.dout(new_net_9192)
	);

	bfr new_net_9193_bfr_after (
		.din(new_net_9192),
		.dout(new_net_9193)
	);

	bfr new_net_9194_bfr_after (
		.din(new_net_9193),
		.dout(new_net_9194)
	);

	bfr N10713_bfr_after (
		.din(new_net_9194),
		.dout(N10713)
	);

	bfr new_net_2362_bfr_after (
		.din(n_1252_),
		.dout(new_net_2362)
	);

	bfr new_net_9195_bfr_after (
		.din(new_net_2499),
		.dout(new_net_9195)
	);

	bfr new_net_9196_bfr_after (
		.din(new_net_9195),
		.dout(new_net_9196)
	);

	bfr new_net_9197_bfr_after (
		.din(new_net_9196),
		.dout(new_net_9197)
	);

	bfr new_net_9198_bfr_after (
		.din(new_net_9197),
		.dout(new_net_9198)
	);

	bfr new_net_9199_bfr_after (
		.din(new_net_9198),
		.dout(new_net_9199)
	);

	bfr new_net_9200_bfr_after (
		.din(new_net_9199),
		.dout(new_net_9200)
	);

	bfr new_net_9201_bfr_after (
		.din(new_net_9200),
		.dout(new_net_9201)
	);

	bfr new_net_9202_bfr_after (
		.din(new_net_9201),
		.dout(new_net_9202)
	);

	bfr new_net_9203_bfr_after (
		.din(new_net_9202),
		.dout(new_net_9203)
	);

	bfr new_net_9204_bfr_after (
		.din(new_net_9203),
		.dout(new_net_9204)
	);

	bfr new_net_9205_bfr_after (
		.din(new_net_9204),
		.dout(new_net_9205)
	);

	bfr new_net_9206_bfr_after (
		.din(new_net_9205),
		.dout(new_net_9206)
	);

	bfr new_net_9207_bfr_after (
		.din(new_net_9206),
		.dout(new_net_9207)
	);

	bfr new_net_9208_bfr_after (
		.din(new_net_9207),
		.dout(new_net_9208)
	);

	bfr new_net_9209_bfr_after (
		.din(new_net_9208),
		.dout(new_net_9209)
	);

	bfr new_net_9210_bfr_after (
		.din(new_net_9209),
		.dout(new_net_9210)
	);

	bfr new_net_9211_bfr_after (
		.din(new_net_9210),
		.dout(new_net_9211)
	);

	bfr new_net_9212_bfr_after (
		.din(new_net_9211),
		.dout(new_net_9212)
	);

	bfr new_net_9213_bfr_after (
		.din(new_net_9212),
		.dout(new_net_9213)
	);

	bfr new_net_9214_bfr_after (
		.din(new_net_9213),
		.dout(new_net_9214)
	);

	bfr new_net_9215_bfr_after (
		.din(new_net_9214),
		.dout(new_net_9215)
	);

	bfr new_net_9216_bfr_after (
		.din(new_net_9215),
		.dout(new_net_9216)
	);

	bfr new_net_9217_bfr_after (
		.din(new_net_9216),
		.dout(new_net_9217)
	);

	bfr new_net_9218_bfr_after (
		.din(new_net_9217),
		.dout(new_net_9218)
	);

	bfr new_net_9219_bfr_after (
		.din(new_net_9218),
		.dout(new_net_9219)
	);

	bfr new_net_9220_bfr_after (
		.din(new_net_9219),
		.dout(new_net_9220)
	);

	bfr new_net_9221_bfr_after (
		.din(new_net_9220),
		.dout(new_net_9221)
	);

	bfr new_net_9222_bfr_after (
		.din(new_net_9221),
		.dout(new_net_9222)
	);

	bfr new_net_9223_bfr_after (
		.din(new_net_9222),
		.dout(new_net_9223)
	);

	bfr new_net_9224_bfr_after (
		.din(new_net_9223),
		.dout(new_net_9224)
	);

	bfr new_net_9225_bfr_after (
		.din(new_net_9224),
		.dout(new_net_9225)
	);

	bfr new_net_9226_bfr_after (
		.din(new_net_9225),
		.dout(new_net_9226)
	);

	bfr new_net_9227_bfr_after (
		.din(new_net_9226),
		.dout(new_net_9227)
	);

	bfr new_net_9228_bfr_after (
		.din(new_net_9227),
		.dout(new_net_9228)
	);

	bfr new_net_9229_bfr_after (
		.din(new_net_9228),
		.dout(new_net_9229)
	);

	bfr new_net_9230_bfr_after (
		.din(new_net_9229),
		.dout(new_net_9230)
	);

	bfr new_net_9231_bfr_after (
		.din(new_net_9230),
		.dout(new_net_9231)
	);

	bfr new_net_9232_bfr_after (
		.din(new_net_9231),
		.dout(new_net_9232)
	);

	bfr new_net_9233_bfr_after (
		.din(new_net_9232),
		.dout(new_net_9233)
	);

	bfr new_net_9234_bfr_after (
		.din(new_net_9233),
		.dout(new_net_9234)
	);

	bfr new_net_9235_bfr_after (
		.din(new_net_9234),
		.dout(new_net_9235)
	);

	bfr new_net_9236_bfr_after (
		.din(new_net_9235),
		.dout(new_net_9236)
	);

	bfr new_net_9237_bfr_after (
		.din(new_net_9236),
		.dout(new_net_9237)
	);

	bfr new_net_9238_bfr_after (
		.din(new_net_9237),
		.dout(new_net_9238)
	);

	bfr new_net_9239_bfr_after (
		.din(new_net_9238),
		.dout(new_net_9239)
	);

	bfr new_net_9240_bfr_after (
		.din(new_net_9239),
		.dout(new_net_9240)
	);

	bfr new_net_9241_bfr_after (
		.din(new_net_9240),
		.dout(new_net_9241)
	);

	bfr new_net_9242_bfr_after (
		.din(new_net_9241),
		.dout(new_net_9242)
	);

	bfr new_net_9243_bfr_after (
		.din(new_net_9242),
		.dout(new_net_9243)
	);

	bfr new_net_9244_bfr_after (
		.din(new_net_9243),
		.dout(new_net_9244)
	);

	bfr new_net_9245_bfr_after (
		.din(new_net_9244),
		.dout(new_net_9245)
	);

	bfr new_net_9246_bfr_after (
		.din(new_net_9245),
		.dout(new_net_9246)
	);

	bfr new_net_9247_bfr_after (
		.din(new_net_9246),
		.dout(new_net_9247)
	);

	bfr new_net_9248_bfr_after (
		.din(new_net_9247),
		.dout(new_net_9248)
	);

	bfr new_net_9249_bfr_after (
		.din(new_net_9248),
		.dout(new_net_9249)
	);

	bfr new_net_9250_bfr_after (
		.din(new_net_9249),
		.dout(new_net_9250)
	);

	bfr new_net_9251_bfr_after (
		.din(new_net_9250),
		.dout(new_net_9251)
	);

	bfr new_net_9252_bfr_after (
		.din(new_net_9251),
		.dout(new_net_9252)
	);

	bfr new_net_9253_bfr_after (
		.din(new_net_9252),
		.dout(new_net_9253)
	);

	bfr new_net_9254_bfr_after (
		.din(new_net_9253),
		.dout(new_net_9254)
	);

	bfr new_net_9255_bfr_after (
		.din(new_net_9254),
		.dout(new_net_9255)
	);

	bfr new_net_9256_bfr_after (
		.din(new_net_9255),
		.dout(new_net_9256)
	);

	bfr new_net_9257_bfr_after (
		.din(new_net_9256),
		.dout(new_net_9257)
	);

	bfr N1781_bfr_after (
		.din(new_net_9257),
		.dout(N1781)
	);

	bfr new_net_2242_bfr_after (
		.din(n_0825_),
		.dout(new_net_2242)
	);

	bfr new_net_9258_bfr_after (
		.din(N234),
		.dout(new_net_9258)
	);

	bfr new_net_9259_bfr_after (
		.din(new_net_9258),
		.dout(new_net_9259)
	);

	bfr new_net_9260_bfr_after (
		.din(new_net_9259),
		.dout(new_net_9260)
	);

	bfr new_net_2237_bfr_after (
		.din(new_net_9260),
		.dout(new_net_2237)
	);

	bfr new_net_9261_bfr_after (
		.din(new_net_2531),
		.dout(new_net_9261)
	);

	bfr new_net_9262_bfr_after (
		.din(new_net_9261),
		.dout(new_net_9262)
	);

	bfr new_net_9263_bfr_after (
		.din(new_net_9262),
		.dout(new_net_9263)
	);

	bfr new_net_9264_bfr_after (
		.din(new_net_9263),
		.dout(new_net_9264)
	);

	bfr new_net_9265_bfr_after (
		.din(new_net_9264),
		.dout(new_net_9265)
	);

	bfr new_net_9266_bfr_after (
		.din(new_net_9265),
		.dout(new_net_9266)
	);

	bfr new_net_9267_bfr_after (
		.din(new_net_9266),
		.dout(new_net_9267)
	);

	bfr new_net_9268_bfr_after (
		.din(new_net_9267),
		.dout(new_net_9268)
	);

	bfr new_net_9269_bfr_after (
		.din(new_net_9268),
		.dout(new_net_9269)
	);

	bfr new_net_9270_bfr_after (
		.din(new_net_9269),
		.dout(new_net_9270)
	);

	bfr new_net_9271_bfr_after (
		.din(new_net_9270),
		.dout(new_net_9271)
	);

	bfr new_net_9272_bfr_after (
		.din(new_net_9271),
		.dout(new_net_9272)
	);

	bfr new_net_9273_bfr_after (
		.din(new_net_9272),
		.dout(new_net_9273)
	);

	bfr new_net_9274_bfr_after (
		.din(new_net_9273),
		.dout(new_net_9274)
	);

	bfr new_net_9275_bfr_after (
		.din(new_net_9274),
		.dout(new_net_9275)
	);

	bfr new_net_9276_bfr_after (
		.din(new_net_9275),
		.dout(new_net_9276)
	);

	bfr new_net_9277_bfr_after (
		.din(new_net_9276),
		.dout(new_net_9277)
	);

	bfr new_net_9278_bfr_after (
		.din(new_net_9277),
		.dout(new_net_9278)
	);

	bfr new_net_9279_bfr_after (
		.din(new_net_9278),
		.dout(new_net_9279)
	);

	bfr new_net_9280_bfr_after (
		.din(new_net_9279),
		.dout(new_net_9280)
	);

	bfr new_net_9281_bfr_after (
		.din(new_net_9280),
		.dout(new_net_9281)
	);

	bfr new_net_9282_bfr_after (
		.din(new_net_9281),
		.dout(new_net_9282)
	);

	bfr new_net_9283_bfr_after (
		.din(new_net_9282),
		.dout(new_net_9283)
	);

	bfr new_net_9284_bfr_after (
		.din(new_net_9283),
		.dout(new_net_9284)
	);

	bfr new_net_9285_bfr_after (
		.din(new_net_9284),
		.dout(new_net_9285)
	);

	bfr new_net_9286_bfr_after (
		.din(new_net_9285),
		.dout(new_net_9286)
	);

	bfr new_net_9287_bfr_after (
		.din(new_net_9286),
		.dout(new_net_9287)
	);

	bfr new_net_9288_bfr_after (
		.din(new_net_9287),
		.dout(new_net_9288)
	);

	bfr new_net_9289_bfr_after (
		.din(new_net_9288),
		.dout(new_net_9289)
	);

	bfr new_net_9290_bfr_after (
		.din(new_net_9289),
		.dout(new_net_9290)
	);

	bfr new_net_9291_bfr_after (
		.din(new_net_9290),
		.dout(new_net_9291)
	);

	bfr new_net_9292_bfr_after (
		.din(new_net_9291),
		.dout(new_net_9292)
	);

	bfr new_net_9293_bfr_after (
		.din(new_net_9292),
		.dout(new_net_9293)
	);

	bfr new_net_9294_bfr_after (
		.din(new_net_9293),
		.dout(new_net_9294)
	);

	bfr new_net_9295_bfr_after (
		.din(new_net_9294),
		.dout(new_net_9295)
	);

	bfr new_net_9296_bfr_after (
		.din(new_net_9295),
		.dout(new_net_9296)
	);

	bfr new_net_9297_bfr_after (
		.din(new_net_9296),
		.dout(new_net_9297)
	);

	bfr new_net_9298_bfr_after (
		.din(new_net_9297),
		.dout(new_net_9298)
	);

	bfr new_net_9299_bfr_after (
		.din(new_net_9298),
		.dout(new_net_9299)
	);

	bfr new_net_9300_bfr_after (
		.din(new_net_9299),
		.dout(new_net_9300)
	);

	bfr new_net_9301_bfr_after (
		.din(new_net_9300),
		.dout(new_net_9301)
	);

	bfr new_net_9302_bfr_after (
		.din(new_net_9301),
		.dout(new_net_9302)
	);

	bfr new_net_9303_bfr_after (
		.din(new_net_9302),
		.dout(new_net_9303)
	);

	bfr new_net_9304_bfr_after (
		.din(new_net_9303),
		.dout(new_net_9304)
	);

	bfr new_net_9305_bfr_after (
		.din(new_net_9304),
		.dout(new_net_9305)
	);

	bfr new_net_9306_bfr_after (
		.din(new_net_9305),
		.dout(new_net_9306)
	);

	bfr new_net_9307_bfr_after (
		.din(new_net_9306),
		.dout(new_net_9307)
	);

	bfr new_net_9308_bfr_after (
		.din(new_net_9307),
		.dout(new_net_9308)
	);

	bfr new_net_9309_bfr_after (
		.din(new_net_9308),
		.dout(new_net_9309)
	);

	bfr new_net_9310_bfr_after (
		.din(new_net_9309),
		.dout(new_net_9310)
	);

	bfr new_net_9311_bfr_after (
		.din(new_net_9310),
		.dout(new_net_9311)
	);

	bfr new_net_9312_bfr_after (
		.din(new_net_9311),
		.dout(new_net_9312)
	);

	bfr N10025_bfr_after (
		.din(new_net_9312),
		.dout(N10025)
	);

	bfr new_net_9313_bfr_after (
		.din(new_net_2562),
		.dout(new_net_9313)
	);

	bfr new_net_9314_bfr_after (
		.din(new_net_9313),
		.dout(new_net_9314)
	);

	bfr new_net_9315_bfr_after (
		.din(new_net_9314),
		.dout(new_net_9315)
	);

	bfr new_net_9316_bfr_after (
		.din(new_net_9315),
		.dout(new_net_9316)
	);

	bfr new_net_9317_bfr_after (
		.din(new_net_9316),
		.dout(new_net_9317)
	);

	bfr new_net_9318_bfr_after (
		.din(new_net_9317),
		.dout(new_net_9318)
	);

	bfr new_net_9319_bfr_after (
		.din(new_net_9318),
		.dout(new_net_9319)
	);

	bfr new_net_9320_bfr_after (
		.din(new_net_9319),
		.dout(new_net_9320)
	);

	bfr new_net_9321_bfr_after (
		.din(new_net_9320),
		.dout(new_net_9321)
	);

	bfr new_net_9322_bfr_after (
		.din(new_net_9321),
		.dout(new_net_9322)
	);

	bfr new_net_9323_bfr_after (
		.din(new_net_9322),
		.dout(new_net_9323)
	);

	bfr new_net_9324_bfr_after (
		.din(new_net_9323),
		.dout(new_net_9324)
	);

	bfr new_net_9325_bfr_after (
		.din(new_net_9324),
		.dout(new_net_9325)
	);

	bfr new_net_9326_bfr_after (
		.din(new_net_9325),
		.dout(new_net_9326)
	);

	bfr new_net_9327_bfr_after (
		.din(new_net_9326),
		.dout(new_net_9327)
	);

	bfr new_net_9328_bfr_after (
		.din(new_net_9327),
		.dout(new_net_9328)
	);

	bfr new_net_9329_bfr_after (
		.din(new_net_9328),
		.dout(new_net_9329)
	);

	bfr new_net_9330_bfr_after (
		.din(new_net_9329),
		.dout(new_net_9330)
	);

	bfr new_net_9331_bfr_after (
		.din(new_net_9330),
		.dout(new_net_9331)
	);

	bfr new_net_9332_bfr_after (
		.din(new_net_9331),
		.dout(new_net_9332)
	);

	bfr new_net_9333_bfr_after (
		.din(new_net_9332),
		.dout(new_net_9333)
	);

	bfr new_net_9334_bfr_after (
		.din(new_net_9333),
		.dout(new_net_9334)
	);

	bfr new_net_9335_bfr_after (
		.din(new_net_9334),
		.dout(new_net_9335)
	);

	bfr new_net_9336_bfr_after (
		.din(new_net_9335),
		.dout(new_net_9336)
	);

	bfr new_net_9337_bfr_after (
		.din(new_net_9336),
		.dout(new_net_9337)
	);

	bfr new_net_9338_bfr_after (
		.din(new_net_9337),
		.dout(new_net_9338)
	);

	bfr new_net_9339_bfr_after (
		.din(new_net_9338),
		.dout(new_net_9339)
	);

	bfr new_net_9340_bfr_after (
		.din(new_net_9339),
		.dout(new_net_9340)
	);

	bfr new_net_9341_bfr_after (
		.din(new_net_9340),
		.dout(new_net_9341)
	);

	bfr new_net_9342_bfr_after (
		.din(new_net_9341),
		.dout(new_net_9342)
	);

	bfr new_net_9343_bfr_after (
		.din(new_net_9342),
		.dout(new_net_9343)
	);

	bfr new_net_9344_bfr_after (
		.din(new_net_9343),
		.dout(new_net_9344)
	);

	bfr new_net_9345_bfr_after (
		.din(new_net_9344),
		.dout(new_net_9345)
	);

	bfr new_net_9346_bfr_after (
		.din(new_net_9345),
		.dout(new_net_9346)
	);

	bfr new_net_9347_bfr_after (
		.din(new_net_9346),
		.dout(new_net_9347)
	);

	bfr new_net_9348_bfr_after (
		.din(new_net_9347),
		.dout(new_net_9348)
	);

	bfr new_net_9349_bfr_after (
		.din(new_net_9348),
		.dout(new_net_9349)
	);

	bfr new_net_9350_bfr_after (
		.din(new_net_9349),
		.dout(new_net_9350)
	);

	bfr new_net_9351_bfr_after (
		.din(new_net_9350),
		.dout(new_net_9351)
	);

	bfr new_net_9352_bfr_after (
		.din(new_net_9351),
		.dout(new_net_9352)
	);

	bfr new_net_9353_bfr_after (
		.din(new_net_9352),
		.dout(new_net_9353)
	);

	bfr new_net_9354_bfr_after (
		.din(new_net_9353),
		.dout(new_net_9354)
	);

	bfr new_net_9355_bfr_after (
		.din(new_net_9354),
		.dout(new_net_9355)
	);

	bfr new_net_9356_bfr_after (
		.din(new_net_9355),
		.dout(new_net_9356)
	);

	bfr new_net_9357_bfr_after (
		.din(new_net_9356),
		.dout(new_net_9357)
	);

	bfr new_net_9358_bfr_after (
		.din(new_net_9357),
		.dout(new_net_9358)
	);

	bfr new_net_9359_bfr_after (
		.din(new_net_9358),
		.dout(new_net_9359)
	);

	bfr new_net_9360_bfr_after (
		.din(new_net_9359),
		.dout(new_net_9360)
	);

	bfr new_net_9361_bfr_after (
		.din(new_net_9360),
		.dout(new_net_9361)
	);

	bfr new_net_9362_bfr_after (
		.din(new_net_9361),
		.dout(new_net_9362)
	);

	bfr new_net_9363_bfr_after (
		.din(new_net_9362),
		.dout(new_net_9363)
	);

	bfr new_net_9364_bfr_after (
		.din(new_net_9363),
		.dout(new_net_9364)
	);

	bfr new_net_9365_bfr_after (
		.din(new_net_9364),
		.dout(new_net_9365)
	);

	bfr new_net_9366_bfr_after (
		.din(new_net_9365),
		.dout(new_net_9366)
	);

	bfr new_net_9367_bfr_after (
		.din(new_net_9366),
		.dout(new_net_9367)
	);

	bfr new_net_9368_bfr_after (
		.din(new_net_9367),
		.dout(new_net_9368)
	);

	bfr new_net_9369_bfr_after (
		.din(new_net_9368),
		.dout(new_net_9369)
	);

	bfr new_net_9370_bfr_after (
		.din(new_net_9369),
		.dout(new_net_9370)
	);

	bfr new_net_9371_bfr_after (
		.din(new_net_9370),
		.dout(new_net_9371)
	);

	bfr new_net_9372_bfr_after (
		.din(new_net_9371),
		.dout(new_net_9372)
	);

	bfr new_net_9373_bfr_after (
		.din(new_net_9372),
		.dout(new_net_9373)
	);

	bfr new_net_9374_bfr_after (
		.din(new_net_9373),
		.dout(new_net_9374)
	);

	bfr new_net_9375_bfr_after (
		.din(new_net_9374),
		.dout(new_net_9375)
	);

	bfr N881_bfr_after (
		.din(new_net_9375),
		.dout(N881)
	);

	bfr new_net_2454_bfr_after (
		.din(n_0430_),
		.dout(new_net_2454)
	);

	bfr new_net_9376_bfr_after (
		.din(N219),
		.dout(new_net_9376)
	);

	bfr new_net_9377_bfr_after (
		.din(new_net_9376),
		.dout(new_net_9377)
	);

	bfr new_net_9378_bfr_after (
		.din(new_net_9377),
		.dout(new_net_9378)
	);

	bfr new_net_2267_bfr_after (
		.din(new_net_9378),
		.dout(new_net_2267)
	);

	bfr new_net_2484_bfr_after (
		.din(n_0617_),
		.dout(new_net_2484)
	);

	bfr new_net_9379_bfr_after (
		.din(n_0594_),
		.dout(new_net_9379)
	);

	bfr new_net_2479_bfr_after (
		.din(new_net_9379),
		.dout(new_net_2479)
	);

	bfr new_net_9380_bfr_after (
		.din(N53),
		.dout(new_net_9380)
	);

	bfr new_net_9381_bfr_after (
		.din(new_net_9380),
		.dout(new_net_9381)
	);

	bfr new_net_9382_bfr_after (
		.din(new_net_9381),
		.dout(new_net_9382)
	);

	bfr new_net_2293_bfr_after (
		.din(new_net_9382),
		.dout(new_net_2293)
	);

	bfr new_net_9383_bfr_after (
		.din(n_1318_),
		.dout(new_net_9383)
	);

	bfr new_net_2377_bfr_after (
		.din(new_net_9383),
		.dout(new_net_2377)
	);

	bfr new_net_9384_bfr_after (
		.din(n_0483_),
		.dout(new_net_9384)
	);

	bfr new_net_9385_bfr_after (
		.din(new_net_9384),
		.dout(new_net_9385)
	);

	bfr new_net_9386_bfr_after (
		.din(new_net_9385),
		.dout(new_net_9386)
	);

	bfr new_net_9387_bfr_after (
		.din(new_net_9386),
		.dout(new_net_9387)
	);

	bfr new_net_9388_bfr_after (
		.din(new_net_9387),
		.dout(new_net_9388)
	);

	bfr new_net_9389_bfr_after (
		.din(new_net_9388),
		.dout(new_net_9389)
	);

	bfr new_net_2461_bfr_after (
		.din(new_net_9389),
		.dout(new_net_2461)
	);

	bfr new_net_2482_bfr_after (
		.din(n_0612_),
		.dout(new_net_2482)
	);

	bfr new_net_9390_bfr_after (
		.din(N83),
		.dout(new_net_9390)
	);

	bfr new_net_9391_bfr_after (
		.din(new_net_9390),
		.dout(new_net_9391)
	);

	bfr new_net_9392_bfr_after (
		.din(new_net_9391),
		.dout(new_net_9392)
	);

	bfr new_net_2314_bfr_after (
		.din(new_net_9392),
		.dout(new_net_2314)
	);

	bfr new_net_2398_bfr_after (
		.din(n_0195_),
		.dout(new_net_2398)
	);

	bfr new_net_2272_bfr_after (
		.din(n_0885_),
		.dout(new_net_2272)
	);

	bfr new_net_9393_bfr_after (
		.din(N193),
		.dout(new_net_9393)
	);

	bfr new_net_9394_bfr_after (
		.din(new_net_9393),
		.dout(new_net_9394)
	);

	bfr new_net_9395_bfr_after (
		.din(new_net_9394),
		.dout(new_net_9395)
	);

	bfr new_net_2335_bfr_after (
		.din(new_net_9395),
		.dout(new_net_2335)
	);

	bfr new_net_9396_bfr_after (
		.din(n_0262_),
		.dout(new_net_9396)
	);

	bfr new_net_2419_bfr_after (
		.din(new_net_9396),
		.dout(new_net_2419)
	);

	bfr new_net_9397_bfr_after (
		.din(n_0313_),
		.dout(new_net_9397)
	);

	bfr new_net_9398_bfr_after (
		.din(new_net_9397),
		.dout(new_net_9398)
	);

	bfr new_net_2440_bfr_after (
		.din(new_net_9398),
		.dout(new_net_2440)
	);

	bfr new_net_9399_bfr_after (
		.din(N205),
		.dout(new_net_9399)
	);

	bfr new_net_9400_bfr_after (
		.din(new_net_9399),
		.dout(new_net_9400)
	);

	bfr new_net_9401_bfr_after (
		.din(new_net_9400),
		.dout(new_net_9401)
	);

	bfr new_net_2365_bfr_after (
		.din(new_net_9401),
		.dout(new_net_2365)
	);

	bfr new_net_2428_bfr_after (
		.din(n_0286_),
		.dout(new_net_2428)
	);

	bfr new_net_2423_bfr_after (
		.din(n_0276_),
		.dout(new_net_2423)
	);

	bfr new_net_2183_bfr_after (
		.din(N57),
		.dout(new_net_2183)
	);

	bfr new_net_9402_bfr_after (
		.din(new_net_2578),
		.dout(new_net_9402)
	);

	bfr new_net_9403_bfr_after (
		.din(new_net_9402),
		.dout(new_net_9403)
	);

	bfr new_net_9404_bfr_after (
		.din(new_net_9403),
		.dout(new_net_9404)
	);

	bfr new_net_9405_bfr_after (
		.din(new_net_9404),
		.dout(new_net_9405)
	);

	bfr new_net_9406_bfr_after (
		.din(new_net_9405),
		.dout(new_net_9406)
	);

	bfr new_net_9407_bfr_after (
		.din(new_net_9406),
		.dout(new_net_9407)
	);

	bfr new_net_9408_bfr_after (
		.din(new_net_9407),
		.dout(new_net_9408)
	);

	bfr new_net_9409_bfr_after (
		.din(new_net_9408),
		.dout(new_net_9409)
	);

	bfr new_net_9410_bfr_after (
		.din(new_net_9409),
		.dout(new_net_9410)
	);

	bfr new_net_9411_bfr_after (
		.din(new_net_9410),
		.dout(new_net_9411)
	);

	bfr new_net_9412_bfr_after (
		.din(new_net_9411),
		.dout(new_net_9412)
	);

	bfr new_net_9413_bfr_after (
		.din(new_net_9412),
		.dout(new_net_9413)
	);

	bfr new_net_9414_bfr_after (
		.din(new_net_9413),
		.dout(new_net_9414)
	);

	bfr new_net_9415_bfr_after (
		.din(new_net_9414),
		.dout(new_net_9415)
	);

	bfr new_net_9416_bfr_after (
		.din(new_net_9415),
		.dout(new_net_9416)
	);

	bfr new_net_9417_bfr_after (
		.din(new_net_9416),
		.dout(new_net_9417)
	);

	bfr new_net_9418_bfr_after (
		.din(new_net_9417),
		.dout(new_net_9418)
	);

	bfr new_net_9419_bfr_after (
		.din(new_net_9418),
		.dout(new_net_9419)
	);

	bfr new_net_9420_bfr_after (
		.din(new_net_9419),
		.dout(new_net_9420)
	);

	bfr N10632_bfr_after (
		.din(new_net_9420),
		.dout(N10632)
	);

	bfr new_net_9421_bfr_after (
		.din(N207),
		.dout(new_net_9421)
	);

	bfr new_net_9422_bfr_after (
		.din(new_net_9421),
		.dout(new_net_9422)
	);

	bfr new_net_9423_bfr_after (
		.din(new_net_9422),
		.dout(new_net_9423)
	);

	bfr new_net_2361_bfr_after (
		.din(new_net_9423),
		.dout(new_net_2361)
	);

	bfr new_net_9424_bfr_after (
		.din(N77),
		.dout(new_net_9424)
	);

	bfr new_net_9425_bfr_after (
		.din(new_net_9424),
		.dout(new_net_9425)
	);

	bfr new_net_9426_bfr_after (
		.din(new_net_9425),
		.dout(new_net_9426)
	);

	bfr new_net_2304_bfr_after (
		.din(new_net_9426),
		.dout(new_net_2304)
	);

	bfr new_net_9427_bfr_after (
		.din(N78),
		.dout(new_net_9427)
	);

	bfr new_net_9428_bfr_after (
		.din(new_net_9427),
		.dout(new_net_9428)
	);

	bfr new_net_9429_bfr_after (
		.din(new_net_9428),
		.dout(new_net_9429)
	);

	bfr new_net_2299_bfr_after (
		.din(new_net_9429),
		.dout(new_net_2299)
	);

	bfr new_net_9430_bfr_after (
		.din(n_0427_),
		.dout(new_net_9430)
	);

	bfr new_net_9431_bfr_after (
		.din(new_net_9430),
		.dout(new_net_9431)
	);

	bfr new_net_9432_bfr_after (
		.din(new_net_9431),
		.dout(new_net_9432)
	);

	bfr new_net_9433_bfr_after (
		.din(new_net_9432),
		.dout(new_net_9433)
	);

	bfr new_net_9434_bfr_after (
		.din(new_net_9433),
		.dout(new_net_9434)
	);

	bfr new_net_9435_bfr_after (
		.din(new_net_9434),
		.dout(new_net_9435)
	);

	bfr new_net_9436_bfr_after (
		.din(new_net_9435),
		.dout(new_net_9436)
	);

	bfr new_net_9437_bfr_after (
		.din(new_net_9436),
		.dout(new_net_9437)
	);

	bfr new_net_9438_bfr_after (
		.din(new_net_9437),
		.dout(new_net_9438)
	);

	bfr new_net_9439_bfr_after (
		.din(new_net_9438),
		.dout(new_net_9439)
	);

	bfr new_net_9440_bfr_after (
		.din(new_net_9439),
		.dout(new_net_9440)
	);

	bfr new_net_9441_bfr_after (
		.din(new_net_9440),
		.dout(new_net_9441)
	);

	bfr new_net_9442_bfr_after (
		.din(new_net_9441),
		.dout(new_net_9442)
	);

	bfr new_net_9443_bfr_after (
		.din(new_net_9442),
		.dout(new_net_9443)
	);

	bfr new_net_9444_bfr_after (
		.din(new_net_9443),
		.dout(new_net_9444)
	);

	bfr new_net_9445_bfr_after (
		.din(new_net_9444),
		.dout(new_net_9445)
	);

	bfr new_net_2453_bfr_after (
		.din(new_net_9445),
		.dout(new_net_2453)
	);

	bfr new_net_2372_bfr_after (
		.din(n_1274_),
		.dout(new_net_2372)
	);

	bfr new_net_9446_bfr_after (
		.din(n_0306_),
		.dout(new_net_9446)
	);

	bfr new_net_9447_bfr_after (
		.din(new_net_9446),
		.dout(new_net_9447)
	);

	bfr new_net_9448_bfr_after (
		.din(new_net_9447),
		.dout(new_net_9448)
	);

	bfr new_net_9449_bfr_after (
		.din(new_net_9448),
		.dout(new_net_9449)
	);

	bfr new_net_9450_bfr_after (
		.din(new_net_9449),
		.dout(new_net_9450)
	);

	bfr new_net_9451_bfr_after (
		.din(new_net_9450),
		.dout(new_net_9451)
	);

	bfr new_net_9452_bfr_after (
		.din(new_net_9451),
		.dout(new_net_9452)
	);

	bfr new_net_9453_bfr_after (
		.din(new_net_9452),
		.dout(new_net_9453)
	);

	bfr new_net_9454_bfr_after (
		.din(new_net_9453),
		.dout(new_net_9454)
	);

	bfr new_net_9455_bfr_after (
		.din(new_net_9454),
		.dout(new_net_9455)
	);

	bfr new_net_2435_bfr_after (
		.din(new_net_9455),
		.dout(new_net_2435)
	);

	bfr new_net_9456_bfr_after (
		.din(n_0448_),
		.dout(new_net_9456)
	);

	bfr new_net_9457_bfr_after (
		.din(new_net_9456),
		.dout(new_net_9457)
	);

	bfr new_net_9458_bfr_after (
		.din(new_net_9457),
		.dout(new_net_9458)
	);

	bfr new_net_9459_bfr_after (
		.din(new_net_9458),
		.dout(new_net_9459)
	);

	bfr new_net_9460_bfr_after (
		.din(new_net_9459),
		.dout(new_net_9460)
	);

	bfr new_net_9461_bfr_after (
		.din(new_net_9460),
		.dout(new_net_9461)
	);

	bfr new_net_9462_bfr_after (
		.din(new_net_9461),
		.dout(new_net_9462)
	);

	bfr new_net_9463_bfr_after (
		.din(new_net_9462),
		.dout(new_net_9463)
	);

	bfr new_net_9464_bfr_after (
		.din(new_net_9463),
		.dout(new_net_9464)
	);

	bfr new_net_9465_bfr_after (
		.din(new_net_9464),
		.dout(new_net_9465)
	);

	bfr new_net_9466_bfr_after (
		.din(new_net_9465),
		.dout(new_net_9466)
	);

	bfr new_net_9467_bfr_after (
		.din(new_net_9466),
		.dout(new_net_9467)
	);

	bfr new_net_9468_bfr_after (
		.din(new_net_9467),
		.dout(new_net_9468)
	);

	bfr new_net_9469_bfr_after (
		.din(new_net_9468),
		.dout(new_net_9469)
	);

	bfr new_net_9470_bfr_after (
		.din(new_net_9469),
		.dout(new_net_9470)
	);

	bfr new_net_9471_bfr_after (
		.din(new_net_9470),
		.dout(new_net_9471)
	);

	bfr new_net_9472_bfr_after (
		.din(new_net_9471),
		.dout(new_net_9472)
	);

	bfr new_net_9473_bfr_after (
		.din(new_net_9472),
		.dout(new_net_9473)
	);

	bfr new_net_9474_bfr_after (
		.din(new_net_9473),
		.dout(new_net_9474)
	);

	bfr new_net_9475_bfr_after (
		.din(new_net_9474),
		.dout(new_net_9475)
	);

	bfr new_net_9476_bfr_after (
		.din(new_net_9475),
		.dout(new_net_9476)
	);

	bfr new_net_9477_bfr_after (
		.din(new_net_9476),
		.dout(new_net_9477)
	);

	bfr new_net_9478_bfr_after (
		.din(new_net_9477),
		.dout(new_net_9478)
	);

	bfr new_net_9479_bfr_after (
		.din(new_net_9478),
		.dout(new_net_9479)
	);

	bfr new_net_9480_bfr_after (
		.din(new_net_9479),
		.dout(new_net_9480)
	);

	bfr new_net_9481_bfr_after (
		.din(new_net_9480),
		.dout(new_net_9481)
	);

	bfr new_net_2456_bfr_after (
		.din(new_net_9481),
		.dout(new_net_2456)
	);

	bfr new_net_2477_bfr_after (
		.din(n_0600_),
		.dout(new_net_2477)
	);

	bfr new_net_9482_bfr_after (
		.din(N82),
		.dout(new_net_9482)
	);

	bfr new_net_9483_bfr_after (
		.din(new_net_9482),
		.dout(new_net_9483)
	);

	bfr new_net_9484_bfr_after (
		.din(new_net_9483),
		.dout(new_net_9484)
	);

	bfr new_net_2309_bfr_after (
		.din(new_net_9484),
		.dout(new_net_2309)
	);

	bfr new_net_9485_bfr_after (
		.din(n_0174_),
		.dout(new_net_9485)
	);

	bfr new_net_9486_bfr_after (
		.din(new_net_9485),
		.dout(new_net_9486)
	);

	bfr new_net_9487_bfr_after (
		.din(new_net_9486),
		.dout(new_net_9487)
	);

	bfr new_net_9488_bfr_after (
		.din(new_net_9487),
		.dout(new_net_9488)
	);

	bfr new_net_9489_bfr_after (
		.din(new_net_9488),
		.dout(new_net_9489)
	);

	bfr new_net_9490_bfr_after (
		.din(new_net_9489),
		.dout(new_net_9490)
	);

	bfr new_net_9491_bfr_after (
		.din(new_net_9490),
		.dout(new_net_9491)
	);

	bfr new_net_9492_bfr_after (
		.din(new_net_9491),
		.dout(new_net_9492)
	);

	bfr new_net_9493_bfr_after (
		.din(new_net_9492),
		.dout(new_net_9493)
	);

	bfr new_net_9494_bfr_after (
		.din(new_net_9493),
		.dout(new_net_9494)
	);

	bfr new_net_9495_bfr_after (
		.din(new_net_9494),
		.dout(new_net_9495)
	);

	bfr new_net_9496_bfr_after (
		.din(new_net_9495),
		.dout(new_net_9496)
	);

	bfr new_net_9497_bfr_after (
		.din(new_net_9496),
		.dout(new_net_9497)
	);

	bfr new_net_9498_bfr_after (
		.din(new_net_9497),
		.dout(new_net_9498)
	);

	bfr new_net_9499_bfr_after (
		.din(new_net_9498),
		.dout(new_net_9499)
	);

	bfr new_net_9500_bfr_after (
		.din(new_net_9499),
		.dout(new_net_9500)
	);

	bfr new_net_9501_bfr_after (
		.din(new_net_9500),
		.dout(new_net_9501)
	);

	bfr new_net_9502_bfr_after (
		.din(new_net_9501),
		.dout(new_net_9502)
	);

	bfr new_net_9503_bfr_after (
		.din(new_net_9502),
		.dout(new_net_9503)
	);

	bfr new_net_9504_bfr_after (
		.din(new_net_9503),
		.dout(new_net_9504)
	);

	bfr new_net_9505_bfr_after (
		.din(new_net_9504),
		.dout(new_net_9505)
	);

	bfr new_net_9506_bfr_after (
		.din(new_net_9505),
		.dout(new_net_9506)
	);

	bfr new_net_9507_bfr_after (
		.din(new_net_9506),
		.dout(new_net_9507)
	);

	bfr new_net_9508_bfr_after (
		.din(new_net_9507),
		.dout(new_net_9508)
	);

	bfr new_net_9509_bfr_after (
		.din(new_net_9508),
		.dout(new_net_9509)
	);

	bfr new_net_9510_bfr_after (
		.din(new_net_9509),
		.dout(new_net_9510)
	);

	bfr new_net_9511_bfr_after (
		.din(new_net_9510),
		.dout(new_net_9511)
	);

	bfr new_net_9512_bfr_after (
		.din(new_net_9511),
		.dout(new_net_9512)
	);

	bfr new_net_9513_bfr_after (
		.din(new_net_9512),
		.dout(new_net_9513)
	);

	bfr new_net_9514_bfr_after (
		.din(new_net_9513),
		.dout(new_net_9514)
	);

	bfr new_net_9515_bfr_after (
		.din(new_net_9514),
		.dout(new_net_9515)
	);

	bfr new_net_9516_bfr_after (
		.din(new_net_9515),
		.dout(new_net_9516)
	);

	bfr new_net_9517_bfr_after (
		.din(new_net_9516),
		.dout(new_net_9517)
	);

	bfr new_net_9518_bfr_after (
		.din(new_net_9517),
		.dout(new_net_9518)
	);

	bfr new_net_9519_bfr_after (
		.din(new_net_9518),
		.dout(new_net_9519)
	);

	bfr new_net_9520_bfr_after (
		.din(new_net_9519),
		.dout(new_net_9520)
	);

	bfr new_net_2393_bfr_after (
		.din(new_net_9520),
		.dout(new_net_2393)
	);

	bfr new_net_2414_bfr_after (
		.din(n_0247_),
		.dout(new_net_2414)
	);

	bfr new_net_9521_bfr_after (
		.din(N155),
		.dout(new_net_9521)
	);

	bfr new_net_9522_bfr_after (
		.din(new_net_9521),
		.dout(new_net_9522)
	);

	bfr new_net_9523_bfr_after (
		.din(new_net_9522),
		.dout(new_net_9523)
	);

	bfr new_net_2204_bfr_after (
		.din(new_net_9523),
		.dout(new_net_2204)
	);

	bfr new_net_9524_bfr_after (
		.din(N215),
		.dout(new_net_9524)
	);

	bfr new_net_9525_bfr_after (
		.din(new_net_9524),
		.dout(new_net_9525)
	);

	bfr new_net_9526_bfr_after (
		.din(new_net_9525),
		.dout(new_net_9526)
	);

	bfr new_net_2225_bfr_after (
		.din(new_net_9526),
		.dout(new_net_2225)
	);

	bfr new_net_9527_bfr_after (
		.din(N224),
		.dout(new_net_9527)
	);

	bfr new_net_9528_bfr_after (
		.din(new_net_9527),
		.dout(new_net_9528)
	);

	bfr new_net_9529_bfr_after (
		.din(new_net_9528),
		.dout(new_net_9529)
	);

	bfr new_net_2246_bfr_after (
		.din(new_net_9529),
		.dout(new_net_2246)
	);

	bfr new_net_9530_bfr_after (
		.din(n_0184_),
		.dout(new_net_9530)
	);

	bfr new_net_9531_bfr_after (
		.din(new_net_9530),
		.dout(new_net_9531)
	);

	bfr new_net_9532_bfr_after (
		.din(new_net_9531),
		.dout(new_net_9532)
	);

	bfr new_net_2396_bfr_after (
		.din(new_net_9532),
		.dout(new_net_2396)
	);

	bfr new_net_9533_bfr_after (
		.din(n_0171_),
		.dout(new_net_9533)
	);

	bfr new_net_9534_bfr_after (
		.din(new_net_9533),
		.dout(new_net_9534)
	);

	bfr new_net_9535_bfr_after (
		.din(new_net_9534),
		.dout(new_net_9535)
	);

	bfr new_net_9536_bfr_after (
		.din(new_net_9535),
		.dout(new_net_9536)
	);

	bfr new_net_9537_bfr_after (
		.din(new_net_9536),
		.dout(new_net_9537)
	);

	bfr new_net_9538_bfr_after (
		.din(new_net_9537),
		.dout(new_net_9538)
	);

	bfr new_net_2392_bfr_after (
		.din(new_net_9538),
		.dout(new_net_2392)
	);

	bfr new_net_2330_bfr_after (
		.din(n_1164_),
		.dout(new_net_2330)
	);

	bfr new_net_2483_bfr_after (
		.din(n_0614_),
		.dout(new_net_2483)
	);

	bfr new_net_2478_bfr_after (
		.din(n_0599_),
		.dout(new_net_2478)
	);

	bfr new_net_2360_bfr_after (
		.din(n_1247_),
		.dout(new_net_2360)
	);

	bfr new_net_9539_bfr_after (
		.din(n_0181_),
		.dout(new_net_9539)
	);

	bfr new_net_9540_bfr_after (
		.din(new_net_9539),
		.dout(new_net_9540)
	);

	bfr new_net_9541_bfr_after (
		.din(new_net_9540),
		.dout(new_net_9541)
	);

	bfr new_net_9542_bfr_after (
		.din(new_net_9541),
		.dout(new_net_9542)
	);

	bfr new_net_2401_bfr_after (
		.din(new_net_9542),
		.dout(new_net_2401)
	);

	bfr new_net_9543_bfr_after (
		.din(new_net_2576),
		.dout(new_net_9543)
	);

	bfr new_net_9544_bfr_after (
		.din(new_net_9543),
		.dout(new_net_9544)
	);

	bfr new_net_9545_bfr_after (
		.din(new_net_9544),
		.dout(new_net_9545)
	);

	bfr new_net_9546_bfr_after (
		.din(new_net_9545),
		.dout(new_net_9546)
	);

	bfr new_net_9547_bfr_after (
		.din(new_net_9546),
		.dout(new_net_9547)
	);

	bfr new_net_9548_bfr_after (
		.din(new_net_9547),
		.dout(new_net_9548)
	);

	bfr new_net_9549_bfr_after (
		.din(new_net_9548),
		.dout(new_net_9549)
	);

	bfr new_net_9550_bfr_after (
		.din(new_net_9549),
		.dout(new_net_9550)
	);

	bfr new_net_9551_bfr_after (
		.din(new_net_9550),
		.dout(new_net_9551)
	);

	bfr new_net_9552_bfr_after (
		.din(new_net_9551),
		.dout(new_net_9552)
	);

	bfr new_net_9553_bfr_after (
		.din(new_net_9552),
		.dout(new_net_9553)
	);

	bfr new_net_9554_bfr_after (
		.din(new_net_9553),
		.dout(new_net_9554)
	);

	bfr new_net_9555_bfr_after (
		.din(new_net_9554),
		.dout(new_net_9555)
	);

	bfr new_net_9556_bfr_after (
		.din(new_net_9555),
		.dout(new_net_9556)
	);

	bfr new_net_9557_bfr_after (
		.din(new_net_9556),
		.dout(new_net_9557)
	);

	bfr new_net_9558_bfr_after (
		.din(new_net_9557),
		.dout(new_net_9558)
	);

	bfr new_net_9559_bfr_after (
		.din(new_net_9558),
		.dout(new_net_9559)
	);

	bfr new_net_9560_bfr_after (
		.din(new_net_9559),
		.dout(new_net_9560)
	);

	bfr new_net_9561_bfr_after (
		.din(new_net_9560),
		.dout(new_net_9561)
	);

	bfr new_net_9562_bfr_after (
		.din(new_net_9561),
		.dout(new_net_9562)
	);

	bfr new_net_9563_bfr_after (
		.din(new_net_9562),
		.dout(new_net_9563)
	);

	bfr new_net_9564_bfr_after (
		.din(new_net_9563),
		.dout(new_net_9564)
	);

	bfr new_net_9565_bfr_after (
		.din(new_net_9564),
		.dout(new_net_9565)
	);

	bfr new_net_9566_bfr_after (
		.din(new_net_9565),
		.dout(new_net_9566)
	);

	bfr new_net_9567_bfr_after (
		.din(new_net_9566),
		.dout(new_net_9567)
	);

	bfr new_net_9568_bfr_after (
		.din(new_net_9567),
		.dout(new_net_9568)
	);

	bfr new_net_9569_bfr_after (
		.din(new_net_9568),
		.dout(new_net_9569)
	);

	bfr N10908_bfr_after (
		.din(new_net_9569),
		.dout(N10908)
	);

	bfr new_net_9570_bfr_after (
		.din(new_net_2511),
		.dout(new_net_9570)
	);

	bfr new_net_9571_bfr_after (
		.din(new_net_9570),
		.dout(new_net_9571)
	);

	bfr new_net_9572_bfr_after (
		.din(new_net_9571),
		.dout(new_net_9572)
	);

	bfr new_net_9573_bfr_after (
		.din(new_net_9572),
		.dout(new_net_9573)
	);

	bfr new_net_9574_bfr_after (
		.din(new_net_9573),
		.dout(new_net_9574)
	);

	bfr new_net_9575_bfr_after (
		.din(new_net_9574),
		.dout(new_net_9575)
	);

	bfr new_net_9576_bfr_after (
		.din(new_net_9575),
		.dout(new_net_9576)
	);

	bfr new_net_9577_bfr_after (
		.din(new_net_9576),
		.dout(new_net_9577)
	);

	bfr new_net_9578_bfr_after (
		.din(new_net_9577),
		.dout(new_net_9578)
	);

	bfr new_net_9579_bfr_after (
		.din(new_net_9578),
		.dout(new_net_9579)
	);

	bfr new_net_9580_bfr_after (
		.din(new_net_9579),
		.dout(new_net_9580)
	);

	bfr new_net_9581_bfr_after (
		.din(new_net_9580),
		.dout(new_net_9581)
	);

	bfr new_net_9582_bfr_after (
		.din(new_net_9581),
		.dout(new_net_9582)
	);

	bfr new_net_9583_bfr_after (
		.din(new_net_9582),
		.dout(new_net_9583)
	);

	bfr new_net_9584_bfr_after (
		.din(new_net_9583),
		.dout(new_net_9584)
	);

	bfr new_net_9585_bfr_after (
		.din(new_net_9584),
		.dout(new_net_9585)
	);

	bfr new_net_9586_bfr_after (
		.din(new_net_9585),
		.dout(new_net_9586)
	);

	bfr new_net_9587_bfr_after (
		.din(new_net_9586),
		.dout(new_net_9587)
	);

	bfr new_net_9588_bfr_after (
		.din(new_net_9587),
		.dout(new_net_9588)
	);

	bfr new_net_9589_bfr_after (
		.din(new_net_9588),
		.dout(new_net_9589)
	);

	bfr new_net_9590_bfr_after (
		.din(new_net_9589),
		.dout(new_net_9590)
	);

	bfr new_net_9591_bfr_after (
		.din(new_net_9590),
		.dout(new_net_9591)
	);

	bfr new_net_9592_bfr_after (
		.din(new_net_9591),
		.dout(new_net_9592)
	);

	bfr new_net_9593_bfr_after (
		.din(new_net_9592),
		.dout(new_net_9593)
	);

	bfr new_net_9594_bfr_after (
		.din(new_net_9593),
		.dout(new_net_9594)
	);

	bfr new_net_9595_bfr_after (
		.din(new_net_9594),
		.dout(new_net_9595)
	);

	bfr new_net_9596_bfr_after (
		.din(new_net_9595),
		.dout(new_net_9596)
	);

	bfr new_net_9597_bfr_after (
		.din(new_net_9596),
		.dout(new_net_9597)
	);

	bfr new_net_9598_bfr_after (
		.din(new_net_9597),
		.dout(new_net_9598)
	);

	bfr N10869_bfr_after (
		.din(new_net_9598),
		.dout(N10869)
	);

	bfr new_net_2283_bfr_after (
		.din(n_0937_),
		.dout(new_net_2283)
	);

	bfr new_net_9599_bfr_after (
		.din(N190),
		.dout(new_net_9599)
	);

	bfr new_net_9600_bfr_after (
		.din(new_net_9599),
		.dout(new_net_9600)
	);

	bfr new_net_9601_bfr_after (
		.din(new_net_9600),
		.dout(new_net_9601)
	);

	bfr new_net_2325_bfr_after (
		.din(new_net_9601),
		.dout(new_net_2325)
	);

	bfr new_net_9602_bfr_after (
		.din(N174),
		.dout(new_net_9602)
	);

	bfr new_net_9603_bfr_after (
		.din(new_net_9602),
		.dout(new_net_9603)
	);

	bfr new_net_9604_bfr_after (
		.din(new_net_9603),
		.dout(new_net_9604)
	);

	bfr new_net_2346_bfr_after (
		.din(new_net_9604),
		.dout(new_net_2346)
	);

	bfr new_net_2220_bfr_after (
		.din(n_0760_),
		.dout(new_net_2220)
	);

	bfr new_net_9605_bfr_after (
		.din(N127),
		.dout(new_net_9605)
	);

	bfr new_net_9606_bfr_after (
		.din(new_net_9605),
		.dout(new_net_9606)
	);

	bfr new_net_9607_bfr_after (
		.din(new_net_9606),
		.dout(new_net_9607)
	);

	bfr new_net_2241_bfr_after (
		.din(new_net_9607),
		.dout(new_net_2241)
	);

	bfr new_net_9608_bfr_after (
		.din(N103),
		.dout(new_net_9608)
	);

	bfr new_net_9609_bfr_after (
		.din(new_net_9608),
		.dout(new_net_9609)
	);

	bfr new_net_9610_bfr_after (
		.din(new_net_9609),
		.dout(new_net_9610)
	);

	bfr new_net_2189_bfr_after (
		.din(new_net_9610),
		.dout(new_net_2189)
	);

	bfr new_net_2199_bfr_after (
		.din(n_0687_),
		.dout(new_net_2199)
	);

	bfr new_net_9611_bfr_after (
		.din(N118),
		.dout(new_net_9611)
	);

	bfr new_net_9612_bfr_after (
		.din(new_net_9611),
		.dout(new_net_9612)
	);

	bfr new_net_9613_bfr_after (
		.din(new_net_9612),
		.dout(new_net_9613)
	);

	bfr new_net_2262_bfr_after (
		.din(new_net_9613),
		.dout(new_net_2262)
	);

	bfr new_net_9614_bfr_after (
		.din(N204),
		.dout(new_net_9614)
	);

	bfr new_net_9615_bfr_after (
		.din(new_net_9614),
		.dout(new_net_9615)
	);

	bfr new_net_9616_bfr_after (
		.din(new_net_9615),
		.dout(new_net_9616)
	);

	bfr new_net_2367_bfr_after (
		.din(new_net_9616),
		.dout(new_net_2367)
	);

	bfr new_net_2430_bfr_after (
		.din(n_0289_),
		.dout(new_net_2430)
	);

	bfr new_net_9617_bfr_after (
		.din(N151),
		.dout(new_net_9617)
	);

	bfr new_net_9618_bfr_after (
		.din(new_net_9617),
		.dout(new_net_9618)
	);

	bfr new_net_9619_bfr_after (
		.din(new_net_9618),
		.dout(new_net_9619)
	);

	bfr new_net_2209_bfr_after (
		.din(new_net_9619),
		.dout(new_net_2209)
	);

	bfr new_net_2185_bfr_after (
		.din(N134),
		.dout(new_net_2185)
	);

	bfr new_net_9620_bfr_after (
		.din(n_1142_),
		.dout(new_net_9620)
	);

	bfr new_net_9621_bfr_after (
		.din(new_net_9620),
		.dout(new_net_9621)
	);

	bfr new_net_9622_bfr_after (
		.din(new_net_9621),
		.dout(new_net_9622)
	);

	bfr new_net_2320_bfr_after (
		.din(new_net_9622),
		.dout(new_net_2320)
	);

	bfr new_net_9623_bfr_after (
		.din(n_0213_),
		.dout(new_net_9623)
	);

	bfr new_net_9624_bfr_after (
		.din(new_net_9623),
		.dout(new_net_9624)
	);

	bfr new_net_9625_bfr_after (
		.din(new_net_9624),
		.dout(new_net_9625)
	);

	bfr new_net_2404_bfr_after (
		.din(new_net_9625),
		.dout(new_net_2404)
	);

	bfr new_net_9626_bfr_after (
		.din(N138),
		.dout(new_net_9626)
	);

	bfr new_net_9627_bfr_after (
		.din(new_net_9626),
		.dout(new_net_9627)
	);

	bfr new_net_9628_bfr_after (
		.din(new_net_9627),
		.dout(new_net_9628)
	);

	bfr new_net_2215_bfr_after (
		.din(new_net_9628),
		.dout(new_net_2215)
	);

	bfr new_net_2236_bfr_after (
		.din(n_0810_),
		.dout(new_net_2236)
	);

	bfr new_net_2257_bfr_after (
		.din(n_0858_),
		.dout(new_net_2257)
	);

	bfr new_net_9629_bfr_after (
		.din(N237),
		.dout(new_net_9629)
	);

	bfr new_net_9630_bfr_after (
		.din(new_net_9629),
		.dout(new_net_9630)
	);

	bfr new_net_9631_bfr_after (
		.din(new_net_9630),
		.dout(new_net_9631)
	);

	bfr new_net_2194_bfr_after (
		.din(new_net_9631),
		.dout(new_net_2194)
	);

	bfr new_net_9632_bfr_after (
		.din(N112),
		.dout(new_net_9632)
	);

	bfr new_net_9633_bfr_after (
		.din(new_net_9632),
		.dout(new_net_9633)
	);

	bfr new_net_9634_bfr_after (
		.din(new_net_9633),
		.dout(new_net_9634)
	);

	bfr new_net_2278_bfr_after (
		.din(new_net_9634),
		.dout(new_net_2278)
	);

	bfr new_net_9635_bfr_after (
		.din(n_1149_),
		.dout(new_net_9635)
	);

	bfr new_net_9636_bfr_after (
		.din(new_net_9635),
		.dout(new_net_9636)
	);

	bfr new_net_2341_bfr_after (
		.din(new_net_9636),
		.dout(new_net_2341)
	);

	bfr new_net_2425_bfr_after (
		.din(n_0281_),
		.dout(new_net_2425)
	);

	bfr new_net_9637_bfr_after (
		.din(n_0337_),
		.dout(new_net_9637)
	);

	bfr new_net_9638_bfr_after (
		.din(new_net_9637),
		.dout(new_net_9638)
	);

	bfr new_net_9639_bfr_after (
		.din(new_net_9638),
		.dout(new_net_9639)
	);

	bfr new_net_9640_bfr_after (
		.din(new_net_9639),
		.dout(new_net_9640)
	);

	bfr new_net_9641_bfr_after (
		.din(new_net_9640),
		.dout(new_net_9641)
	);

	bfr new_net_9642_bfr_after (
		.din(new_net_9641),
		.dout(new_net_9642)
	);

	bfr new_net_2446_bfr_after (
		.din(new_net_9642),
		.dout(new_net_2446)
	);

	bfr new_net_9643_bfr_after (
		.din(new_net_2493),
		.dout(new_net_9643)
	);

	bfr new_net_9644_bfr_after (
		.din(new_net_9643),
		.dout(new_net_9644)
	);

	bfr new_net_9645_bfr_after (
		.din(new_net_9644),
		.dout(new_net_9645)
	);

	bfr new_net_9646_bfr_after (
		.din(new_net_9645),
		.dout(new_net_9646)
	);

	bfr new_net_9647_bfr_after (
		.din(new_net_9646),
		.dout(new_net_9647)
	);

	bfr new_net_9648_bfr_after (
		.din(new_net_9647),
		.dout(new_net_9648)
	);

	bfr new_net_9649_bfr_after (
		.din(new_net_9648),
		.dout(new_net_9649)
	);

	bfr new_net_9650_bfr_after (
		.din(new_net_9649),
		.dout(new_net_9650)
	);

	bfr new_net_9651_bfr_after (
		.din(new_net_9650),
		.dout(new_net_9651)
	);

	bfr new_net_9652_bfr_after (
		.din(new_net_9651),
		.dout(new_net_9652)
	);

	bfr new_net_9653_bfr_after (
		.din(new_net_9652),
		.dout(new_net_9653)
	);

	bfr new_net_9654_bfr_after (
		.din(new_net_9653),
		.dout(new_net_9654)
	);

	bfr new_net_9655_bfr_after (
		.din(new_net_9654),
		.dout(new_net_9655)
	);

	bfr new_net_9656_bfr_after (
		.din(new_net_9655),
		.dout(new_net_9656)
	);

	bfr new_net_9657_bfr_after (
		.din(new_net_9656),
		.dout(new_net_9657)
	);

	bfr new_net_9658_bfr_after (
		.din(new_net_9657),
		.dout(new_net_9658)
	);

	bfr new_net_9659_bfr_after (
		.din(new_net_9658),
		.dout(new_net_9659)
	);

	bfr new_net_9660_bfr_after (
		.din(new_net_9659),
		.dout(new_net_9660)
	);

	bfr new_net_9661_bfr_after (
		.din(new_net_9660),
		.dout(new_net_9661)
	);

	bfr new_net_9662_bfr_after (
		.din(new_net_9661),
		.dout(new_net_9662)
	);

	bfr new_net_9663_bfr_after (
		.din(new_net_9662),
		.dout(new_net_9663)
	);

	bfr new_net_9664_bfr_after (
		.din(new_net_9663),
		.dout(new_net_9664)
	);

	bfr new_net_9665_bfr_after (
		.din(new_net_9664),
		.dout(new_net_9665)
	);

	bfr new_net_9666_bfr_after (
		.din(new_net_9665),
		.dout(new_net_9666)
	);

	bfr new_net_9667_bfr_after (
		.din(new_net_9666),
		.dout(new_net_9667)
	);

	bfr new_net_9668_bfr_after (
		.din(new_net_9667),
		.dout(new_net_9668)
	);

	bfr new_net_9669_bfr_after (
		.din(new_net_9668),
		.dout(new_net_9669)
	);

	bfr new_net_9670_bfr_after (
		.din(new_net_9669),
		.dout(new_net_9670)
	);

	bfr new_net_9671_bfr_after (
		.din(new_net_9670),
		.dout(new_net_9671)
	);

	bfr new_net_9672_bfr_after (
		.din(new_net_9671),
		.dout(new_net_9672)
	);

	bfr new_net_9673_bfr_after (
		.din(new_net_9672),
		.dout(new_net_9673)
	);

	bfr new_net_9674_bfr_after (
		.din(new_net_9673),
		.dout(new_net_9674)
	);

	bfr new_net_9675_bfr_after (
		.din(new_net_9674),
		.dout(new_net_9675)
	);

	bfr new_net_9676_bfr_after (
		.din(new_net_9675),
		.dout(new_net_9676)
	);

	bfr new_net_9677_bfr_after (
		.din(new_net_9676),
		.dout(new_net_9677)
	);

	bfr new_net_9678_bfr_after (
		.din(new_net_9677),
		.dout(new_net_9678)
	);

	bfr N10353_bfr_after (
		.din(new_net_9678),
		.dout(N10353)
	);

	bfr new_net_9679_bfr_after (
		.din(new_net_2505),
		.dout(new_net_9679)
	);

	bfr new_net_9680_bfr_after (
		.din(new_net_9679),
		.dout(new_net_9680)
	);

	bfr new_net_9681_bfr_after (
		.din(new_net_9680),
		.dout(new_net_9681)
	);

	bfr new_net_9682_bfr_after (
		.din(new_net_9681),
		.dout(new_net_9682)
	);

	bfr new_net_9683_bfr_after (
		.din(new_net_9682),
		.dout(new_net_9683)
	);

	bfr new_net_9684_bfr_after (
		.din(new_net_9683),
		.dout(new_net_9684)
	);

	bfr new_net_9685_bfr_after (
		.din(new_net_9684),
		.dout(new_net_9685)
	);

	bfr new_net_9686_bfr_after (
		.din(new_net_9685),
		.dout(new_net_9686)
	);

	bfr new_net_9687_bfr_after (
		.din(new_net_9686),
		.dout(new_net_9687)
	);

	bfr new_net_9688_bfr_after (
		.din(new_net_9687),
		.dout(new_net_9688)
	);

	bfr new_net_9689_bfr_after (
		.din(new_net_9688),
		.dout(new_net_9689)
	);

	bfr new_net_9690_bfr_after (
		.din(new_net_9689),
		.dout(new_net_9690)
	);

	bfr new_net_9691_bfr_after (
		.din(new_net_9690),
		.dout(new_net_9691)
	);

	bfr new_net_9692_bfr_after (
		.din(new_net_9691),
		.dout(new_net_9692)
	);

	bfr new_net_9693_bfr_after (
		.din(new_net_9692),
		.dout(new_net_9693)
	);

	bfr N10711_bfr_after (
		.din(new_net_9693),
		.dout(N10711)
	);

	bfr new_net_9694_bfr_after (
		.din(n_0415_),
		.dout(new_net_9694)
	);

	bfr new_net_9695_bfr_after (
		.din(new_net_9694),
		.dout(new_net_9695)
	);

	bfr new_net_9696_bfr_after (
		.din(new_net_9695),
		.dout(new_net_9696)
	);

	bfr new_net_9697_bfr_after (
		.din(new_net_9696),
		.dout(new_net_9697)
	);

	bfr new_net_9698_bfr_after (
		.din(new_net_9697),
		.dout(new_net_9698)
	);

	bfr new_net_9699_bfr_after (
		.din(new_net_9698),
		.dout(new_net_9699)
	);

	bfr new_net_9700_bfr_after (
		.din(new_net_9699),
		.dout(new_net_9700)
	);

	bfr new_net_9701_bfr_after (
		.din(new_net_9700),
		.dout(new_net_9701)
	);

	bfr new_net_9702_bfr_after (
		.din(new_net_9701),
		.dout(new_net_9702)
	);

	bfr new_net_9703_bfr_after (
		.din(new_net_9702),
		.dout(new_net_9703)
	);

	bfr new_net_9704_bfr_after (
		.din(new_net_9703),
		.dout(new_net_9704)
	);

	bfr new_net_9705_bfr_after (
		.din(new_net_9704),
		.dout(new_net_9705)
	);

	bfr new_net_9706_bfr_after (
		.din(new_net_9705),
		.dout(new_net_9706)
	);

	bfr new_net_9707_bfr_after (
		.din(new_net_9706),
		.dout(new_net_9707)
	);

	bfr new_net_2451_bfr_after (
		.din(new_net_9707),
		.dout(new_net_2451)
	);

	bfr new_net_9708_bfr_after (
		.din(new_net_2517),
		.dout(new_net_9708)
	);

	bfr new_net_9709_bfr_after (
		.din(new_net_9708),
		.dout(new_net_9709)
	);

	bfr new_net_9710_bfr_after (
		.din(new_net_9709),
		.dout(new_net_9710)
	);

	bfr new_net_9711_bfr_after (
		.din(new_net_9710),
		.dout(new_net_9711)
	);

	bfr new_net_9712_bfr_after (
		.din(new_net_9711),
		.dout(new_net_9712)
	);

	bfr new_net_9713_bfr_after (
		.din(new_net_9712),
		.dout(new_net_9713)
	);

	bfr new_net_9714_bfr_after (
		.din(new_net_9713),
		.dout(new_net_9714)
	);

	bfr new_net_9715_bfr_after (
		.din(new_net_9714),
		.dout(new_net_9715)
	);

	bfr new_net_9716_bfr_after (
		.din(new_net_9715),
		.dout(new_net_9716)
	);

	bfr new_net_9717_bfr_after (
		.din(new_net_9716),
		.dout(new_net_9717)
	);

	bfr new_net_9718_bfr_after (
		.din(new_net_9717),
		.dout(new_net_9718)
	);

	bfr new_net_9719_bfr_after (
		.din(new_net_9718),
		.dout(new_net_9719)
	);

	bfr new_net_9720_bfr_after (
		.din(new_net_9719),
		.dout(new_net_9720)
	);

	bfr new_net_9721_bfr_after (
		.din(new_net_9720),
		.dout(new_net_9721)
	);

	bfr new_net_9722_bfr_after (
		.din(new_net_9721),
		.dout(new_net_9722)
	);

	bfr new_net_9723_bfr_after (
		.din(new_net_9722),
		.dout(new_net_9723)
	);

	bfr N10712_bfr_after (
		.din(new_net_9723),
		.dout(N10712)
	);

	bfr new_net_9724_bfr_after (
		.din(new_net_2523),
		.dout(new_net_9724)
	);

	bfr new_net_9725_bfr_after (
		.din(new_net_9724),
		.dout(new_net_9725)
	);

	bfr new_net_9726_bfr_after (
		.din(new_net_9725),
		.dout(new_net_9726)
	);

	bfr new_net_9727_bfr_after (
		.din(new_net_9726),
		.dout(new_net_9727)
	);

	bfr new_net_9728_bfr_after (
		.din(new_net_9727),
		.dout(new_net_9728)
	);

	bfr new_net_9729_bfr_after (
		.din(new_net_9728),
		.dout(new_net_9729)
	);

	bfr new_net_9730_bfr_after (
		.din(new_net_9729),
		.dout(new_net_9730)
	);

	bfr new_net_9731_bfr_after (
		.din(new_net_9730),
		.dout(new_net_9731)
	);

	bfr new_net_9732_bfr_after (
		.din(new_net_9731),
		.dout(new_net_9732)
	);

	bfr new_net_9733_bfr_after (
		.din(new_net_9732),
		.dout(new_net_9733)
	);

	bfr new_net_9734_bfr_after (
		.din(new_net_9733),
		.dout(new_net_9734)
	);

	bfr new_net_9735_bfr_after (
		.din(new_net_9734),
		.dout(new_net_9735)
	);

	bfr new_net_9736_bfr_after (
		.din(new_net_9735),
		.dout(new_net_9736)
	);

	bfr new_net_9737_bfr_after (
		.din(new_net_9736),
		.dout(new_net_9737)
	);

	bfr new_net_9738_bfr_after (
		.din(new_net_9737),
		.dout(new_net_9738)
	);

	bfr new_net_9739_bfr_after (
		.din(new_net_9738),
		.dout(new_net_9739)
	);

	bfr new_net_9740_bfr_after (
		.din(new_net_9739),
		.dout(new_net_9740)
	);

	bfr new_net_9741_bfr_after (
		.din(new_net_9740),
		.dout(new_net_9741)
	);

	bfr new_net_9742_bfr_after (
		.din(new_net_9741),
		.dout(new_net_9742)
	);

	bfr new_net_9743_bfr_after (
		.din(new_net_9742),
		.dout(new_net_9743)
	);

	bfr new_net_9744_bfr_after (
		.din(new_net_9743),
		.dout(new_net_9744)
	);

	bfr new_net_9745_bfr_after (
		.din(new_net_9744),
		.dout(new_net_9745)
	);

	bfr new_net_9746_bfr_after (
		.din(new_net_9745),
		.dout(new_net_9746)
	);

	bfr new_net_9747_bfr_after (
		.din(new_net_9746),
		.dout(new_net_9747)
	);

	bfr new_net_9748_bfr_after (
		.din(new_net_9747),
		.dout(new_net_9748)
	);

	bfr new_net_9749_bfr_after (
		.din(new_net_9748),
		.dout(new_net_9749)
	);

	bfr new_net_9750_bfr_after (
		.din(new_net_9749),
		.dout(new_net_9750)
	);

	bfr N10870_bfr_after (
		.din(new_net_9750),
		.dout(N10870)
	);

	bfr N11334_bfr_after (
		.din(new_net_2529),
		.dout(N11334)
	);

	bfr new_net_9751_bfr_after (
		.din(new_net_2541),
		.dout(new_net_9751)
	);

	bfr new_net_9752_bfr_after (
		.din(new_net_9751),
		.dout(new_net_9752)
	);

	bfr new_net_9753_bfr_after (
		.din(new_net_9752),
		.dout(new_net_9753)
	);

	bfr new_net_9754_bfr_after (
		.din(new_net_9753),
		.dout(new_net_9754)
	);

	bfr new_net_9755_bfr_after (
		.din(new_net_9754),
		.dout(new_net_9755)
	);

	bfr new_net_9756_bfr_after (
		.din(new_net_9755),
		.dout(new_net_9756)
	);

	bfr new_net_9757_bfr_after (
		.din(new_net_9756),
		.dout(new_net_9757)
	);

	bfr new_net_9758_bfr_after (
		.din(new_net_9757),
		.dout(new_net_9758)
	);

	bfr new_net_9759_bfr_after (
		.din(new_net_9758),
		.dout(new_net_9759)
	);

	bfr new_net_9760_bfr_after (
		.din(new_net_9759),
		.dout(new_net_9760)
	);

	bfr new_net_9761_bfr_after (
		.din(new_net_9760),
		.dout(new_net_9761)
	);

	bfr new_net_9762_bfr_after (
		.din(new_net_9761),
		.dout(new_net_9762)
	);

	bfr new_net_9763_bfr_after (
		.din(new_net_9762),
		.dout(new_net_9763)
	);

	bfr new_net_9764_bfr_after (
		.din(new_net_9763),
		.dout(new_net_9764)
	);

	bfr new_net_9765_bfr_after (
		.din(new_net_9764),
		.dout(new_net_9765)
	);

	bfr new_net_9766_bfr_after (
		.din(new_net_9765),
		.dout(new_net_9766)
	);

	bfr new_net_9767_bfr_after (
		.din(new_net_9766),
		.dout(new_net_9767)
	);

	bfr new_net_9768_bfr_after (
		.din(new_net_9767),
		.dout(new_net_9768)
	);

	bfr new_net_9769_bfr_after (
		.din(new_net_9768),
		.dout(new_net_9769)
	);

	bfr new_net_9770_bfr_after (
		.din(new_net_9769),
		.dout(new_net_9770)
	);

	bfr new_net_9771_bfr_after (
		.din(new_net_9770),
		.dout(new_net_9771)
	);

	bfr new_net_9772_bfr_after (
		.din(new_net_9771),
		.dout(new_net_9772)
	);

	bfr new_net_9773_bfr_after (
		.din(new_net_9772),
		.dout(new_net_9773)
	);

	bfr new_net_9774_bfr_after (
		.din(new_net_9773),
		.dout(new_net_9774)
	);

	bfr new_net_9775_bfr_after (
		.din(new_net_9774),
		.dout(new_net_9775)
	);

	bfr new_net_9776_bfr_after (
		.din(new_net_9775),
		.dout(new_net_9776)
	);

	bfr new_net_9777_bfr_after (
		.din(new_net_9776),
		.dout(new_net_9777)
	);

	bfr new_net_9778_bfr_after (
		.din(new_net_9777),
		.dout(new_net_9778)
	);

	bfr new_net_9779_bfr_after (
		.din(new_net_9778),
		.dout(new_net_9779)
	);

	bfr new_net_9780_bfr_after (
		.din(new_net_9779),
		.dout(new_net_9780)
	);

	bfr new_net_9781_bfr_after (
		.din(new_net_9780),
		.dout(new_net_9781)
	);

	bfr N11342_bfr_after (
		.din(new_net_9781),
		.dout(N11342)
	);

	bfr new_net_9782_bfr_after (
		.din(new_net_2543),
		.dout(new_net_9782)
	);

	bfr new_net_9783_bfr_after (
		.din(new_net_9782),
		.dout(new_net_9783)
	);

	bfr new_net_9784_bfr_after (
		.din(new_net_9783),
		.dout(new_net_9784)
	);

	bfr new_net_9785_bfr_after (
		.din(new_net_9784),
		.dout(new_net_9785)
	);

	bfr new_net_9786_bfr_after (
		.din(new_net_9785),
		.dout(new_net_9786)
	);

	bfr new_net_9787_bfr_after (
		.din(new_net_9786),
		.dout(new_net_9787)
	);

	bfr new_net_9788_bfr_after (
		.din(new_net_9787),
		.dout(new_net_9788)
	);

	bfr new_net_9789_bfr_after (
		.din(new_net_9788),
		.dout(new_net_9789)
	);

	bfr new_net_9790_bfr_after (
		.din(new_net_9789),
		.dout(new_net_9790)
	);

	bfr new_net_9791_bfr_after (
		.din(new_net_9790),
		.dout(new_net_9791)
	);

	bfr new_net_9792_bfr_after (
		.din(new_net_9791),
		.dout(new_net_9792)
	);

	bfr new_net_9793_bfr_after (
		.din(new_net_9792),
		.dout(new_net_9793)
	);

	bfr new_net_9794_bfr_after (
		.din(new_net_9793),
		.dout(new_net_9794)
	);

	bfr new_net_9795_bfr_after (
		.din(new_net_9794),
		.dout(new_net_9795)
	);

	bfr new_net_9796_bfr_after (
		.din(new_net_9795),
		.dout(new_net_9796)
	);

	bfr new_net_9797_bfr_after (
		.din(new_net_9796),
		.dout(new_net_9797)
	);

	bfr new_net_9798_bfr_after (
		.din(new_net_9797),
		.dout(new_net_9798)
	);

	bfr new_net_9799_bfr_after (
		.din(new_net_9798),
		.dout(new_net_9799)
	);

	bfr new_net_9800_bfr_after (
		.din(new_net_9799),
		.dout(new_net_9800)
	);

	bfr new_net_9801_bfr_after (
		.din(new_net_9800),
		.dout(new_net_9801)
	);

	bfr new_net_9802_bfr_after (
		.din(new_net_9801),
		.dout(new_net_9802)
	);

	bfr new_net_9803_bfr_after (
		.din(new_net_9802),
		.dout(new_net_9803)
	);

	bfr new_net_9804_bfr_after (
		.din(new_net_9803),
		.dout(new_net_9804)
	);

	bfr new_net_9805_bfr_after (
		.din(new_net_9804),
		.dout(new_net_9805)
	);

	bfr new_net_9806_bfr_after (
		.din(new_net_9805),
		.dout(new_net_9806)
	);

	bfr new_net_9807_bfr_after (
		.din(new_net_9806),
		.dout(new_net_9807)
	);

	bfr new_net_9808_bfr_after (
		.din(new_net_9807),
		.dout(new_net_9808)
	);

	bfr new_net_9809_bfr_after (
		.din(new_net_9808),
		.dout(new_net_9809)
	);

	bfr new_net_9810_bfr_after (
		.din(new_net_9809),
		.dout(new_net_9810)
	);

	bfr new_net_9811_bfr_after (
		.din(new_net_9810),
		.dout(new_net_9811)
	);

	bfr new_net_9812_bfr_after (
		.din(new_net_9811),
		.dout(new_net_9812)
	);

	bfr N10868_bfr_after (
		.din(new_net_9812),
		.dout(N10868)
	);

	bfr new_net_9813_bfr_after (
		.din(n_0597_),
		.dout(new_net_9813)
	);

	bfr new_net_2476_bfr_after (
		.din(new_net_9813),
		.dout(new_net_2476)
	);

	bfr new_net_2233_bfr_after (
		.din(n_0805_),
		.dout(new_net_2233)
	);

	bfr new_net_9814_bfr_after (
		.din(N170),
		.dout(new_net_9814)
	);

	bfr new_net_9815_bfr_after (
		.din(new_net_9814),
		.dout(new_net_9815)
	);

	bfr new_net_9816_bfr_after (
		.din(new_net_9815),
		.dout(new_net_9816)
	);

	bfr new_net_9817_bfr_after (
		.din(new_net_9816),
		.dout(new_net_9817)
	);

	bfr new_net_9818_bfr_after (
		.din(new_net_9817),
		.dout(new_net_9818)
	);

	bfr new_net_9819_bfr_after (
		.din(new_net_9818),
		.dout(new_net_9819)
	);

	bfr new_net_2315_bfr_after (
		.din(new_net_9819),
		.dout(new_net_2315)
	);

	bfr new_net_9820_bfr_after (
		.din(n_0199_),
		.dout(new_net_9820)
	);

	bfr new_net_2399_bfr_after (
		.din(new_net_9820),
		.dout(new_net_2399)
	);

	bfr new_net_2336_bfr_after (
		.din(n_1179_),
		.dout(new_net_2336)
	);

	bfr new_net_9821_bfr_after (
		.din(n_0263_),
		.dout(new_net_9821)
	);

	bfr new_net_9822_bfr_after (
		.din(new_net_9821),
		.dout(new_net_9822)
	);

	bfr new_net_9823_bfr_after (
		.din(new_net_9822),
		.dout(new_net_9823)
	);

	bfr new_net_9824_bfr_after (
		.din(new_net_9823),
		.dout(new_net_9824)
	);

	bfr new_net_9825_bfr_after (
		.din(new_net_9824),
		.dout(new_net_9825)
	);

	bfr new_net_2420_bfr_after (
		.din(new_net_9825),
		.dout(new_net_2420)
	);

	bfr new_net_2441_bfr_after (
		.din(n_0322_),
		.dout(new_net_2441)
	);

	bfr new_net_2231_bfr_after (
		.din(n_0802_),
		.dout(new_net_2231)
	);

	bfr new_net_9826_bfr_after (
		.din(N226),
		.dout(new_net_9826)
	);

	bfr new_net_9827_bfr_after (
		.din(new_net_9826),
		.dout(new_net_9827)
	);

	bfr new_net_9828_bfr_after (
		.din(new_net_9827),
		.dout(new_net_9828)
	);

	bfr new_net_2252_bfr_after (
		.din(new_net_9828),
		.dout(new_net_2252)
	);

	bfr new_net_2210_bfr_after (
		.din(n_0737_),
		.dout(new_net_2210)
	);

	bfr new_net_9829_bfr_after (
		.din(N221),
		.dout(new_net_9829)
	);

	bfr new_net_9830_bfr_after (
		.din(new_net_9829),
		.dout(new_net_9830)
	);

	bfr new_net_9831_bfr_after (
		.din(new_net_9830),
		.dout(new_net_9831)
	);

	bfr new_net_2273_bfr_after (
		.din(new_net_9831),
		.dout(new_net_2273)
	);

	bfr new_net_9832_bfr_after (
		.din(n_0948_),
		.dout(new_net_9832)
	);

	bfr new_net_9833_bfr_after (
		.din(new_net_9832),
		.dout(new_net_9833)
	);

	bfr new_net_2294_bfr_after (
		.din(new_net_9833),
		.dout(new_net_2294)
	);

	bfr new_net_2450_bfr_after (
		.din(n_0397_),
		.dout(new_net_2450)
	);

	bfr new_net_2445_bfr_after (
		.din(n_0334_),
		.dout(new_net_2445)
	);

	bfr new_net_2263_bfr_after (
		.din(n_0870_),
		.dout(new_net_2263)
	);

	bfr N10104_bfr_after (
		.din(new_net_2554),
		.dout(N10104)
	);

	bfr new_net_9834_bfr_after (
		.din(N66),
		.dout(new_net_9834)
	);

	bfr new_net_9835_bfr_after (
		.din(new_net_9834),
		.dout(new_net_9835)
	);

	bfr new_net_9836_bfr_after (
		.din(new_net_9835),
		.dout(new_net_9836)
	);

	bfr new_net_2268_bfr_after (
		.din(new_net_9836),
		.dout(new_net_2268)
	);

	bfr new_net_9837_bfr_after (
		.din(N65),
		.dout(new_net_9837)
	);

	bfr new_net_9838_bfr_after (
		.din(new_net_9837),
		.dout(new_net_9838)
	);

	bfr new_net_9839_bfr_after (
		.din(new_net_9838),
		.dout(new_net_9839)
	);

	bfr new_net_2310_bfr_after (
		.din(new_net_9839),
		.dout(new_net_2310)
	);

	bfr new_net_9840_bfr_after (
		.din(n_0165_),
		.dout(new_net_9840)
	);

	bfr new_net_9841_bfr_after (
		.din(new_net_9840),
		.dout(new_net_9841)
	);

	bfr new_net_9842_bfr_after (
		.din(new_net_9841),
		.dout(new_net_9842)
	);

	bfr new_net_9843_bfr_after (
		.din(new_net_9842),
		.dout(new_net_9843)
	);

	bfr new_net_9844_bfr_after (
		.din(new_net_9843),
		.dout(new_net_9844)
	);

	bfr new_net_9845_bfr_after (
		.din(new_net_9844),
		.dout(new_net_9845)
	);

	bfr new_net_9846_bfr_after (
		.din(new_net_9845),
		.dout(new_net_9846)
	);

	bfr new_net_9847_bfr_after (
		.din(new_net_9846),
		.dout(new_net_9847)
	);

	bfr new_net_9848_bfr_after (
		.din(new_net_9847),
		.dout(new_net_9848)
	);

	bfr new_net_9849_bfr_after (
		.din(new_net_9848),
		.dout(new_net_9849)
	);

	bfr new_net_9850_bfr_after (
		.din(new_net_9849),
		.dout(new_net_9850)
	);

	bfr new_net_9851_bfr_after (
		.din(new_net_9850),
		.dout(new_net_9851)
	);

	bfr new_net_9852_bfr_after (
		.din(new_net_9851),
		.dout(new_net_9852)
	);

	bfr new_net_9853_bfr_after (
		.din(new_net_9852),
		.dout(new_net_9853)
	);

	bfr new_net_9854_bfr_after (
		.din(new_net_9853),
		.dout(new_net_9854)
	);

	bfr new_net_9855_bfr_after (
		.din(new_net_9854),
		.dout(new_net_9855)
	);

	bfr new_net_9856_bfr_after (
		.din(new_net_9855),
		.dout(new_net_9856)
	);

	bfr new_net_9857_bfr_after (
		.din(new_net_9856),
		.dout(new_net_9857)
	);

	bfr new_net_9858_bfr_after (
		.din(new_net_9857),
		.dout(new_net_9858)
	);

	bfr new_net_9859_bfr_after (
		.din(new_net_9858),
		.dout(new_net_9859)
	);

	bfr new_net_9860_bfr_after (
		.din(new_net_9859),
		.dout(new_net_9860)
	);

	bfr new_net_9861_bfr_after (
		.din(new_net_9860),
		.dout(new_net_9861)
	);

	bfr new_net_9862_bfr_after (
		.din(new_net_9861),
		.dout(new_net_9862)
	);

	bfr new_net_9863_bfr_after (
		.din(new_net_9862),
		.dout(new_net_9863)
	);

	bfr new_net_9864_bfr_after (
		.din(new_net_9863),
		.dout(new_net_9864)
	);

	bfr new_net_9865_bfr_after (
		.din(new_net_9864),
		.dout(new_net_9865)
	);

	bfr new_net_9866_bfr_after (
		.din(new_net_9865),
		.dout(new_net_9866)
	);

	bfr new_net_9867_bfr_after (
		.din(new_net_9866),
		.dout(new_net_9867)
	);

	bfr new_net_9868_bfr_after (
		.din(new_net_9867),
		.dout(new_net_9868)
	);

	bfr new_net_9869_bfr_after (
		.din(new_net_9868),
		.dout(new_net_9869)
	);

	bfr new_net_9870_bfr_after (
		.din(new_net_9869),
		.dout(new_net_9870)
	);

	bfr new_net_9871_bfr_after (
		.din(new_net_9870),
		.dout(new_net_9871)
	);

	bfr new_net_9872_bfr_after (
		.din(new_net_9871),
		.dout(new_net_9872)
	);

	bfr new_net_9873_bfr_after (
		.din(new_net_9872),
		.dout(new_net_9873)
	);

	bfr new_net_9874_bfr_after (
		.din(new_net_9873),
		.dout(new_net_9874)
	);

	bfr new_net_9875_bfr_after (
		.din(new_net_9874),
		.dout(new_net_9875)
	);

	bfr new_net_9876_bfr_after (
		.din(new_net_9875),
		.dout(new_net_9876)
	);

	bfr new_net_9877_bfr_after (
		.din(new_net_9876),
		.dout(new_net_9877)
	);

	bfr new_net_9878_bfr_after (
		.din(new_net_9877),
		.dout(new_net_9878)
	);

	bfr new_net_9879_bfr_after (
		.din(new_net_9878),
		.dout(new_net_9879)
	);

	bfr new_net_9880_bfr_after (
		.din(new_net_9879),
		.dout(new_net_9880)
	);

	bfr new_net_9881_bfr_after (
		.din(new_net_9880),
		.dout(new_net_9881)
	);

	bfr new_net_9882_bfr_after (
		.din(new_net_9881),
		.dout(new_net_9882)
	);

	bfr new_net_9883_bfr_after (
		.din(new_net_9882),
		.dout(new_net_9883)
	);

	bfr new_net_9884_bfr_after (
		.din(new_net_9883),
		.dout(new_net_9884)
	);

	bfr new_net_9885_bfr_after (
		.din(new_net_9884),
		.dout(new_net_9885)
	);

	bfr new_net_9886_bfr_after (
		.din(new_net_9885),
		.dout(new_net_9886)
	);

	bfr new_net_9887_bfr_after (
		.din(new_net_9886),
		.dout(new_net_9887)
	);

	bfr new_net_9888_bfr_after (
		.din(new_net_9887),
		.dout(new_net_9888)
	);

	bfr new_net_9889_bfr_after (
		.din(new_net_9888),
		.dout(new_net_9889)
	);

	bfr new_net_9890_bfr_after (
		.din(new_net_9889),
		.dout(new_net_9890)
	);

	bfr new_net_9891_bfr_after (
		.din(new_net_9890),
		.dout(new_net_9891)
	);

	bfr new_net_9892_bfr_after (
		.din(new_net_9891),
		.dout(new_net_9892)
	);

	bfr new_net_9893_bfr_after (
		.din(new_net_9892),
		.dout(new_net_9893)
	);

	bfr new_net_9894_bfr_after (
		.din(new_net_9893),
		.dout(new_net_9894)
	);

	bfr new_net_9895_bfr_after (
		.din(new_net_9894),
		.dout(new_net_9895)
	);

	bfr new_net_2394_bfr_after (
		.din(new_net_9895),
		.dout(new_net_2394)
	);

	bfr new_net_2415_bfr_after (
		.din(n_0254_),
		.dout(new_net_2415)
	);

	bfr new_net_9896_bfr_after (
		.din(N141),
		.dout(new_net_9896)
	);

	bfr new_net_9897_bfr_after (
		.din(new_net_9896),
		.dout(new_net_9897)
	);

	bfr new_net_9898_bfr_after (
		.din(new_net_9897),
		.dout(new_net_9898)
	);

	bfr new_net_2205_bfr_after (
		.din(new_net_9898),
		.dout(new_net_2205)
	);

	bfr new_net_9899_bfr_after (
		.din(n_0791_),
		.dout(new_net_9899)
	);

	bfr new_net_9900_bfr_after (
		.din(new_net_9899),
		.dout(new_net_9900)
	);

	bfr new_net_9901_bfr_after (
		.din(new_net_9900),
		.dout(new_net_9901)
	);

	bfr new_net_2226_bfr_after (
		.din(new_net_9901),
		.dout(new_net_2226)
	);

	bfr new_net_9902_bfr_after (
		.din(N121),
		.dout(new_net_9902)
	);

	bfr new_net_9903_bfr_after (
		.din(new_net_9902),
		.dout(new_net_9903)
	);

	bfr new_net_9904_bfr_after (
		.din(new_net_9903),
		.dout(new_net_9904)
	);

	bfr new_net_2247_bfr_after (
		.din(new_net_9904),
		.dout(new_net_2247)
	);

	bfr new_net_2475_bfr_after (
		.din(n_0586_),
		.dout(new_net_2475)
	);

	bfr new_net_9905_bfr_after (
		.din(N56),
		.dout(new_net_9905)
	);

	bfr new_net_9906_bfr_after (
		.din(new_net_9905),
		.dout(new_net_9906)
	);

	bfr new_net_9907_bfr_after (
		.din(new_net_9906),
		.dout(new_net_9907)
	);

	bfr new_net_2289_bfr_after (
		.din(new_net_9907),
		.dout(new_net_2289)
	);

	bfr new_net_9908_bfr_after (
		.din(N191),
		.dout(new_net_9908)
	);

	bfr new_net_9909_bfr_after (
		.din(new_net_9908),
		.dout(new_net_9909)
	);

	bfr new_net_9910_bfr_after (
		.din(new_net_9909),
		.dout(new_net_9910)
	);

	bfr new_net_2331_bfr_after (
		.din(new_net_9910),
		.dout(new_net_2331)
	);

	bfr new_net_9911_bfr_after (
		.din(N208),
		.dout(new_net_9911)
	);

	bfr new_net_9912_bfr_after (
		.din(new_net_9911),
		.dout(new_net_9912)
	);

	bfr new_net_9913_bfr_after (
		.din(new_net_9912),
		.dout(new_net_9913)
	);

	bfr new_net_2357_bfr_after (
		.din(new_net_9913),
		.dout(new_net_2357)
	);

	bfr new_net_9914_bfr_after (
		.din(N177),
		.dout(new_net_9914)
	);

	bfr new_net_9915_bfr_after (
		.din(new_net_9914),
		.dout(new_net_9915)
	);

	bfr new_net_9916_bfr_after (
		.din(new_net_9915),
		.dout(new_net_9916)
	);

	bfr new_net_2352_bfr_after (
		.din(new_net_9916),
		.dout(new_net_2352)
	);

	bfr new_net_9917_bfr_after (
		.din(new_net_2568),
		.dout(new_net_9917)
	);

	bfr new_net_9918_bfr_after (
		.din(new_net_9917),
		.dout(new_net_9918)
	);

	bfr new_net_9919_bfr_after (
		.din(new_net_9918),
		.dout(new_net_9919)
	);

	bfr new_net_9920_bfr_after (
		.din(new_net_9919),
		.dout(new_net_9920)
	);

	bfr new_net_9921_bfr_after (
		.din(new_net_9920),
		.dout(new_net_9921)
	);

	bfr new_net_9922_bfr_after (
		.din(new_net_9921),
		.dout(new_net_9922)
	);

	bfr new_net_9923_bfr_after (
		.din(new_net_9922),
		.dout(new_net_9923)
	);

	bfr new_net_9924_bfr_after (
		.din(new_net_9923),
		.dout(new_net_9924)
	);

	bfr new_net_9925_bfr_after (
		.din(new_net_9924),
		.dout(new_net_9925)
	);

	bfr new_net_9926_bfr_after (
		.din(new_net_9925),
		.dout(new_net_9926)
	);

	bfr new_net_9927_bfr_after (
		.din(new_net_9926),
		.dout(new_net_9927)
	);

	bfr new_net_9928_bfr_after (
		.din(new_net_9927),
		.dout(new_net_9928)
	);

	bfr new_net_9929_bfr_after (
		.din(new_net_9928),
		.dout(new_net_9929)
	);

	bfr new_net_9930_bfr_after (
		.din(new_net_9929),
		.dout(new_net_9930)
	);

	bfr new_net_9931_bfr_after (
		.din(new_net_9930),
		.dout(new_net_9931)
	);

	bfr new_net_9932_bfr_after (
		.din(new_net_9931),
		.dout(new_net_9932)
	);

	bfr new_net_9933_bfr_after (
		.din(new_net_9932),
		.dout(new_net_9933)
	);

	bfr new_net_9934_bfr_after (
		.din(new_net_9933),
		.dout(new_net_9934)
	);

	bfr new_net_9935_bfr_after (
		.din(new_net_9934),
		.dout(new_net_9935)
	);

	bfr new_net_9936_bfr_after (
		.din(new_net_9935),
		.dout(new_net_9936)
	);

	bfr new_net_9937_bfr_after (
		.din(new_net_9936),
		.dout(new_net_9937)
	);

	bfr new_net_9938_bfr_after (
		.din(new_net_9937),
		.dout(new_net_9938)
	);

	bfr new_net_9939_bfr_after (
		.din(new_net_9938),
		.dout(new_net_9939)
	);

	bfr new_net_9940_bfr_after (
		.din(new_net_9939),
		.dout(new_net_9940)
	);

	bfr new_net_9941_bfr_after (
		.din(new_net_9940),
		.dout(new_net_9941)
	);

	bfr new_net_9942_bfr_after (
		.din(new_net_9941),
		.dout(new_net_9942)
	);

	bfr new_net_9943_bfr_after (
		.din(new_net_9942),
		.dout(new_net_9943)
	);

	bfr new_net_9944_bfr_after (
		.din(new_net_9943),
		.dout(new_net_9944)
	);

	bfr new_net_9945_bfr_after (
		.din(new_net_9944),
		.dout(new_net_9945)
	);

	bfr new_net_9946_bfr_after (
		.din(new_net_9945),
		.dout(new_net_9946)
	);

	bfr new_net_9947_bfr_after (
		.din(new_net_9946),
		.dout(new_net_9947)
	);

	bfr new_net_9948_bfr_after (
		.din(new_net_9947),
		.dout(new_net_9948)
	);

	bfr new_net_9949_bfr_after (
		.din(new_net_9948),
		.dout(new_net_9949)
	);

	bfr new_net_9950_bfr_after (
		.din(new_net_9949),
		.dout(new_net_9950)
	);

	bfr new_net_9951_bfr_after (
		.din(new_net_9950),
		.dout(new_net_9951)
	);

	bfr new_net_9952_bfr_after (
		.din(new_net_9951),
		.dout(new_net_9952)
	);

	bfr new_net_9953_bfr_after (
		.din(new_net_9952),
		.dout(new_net_9953)
	);

	bfr new_net_9954_bfr_after (
		.din(new_net_9953),
		.dout(new_net_9954)
	);

	bfr new_net_9955_bfr_after (
		.din(new_net_9954),
		.dout(new_net_9955)
	);

	bfr new_net_9956_bfr_after (
		.din(new_net_9955),
		.dout(new_net_9956)
	);

	bfr new_net_9957_bfr_after (
		.din(new_net_9956),
		.dout(new_net_9957)
	);

	bfr new_net_9958_bfr_after (
		.din(new_net_9957),
		.dout(new_net_9958)
	);

	bfr N10109_bfr_after (
		.din(new_net_9958),
		.dout(N10109)
	);

	bfr new_net_2449_bfr_after (
		.din(n_0381_),
		.dout(new_net_2449)
	);

	bfr new_net_9959_bfr_after (
		.din(n_0331_),
		.dout(new_net_9959)
	);

	bfr new_net_9960_bfr_after (
		.din(new_net_9959),
		.dout(new_net_9960)
	);

	bfr new_net_9961_bfr_after (
		.din(new_net_9960),
		.dout(new_net_9961)
	);

	bfr new_net_9962_bfr_after (
		.din(new_net_9961),
		.dout(new_net_9962)
	);

	bfr new_net_9963_bfr_after (
		.din(new_net_9962),
		.dout(new_net_9963)
	);

	bfr new_net_9964_bfr_after (
		.din(new_net_9963),
		.dout(new_net_9964)
	);

	bfr new_net_9965_bfr_after (
		.din(new_net_9964),
		.dout(new_net_9965)
	);

	bfr new_net_9966_bfr_after (
		.din(new_net_9965),
		.dout(new_net_9966)
	);

	bfr new_net_9967_bfr_after (
		.din(new_net_9966),
		.dout(new_net_9967)
	);

	bfr new_net_9968_bfr_after (
		.din(new_net_9967),
		.dout(new_net_9968)
	);

	bfr new_net_9969_bfr_after (
		.din(new_net_9968),
		.dout(new_net_9969)
	);

	bfr new_net_2444_bfr_after (
		.din(new_net_9969),
		.dout(new_net_2444)
	);

	bfr new_net_9970_bfr_after (
		.din(new_net_2560),
		.dout(new_net_9970)
	);

	bfr new_net_9971_bfr_after (
		.din(new_net_9970),
		.dout(new_net_9971)
	);

	bfr new_net_9972_bfr_after (
		.din(new_net_9971),
		.dout(new_net_9972)
	);

	bfr new_net_9973_bfr_after (
		.din(new_net_9972),
		.dout(new_net_9973)
	);

	bfr new_net_9974_bfr_after (
		.din(new_net_9973),
		.dout(new_net_9974)
	);

	bfr new_net_9975_bfr_after (
		.din(new_net_9974),
		.dout(new_net_9975)
	);

	bfr new_net_9976_bfr_after (
		.din(new_net_9975),
		.dout(new_net_9976)
	);

	bfr new_net_9977_bfr_after (
		.din(new_net_9976),
		.dout(new_net_9977)
	);

	bfr new_net_9978_bfr_after (
		.din(new_net_9977),
		.dout(new_net_9978)
	);

	bfr new_net_9979_bfr_after (
		.din(new_net_9978),
		.dout(new_net_9979)
	);

	bfr new_net_9980_bfr_after (
		.din(new_net_9979),
		.dout(new_net_9980)
	);

	bfr new_net_9981_bfr_after (
		.din(new_net_9980),
		.dout(new_net_9981)
	);

	bfr new_net_9982_bfr_after (
		.din(new_net_9981),
		.dout(new_net_9982)
	);

	bfr new_net_9983_bfr_after (
		.din(new_net_9982),
		.dout(new_net_9983)
	);

	bfr new_net_9984_bfr_after (
		.din(new_net_9983),
		.dout(new_net_9984)
	);

	bfr new_net_9985_bfr_after (
		.din(new_net_9984),
		.dout(new_net_9985)
	);

	bfr new_net_9986_bfr_after (
		.din(new_net_9985),
		.dout(new_net_9986)
	);

	bfr new_net_9987_bfr_after (
		.din(new_net_9986),
		.dout(new_net_9987)
	);

	bfr new_net_9988_bfr_after (
		.din(new_net_9987),
		.dout(new_net_9988)
	);

	bfr new_net_9989_bfr_after (
		.din(new_net_9988),
		.dout(new_net_9989)
	);

	bfr new_net_9990_bfr_after (
		.din(new_net_9989),
		.dout(new_net_9990)
	);

	bfr new_net_9991_bfr_after (
		.din(new_net_9990),
		.dout(new_net_9991)
	);

	bfr new_net_9992_bfr_after (
		.din(new_net_9991),
		.dout(new_net_9992)
	);

	bfr new_net_9993_bfr_after (
		.din(new_net_9992),
		.dout(new_net_9993)
	);

	bfr new_net_9994_bfr_after (
		.din(new_net_9993),
		.dout(new_net_9994)
	);

	bfr new_net_9995_bfr_after (
		.din(new_net_9994),
		.dout(new_net_9995)
	);

	bfr new_net_9996_bfr_after (
		.din(new_net_9995),
		.dout(new_net_9996)
	);

	bfr new_net_9997_bfr_after (
		.din(new_net_9996),
		.dout(new_net_9997)
	);

	bfr new_net_9998_bfr_after (
		.din(new_net_9997),
		.dout(new_net_9998)
	);

	bfr new_net_9999_bfr_after (
		.din(new_net_9998),
		.dout(new_net_9999)
	);

	bfr new_net_10000_bfr_after (
		.din(new_net_9999),
		.dout(new_net_10000)
	);

	bfr new_net_10001_bfr_after (
		.din(new_net_10000),
		.dout(new_net_10001)
	);

	bfr new_net_10002_bfr_after (
		.din(new_net_10001),
		.dout(new_net_10002)
	);

	bfr new_net_10003_bfr_after (
		.din(new_net_10002),
		.dout(new_net_10003)
	);

	bfr new_net_10004_bfr_after (
		.din(new_net_10003),
		.dout(new_net_10004)
	);

	bfr new_net_10005_bfr_after (
		.din(new_net_10004),
		.dout(new_net_10005)
	);

	bfr new_net_10006_bfr_after (
		.din(new_net_10005),
		.dout(new_net_10006)
	);

	bfr new_net_10007_bfr_after (
		.din(new_net_10006),
		.dout(new_net_10007)
	);

	bfr new_net_10008_bfr_after (
		.din(new_net_10007),
		.dout(new_net_10008)
	);

	bfr new_net_10009_bfr_after (
		.din(new_net_10008),
		.dout(new_net_10009)
	);

	bfr new_net_10010_bfr_after (
		.din(new_net_10009),
		.dout(new_net_10010)
	);

	bfr N10729_bfr_after (
		.din(new_net_10010),
		.dout(N10729)
	);

	bfr new_net_10011_bfr_after (
		.din(n_0101_),
		.dout(new_net_10011)
	);

	bfr new_net_10012_bfr_after (
		.din(new_net_10011),
		.dout(new_net_10012)
	);

	bfr new_net_10013_bfr_after (
		.din(new_net_10012),
		.dout(new_net_10013)
	);

	bfr new_net_2388_bfr_after (
		.din(new_net_10013),
		.dout(new_net_2388)
	);

	bfr new_net_2383_bfr_after (
		.din(n_0021_),
		.dout(new_net_2383)
	);

	bfr new_net_10014_bfr_after (
		.din(new_net_2535),
		.dout(new_net_10014)
	);

	bfr new_net_10015_bfr_after (
		.din(new_net_10014),
		.dout(new_net_10015)
	);

	bfr new_net_10016_bfr_after (
		.din(new_net_10015),
		.dout(new_net_10016)
	);

	bfr new_net_10017_bfr_after (
		.din(new_net_10016),
		.dout(new_net_10017)
	);

	bfr new_net_10018_bfr_after (
		.din(new_net_10017),
		.dout(new_net_10018)
	);

	bfr new_net_10019_bfr_after (
		.din(new_net_10018),
		.dout(new_net_10019)
	);

	bfr new_net_10020_bfr_after (
		.din(new_net_10019),
		.dout(new_net_10020)
	);

	bfr new_net_10021_bfr_after (
		.din(new_net_10020),
		.dout(new_net_10021)
	);

	bfr new_net_10022_bfr_after (
		.din(new_net_10021),
		.dout(new_net_10022)
	);

	bfr new_net_10023_bfr_after (
		.din(new_net_10022),
		.dout(new_net_10023)
	);

	bfr new_net_10024_bfr_after (
		.din(new_net_10023),
		.dout(new_net_10024)
	);

	bfr new_net_10025_bfr_after (
		.din(new_net_10024),
		.dout(new_net_10025)
	);

	bfr new_net_10026_bfr_after (
		.din(new_net_10025),
		.dout(new_net_10026)
	);

	bfr new_net_10027_bfr_after (
		.din(new_net_10026),
		.dout(new_net_10027)
	);

	bfr new_net_10028_bfr_after (
		.din(new_net_10027),
		.dout(new_net_10028)
	);

	bfr new_net_10029_bfr_after (
		.din(new_net_10028),
		.dout(new_net_10029)
	);

	bfr new_net_10030_bfr_after (
		.din(new_net_10029),
		.dout(new_net_10030)
	);

	bfr new_net_10031_bfr_after (
		.din(new_net_10030),
		.dout(new_net_10031)
	);

	bfr new_net_10032_bfr_after (
		.din(new_net_10031),
		.dout(new_net_10032)
	);

	bfr new_net_10033_bfr_after (
		.din(new_net_10032),
		.dout(new_net_10033)
	);

	bfr new_net_10034_bfr_after (
		.din(new_net_10033),
		.dout(new_net_10034)
	);

	bfr new_net_10035_bfr_after (
		.din(new_net_10034),
		.dout(new_net_10035)
	);

	bfr new_net_10036_bfr_after (
		.din(new_net_10035),
		.dout(new_net_10036)
	);

	bfr new_net_10037_bfr_after (
		.din(new_net_10036),
		.dout(new_net_10037)
	);

	bfr new_net_10038_bfr_after (
		.din(new_net_10037),
		.dout(new_net_10038)
	);

	bfr new_net_10039_bfr_after (
		.din(new_net_10038),
		.dout(new_net_10039)
	);

	bfr new_net_10040_bfr_after (
		.din(new_net_10039),
		.dout(new_net_10040)
	);

	bfr new_net_10041_bfr_after (
		.din(new_net_10040),
		.dout(new_net_10041)
	);

	bfr new_net_10042_bfr_after (
		.din(new_net_10041),
		.dout(new_net_10042)
	);

	bfr new_net_10043_bfr_after (
		.din(new_net_10042),
		.dout(new_net_10043)
	);

	bfr new_net_10044_bfr_after (
		.din(new_net_10043),
		.dout(new_net_10044)
	);

	bfr new_net_10045_bfr_after (
		.din(new_net_10044),
		.dout(new_net_10045)
	);

	bfr N10352_bfr_after (
		.din(new_net_10045),
		.dout(N10352)
	);

	bfr new_net_10046_bfr_after (
		.din(new_net_2566),
		.dout(new_net_10046)
	);

	bfr new_net_10047_bfr_after (
		.din(new_net_10046),
		.dout(new_net_10047)
	);

	bfr new_net_10048_bfr_after (
		.din(new_net_10047),
		.dout(new_net_10048)
	);

	bfr new_net_10049_bfr_after (
		.din(new_net_10048),
		.dout(new_net_10049)
	);

	bfr new_net_10050_bfr_after (
		.din(new_net_10049),
		.dout(new_net_10050)
	);

	bfr new_net_10051_bfr_after (
		.din(new_net_10050),
		.dout(new_net_10051)
	);

	bfr new_net_10052_bfr_after (
		.din(new_net_10051),
		.dout(new_net_10052)
	);

	bfr new_net_10053_bfr_after (
		.din(new_net_10052),
		.dout(new_net_10053)
	);

	bfr new_net_10054_bfr_after (
		.din(new_net_10053),
		.dout(new_net_10054)
	);

	bfr new_net_10055_bfr_after (
		.din(new_net_10054),
		.dout(new_net_10055)
	);

	bfr new_net_10056_bfr_after (
		.din(new_net_10055),
		.dout(new_net_10056)
	);

	bfr new_net_10057_bfr_after (
		.din(new_net_10056),
		.dout(new_net_10057)
	);

	bfr new_net_10058_bfr_after (
		.din(new_net_10057),
		.dout(new_net_10058)
	);

	bfr N10762_bfr_after (
		.din(new_net_10058),
		.dout(N10762)
	);

	bfr new_net_10059_bfr_after (
		.din(N227),
		.dout(new_net_10059)
	);

	bfr new_net_10060_bfr_after (
		.din(new_net_10059),
		.dout(new_net_10060)
	);

	bfr new_net_10061_bfr_after (
		.din(new_net_10060),
		.dout(new_net_10061)
	);

	bfr new_net_2258_bfr_after (
		.din(new_net_10061),
		.dout(new_net_2258)
	);

	bfr new_net_10062_bfr_after (
		.din(n_0581_),
		.dout(new_net_10062)
	);

	bfr new_net_10063_bfr_after (
		.din(new_net_10062),
		.dout(new_net_10063)
	);

	bfr new_net_10064_bfr_after (
		.din(new_net_10063),
		.dout(new_net_10064)
	);

	bfr new_net_2474_bfr_after (
		.din(new_net_10064),
		.dout(new_net_2474)
	);

	bfr new_net_2368_bfr_after (
		.din(n_1261_),
		.dout(new_net_2368)
	);

	bfr new_net_10065_bfr_after (
		.din(n_0290_),
		.dout(new_net_10065)
	);

	bfr new_net_10066_bfr_after (
		.din(new_net_10065),
		.dout(new_net_10066)
	);

	bfr new_net_10067_bfr_after (
		.din(new_net_10066),
		.dout(new_net_10067)
	);

	bfr new_net_10068_bfr_after (
		.din(new_net_10067),
		.dout(new_net_10068)
	);

	bfr new_net_10069_bfr_after (
		.din(new_net_10068),
		.dout(new_net_10069)
	);

	bfr new_net_10070_bfr_after (
		.din(new_net_10069),
		.dout(new_net_10070)
	);

	bfr new_net_2431_bfr_after (
		.din(new_net_10070),
		.dout(new_net_2431)
	);

	bfr new_net_2452_bfr_after (
		.din(n_0417_),
		.dout(new_net_2452)
	);

	bfr new_net_2473_bfr_after (
		.din(n_0573_),
		.dout(new_net_2473)
	);

	bfr new_net_10071_bfr_after (
		.din(N85),
		.dout(new_net_10071)
	);

	bfr new_net_10072_bfr_after (
		.din(new_net_10071),
		.dout(new_net_10072)
	);

	bfr new_net_10073_bfr_after (
		.din(new_net_10072),
		.dout(new_net_10073)
	);

	bfr new_net_2305_bfr_after (
		.din(new_net_10073),
		.dout(new_net_2305)
	);

	bfr new_net_10074_bfr_after (
		.din(n_0136_),
		.dout(new_net_10074)
	);

	bfr new_net_10075_bfr_after (
		.din(new_net_10074),
		.dout(new_net_10075)
	);

	bfr new_net_10076_bfr_after (
		.din(new_net_10075),
		.dout(new_net_10076)
	);

	bfr new_net_10077_bfr_after (
		.din(new_net_10076),
		.dout(new_net_10077)
	);

	bfr new_net_10078_bfr_after (
		.din(new_net_10077),
		.dout(new_net_10078)
	);

	bfr new_net_10079_bfr_after (
		.din(new_net_10078),
		.dout(new_net_10079)
	);

	bfr new_net_10080_bfr_after (
		.din(new_net_10079),
		.dout(new_net_10080)
	);

	bfr new_net_10081_bfr_after (
		.din(new_net_10080),
		.dout(new_net_10081)
	);

	bfr new_net_10082_bfr_after (
		.din(new_net_10081),
		.dout(new_net_10082)
	);

	bfr new_net_10083_bfr_after (
		.din(new_net_10082),
		.dout(new_net_10083)
	);

	bfr new_net_10084_bfr_after (
		.din(new_net_10083),
		.dout(new_net_10084)
	);

	bfr new_net_10085_bfr_after (
		.din(new_net_10084),
		.dout(new_net_10085)
	);

	bfr new_net_10086_bfr_after (
		.din(new_net_10085),
		.dout(new_net_10086)
	);

	bfr new_net_10087_bfr_after (
		.din(new_net_10086),
		.dout(new_net_10087)
	);

	bfr new_net_10088_bfr_after (
		.din(new_net_10087),
		.dout(new_net_10088)
	);

	bfr new_net_10089_bfr_after (
		.din(new_net_10088),
		.dout(new_net_10089)
	);

	bfr new_net_2389_bfr_after (
		.din(new_net_10089),
		.dout(new_net_2389)
	);

	bfr new_net_10090_bfr_after (
		.din(n_0236_),
		.dout(new_net_10090)
	);

	bfr new_net_2410_bfr_after (
		.din(new_net_10090),
		.dout(new_net_2410)
	);

	bfr new_net_2326_bfr_after (
		.din(n_1157_),
		.dout(new_net_2326)
	);

	bfr new_net_10091_bfr_after (
		.din(N173),
		.dout(new_net_10091)
	);

	bfr new_net_10092_bfr_after (
		.din(new_net_10091),
		.dout(new_net_10092)
	);

	bfr new_net_10093_bfr_after (
		.din(new_net_10092),
		.dout(new_net_10093)
	);

	bfr new_net_2347_bfr_after (
		.din(new_net_10093),
		.dout(new_net_2347)
	);

	bfr new_net_10094_bfr_after (
		.din(N209),
		.dout(new_net_10094)
	);

	bfr new_net_10095_bfr_after (
		.din(new_net_10094),
		.dout(new_net_10095)
	);

	bfr new_net_10096_bfr_after (
		.din(new_net_10095),
		.dout(new_net_10096)
	);

	bfr new_net_2221_bfr_after (
		.din(new_net_10096),
		.dout(new_net_2221)
	);

	bfr new_net_2418_bfr_after (
		.din(n_0259_),
		.dout(new_net_2418)
	);

	bfr new_net_10097_bfr_after (
		.din(n_0241_),
		.dout(new_net_10097)
	);

	bfr new_net_10098_bfr_after (
		.din(new_net_10097),
		.dout(new_net_10098)
	);

	bfr new_net_2413_bfr_after (
		.din(new_net_10098),
		.dout(new_net_2413)
	);

	bfr new_net_10099_bfr_after (
		.din(N236),
		.dout(new_net_10099)
	);

	bfr new_net_10100_bfr_after (
		.din(new_net_10099),
		.dout(new_net_10100)
	);

	bfr new_net_10101_bfr_after (
		.din(new_net_10100),
		.dout(new_net_10101)
	);

	bfr new_net_2191_bfr_after (
		.din(new_net_10101),
		.dout(new_net_2191)
	);

	bfr new_net_2356_bfr_after (
		.din(n_1234_),
		.dout(new_net_2356)
	);

	bfr new_net_10102_bfr_after (
		.din(N55),
		.dout(new_net_10102)
	);

	bfr new_net_10103_bfr_after (
		.din(new_net_10102),
		.dout(new_net_10103)
	);

	bfr new_net_10104_bfr_after (
		.din(new_net_10103),
		.dout(new_net_10104)
	);

	bfr new_net_2288_bfr_after (
		.din(new_net_10104),
		.dout(new_net_2288)
	);

	bfr new_net_2351_bfr_after (
		.din(n_1225_),
		.dout(new_net_2351)
	);

	bfr new_net_10105_bfr_after (
		.din(N88),
		.dout(new_net_10105)
	);

	bfr new_net_10106_bfr_after (
		.din(new_net_10105),
		.dout(new_net_10106)
	);

	bfr new_net_10107_bfr_after (
		.din(new_net_10106),
		.dout(new_net_10107)
	);

	bfr new_net_2279_bfr_after (
		.din(new_net_10107),
		.dout(new_net_2279)
	);

	bfr new_net_10108_bfr_after (
		.din(N181),
		.dout(new_net_10108)
	);

	bfr new_net_10109_bfr_after (
		.din(new_net_10108),
		.dout(new_net_10109)
	);

	bfr new_net_10110_bfr_after (
		.din(new_net_10109),
		.dout(new_net_10110)
	);

	bfr new_net_2342_bfr_after (
		.din(new_net_10110),
		.dout(new_net_2342)
	);

	bfr new_net_10111_bfr_after (
		.din(n_0282_),
		.dout(new_net_10111)
	);

	bfr new_net_10112_bfr_after (
		.din(new_net_10111),
		.dout(new_net_10112)
	);

	bfr new_net_10113_bfr_after (
		.din(new_net_10112),
		.dout(new_net_10113)
	);

	bfr new_net_2426_bfr_after (
		.din(new_net_10113),
		.dout(new_net_2426)
	);

	bfr new_net_10114_bfr_after (
		.din(n_0340_),
		.dout(new_net_10114)
	);

	bfr new_net_2447_bfr_after (
		.din(new_net_10114),
		.dout(new_net_2447)
	);

	bfr new_net_10115_bfr_after (
		.din(N206),
		.dout(new_net_10115)
	);

	bfr new_net_10116_bfr_after (
		.din(new_net_10115),
		.dout(new_net_10116)
	);

	bfr new_net_10117_bfr_after (
		.din(new_net_10116),
		.dout(new_net_10117)
	);

	bfr new_net_2363_bfr_after (
		.din(new_net_10117),
		.dout(new_net_2363)
	);

	bfr new_net_10118_bfr_after (
		.din(N59),
		.dout(new_net_10118)
	);

	bfr new_net_10119_bfr_after (
		.din(new_net_10118),
		.dout(new_net_10119)
	);

	bfr new_net_10120_bfr_after (
		.din(new_net_10119),
		.dout(new_net_10120)
	);

	bfr new_net_2300_bfr_after (
		.din(new_net_10120),
		.dout(new_net_2300)
	);

	bfr new_net_10121_bfr_after (
		.din(n_0042_),
		.dout(new_net_10121)
	);

	bfr new_net_10122_bfr_after (
		.din(new_net_10121),
		.dout(new_net_10122)
	);

	bfr new_net_2384_bfr_after (
		.din(new_net_10122),
		.dout(new_net_2384)
	);

	bfr new_net_10123_bfr_after (
		.din(n_0544_),
		.dout(new_net_10123)
	);

	bfr new_net_10124_bfr_after (
		.din(new_net_10123),
		.dout(new_net_10124)
	);

	bfr new_net_10125_bfr_after (
		.din(new_net_10124),
		.dout(new_net_10125)
	);

	bfr new_net_10126_bfr_after (
		.din(new_net_10125),
		.dout(new_net_10126)
	);

	bfr new_net_10127_bfr_after (
		.din(new_net_10126),
		.dout(new_net_10127)
	);

	bfr new_net_10128_bfr_after (
		.din(new_net_10127),
		.dout(new_net_10128)
	);

	bfr new_net_10129_bfr_after (
		.din(new_net_10128),
		.dout(new_net_10129)
	);

	bfr new_net_10130_bfr_after (
		.din(new_net_10129),
		.dout(new_net_10130)
	);

	bfr new_net_10131_bfr_after (
		.din(new_net_10130),
		.dout(new_net_10131)
	);

	bfr new_net_10132_bfr_after (
		.din(new_net_10131),
		.dout(new_net_10132)
	);

	bfr new_net_10133_bfr_after (
		.din(new_net_10132),
		.dout(new_net_10133)
	);

	bfr new_net_10134_bfr_after (
		.din(new_net_10133),
		.dout(new_net_10134)
	);

	bfr new_net_10135_bfr_after (
		.din(new_net_10134),
		.dout(new_net_10135)
	);

	bfr new_net_2468_bfr_after (
		.din(new_net_10135),
		.dout(new_net_2468)
	);

	bfr new_net_10136_bfr_after (
		.din(N196),
		.dout(new_net_10136)
	);

	bfr new_net_10137_bfr_after (
		.din(new_net_10136),
		.dout(new_net_10137)
	);

	bfr new_net_10138_bfr_after (
		.din(new_net_10137),
		.dout(new_net_10138)
	);

	bfr new_net_2321_bfr_after (
		.din(new_net_10138),
		.dout(new_net_2321)
	);

	bfr new_net_2405_bfr_after (
		.din(n_0218_),
		.dout(new_net_2405)
	);

	bfr new_net_2200_bfr_after (
		.din(n_0698_),
		.dout(new_net_2200)
	);

	bfr new_net_10139_bfr_after (
		.din(N133),
		.dout(new_net_10139)
	);

	bfr new_net_2186_bfr_after (
		.din(new_net_10139),
		.dout(new_net_2186)
	);

	bfr new_net_10140_bfr_after (
		.din(new_net_2572),
		.dout(new_net_10140)
	);

	bfr new_net_10141_bfr_after (
		.din(new_net_10140),
		.dout(new_net_10141)
	);

	bfr new_net_10142_bfr_after (
		.din(new_net_10141),
		.dout(new_net_10142)
	);

	bfr new_net_10143_bfr_after (
		.din(new_net_10142),
		.dout(new_net_10143)
	);

	bfr new_net_10144_bfr_after (
		.din(new_net_10143),
		.dout(new_net_10144)
	);

	bfr N10718_bfr_after (
		.din(new_net_10144),
		.dout(N10718)
	);

	bfr new_net_10145_bfr_after (
		.din(N241_I),
		.dout(new_net_10145)
	);

	bfr new_net_10146_bfr_after (
		.din(new_net_10145),
		.dout(new_net_10146)
	);

	bfr new_net_10147_bfr_after (
		.din(new_net_10146),
		.dout(new_net_10147)
	);

	bfr new_net_10148_bfr_after (
		.din(new_net_10147),
		.dout(new_net_10148)
	);

	bfr new_net_10149_bfr_after (
		.din(new_net_10148),
		.dout(new_net_10149)
	);

	bfr new_net_10150_bfr_after (
		.din(new_net_10149),
		.dout(new_net_10150)
	);

	bfr new_net_10151_bfr_after (
		.din(new_net_10150),
		.dout(new_net_10151)
	);

	bfr new_net_10152_bfr_after (
		.din(new_net_10151),
		.dout(new_net_10152)
	);

	bfr new_net_10153_bfr_after (
		.din(new_net_10152),
		.dout(new_net_10153)
	);

	bfr new_net_10154_bfr_after (
		.din(new_net_10153),
		.dout(new_net_10154)
	);

	bfr new_net_10155_bfr_after (
		.din(new_net_10154),
		.dout(new_net_10155)
	);

	bfr new_net_10156_bfr_after (
		.din(new_net_10155),
		.dout(new_net_10156)
	);

	bfr new_net_10157_bfr_after (
		.din(new_net_10156),
		.dout(new_net_10157)
	);

	bfr new_net_10158_bfr_after (
		.din(new_net_10157),
		.dout(new_net_10158)
	);

	bfr new_net_10159_bfr_after (
		.din(new_net_10158),
		.dout(new_net_10159)
	);

	bfr new_net_10160_bfr_after (
		.din(new_net_10159),
		.dout(new_net_10160)
	);

	bfr new_net_10161_bfr_after (
		.din(new_net_10160),
		.dout(new_net_10161)
	);

	bfr new_net_10162_bfr_after (
		.din(new_net_10161),
		.dout(new_net_10162)
	);

	bfr new_net_10163_bfr_after (
		.din(new_net_10162),
		.dout(new_net_10163)
	);

	bfr new_net_10164_bfr_after (
		.din(new_net_10163),
		.dout(new_net_10164)
	);

	bfr new_net_10165_bfr_after (
		.din(new_net_10164),
		.dout(new_net_10165)
	);

	bfr new_net_10166_bfr_after (
		.din(new_net_10165),
		.dout(new_net_10166)
	);

	bfr new_net_10167_bfr_after (
		.din(new_net_10166),
		.dout(new_net_10167)
	);

	bfr new_net_10168_bfr_after (
		.din(new_net_10167),
		.dout(new_net_10168)
	);

	bfr new_net_10169_bfr_after (
		.din(new_net_10168),
		.dout(new_net_10169)
	);

	bfr new_net_10170_bfr_after (
		.din(new_net_10169),
		.dout(new_net_10170)
	);

	bfr new_net_10171_bfr_after (
		.din(new_net_10170),
		.dout(new_net_10171)
	);

	bfr new_net_10172_bfr_after (
		.din(new_net_10171),
		.dout(new_net_10172)
	);

	bfr new_net_10173_bfr_after (
		.din(new_net_10172),
		.dout(new_net_10173)
	);

	bfr new_net_10174_bfr_after (
		.din(new_net_10173),
		.dout(new_net_10174)
	);

	bfr new_net_10175_bfr_after (
		.din(new_net_10174),
		.dout(new_net_10175)
	);

	bfr new_net_10176_bfr_after (
		.din(new_net_10175),
		.dout(new_net_10176)
	);

	bfr new_net_10177_bfr_after (
		.din(new_net_10176),
		.dout(new_net_10177)
	);

	bfr new_net_10178_bfr_after (
		.din(new_net_10177),
		.dout(new_net_10178)
	);

	bfr new_net_10179_bfr_after (
		.din(new_net_10178),
		.dout(new_net_10179)
	);

	bfr new_net_10180_bfr_after (
		.din(new_net_10179),
		.dout(new_net_10180)
	);

	bfr new_net_10181_bfr_after (
		.din(new_net_10180),
		.dout(new_net_10181)
	);

	bfr new_net_10182_bfr_after (
		.din(new_net_10181),
		.dout(new_net_10182)
	);

	bfr new_net_10183_bfr_after (
		.din(new_net_10182),
		.dout(new_net_10183)
	);

	bfr new_net_10184_bfr_after (
		.din(new_net_10183),
		.dout(new_net_10184)
	);

	bfr new_net_10185_bfr_after (
		.din(new_net_10184),
		.dout(new_net_10185)
	);

	bfr new_net_10186_bfr_after (
		.din(new_net_10185),
		.dout(new_net_10186)
	);

	bfr new_net_10187_bfr_after (
		.din(new_net_10186),
		.dout(new_net_10187)
	);

	bfr new_net_10188_bfr_after (
		.din(new_net_10187),
		.dout(new_net_10188)
	);

	bfr new_net_10189_bfr_after (
		.din(new_net_10188),
		.dout(new_net_10189)
	);

	bfr new_net_10190_bfr_after (
		.din(new_net_10189),
		.dout(new_net_10190)
	);

	bfr new_net_10191_bfr_after (
		.din(new_net_10190),
		.dout(new_net_10191)
	);

	bfr new_net_10192_bfr_after (
		.din(new_net_10191),
		.dout(new_net_10192)
	);

	bfr new_net_10193_bfr_after (
		.din(new_net_10192),
		.dout(new_net_10193)
	);

	bfr new_net_10194_bfr_after (
		.din(new_net_10193),
		.dout(new_net_10194)
	);

	bfr new_net_10195_bfr_after (
		.din(new_net_10194),
		.dout(new_net_10195)
	);

	bfr new_net_10196_bfr_after (
		.din(new_net_10195),
		.dout(new_net_10196)
	);

	bfr new_net_10197_bfr_after (
		.din(new_net_10196),
		.dout(new_net_10197)
	);

	bfr new_net_10198_bfr_after (
		.din(new_net_10197),
		.dout(new_net_10198)
	);

	bfr new_net_10199_bfr_after (
		.din(new_net_10198),
		.dout(new_net_10199)
	);

	bfr new_net_10200_bfr_after (
		.din(new_net_10199),
		.dout(new_net_10200)
	);

	bfr new_net_10201_bfr_after (
		.din(new_net_10200),
		.dout(new_net_10201)
	);

	bfr new_net_10202_bfr_after (
		.din(new_net_10201),
		.dout(new_net_10202)
	);

	bfr new_net_10203_bfr_after (
		.din(new_net_10202),
		.dout(new_net_10203)
	);

	bfr new_net_10204_bfr_after (
		.din(new_net_10203),
		.dout(new_net_10204)
	);

	bfr new_net_10205_bfr_after (
		.din(new_net_10204),
		.dout(new_net_10205)
	);

	bfr new_net_10206_bfr_after (
		.din(new_net_10205),
		.dout(new_net_10206)
	);

	bfr new_net_10207_bfr_after (
		.din(new_net_10206),
		.dout(new_net_10207)
	);

	bfr new_net_10208_bfr_after (
		.din(new_net_10207),
		.dout(new_net_10208)
	);

	bfr new_net_10209_bfr_after (
		.din(new_net_10208),
		.dout(new_net_10209)
	);

	bfr N241_O_bfr_after (
		.din(new_net_10209),
		.dout(N241_O)
	);

	bfr new_net_10210_bfr_after (
		.din(n_0257_),
		.dout(new_net_10210)
	);

	bfr new_net_10211_bfr_after (
		.din(new_net_10210),
		.dout(new_net_10211)
	);

	bfr new_net_10212_bfr_after (
		.din(new_net_10211),
		.dout(new_net_10212)
	);

	bfr new_net_10213_bfr_after (
		.din(new_net_10212),
		.dout(new_net_10213)
	);

	bfr new_net_10214_bfr_after (
		.din(new_net_10213),
		.dout(new_net_10214)
	);

	bfr new_net_2417_bfr_after (
		.din(new_net_10214),
		.dout(new_net_2417)
	);

	bfr new_net_10215_bfr_after (
		.din(new_net_2491),
		.dout(new_net_10215)
	);

	bfr new_net_10216_bfr_after (
		.din(new_net_10215),
		.dout(new_net_10216)
	);

	bfr new_net_10217_bfr_after (
		.din(new_net_10216),
		.dout(new_net_10217)
	);

	bfr new_net_10218_bfr_after (
		.din(new_net_10217),
		.dout(new_net_10218)
	);

	bfr new_net_10219_bfr_after (
		.din(new_net_10218),
		.dout(new_net_10219)
	);

	bfr new_net_10220_bfr_after (
		.din(new_net_10219),
		.dout(new_net_10220)
	);

	bfr new_net_10221_bfr_after (
		.din(new_net_10220),
		.dout(new_net_10221)
	);

	bfr new_net_10222_bfr_after (
		.din(new_net_10221),
		.dout(new_net_10222)
	);

	bfr new_net_10223_bfr_after (
		.din(new_net_10222),
		.dout(new_net_10223)
	);

	bfr new_net_10224_bfr_after (
		.din(new_net_10223),
		.dout(new_net_10224)
	);

	bfr new_net_10225_bfr_after (
		.din(new_net_10224),
		.dout(new_net_10225)
	);

	bfr new_net_10226_bfr_after (
		.din(new_net_10225),
		.dout(new_net_10226)
	);

	bfr new_net_10227_bfr_after (
		.din(new_net_10226),
		.dout(new_net_10227)
	);

	bfr N10760_bfr_after (
		.din(new_net_10227),
		.dout(N10760)
	);

	bfr new_net_10228_bfr_after (
		.din(N124),
		.dout(new_net_10228)
	);

	bfr new_net_10229_bfr_after (
		.din(new_net_10228),
		.dout(new_net_10229)
	);

	bfr new_net_10230_bfr_after (
		.din(new_net_10229),
		.dout(new_net_10230)
	);

	bfr new_net_2230_bfr_after (
		.din(new_net_10230),
		.dout(new_net_2230)
	);

	bfr new_net_10231_bfr_after (
		.din(N32),
		.dout(new_net_10231)
	);

	bfr new_net_10232_bfr_after (
		.din(new_net_10231),
		.dout(new_net_10232)
	);

	bfr new_net_10233_bfr_after (
		.din(new_net_10232),
		.dout(new_net_10233)
	);

	bfr new_net_2274_bfr_after (
		.din(new_net_10233),
		.dout(new_net_2274)
	);

	bfr new_net_10234_bfr_after (
		.din(N197),
		.dout(new_net_10234)
	);

	bfr new_net_10235_bfr_after (
		.din(new_net_10234),
		.dout(new_net_10235)
	);

	bfr new_net_10236_bfr_after (
		.din(new_net_10235),
		.dout(new_net_10236)
	);

	bfr new_net_2337_bfr_after (
		.din(new_net_10236),
		.dout(new_net_2337)
	);

	bfr new_net_2421_bfr_after (
		.din(n_0265_),
		.dout(new_net_2421)
	);

	bfr new_net_10237_bfr_after (
		.din(n_0325_),
		.dout(new_net_10237)
	);

	bfr new_net_10238_bfr_after (
		.din(new_net_10237),
		.dout(new_net_10238)
	);

	bfr new_net_2442_bfr_after (
		.din(new_net_10238),
		.dout(new_net_2442)
	);

	bfr new_net_10239_bfr_after (
		.din(N135),
		.dout(new_net_10239)
	);

	bfr new_net_10240_bfr_after (
		.din(new_net_10239),
		.dout(new_net_10240)
	);

	bfr new_net_10241_bfr_after (
		.din(new_net_10240),
		.dout(new_net_10241)
	);

	bfr new_net_2211_bfr_after (
		.din(new_net_10241),
		.dout(new_net_2211)
	);

	bfr new_net_10242_bfr_after (
		.din(N229),
		.dout(new_net_10242)
	);

	bfr new_net_10243_bfr_after (
		.din(new_net_10242),
		.dout(new_net_10243)
	);

	bfr new_net_10244_bfr_after (
		.din(new_net_10243),
		.dout(new_net_10244)
	);

	bfr new_net_2232_bfr_after (
		.din(new_net_10244),
		.dout(new_net_2232)
	);

	bfr new_net_10245_bfr_after (
		.din(N97),
		.dout(new_net_10245)
	);

	bfr new_net_10246_bfr_after (
		.din(new_net_10245),
		.dout(new_net_10246)
	);

	bfr new_net_10247_bfr_after (
		.din(new_net_10246),
		.dout(new_net_10247)
	);

	bfr new_net_2253_bfr_after (
		.din(new_net_10247),
		.dout(new_net_2253)
	);

	bfr new_net_2358_bfr_after (
		.din(n_1245_),
		.dout(new_net_2358)
	);

	bfr new_net_10248_bfr_after (
		.din(N81),
		.dout(new_net_10248)
	);

	bfr new_net_10249_bfr_after (
		.din(new_net_10248),
		.dout(new_net_10249)
	);

	bfr new_net_10250_bfr_after (
		.din(new_net_10249),
		.dout(new_net_10250)
	);

	bfr new_net_2295_bfr_after (
		.din(new_net_10250),
		.dout(new_net_2295)
	);

	bfr new_net_10251_bfr_after (
		.din(n_1363_),
		.dout(new_net_10251)
	);

	bfr new_net_2379_bfr_after (
		.din(new_net_10251),
		.dout(new_net_2379)
	);

	bfr new_net_10252_bfr_after (
		.din(n_0570_),
		.dout(new_net_10252)
	);

	bfr new_net_2472_bfr_after (
		.din(new_net_10252),
		.dout(new_net_2472)
	);

	bfr new_net_2190_bfr_after (
		.din(n_0671_),
		.dout(new_net_2190)
	);

	bfr new_net_2269_bfr_after (
		.din(n_0879_),
		.dout(new_net_2269)
	);

	bfr new_net_10253_bfr_after (
		.din(N84),
		.dout(new_net_10253)
	);

	bfr new_net_10254_bfr_after (
		.din(new_net_10253),
		.dout(new_net_10254)
	);

	bfr new_net_10255_bfr_after (
		.din(new_net_10254),
		.dout(new_net_10255)
	);

	bfr new_net_2311_bfr_after (
		.din(new_net_10255),
		.dout(new_net_2311)
	);

	bfr new_net_2395_bfr_after (
		.din(n_0179_),
		.dout(new_net_2395)
	);

	bfr new_net_2416_bfr_after (
		.din(n_0256_),
		.dout(new_net_2416)
	);

	bfr new_net_10256_bfr_after (
		.din(N161),
		.dout(new_net_10256)
	);

	bfr new_net_10257_bfr_after (
		.din(new_net_10256),
		.dout(new_net_10257)
	);

	bfr new_net_10258_bfr_after (
		.din(new_net_10257),
		.dout(new_net_10258)
	);

	bfr new_net_2206_bfr_after (
		.din(new_net_10258),
		.dout(new_net_2206)
	);

	bfr new_net_10259_bfr_after (
		.din(n_0798_),
		.dout(new_net_10259)
	);

	bfr new_net_2227_bfr_after (
		.din(new_net_10259),
		.dout(new_net_2227)
	);

	bfr new_net_2248_bfr_after (
		.din(n_0846_),
		.dout(new_net_2248)
	);

	bfr new_net_10260_bfr_after (
		.din(N54),
		.dout(new_net_10260)
	);

	bfr new_net_10261_bfr_after (
		.din(new_net_10260),
		.dout(new_net_10261)
	);

	bfr new_net_10262_bfr_after (
		.din(new_net_10261),
		.dout(new_net_10262)
	);

	bfr new_net_2290_bfr_after (
		.din(new_net_10262),
		.dout(new_net_2290)
	);

	bfr new_net_2332_bfr_after (
		.din(n_1166_),
		.dout(new_net_2332)
	);

	bfr new_net_10263_bfr_after (
		.din(N180),
		.dout(new_net_10263)
	);

	bfr new_net_10264_bfr_after (
		.din(new_net_10263),
		.dout(new_net_10264)
	);

	bfr new_net_10265_bfr_after (
		.din(new_net_10264),
		.dout(new_net_10265)
	);

	bfr new_net_2353_bfr_after (
		.din(new_net_10265),
		.dout(new_net_2353)
	);

	bfr new_net_10266_bfr_after (
		.din(N232),
		.dout(new_net_10266)
	);

	bfr new_net_10267_bfr_after (
		.din(new_net_10266),
		.dout(new_net_10267)
	);

	bfr new_net_10268_bfr_after (
		.din(new_net_10267),
		.dout(new_net_10268)
	);

	bfr new_net_2229_bfr_after (
		.din(new_net_10268),
		.dout(new_net_2229)
	);

	bfr new_net_2184_bfr_after (
		.din(N242),
		.dout(new_net_2184)
	);

	bfr new_net_10269_bfr_after (
		.din(n_0562_),
		.dout(new_net_10269)
	);

	bfr new_net_2471_bfr_after (
		.din(new_net_10269),
		.dout(new_net_2471)
	);

	bfr N10101_bfr_after (
		.din(new_net_2489),
		.dout(N10101)
	);

	bfr new_net_10270_bfr_after (
		.din(new_net_2501),
		.dout(new_net_10270)
	);

	bfr new_net_10271_bfr_after (
		.din(new_net_10270),
		.dout(new_net_10271)
	);

	bfr new_net_10272_bfr_after (
		.din(new_net_10271),
		.dout(new_net_10272)
	);

	bfr new_net_10273_bfr_after (
		.din(new_net_10272),
		.dout(new_net_10273)
	);

	bfr new_net_10274_bfr_after (
		.din(new_net_10273),
		.dout(new_net_10274)
	);

	bfr new_net_10275_bfr_after (
		.din(new_net_10274),
		.dout(new_net_10275)
	);

	bfr new_net_10276_bfr_after (
		.din(new_net_10275),
		.dout(new_net_10276)
	);

	bfr new_net_10277_bfr_after (
		.din(new_net_10276),
		.dout(new_net_10277)
	);

	bfr new_net_10278_bfr_after (
		.din(new_net_10277),
		.dout(new_net_10278)
	);

	bfr new_net_10279_bfr_after (
		.din(new_net_10278),
		.dout(new_net_10279)
	);

	bfr new_net_10280_bfr_after (
		.din(new_net_10279),
		.dout(new_net_10280)
	);

	bfr new_net_10281_bfr_after (
		.din(new_net_10280),
		.dout(new_net_10281)
	);

	bfr new_net_10282_bfr_after (
		.din(new_net_10281),
		.dout(new_net_10282)
	);

	bfr new_net_10283_bfr_after (
		.din(new_net_10282),
		.dout(new_net_10283)
	);

	bfr new_net_10284_bfr_after (
		.din(new_net_10283),
		.dout(new_net_10284)
	);

	bfr new_net_10285_bfr_after (
		.din(new_net_10284),
		.dout(new_net_10285)
	);

	bfr new_net_10286_bfr_after (
		.din(new_net_10285),
		.dout(new_net_10286)
	);

	bfr new_net_10287_bfr_after (
		.din(new_net_10286),
		.dout(new_net_10287)
	);

	bfr new_net_10288_bfr_after (
		.din(new_net_10287),
		.dout(new_net_10288)
	);

	bfr new_net_10289_bfr_after (
		.din(new_net_10288),
		.dout(new_net_10289)
	);

	bfr new_net_10290_bfr_after (
		.din(new_net_10289),
		.dout(new_net_10290)
	);

	bfr new_net_10291_bfr_after (
		.din(new_net_10290),
		.dout(new_net_10291)
	);

	bfr new_net_10292_bfr_after (
		.din(new_net_10291),
		.dout(new_net_10292)
	);

	bfr new_net_10293_bfr_after (
		.din(new_net_10292),
		.dout(new_net_10293)
	);

	bfr new_net_10294_bfr_after (
		.din(new_net_10293),
		.dout(new_net_10294)
	);

	bfr new_net_10295_bfr_after (
		.din(new_net_10294),
		.dout(new_net_10295)
	);

	bfr new_net_10296_bfr_after (
		.din(new_net_10295),
		.dout(new_net_10296)
	);

	bfr new_net_10297_bfr_after (
		.din(new_net_10296),
		.dout(new_net_10297)
	);

	bfr new_net_10298_bfr_after (
		.din(new_net_10297),
		.dout(new_net_10298)
	);

	bfr new_net_10299_bfr_after (
		.din(new_net_10298),
		.dout(new_net_10299)
	);

	bfr new_net_10300_bfr_after (
		.din(new_net_10299),
		.dout(new_net_10300)
	);

	bfr new_net_10301_bfr_after (
		.din(new_net_10300),
		.dout(new_net_10301)
	);

	bfr new_net_10302_bfr_after (
		.din(new_net_10301),
		.dout(new_net_10302)
	);

	bfr N10350_bfr_after (
		.din(new_net_10302),
		.dout(N10350)
	);

	bfr new_net_10303_bfr_after (
		.din(new_net_2513),
		.dout(new_net_10303)
	);

	bfr new_net_10304_bfr_after (
		.din(new_net_10303),
		.dout(new_net_10304)
	);

	bfr new_net_10305_bfr_after (
		.din(new_net_10304),
		.dout(new_net_10305)
	);

	bfr new_net_10306_bfr_after (
		.din(new_net_10305),
		.dout(new_net_10306)
	);

	bfr new_net_10307_bfr_after (
		.din(new_net_10306),
		.dout(new_net_10307)
	);

	bfr new_net_10308_bfr_after (
		.din(new_net_10307),
		.dout(new_net_10308)
	);

	bfr new_net_10309_bfr_after (
		.din(new_net_10308),
		.dout(new_net_10309)
	);

	bfr new_net_10310_bfr_after (
		.din(new_net_10309),
		.dout(new_net_10310)
	);

	bfr new_net_10311_bfr_after (
		.din(new_net_10310),
		.dout(new_net_10311)
	);

	bfr new_net_10312_bfr_after (
		.din(new_net_10311),
		.dout(new_net_10312)
	);

	bfr new_net_10313_bfr_after (
		.din(new_net_10312),
		.dout(new_net_10313)
	);

	bfr new_net_10314_bfr_after (
		.din(new_net_10313),
		.dout(new_net_10314)
	);

	bfr new_net_10315_bfr_after (
		.din(new_net_10314),
		.dout(new_net_10315)
	);

	bfr new_net_10316_bfr_after (
		.din(new_net_10315),
		.dout(new_net_10316)
	);

	bfr new_net_10317_bfr_after (
		.din(new_net_10316),
		.dout(new_net_10317)
	);

	bfr new_net_10318_bfr_after (
		.din(new_net_10317),
		.dout(new_net_10318)
	);

	bfr new_net_10319_bfr_after (
		.din(new_net_10318),
		.dout(new_net_10319)
	);

	bfr new_net_10320_bfr_after (
		.din(new_net_10319),
		.dout(new_net_10320)
	);

	bfr new_net_10321_bfr_after (
		.din(new_net_10320),
		.dout(new_net_10321)
	);

	bfr new_net_10322_bfr_after (
		.din(new_net_10321),
		.dout(new_net_10322)
	);

	bfr new_net_10323_bfr_after (
		.din(new_net_10322),
		.dout(new_net_10323)
	);

	bfr new_net_10324_bfr_after (
		.din(new_net_10323),
		.dout(new_net_10324)
	);

	bfr new_net_10325_bfr_after (
		.din(new_net_10324),
		.dout(new_net_10325)
	);

	bfr new_net_10326_bfr_after (
		.din(new_net_10325),
		.dout(new_net_10326)
	);

	bfr new_net_10327_bfr_after (
		.din(new_net_10326),
		.dout(new_net_10327)
	);

	bfr new_net_10328_bfr_after (
		.din(new_net_10327),
		.dout(new_net_10328)
	);

	bfr new_net_10329_bfr_after (
		.din(new_net_10328),
		.dout(new_net_10329)
	);

	bfr new_net_10330_bfr_after (
		.din(new_net_10329),
		.dout(new_net_10330)
	);

	bfr new_net_10331_bfr_after (
		.din(new_net_10330),
		.dout(new_net_10331)
	);

	bfr new_net_10332_bfr_after (
		.din(new_net_10331),
		.dout(new_net_10332)
	);

	bfr new_net_10333_bfr_after (
		.din(new_net_10332),
		.dout(new_net_10333)
	);

	bfr new_net_10334_bfr_after (
		.din(new_net_10333),
		.dout(new_net_10334)
	);

	bfr new_net_10335_bfr_after (
		.din(new_net_10334),
		.dout(new_net_10335)
	);

	bfr new_net_10336_bfr_after (
		.din(new_net_10335),
		.dout(new_net_10336)
	);

	bfr new_net_10337_bfr_after (
		.din(new_net_10336),
		.dout(new_net_10337)
	);

	bfr new_net_10338_bfr_after (
		.din(new_net_10337),
		.dout(new_net_10338)
	);

	bfr new_net_10339_bfr_after (
		.din(new_net_10338),
		.dout(new_net_10339)
	);

	bfr new_net_10340_bfr_after (
		.din(new_net_10339),
		.dout(new_net_10340)
	);

	bfr new_net_10341_bfr_after (
		.din(new_net_10340),
		.dout(new_net_10341)
	);

	bfr new_net_10342_bfr_after (
		.din(new_net_10341),
		.dout(new_net_10342)
	);

	bfr new_net_10343_bfr_after (
		.din(new_net_10342),
		.dout(new_net_10343)
	);

	bfr new_net_10344_bfr_after (
		.din(new_net_10343),
		.dout(new_net_10344)
	);

	bfr new_net_10345_bfr_after (
		.din(new_net_10344),
		.dout(new_net_10345)
	);

	bfr N10110_bfr_after (
		.din(new_net_10345),
		.dout(N10110)
	);

	bfr new_net_10346_bfr_after (
		.din(new_net_2525),
		.dout(new_net_10346)
	);

	bfr new_net_10347_bfr_after (
		.din(new_net_10346),
		.dout(new_net_10347)
	);

	bfr new_net_10348_bfr_after (
		.din(new_net_10347),
		.dout(new_net_10348)
	);

	bfr new_net_10349_bfr_after (
		.din(new_net_10348),
		.dout(new_net_10349)
	);

	bfr new_net_10350_bfr_after (
		.din(new_net_10349),
		.dout(new_net_10350)
	);

	bfr new_net_10351_bfr_after (
		.din(new_net_10350),
		.dout(new_net_10351)
	);

	bfr new_net_10352_bfr_after (
		.din(new_net_10351),
		.dout(new_net_10352)
	);

	bfr new_net_10353_bfr_after (
		.din(new_net_10352),
		.dout(new_net_10353)
	);

	bfr new_net_10354_bfr_after (
		.din(new_net_10353),
		.dout(new_net_10354)
	);

	bfr new_net_10355_bfr_after (
		.din(new_net_10354),
		.dout(new_net_10355)
	);

	bfr new_net_10356_bfr_after (
		.din(new_net_10355),
		.dout(new_net_10356)
	);

	bfr new_net_10357_bfr_after (
		.din(new_net_10356),
		.dout(new_net_10357)
	);

	bfr new_net_10358_bfr_after (
		.din(new_net_10357),
		.dout(new_net_10358)
	);

	bfr new_net_10359_bfr_after (
		.din(new_net_10358),
		.dout(new_net_10359)
	);

	bfr new_net_10360_bfr_after (
		.din(new_net_10359),
		.dout(new_net_10360)
	);

	bfr new_net_10361_bfr_after (
		.din(new_net_10360),
		.dout(new_net_10361)
	);

	bfr new_net_10362_bfr_after (
		.din(new_net_10361),
		.dout(new_net_10362)
	);

	bfr new_net_10363_bfr_after (
		.din(new_net_10362),
		.dout(new_net_10363)
	);

	bfr new_net_10364_bfr_after (
		.din(new_net_10363),
		.dout(new_net_10364)
	);

	bfr new_net_10365_bfr_after (
		.din(new_net_10364),
		.dout(new_net_10365)
	);

	bfr new_net_10366_bfr_after (
		.din(new_net_10365),
		.dout(new_net_10366)
	);

	bfr new_net_10367_bfr_after (
		.din(new_net_10366),
		.dout(new_net_10367)
	);

	bfr new_net_10368_bfr_after (
		.din(new_net_10367),
		.dout(new_net_10368)
	);

	bfr new_net_10369_bfr_after (
		.din(new_net_10368),
		.dout(new_net_10369)
	);

	bfr new_net_10370_bfr_after (
		.din(new_net_10369),
		.dout(new_net_10370)
	);

	bfr new_net_10371_bfr_after (
		.din(new_net_10370),
		.dout(new_net_10371)
	);

	bfr new_net_10372_bfr_after (
		.din(new_net_10371),
		.dout(new_net_10372)
	);

	bfr new_net_10373_bfr_after (
		.din(new_net_10372),
		.dout(new_net_10373)
	);

	bfr new_net_10374_bfr_after (
		.din(new_net_10373),
		.dout(new_net_10374)
	);

	bfr new_net_10375_bfr_after (
		.din(new_net_10374),
		.dout(new_net_10375)
	);

	bfr new_net_10376_bfr_after (
		.din(new_net_10375),
		.dout(new_net_10376)
	);

	bfr N10827_bfr_after (
		.din(new_net_10376),
		.dout(N10827)
	);

	bfr new_net_10377_bfr_after (
		.din(new_net_2537),
		.dout(new_net_10377)
	);

	bfr new_net_10378_bfr_after (
		.din(new_net_10377),
		.dout(new_net_10378)
	);

	bfr new_net_10379_bfr_after (
		.din(new_net_10378),
		.dout(new_net_10379)
	);

	bfr new_net_10380_bfr_after (
		.din(new_net_10379),
		.dout(new_net_10380)
	);

	bfr new_net_10381_bfr_after (
		.din(new_net_10380),
		.dout(new_net_10381)
	);

	bfr new_net_10382_bfr_after (
		.din(new_net_10381),
		.dout(new_net_10382)
	);

	bfr N10717_bfr_after (
		.din(new_net_10382),
		.dout(N10717)
	);

	bfr new_net_10383_bfr_after (
		.din(new_net_2547),
		.dout(new_net_10383)
	);

	bfr new_net_10384_bfr_after (
		.din(new_net_10383),
		.dout(new_net_10384)
	);

	bfr new_net_10385_bfr_after (
		.din(new_net_10384),
		.dout(new_net_10385)
	);

	bfr new_net_10386_bfr_after (
		.din(new_net_10385),
		.dout(new_net_10386)
	);

	bfr new_net_10387_bfr_after (
		.din(new_net_10386),
		.dout(new_net_10387)
	);

	bfr new_net_10388_bfr_after (
		.din(new_net_10387),
		.dout(new_net_10388)
	);

	bfr new_net_10389_bfr_after (
		.din(new_net_10388),
		.dout(new_net_10389)
	);

	bfr new_net_10390_bfr_after (
		.din(new_net_10389),
		.dout(new_net_10390)
	);

	bfr new_net_10391_bfr_after (
		.din(new_net_10390),
		.dout(new_net_10391)
	);

	bfr new_net_10392_bfr_after (
		.din(new_net_10391),
		.dout(new_net_10392)
	);

	bfr new_net_10393_bfr_after (
		.din(new_net_10392),
		.dout(new_net_10393)
	);

	bfr new_net_10394_bfr_after (
		.din(new_net_10393),
		.dout(new_net_10394)
	);

	bfr new_net_10395_bfr_after (
		.din(new_net_10394),
		.dout(new_net_10395)
	);

	bfr new_net_10396_bfr_after (
		.din(new_net_10395),
		.dout(new_net_10396)
	);

	bfr new_net_10397_bfr_after (
		.din(new_net_10396),
		.dout(new_net_10397)
	);

	bfr new_net_10398_bfr_after (
		.din(new_net_10397),
		.dout(new_net_10398)
	);

	bfr new_net_10399_bfr_after (
		.din(new_net_10398),
		.dout(new_net_10399)
	);

	bfr new_net_10400_bfr_after (
		.din(new_net_10399),
		.dout(new_net_10400)
	);

	bfr new_net_10401_bfr_after (
		.din(new_net_10400),
		.dout(new_net_10401)
	);

	bfr new_net_10402_bfr_after (
		.din(new_net_10401),
		.dout(new_net_10402)
	);

	bfr new_net_10403_bfr_after (
		.din(new_net_10402),
		.dout(new_net_10403)
	);

	bfr new_net_10404_bfr_after (
		.din(new_net_10403),
		.dout(new_net_10404)
	);

	bfr new_net_10405_bfr_after (
		.din(new_net_10404),
		.dout(new_net_10405)
	);

	bfr new_net_10406_bfr_after (
		.din(new_net_10405),
		.dout(new_net_10406)
	);

	bfr new_net_10407_bfr_after (
		.din(new_net_10406),
		.dout(new_net_10407)
	);

	bfr new_net_10408_bfr_after (
		.din(new_net_10407),
		.dout(new_net_10408)
	);

	bfr new_net_10409_bfr_after (
		.din(new_net_10408),
		.dout(new_net_10409)
	);

	bfr new_net_10410_bfr_after (
		.din(new_net_10409),
		.dout(new_net_10410)
	);

	bfr N10871_bfr_after (
		.din(new_net_10410),
		.dout(N10871)
	);

	bfr new_net_10411_bfr_after (
		.din(new_net_2549),
		.dout(new_net_10411)
	);

	bfr new_net_10412_bfr_after (
		.din(new_net_10411),
		.dout(new_net_10412)
	);

	bfr new_net_10413_bfr_after (
		.din(new_net_10412),
		.dout(new_net_10413)
	);

	bfr new_net_10414_bfr_after (
		.din(new_net_10413),
		.dout(new_net_10414)
	);

	bfr new_net_10415_bfr_after (
		.din(new_net_10414),
		.dout(new_net_10415)
	);

	bfr new_net_10416_bfr_after (
		.din(new_net_10415),
		.dout(new_net_10416)
	);

	bfr new_net_10417_bfr_after (
		.din(new_net_10416),
		.dout(new_net_10417)
	);

	bfr new_net_10418_bfr_after (
		.din(new_net_10417),
		.dout(new_net_10418)
	);

	bfr new_net_10419_bfr_after (
		.din(new_net_10418),
		.dout(new_net_10419)
	);

	bfr new_net_10420_bfr_after (
		.din(new_net_10419),
		.dout(new_net_10420)
	);

	bfr new_net_10421_bfr_after (
		.din(new_net_10420),
		.dout(new_net_10421)
	);

	bfr new_net_10422_bfr_after (
		.din(new_net_10421),
		.dout(new_net_10422)
	);

	bfr new_net_10423_bfr_after (
		.din(new_net_10422),
		.dout(new_net_10423)
	);

	bfr new_net_10424_bfr_after (
		.din(new_net_10423),
		.dout(new_net_10424)
	);

	bfr new_net_10425_bfr_after (
		.din(new_net_10424),
		.dout(new_net_10425)
	);

	bfr new_net_10426_bfr_after (
		.din(new_net_10425),
		.dout(new_net_10426)
	);

	bfr N10763_bfr_after (
		.din(new_net_10426),
		.dout(N10763)
	);

	bfr new_net_10427_bfr_after (
		.din(N220),
		.dout(new_net_10427)
	);

	bfr new_net_10428_bfr_after (
		.din(new_net_10427),
		.dout(new_net_10428)
	);

	bfr new_net_10429_bfr_after (
		.din(new_net_10428),
		.dout(new_net_10429)
	);

	bfr new_net_2264_bfr_after (
		.din(new_net_10429),
		.dout(new_net_2264)
	);

	bfr new_net_10430_bfr_after (
		.din(N64),
		.dout(new_net_10430)
	);

	bfr new_net_10431_bfr_after (
		.din(new_net_10430),
		.dout(new_net_10431)
	);

	bfr new_net_10432_bfr_after (
		.din(new_net_10431),
		.dout(new_net_10432)
	);

	bfr new_net_2306_bfr_after (
		.din(new_net_10432),
		.dout(new_net_2306)
	);

	bfr new_net_2390_bfr_after (
		.din(n_0141_),
		.dout(new_net_2390)
	);

	bfr new_net_10433_bfr_after (
		.din(n_0237_),
		.dout(new_net_10433)
	);

	bfr new_net_10434_bfr_after (
		.din(new_net_10433),
		.dout(new_net_10434)
	);

	bfr new_net_2411_bfr_after (
		.din(new_net_10434),
		.dout(new_net_2411)
	);

	bfr new_net_10435_bfr_after (
		.din(N69),
		.dout(new_net_10435)
	);

	bfr new_net_10436_bfr_after (
		.din(new_net_10435),
		.dout(new_net_10436)
	);

	bfr new_net_10437_bfr_after (
		.din(new_net_10436),
		.dout(new_net_10437)
	);

	bfr new_net_2285_bfr_after (
		.din(new_net_10437),
		.dout(new_net_2285)
	);

	bfr new_net_10438_bfr_after (
		.din(N189),
		.dout(new_net_10438)
	);

	bfr new_net_10439_bfr_after (
		.din(new_net_10438),
		.dout(new_net_10439)
	);

	bfr new_net_10440_bfr_after (
		.din(new_net_10439),
		.dout(new_net_10440)
	);

	bfr new_net_2327_bfr_after (
		.din(new_net_10440),
		.dout(new_net_2327)
	);

	bfr new_net_10441_bfr_after (
		.din(N176),
		.dout(new_net_10441)
	);

	bfr new_net_10442_bfr_after (
		.din(new_net_10441),
		.dout(new_net_10442)
	);

	bfr new_net_10443_bfr_after (
		.din(new_net_10442),
		.dout(new_net_10443)
	);

	bfr new_net_2348_bfr_after (
		.din(new_net_10443),
		.dout(new_net_2348)
	);

	bfr new_net_10444_bfr_after (
		.din(N214),
		.dout(new_net_10444)
	);

	bfr new_net_10445_bfr_after (
		.din(new_net_10444),
		.dout(new_net_10445)
	);

	bfr new_net_10446_bfr_after (
		.din(new_net_10445),
		.dout(new_net_10446)
	);

	bfr new_net_2222_bfr_after (
		.din(new_net_10446),
		.dout(new_net_2222)
	);

	bfr new_net_10447_bfr_after (
		.din(N239),
		.dout(new_net_10447)
	);

	bfr new_net_10448_bfr_after (
		.din(new_net_10447),
		.dout(new_net_10448)
	);

	bfr new_net_10449_bfr_after (
		.din(new_net_10448),
		.dout(new_net_10449)
	);

	bfr new_net_2243_bfr_after (
		.din(new_net_10449),
		.dout(new_net_2243)
	);

	bfr new_net_10450_bfr_after (
		.din(N154),
		.dout(new_net_10450)
	);

	bfr new_net_10451_bfr_after (
		.din(new_net_10450),
		.dout(new_net_10451)
	);

	bfr new_net_10452_bfr_after (
		.din(new_net_10451),
		.dout(new_net_10452)
	);

	bfr new_net_2201_bfr_after (
		.din(new_net_10452),
		.dout(new_net_2201)
	);

	bfr new_net_10453_bfr_after (
		.din(new_net_2503),
		.dout(new_net_10453)
	);

	bfr new_net_10454_bfr_after (
		.din(new_net_10453),
		.dout(new_net_10454)
	);

	bfr new_net_10455_bfr_after (
		.din(new_net_10454),
		.dout(new_net_10455)
	);

	bfr new_net_10456_bfr_after (
		.din(new_net_10455),
		.dout(new_net_10456)
	);

	bfr new_net_10457_bfr_after (
		.din(new_net_10456),
		.dout(new_net_10457)
	);

	bfr new_net_10458_bfr_after (
		.din(new_net_10457),
		.dout(new_net_10458)
	);

	bfr new_net_10459_bfr_after (
		.din(new_net_10458),
		.dout(new_net_10459)
	);

	bfr new_net_10460_bfr_after (
		.din(new_net_10459),
		.dout(new_net_10460)
	);

	bfr new_net_10461_bfr_after (
		.din(new_net_10460),
		.dout(new_net_10461)
	);

	bfr new_net_10462_bfr_after (
		.din(new_net_10461),
		.dout(new_net_10462)
	);

	bfr new_net_10463_bfr_after (
		.din(new_net_10462),
		.dout(new_net_10463)
	);

	bfr new_net_10464_bfr_after (
		.din(new_net_10463),
		.dout(new_net_10464)
	);

	bfr new_net_10465_bfr_after (
		.din(new_net_10464),
		.dout(new_net_10465)
	);

	bfr new_net_10466_bfr_after (
		.din(new_net_10465),
		.dout(new_net_10466)
	);

	bfr new_net_10467_bfr_after (
		.din(new_net_10466),
		.dout(new_net_10467)
	);

	bfr new_net_10468_bfr_after (
		.din(new_net_10467),
		.dout(new_net_10468)
	);

	bfr new_net_10469_bfr_after (
		.din(new_net_10468),
		.dout(new_net_10469)
	);

	bfr new_net_10470_bfr_after (
		.din(new_net_10469),
		.dout(new_net_10470)
	);

	bfr new_net_10471_bfr_after (
		.din(new_net_10470),
		.dout(new_net_10471)
	);

	bfr new_net_10472_bfr_after (
		.din(new_net_10471),
		.dout(new_net_10472)
	);

	bfr new_net_10473_bfr_after (
		.din(new_net_10472),
		.dout(new_net_10473)
	);

	bfr new_net_10474_bfr_after (
		.din(new_net_10473),
		.dout(new_net_10474)
	);

	bfr new_net_10475_bfr_after (
		.din(new_net_10474),
		.dout(new_net_10475)
	);

	bfr new_net_10476_bfr_after (
		.din(new_net_10475),
		.dout(new_net_10476)
	);

	bfr N10906_bfr_after (
		.din(new_net_10476),
		.dout(N10906)
	);

	bfr new_net_2374_bfr_after (
		.din(n_1279_),
		.dout(new_net_2374)
	);

	bfr new_net_10477_bfr_after (
		.din(n_0310_),
		.dout(new_net_10477)
	);

	bfr new_net_2437_bfr_after (
		.din(new_net_10477),
		.dout(new_net_2437)
	);

	bfr new_net_2364_bfr_after (
		.din(n_1254_),
		.dout(new_net_2364)
	);

	bfr new_net_2469_bfr_after (
		.din(n_0547_),
		.dout(new_net_2469)
	);

	bfr new_net_10478_bfr_after (
		.din(N79),
		.dout(new_net_10478)
	);

	bfr new_net_10479_bfr_after (
		.din(new_net_10478),
		.dout(new_net_10479)
	);

	bfr new_net_10480_bfr_after (
		.din(new_net_10479),
		.dout(new_net_10480)
	);

	bfr new_net_2301_bfr_after (
		.din(new_net_10480),
		.dout(new_net_2301)
	);

	bfr new_net_10481_bfr_after (
		.din(n_0050_),
		.dout(new_net_10481)
	);

	bfr new_net_10482_bfr_after (
		.din(new_net_10481),
		.dout(new_net_10482)
	);

	bfr new_net_10483_bfr_after (
		.din(new_net_10482),
		.dout(new_net_10483)
	);

	bfr new_net_2385_bfr_after (
		.din(new_net_10483),
		.dout(new_net_2385)
	);

	bfr new_net_2322_bfr_after (
		.din(n_1150_),
		.dout(new_net_2322)
	);

	bfr new_net_10484_bfr_after (
		.din(n_0219_),
		.dout(new_net_10484)
	);

	bfr new_net_10485_bfr_after (
		.din(new_net_10484),
		.dout(new_net_10485)
	);

	bfr new_net_10486_bfr_after (
		.din(new_net_10485),
		.dout(new_net_10486)
	);

	bfr new_net_10487_bfr_after (
		.din(new_net_10486),
		.dout(new_net_10487)
	);

	bfr new_net_2406_bfr_after (
		.din(new_net_10487),
		.dout(new_net_2406)
	);

	bfr new_net_10488_bfr_after (
		.din(n_0341_),
		.dout(new_net_10488)
	);

	bfr new_net_10489_bfr_after (
		.din(new_net_10488),
		.dout(new_net_10489)
	);

	bfr new_net_10490_bfr_after (
		.din(new_net_10489),
		.dout(new_net_10490)
	);

	bfr new_net_10491_bfr_after (
		.din(new_net_10490),
		.dout(new_net_10491)
	);

	bfr new_net_10492_bfr_after (
		.din(new_net_10491),
		.dout(new_net_10492)
	);

	bfr new_net_10493_bfr_after (
		.din(new_net_10492),
		.dout(new_net_10493)
	);

	bfr new_net_10494_bfr_after (
		.din(new_net_10493),
		.dout(new_net_10494)
	);

	bfr new_net_10495_bfr_after (
		.din(new_net_10494),
		.dout(new_net_10495)
	);

	bfr new_net_10496_bfr_after (
		.din(new_net_10495),
		.dout(new_net_10496)
	);

	bfr new_net_10497_bfr_after (
		.din(new_net_10496),
		.dout(new_net_10497)
	);

	bfr new_net_10498_bfr_after (
		.din(new_net_10497),
		.dout(new_net_10498)
	);

	bfr new_net_2448_bfr_after (
		.din(new_net_10498),
		.dout(new_net_2448)
	);

	bfr new_net_2217_bfr_after (
		.din(n_0757_),
		.dout(new_net_2217)
	);

	bfr new_net_10499_bfr_after (
		.din(N130),
		.dout(new_net_10499)
	);

	bfr new_net_10500_bfr_after (
		.din(new_net_10499),
		.dout(new_net_10500)
	);

	bfr new_net_10501_bfr_after (
		.din(new_net_10500),
		.dout(new_net_10501)
	);

	bfr new_net_2238_bfr_after (
		.din(new_net_10501),
		.dout(new_net_2238)
	);

	bfr new_net_10502_bfr_after (
		.din(N115),
		.dout(new_net_10502)
	);

	bfr new_net_10503_bfr_after (
		.din(new_net_10502),
		.dout(new_net_10503)
	);

	bfr new_net_10504_bfr_after (
		.din(new_net_10503),
		.dout(new_net_10504)
	);

	bfr new_net_2259_bfr_after (
		.din(new_net_10504),
		.dout(new_net_2259)
	);

	bfr new_net_10505_bfr_after (
		.din(n_0557_),
		.dout(new_net_10505)
	);

	bfr new_net_10506_bfr_after (
		.din(new_net_10505),
		.dout(new_net_10506)
	);

	bfr new_net_10507_bfr_after (
		.din(new_net_10506),
		.dout(new_net_10507)
	);

	bfr new_net_10508_bfr_after (
		.din(new_net_10507),
		.dout(new_net_10508)
	);

	bfr new_net_2470_bfr_after (
		.din(new_net_10508),
		.dout(new_net_2470)
	);

	bfr new_net_10509_bfr_after (
		.din(N235),
		.dout(new_net_10509)
	);

	bfr new_net_10510_bfr_after (
		.din(new_net_10509),
		.dout(new_net_10510)
	);

	bfr new_net_10511_bfr_after (
		.din(new_net_10510),
		.dout(new_net_10511)
	);

	bfr new_net_2188_bfr_after (
		.din(new_net_10511),
		.dout(new_net_2188)
	);

	bfr new_net_10512_bfr_after (
		.din(new_net_2558),
		.dout(new_net_10512)
	);

	bfr new_net_10513_bfr_after (
		.din(new_net_10512),
		.dout(new_net_10513)
	);

	bfr new_net_10514_bfr_after (
		.din(new_net_10513),
		.dout(new_net_10514)
	);

	bfr new_net_10515_bfr_after (
		.din(new_net_10514),
		.dout(new_net_10515)
	);

	bfr new_net_10516_bfr_after (
		.din(new_net_10515),
		.dout(new_net_10516)
	);

	bfr new_net_10517_bfr_after (
		.din(new_net_10516),
		.dout(new_net_10517)
	);

	bfr new_net_10518_bfr_after (
		.din(new_net_10517),
		.dout(new_net_10518)
	);

	bfr new_net_10519_bfr_after (
		.din(new_net_10518),
		.dout(new_net_10519)
	);

	bfr new_net_10520_bfr_after (
		.din(new_net_10519),
		.dout(new_net_10520)
	);

	bfr new_net_10521_bfr_after (
		.din(new_net_10520),
		.dout(new_net_10521)
	);

	bfr new_net_10522_bfr_after (
		.din(new_net_10521),
		.dout(new_net_10522)
	);

	bfr new_net_10523_bfr_after (
		.din(new_net_10522),
		.dout(new_net_10523)
	);

	bfr new_net_10524_bfr_after (
		.din(new_net_10523),
		.dout(new_net_10524)
	);

	bfr new_net_10525_bfr_after (
		.din(new_net_10524),
		.dout(new_net_10525)
	);

	bfr new_net_10526_bfr_after (
		.din(new_net_10525),
		.dout(new_net_10526)
	);

	bfr new_net_10527_bfr_after (
		.din(new_net_10526),
		.dout(new_net_10527)
	);

	bfr new_net_10528_bfr_after (
		.din(new_net_10527),
		.dout(new_net_10528)
	);

	bfr new_net_10529_bfr_after (
		.din(new_net_10528),
		.dout(new_net_10529)
	);

	bfr new_net_10530_bfr_after (
		.din(new_net_10529),
		.dout(new_net_10530)
	);

	bfr new_net_10531_bfr_after (
		.din(new_net_10530),
		.dout(new_net_10531)
	);

	bfr new_net_10532_bfr_after (
		.din(new_net_10531),
		.dout(new_net_10532)
	);

	bfr new_net_10533_bfr_after (
		.din(new_net_10532),
		.dout(new_net_10533)
	);

	bfr new_net_10534_bfr_after (
		.din(new_net_10533),
		.dout(new_net_10534)
	);

	bfr new_net_10535_bfr_after (
		.din(new_net_10534),
		.dout(new_net_10535)
	);

	bfr new_net_10536_bfr_after (
		.din(new_net_10535),
		.dout(new_net_10536)
	);

	bfr new_net_10537_bfr_after (
		.din(new_net_10536),
		.dout(new_net_10537)
	);

	bfr new_net_10538_bfr_after (
		.din(new_net_10537),
		.dout(new_net_10538)
	);

	bfr new_net_10539_bfr_after (
		.din(new_net_10538),
		.dout(new_net_10539)
	);

	bfr new_net_10540_bfr_after (
		.din(new_net_10539),
		.dout(new_net_10540)
	);

	bfr new_net_10541_bfr_after (
		.din(new_net_10540),
		.dout(new_net_10541)
	);

	bfr new_net_10542_bfr_after (
		.din(new_net_10541),
		.dout(new_net_10542)
	);

	bfr new_net_10543_bfr_after (
		.din(new_net_10542),
		.dout(new_net_10543)
	);

	bfr new_net_10544_bfr_after (
		.din(new_net_10543),
		.dout(new_net_10544)
	);

	bfr new_net_10545_bfr_after (
		.din(new_net_10544),
		.dout(new_net_10545)
	);

	bfr new_net_10546_bfr_after (
		.din(new_net_10545),
		.dout(new_net_10546)
	);

	bfr new_net_10547_bfr_after (
		.din(new_net_10546),
		.dout(new_net_10547)
	);

	bfr new_net_10548_bfr_after (
		.din(new_net_10547),
		.dout(new_net_10548)
	);

	bfr new_net_10549_bfr_after (
		.din(new_net_10548),
		.dout(new_net_10549)
	);

	bfr new_net_10550_bfr_after (
		.din(new_net_10549),
		.dout(new_net_10550)
	);

	bfr new_net_10551_bfr_after (
		.din(new_net_10550),
		.dout(new_net_10551)
	);

	bfr new_net_10552_bfr_after (
		.din(new_net_10551),
		.dout(new_net_10552)
	);

	bfr new_net_10553_bfr_after (
		.din(new_net_10552),
		.dout(new_net_10553)
	);

	bfr new_net_10554_bfr_after (
		.din(new_net_10553),
		.dout(new_net_10554)
	);

	bfr new_net_10555_bfr_after (
		.din(new_net_10554),
		.dout(new_net_10555)
	);

	bfr new_net_10556_bfr_after (
		.din(new_net_10555),
		.dout(new_net_10556)
	);

	bfr new_net_10557_bfr_after (
		.din(new_net_10556),
		.dout(new_net_10557)
	);

	bfr new_net_10558_bfr_after (
		.din(new_net_10557),
		.dout(new_net_10558)
	);

	bfr new_net_10559_bfr_after (
		.din(new_net_10558),
		.dout(new_net_10559)
	);

	bfr N10111_bfr_after (
		.din(new_net_10559),
		.dout(N10111)
	);

	bfr new_net_2409_bfr_after (
		.din(n_0235_),
		.dout(new_net_2409)
	);

	bfr new_net_10560_bfr_after (
		.din(n_0537_),
		.dout(new_net_10560)
	);

	bfr new_net_10561_bfr_after (
		.din(new_net_10560),
		.dout(new_net_10561)
	);

	bfr new_net_10562_bfr_after (
		.din(new_net_10561),
		.dout(new_net_10562)
	);

	bfr new_net_2467_bfr_after (
		.din(new_net_10562),
		.dout(new_net_2467)
	);

	bfr new_net_2284_bfr_after (
		.din(n_0949_),
		.dout(new_net_2284)
	);

	bfr new_net_2196_bfr_after (
		.din(n_0681_),
		.dout(new_net_2196)
	);

	bfr new_net_10563_bfr_after (
		.din(N111),
		.dout(new_net_10563)
	);

	bfr new_net_10564_bfr_after (
		.din(new_net_10563),
		.dout(new_net_10564)
	);

	bfr new_net_10565_bfr_after (
		.din(new_net_10564),
		.dout(new_net_10565)
	);

	bfr new_net_2280_bfr_after (
		.din(new_net_10565),
		.dout(new_net_2280)
	);

	bfr new_net_2343_bfr_after (
		.din(n_1198_),
		.dout(new_net_2343)
	);

	bfr new_net_2439_bfr_after (
		.din(n_0318_),
		.dout(new_net_2439)
	);

	bfr new_net_10566_bfr_after (
		.din(new_net_2515),
		.dout(new_net_10566)
	);

	bfr new_net_10567_bfr_after (
		.din(new_net_10566),
		.dout(new_net_10567)
	);

	bfr new_net_10568_bfr_after (
		.din(new_net_10567),
		.dout(new_net_10568)
	);

	bfr new_net_10569_bfr_after (
		.din(new_net_10568),
		.dout(new_net_10569)
	);

	bfr new_net_10570_bfr_after (
		.din(new_net_10569),
		.dout(new_net_10570)
	);

	bfr new_net_10571_bfr_after (
		.din(new_net_10570),
		.dout(new_net_10571)
	);

	bfr new_net_10572_bfr_after (
		.din(new_net_10571),
		.dout(new_net_10572)
	);

	bfr new_net_10573_bfr_after (
		.din(new_net_10572),
		.dout(new_net_10573)
	);

	bfr new_net_10574_bfr_after (
		.din(new_net_10573),
		.dout(new_net_10574)
	);

	bfr new_net_10575_bfr_after (
		.din(new_net_10574),
		.dout(new_net_10575)
	);

	bfr new_net_10576_bfr_after (
		.din(new_net_10575),
		.dout(new_net_10576)
	);

	bfr new_net_10577_bfr_after (
		.din(new_net_10576),
		.dout(new_net_10577)
	);

	bfr new_net_10578_bfr_after (
		.din(new_net_10577),
		.dout(new_net_10578)
	);

	bfr new_net_10579_bfr_after (
		.din(new_net_10578),
		.dout(new_net_10579)
	);

	bfr new_net_10580_bfr_after (
		.din(new_net_10579),
		.dout(new_net_10580)
	);

	bfr new_net_10581_bfr_after (
		.din(new_net_10580),
		.dout(new_net_10581)
	);

	bfr new_net_10582_bfr_after (
		.din(new_net_10581),
		.dout(new_net_10582)
	);

	bfr new_net_10583_bfr_after (
		.din(new_net_10582),
		.dout(new_net_10583)
	);

	bfr new_net_10584_bfr_after (
		.din(new_net_10583),
		.dout(new_net_10584)
	);

	bfr new_net_10585_bfr_after (
		.din(new_net_10584),
		.dout(new_net_10585)
	);

	bfr new_net_10586_bfr_after (
		.din(new_net_10585),
		.dout(new_net_10586)
	);

	bfr new_net_10587_bfr_after (
		.din(new_net_10586),
		.dout(new_net_10587)
	);

	bfr new_net_10588_bfr_after (
		.din(new_net_10587),
		.dout(new_net_10588)
	);

	bfr new_net_10589_bfr_after (
		.din(new_net_10588),
		.dout(new_net_10589)
	);

	bfr new_net_10590_bfr_after (
		.din(new_net_10589),
		.dout(new_net_10590)
	);

	bfr new_net_10591_bfr_after (
		.din(new_net_10590),
		.dout(new_net_10591)
	);

	bfr new_net_10592_bfr_after (
		.din(new_net_10591),
		.dout(new_net_10592)
	);

	bfr new_net_10593_bfr_after (
		.din(new_net_10592),
		.dout(new_net_10593)
	);

	bfr new_net_10594_bfr_after (
		.din(new_net_10593),
		.dout(new_net_10594)
	);

	bfr new_net_10595_bfr_after (
		.din(new_net_10594),
		.dout(new_net_10595)
	);

	bfr new_net_10596_bfr_after (
		.din(new_net_10595),
		.dout(new_net_10596)
	);

	bfr N10351_bfr_after (
		.din(new_net_10596),
		.dout(N10351)
	);

	bfr new_net_10597_bfr_after (
		.din(new_net_2570),
		.dout(new_net_10597)
	);

	bfr new_net_10598_bfr_after (
		.din(new_net_10597),
		.dout(new_net_10598)
	);

	bfr new_net_10599_bfr_after (
		.din(new_net_10598),
		.dout(new_net_10599)
	);

	bfr new_net_10600_bfr_after (
		.din(new_net_10599),
		.dout(new_net_10600)
	);

	bfr new_net_10601_bfr_after (
		.din(new_net_10600),
		.dout(new_net_10601)
	);

	bfr new_net_10602_bfr_after (
		.din(new_net_10601),
		.dout(new_net_10602)
	);

	bfr new_net_10603_bfr_after (
		.din(new_net_10602),
		.dout(new_net_10603)
	);

	bfr new_net_10604_bfr_after (
		.din(new_net_10603),
		.dout(new_net_10604)
	);

	bfr new_net_10605_bfr_after (
		.din(new_net_10604),
		.dout(new_net_10605)
	);

	bfr new_net_10606_bfr_after (
		.din(new_net_10605),
		.dout(new_net_10606)
	);

	bfr new_net_10607_bfr_after (
		.din(new_net_10606),
		.dout(new_net_10607)
	);

	bfr new_net_10608_bfr_after (
		.din(new_net_10607),
		.dout(new_net_10608)
	);

	bfr new_net_10609_bfr_after (
		.din(new_net_10608),
		.dout(new_net_10609)
	);

	bfr new_net_10610_bfr_after (
		.din(new_net_10609),
		.dout(new_net_10610)
	);

	bfr new_net_10611_bfr_after (
		.din(new_net_10610),
		.dout(new_net_10611)
	);

	bfr new_net_10612_bfr_after (
		.din(new_net_10611),
		.dout(new_net_10612)
	);

	bfr new_net_10613_bfr_after (
		.din(new_net_10612),
		.dout(new_net_10613)
	);

	bfr new_net_10614_bfr_after (
		.din(new_net_10613),
		.dout(new_net_10614)
	);

	bfr new_net_10615_bfr_after (
		.din(new_net_10614),
		.dout(new_net_10615)
	);

	bfr new_net_10616_bfr_after (
		.din(new_net_10615),
		.dout(new_net_10616)
	);

	bfr new_net_10617_bfr_after (
		.din(new_net_10616),
		.dout(new_net_10617)
	);

	bfr new_net_10618_bfr_after (
		.din(new_net_10617),
		.dout(new_net_10618)
	);

	bfr new_net_10619_bfr_after (
		.din(new_net_10618),
		.dout(new_net_10619)
	);

	bfr new_net_10620_bfr_after (
		.din(new_net_10619),
		.dout(new_net_10620)
	);

	bfr new_net_10621_bfr_after (
		.din(new_net_10620),
		.dout(new_net_10621)
	);

	bfr new_net_10622_bfr_after (
		.din(new_net_10621),
		.dout(new_net_10622)
	);

	bfr new_net_10623_bfr_after (
		.din(new_net_10622),
		.dout(new_net_10623)
	);

	bfr new_net_10624_bfr_after (
		.din(new_net_10623),
		.dout(new_net_10624)
	);

	bfr new_net_10625_bfr_after (
		.din(new_net_10624),
		.dout(new_net_10625)
	);

	bfr new_net_10626_bfr_after (
		.din(new_net_10625),
		.dout(new_net_10626)
	);

	bfr new_net_10627_bfr_after (
		.din(new_net_10626),
		.dout(new_net_10627)
	);

	bfr new_net_10628_bfr_after (
		.din(new_net_10627),
		.dout(new_net_10628)
	);

	bfr new_net_10629_bfr_after (
		.din(new_net_10628),
		.dout(new_net_10629)
	);

	bfr new_net_10630_bfr_after (
		.din(new_net_10629),
		.dout(new_net_10630)
	);

	bfr new_net_10631_bfr_after (
		.din(new_net_10630),
		.dout(new_net_10631)
	);

	bfr new_net_10632_bfr_after (
		.din(new_net_10631),
		.dout(new_net_10632)
	);

	bfr new_net_10633_bfr_after (
		.din(new_net_10632),
		.dout(new_net_10633)
	);

	bfr new_net_10634_bfr_after (
		.din(new_net_10633),
		.dout(new_net_10634)
	);

	bfr new_net_10635_bfr_after (
		.din(new_net_10634),
		.dout(new_net_10635)
	);

	bfr new_net_10636_bfr_after (
		.din(new_net_10635),
		.dout(new_net_10636)
	);

	bfr new_net_10637_bfr_after (
		.din(new_net_10636),
		.dout(new_net_10637)
	);

	bfr N10704_bfr_after (
		.din(new_net_10637),
		.dout(N10704)
	);

	bfr new_net_10638_bfr_after (
		.din(n_1346_),
		.dout(new_net_10638)
	);

	bfr new_net_10639_bfr_after (
		.din(new_net_10638),
		.dout(new_net_10639)
	);

	bfr new_net_10640_bfr_after (
		.din(new_net_10639),
		.dout(new_net_10640)
	);

	bfr new_net_2378_bfr_after (
		.din(new_net_10640),
		.dout(new_net_2378)
	);

	bfr new_net_10641_bfr_after (
		.din(N203),
		.dout(new_net_10641)
	);

	bfr new_net_10642_bfr_after (
		.din(new_net_10641),
		.dout(new_net_10642)
	);

	bfr new_net_10643_bfr_after (
		.din(new_net_10642),
		.dout(new_net_10643)
	);

	bfr new_net_2373_bfr_after (
		.din(new_net_10643),
		.dout(new_net_2373)
	);

	bfr new_net_2436_bfr_after (
		.din(n_0308_),
		.dout(new_net_2436)
	);

	bfr new_net_10644_bfr_after (
		.din(N167),
		.dout(new_net_10644)
	);

	bfr new_net_10645_bfr_after (
		.din(new_net_10644),
		.dout(new_net_10645)
	);

	bfr new_net_10646_bfr_after (
		.din(new_net_10645),
		.dout(new_net_10646)
	);

	bfr new_net_2316_bfr_after (
		.din(new_net_10646),
		.dout(new_net_2316)
	);

	bfr new_net_2275_bfr_after (
		.din(n_0888_),
		.dout(new_net_2275)
	);

	bfr new_net_2338_bfr_after (
		.din(n_1184_),
		.dout(new_net_2338)
	);

	bfr new_net_2422_bfr_after (
		.din(n_0270_),
		.dout(new_net_2422)
	);

	bfr new_net_2443_bfr_after (
		.din(n_0330_),
		.dout(new_net_2443)
	);

	bfr new_net_10647_bfr_after (
		.din(N198),
		.dout(new_net_10647)
	);

	bfr new_net_10648_bfr_after (
		.din(new_net_10647),
		.dout(new_net_10648)
	);

	bfr new_net_10649_bfr_after (
		.din(new_net_10648),
		.dout(new_net_10649)
	);

	bfr new_net_2359_bfr_after (
		.din(new_net_10649),
		.dout(new_net_2359)
	);

	bfr new_net_10650_bfr_after (
		.din(N80),
		.dout(new_net_10650)
	);

	bfr new_net_10651_bfr_after (
		.din(new_net_10650),
		.dout(new_net_10651)
	);

	bfr new_net_10652_bfr_after (
		.din(new_net_10651),
		.dout(new_net_10652)
	);

	bfr new_net_2296_bfr_after (
		.din(new_net_10652),
		.dout(new_net_2296)
	);

	bfr new_net_10653_bfr_after (
		.din(n_0003_),
		.dout(new_net_10653)
	);

	bfr new_net_10654_bfr_after (
		.din(new_net_10653),
		.dout(new_net_10654)
	);

	bfr new_net_10655_bfr_after (
		.din(new_net_10654),
		.dout(new_net_10655)
	);

	bfr new_net_10656_bfr_after (
		.din(new_net_10655),
		.dout(new_net_10656)
	);

	bfr new_net_10657_bfr_after (
		.din(new_net_10656),
		.dout(new_net_10657)
	);

	bfr new_net_10658_bfr_after (
		.din(new_net_10657),
		.dout(new_net_10658)
	);

	bfr new_net_10659_bfr_after (
		.din(new_net_10658),
		.dout(new_net_10659)
	);

	bfr new_net_10660_bfr_after (
		.din(new_net_10659),
		.dout(new_net_10660)
	);

	bfr new_net_10661_bfr_after (
		.din(new_net_10660),
		.dout(new_net_10661)
	);

	bfr new_net_10662_bfr_after (
		.din(new_net_10661),
		.dout(new_net_10662)
	);

	bfr new_net_2380_bfr_after (
		.din(new_net_10662),
		.dout(new_net_2380)
	);

	bfr new_net_10663_bfr_after (
		.din(N166),
		.dout(new_net_10663)
	);

	bfr new_net_10664_bfr_after (
		.din(new_net_10663),
		.dout(new_net_10664)
	);

	bfr new_net_10665_bfr_after (
		.din(new_net_10664),
		.dout(new_net_10665)
	);

	bfr new_net_2317_bfr_after (
		.din(new_net_10665),
		.dout(new_net_2317)
	);

	bfr new_net_10666_bfr_after (
		.din(n_0509_),
		.dout(new_net_10666)
	);

	bfr new_net_10667_bfr_after (
		.din(new_net_10666),
		.dout(new_net_10667)
	);

	bfr new_net_10668_bfr_after (
		.din(new_net_10667),
		.dout(new_net_10668)
	);

	bfr new_net_10669_bfr_after (
		.din(new_net_10668),
		.dout(new_net_10669)
	);

	bfr new_net_10670_bfr_after (
		.din(new_net_10669),
		.dout(new_net_10670)
	);

	bfr new_net_10671_bfr_after (
		.din(new_net_10670),
		.dout(new_net_10671)
	);

	bfr new_net_10672_bfr_after (
		.din(new_net_10671),
		.dout(new_net_10672)
	);

	bfr new_net_10673_bfr_after (
		.din(new_net_10672),
		.dout(new_net_10673)
	);

	bfr new_net_10674_bfr_after (
		.din(new_net_10673),
		.dout(new_net_10674)
	);

	bfr new_net_10675_bfr_after (
		.din(new_net_10674),
		.dout(new_net_10675)
	);

	bfr new_net_10676_bfr_after (
		.din(new_net_10675),
		.dout(new_net_10676)
	);

	bfr new_net_10677_bfr_after (
		.din(new_net_10676),
		.dout(new_net_10677)
	);

	bfr new_net_10678_bfr_after (
		.din(new_net_10677),
		.dout(new_net_10678)
	);

	bfr new_net_10679_bfr_after (
		.din(new_net_10678),
		.dout(new_net_10679)
	);

	bfr new_net_10680_bfr_after (
		.din(new_net_10679),
		.dout(new_net_10680)
	);

	bfr new_net_10681_bfr_after (
		.din(new_net_10680),
		.dout(new_net_10681)
	);

	bfr new_net_10682_bfr_after (
		.din(new_net_10681),
		.dout(new_net_10682)
	);

	bfr new_net_10683_bfr_after (
		.din(new_net_10682),
		.dout(new_net_10683)
	);

	bfr new_net_10684_bfr_after (
		.din(new_net_10683),
		.dout(new_net_10684)
	);

	bfr new_net_10685_bfr_after (
		.din(new_net_10684),
		.dout(new_net_10685)
	);

	bfr new_net_10686_bfr_after (
		.din(new_net_10685),
		.dout(new_net_10686)
	);

	bfr new_net_10687_bfr_after (
		.din(new_net_10686),
		.dout(new_net_10687)
	);

	bfr new_net_10688_bfr_after (
		.din(new_net_10687),
		.dout(new_net_10688)
	);

	bfr new_net_10689_bfr_after (
		.din(new_net_10688),
		.dout(new_net_10689)
	);

	bfr new_net_10690_bfr_after (
		.din(new_net_10689),
		.dout(new_net_10690)
	);

	bfr new_net_10691_bfr_after (
		.din(new_net_10690),
		.dout(new_net_10691)
	);

	bfr new_net_10692_bfr_after (
		.din(new_net_10691),
		.dout(new_net_10692)
	);

	bfr new_net_2464_bfr_after (
		.din(new_net_10692),
		.dout(new_net_2464)
	);

	bfr new_net_2485_bfr_after (
		.din(n_0625_),
		.dout(new_net_2485)
	);

endmodule