module multi(a, b, s);
  wire n_000_;
  wire n_001_;
  wire n_002_;
  wire n_003_;
  wire n_004_;
  wire n_005_;
  wire n_006_;
  wire n_007_;
  wire n_008_;
  wire n_009_;
  wire n_010_;
  wire n_011_;
  wire n_012_;
  wire n_013_;
  wire n_014_;
  wire n_015_;
  wire n_016_;
  wire n_017_;
  wire n_018_;
  wire n_019_;
  wire n_020_;
  wire n_021_;
  wire n_022_;
  wire n_023_;
  wire n_024_;
  wire n_025_;
  wire n_026_;
  wire n_027_;
  wire n_028_;
  wire n_029_;
  wire n_030_;
  wire n_031_;
  wire n_032_;
  wire n_033_;
  wire n_034_;
  wire n_035_;
  wire n_036_;
  wire n_037_;
  wire n_038_;
  wire n_039_;
  wire n_040_;
  wire n_041_;
  wire n_042_;
  wire n_043_;
  wire n_044_;
  wire n_045_;
  wire n_046_;
  wire n_047_;
  wire n_048_;
  wire n_049_;
  wire n_050_;
  wire n_051_;
  wire n_052_;
  wire n_053_;
  wire n_054_;
  wire n_055_;
  wire n_056_;
  wire n_057_;
  wire n_058_;
  wire n_059_;
  wire n_060_;
  wire n_061_;
  wire n_062_;
  wire n_063_;
  wire n_064_;
  wire n_065_;
  wire n_066_;
  wire n_067_;
  wire n_068_;
  wire n_069_;
  wire n_070_;
  wire n_071_;
  wire n_072_;
  wire n_073_;
  wire n_074_;
  wire n_075_;
  wire n_076_;
  wire n_077_;
  wire n_078_;
  wire n_079_;
  wire n_080_;
  wire n_081_;
  wire n_082_;
  wire n_083_;
  wire n_084_;
  wire n_085_;
  wire n_086_;
  wire n_087_;
  wire n_088_;
  wire n_089_;
  wire n_090_;
  wire n_091_;
  wire n_092_;
  wire n_093_;
  wire n_094_;
  wire n_095_;
  wire n_096_;
  wire n_097_;
  wire n_098_;
  wire n_099_;
  wire n_100_;
  wire n_101_;
  wire n_102_;
  wire n_103_;
  wire n_104_;
  wire n_105_;
  wire n_106_;
  wire n_107_;
  wire n_108_;
  wire n_109_;
  wire n_110_;
  wire n_111_;
  wire n_112_;
  wire n_113_;
  wire n_114_;
  wire n_115_;
  wire n_116_;
  wire n_117_;
  wire n_118_;
  wire n_119_;
  wire n_120_;
  wire n_121_;
  wire n_122_;
  wire n_123_;
  wire n_124_;
  wire n_125_;
  wire n_126_;
  wire n_127_;
  wire n_128_;
  wire n_129_;
  wire n_130_;
  wire n_131_;
  wire n_132_;
  wire n_133_;
  wire n_134_;
  wire n_135_;
  wire n_136_;
  wire n_137_;
  wire n_138_;
  wire n_139_;
  wire n_140_;
  wire n_141_;
  wire n_142_;
  wire n_143_;
  wire n_144_;
  wire n_145_;
  wire n_146_;
  wire n_147_;
  wire n_148_;
  wire n_149_;
  wire n_150_;
  wire n_151_;
  wire n_152_;
  wire n_153_;
  wire n_154_;
  wire n_155_;
  wire n_156_;
  wire n_157_;
  wire n_158_;
  wire n_159_;
  wire n_160_;
  wire n_161_;
  wire n_162_;
  wire n_163_;
  wire n_164_;
  wire n_165_;
  wire n_166_;
  wire n_167_;
  wire n_168_;
  wire n_169_;
  wire n_170_;
  wire n_171_;
  wire n_172_;
  wire n_173_;
  wire n_174_;
  wire n_175_;
  wire n_176_;
  wire n_177_;
  wire n_178_;
  wire n_179_;
  wire n_180_;
  wire n_181_;
  wire n_182_;
  wire n_183_;
  wire n_184_;
  wire n_185_;
  wire n_186_;
  wire n_187_;
  wire n_188_;
  wire n_189_;
  wire n_190_;
  wire n_191_;
  wire n_192_;
  wire n_193_;
  wire n_194_;
  wire n_195_;
  wire n_196_;
  wire n_197_;
  wire n_198_;
  wire n_199_;
  wire n_200_;
  wire n_201_;
  wire n_202_;
  wire n_203_;
  wire n_204_;
  wire n_205_;
  wire n_206_;
  wire n_207_;
  wire n_208_;
  wire n_209_;
  wire n_210_;
  wire n_211_;
  wire n_212_;
  wire n_213_;
  wire n_214_;
  wire n_215_;
  wire n_216_;
  wire n_217_;
  wire n_218_;
  wire n_219_;
  wire n_220_;
  wire n_221_;
  wire n_222_;
  wire n_223_;
  wire n_224_;
  wire n_225_;
  wire n_226_;
  wire n_227_;
  wire n_228_;
  wire n_229_;
  wire n_230_;
  wire n_231_;
  wire n_232_;
  wire n_233_;
  wire n_234_;
  wire n_235_;
  wire n_236_;
  wire n_237_;
  wire n_238_;
  wire n_239_;
  wire n_240_;
  wire n_241_;
  wire n_242_;
  wire n_243_;
  wire n_244_;
  wire n_245_;
  wire n_246_;
  wire n_247_;
  wire n_248_;
  wire n_249_;
  wire n_250_;
  wire n_251_;
  wire n_252_;
  wire n_253_;
  wire n_254_;
  wire n_255_;
  wire n_256_;
  wire n_257_;
  wire n_258_;
  wire n_259_;
  wire n_260_;
  wire n_261_;
  wire n_262_;
  wire n_263_;
  wire n_264_;
  wire n_265_;
  wire n_266_;
  wire n_267_;
  wire n_268_;
  wire n_269_;
  wire n_270_;
  wire n_271_;
  wire n_272_;
  wire n_273_;
  wire n_274_;
  wire n_275_;
  wire n_276_;
  wire n_277_;
  wire n_278_;
  wire n_279_;
  wire n_280_;
  wire n_281_;
  wire n_282_;
  wire n_283_;
  wire n_284_;
  wire n_285_;
  wire n_286_;
  wire n_287_;
  wire n_288_;
  wire n_289_;
  wire n_290_;
  wire n_291_;
  wire n_292_;
  wire n_293_;
  wire n_294_;
  wire n_295_;
  wire n_296_;
  wire n_297_;
  wire n_298_;
  wire n_299_;
  wire n_300_;
  wire n_301_;
  wire n_302_;
  wire n_303_;
  wire n_304_;
  wire n_305_;
  wire n_306_;
  wire n_307_;
  wire n_308_;
  wire n_309_;
  wire n_310_;
  wire n_311_;
  wire n_312_;
  wire n_313_;
  wire n_314_;
  wire n_315_;
  wire n_316_;
  wire n_317_;
  wire n_318_;
  wire n_319_;
  wire n_320_;
  wire n_321_;
  wire n_322_;
  wire n_323_;
  wire n_324_;
  wire n_325_;
  wire n_326_;
  wire n_327_;
  wire n_328_;
  wire n_329_;
  wire n_330_;
  wire n_331_;
  wire n_332_;
  wire n_333_;
  wire n_334_;
  wire n_335_;
  wire n_336_;
  wire n_337_;
  wire n_338_;
  wire n_339_;
  wire n_340_;
  wire n_341_;
  wire n_342_;
  wire n_343_;
  wire n_344_;
  wire n_345_;
  wire n_346_;
  wire n_347_;
  wire n_348_;
  wire n_349_;
  wire n_350_;
  wire n_351_;
  wire n_352_;
  wire n_353_;
  wire n_354_;
  wire n_355_;
  wire n_356_;
  wire n_357_;
  wire n_358_;
  wire n_359_;
  wire n_360_;
  wire n_361_;
  wire n_362_;
  wire n_363_;
  wire n_364_;
  wire n_365_;
  wire n_366_;
  wire n_367_;
  wire n_368_;
  wire n_369_;
  wire n_370_;
  wire n_371_;
  wire n_372_;
  wire n_373_;
  wire n_374_;
  wire n_375_;
  wire n_376_;
  wire n_377_;
  wire n_378_;
  wire n_379_;
  wire n_380_;
  wire n_381_;
  wire n_382_;
  wire n_383_;
  wire n_384_;
  wire n_385_;
  wire n_386_;
  wire n_387_;
  wire n_388_;
  wire n_389_;
  wire n_390_;
  wire n_391_;
  wire n_392_;
  wire n_393_;
  wire n_394_;
  wire n_395_;
  wire n_396_;
  wire n_397_;
  wire n_398_;
  wire n_399_;
  wire n_400_;
  wire n_401_;
  wire n_402_;
  wire n_403_;
  wire n_404_;
  wire n_405_;
  wire n_406_;
  wire n_407_;
  wire n_408_;
  wire n_409_;
  wire n_410_;
  wire n_411_;
  wire n_412_;
  wire n_413_;
  wire n_414_;
  wire n_415_;
  wire n_416_;
  wire n_417_;
  wire n_418_;
  wire n_419_;
  wire n_420_;
  wire n_421_;
  wire n_422_;
  input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input b_0_;
  input b_1_;
  input b_2_;
  input b_3_;
  input b_4_;
  input b_5_;
  input b_6_;
  input b_7_;
  output s_0_;
  output s_1_;
  output s_2_;
  output s_3_;
  output s_4_;
  output s_5_;
  output s_6_;
  output s_7_;
  output s_8_;
  output s_9_;
  output s_10_;
  output s_11_;
  output s_12_;
  output s_13_;
  output s_14_;
  output s_15_;
  and_bb n_423_ (
    .a(n_391_),
    .b(n_373_),
    .c(n_393_)
  );
  and_bi n_424_ (
    .a(n_392_),
    .b(n_393_),
    .c(s_3_)
  );
  and_ii n_425_ (
    .a(n_389_),
    .b(n_386_),
    .c(n_394_)
  );
  and_bi n_426_ (
    .a(n_380_),
    .b(n_383_),
    .c(n_395_)
  );
  or_ii n_427_ (
    .a(b_2_),
    .b(a_2_),
    .c(n_396_)
  );
  or_ii n_428_ (
    .a(a_3_),
    .b(b_1_),
    .c(n_397_)
  );
  or_ii n_429_ (
    .a(b_0_),
    .b(a_4_),
    .c(n_398_)
  );
  or_bb n_430_ (
    .a(n_398_),
    .b(n_397_),
    .c(n_399_)
  );
  or_ii n_431_ (
    .a(n_398_),
    .b(n_397_),
    .c(n_400_)
  );
  or_ii n_432_ (
    .a(n_400_),
    .b(n_399_),
    .c(n_401_)
  );
  and_ii n_433_ (
    .a(n_401_),
    .b(n_396_),
    .c(n_402_)
  );
  and_bb n_434_ (
    .a(n_401_),
    .b(n_396_),
    .c(n_403_)
  );
  or_bb n_435_ (
    .a(n_403_),
    .b(n_402_),
    .c(n_404_)
  );
  or_bb n_436_ (
    .a(n_404_),
    .b(n_395_),
    .c(n_405_)
  );
  or_ii n_437_ (
    .a(n_404_),
    .b(n_395_),
    .c(n_406_)
  );
  or_ii n_438_ (
    .a(n_406_),
    .b(n_405_),
    .c(n_407_)
  );
  or_ii n_439_ (
    .a(b_4_),
    .b(a_1_),
    .c(n_408_)
  );
  or_bb n_440_ (
    .a(n_408_),
    .b(n_375_),
    .c(n_409_)
  );
  or_ii n_441_ (
    .a(b_3_),
    .b(a_1_),
    .c(n_410_)
  );
  and_bb n_442_ (
    .a(b_4_),
    .b(a_0_),
    .c(n_411_)
  );
  and_bi n_443_ (
    .a(n_410_),
    .b(n_411_),
    .c(n_412_)
  );
  or_bi n_444_ (
    .a(n_412_),
    .b(n_409_),
    .c(n_413_)
  );
  and_ii n_445_ (
    .a(n_413_),
    .b(n_407_),
    .c(n_414_)
  );
  and_bb n_446_ (
    .a(n_413_),
    .b(n_407_),
    .c(n_415_)
  );
  or_bb n_447_ (
    .a(n_415_),
    .b(n_414_),
    .c(n_416_)
  );
  or_bb n_448_ (
    .a(n_416_),
    .b(n_394_),
    .c(n_417_)
  );
  and_bb n_449_ (
    .a(n_416_),
    .b(n_394_),
    .c(n_418_)
  );
  or_bi n_450_ (
    .a(n_418_),
    .b(n_417_),
    .c(n_419_)
  );
  or_bb n_451_ (
    .a(n_419_),
    .b(n_392_),
    .c(n_420_)
  );
  and_bb n_452_ (
    .a(n_419_),
    .b(n_392_),
    .c(n_421_)
  );
  and_bi n_453_ (
    .a(n_420_),
    .b(n_421_),
    .c(s_4_)
  );
  and_bi n_454_ (
    .a(n_405_),
    .b(n_414_),
    .c(n_422_)
  );
  and_bi n_455_ (
    .a(n_399_),
    .b(n_402_),
    .c(n_000_)
  );
  or_ii n_456_ (
    .a(b_2_),
    .b(a_3_),
    .c(n_001_)
  );
  or_ii n_457_ (
    .a(a_4_),
    .b(b_1_),
    .c(n_002_)
  );
  or_ii n_458_ (
    .a(b_0_),
    .b(a_5_),
    .c(n_003_)
  );
  or_bb n_459_ (
    .a(n_003_),
    .b(n_002_),
    .c(n_004_)
  );
  or_ii n_460_ (
    .a(n_003_),
    .b(n_002_),
    .c(n_005_)
  );
  or_ii n_461_ (
    .a(n_005_),
    .b(n_004_),
    .c(n_006_)
  );
  and_ii n_462_ (
    .a(n_006_),
    .b(n_001_),
    .c(n_007_)
  );
  and_bb n_463_ (
    .a(n_006_),
    .b(n_001_),
    .c(n_008_)
  );
  or_bb n_464_ (
    .a(n_008_),
    .b(n_007_),
    .c(n_009_)
  );
  or_bb n_465_ (
    .a(n_009_),
    .b(n_000_),
    .c(n_010_)
  );
  or_ii n_466_ (
    .a(n_009_),
    .b(n_000_),
    .c(n_011_)
  );
  or_ii n_467_ (
    .a(n_011_),
    .b(n_010_),
    .c(n_012_)
  );
  or_ii n_468_ (
    .a(b_5_),
    .b(a_0_),
    .c(n_013_)
  );
  and_bb n_469_ (
    .a(b_3_),
    .b(a_2_),
    .c(n_014_)
  );
  and_bi n_470_ (
    .a(n_014_),
    .b(n_408_),
    .c(n_015_)
  );
  and_bi n_471_ (
    .a(n_408_),
    .b(n_014_),
    .c(n_016_)
  );
  or_bb n_472_ (
    .a(n_016_),
    .b(n_015_),
    .c(n_017_)
  );
  and_ii n_473_ (
    .a(n_017_),
    .b(n_013_),
    .c(n_018_)
  );
  and_bb n_474_ (
    .a(n_017_),
    .b(n_013_),
    .c(n_019_)
  );
  or_bb n_475_ (
    .a(n_019_),
    .b(n_018_),
    .c(n_020_)
  );
  and_ii n_476_ (
    .a(n_020_),
    .b(n_012_),
    .c(n_021_)
  );
  and_bb n_477_ (
    .a(n_020_),
    .b(n_012_),
    .c(n_022_)
  );
  or_bb n_478_ (
    .a(n_022_),
    .b(n_021_),
    .c(n_023_)
  );
  or_bb n_479_ (
    .a(n_023_),
    .b(n_422_),
    .c(n_024_)
  );
  or_ii n_480_ (
    .a(n_023_),
    .b(n_422_),
    .c(n_025_)
  );
  or_ii n_481_ (
    .a(n_025_),
    .b(n_024_),
    .c(n_026_)
  );
  and_ii n_482_ (
    .a(n_026_),
    .b(n_409_),
    .c(n_027_)
  );
  and_bb n_483_ (
    .a(n_026_),
    .b(n_409_),
    .c(n_028_)
  );
  or_bb n_484_ (
    .a(n_028_),
    .b(n_027_),
    .c(n_029_)
  );
  or_bb n_485_ (
    .a(n_029_),
    .b(n_417_),
    .c(n_030_)
  );
  and_bb n_486_ (
    .a(n_029_),
    .b(n_417_),
    .c(n_031_)
  );
  or_bi n_487_ (
    .a(n_031_),
    .b(n_030_),
    .c(n_032_)
  );
  or_bb n_488_ (
    .a(n_032_),
    .b(n_420_),
    .c(n_033_)
  );
  and_bb n_489_ (
    .a(n_032_),
    .b(n_420_),
    .c(n_034_)
  );
  and_bi n_490_ (
    .a(n_033_),
    .b(n_034_),
    .c(s_5_)
  );
  and_bi n_491_ (
    .a(n_024_),
    .b(n_027_),
    .c(n_035_)
  );
  and_bi n_492_ (
    .a(n_010_),
    .b(n_021_),
    .c(n_036_)
  );
  and_bi n_493_ (
    .a(n_004_),
    .b(n_007_),
    .c(n_037_)
  );
  or_ii n_494_ (
    .a(b_2_),
    .b(a_4_),
    .c(n_038_)
  );
  or_ii n_495_ (
    .a(a_6_),
    .b(b_1_),
    .c(n_039_)
  );
  or_bb n_496_ (
    .a(n_039_),
    .b(n_003_),
    .c(n_040_)
  );
  or_ii n_497_ (
    .a(a_5_),
    .b(b_1_),
    .c(n_041_)
  );
  and_bb n_498_ (
    .a(b_0_),
    .b(a_6_),
    .c(n_042_)
  );
  or_bi n_499_ (
    .a(n_042_),
    .b(n_041_),
    .c(n_043_)
  );
  or_ii n_500_ (
    .a(n_043_),
    .b(n_040_),
    .c(n_044_)
  );
  and_ii n_501_ (
    .a(n_044_),
    .b(n_038_),
    .c(n_045_)
  );
  and_bb n_502_ (
    .a(n_044_),
    .b(n_038_),
    .c(n_046_)
  );
  or_bb n_503_ (
    .a(n_046_),
    .b(n_045_),
    .c(n_047_)
  );
  or_bb n_504_ (
    .a(n_047_),
    .b(n_037_),
    .c(n_048_)
  );
  or_ii n_505_ (
    .a(n_047_),
    .b(n_037_),
    .c(n_049_)
  );
  or_ii n_506_ (
    .a(n_049_),
    .b(n_048_),
    .c(n_050_)
  );
  or_ii n_507_ (
    .a(b_5_),
    .b(a_1_),
    .c(n_051_)
  );
  or_ii n_508_ (
    .a(b_4_),
    .b(a_2_),
    .c(n_052_)
  );
  or_ii n_509_ (
    .a(b_3_),
    .b(a_3_),
    .c(n_053_)
  );
  or_bb n_510_ (
    .a(n_053_),
    .b(n_052_),
    .c(n_054_)
  );
  or_ii n_511_ (
    .a(n_053_),
    .b(n_052_),
    .c(n_055_)
  );
  or_ii n_512_ (
    .a(n_055_),
    .b(n_054_),
    .c(n_056_)
  );
  and_ii n_513_ (
    .a(n_056_),
    .b(n_051_),
    .c(n_057_)
  );
  and_bb n_514_ (
    .a(n_056_),
    .b(n_051_),
    .c(n_058_)
  );
  or_bb n_515_ (
    .a(n_058_),
    .b(n_057_),
    .c(n_059_)
  );
  and_ii n_516_ (
    .a(n_059_),
    .b(n_050_),
    .c(n_060_)
  );
  and_bb n_517_ (
    .a(n_059_),
    .b(n_050_),
    .c(n_061_)
  );
  or_bb n_518_ (
    .a(n_061_),
    .b(n_060_),
    .c(n_062_)
  );
  or_bb n_519_ (
    .a(n_062_),
    .b(n_036_),
    .c(n_063_)
  );
  or_ii n_520_ (
    .a(n_062_),
    .b(n_036_),
    .c(n_064_)
  );
  or_ii n_521_ (
    .a(n_064_),
    .b(n_063_),
    .c(n_065_)
  );
  and_ii n_522_ (
    .a(n_018_),
    .b(n_015_),
    .c(n_066_)
  );
  or_ii n_523_ (
    .a(b_6_),
    .b(a_0_),
    .c(n_067_)
  );
  or_bb n_524_ (
    .a(n_067_),
    .b(n_066_),
    .c(n_068_)
  );
  and_bb n_525_ (
    .a(n_067_),
    .b(n_066_),
    .c(n_069_)
  );
  or_bi n_526_ (
    .a(n_069_),
    .b(n_068_),
    .c(n_070_)
  );
  and_ii n_527_ (
    .a(n_070_),
    .b(n_065_),
    .c(n_071_)
  );
  and_bb n_528_ (
    .a(n_070_),
    .b(n_065_),
    .c(n_072_)
  );
  or_bb n_529_ (
    .a(n_072_),
    .b(n_071_),
    .c(n_073_)
  );
  or_bb n_530_ (
    .a(n_073_),
    .b(n_035_),
    .c(n_074_)
  );
  and_bb n_531_ (
    .a(n_073_),
    .b(n_035_),
    .c(n_075_)
  );
  or_bi n_532_ (
    .a(n_075_),
    .b(n_074_),
    .c(n_076_)
  );
  or_bb n_533_ (
    .a(n_076_),
    .b(n_030_),
    .c(n_077_)
  );
  or_ii n_534_ (
    .a(n_076_),
    .b(n_030_),
    .c(n_078_)
  );
  or_ii n_535_ (
    .a(n_078_),
    .b(n_077_),
    .c(n_079_)
  );
  and_ii n_536_ (
    .a(n_079_),
    .b(n_033_),
    .c(n_080_)
  );
  and_bb n_537_ (
    .a(n_079_),
    .b(n_033_),
    .c(n_081_)
  );
  and_ii n_538_ (
    .a(n_081_),
    .b(n_080_),
    .c(s_6_)
  );
  and_bi n_539_ (
    .a(n_077_),
    .b(n_080_),
    .c(n_082_)
  );
  and_bi n_540_ (
    .a(n_063_),
    .b(n_071_),
    .c(n_083_)
  );
  and_bi n_541_ (
    .a(n_048_),
    .b(n_060_),
    .c(n_084_)
  );
  and_bi n_542_ (
    .a(n_040_),
    .b(n_045_),
    .c(n_085_)
  );
  or_ii n_543_ (
    .a(b_2_),
    .b(a_5_),
    .c(n_086_)
  );
  or_ii n_544_ (
    .a(b_0_),
    .b(a_7_),
    .c(n_087_)
  );
  or_bb n_545_ (
    .a(n_087_),
    .b(n_039_),
    .c(n_088_)
  );
  or_ii n_546_ (
    .a(n_087_),
    .b(n_039_),
    .c(n_089_)
  );
  or_ii n_547_ (
    .a(n_089_),
    .b(n_088_),
    .c(n_090_)
  );
  and_ii n_548_ (
    .a(n_090_),
    .b(n_086_),
    .c(n_091_)
  );
  and_bb n_549_ (
    .a(n_090_),
    .b(n_086_),
    .c(n_092_)
  );
  or_bb n_550_ (
    .a(n_092_),
    .b(n_091_),
    .c(n_093_)
  );
  or_bb n_551_ (
    .a(n_093_),
    .b(n_085_),
    .c(n_094_)
  );
  or_ii n_552_ (
    .a(n_093_),
    .b(n_085_),
    .c(n_095_)
  );
  or_ii n_553_ (
    .a(n_095_),
    .b(n_094_),
    .c(n_096_)
  );
  or_ii n_554_ (
    .a(b_5_),
    .b(a_2_),
    .c(n_097_)
  );
  or_ii n_555_ (
    .a(b_4_),
    .b(a_3_),
    .c(n_098_)
  );
  and_bb n_556_ (
    .a(b_3_),
    .b(a_4_),
    .c(n_099_)
  );
  and_bi n_557_ (
    .a(n_099_),
    .b(n_098_),
    .c(n_100_)
  );
  and_bi n_558_ (
    .a(n_098_),
    .b(n_099_),
    .c(n_101_)
  );
  or_bb n_559_ (
    .a(n_101_),
    .b(n_100_),
    .c(n_102_)
  );
  and_ii n_560_ (
    .a(n_102_),
    .b(n_097_),
    .c(n_103_)
  );
  and_bb n_561_ (
    .a(n_102_),
    .b(n_097_),
    .c(n_104_)
  );
  or_bb n_562_ (
    .a(n_104_),
    .b(n_103_),
    .c(n_105_)
  );
  and_ii n_563_ (
    .a(n_105_),
    .b(n_096_),
    .c(n_106_)
  );
  and_bb n_564_ (
    .a(n_105_),
    .b(n_096_),
    .c(n_107_)
  );
  or_bb n_565_ (
    .a(n_107_),
    .b(n_106_),
    .c(n_108_)
  );
  or_bb n_566_ (
    .a(n_108_),
    .b(n_084_),
    .c(n_109_)
  );
  or_ii n_567_ (
    .a(n_108_),
    .b(n_084_),
    .c(n_110_)
  );
  or_ii n_568_ (
    .a(n_110_),
    .b(n_109_),
    .c(n_111_)
  );
  or_ii n_569_ (
    .a(b_7_),
    .b(a_0_),
    .c(n_112_)
  );
  and_bi n_570_ (
    .a(n_054_),
    .b(n_057_),
    .c(n_113_)
  );
  or_ii n_571_ (
    .a(b_6_),
    .b(a_1_),
    .c(n_114_)
  );
  and_ii n_572_ (
    .a(n_114_),
    .b(n_113_),
    .c(n_115_)
  );
  and_bb n_573_ (
    .a(n_114_),
    .b(n_113_),
    .c(n_116_)
  );
  or_bb n_574_ (
    .a(n_116_),
    .b(n_115_),
    .c(n_117_)
  );
  and_ii n_575_ (
    .a(n_117_),
    .b(n_112_),
    .c(n_118_)
  );
  and_bb n_576_ (
    .a(n_117_),
    .b(n_112_),
    .c(n_119_)
  );
  or_bb n_577_ (
    .a(n_119_),
    .b(n_118_),
    .c(n_120_)
  );
  and_ii n_578_ (
    .a(n_120_),
    .b(n_111_),
    .c(n_121_)
  );
  and_bb n_579_ (
    .a(n_120_),
    .b(n_111_),
    .c(n_122_)
  );
  or_bb n_580_ (
    .a(n_122_),
    .b(n_121_),
    .c(n_123_)
  );
  or_bb n_581_ (
    .a(n_123_),
    .b(n_083_),
    .c(n_124_)
  );
  or_ii n_582_ (
    .a(n_123_),
    .b(n_083_),
    .c(n_125_)
  );
  or_ii n_583_ (
    .a(n_125_),
    .b(n_124_),
    .c(n_126_)
  );
  and_ii n_584_ (
    .a(n_126_),
    .b(n_068_),
    .c(n_127_)
  );
  and_bb n_585_ (
    .a(n_126_),
    .b(n_068_),
    .c(n_128_)
  );
  or_bb n_586_ (
    .a(n_128_),
    .b(n_127_),
    .c(n_129_)
  );
  or_bb n_587_ (
    .a(n_129_),
    .b(n_074_),
    .c(n_130_)
  );
  or_ii n_588_ (
    .a(n_129_),
    .b(n_074_),
    .c(n_131_)
  );
  or_ii n_589_ (
    .a(n_131_),
    .b(n_130_),
    .c(n_132_)
  );
  and_ii n_590_ (
    .a(n_132_),
    .b(n_082_),
    .c(n_133_)
  );
  and_bb n_591_ (
    .a(n_132_),
    .b(n_082_),
    .c(n_134_)
  );
  and_ii n_592_ (
    .a(n_134_),
    .b(n_133_),
    .c(s_7_)
  );
  and_bi n_593_ (
    .a(n_130_),
    .b(n_133_),
    .c(n_135_)
  );
  and_bi n_594_ (
    .a(n_124_),
    .b(n_127_),
    .c(n_136_)
  );
  and_ii n_595_ (
    .a(n_118_),
    .b(n_115_),
    .c(n_137_)
  );
  and_bi n_596_ (
    .a(n_109_),
    .b(n_121_),
    .c(n_138_)
  );
  and_bi n_597_ (
    .a(n_094_),
    .b(n_106_),
    .c(n_139_)
  );
  and_bi n_598_ (
    .a(n_088_),
    .b(n_091_),
    .c(n_140_)
  );
  or_ii n_599_ (
    .a(b_2_),
    .b(a_7_),
    .c(n_141_)
  );
  and_ii n_600_ (
    .a(n_141_),
    .b(n_039_),
    .c(n_142_)
  );
  or_ii n_601_ (
    .a(a_7_),
    .b(b_1_),
    .c(n_143_)
  );
  and_bb n_602_ (
    .a(b_2_),
    .b(a_6_),
    .c(n_144_)
  );
  and_bi n_603_ (
    .a(n_143_),
    .b(n_144_),
    .c(n_145_)
  );
  or_bb n_604_ (
    .a(n_145_),
    .b(n_142_),
    .c(n_146_)
  );
  and_ii n_605_ (
    .a(n_146_),
    .b(n_140_),
    .c(n_147_)
  );
  and_bb n_606_ (
    .a(n_146_),
    .b(n_140_),
    .c(n_148_)
  );
  or_bb n_607_ (
    .a(n_148_),
    .b(n_147_),
    .c(n_149_)
  );
  or_ii n_608_ (
    .a(b_5_),
    .b(a_3_),
    .c(n_150_)
  );
  or_ii n_609_ (
    .a(b_4_),
    .b(a_4_),
    .c(n_151_)
  );
  and_bb n_610_ (
    .a(b_3_),
    .b(a_5_),
    .c(n_152_)
  );
  and_bi n_611_ (
    .a(n_152_),
    .b(n_151_),
    .c(n_153_)
  );
  and_bi n_612_ (
    .a(n_151_),
    .b(n_152_),
    .c(n_154_)
  );
  or_bb n_613_ (
    .a(n_154_),
    .b(n_153_),
    .c(n_155_)
  );
  and_ii n_614_ (
    .a(n_155_),
    .b(n_150_),
    .c(n_156_)
  );
  and_bb n_615_ (
    .a(n_155_),
    .b(n_150_),
    .c(n_157_)
  );
  or_bb n_616_ (
    .a(n_157_),
    .b(n_156_),
    .c(n_158_)
  );
  and_ii n_617_ (
    .a(n_158_),
    .b(n_149_),
    .c(n_159_)
  );
  and_bb n_618_ (
    .a(n_158_),
    .b(n_149_),
    .c(n_160_)
  );
  or_bb n_619_ (
    .a(n_160_),
    .b(n_159_),
    .c(n_161_)
  );
  and_ii n_620_ (
    .a(n_161_),
    .b(n_139_),
    .c(n_162_)
  );
  and_bb n_621_ (
    .a(n_161_),
    .b(n_139_),
    .c(n_163_)
  );
  or_bb n_622_ (
    .a(n_163_),
    .b(n_162_),
    .c(n_164_)
  );
  or_ii n_623_ (
    .a(b_7_),
    .b(a_1_),
    .c(n_165_)
  );
  and_ii n_624_ (
    .a(n_103_),
    .b(n_100_),
    .c(n_166_)
  );
  or_ii n_625_ (
    .a(b_6_),
    .b(a_2_),
    .c(n_167_)
  );
  and_ii n_626_ (
    .a(n_167_),
    .b(n_166_),
    .c(n_168_)
  );
  and_bb n_627_ (
    .a(n_167_),
    .b(n_166_),
    .c(n_169_)
  );
  or_bb n_628_ (
    .a(n_169_),
    .b(n_168_),
    .c(n_170_)
  );
  and_ii n_629_ (
    .a(n_170_),
    .b(n_165_),
    .c(n_171_)
  );
  and_bb n_630_ (
    .a(n_170_),
    .b(n_165_),
    .c(n_172_)
  );
  or_bb n_631_ (
    .a(n_172_),
    .b(n_171_),
    .c(n_173_)
  );
  and_ii n_632_ (
    .a(n_173_),
    .b(n_164_),
    .c(n_174_)
  );
  and_bb n_633_ (
    .a(n_173_),
    .b(n_164_),
    .c(n_175_)
  );
  or_bb n_634_ (
    .a(n_175_),
    .b(n_174_),
    .c(n_176_)
  );
  and_ii n_635_ (
    .a(n_176_),
    .b(n_138_),
    .c(n_177_)
  );
  and_bb n_636_ (
    .a(n_176_),
    .b(n_138_),
    .c(n_178_)
  );
  or_bb n_637_ (
    .a(n_178_),
    .b(n_177_),
    .c(n_179_)
  );
  and_ii n_638_ (
    .a(n_179_),
    .b(n_137_),
    .c(n_180_)
  );
  and_bb n_639_ (
    .a(n_179_),
    .b(n_137_),
    .c(n_181_)
  );
  or_bb n_640_ (
    .a(n_181_),
    .b(n_180_),
    .c(n_182_)
  );
  and_ii n_641_ (
    .a(n_182_),
    .b(n_136_),
    .c(n_183_)
  );
  and_bb n_642_ (
    .a(n_182_),
    .b(n_136_),
    .c(n_184_)
  );
  or_bb n_643_ (
    .a(n_184_),
    .b(n_183_),
    .c(n_185_)
  );
  and_ii n_644_ (
    .a(n_185_),
    .b(n_135_),
    .c(n_186_)
  );
  and_bb n_645_ (
    .a(n_185_),
    .b(n_135_),
    .c(n_187_)
  );
  and_ii n_646_ (
    .a(n_187_),
    .b(n_186_),
    .c(s_8_)
  );
  or_bb n_647_ (
    .a(n_186_),
    .b(n_183_),
    .c(n_188_)
  );
  and_ii n_648_ (
    .a(n_180_),
    .b(n_177_),
    .c(n_189_)
  );
  and_ii n_649_ (
    .a(n_171_),
    .b(n_168_),
    .c(n_190_)
  );
  and_ii n_650_ (
    .a(n_174_),
    .b(n_162_),
    .c(n_191_)
  );
  and_ii n_651_ (
    .a(n_159_),
    .b(n_147_),
    .c(n_192_)
  );
  or_bi n_652_ (
    .a(n_141_),
    .b(n_039_),
    .c(n_193_)
  );
  or_ii n_653_ (
    .a(b_5_),
    .b(a_4_),
    .c(n_194_)
  );
  or_ii n_654_ (
    .a(b_4_),
    .b(a_6_),
    .c(n_195_)
  );
  and_bi n_655_ (
    .a(n_152_),
    .b(n_195_),
    .c(n_196_)
  );
  or_ii n_656_ (
    .a(b_4_),
    .b(a_5_),
    .c(n_197_)
  );
  and_bb n_657_ (
    .a(b_3_),
    .b(a_6_),
    .c(n_198_)
  );
  and_bi n_658_ (
    .a(n_197_),
    .b(n_198_),
    .c(n_199_)
  );
  or_bb n_659_ (
    .a(n_199_),
    .b(n_196_),
    .c(n_200_)
  );
  and_ii n_660_ (
    .a(n_200_),
    .b(n_194_),
    .c(n_201_)
  );
  and_bb n_661_ (
    .a(n_200_),
    .b(n_194_),
    .c(n_202_)
  );
  or_bb n_662_ (
    .a(n_202_),
    .b(n_201_),
    .c(n_203_)
  );
  and_ii n_663_ (
    .a(n_203_),
    .b(n_193_),
    .c(n_204_)
  );
  and_bb n_664_ (
    .a(n_203_),
    .b(n_193_),
    .c(n_205_)
  );
  or_bb n_665_ (
    .a(n_205_),
    .b(n_204_),
    .c(n_206_)
  );
  and_ii n_666_ (
    .a(n_206_),
    .b(n_192_),
    .c(n_207_)
  );
  and_bb n_667_ (
    .a(n_206_),
    .b(n_192_),
    .c(n_208_)
  );
  or_bb n_668_ (
    .a(n_208_),
    .b(n_207_),
    .c(n_209_)
  );
  or_ii n_669_ (
    .a(b_7_),
    .b(a_2_),
    .c(n_210_)
  );
  and_ii n_670_ (
    .a(n_156_),
    .b(n_153_),
    .c(n_211_)
  );
  or_ii n_671_ (
    .a(b_6_),
    .b(a_3_),
    .c(n_212_)
  );
  and_ii n_672_ (
    .a(n_212_),
    .b(n_211_),
    .c(n_213_)
  );
  and_bb n_673_ (
    .a(n_212_),
    .b(n_211_),
    .c(n_214_)
  );
  or_bb n_674_ (
    .a(n_214_),
    .b(n_213_),
    .c(n_215_)
  );
  and_ii n_675_ (
    .a(n_215_),
    .b(n_210_),
    .c(n_216_)
  );
  and_bb n_676_ (
    .a(n_215_),
    .b(n_210_),
    .c(n_217_)
  );
  or_bb n_677_ (
    .a(n_217_),
    .b(n_216_),
    .c(n_218_)
  );
  and_ii n_678_ (
    .a(n_218_),
    .b(n_209_),
    .c(n_219_)
  );
  and_bb n_679_ (
    .a(n_218_),
    .b(n_209_),
    .c(n_220_)
  );
  or_bb n_680_ (
    .a(n_220_),
    .b(n_219_),
    .c(n_221_)
  );
  and_ii n_681_ (
    .a(n_221_),
    .b(n_191_),
    .c(n_222_)
  );
  and_bb n_682_ (
    .a(n_221_),
    .b(n_191_),
    .c(n_223_)
  );
  or_bb n_683_ (
    .a(n_223_),
    .b(n_222_),
    .c(n_224_)
  );
  and_ii n_684_ (
    .a(n_224_),
    .b(n_190_),
    .c(n_225_)
  );
  and_bb n_685_ (
    .a(n_224_),
    .b(n_190_),
    .c(n_227_)
  );
  and_ii n_686_ (
    .a(n_227_),
    .b(n_225_),
    .c(n_228_)
  );
  and_bi n_687_ (
    .a(n_228_),
    .b(n_189_),
    .c(n_229_)
  );
  and_bi n_688_ (
    .a(n_189_),
    .b(n_228_),
    .c(n_230_)
  );
  and_ii n_689_ (
    .a(n_230_),
    .b(n_229_),
    .c(n_231_)
  );
  or_bb n_690_ (
    .a(n_231_),
    .b(n_188_),
    .c(n_232_)
  );
  and_bb n_691_ (
    .a(n_231_),
    .b(n_188_),
    .c(n_233_)
  );
  and_bi n_692_ (
    .a(n_232_),
    .b(n_233_),
    .c(s_9_)
  );
  and_ii n_693_ (
    .a(n_225_),
    .b(n_222_),
    .c(n_234_)
  );
  and_ii n_694_ (
    .a(n_216_),
    .b(n_213_),
    .c(n_235_)
  );
  and_ii n_695_ (
    .a(n_219_),
    .b(n_207_),
    .c(n_237_)
  );
  and_ii n_696_ (
    .a(n_204_),
    .b(n_142_),
    .c(n_238_)
  );
  or_ii n_697_ (
    .a(b_5_),
    .b(a_5_),
    .c(n_239_)
  );
  or_ii n_698_ (
    .a(b_4_),
    .b(a_7_),
    .c(n_240_)
  );
  and_bi n_699_ (
    .a(n_198_),
    .b(n_240_),
    .c(n_241_)
  );
  and_bb n_700_ (
    .a(b_3_),
    .b(a_7_),
    .c(n_242_)
  );
  and_bi n_701_ (
    .a(n_195_),
    .b(n_242_),
    .c(n_243_)
  );
  or_bb n_702_ (
    .a(n_243_),
    .b(n_241_),
    .c(n_244_)
  );
  and_ii n_703_ (
    .a(n_244_),
    .b(n_239_),
    .c(n_245_)
  );
  and_bb n_704_ (
    .a(n_244_),
    .b(n_239_),
    .c(n_246_)
  );
  or_bb n_705_ (
    .a(n_246_),
    .b(n_245_),
    .c(n_247_)
  );
  and_ii n_706_ (
    .a(n_247_),
    .b(n_238_),
    .c(n_248_)
  );
  and_bb n_707_ (
    .a(n_247_),
    .b(n_238_),
    .c(n_249_)
  );
  or_bb n_708_ (
    .a(n_249_),
    .b(n_248_),
    .c(n_250_)
  );
  or_ii n_709_ (
    .a(b_7_),
    .b(a_3_),
    .c(n_251_)
  );
  and_ii n_710_ (
    .a(n_201_),
    .b(n_196_),
    .c(n_252_)
  );
  or_ii n_711_ (
    .a(b_6_),
    .b(a_4_),
    .c(n_253_)
  );
  and_ii n_712_ (
    .a(n_253_),
    .b(n_252_),
    .c(n_254_)
  );
  and_bb n_713_ (
    .a(n_253_),
    .b(n_252_),
    .c(n_255_)
  );
  or_bb n_714_ (
    .a(n_255_),
    .b(n_254_),
    .c(n_256_)
  );
  and_ii n_715_ (
    .a(n_256_),
    .b(n_251_),
    .c(n_259_)
  );
  and_bb n_716_ (
    .a(n_256_),
    .b(n_251_),
    .c(n_260_)
  );
  or_bb n_717_ (
    .a(n_260_),
    .b(n_259_),
    .c(n_261_)
  );
  and_ii n_718_ (
    .a(n_261_),
    .b(n_250_),
    .c(n_262_)
  );
  and_bb n_719_ (
    .a(n_261_),
    .b(n_250_),
    .c(n_263_)
  );
  or_bb n_720_ (
    .a(n_263_),
    .b(n_262_),
    .c(n_264_)
  );
  and_ii n_721_ (
    .a(n_264_),
    .b(n_237_),
    .c(n_265_)
  );
  and_bb n_722_ (
    .a(n_264_),
    .b(n_237_),
    .c(n_266_)
  );
  or_bb n_723_ (
    .a(n_266_),
    .b(n_265_),
    .c(n_267_)
  );
  and_ii n_724_ (
    .a(n_267_),
    .b(n_235_),
    .c(n_268_)
  );
  and_bb n_725_ (
    .a(n_267_),
    .b(n_235_),
    .c(n_269_)
  );
  or_bb n_726_ (
    .a(n_269_),
    .b(n_268_),
    .c(n_270_)
  );
  and_ii n_727_ (
    .a(n_270_),
    .b(n_234_),
    .c(n_271_)
  );
  and_bb n_728_ (
    .a(n_270_),
    .b(n_234_),
    .c(n_272_)
  );
  or_bb n_729_ (
    .a(n_272_),
    .b(n_271_),
    .c(n_273_)
  );
  and_ii n_730_ (
    .a(n_229_),
    .b(n_188_),
    .c(n_274_)
  );
  or_bb n_731_ (
    .a(n_274_),
    .b(n_230_),
    .c(n_275_)
  );
  and_ii n_732_ (
    .a(n_275_),
    .b(n_273_),
    .c(n_276_)
  );
  and_bb n_733_ (
    .a(n_275_),
    .b(n_273_),
    .c(n_277_)
  );
  and_ii n_734_ (
    .a(n_277_),
    .b(n_276_),
    .c(s_10_)
  );
  and_ii n_735_ (
    .a(n_276_),
    .b(n_271_),
    .c(n_279_)
  );
  and_ii n_736_ (
    .a(n_268_),
    .b(n_265_),
    .c(n_280_)
  );
  and_ii n_737_ (
    .a(n_259_),
    .b(n_254_),
    .c(n_281_)
  );
  and_ii n_738_ (
    .a(n_262_),
    .b(n_248_),
    .c(n_282_)
  );
  or_ii n_739_ (
    .a(b_5_),
    .b(a_7_),
    .c(n_283_)
  );
  or_bb n_740_ (
    .a(n_283_),
    .b(n_195_),
    .c(n_284_)
  );
  and_bb n_741_ (
    .a(b_5_),
    .b(a_6_),
    .c(n_285_)
  );
  and_bi n_742_ (
    .a(n_240_),
    .b(n_285_),
    .c(n_286_)
  );
  or_bi n_743_ (
    .a(n_286_),
    .b(n_284_),
    .c(n_287_)
  );
  or_ii n_744_ (
    .a(b_7_),
    .b(a_4_),
    .c(n_288_)
  );
  and_ii n_745_ (
    .a(n_245_),
    .b(n_241_),
    .c(n_290_)
  );
  or_ii n_746_ (
    .a(b_6_),
    .b(a_5_),
    .c(n_291_)
  );
  and_ii n_747_ (
    .a(n_291_),
    .b(n_290_),
    .c(n_292_)
  );
  and_bb n_748_ (
    .a(n_291_),
    .b(n_290_),
    .c(n_293_)
  );
  or_bb n_749_ (
    .a(n_293_),
    .b(n_292_),
    .c(n_294_)
  );
  and_ii n_750_ (
    .a(n_294_),
    .b(n_288_),
    .c(n_295_)
  );
  and_bb n_751_ (
    .a(n_294_),
    .b(n_288_),
    .c(n_296_)
  );
  or_bb n_752_ (
    .a(n_296_),
    .b(n_295_),
    .c(n_297_)
  );
  or_bb n_753_ (
    .a(n_297_),
    .b(n_287_),
    .c(n_298_)
  );
  and_bb n_754_ (
    .a(n_297_),
    .b(n_287_),
    .c(n_299_)
  );
  or_bi n_755_ (
    .a(n_299_),
    .b(n_298_),
    .c(n_301_)
  );
  and_ii n_756_ (
    .a(n_301_),
    .b(n_282_),
    .c(n_302_)
  );
  and_bb n_757_ (
    .a(n_301_),
    .b(n_282_),
    .c(n_303_)
  );
  or_bb n_758_ (
    .a(n_303_),
    .b(n_302_),
    .c(n_304_)
  );
  and_ii n_759_ (
    .a(n_304_),
    .b(n_281_),
    .c(n_305_)
  );
  and_bb n_760_ (
    .a(n_304_),
    .b(n_281_),
    .c(n_306_)
  );
  or_bb n_761_ (
    .a(n_306_),
    .b(n_305_),
    .c(n_307_)
  );
  and_ii n_762_ (
    .a(n_307_),
    .b(n_280_),
    .c(n_308_)
  );
  and_bb n_763_ (
    .a(n_307_),
    .b(n_280_),
    .c(n_309_)
  );
  or_bb n_764_ (
    .a(n_309_),
    .b(n_308_),
    .c(n_310_)
  );
  and_ii n_765_ (
    .a(n_310_),
    .b(n_279_),
    .c(n_312_)
  );
  and_bb n_766_ (
    .a(n_310_),
    .b(n_279_),
    .c(n_313_)
  );
  and_ii n_767_ (
    .a(n_313_),
    .b(n_312_),
    .c(s_11_)
  );
  and_ii n_768_ (
    .a(n_312_),
    .b(n_308_),
    .c(n_314_)
  );
  and_ii n_769_ (
    .a(n_305_),
    .b(n_302_),
    .c(n_315_)
  );
  and_ii n_770_ (
    .a(n_295_),
    .b(n_292_),
    .c(n_316_)
  );
  or_ii n_771_ (
    .a(b_7_),
    .b(a_5_),
    .c(n_317_)
  );
  and_bi n_772_ (
    .a(b_6_),
    .b(n_284_),
    .c(n_318_)
  );
  and_bb n_773_ (
    .a(b_6_),
    .b(a_6_),
    .c(n_319_)
  );
  and_bi n_774_ (
    .a(n_284_),
    .b(n_319_),
    .c(n_320_)
  );
  or_bb n_775_ (
    .a(n_320_),
    .b(n_318_),
    .c(n_322_)
  );
  and_ii n_776_ (
    .a(n_322_),
    .b(n_317_),
    .c(n_323_)
  );
  and_bb n_777_ (
    .a(n_322_),
    .b(n_317_),
    .c(n_324_)
  );
  or_bb n_778_ (
    .a(n_324_),
    .b(n_323_),
    .c(n_325_)
  );
  or_bb n_779_ (
    .a(n_325_),
    .b(n_283_),
    .c(n_326_)
  );
  and_bb n_780_ (
    .a(n_325_),
    .b(n_283_),
    .c(n_327_)
  );
  or_bi n_781_ (
    .a(n_327_),
    .b(n_326_),
    .c(n_328_)
  );
  and_ii n_782_ (
    .a(n_328_),
    .b(n_298_),
    .c(n_329_)
  );
  and_bb n_783_ (
    .a(n_328_),
    .b(n_298_),
    .c(n_330_)
  );
  or_bb n_784_ (
    .a(n_330_),
    .b(n_329_),
    .c(n_331_)
  );
  and_ii n_785_ (
    .a(n_331_),
    .b(n_316_),
    .c(n_333_)
  );
  and_bb n_786_ (
    .a(n_331_),
    .b(n_316_),
    .c(n_334_)
  );
  or_bb n_787_ (
    .a(n_334_),
    .b(n_333_),
    .c(n_335_)
  );
  and_ii n_788_ (
    .a(n_335_),
    .b(n_315_),
    .c(n_336_)
  );
  and_bb n_789_ (
    .a(n_335_),
    .b(n_315_),
    .c(n_337_)
  );
  or_bb n_790_ (
    .a(n_337_),
    .b(n_336_),
    .c(n_338_)
  );
  and_ii n_791_ (
    .a(n_338_),
    .b(n_314_),
    .c(n_339_)
  );
  and_bb n_792_ (
    .a(n_338_),
    .b(n_314_),
    .c(n_340_)
  );
  and_ii n_793_ (
    .a(n_340_),
    .b(n_339_),
    .c(s_12_)
  );
  and_ii n_794_ (
    .a(n_339_),
    .b(n_336_),
    .c(n_341_)
  );
  and_ii n_795_ (
    .a(n_333_),
    .b(n_329_),
    .c(n_342_)
  );
  and_ii n_796_ (
    .a(n_323_),
    .b(n_318_),
    .c(n_343_)
  );
  or_ii n_797_ (
    .a(b_7_),
    .b(a_7_),
    .c(n_344_)
  );
  and_bi n_798_ (
    .a(n_319_),
    .b(n_344_),
    .c(n_345_)
  );
  or_ii n_799_ (
    .a(b_6_),
    .b(a_7_),
    .c(n_346_)
  );
  and_bb n_800_ (
    .a(b_7_),
    .b(a_6_),
    .c(n_347_)
  );
  and_bi n_801_ (
    .a(n_346_),
    .b(n_347_),
    .c(n_348_)
  );
  or_bb n_802_ (
    .a(n_348_),
    .b(n_345_),
    .c(n_349_)
  );
  and_ii n_803_ (
    .a(n_349_),
    .b(n_326_),
    .c(n_350_)
  );
  and_bb n_804_ (
    .a(n_349_),
    .b(n_326_),
    .c(n_351_)
  );
  or_bb n_805_ (
    .a(n_351_),
    .b(n_350_),
    .c(n_354_)
  );
  and_ii n_806_ (
    .a(n_354_),
    .b(n_343_),
    .c(n_355_)
  );
  and_bb n_807_ (
    .a(n_354_),
    .b(n_343_),
    .c(n_356_)
  );
  or_bb n_808_ (
    .a(n_356_),
    .b(n_355_),
    .c(n_357_)
  );
  and_ii n_809_ (
    .a(n_357_),
    .b(n_342_),
    .c(n_358_)
  );
  and_bb n_810_ (
    .a(n_357_),
    .b(n_342_),
    .c(n_359_)
  );
  or_bb n_811_ (
    .a(n_359_),
    .b(n_358_),
    .c(n_360_)
  );
  and_ii n_812_ (
    .a(n_360_),
    .b(n_341_),
    .c(n_361_)
  );
  and_bb n_813_ (
    .a(n_360_),
    .b(n_341_),
    .c(n_362_)
  );
  and_ii n_814_ (
    .a(n_362_),
    .b(n_361_),
    .c(s_13_)
  );
  and_ii n_815_ (
    .a(n_361_),
    .b(n_358_),
    .c(n_364_)
  );
  or_bb n_816_ (
    .a(n_344_),
    .b(n_319_),
    .c(n_365_)
  );
  and_ii n_817_ (
    .a(n_355_),
    .b(n_350_),
    .c(n_366_)
  );
  and_ii n_818_ (
    .a(n_366_),
    .b(n_365_),
    .c(n_367_)
  );
  and_bb n_819_ (
    .a(n_366_),
    .b(n_365_),
    .c(n_368_)
  );
  or_bb n_820_ (
    .a(n_368_),
    .b(n_367_),
    .c(n_369_)
  );
  and_ii n_821_ (
    .a(n_369_),
    .b(n_364_),
    .c(n_370_)
  );
  or_ii n_822_ (
    .a(n_369_),
    .b(n_364_),
    .c(n_371_)
  );
  and_bi n_823_ (
    .a(n_371_),
    .b(n_370_),
    .c(s_14_)
  );
  or_bb n_824_ (
    .a(n_367_),
    .b(n_345_),
    .c(n_372_)
  );
  or_bb n_825_ (
    .a(n_372_),
    .b(n_370_),
    .c(s_15_)
  );
  and_bb n_826_ (
    .a(b_0_),
    .b(a_0_),
    .c(s_0_)
  );
  or_ii n_827_ (
    .a(b_0_),
    .b(a_1_),
    .c(n_226_)
  );
  and_bb n_828_ (
    .a(b_1_),
    .b(a_0_),
    .c(n_236_)
  );
  or_bi n_829_ (
    .a(n_226_),
    .b(n_236_),
    .c(n_257_)
  );
  and_bi n_830_ (
    .a(n_226_),
    .b(n_236_),
    .c(n_258_)
  );
  and_bi n_831_ (
    .a(n_257_),
    .b(n_258_),
    .c(s_1_)
  );
  or_ii n_832_ (
    .a(b_2_),
    .b(a_0_),
    .c(n_278_)
  );
  or_ii n_833_ (
    .a(a_1_),
    .b(b_1_),
    .c(n_289_)
  );
  and_bb n_834_ (
    .a(b_0_),
    .b(a_2_),
    .c(n_300_)
  );
  and_bi n_835_ (
    .a(n_300_),
    .b(n_289_),
    .c(n_311_)
  );
  and_bi n_836_ (
    .a(n_289_),
    .b(n_300_),
    .c(n_321_)
  );
  or_bb n_837_ (
    .a(n_321_),
    .b(n_311_),
    .c(n_332_)
  );
  and_ii n_838_ (
    .a(n_332_),
    .b(n_278_),
    .c(n_352_)
  );
  and_bb n_839_ (
    .a(n_332_),
    .b(n_278_),
    .c(n_353_)
  );
  or_bb n_840_ (
    .a(n_353_),
    .b(n_352_),
    .c(n_363_)
  );
  or_bb n_841_ (
    .a(n_363_),
    .b(n_257_),
    .c(n_373_)
  );
  and_bb n_842_ (
    .a(n_363_),
    .b(n_257_),
    .c(n_374_)
  );
  and_bi n_843_ (
    .a(n_373_),
    .b(n_374_),
    .c(s_2_)
  );
  or_ii n_844_ (
    .a(b_3_),
    .b(a_0_),
    .c(n_375_)
  );
  and_ii n_845_ (
    .a(n_352_),
    .b(n_311_),
    .c(n_376_)
  );
  or_ii n_846_ (
    .a(b_2_),
    .b(a_1_),
    .c(n_377_)
  );
  or_ii n_847_ (
    .a(a_2_),
    .b(b_1_),
    .c(n_378_)
  );
  or_ii n_848_ (
    .a(b_0_),
    .b(a_3_),
    .c(n_379_)
  );
  or_bb n_849_ (
    .a(n_379_),
    .b(n_378_),
    .c(n_380_)
  );
  or_ii n_850_ (
    .a(n_379_),
    .b(n_378_),
    .c(n_381_)
  );
  or_ii n_851_ (
    .a(n_381_),
    .b(n_380_),
    .c(n_382_)
  );
  and_ii n_852_ (
    .a(n_382_),
    .b(n_377_),
    .c(n_383_)
  );
  and_bb n_853_ (
    .a(n_382_),
    .b(n_377_),
    .c(n_384_)
  );
  or_bb n_854_ (
    .a(n_384_),
    .b(n_383_),
    .c(n_385_)
  );
  and_ii n_855_ (
    .a(n_385_),
    .b(n_376_),
    .c(n_386_)
  );
  and_bb n_856_ (
    .a(n_385_),
    .b(n_376_),
    .c(n_387_)
  );
  or_bb n_857_ (
    .a(n_387_),
    .b(n_386_),
    .c(n_388_)
  );
  and_ii n_858_ (
    .a(n_388_),
    .b(n_375_),
    .c(n_389_)
  );
  and_bb n_859_ (
    .a(n_388_),
    .b(n_375_),
    .c(n_390_)
  );
  or_bb n_860_ (
    .a(n_390_),
    .b(n_389_),
    .c(n_391_)
  );
  or_bb n_861_ (
    .a(n_391_),
    .b(n_373_),
    .c(n_392_)
  );
endmodule
