module c880(N259,N268,N153,N42,N201,N255,N207,N72,N183,N75,N267,N146,N111,N101,N177,N195,N171,N59,N106,N126,N8,N96,N17,N260,N1,N143,N165,N261,N86,N91,N36,N246,N189,N219,N228,N138,N13,N90,N156,N88,N51,N149,N74,N152,N210,N135,N237,N29,N85,N89,N116,N80,N73,N130,N87,N68,N121,N55,N159,N26);
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_181;
    wire _245_;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_1118;
    wire _015_;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_1487;
    wire _216_;
    wire _279_;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_106;
    wire _143_;
    wire new_Jinkela_wire_1987;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_1870;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_1843;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_1884;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_1620;
    wire _149_;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_1763;
    wire new_Jinkela_wire_0;
    wire _025_;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_1349;
    wire _238_;
    wire new_Jinkela_wire_1137;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_1396;
    wire _127_;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_1855;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_1195;
    wire _126_;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_619;
    wire _260_;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_877;
    wire _145_;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_1657;
    wire new_net_566;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_1156;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_628;
    wire new_net_530;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_1874;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_1691;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_1742;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_1853;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_1516;
    wire _178_;
    wire new_Jinkela_wire_1145;
    wire _205_;
    wire new_Jinkela_wire_1245;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_2030;
    wire _165_;
    wire _168_;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_2028;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_1748;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_914;
    wire _161_;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_1955;
    wire new_Jinkela_wire_1655;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_1929;
    wire _072_;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_1209;
    wire _241_;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_263;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_623;
    wire _019_;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_1185;
    wire _244_;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_601;
    wire _235_;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_1675;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_1883;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_208;
    wire _247_;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_1818;
    wire _105_;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_878;
    wire _000_;
    wire _185_;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_1820;
    wire _259_;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_2016;
    wire new_Jinkela_wire_2044;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_1315;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_1630;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_1123;
    wire _024_;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_1978;
    wire _049_;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_1682;
    wire _256_;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_1797;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_1688;
    wire _009_;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_483;
    wire _200_;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_1567;
    wire _286_;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_477;
    wire _179_;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_1262;
    wire _041_;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_1749;
    wire _199_;
    wire new_net_522;
    wire new_Jinkela_wire_1066;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_1510;
    wire _104_;
    wire new_Jinkela_wire_930;
    wire _232_;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_837;
    wire _064_;
    wire new_Jinkela_wire_1486;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_1832;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_1771;
    wire _036_;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_1437;
    wire _192_;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_1893;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_771;
    wire _092_;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_1862;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_1809;
    wire new_Jinkela_wire_2027;
    wire new_Jinkela_wire_2037;
    wire new_Jinkela_wire_363;
    wire _027_;
    wire _196_;
    wire _096_;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_1750;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_1705;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_1595;
    wire _140_;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_1800;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_151;
    wire new_net_552;
    wire _124_;
    wire new_Jinkela_wire_2014;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_121;
    wire _119_;
    wire new_Jinkela_wire_516;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_1856;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_1900;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_1866;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_918;
    wire _128_;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_1702;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_339;
    wire _176_;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_1252;
    wire new_Jinkela_wire_1852;
    wire _187_;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_310;
    wire _086_;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_115;
    wire _089_;
    wire _135_;
    wire new_Jinkela_wire_1755;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_1734;
    wire _226_;
    wire new_Jinkela_wire_1785;
    wire _280_;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_1945;
    wire new_Jinkela_wire_1618;
    wire _162_;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_1867;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_1989;
    wire _074_;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_1828;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_866;
    wire _172_;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_852;
    wire _188_;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_158;
    wire _035_;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_408;
    wire _110_;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_1745;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_1114;
    wire new_Jinkela_wire_1975;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_1757;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_1871;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_1726;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_1284;
    wire _284_;
    wire new_Jinkela_wire_1787;
    wire _103_;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_828;
    wire _102_;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_1404;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_1672;
    wire _222_;
    wire _047_;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_903;
    wire _234_;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_1689;
    wire new_Jinkela_wire_1713;
    wire _252_;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_1661;
    wire _182_;
    wire new_Jinkela_wire_198;
    wire _050_;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_1212;
    wire _177_;
    wire new_Jinkela_wire_1819;
    wire _203_;
    wire _156_;
    wire new_Jinkela_wire_1451;
    wire _084_;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_1403;
    wire _045_;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_1720;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_1990;
    wire _228_;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_690;
    wire _159_;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_1273;
    wire _087_;
    wire _148_;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_1807;
    wire _189_;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_1847;
    wire _249_;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_1415;
    wire _275_;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_307;
    wire _266_;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_248;
    wire _268_;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_800;
    wire _012_;
    wire _031_;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_1391;
    wire _173_;
    wire new_Jinkela_wire_1372;
    wire _056_;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_86;
    wire _032_;
    wire new_Jinkela_wire_698;
    wire _052_;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_1776;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_1627;
    wire _278_;
    wire new_Jinkela_wire_582;
    wire _229_;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_1359;
    wire _276_;
    wire _061_;
    wire new_Jinkela_wire_1132;
    wire _026_;
    wire new_net_558;
    wire new_Jinkela_wire_1991;
    wire _131_;
    wire _195_;
    wire new_Jinkela_wire_411;
    wire _230_;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_1450;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_1057;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_1140;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_2039;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_1761;
    wire new_Jinkela_wire_280;
    wire _186_;
    wire new_Jinkela_wire_1747;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_1134;
    wire _242_;
    wire new_Jinkela_wire_1258;
    wire new_Jinkela_wire_536;
    wire new_net_548;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_441;
    wire _018_;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_1904;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_1685;
    wire _236_;
    wire new_Jinkela_wire_1015;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_1583;
    wire new_Jinkela_wire_2015;
    wire _267_;
    wire new_Jinkela_wire_1358;
    wire _121_;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_1782;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_1110;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_925;
    wire _057_;
    wire _101_;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_1038;
    wire _270_;
    wire _251_;
    wire _022_;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_1848;
    wire new_Jinkela_wire_178;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_74;
    wire _014_;
    wire _184_;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_1371;
    wire _151_;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_325;
    wire _043_;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_1759;
    wire new_Jinkela_wire_189;
    wire _060_;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_1882;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_1764;
    wire _243_;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_1995;
    wire new_Jinkela_wire_1309;
    wire new_Jinkela_wire_279;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_1746;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_1668;
    wire _214_;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_1530;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_1407;
    wire _261_;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_1005;
    wire _034_;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_377;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_1972;
    wire new_Jinkela_wire_1997;
    wire new_Jinkela_wire_1268;
    wire _091_;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_1786;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_1326;
    wire _144_;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_1917;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_1203;
    wire _217_;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_1078;
    wire _277_;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_314;
    wire _138_;
    wire _254_;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_1073;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_1934;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_1915;
    wire new_net_534;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_274;
    wire _150_;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_1888;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_1963;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_713;
    wire _093_;
    wire new_Jinkela_wire_1804;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_1428;
    wire new_net_528;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_1398;
    wire _125_;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_1089;
    wire new_Jinkela_wire_1272;
    wire _158_;
    wire _106_;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_1846;
    wire new_Jinkela_wire_1872;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_1234;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_1777;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_1773;
    wire _046_;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_1833;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_845;
    wire new_net_0;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_1266;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_1131;
    wire _077_;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_2004;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_1485;
    wire _263_;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_2;
    wire _130_;
    wire _273_;
    wire _044_;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_1094;
    wire _274_;
    wire new_Jinkela_wire_1723;
    wire _210_;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_1724;
    wire new_Jinkela_wire_1817;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_681;
    wire _154_;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_993;
    wire _122_;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_1823;
    wire new_Jinkela_wire_1088;
    wire _083_;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_850;
    wire _227_;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_1160;
    wire _197_;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_1865;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_1652;
    wire _109_;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_236;
    wire new_net_524;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_1939;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_1406;
    wire _117_;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_14;
    wire _166_;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_1656;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_23;
    wire _271_;
    wire new_Jinkela_wire_1721;
    wire _272_;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_1984;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_1617;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_1106;
    wire _118_;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_1055;
    wire new_Jinkela_wire_598;
    wire _193_;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_1908;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_608;
    wire _194_;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_1722;
    wire _212_;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_1408;
    wire _066_;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_2001;
    wire _097_;
    wire _153_;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_895;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_1133;
    wire new_net_550;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_1141;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_921;
    wire _008_;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_1553;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_1333;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_1036;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_372;
    wire new_Jinkela_wire_737;
    wire _099_;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_407;
    wire _183_;
    wire new_Jinkela_wire_2012;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_1612;
    wire new_Jinkela_wire_589;
    wire _257_;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_1947;
    wire new_net_538;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_1741;
    wire _170_;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_1300;
    wire _003_;
    wire new_Jinkela_wire_12;
    wire _269_;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_395;
    wire _011_;
    wire new_net_520;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_1869;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_1421;
    wire _062_;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_592;
    wire new_net_554;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_39;
    wire _042_;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_1197;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_1948;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_1993;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_1285;
    wire _258_;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_1806;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_1949;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_1967;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_901;
    wire new_net_556;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_1951;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_1671;
    wire new_Jinkela_wire_760;
    wire new_net_532;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_1815;
    wire _213_;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_728;
    wire _081_;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_232;
    wire _111_;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_1844;
    wire _023_;
    wire _094_;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_1164;
    wire _146_;
    wire _082_;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_340;
    wire _223_;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_1009;
    wire _239_;
    wire _134_;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_1954;
    wire _157_;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_816;
    wire _147_;
    wire _007_;
    wire _171_;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_739;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_1857;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_1889;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_1037;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_1916;
    wire _113_;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_1829;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_1861;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_1420;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_1728;
    wire _071_;
    wire new_Jinkela_wire_1439;
    wire _255_;
    wire new_Jinkela_wire_2035;
    wire _224_;
    wire new_Jinkela_wire_385;
    wire _209_;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_56;
    wire new_Jinkela_wire_1751;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_145;
    wire new_net_540;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_1880;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_1163;
    wire _240_;
    wire _029_;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_1788;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_1802;
    wire new_Jinkela_wire_1943;
    wire _174_;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_547;
    wire _198_;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_1792;
    wire _208_;
    wire new_Jinkela_wire_1224;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_1666;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_79;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_1737;
    wire new_Jinkela_wire_1202;
    wire _112_;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_1715;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_1966;
    wire new_Jinkela_wire_1941;
    wire new_Jinkela_wire_1374;
    wire _075_;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_532;
    wire _069_;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_1924;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_2018;
    wire new_Jinkela_wire_624;
    wire _065_;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_119;
    wire _181_;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_1074;
    wire _078_;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_1781;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_1918;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_335;
    wire _265_;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_1753;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_2033;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_1646;
    wire _090_;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_1911;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_1765;
    wire _163_;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_1135;
    wire _053_;
    wire new_Jinkela_wire_2043;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_1192;
    wire _017_;
    wire _264_;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_1725;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_499;
    wire _129_;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_1860;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_1740;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_1240;
    wire new_net_546;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_1340;
    wire _004_;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_1897;
    wire _040_;
    wire new_Jinkela_wire_1950;
    wire new_Jinkela_wire_1549;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_1479;
    wire _285_;
    wire _028_;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_987;
    wire _002_;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_1779;
    wire _282_;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_150;
    wire _037_;
    wire new_Jinkela_wire_1931;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_1906;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_1913;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_1016;
    wire new_Jinkela_wire_1647;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_1151;
    wire new_Jinkela_wire_1892;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_1775;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_714;
    wire _108_;
    wire _048_;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_571;
    wire _107_;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_1286;
    wire _152_;
    wire new_Jinkela_wire_1962;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_1475;
    wire new_Jinkela_wire_1816;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_1719;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_1878;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_1953;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_2013;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_403;
    wire _207_;
    wire _225_;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_272;
    wire _115_;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_61;
    wire _169_;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_2034;
    wire new_Jinkela_wire_1248;
    wire new_net_564;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_2005;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_1886;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_1754;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_1994;
    wire new_Jinkela_wire_204;
    wire _016_;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_813;
    wire _218_;
    wire new_Jinkela_wire_755;
    wire _133_;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_1693;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_1178;
    wire _051_;
    wire new_Jinkela_wire_1351;
    wire _039_;
    wire _202_;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_1445;
    wire _204_;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_64;
    wire new_net_542;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_1979;
    wire new_Jinkela_wire_1004;
    wire _262_;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_233;
    wire _076_;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_1854;
    wire _160_;
    wire new_Jinkela_wire_1717;
    wire new_Jinkela_wire_847;
    wire _068_;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_1729;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_1985;
    wire _013_;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_1698;
    wire _246_;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_1086;
    wire new_Jinkela_wire_2002;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_1895;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_1584;
    wire _010_;
    wire new_Jinkela_wire_431;
    wire _211_;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_1261;
    wire _006_;
    wire _175_;
    wire _020_;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_1334;
    wire _001_;
    wire _070_;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_1780;
    wire _038_;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_1921;
    wire _088_;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_1712;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_1930;
    wire _067_;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_1436;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_1076;
    wire _059_;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_1907;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_1803;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_430;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_1935;
    wire new_Jinkela_wire_1977;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_1591;
    wire _142_;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_1113;
    wire _073_;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_122;
    wire _283_;
    wire _281_;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_1063;
    wire new_Jinkela_wire_1840;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_1957;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_1093;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_1643;
    wire new_Jinkela_wire_480;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_1294;
    wire _190_;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_1973;
    wire _021_;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_1626;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_1007;
    wire _136_;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_1801;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_161;
    wire _201_;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_1996;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_93;
    wire _123_;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_1942;
    wire new_Jinkela_wire_1739;
    wire _055_;
    wire new_Jinkela_wire_814;
    wire new_net_536;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_1201;
    wire new_net_560;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_482;
    wire new_net_544;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_2009;
    wire new_Jinkela_wire_1960;
    wire new_net_562;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_249;
    wire _120_;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_2017;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_1097;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_1899;
    wire new_Jinkela_wire_1514;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_964;
    wire _164_;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_173;
    wire _030_;
    wire new_Jinkela_wire_104;
    wire _220_;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_2046;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_120;
    wire new_net_526;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_1506;
    wire _233_;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_1971;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_1744;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_767;
    wire _248_;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_2003;
    wire _139_;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_1040;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_22;
    wire _063_;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_40;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_999;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_2010;
    wire _215_;
    wire new_Jinkela_wire_2038;
    wire new_Jinkela_wire_370;
    wire _085_;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_1767;
    wire _033_;
    wire new_Jinkela_wire_1166;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_1090;
    wire _221_;
    wire new_Jinkela_wire_1822;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_1727;
    wire _132_;
    wire new_Jinkela_wire_1241;
    wire _095_;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_1405;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_835;
    wire _100_;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_1482;
    wire _250_;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_1896;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_981;
    wire _253_;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_1774;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_1697;
    wire _219_;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_254;
    wire _167_;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_1743;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_2045;
    wire _114_;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_1881;
    wire new_Jinkela_wire_1677;
    wire _141_;
    wire _054_;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_1938;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_1859;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_1503;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_1709;
    wire _058_;
    wire _116_;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_304;
    wire _206_;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_241;
    wire _079_;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_1687;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_505;
    wire _005_;
    wire new_Jinkela_wire_1028;
    wire _080_;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_364;
    wire _098_;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_268;
    wire _191_;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_180;
    wire _180_;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_2025;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_928;
    wire _137_;
    wire new_Jinkela_wire_1096;
    wire _237_;
    wire new_Jinkela_wire_661;
    wire _231_;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_1969;
    wire new_Jinkela_wire_365;
    wire _155_;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_1354;
    input N259;
    input N268;
    input N153;
    input N42;
    input N201;
    input N255;
    input N207;
    input N72;
    input N183;
    input N75;
    input N267;
    input N146;
    input N111;
    input N101;
    input N177;
    input N195;
    input N171;
    input N59;
    input N106;
    input N126;
    input N8;
    input N96;
    input N17;
    input N260;
    input N1;
    input N143;
    input N165;
    input N261;
    input N86;
    input N91;
    input N36;
    input N246;
    input N189;
    input N219;
    input N228;
    input N138;
    input N13;
    input N90;
    input N156;
    input N88;
    input N51;
    input N149;
    input N74;
    input N152;
    input N210;
    input N135;
    input N237;
    input N29;
    input N85;
    input N89;
    input N116;
    input N80;
    input N73;
    input N130;
    input N87;
    input N68;
    input N121;
    input N55;
    input N159;
    input N26;
    output N419;
    output N447;
    output N448;
    output N866;
    output N389;
    output N446;
    output N449;
    output N418;
    output N768;
    output N420;
    output N874;
    output N421;
    output N880;
    output N390;
    output N865;
    output N767;
    output N450;
    output N391;
    output N863;
    output N878;
    output N422;
    output N864;
    output N879;
    output N423;
    output N388;
    output N850;

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_1446),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_1470),
        .dout(new_Jinkela_wire_1471)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(new_Jinkela_wire_1447),
        .dout(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_1471),
        .dout(new_Jinkela_wire_1472)
    );

    spl2 new_Jinkela_splitter_142 (
        .a(new_Jinkela_wire_1448),
        .b(new_Jinkela_wire_1449),
        .c(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_1450),
        .dout(new_Jinkela_wire_1451)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(_255_),
        .b(new_Jinkela_wire_1500),
        .c(new_Jinkela_wire_1501)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_1472),
        .dout(new_Jinkela_wire_1473)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_1451),
        .dout(new_Jinkela_wire_1452)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(_209_),
        .dout(new_Jinkela_wire_1502)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(new_Jinkela_wire_1493),
        .dout(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_1452),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_1473),
        .dout(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_1474),
        .dout(new_Jinkela_wire_1475)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_1502),
        .dout(new_Jinkela_wire_1503)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_1494),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_1475),
        .dout(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_1495),
        .dout(new_Jinkela_wire_1496)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(new_net_540),
        .dout(new_Jinkela_wire_1507)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(new_Jinkela_wire_1496),
        .dout(new_Jinkela_wire_1497)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(_029_),
        .b(new_Jinkela_wire_1543),
        .c(new_Jinkela_wire_1544)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(_198_),
        .b(new_Jinkela_wire_1553),
        .c(new_Jinkela_wire_1554)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_Jinkela_wire_1497),
        .dout(new_Jinkela_wire_1498)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_1503),
        .dout(new_Jinkela_wire_1504)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_1504),
        .dout(new_Jinkela_wire_1505)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(new_Jinkela_wire_1544),
        .dout(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(new_Jinkela_wire_1505),
        .dout(new_Jinkela_wire_1506)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(_075_),
        .dout(new_Jinkela_wire_1557)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    spl2 new_Jinkela_splitter_148 (
        .a(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_1555),
        .c(new_Jinkela_wire_1556)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_1545),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_1511),
        .dout(new_Jinkela_wire_1512)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(_181_),
        .dout(new_Jinkela_wire_1561)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_1512),
        .dout(new_Jinkela_wire_1513)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_1513),
        .dout(new_Jinkela_wire_1514)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(new_Jinkela_wire_1514),
        .dout(new_Jinkela_wire_1515)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(new_Jinkela_wire_1557),
        .dout(new_Jinkela_wire_1558)
    );

    spl2 new_Jinkela_splitter_133 (
        .a(new_Jinkela_wire_1195),
        .b(new_Jinkela_wire_1196),
        .c(new_Jinkela_wire_1197)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1163),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1203),
        .dout(new_Jinkela_wire_1204)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1164),
        .dout(new_Jinkela_wire_1165)
    );

    bfr new_Jinkela_buffer_873 (
        .din(_212_),
        .dout(new_Jinkela_wire_1212)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1165),
        .dout(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1207),
        .dout(new_Jinkela_wire_1208)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_1166),
        .dout(new_Jinkela_wire_1167)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1204),
        .dout(new_Jinkela_wire_1205)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1167),
        .dout(new_Jinkela_wire_1168)
    );

    bfr new_Jinkela_buffer_874 (
        .din(_066_),
        .dout(new_Jinkela_wire_1213)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1168),
        .dout(new_Jinkela_wire_1169)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1205),
        .dout(new_Jinkela_wire_1206)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_1169),
        .dout(new_Jinkela_wire_1170)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1208),
        .dout(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1170),
        .dout(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_net_550),
        .dout(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_1171),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1209),
        .dout(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_1172),
        .dout(new_Jinkela_wire_1173)
    );

    spl3L new_Jinkela_splitter_136 (
        .a(_008_),
        .b(new_Jinkela_wire_1249),
        .c(new_Jinkela_wire_1250),
        .d(new_Jinkela_wire_1251)
    );

    bfr new_Jinkela_buffer_910 (
        .din(_183_),
        .dout(new_Jinkela_wire_1252)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1173),
        .dout(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_872 (
        .din(new_Jinkela_wire_1210),
        .dout(new_Jinkela_wire_1211)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1174),
        .dout(new_Jinkela_wire_1175)
    );

    bfr new_Jinkela_buffer_876 (
        .din(new_Jinkela_wire_1214),
        .dout(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1175),
        .dout(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_net_538),
        .dout(new_Jinkela_wire_1253)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1176),
        .dout(new_Jinkela_wire_1177)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1215),
        .dout(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1177),
        .dout(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_net_520),
        .dout(new_Jinkela_wire_1293)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1178),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_1179),
        .dout(new_Jinkela_wire_1180)
    );

    spl2 new_Jinkela_splitter_137 (
        .a(_011_),
        .b(new_Jinkela_wire_1291),
        .c(new_Jinkela_wire_1292)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1217),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1181),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1253),
        .dout(new_Jinkela_wire_1254)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1182),
        .dout(new_Jinkela_wire_1183)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1218),
        .dout(new_Jinkela_wire_1219)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1183),
        .dout(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    spl3L new_Jinkela_splitter_110 (
        .a(_182_),
        .b(new_Jinkela_wire_830),
        .c(new_Jinkela_wire_831),
        .d(new_Jinkela_wire_832)
    );

    spl3L new_Jinkela_splitter_111 (
        .a(_084_),
        .b(new_Jinkela_wire_838),
        .c(new_Jinkela_wire_839),
        .d(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(_087_),
        .b(new_Jinkela_wire_841),
        .c(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_555 (
        .din(_177_),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    bfr new_Jinkela_buffer_579 (
        .din(_148_),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_803),
        .dout(new_Jinkela_wire_804)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    bfr new_Jinkela_buffer_583 (
        .din(_249_),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_835),
        .dout(new_Jinkela_wire_836)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_836),
        .dout(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_842),
        .dout(new_Jinkela_wire_843)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    bfr new_Jinkela_buffer_586 (
        .din(_012_),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_843),
        .dout(new_Jinkela_wire_844)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_821),
        .dout(new_Jinkela_wire_822)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_822),
        .dout(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_844),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_2001),
        .dout(new_Jinkela_wire_2002)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_1979),
        .dout(new_Jinkela_wire_1980)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_Jinkela_wire_2023),
        .dout(new_Jinkela_wire_2024)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_1980),
        .dout(new_Jinkela_wire_1981)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_2002),
        .dout(new_Jinkela_wire_2003)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(new_Jinkela_wire_1981),
        .dout(new_Jinkela_wire_1982)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(_137_),
        .dout(new_Jinkela_wire_2030)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(new_Jinkela_wire_1982),
        .dout(new_Jinkela_wire_1983)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_2003),
        .dout(new_Jinkela_wire_2004)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(new_Jinkela_wire_1983),
        .dout(new_Jinkela_wire_1984)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(new_Jinkela_wire_2024),
        .dout(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(new_Jinkela_wire_1984),
        .dout(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_2004),
        .dout(new_Jinkela_wire_2005)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_1985),
        .dout(new_Jinkela_wire_1986)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_Jinkela_wire_1986),
        .dout(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_2005),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(new_Jinkela_wire_2025),
        .dout(new_Jinkela_wire_2026)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_2006),
        .dout(new_Jinkela_wire_2007)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_2030),
        .dout(new_Jinkela_wire_2031)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_2007),
        .dout(new_Jinkela_wire_2008)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(new_Jinkela_wire_2008),
        .dout(new_Jinkela_wire_2009)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(new_Jinkela_wire_2009),
        .dout(new_Jinkela_wire_2010)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(new_Jinkela_wire_2031),
        .dout(new_Jinkela_wire_2032)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_2010),
        .dout(new_Jinkela_wire_2011)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_2011),
        .dout(new_Jinkela_wire_2012)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_2032),
        .dout(new_Jinkela_wire_2033)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_2012),
        .dout(new_Jinkela_wire_2013)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(new_Jinkela_wire_2013),
        .dout(new_Jinkela_wire_2014)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_2033),
        .dout(new_Jinkela_wire_2034)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_2014),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(new_Jinkela_wire_2015),
        .dout(new_Jinkela_wire_2016)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(new_Jinkela_wire_2034),
        .dout(new_Jinkela_wire_2035)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_2016),
        .dout(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_Jinkela_wire_2035),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_158),
        .dout(new_Jinkela_wire_159)
    );

    or_bb _484_ (
        .a(new_Jinkela_wire_571),
        .b(_173_),
        .c(_179_)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_1759),
        .dout(new_Jinkela_wire_1760)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_196),
        .b(new_Jinkela_wire_197),
        .c(new_Jinkela_wire_198)
    );

    and_bi _334_ (
        .a(new_Jinkela_wire_337),
        .b(new_Jinkela_wire_1989),
        .c(_034_)
    );

    or_bb _485_ (
        .a(new_Jinkela_wire_630),
        .b(_172_),
        .c(_180_)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1184),
        .dout(new_Jinkela_wire_1185)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_159),
        .dout(new_Jinkela_wire_160)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(new_Jinkela_wire_1775),
        .dout(new_Jinkela_wire_1776)
    );

    or_bb _486_ (
        .a(new_Jinkela_wire_2029),
        .b(_171_),
        .c(_181_)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_1219),
        .dout(new_Jinkela_wire_1220)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_1760),
        .dout(new_Jinkela_wire_1761)
    );

    or_bb _487_ (
        .a(new_Jinkela_wire_1565),
        .b(_170_),
        .c(new_net_530)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1185),
        .dout(new_Jinkela_wire_1186)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(_120_),
        .dout(new_Jinkela_wire_1889)
    );

    spl2 new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_160),
        .b(new_Jinkela_wire_161),
        .c(new_Jinkela_wire_162)
    );

    and_ii _488_ (
        .a(new_Jinkela_wire_621),
        .b(new_Jinkela_wire_825),
        .c(_182_)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1254),
        .dout(new_Jinkela_wire_1255)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_1761),
        .dout(new_Jinkela_wire_1762)
    );

    or_ii _489_ (
        .a(new_Jinkela_wire_831),
        .b(new_Jinkela_wire_281),
        .c(_183_)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1186),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_1776),
        .dout(new_Jinkela_wire_1777)
    );

    spl3L new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_182),
        .b(new_Jinkela_wire_183),
        .c(new_Jinkela_wire_184),
        .d(new_Jinkela_wire_185)
    );

    and_bi _490_ (
        .a(new_Jinkela_wire_1678),
        .b(new_Jinkela_wire_832),
        .c(_184_)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_1762),
        .dout(new_Jinkela_wire_1763)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    or_bb _491_ (
        .a(_184_),
        .b(new_Jinkela_wire_1431),
        .c(_185_)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_176),
        .dout(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1187),
        .dout(new_Jinkela_wire_1188)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    and_bi _492_ (
        .a(new_Jinkela_wire_1252),
        .b(_185_),
        .c(_186_)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1293),
        .dout(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_1763),
        .dout(new_Jinkela_wire_1764)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    and_bb _493_ (
        .a(new_Jinkela_wire_830),
        .b(new_Jinkela_wire_391),
        .c(_187_)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1188),
        .dout(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_1777),
        .dout(new_Jinkela_wire_1778)
    );

    and_bi _494_ (
        .a(new_Jinkela_wire_623),
        .b(new_Jinkela_wire_1956),
        .c(_188_)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_1764),
        .dout(new_Jinkela_wire_1765)
    );

    and_bi _495_ (
        .a(new_Jinkela_wire_315),
        .b(new_Jinkela_wire_1090),
        .c(_189_)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_178),
        .dout(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1189),
        .dout(new_Jinkela_wire_1190)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_1834),
        .dout(new_Jinkela_wire_1835)
    );

    and_bi _496_ (
        .a(new_Jinkela_wire_40),
        .b(new_Jinkela_wire_592),
        .c(_190_)
    );

    spl4L new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_211),
        .b(new_Jinkela_wire_212),
        .c(new_Jinkela_wire_213),
        .d(new_Jinkela_wire_214),
        .e(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1255),
        .dout(new_Jinkela_wire_1256)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(new_Jinkela_wire_1778),
        .dout(new_Jinkela_wire_1779)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    and_bb _497_ (
        .a(new_Jinkela_wire_79),
        .b(new_Jinkela_wire_49),
        .c(_191_)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1222),
        .dout(new_Jinkela_wire_1223)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    and_bb _498_ (
        .a(new_Jinkela_wire_447),
        .b(new_Jinkela_wire_504),
        .c(_192_)
    );

    spl3L new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_207),
        .b(new_Jinkela_wire_208),
        .c(new_Jinkela_wire_209),
        .d(new_Jinkela_wire_210)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_net_554),
        .dout(new_Jinkela_wire_1322)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_1779),
        .dout(new_Jinkela_wire_1780)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    or_bb _499_ (
        .a(_192_),
        .b(new_Jinkela_wire_2028),
        .c(_193_)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1223),
        .dout(new_Jinkela_wire_1224)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(new_Jinkela_wire_1852),
        .dout(new_Jinkela_wire_1853)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_215),
        .dout(new_Jinkela_wire_216)
    );

    or_bb _500_ (
        .a(new_Jinkela_wire_1206),
        .b(_190_),
        .c(_194_)
    );

    spl3L new_Jinkela_splitter_36 (
        .a(N1),
        .b(new_Jinkela_wire_223),
        .c(new_Jinkela_wire_224),
        .d(new_Jinkela_wire_225)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1256),
        .dout(new_Jinkela_wire_1257)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_1780),
        .dout(new_Jinkela_wire_1781)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    or_bb _501_ (
        .a(new_Jinkela_wire_1211),
        .b(_189_),
        .c(_195_)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1224),
        .dout(new_Jinkela_wire_1225)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    or_bb _502_ (
        .a(new_Jinkela_wire_933),
        .b(_188_),
        .c(_196_)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_199),
        .dout(new_Jinkela_wire_200)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(_042_),
        .b(new_Jinkela_wire_1359),
        .c(new_Jinkela_wire_1360)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(_258_),
        .b(new_Jinkela_wire_1364),
        .c(new_Jinkela_wire_1365)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_1781),
        .dout(new_Jinkela_wire_1782)
    );

    or_bb _503_ (
        .a(new_Jinkela_wire_674),
        .b(_187_),
        .c(_197_)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1225),
        .dout(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    or_bb _504_ (
        .a(new_Jinkela_wire_1150),
        .b(_186_),
        .c(new_net_544)
    );

    bfr new_Jinkela_buffer_130 (
        .din(N260),
        .dout(new_Jinkela_wire_222)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1257),
        .dout(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_1782),
        .dout(new_Jinkela_wire_1783)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_190),
        .dout(new_Jinkela_wire_191)
    );

    and_bb _505_ (
        .a(new_Jinkela_wire_1359),
        .b(new_Jinkela_wire_632),
        .c(_198_)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1226),
        .dout(new_Jinkela_wire_1227)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_1810),
        .dout(new_Jinkela_wire_1811)
    );

    and_bi _506_ (
        .a(new_Jinkela_wire_1709),
        .b(new_Jinkela_wire_1556),
        .c(_199_)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1294),
        .dout(new_Jinkela_wire_1295)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    and_bi _507_ (
        .a(new_Jinkela_wire_1555),
        .b(new_Jinkela_wire_1707),
        .c(_200_)
    );

    spl3L new_Jinkela_splitter_38 (
        .a(N165),
        .b(new_Jinkela_wire_246),
        .c(new_Jinkela_wire_247),
        .d(new_Jinkela_wire_248)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_1227),
        .dout(new_Jinkela_wire_1228)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(_164_),
        .dout(new_Jinkela_wire_1893)
    );

    or_bb _508_ (
        .a(_200_),
        .b(_199_),
        .c(_201_)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1258),
        .dout(new_Jinkela_wire_1259)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    and_bi _509_ (
        .a(new_Jinkela_wire_360),
        .b(_201_),
        .c(_202_)
    );

    bfr new_Jinkela_buffer_139 (
        .din(N143),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1228),
        .dout(new_Jinkela_wire_1229)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_1811),
        .dout(new_Jinkela_wire_1812)
    );

    and_bb _510_ (
        .a(new_Jinkela_wire_1553),
        .b(new_Jinkela_wire_392),
        .c(_203_)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(new_Jinkela_wire_1785),
        .dout(new_Jinkela_wire_1786)
    );

    and_bi _511_ (
        .a(new_Jinkela_wire_467),
        .b(new_Jinkela_wire_631),
        .c(_204_)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1229),
        .dout(new_Jinkela_wire_1230)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    and_bi _512_ (
        .a(new_Jinkela_wire_317),
        .b(new_Jinkela_wire_1635),
        .c(_205_)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_203),
        .dout(new_Jinkela_wire_204)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1259),
        .dout(new_Jinkela_wire_1260)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_1786),
        .dout(new_Jinkela_wire_1787)
    );

    and_bi _513_ (
        .a(new_Jinkela_wire_145),
        .b(new_Jinkela_wire_588),
        .c(_206_)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1230),
        .dout(new_Jinkela_wire_1231)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_216),
        .dout(new_Jinkela_wire_217)
    );

    and_bb _514_ (
        .a(new_Jinkela_wire_222),
        .b(new_Jinkela_wire_51),
        .c(_207_)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_204),
        .dout(new_Jinkela_wire_205)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1295),
        .dout(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_1787),
        .dout(new_Jinkela_wire_1788)
    );

    and_bb _515_ (
        .a(new_Jinkela_wire_442),
        .b(new_Jinkela_wire_476),
        .c(_208_)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1231),
        .dout(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(new_Jinkela_wire_1853),
        .dout(new_Jinkela_wire_1854)
    );

    or_bb _516_ (
        .a(_208_),
        .b(new_Jinkela_wire_1691),
        .c(_209_)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_205),
        .dout(new_Jinkela_wire_206)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_1260),
        .dout(new_Jinkela_wire_1261)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(new_Jinkela_wire_1788),
        .dout(new_Jinkela_wire_1789)
    );

    or_bb _517_ (
        .a(new_Jinkela_wire_1506),
        .b(_206_),
        .c(_210_)
    );

    spl2 new_Jinkela_splitter_41 (
        .a(N261),
        .b(new_Jinkela_wire_263),
        .c(new_Jinkela_wire_264)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1232),
        .dout(new_Jinkela_wire_1233)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    or_bb _518_ (
        .a(new_Jinkela_wire_1148),
        .b(_205_),
        .c(_211_)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1360),
        .dout(new_Jinkela_wire_1361)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(new_Jinkela_wire_1789),
        .dout(new_Jinkela_wire_1790)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_226),
        .dout(new_Jinkela_wire_227)
    );

    or_bb _519_ (
        .a(new_Jinkela_wire_1729),
        .b(_204_),
        .c(_212_)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1233),
        .dout(new_Jinkela_wire_1234)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    or_bb _520_ (
        .a(new_Jinkela_wire_1212),
        .b(_203_),
        .c(_213_)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1261),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_1790),
        .dout(new_Jinkela_wire_1791)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    or_bb _521_ (
        .a(new_Jinkela_wire_1407),
        .b(_202_),
        .c(new_net_522)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1234),
        .dout(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_1814),
        .dout(new_Jinkela_wire_1815)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    and_ii _522_ (
        .a(new_Jinkela_wire_1151),
        .b(new_Jinkela_wire_762),
        .c(_214_)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1296),
        .dout(new_Jinkela_wire_1297)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_1791),
        .dout(new_Jinkela_wire_1792)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    or_bb _523_ (
        .a(_214_),
        .b(new_Jinkela_wire_1987),
        .c(new_net_566)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1235),
        .dout(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_1889),
        .dout(new_Jinkela_wire_1890)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    or_ii _524_ (
        .a(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_468),
        .c(_215_)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_1792),
        .dout(new_Jinkela_wire_1793)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    and_bi _525_ (
        .a(new_Jinkela_wire_1734),
        .b(new_Jinkela_wire_1961),
        .c(new_net_550)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_1236),
        .dout(new_Jinkela_wire_1237)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_1815),
        .dout(new_Jinkela_wire_1816)
    );

    and_bi _313_ (
        .a(new_Jinkela_wire_876),
        .b(new_Jinkela_wire_1292),
        .c(_013_)
    );

    spl3L new_Jinkela_splitter_69 (
        .a(N29),
        .b(new_Jinkela_wire_468),
        .c(new_Jinkela_wire_469),
        .d(new_Jinkela_wire_470)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_405),
        .dout(new_Jinkela_wire_406)
    );

    or_bb _314_ (
        .a(new_Jinkela_wire_1725),
        .b(new_Jinkela_wire_1498),
        .c(_014_)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_845),
        .dout(new_Jinkela_wire_846)
    );

    bfr new_Jinkela_buffer_292 (
        .din(N89),
        .dout(new_Jinkela_wire_471)
    );

    or_bb _315_ (
        .a(_014_),
        .b(_006_),
        .c(_015_)
    );

    spl4L new_Jinkela_splitter_115 (
        .a(_278_),
        .b(new_Jinkela_wire_877),
        .c(new_Jinkela_wire_878),
        .d(new_Jinkela_wire_879),
        .e(new_Jinkela_wire_880)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_433),
        .dout(new_Jinkela_wire_434)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    and_bi _316_ (
        .a(_003_),
        .b(_015_),
        .c(_016_)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_846),
        .dout(new_Jinkela_wire_847)
    );

    or_bi _317_ (
        .a(new_Jinkela_wire_134),
        .b(new_Jinkela_wire_1705),
        .c(_017_)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    spl3L new_Jinkela_splitter_70 (
        .a(N116),
        .b(new_Jinkela_wire_473),
        .c(new_Jinkela_wire_474),
        .d(new_Jinkela_wire_475)
    );

    and_bi _318_ (
        .a(new_Jinkela_wire_133),
        .b(new_Jinkela_wire_1706),
        .c(_018_)
    );

    spl2 new_Jinkela_splitter_72 (
        .a(N80),
        .b(new_Jinkela_wire_486),
        .c(new_Jinkela_wire_487)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_453),
        .dout(new_Jinkela_wire_454)
    );

    and_bi _319_ (
        .a(new_Jinkela_wire_1578),
        .b(new_Jinkela_wire_937),
        .c(_019_)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(_229_),
        .b(new_Jinkela_wire_881),
        .c(new_Jinkela_wire_882)
    );

    and_bi _320_ (
        .a(new_Jinkela_wire_521),
        .b(new_Jinkela_wire_1291),
        .c(_020_)
    );

    bfr new_Jinkela_buffer_304 (
        .din(N73),
        .dout(new_Jinkela_wire_490)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_454),
        .dout(new_Jinkela_wire_455)
    );

    and_bi _321_ (
        .a(_020_),
        .b(new_Jinkela_wire_10),
        .c(_021_)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    and_bi _322_ (
        .a(new_Jinkela_wire_104),
        .b(new_Jinkela_wire_1653),
        .c(_022_)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    and_bi _323_ (
        .a(new_Jinkela_wire_221),
        .b(new_Jinkela_wire_1634),
        .c(_023_)
    );

    and_bi _324_ (
        .a(new_Jinkela_wire_233),
        .b(_023_),
        .c(_024_)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    and_bi _325_ (
        .a(new_Jinkela_wire_245),
        .b(new_Jinkela_wire_620),
        .c(_025_)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(new_Jinkela_wire_870),
        .b(new_Jinkela_wire_871),
        .c(new_Jinkela_wire_872)
    );

    or_bb _326_ (
        .a(_025_),
        .b(new_Jinkela_wire_964),
        .c(_026_)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_475),
        .b(new_Jinkela_wire_476),
        .c(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    and_ii _327_ (
        .a(_026_),
        .b(new_Jinkela_wire_1743),
        .c(_027_)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    and_bi _328_ (
        .a(new_Jinkela_wire_76),
        .b(new_Jinkela_wire_672),
        .c(_028_)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    and_bi _329_ (
        .a(new_Jinkela_wire_671),
        .b(new_Jinkela_wire_75),
        .c(_029_)
    );

    bfr new_Jinkela_buffer_592 (
        .din(_061_),
        .dout(new_Jinkela_wire_885)
    );

    or_bi _330_ (
        .a(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_91),
        .c(_030_)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    and_bi _331_ (
        .a(new_Jinkela_wire_485),
        .b(new_Jinkela_wire_1656),
        .c(_031_)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    spl3L new_Jinkela_splitter_73 (
        .a(N130),
        .b(new_Jinkela_wire_492),
        .c(new_Jinkela_wire_493),
        .d(new_Jinkela_wire_494)
    );

    or_bb _332_ (
        .a(_031_),
        .b(new_Jinkela_wire_1740),
        .c(_032_)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_854),
        .dout(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    inv _336_ (
        .din(new_Jinkela_wire_137),
        .dout(_036_)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    spl2 new_Jinkela_splitter_75 (
        .a(N68),
        .b(new_Jinkela_wire_499),
        .c(new_Jinkela_wire_500)
    );

    or_bi _337_ (
        .a(new_Jinkela_wire_617),
        .b(new_Jinkela_wire_434),
        .c(_037_)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    and_bi _338_ (
        .a(new_Jinkela_wire_513),
        .b(new_Jinkela_wire_1657),
        .c(_038_)
    );

    bfr new_Jinkela_buffer_590 (
        .din(_276_),
        .dout(new_Jinkela_wire_883)
    );

    or_bb _339_ (
        .a(_038_),
        .b(new_Jinkela_wire_1739),
        .c(_039_)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_490),
        .dout(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    and_bi _340_ (
        .a(_037_),
        .b(_039_),
        .c(_040_)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_488),
        .dout(new_Jinkela_wire_489)
    );

    or_bb _341_ (
        .a(new_Jinkela_wire_1636),
        .b(new_Jinkela_wire_670),
        .c(_041_)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    or_ii _342_ (
        .a(new_Jinkela_wire_1637),
        .b(new_Jinkela_wire_669),
        .c(_042_)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_net_558),
        .dout(new_Jinkela_wire_895)
    );

    or_bi _343_ (
        .a(new_Jinkela_wire_619),
        .b(new_Jinkela_wire_22),
        .c(_043_)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    and_bi _344_ (
        .a(new_Jinkela_wire_191),
        .b(new_Jinkela_wire_1652),
        .c(_044_)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    or_bb _345_ (
        .a(_044_),
        .b(new_Jinkela_wire_1738),
        .c(_045_)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    and_bi _346_ (
        .a(_043_),
        .b(_045_),
        .c(_046_)
    );

    bfr new_Jinkela_buffer_640 (
        .din(_195_),
        .dout(new_Jinkela_wire_933)
    );

    and_bi _347_ (
        .a(new_Jinkela_wire_1089),
        .b(new_Jinkela_wire_48),
        .c(_047_)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    inv _348_ (
        .din(new_Jinkela_wire_263),
        .dout(_048_)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    spl3L new_Jinkela_splitter_76 (
        .a(N121),
        .b(new_Jinkela_wire_501),
        .c(new_Jinkela_wire_502),
        .d(new_Jinkela_wire_503)
    );

    and_bi _349_ (
        .a(new_Jinkela_wire_47),
        .b(new_Jinkela_wire_1088),
        .c(_049_)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(new_Jinkela_wire_861),
        .b(new_Jinkela_wire_862),
        .c(new_Jinkela_wire_863)
    );

    and_bi _350_ (
        .a(new_Jinkela_wire_1675),
        .b(new_Jinkela_wire_622),
        .c(_050_)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_887),
        .dout(new_Jinkela_wire_888)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_515),
        .dout(new_Jinkela_wire_516)
    );

    or_bb _351_ (
        .a(_050_),
        .b(new_Jinkela_wire_827),
        .c(_051_)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    and_bi _352_ (
        .a(new_Jinkela_wire_1363),
        .b(new_Jinkela_wire_1708),
        .c(_052_)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_494),
        .dout(new_Jinkela_wire_495)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_net_548),
        .dout(new_Jinkela_wire_934)
    );

    and_bi _353_ (
        .a(new_Jinkela_wire_637),
        .b(_052_),
        .c(_053_)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_483),
        .dout(new_Jinkela_wire_484)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_888),
        .dout(new_Jinkela_wire_889)
    );

    or_bi _354_ (
        .a(new_Jinkela_wire_1576),
        .b(new_Jinkela_wire_785),
        .c(_054_)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_495),
        .dout(new_Jinkela_wire_496)
    );

    and_bi _355_ (
        .a(_054_),
        .b(new_Jinkela_wire_991),
        .c(_055_)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_484),
        .dout(new_Jinkela_wire_485)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_889),
        .dout(new_Jinkela_wire_890)
    );

    or_bb _356_ (
        .a(new_Jinkela_wire_1767),
        .b(new_Jinkela_wire_1552),
        .c(_056_)
    );

    spl3L new_Jinkela_splitter_117 (
        .a(_018_),
        .b(new_Jinkela_wire_937),
        .c(new_Jinkela_wire_938),
        .d(new_Jinkela_wire_939)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(_267_),
        .b(new_Jinkela_wire_954),
        .c(new_Jinkela_wire_955)
    );

    and_bi _357_ (
        .a(_056_),
        .b(new_Jinkela_wire_1649),
        .c(_057_)
    );

    spl2 new_Jinkela_splitter_78 (
        .a(N55),
        .b(new_Jinkela_wire_514),
        .c(new_Jinkela_wire_515)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_Jinkela_wire_2036),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(new_Jinkela_wire_2041),
        .dout(new_Jinkela_wire_2042)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(new_Jinkela_wire_2042),
        .dout(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_2044),
        .dout(new_Jinkela_wire_2045)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_2046),
        .dout(new_Jinkela_wire_2047)
    );

    bfr new_Jinkela_buffer_1 (
        .din(N268),
        .dout(new_Jinkela_wire_1)
    );

    bfr new_Jinkela_buffer_0 (
        .din(N259),
        .dout(new_Jinkela_wire_0)
    );

    bfr new_Jinkela_buffer_8 (
        .din(N153),
        .dout(new_Jinkela_wire_11)
    );

    spl3L new_Jinkela_splitter_2 (
        .a(N42),
        .b(new_Jinkela_wire_23),
        .c(new_Jinkela_wire_24),
        .d(new_Jinkela_wire_25)
    );

    spl3L new_Jinkela_splitter_5 (
        .a(N201),
        .b(new_Jinkela_wire_31),
        .c(new_Jinkela_wire_32),
        .d(new_Jinkela_wire_33)
    );

    spl3L new_Jinkela_splitter_0 (
        .a(new_Jinkela_wire_1),
        .b(new_Jinkela_wire_2),
        .c(new_Jinkela_wire_3),
        .d(new_Jinkela_wire_4)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_4),
        .dout(new_Jinkela_wire_5)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_259 (
        .din(N90),
        .dout(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1323),
        .dout(new_Jinkela_wire_1324)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(new_Jinkela_wire_1515),
        .dout(new_Jinkela_wire_1516)
    );

    spl2 new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_328),
        .b(new_Jinkela_wire_329),
        .c(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1237),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_1516),
        .dout(new_Jinkela_wire_1517)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_341),
        .dout(new_Jinkela_wire_342)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1238),
        .dout(new_Jinkela_wire_1239)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1297),
        .dout(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(new_Jinkela_wire_1517),
        .dout(new_Jinkela_wire_1518)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_331),
        .dout(new_Jinkela_wire_332)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1239),
        .dout(new_Jinkela_wire_1240)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_342),
        .dout(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(_078_),
        .dout(new_Jinkela_wire_1566)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_1264),
        .dout(new_Jinkela_wire_1265)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_1518),
        .dout(new_Jinkela_wire_1519)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1240),
        .dout(new_Jinkela_wire_1241)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_1558),
        .dout(new_Jinkela_wire_1559)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_1549),
        .dout(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_1519),
        .dout(new_Jinkela_wire_1520)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1241),
        .dout(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_343),
        .dout(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1265),
        .dout(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(new_Jinkela_wire_1520),
        .dout(new_Jinkela_wire_1521)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1242),
        .dout(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1298),
        .dout(new_Jinkela_wire_1299)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_1521),
        .dout(new_Jinkela_wire_1522)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_335),
        .b(new_Jinkela_wire_336),
        .c(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1243),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_1266),
        .dout(new_Jinkela_wire_1267)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(new_Jinkela_wire_1522),
        .dout(new_Jinkela_wire_1523)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_1559),
        .dout(new_Jinkela_wire_1560)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(new_Jinkela_wire_1551),
        .dout(new_Jinkela_wire_1552)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_413),
        .dout(new_Jinkela_wire_414)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1324),
        .dout(new_Jinkela_wire_1325)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_1523),
        .dout(new_Jinkela_wire_1524)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_261 (
        .din(N156),
        .dout(new_Jinkela_wire_417)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1267),
        .dout(new_Jinkela_wire_1268)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_1524),
        .dout(new_Jinkela_wire_1525)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_1246),
        .dout(new_Jinkela_wire_1247)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(_090_),
        .dout(new_Jinkela_wire_1567)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1299),
        .dout(new_Jinkela_wire_1300)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    spl2 new_Jinkela_splitter_61 (
        .a(N51),
        .b(new_Jinkela_wire_418),
        .c(new_Jinkela_wire_419)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1247),
        .dout(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_348),
        .dout(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1268),
        .dout(new_Jinkela_wire_1269)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    bfr new_Jinkela_buffer_263 (
        .din(N149),
        .dout(new_Jinkela_wire_423)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_net_556),
        .dout(new_Jinkela_wire_1366)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(_163_),
        .dout(new_Jinkela_wire_1574)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1269),
        .dout(new_Jinkela_wire_1270)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(new_Jinkela_wire_1527),
        .dout(new_Jinkela_wire_1528)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1300),
        .dout(new_Jinkela_wire_1301)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_350),
        .dout(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1270),
        .dout(new_Jinkela_wire_1271)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(new_Jinkela_wire_1528),
        .dout(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1325),
        .dout(new_Jinkela_wire_1326)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_1567),
        .dout(new_Jinkela_wire_1568)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1271),
        .dout(new_Jinkela_wire_1272)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_1529),
        .dout(new_Jinkela_wire_1530)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1301),
        .dout(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_1564),
        .dout(new_Jinkela_wire_1565)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1272),
        .dout(new_Jinkela_wire_1273)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(new_Jinkela_wire_1530),
        .dout(new_Jinkela_wire_1531)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_419),
        .b(new_Jinkela_wire_420),
        .c(new_Jinkela_wire_421)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    spl3L new_Jinkela_splitter_149 (
        .a(_053_),
        .b(new_Jinkela_wire_1575),
        .c(new_Jinkela_wire_1576),
        .d(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1361),
        .dout(new_Jinkela_wire_1362)
    );

    spl2 new_Jinkela_splitter_150 (
        .a(_017_),
        .b(new_Jinkela_wire_1578),
        .c(new_Jinkela_wire_1579)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1273),
        .dout(new_Jinkela_wire_1274)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_1531),
        .dout(new_Jinkela_wire_1532)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1302),
        .dout(new_Jinkela_wire_1303)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_1568),
        .dout(new_Jinkela_wire_1569)
    );

    spl2 new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_354),
        .b(new_Jinkela_wire_355),
        .c(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1274),
        .dout(new_Jinkela_wire_1275)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(new_Jinkela_wire_1532),
        .dout(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1326),
        .dout(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_273 (
        .din(N74),
        .dout(new_Jinkela_wire_435)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1275),
        .dout(new_Jinkela_wire_1276)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_1533),
        .dout(new_Jinkela_wire_1534)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1303),
        .dout(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(new_Jinkela_wire_1569),
        .dout(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1276),
        .dout(new_Jinkela_wire_1277)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_421),
        .dout(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(new_net_532),
        .dout(new_Jinkela_wire_1400)
    );

    spl2 new_Jinkela_splitter_151 (
        .a(_264_),
        .b(new_Jinkela_wire_1593),
        .c(new_Jinkela_wire_1594)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1277),
        .dout(new_Jinkela_wire_1278)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1304),
        .dout(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(new_Jinkela_wire_1838),
        .dout(new_Jinkela_wire_1839)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(new_Jinkela_wire_1794),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_1795),
        .dout(new_Jinkela_wire_1796)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(new_Jinkela_wire_1854),
        .dout(new_Jinkela_wire_1855)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(new_Jinkela_wire_1796),
        .dout(new_Jinkela_wire_1797)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_1817),
        .dout(new_Jinkela_wire_1818)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(new_Jinkela_wire_1797),
        .dout(new_Jinkela_wire_1798)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_Jinkela_wire_1839),
        .dout(new_Jinkela_wire_1840)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(new_Jinkela_wire_1798),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_1818),
        .dout(new_Jinkela_wire_1819)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(_220_),
        .b(new_Jinkela_wire_1894),
        .c(new_Jinkela_wire_1895)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_net_526),
        .dout(new_Jinkela_wire_1896)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(new_Jinkela_wire_1819),
        .dout(new_Jinkela_wire_1820)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_1840),
        .dout(new_Jinkela_wire_1841)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(new_Jinkela_wire_1802),
        .dout(new_Jinkela_wire_1803)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_1820),
        .dout(new_Jinkela_wire_1821)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(new_Jinkela_wire_1855),
        .dout(new_Jinkela_wire_1856)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_1841),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_1822),
        .dout(new_Jinkela_wire_1823)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(new_Jinkela_wire_1890),
        .dout(new_Jinkela_wire_1891)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_1823),
        .dout(new_Jinkela_wire_1824)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_1842),
        .dout(new_Jinkela_wire_1843)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_1824),
        .dout(new_Jinkela_wire_1825)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(new_Jinkela_wire_1856),
        .dout(new_Jinkela_wire_1857)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_1843),
        .dout(new_Jinkela_wire_1844)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_1826),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_1844),
        .dout(new_Jinkela_wire_1845)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(new_Jinkela_wire_1857),
        .dout(new_Jinkela_wire_1858)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(new_Jinkela_wire_1845),
        .dout(new_Jinkela_wire_1846)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(new_Jinkela_wire_1830),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(new_Jinkela_wire_1891),
        .dout(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    spl2 new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_503),
        .b(new_Jinkela_wire_504),
        .c(new_Jinkela_wire_505)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_496),
        .b(new_Jinkela_wire_497),
        .c(new_Jinkela_wire_498)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_891),
        .dout(new_Jinkela_wire_892)
    );

    spl3L new_Jinkela_splitter_80 (
        .a(N159),
        .b(new_Jinkela_wire_523),
        .c(new_Jinkela_wire_524),
        .d(new_Jinkela_wire_525)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    spl2 new_Jinkela_splitter_83 (
        .a(_216_),
        .b(new_Jinkela_wire_541),
        .c(new_Jinkela_wire_542)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_525),
        .dout(new_Jinkela_wire_526)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_332 (
        .din(_279_),
        .dout(new_Jinkela_wire_543)
    );

    bfr new_Jinkela_buffer_658 (
        .din(_121_),
        .dout(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_644 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_526),
        .dout(new_Jinkela_wire_527)
    );

    spl3L new_Jinkela_splitter_120 (
        .a(_101_),
        .b(new_Jinkela_wire_960),
        .c(new_Jinkela_wire_961),
        .d(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_331 (
        .din(N26),
        .dout(new_Jinkela_wire_540)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    spl2 new_Jinkela_splitter_85 (
        .a(_238_),
        .b(new_Jinkela_wire_548),
        .c(new_Jinkela_wire_549)
    );

    or_bi _335_ (
        .a(new_Jinkela_wire_336),
        .b(new_Jinkela_wire_1990),
        .c(_035_)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_527),
        .dout(new_Jinkela_wire_528)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    spl3L new_Jinkela_splitter_119 (
        .a(_057_),
        .b(new_Jinkela_wire_957),
        .c(new_Jinkela_wire_958),
        .d(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_519),
        .dout(new_Jinkela_wire_520)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_659 (
        .din(_270_),
        .dout(new_Jinkela_wire_963)
    );

    spl2 new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_520),
        .b(new_Jinkela_wire_521),
        .c(new_Jinkela_wire_522)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_660 (
        .din(_022_),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_net_566),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_334 (
        .din(_149_),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    bfr new_Jinkela_buffer_661 (
        .din(_151_),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    spl2 new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_544),
        .b(new_Jinkela_wire_545),
        .c(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_530),
        .dout(new_Jinkela_wire_531)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_net_530),
        .dout(new_Jinkela_wire_552)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(_261_),
        .b(new_Jinkela_wire_980),
        .c(new_Jinkela_wire_981)
    );

    spl2 new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_531),
        .b(new_Jinkela_wire_532),
        .c(new_Jinkela_wire_533)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_352 (
        .din(_178_),
        .dout(new_Jinkela_wire_567)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_534),
        .dout(new_Jinkela_wire_535)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_535),
        .dout(new_Jinkela_wire_536)
    );

    spl3L new_Jinkela_splitter_122 (
        .a(_034_),
        .b(new_Jinkela_wire_982),
        .c(new_Jinkela_wire_983),
        .d(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_357 (
        .din(_165_),
        .dout(new_Jinkela_wire_572)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    spl2 new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_537),
        .b(new_Jinkela_wire_538),
        .c(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    bfr new_Jinkela_buffer_184 (
        .din(N246),
        .dout(new_Jinkela_wire_297)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_231),
        .dout(new_Jinkela_wire_232)
    );

    spl2 new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_282),
        .b(new_Jinkela_wire_283),
        .c(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_232),
        .dout(new_Jinkela_wire_233)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_237),
        .dout(new_Jinkela_wire_238)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_248),
        .dout(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_238),
        .dout(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_240),
        .dout(new_Jinkela_wire_241)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    spl2 new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_241),
        .b(new_Jinkela_wire_242),
        .c(new_Jinkela_wire_243)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    bfr new_Jinkela_buffer_176 (
        .din(N91),
        .dout(new_Jinkela_wire_282)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_251),
        .dout(new_Jinkela_wire_252)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_244),
        .dout(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_266),
        .dout(new_Jinkela_wire_267)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_253),
        .dout(new_Jinkela_wire_254)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(N36),
        .b(new_Jinkela_wire_295),
        .c(new_Jinkela_wire_296)
    );

    spl2 new_Jinkela_splitter_39 (
        .a(new_Jinkela_wire_254),
        .b(new_Jinkela_wire_255),
        .c(new_Jinkela_wire_256)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_256),
        .dout(new_Jinkela_wire_257)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_267),
        .dout(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_257),
        .dout(new_Jinkela_wire_258)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_268),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_258),
        .dout(new_Jinkela_wire_259)
    );

    spl3L new_Jinkela_splitter_48 (
        .a(N189),
        .b(new_Jinkela_wire_320),
        .c(new_Jinkela_wire_321),
        .d(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_259),
        .dout(new_Jinkela_wire_260)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    spl2 new_Jinkela_splitter_40 (
        .a(new_Jinkela_wire_260),
        .b(new_Jinkela_wire_261),
        .c(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_270),
        .dout(new_Jinkela_wire_271)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(N219),
        .b(new_Jinkela_wire_338),
        .c(new_Jinkela_wire_339)
    );

    spl3L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_285),
        .b(new_Jinkela_wire_286),
        .c(new_Jinkela_wire_287),
        .d(new_Jinkela_wire_288)
    );

    bfr new_Jinkela_buffer_231 (
        .din(N228),
        .dout(new_Jinkela_wire_371)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_271),
        .dout(new_Jinkela_wire_272)
    );

    or_ii _526_ (
        .a(new_Jinkela_wire_164),
        .b(new_Jinkela_wire_296),
        .c(_216_)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1278),
        .dout(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_1536),
        .dout(new_Jinkela_wire_1537)
    );

    or_bb _527_ (
        .a(new_Jinkela_wire_542),
        .b(new_Jinkela_wire_1660),
        .c(new_net_554)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1327),
        .dout(new_Jinkela_wire_1328)
    );

    or_bb _528_ (
        .a(new_Jinkela_wire_541),
        .b(new_Jinkela_wire_1249),
        .c(new_net_524)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1279),
        .dout(new_Jinkela_wire_1280)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_1537),
        .dout(new_Jinkela_wire_1538)
    );

    or_bb _529_ (
        .a(new_Jinkela_wire_1735),
        .b(new_Jinkela_wire_1251),
        .c(new_net_562)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1305),
        .dout(new_Jinkela_wire_1306)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(new_Jinkela_wire_1571),
        .dout(new_Jinkela_wire_1572)
    );

    or_ii _530_ (
        .a(new_Jinkela_wire_295),
        .b(new_Jinkela_wire_470),
        .c(_217_)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1280),
        .dout(new_Jinkela_wire_1281)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(new_Jinkela_wire_1538),
        .dout(new_Jinkela_wire_1539)
    );

    and_bi _531_ (
        .a(new_Jinkela_wire_30),
        .b(new_Jinkela_wire_993),
        .c(new_net_0)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1366),
        .dout(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_net_546),
        .dout(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1362),
        .dout(new_Jinkela_wire_1363)
    );

    or_bb _532_ (
        .a(new_Jinkela_wire_119),
        .b(new_Jinkela_wire_524),
        .c(_218_)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1281),
        .dout(new_Jinkela_wire_1282)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_1539),
        .dout(new_Jinkela_wire_1540)
    );

    and_bb _533_ (
        .a(new_Jinkela_wire_118),
        .b(new_Jinkela_wire_523),
        .c(_219_)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1306),
        .dout(new_Jinkela_wire_1307)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_1572),
        .dout(new_Jinkela_wire_1573)
    );

    and_bi _534_ (
        .a(_218_),
        .b(_219_),
        .c(_220_)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1282),
        .dout(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(new_Jinkela_wire_1540),
        .dout(new_Jinkela_wire_1541)
    );

    and_bi _535_ (
        .a(new_Jinkela_wire_498),
        .b(new_Jinkela_wire_1895),
        .c(_221_)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1328),
        .dout(new_Jinkela_wire_1329)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    and_bi _536_ (
        .a(new_Jinkela_wire_1894),
        .b(new_Jinkela_wire_497),
        .c(_222_)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1283),
        .dout(new_Jinkela_wire_1284)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_1541),
        .dout(new_Jinkela_wire_1542)
    );

    and_ii _537_ (
        .a(_222_),
        .b(_221_),
        .c(_223_)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1307),
        .dout(new_Jinkela_wire_1308)
    );

    spl3L new_Jinkela_splitter_153 (
        .a(_040_),
        .b(new_Jinkela_wire_1635),
        .c(new_Jinkela_wire_1636),
        .d(new_Jinkela_wire_1637)
    );

    and_ii _538_ (
        .a(new_Jinkela_wire_135),
        .b(new_Jinkela_wire_320),
        .c(_224_)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1284),
        .dout(new_Jinkela_wire_1285)
    );

    spl2 new_Jinkela_splitter_152 (
        .a(_004_),
        .b(new_Jinkela_wire_1632),
        .c(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    and_bb _539_ (
        .a(new_Jinkela_wire_136),
        .b(new_Jinkela_wire_321),
        .c(_225_)
    );

    and_ii _540_ (
        .a(_225_),
        .b(_224_),
        .c(_226_)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1285),
        .dout(new_Jinkela_wire_1286)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_1582),
        .dout(new_Jinkela_wire_1583)
    );

    and_bi _541_ (
        .a(new_Jinkela_wire_56),
        .b(new_Jinkela_wire_765),
        .c(_227_)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1308),
        .dout(new_Jinkela_wire_1309)
    );

    and_bi _542_ (
        .a(new_Jinkela_wire_764),
        .b(new_Jinkela_wire_55),
        .c(_228_)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1286),
        .dout(new_Jinkela_wire_1287)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_1583),
        .dout(new_Jinkela_wire_1584)
    );

    or_bb _543_ (
        .a(_228_),
        .b(_227_),
        .c(_229_)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1329),
        .dout(new_Jinkela_wire_1330)
    );

    or_bi _544_ (
        .a(new_Jinkela_wire_246),
        .b(new_Jinkela_wire_31),
        .c(_230_)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1287),
        .dout(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(new_Jinkela_wire_1584),
        .dout(new_Jinkela_wire_1585)
    );

    and_bi _545_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_32),
        .c(_231_)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1309),
        .dout(new_Jinkela_wire_1310)
    );

    and_bi _546_ (
        .a(_230_),
        .b(_231_),
        .c(_232_)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1288),
        .dout(new_Jinkela_wire_1289)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_Jinkela_wire_1585),
        .dout(new_Jinkela_wire_1586)
    );

    and_bi _547_ (
        .a(new_Jinkela_wire_146),
        .b(new_Jinkela_wire_59),
        .c(_233_)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(_213_),
        .dout(new_Jinkela_wire_1406)
    );

    and_bi _548_ (
        .a(new_Jinkela_wire_58),
        .b(new_Jinkela_wire_147),
        .c(_234_)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1289),
        .dout(new_Jinkela_wire_1290)
    );

    spl3L new_Jinkela_splitter_154 (
        .a(_028_),
        .b(new_Jinkela_wire_1638),
        .c(new_Jinkela_wire_1639),
        .d(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(new_Jinkela_wire_1586),
        .dout(new_Jinkela_wire_1587)
    );

    or_bb _549_ (
        .a(_234_),
        .b(_233_),
        .c(_235_)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1310),
        .dout(new_Jinkela_wire_1311)
    );

    and_ii _550_ (
        .a(new_Jinkela_wire_613),
        .b(new_Jinkela_wire_657),
        .c(_236_)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1330),
        .dout(new_Jinkela_wire_1331)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(new_Jinkela_wire_1587),
        .dout(new_Jinkela_wire_1588)
    );

    and_bb _551_ (
        .a(new_Jinkela_wire_612),
        .b(new_Jinkela_wire_656),
        .c(_237_)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1311),
        .dout(new_Jinkela_wire_1312)
    );

    and_ii _552_ (
        .a(_237_),
        .b(_236_),
        .c(_238_)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1367),
        .dout(new_Jinkela_wire_1368)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(new_Jinkela_wire_1588),
        .dout(new_Jinkela_wire_1589)
    );

    and_ii _553_ (
        .a(new_Jinkela_wire_549),
        .b(new_Jinkela_wire_882),
        .c(_239_)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1312),
        .dout(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(new_Jinkela_wire_1640),
        .dout(new_Jinkela_wire_1641)
    );

    and_bb _554_ (
        .a(new_Jinkela_wire_548),
        .b(new_Jinkela_wire_881),
        .c(_240_)
    );

    bfr new_Jinkela_buffer_988 (
        .din(new_Jinkela_wire_1331),
        .dout(new_Jinkela_wire_1332)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_Jinkela_wire_1589),
        .dout(new_Jinkela_wire_1590)
    );

    and_ii _555_ (
        .a(_240_),
        .b(_239_),
        .c(_241_)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1313),
        .dout(new_Jinkela_wire_1314)
    );

    and_bi _556_ (
        .a(new_Jinkela_wire_596),
        .b(new_Jinkela_wire_1487),
        .c(_242_)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1400),
        .dout(new_Jinkela_wire_1401)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_1590),
        .dout(new_Jinkela_wire_1591)
    );

    and_bi _557_ (
        .a(new_Jinkela_wire_1486),
        .b(new_Jinkela_wire_595),
        .c(_243_)
    );

    bfr new_Jinkela_buffer_971 (
        .din(new_Jinkela_wire_1314),
        .dout(new_Jinkela_wire_1315)
    );

    spl2 new_Jinkela_splitter_158 (
        .a(_282_),
        .b(new_Jinkela_wire_1660),
        .c(new_Jinkela_wire_1661)
    );

    or_bb _558_ (
        .a(_243_),
        .b(_242_),
        .c(new_net_560)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1332),
        .dout(new_Jinkela_wire_1333)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_1591),
        .dout(new_Jinkela_wire_1592)
    );

    and_ii _559_ (
        .a(new_Jinkela_wire_493),
        .b(new_Jinkela_wire_194),
        .c(_244_)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1315),
        .dout(new_Jinkela_wire_1316)
    );

    and_bb _560_ (
        .a(new_Jinkela_wire_492),
        .b(new_Jinkela_wire_195),
        .c(_245_)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1368),
        .dout(new_Jinkela_wire_1369)
    );

    spl2 new_Jinkela_splitter_155 (
        .a(_002_),
        .b(new_Jinkela_wire_1650),
        .c(new_Jinkela_wire_1655)
    );

    or_bb _561_ (
        .a(_245_),
        .b(_244_),
        .c(_246_)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1316),
        .dout(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(new_Jinkela_wire_1601),
        .dout(new_Jinkela_wire_1602)
    );

    and_bi _562_ (
        .a(new_Jinkela_wire_287),
        .b(new_Jinkela_wire_1727),
        .c(_247_)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1333),
        .dout(new_Jinkela_wire_1334)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_1641),
        .dout(new_Jinkela_wire_1642)
    );

    and_bi _563_ (
        .a(new_Jinkela_wire_1726),
        .b(new_Jinkela_wire_286),
        .c(_248_)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1317),
        .dout(new_Jinkela_wire_1318)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    and_ii _564_ (
        .a(_248_),
        .b(_247_),
        .c(_249_)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(_081_),
        .dout(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(_048_),
        .dout(new_Jinkela_wire_1662)
    );

    and_ii _565_ (
        .a(new_Jinkela_wire_450),
        .b(new_Jinkela_wire_501),
        .c(_250_)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1318),
        .dout(new_Jinkela_wire_1319)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    and_bb _566_ (
        .a(new_Jinkela_wire_449),
        .b(new_Jinkela_wire_502),
        .c(_251_)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1334),
        .dout(new_Jinkela_wire_1335)
    );

    spl4L new_Jinkela_splitter_157 (
        .a(new_Jinkela_wire_1655),
        .b(new_Jinkela_wire_1656),
        .c(new_Jinkela_wire_1657),
        .d(new_Jinkela_wire_1658),
        .e(new_Jinkela_wire_1659)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_1642),
        .dout(new_Jinkela_wire_1643)
    );

    and_ii _567_ (
        .a(_251_),
        .b(_250_),
        .c(_252_)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1319),
        .dout(new_Jinkela_wire_1320)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_359),
        .b(new_Jinkela_wire_360),
        .c(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_276 (
        .din(N152),
        .dout(new_Jinkela_wire_438)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_381),
        .dout(new_Jinkela_wire_382)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_423),
        .dout(new_Jinkela_wire_424)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_948),
        .dout(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    spl2 new_Jinkela_splitter_54 (
        .a(new_Jinkela_wire_363),
        .b(new_Jinkela_wire_364),
        .c(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    spl2 new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_367),
        .b(new_Jinkela_wire_368),
        .c(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_424),
        .dout(new_Jinkela_wire_425)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    spl2 new_Jinkela_splitter_64 (
        .a(N210),
        .b(new_Jinkela_wire_439),
        .c(new_Jinkela_wire_444)
    );

    spl2 new_Jinkela_splitter_123 (
        .a(_217_),
        .b(new_Jinkela_wire_992),
        .c(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_385),
        .dout(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_951),
        .dout(new_Jinkela_wire_952)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_425),
        .dout(new_Jinkela_wire_426)
    );

    spl4L new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_386),
        .b(new_Jinkela_wire_387),
        .c(new_Jinkela_wire_388),
        .d(new_Jinkela_wire_389),
        .e(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    spl4L new_Jinkela_splitter_57 (
        .a(new_Jinkela_wire_390),
        .b(new_Jinkela_wire_391),
        .c(new_Jinkela_wire_392),
        .d(new_Jinkela_wire_393),
        .e(new_Jinkela_wire_394)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_952),
        .dout(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_436),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    spl2 new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_394),
        .b(new_Jinkela_wire_395),
        .c(new_Jinkela_wire_396)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_426),
        .dout(new_Jinkela_wire_427)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_net_534),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_427),
        .dout(new_Jinkela_wire_428)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_969),
        .dout(new_Jinkela_wire_970)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    spl4L new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_444),
        .b(new_Jinkela_wire_445),
        .c(new_Jinkela_wire_446),
        .d(new_Jinkela_wire_447),
        .e(new_Jinkela_wire_448)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(_277_),
        .b(new_Jinkela_wire_994),
        .c(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_399),
        .dout(new_Jinkela_wire_400)
    );

    spl4L new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_439),
        .b(new_Jinkela_wire_440),
        .c(new_Jinkela_wire_441),
        .d(new_Jinkela_wire_442),
        .e(new_Jinkela_wire_443)
    );

    spl2 new_Jinkela_splitter_67 (
        .a(N135),
        .b(new_Jinkela_wire_449),
        .c(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_400),
        .dout(new_Jinkela_wire_401)
    );

    spl2 new_Jinkela_splitter_125 (
        .a(_138_),
        .b(new_Jinkela_wire_997),
        .c(new_Jinkela_wire_998)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_972),
        .dout(new_Jinkela_wire_973)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    spl2 new_Jinkela_splitter_68 (
        .a(N237),
        .b(new_Jinkela_wire_451),
        .c(new_Jinkela_wire_452)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_431),
        .c(new_Jinkela_wire_432)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_403),
        .dout(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_432),
        .dout(new_Jinkela_wire_433)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_404),
        .dout(new_Jinkela_wire_405)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_5),
        .dout(new_Jinkela_wire_6)
    );

    or_ii _358_ (
        .a(new_Jinkela_wire_958),
        .b(new_Jinkela_wire_370),
        .c(_058_)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(new_Jinkela_wire_1846),
        .dout(new_Jinkela_wire_1847)
    );

    and_bi _359_ (
        .a(_058_),
        .b(new_Jinkela_wire_406),
        .c(_059_)
    );

    bfr new_Jinkela_buffer_29 (
        .din(N207),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_1858),
        .dout(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    and_bi _360_ (
        .a(new_Jinkela_wire_611),
        .b(_059_),
        .c(_060_)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_1847),
        .dout(new_Jinkela_wire_1848)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    and_bi _361_ (
        .a(new_Jinkela_wire_355),
        .b(new_Jinkela_wire_597),
        .c(_061_)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(new_Jinkela_wire_1896),
        .dout(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(_139_),
        .dout(new_Jinkela_wire_1936)
    );

    and_bi _362_ (
        .a(new_Jinkela_wire_894),
        .b(new_Jinkela_wire_957),
        .c(_062_)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_1848),
        .dout(new_Jinkela_wire_1849)
    );

    inv _363_ (
        .din(new_Jinkela_wire_451),
        .dout(_063_)
    );

    spl3L new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_25),
        .b(new_Jinkela_wire_26),
        .c(new_Jinkela_wire_27),
        .d(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(new_Jinkela_wire_1859),
        .dout(new_Jinkela_wire_1860)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    and_bi _364_ (
        .a(new_Jinkela_wire_938),
        .b(new_Jinkela_wire_1949),
        .c(_064_)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_1849),
        .dout(new_Jinkela_wire_1850)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    and_bi _365_ (
        .a(new_Jinkela_wire_313),
        .b(new_Jinkela_wire_1704),
        .c(_065_)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    or_ii _366_ (
        .a(new_Jinkela_wire_412),
        .b(new_Jinkela_wire_514),
        .c(_066_)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(new_Jinkela_wire_1850),
        .dout(new_Jinkela_wire_1851)
    );

    spl3L new_Jinkela_splitter_8 (
        .a(N255),
        .b(new_Jinkela_wire_49),
        .c(new_Jinkela_wire_50),
        .d(new_Jinkela_wire_51)
    );

    and_ii _367_ (
        .a(new_Jinkela_wire_1213),
        .b(new_Jinkela_wire_626),
        .c(_067_)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_1860),
        .dout(new_Jinkela_wire_1861)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    or_ii _368_ (
        .a(new_Jinkela_wire_500),
        .b(new_Jinkela_wire_165),
        .c(_068_)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(_063_),
        .dout(new_Jinkela_wire_1937)
    );

    and_bb _369_ (
        .a(new_Jinkela_wire_57),
        .b(new_Jinkela_wire_24),
        .c(_069_)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_1861),
        .dout(new_Jinkela_wire_1862)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    or_ii _370_ (
        .a(_069_),
        .b(new_Jinkela_wire_491),
        .c(_070_)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(new_Jinkela_wire_1897),
        .dout(new_Jinkela_wire_1898)
    );

    spl2 new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_28),
        .b(new_Jinkela_wire_29),
        .c(new_Jinkela_wire_30)
    );

    and_ii _371_ (
        .a(_070_),
        .b(new_Jinkela_wire_1721),
        .c(_071_)
    );

    spl3L new_Jinkela_splitter_10 (
        .a(N183),
        .b(new_Jinkela_wire_58),
        .c(new_Jinkela_wire_59),
        .d(new_Jinkela_wire_60)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_1862),
        .dout(new_Jinkela_wire_1863)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    or_ii _372_ (
        .a(new_Jinkela_wire_1499),
        .b(new_Jinkela_wire_1733),
        .c(_072_)
    );

    spl3L new_Jinkela_splitter_176 (
        .a(_085_),
        .b(new_Jinkela_wire_1962),
        .c(new_Jinkela_wire_1963),
        .d(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_32 (
        .din(N72),
        .dout(new_Jinkela_wire_57)
    );

    spl3L new_Jinkela_splitter_177 (
        .a(_033_),
        .b(new_Jinkela_wire_1988),
        .c(new_Jinkela_wire_1989),
        .d(new_Jinkela_wire_1990)
    );

    and_bi _373_ (
        .a(new_Jinkela_wire_127),
        .b(new_Jinkela_wire_594),
        .c(_073_)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_1863),
        .dout(new_Jinkela_wire_1864)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    and_bb _374_ (
        .a(new_Jinkela_wire_445),
        .b(new_Jinkela_wire_108),
        .c(_074_)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_1898),
        .dout(new_Jinkela_wire_1899)
    );

    or_bb _375_ (
        .a(new_Jinkela_wire_777),
        .b(_073_),
        .c(_075_)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_1864),
        .dout(new_Jinkela_wire_1865)
    );

    spl2 new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_18),
        .b(new_Jinkela_wire_19),
        .c(new_Jinkela_wire_20)
    );

    or_bb _376_ (
        .a(new_Jinkela_wire_1560),
        .b(_065_),
        .c(_076_)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(_215_),
        .dout(new_Jinkela_wire_1959)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_20),
        .dout(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_1959),
        .dout(new_Jinkela_wire_1960)
    );

    or_bb _377_ (
        .a(new_Jinkela_wire_1719),
        .b(_064_),
        .c(_077_)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_1865),
        .dout(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_33),
        .dout(new_Jinkela_wire_34)
    );

    or_bb _378_ (
        .a(new_Jinkela_wire_1141),
        .b(_062_),
        .c(_078_)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(new_Jinkela_wire_1899),
        .dout(new_Jinkela_wire_1900)
    );

    or_bb _379_ (
        .a(new_Jinkela_wire_1566),
        .b(_060_),
        .c(new_net_542)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(new_Jinkela_wire_1866),
        .dout(new_Jinkela_wire_1867)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    or_bi _380_ (
        .a(new_Jinkela_wire_1651),
        .b(new_Jinkela_wire_294),
        .c(_079_)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_1937),
        .dout(new_Jinkela_wire_1938)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_35),
        .dout(new_Jinkela_wire_36)
    );

    and_bi _381_ (
        .a(new_Jinkela_wire_242),
        .b(new_Jinkela_wire_2019),
        .c(_080_)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_1867),
        .dout(new_Jinkela_wire_1868)
    );

    and_bb _382_ (
        .a(new_Jinkela_wire_408),
        .b(new_Jinkela_wire_192),
        .c(_081_)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_36),
        .dout(new_Jinkela_wire_37)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    or_bb _383_ (
        .a(new_Jinkela_wire_1414),
        .b(new_Jinkela_wire_1723),
        .c(_082_)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_1868),
        .dout(new_Jinkela_wire_1869)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    or_bb _384_ (
        .a(_082_),
        .b(_080_),
        .c(_083_)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_37),
        .dout(new_Jinkela_wire_38)
    );

    and_bi _385_ (
        .a(_079_),
        .b(_083_),
        .c(_084_)
    );

    bfr new_Jinkela_buffer_45 (
        .din(N267),
        .dout(new_Jinkela_wire_79)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(new_Jinkela_wire_1869),
        .dout(new_Jinkela_wire_1870)
    );

    spl2 new_Jinkela_splitter_13 (
        .a(N75),
        .b(new_Jinkela_wire_77),
        .c(new_Jinkela_wire_78)
    );

    and_bi _386_ (
        .a(new_Jinkela_wire_539),
        .b(new_Jinkela_wire_839),
        .c(_085_)
    );

    bfr new_Jinkela_buffer_46 (
        .din(N146),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_38),
        .dout(new_Jinkela_wire_39)
    );

    and_bi _387_ (
        .a(new_Jinkela_wire_838),
        .b(new_Jinkela_wire_538),
        .c(_086_)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(new_Jinkela_wire_1870),
        .dout(new_Jinkela_wire_1871)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(new_Jinkela_wire_54),
        .b(new_Jinkela_wire_55),
        .c(new_Jinkela_wire_56)
    );

    and_ii _388_ (
        .a(new_Jinkela_wire_739),
        .b(new_Jinkela_wire_1963),
        .c(_087_)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_1938),
        .dout(new_Jinkela_wire_1939)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(new_Jinkela_wire_39),
        .b(new_Jinkela_wire_40),
        .c(new_Jinkela_wire_41)
    );

    or_bi _389_ (
        .a(new_Jinkela_wire_1658),
        .b(new_Jinkela_wire_206),
        .c(_088_)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(new_Jinkela_wire_1871),
        .dout(new_Jinkela_wire_1872)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_41),
        .dout(new_Jinkela_wire_42)
    );

    and_bi _390_ (
        .a(new_Jinkela_wire_88),
        .b(new_Jinkela_wire_2020),
        .c(_089_)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    and_bb _391_ (
        .a(new_Jinkela_wire_407),
        .b(new_Jinkela_wire_418),
        .c(_090_)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(new_Jinkela_wire_1872),
        .dout(new_Jinkela_wire_1873)
    );

    spl3L new_Jinkela_splitter_15 (
        .a(N111),
        .b(new_Jinkela_wire_92),
        .c(new_Jinkela_wire_93),
        .d(new_Jinkela_wire_94)
    );

    or_bb _392_ (
        .a(new_Jinkela_wire_1573),
        .b(new_Jinkela_wire_1724),
        .c(_091_)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_42),
        .dout(new_Jinkela_wire_43)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_1960),
        .dout(new_Jinkela_wire_1961)
    );

    or_bb _393_ (
        .a(_091_),
        .b(_089_),
        .c(_092_)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_1873),
        .dout(new_Jinkela_wire_1874)
    );

    and_bi _394_ (
        .a(_088_),
        .b(_092_),
        .c(_093_)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(new_Jinkela_wire_1903),
        .dout(new_Jinkela_wire_1904)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_43),
        .dout(new_Jinkela_wire_44)
    );

    and_bi _395_ (
        .a(new_Jinkela_wire_262),
        .b(new_Jinkela_wire_1051),
        .c(_094_)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(new_Jinkela_wire_1874),
        .dout(new_Jinkela_wire_1875)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    and_bi _396_ (
        .a(new_Jinkela_wire_1052),
        .b(new_Jinkela_wire_261),
        .c(_095_)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_1939),
        .dout(new_Jinkela_wire_1940)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_44),
        .dout(new_Jinkela_wire_45)
    );

    or_bi _397_ (
        .a(new_Jinkela_wire_1654),
        .b(new_Jinkela_wire_117),
        .c(_096_)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_1875),
        .dout(new_Jinkela_wire_1876)
    );

    and_bi _398_ (
        .a(new_Jinkela_wire_431),
        .b(new_Jinkela_wire_2018),
        .c(_097_)
    );

    spl3L new_Jinkela_splitter_17 (
        .a(N101),
        .b(new_Jinkela_wire_105),
        .c(new_Jinkela_wire_106),
        .d(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(new_Jinkela_wire_1904),
        .dout(new_Jinkela_wire_1905)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    and_bb _399_ (
        .a(new_Jinkela_wire_411),
        .b(new_Jinkela_wire_212),
        .c(_098_)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_Jinkela_wire_1876),
        .dout(new_Jinkela_wire_1877)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_567),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    bfr new_Jinkela_buffer_364 (
        .din(_161_),
        .dout(new_Jinkela_wire_579)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_555),
        .dout(new_Jinkela_wire_556)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_568),
        .dout(new_Jinkela_wire_569)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_557),
        .dout(new_Jinkela_wire_558)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_558),
        .dout(new_Jinkela_wire_559)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(_072_),
        .b(new_Jinkela_wire_585),
        .c(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_561),
        .dout(new_Jinkela_wire_562)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_562),
        .dout(new_Jinkela_wire_563)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_574),
        .dout(new_Jinkela_wire_575)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_563),
        .dout(new_Jinkela_wire_564)
    );

    spl4L new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_585),
        .b(new_Jinkela_wire_586),
        .c(new_Jinkela_wire_587),
        .d(new_Jinkela_wire_588),
        .e(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_564),
        .dout(new_Jinkela_wire_565)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_565),
        .dout(new_Jinkela_wire_566)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_581),
        .dout(new_Jinkela_wire_582)
    );

    spl3L new_Jinkela_splitter_92 (
        .a(_105_),
        .b(new_Jinkela_wire_614),
        .c(new_Jinkela_wire_615),
        .d(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    spl4L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_590),
        .b(new_Jinkela_wire_591),
        .c(new_Jinkela_wire_592),
        .d(new_Jinkela_wire_593),
        .e(new_Jinkela_wire_594)
    );

    spl2 new_Jinkela_splitter_89 (
        .a(_241_),
        .b(new_Jinkela_wire_595),
        .c(new_Jinkela_wire_596)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    spl2 new_Jinkela_splitter_90 (
        .a(_019_),
        .b(new_Jinkela_wire_597),
        .c(new_Jinkela_wire_598)
    );

    spl2 new_Jinkela_splitter_91 (
        .a(_235_),
        .b(new_Jinkela_wire_612),
        .c(new_Jinkela_wire_613)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_598),
        .dout(new_Jinkela_wire_599)
    );

    spl2 new_Jinkela_splitter_95 (
        .a(_009_),
        .b(new_Jinkela_wire_624),
        .c(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_599),
        .dout(new_Jinkela_wire_600)
    );

    spl4L new_Jinkela_splitter_93 (
        .a(_024_),
        .b(new_Jinkela_wire_617),
        .c(new_Jinkela_wire_618),
        .d(new_Jinkela_wire_619),
        .e(new_Jinkela_wire_620)
    );

    spl3L new_Jinkela_splitter_94 (
        .a(_049_),
        .b(new_Jinkela_wire_621),
        .c(new_Jinkela_wire_622),
        .d(new_Jinkela_wire_623)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_600),
        .dout(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1369),
        .dout(new_Jinkela_wire_1370)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1320),
        .dout(new_Jinkela_wire_1321)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1335),
        .dout(new_Jinkela_wire_1336)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_273),
        .dout(new_Jinkela_wire_274)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(new_Jinkela_wire_1401),
        .dout(new_Jinkela_wire_1402)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1336),
        .dout(new_Jinkela_wire_1337)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_274),
        .dout(new_Jinkela_wire_275)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1370),
        .dout(new_Jinkela_wire_1371)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_322),
        .dout(new_Jinkela_wire_323)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1337),
        .dout(new_Jinkela_wire_1338)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_275),
        .dout(new_Jinkela_wire_276)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1406),
        .dout(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_290),
        .dout(new_Jinkela_wire_291)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1338),
        .dout(new_Jinkela_wire_1339)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_276),
        .dout(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1371),
        .dout(new_Jinkela_wire_1372)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1339),
        .dout(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1402),
        .dout(new_Jinkela_wire_1403)
    );

    spl4L new_Jinkela_splitter_59 (
        .a(N138),
        .b(new_Jinkela_wire_407),
        .c(new_Jinkela_wire_408),
        .d(new_Jinkela_wire_409),
        .e(new_Jinkela_wire_410)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1340),
        .dout(new_Jinkela_wire_1341)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_278),
        .dout(new_Jinkela_wire_279)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1372),
        .dout(new_Jinkela_wire_1373)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1341),
        .dout(new_Jinkela_wire_1342)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_279),
        .dout(new_Jinkela_wire_280)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(_111_),
        .dout(new_Jinkela_wire_1415)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1342),
        .dout(new_Jinkela_wire_1343)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_280),
        .dout(new_Jinkela_wire_281)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1373),
        .dout(new_Jinkela_wire_1374)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1343),
        .dout(new_Jinkela_wire_1344)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1403),
        .dout(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1344),
        .dout(new_Jinkela_wire_1345)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_299),
        .dout(new_Jinkela_wire_300)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1374),
        .dout(new_Jinkela_wire_1375)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1345),
        .dout(new_Jinkela_wire_1346)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_323),
        .dout(new_Jinkela_wire_324)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(N13),
        .b(new_Jinkela_wire_412),
        .c(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1346),
        .dout(new_Jinkela_wire_1347)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1375),
        .dout(new_Jinkela_wire_1376)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_324),
        .dout(new_Jinkela_wire_325)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1347),
        .dout(new_Jinkela_wire_1348)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_Jinkela_wire_1404),
        .dout(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_325),
        .dout(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(new_Jinkela_wire_1348),
        .dout(new_Jinkela_wire_1349)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1376),
        .dout(new_Jinkela_wire_1377)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1349),
        .dout(new_Jinkela_wire_1350)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_305),
        .dout(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(_146_),
        .dout(new_Jinkela_wire_1477)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_340),
        .dout(new_Jinkela_wire_341)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(new_Jinkela_wire_1350),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_326),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1351),
        .dout(new_Jinkela_wire_1352)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(new_Jinkela_wire_307),
        .b(new_Jinkela_wire_308),
        .c(new_Jinkela_wire_310)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_311),
        .c(new_Jinkela_wire_312),
        .d(new_Jinkela_wire_313),
        .e(new_Jinkela_wire_314)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(new_Jinkela_wire_1352),
        .dout(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1378),
        .dout(new_Jinkela_wire_1379)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1353),
        .dout(new_Jinkela_wire_1354)
    );

    spl4L new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_314),
        .b(new_Jinkela_wire_315),
        .c(new_Jinkela_wire_316),
        .d(new_Jinkela_wire_317),
        .e(new_Jinkela_wire_318)
    );

    spl3L new_Jinkela_splitter_143 (
        .a(_094_),
        .b(new_Jinkela_wire_1454),
        .c(new_Jinkela_wire_1455),
        .d(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1354),
        .dout(new_Jinkela_wire_1355)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_318),
        .dout(new_Jinkela_wire_319)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1379),
        .dout(new_Jinkela_wire_1380)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_976),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_732 (
        .din(_150_),
        .dout(new_Jinkela_wire_1049)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    spl3L new_Jinkela_splitter_127 (
        .a(_093_),
        .b(new_Jinkela_wire_1050),
        .c(new_Jinkela_wire_1051),
        .d(new_Jinkela_wire_1052)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_net_528),
        .dout(new_Jinkela_wire_1053)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_767 (
        .din(_125_),
        .dout(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_1016),
        .dout(new_Jinkela_wire_1017)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_1017),
        .dout(new_Jinkela_wire_1018)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_1053),
        .dout(new_Jinkela_wire_1054)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_1018),
        .dout(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    spl3L new_Jinkela_splitter_128 (
        .a(_046_),
        .b(new_Jinkela_wire_1088),
        .c(new_Jinkela_wire_1089),
        .d(new_Jinkela_wire_1090)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_net_0),
        .dout(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_1054),
        .dout(new_Jinkela_wire_1055)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    spl2 new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_1011),
        .b(new_Jinkela_wire_1012),
        .c(new_Jinkela_wire_1013)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_1055),
        .dout(new_Jinkela_wire_1056)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_1022),
        .dout(new_Jinkela_wire_1023)
    );

    spl2 new_Jinkela_splitter_130 (
        .a(_273_),
        .b(new_Jinkela_wire_1142),
        .c(new_Jinkela_wire_1143)
    );

    bfr new_Jinkela_buffer_804 (
        .din(_077_),
        .dout(new_Jinkela_wire_1130)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_1023),
        .dout(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_1056),
        .dout(new_Jinkela_wire_1057)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    and_bi _568_ (
        .a(new_Jinkela_wire_183),
        .b(new_Jinkela_wire_829),
        .c(_253_)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_628),
        .dout(new_Jinkela_wire_629)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    and_bi _569_ (
        .a(new_Jinkela_wire_828),
        .b(new_Jinkela_wire_184),
        .c(_254_)
    );

    or_bb _570_ (
        .a(_254_),
        .b(_253_),
        .c(_255_)
    );

    spl3L new_Jinkela_splitter_97 (
        .a(_041_),
        .b(new_Jinkela_wire_631),
        .c(new_Jinkela_wire_632),
        .d(new_Jinkela_wire_633)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    and_bi _571_ (
        .a(new_Jinkela_wire_105),
        .b(new_Jinkela_wire_167),
        .c(_256_)
    );

    bfr new_Jinkela_buffer_384 (
        .din(_179_),
        .dout(new_Jinkela_wire_630)
    );

    and_bi _572_ (
        .a(new_Jinkela_wire_168),
        .b(new_Jinkela_wire_106),
        .c(_257_)
    );

    spl3L new_Jinkela_splitter_96 (
        .a(_286_),
        .b(new_Jinkela_wire_626),
        .c(new_Jinkela_wire_627),
        .d(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    and_ii _573_ (
        .a(_257_),
        .b(_256_),
        .c(_258_)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_net_522),
        .dout(new_Jinkela_wire_638)
    );

    and_ii _574_ (
        .a(new_Jinkela_wire_93),
        .b(new_Jinkela_wire_473),
        .c(_259_)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    and_bb _575_ (
        .a(new_Jinkela_wire_92),
        .b(new_Jinkela_wire_474),
        .c(_260_)
    );

    and_ii _576_ (
        .a(_260_),
        .b(_259_),
        .c(_261_)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    and_bi _577_ (
        .a(new_Jinkela_wire_1365),
        .b(new_Jinkela_wire_981),
        .c(_262_)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(_232_),
        .b(new_Jinkela_wire_656),
        .c(new_Jinkela_wire_657)
    );

    and_bi _578_ (
        .a(new_Jinkela_wire_980),
        .b(new_Jinkela_wire_1364),
        .c(_263_)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_633),
        .dout(new_Jinkela_wire_634)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    and_ii _579_ (
        .a(_263_),
        .b(_262_),
        .c(_264_)
    );

    bfr new_Jinkela_buffer_407 (
        .din(_036_),
        .dout(new_Jinkela_wire_658)
    );

    and_ii _580_ (
        .a(new_Jinkela_wire_1594),
        .b(new_Jinkela_wire_1501),
        .c(_265_)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    and_bb _581_ (
        .a(new_Jinkela_wire_1593),
        .b(new_Jinkela_wire_1500),
        .c(_266_)
    );

    and_ii _582_ (
        .a(_266_),
        .b(_265_),
        .c(_267_)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    and_bi _583_ (
        .a(new_Jinkela_wire_955),
        .b(new_Jinkela_wire_872),
        .c(_268_)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_634),
        .dout(new_Jinkela_wire_635)
    );

    and_bi _584_ (
        .a(new_Jinkela_wire_871),
        .b(new_Jinkela_wire_954),
        .c(_269_)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    or_bb _585_ (
        .a(_269_),
        .b(_268_),
        .c(new_net_520)
    );

    or_bi _586_ (
        .a(new_Jinkela_wire_1720),
        .b(new_Jinkela_wire_437),
        .c(_270_)
    );

    bfr new_Jinkela_buffer_418 (
        .din(_196_),
        .dout(new_Jinkela_wire_674)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    and_bi _587_ (
        .a(new_Jinkela_wire_1732),
        .b(new_Jinkela_wire_963),
        .c(new_net_534)
    );

    and_bi _588_ (
        .a(new_Jinkela_wire_29),
        .b(new_Jinkela_wire_624),
        .c(new_net_546)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    and_bi _589_ (
        .a(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_992),
        .c(new_net_552)
    );

    and_bb _590_ (
        .a(N86),
        .b(N85),
        .c(new_net_526)
    );

    spl3L new_Jinkela_splitter_100 (
        .a(_027_),
        .b(new_Jinkela_wire_671),
        .c(new_Jinkela_wire_672),
        .d(new_Jinkela_wire_673)
    );

    inv _591_ (
        .din(new_Jinkela_wire_879),
        .dout(new_net_536)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    or_ii _592_ (
        .a(new_Jinkela_wire_414),
        .b(new_Jinkela_wire_210),
        .c(_271_)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    and_ii _593_ (
        .a(new_Jinkela_wire_1199),
        .b(new_Jinkela_wire_629),
        .c(new_net_540)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    or_bb _594_ (
        .a(new_Jinkela_wire_1198),
        .b(new_Jinkela_wire_996),
        .c(_272_)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_net_552),
        .dout(new_Jinkela_wire_675)
    );

    or_bi _595_ (
        .a(new_Jinkela_wire_1201),
        .b(new_Jinkela_wire_1093),
        .c(new_net_556)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    and_ii _596_ (
        .a(N88),
        .b(N87),
        .c(_273_)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    and_bi _597_ (
        .a(new_Jinkela_wire_416),
        .b(new_Jinkela_wire_1143),
        .c(new_net_558)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    and_bi _598_ (
        .a(new_Jinkela_wire_472),
        .b(new_Jinkela_wire_1142),
        .c(new_net_538)
    );

    bfr new_Jinkela_buffer_472 (
        .din(_119_),
        .dout(new_Jinkela_wire_732)
    );

    or_bb _599_ (
        .a(new_Jinkela_wire_1200),
        .b(new_Jinkela_wire_1092),
        .c(new_net_528)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    spl2 new_Jinkela_splitter_101 (
        .a(_124_),
        .b(new_Jinkela_wire_712),
        .c(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_660),
        .dout(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_662),
        .dout(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1355),
        .dout(new_Jinkela_wire_1356)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1410),
        .dout(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_1605),
        .dout(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_1877),
        .dout(new_Jinkela_wire_1878)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1356),
        .dout(new_Jinkela_wire_1357)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_1905),
        .dout(new_Jinkela_wire_1906)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_1606),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(new_Jinkela_wire_1878),
        .dout(new_Jinkela_wire_1879)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1357),
        .dout(new_Jinkela_wire_1358)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(new_Jinkela_wire_1607),
        .dout(new_Jinkela_wire_1608)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(new_Jinkela_wire_1879),
        .dout(new_Jinkela_wire_1880)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    spl4L new_Jinkela_splitter_156 (
        .a(new_Jinkela_wire_1650),
        .b(new_Jinkela_wire_1651),
        .c(new_Jinkela_wire_1652),
        .d(new_Jinkela_wire_1653),
        .e(new_Jinkela_wire_1654)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_1906),
        .dout(new_Jinkela_wire_1907)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(new_Jinkela_wire_1644),
        .dout(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1411),
        .dout(new_Jinkela_wire_1412)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_1608),
        .dout(new_Jinkela_wire_1609)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(new_Jinkela_wire_1880),
        .dout(new_Jinkela_wire_1881)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_1940),
        .dout(new_Jinkela_wire_1941)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(_152_),
        .b(new_Jinkela_wire_1682),
        .c(new_Jinkela_wire_1683)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_1941),
        .dout(new_Jinkela_wire_1942)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_1609),
        .dout(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(new_Jinkela_wire_1881),
        .dout(new_Jinkela_wire_1882)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(_223_),
        .dout(new_Jinkela_wire_1483)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(new_Jinkela_wire_1383),
        .dout(new_Jinkela_wire_1384)
    );

    spl3L new_Jinkela_splitter_160 (
        .a(_107_),
        .b(new_Jinkela_wire_1679),
        .c(new_Jinkela_wire_1680),
        .d(new_Jinkela_wire_1681)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_1907),
        .dout(new_Jinkela_wire_1908)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(new_Jinkela_wire_1645),
        .dout(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1412),
        .dout(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_1610),
        .dout(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(new_Jinkela_wire_1882),
        .dout(new_Jinkela_wire_1883)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(new_Jinkela_wire_1384),
        .dout(new_Jinkela_wire_1385)
    );

    spl2 new_Jinkela_splitter_178 (
        .a(_095_),
        .b(new_Jinkela_wire_1997),
        .c(new_Jinkela_wire_1998)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(_132_),
        .dout(new_Jinkela_wire_1991)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(_134_),
        .dout(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(new_Jinkela_wire_1611),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(new_Jinkela_wire_1883),
        .dout(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1385),
        .dout(new_Jinkela_wire_1386)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_1662),
        .dout(new_Jinkela_wire_1663)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(new_Jinkela_wire_1908),
        .dout(new_Jinkela_wire_1909)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1413),
        .dout(new_Jinkela_wire_1414)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_1884),
        .dout(new_Jinkela_wire_1885)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1386),
        .dout(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(_207_),
        .dout(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_1964),
        .dout(new_Jinkela_wire_1965)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(new_Jinkela_wire_1613),
        .dout(new_Jinkela_wire_1614)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_1885),
        .dout(new_Jinkela_wire_1886)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1387),
        .dout(new_Jinkela_wire_1388)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(new_Jinkela_wire_1909),
        .dout(new_Jinkela_wire_1910)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_1647),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(new_Jinkela_wire_1614),
        .dout(new_Jinkela_wire_1615)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(new_Jinkela_wire_1886),
        .dout(new_Jinkela_wire_1887)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1388),
        .dout(new_Jinkela_wire_1389)
    );

    spl4L new_Jinkela_splitter_179 (
        .a(_005_),
        .b(new_Jinkela_wire_2018),
        .c(new_Jinkela_wire_2019),
        .d(new_Jinkela_wire_2020),
        .e(new_Jinkela_wire_2021)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_1663),
        .dout(new_Jinkela_wire_1664)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_1942),
        .dout(new_Jinkela_wire_1943)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(new_Jinkela_wire_1615),
        .dout(new_Jinkela_wire_1616)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_Jinkela_wire_1887),
        .dout(new_Jinkela_wire_1888)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1389),
        .dout(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_1910),
        .dout(new_Jinkela_wire_1911)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_1616),
        .dout(new_Jinkela_wire_1617)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1390),
        .dout(new_Jinkela_wire_1391)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(new_Jinkela_wire_1911),
        .dout(new_Jinkela_wire_1912)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(new_net_564),
        .dout(new_Jinkela_wire_1692)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(new_Jinkela_wire_1617),
        .dout(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_1943),
        .dout(new_Jinkela_wire_1944)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1391),
        .dout(new_Jinkela_wire_1392)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(new_Jinkela_wire_1912),
        .dout(new_Jinkela_wire_1913)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(new_Jinkela_wire_1664),
        .dout(new_Jinkela_wire_1665)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_1618),
        .dout(new_Jinkela_wire_1619)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_1991),
        .dout(new_Jinkela_wire_1992)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1392),
        .dout(new_Jinkela_wire_1393)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(new_Jinkela_wire_1913),
        .dout(new_Jinkela_wire_1914)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(new_Jinkela_wire_1683),
        .dout(new_Jinkela_wire_1684)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_1619),
        .dout(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_1944),
        .dout(new_Jinkela_wire_1945)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1393),
        .dout(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_1665),
        .dout(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_1914),
        .dout(new_Jinkela_wire_1915)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_1620),
        .dout(new_Jinkela_wire_1621)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_1966),
        .dout(new_Jinkela_wire_1967)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1394),
        .dout(new_Jinkela_wire_1395)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(new_Jinkela_wire_1915),
        .dout(new_Jinkela_wire_1916)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(new_Jinkela_wire_1621),
        .dout(new_Jinkela_wire_1622)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_1945),
        .dout(new_Jinkela_wire_1946)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    spl3L new_Jinkela_splitter_163 (
        .a(_016_),
        .b(new_Jinkela_wire_1704),
        .c(new_Jinkela_wire_1705),
        .d(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(new_Jinkela_wire_1916),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_1666),
        .dout(new_Jinkela_wire_1667)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_1622),
        .dout(new_Jinkela_wire_1623)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(new_Jinkela_wire_1396),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(new_Jinkela_wire_1917),
        .dout(new_Jinkela_wire_1918)
    );

    spl3L new_Jinkela_splitter_164 (
        .a(_051_),
        .b(new_Jinkela_wire_1707),
        .c(new_Jinkela_wire_1708),
        .d(new_Jinkela_wire_1709)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(new_Jinkela_wire_1623),
        .dout(new_Jinkela_wire_1624)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_1946),
        .dout(new_Jinkela_wire_1947)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(new_Jinkela_wire_1684),
        .dout(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(new_Jinkela_wire_1918),
        .dout(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_1667),
        .dout(new_Jinkela_wire_1668)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_1624),
        .dout(new_Jinkela_wire_1625)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_1422),
        .dout(new_Jinkela_wire_1423)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_1967),
        .dout(new_Jinkela_wire_1968)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1398),
        .dout(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_1919),
        .dout(new_Jinkela_wire_1920)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_1625),
        .dout(new_Jinkela_wire_1626)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_1057),
        .dout(new_Jinkela_wire_1058)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    bfr new_Jinkela_buffer_816 (
        .din(_210_),
        .dout(new_Jinkela_wire_1144)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_1058),
        .dout(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1130),
        .dout(new_Jinkela_wire_1131)
    );

    spl3L new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_1091),
        .b(new_Jinkela_wire_1092),
        .c(new_Jinkela_wire_1093),
        .d(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_1059),
        .dout(new_Jinkela_wire_1060)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_1030),
        .dout(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_1060),
        .dout(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_821 (
        .din(_122_),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_1095),
        .dout(new_Jinkela_wire_1096)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_1061),
        .dout(new_Jinkela_wire_1062)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_1062),
        .dout(new_Jinkela_wire_1063)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1131),
        .dout(new_Jinkela_wire_1132)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_1039),
        .dout(new_Jinkela_wire_1040)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_1040),
        .dout(new_Jinkela_wire_1041)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_1097),
        .dout(new_Jinkela_wire_1098)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_1041),
        .dout(new_Jinkela_wire_1042)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_1042),
        .dout(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_1044),
        .dout(new_Jinkela_wire_1045)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1132),
        .dout(new_Jinkela_wire_1133)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1098),
        .dout(new_Jinkela_wire_1099)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_1045),
        .dout(new_Jinkela_wire_1046)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    or_bb _400_ (
        .a(new_Jinkela_wire_2027),
        .b(new_Jinkela_wire_1722),
        .c(_099_)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    or_bb _401_ (
        .a(_099_),
        .b(_097_),
        .c(_100_)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    and_bi _402_ (
        .a(_096_),
        .b(_100_),
        .c(_101_)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_676),
        .dout(new_Jinkela_wire_677)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    and_bi _403_ (
        .a(new_Jinkela_wire_162),
        .b(new_Jinkela_wire_961),
        .c(_102_)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    and_bi _404_ (
        .a(new_Jinkela_wire_960),
        .b(new_Jinkela_wire_161),
        .c(_103_)
    );

    or_bi _405_ (
        .a(new_Jinkela_wire_959),
        .b(new_Jinkela_wire_1592),
        .c(_104_)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    and_bi _406_ (
        .a(_104_),
        .b(new_Jinkela_wire_953),
        .c(_105_)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_664),
        .dout(new_Jinkela_wire_665)
    );

    or_bb _407_ (
        .a(new_Jinkela_wire_615),
        .b(new_Jinkela_wire_804),
        .c(_106_)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    and_bi _408_ (
        .a(_106_),
        .b(new_Jinkela_wire_824),
        .c(_107_)
    );

    bfr new_Jinkela_buffer_478 (
        .din(_176_),
        .dout(new_Jinkela_wire_738)
    );

    or_bb _409_ (
        .a(new_Jinkela_wire_1680),
        .b(new_Jinkela_wire_2017),
        .c(_108_)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    and_bi _410_ (
        .a(_108_),
        .b(new_Jinkela_wire_1476),
        .c(_109_)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_665),
        .dout(new_Jinkela_wire_666)
    );

    or_bi _411_ (
        .a(new_Jinkela_wire_863),
        .b(new_Jinkela_wire_1152),
        .c(_110_)
    );

    inv _412_ (
        .din(new_Jinkela_wire_338),
        .dout(_111_)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_666),
        .dout(new_Jinkela_wire_667)
    );

    and_bi _413_ (
        .a(new_Jinkela_wire_862),
        .b(new_Jinkela_wire_1153),
        .c(_112_)
    );

    or_bb _414_ (
        .a(_112_),
        .b(new_Jinkela_wire_1453),
        .c(_113_)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_678),
        .dout(new_Jinkela_wire_679)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_667),
        .dout(new_Jinkela_wire_668)
    );

    and_bi _415_ (
        .a(new_Jinkela_wire_786),
        .b(_113_),
        .c(_114_)
    );

    and_bb _416_ (
        .a(new_Jinkela_wire_841),
        .b(new_Jinkela_wire_387),
        .c(_115_)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    spl2 new_Jinkela_splitter_99 (
        .a(new_Jinkela_wire_668),
        .b(new_Jinkela_wire_669),
        .c(new_Jinkela_wire_670)
    );

    and_bi _417_ (
        .a(new_Jinkela_wire_1962),
        .b(new_Jinkela_wire_1953),
        .c(_116_)
    );

    and_bi _418_ (
        .a(new_Jinkela_wire_309),
        .b(new_Jinkela_wire_840),
        .c(_117_)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    and_bi _419_ (
        .a(new_Jinkela_wire_532),
        .b(new_Jinkela_wire_591),
        .c(_118_)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    and_bb _420_ (
        .a(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_2),
        .c(_119_)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    or_bb _421_ (
        .a(new_Jinkela_wire_737),
        .b(_118_),
        .c(_120_)
    );

    bfr new_Jinkela_buffer_501 (
        .din(_135_),
        .dout(new_Jinkela_wire_763)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(_086_),
        .b(new_Jinkela_wire_739),
        .c(new_Jinkela_wire_740)
    );

    or_bb _422_ (
        .a(new_Jinkela_wire_1892),
        .b(_117_),
        .c(_121_)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    or_bb _423_ (
        .a(new_Jinkela_wire_956),
        .b(_116_),
        .c(_122_)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    or_bb _424_ (
        .a(new_Jinkela_wire_1149),
        .b(_115_),
        .c(_123_)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_682),
        .dout(new_Jinkela_wire_683)
    );

    or_bb _425_ (
        .a(new_Jinkela_wire_1765),
        .b(_114_),
        .c(N878)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    and_ii _426_ (
        .a(new_Jinkela_wire_1997),
        .b(new_Jinkela_wire_1455),
        .c(_124_)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    or_bi _427_ (
        .a(new_Jinkela_wire_1679),
        .b(new_Jinkela_wire_731),
        .c(_125_)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_716),
        .dout(new_Jinkela_wire_717)
    );

    and_bi _428_ (
        .a(new_Jinkela_wire_1681),
        .b(new_Jinkela_wire_730),
        .c(_126_)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    or_bb _429_ (
        .a(_126_),
        .b(new_Jinkela_wire_1449),
        .c(_127_)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    and_bi _430_ (
        .a(new_Jinkela_wire_1087),
        .b(_127_),
        .c(_128_)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    and_bb _431_ (
        .a(new_Jinkela_wire_712),
        .b(new_Jinkela_wire_389),
        .c(_129_)
    );

    and_bi _432_ (
        .a(new_Jinkela_wire_1454),
        .b(new_Jinkela_wire_1951),
        .c(_130_)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_686),
        .dout(new_Jinkela_wire_687)
    );

    and_bi _433_ (
        .a(new_Jinkela_wire_311),
        .b(new_Jinkela_wire_1050),
        .c(_131_)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    and_bb _434_ (
        .a(new_Jinkela_wire_448),
        .b(new_Jinkela_wire_283),
        .c(_132_)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    and_bi _435_ (
        .a(new_Jinkela_wire_255),
        .b(new_Jinkela_wire_586),
        .c(_133_)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    or_bb _436_ (
        .a(_133_),
        .b(new_Jinkela_wire_1996),
        .c(_134_)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    or_bb _437_ (
        .a(new_Jinkela_wire_1491),
        .b(_131_),
        .c(_135_)
    );

    or_bb _438_ (
        .a(new_Jinkela_wire_763),
        .b(_130_),
        .c(_136_)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    or_bb _439_ (
        .a(new_Jinkela_wire_1744),
        .b(_129_),
        .c(_137_)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    or_bb _440_ (
        .a(new_Jinkela_wire_2047),
        .b(_128_),
        .c(new_net_548)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    and_ii _441_ (
        .a(new_Jinkela_wire_787),
        .b(new_Jinkela_wire_806),
        .c(_138_)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_1046),
        .dout(new_Jinkela_wire_1047)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(new_Jinkela_wire_1692),
        .dout(new_Jinkela_wire_1693)
    );

    spl2 new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_46),
        .b(new_Jinkela_wire_47),
        .c(new_Jinkela_wire_48)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_1668),
        .dout(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_1626),
        .dout(new_Jinkela_wire_1627)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_1047),
        .dout(new_Jinkela_wire_1048)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_80),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_1068),
        .dout(new_Jinkela_wire_1069)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_1627),
        .dout(new_Jinkela_wire_1628)
    );

    spl2 new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_94),
        .b(new_Jinkela_wire_95),
        .c(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1144),
        .dout(new_Jinkela_wire_1145)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1099),
        .dout(new_Jinkela_wire_1100)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_1069),
        .dout(new_Jinkela_wire_1070)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_1628),
        .dout(new_Jinkela_wire_1629)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_65),
        .dout(new_Jinkela_wire_66)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_1070),
        .dout(new_Jinkela_wire_1071)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(new_Jinkela_wire_1629),
        .dout(new_Jinkela_wire_1630)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1133),
        .dout(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_net_542),
        .dout(new_Jinkela_wire_1710)
    );

    spl2 new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_66),
        .b(new_Jinkela_wire_67),
        .c(new_Jinkela_wire_68)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1100),
        .dout(new_Jinkela_wire_1101)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(new_Jinkela_wire_1670),
        .dout(new_Jinkela_wire_1671)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_1630),
        .dout(new_Jinkela_wire_1631)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(_076_),
        .dout(new_Jinkela_wire_1719)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_1072),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(new_Jinkela_wire_1686),
        .dout(new_Jinkela_wire_1687)
    );

    spl3L new_Jinkela_splitter_19 (
        .a(N177),
        .b(new_Jinkela_wire_118),
        .c(new_Jinkela_wire_119),
        .d(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_1671),
        .dout(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_822 (
        .din(_197_),
        .dout(new_Jinkela_wire_1150)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1101),
        .dout(new_Jinkela_wire_1102)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_1073),
        .dout(new_Jinkela_wire_1074)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(new_Jinkela_wire_1693),
        .dout(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_1672),
        .dout(new_Jinkela_wire_1673)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_70),
        .dout(new_Jinkela_wire_71)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_1074),
        .dout(new_Jinkela_wire_1075)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(new_Jinkela_wire_1687),
        .dout(new_Jinkela_wire_1688)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(new_Jinkela_wire_1673),
        .dout(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1134),
        .dout(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_71),
        .dout(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_1075),
        .dout(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    spl2 new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_1674),
        .b(new_Jinkela_wire_1675),
        .c(new_Jinkela_wire_1676)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_1676),
        .dout(new_Jinkela_wire_1677)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_1076),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_1145),
        .dout(new_Jinkela_wire_1146)
    );

    spl2 new_Jinkela_splitter_162 (
        .a(new_Jinkela_wire_1688),
        .b(new_Jinkela_wire_1689),
        .c(new_Jinkela_wire_1690)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_73),
        .dout(new_Jinkela_wire_74)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_1677),
        .dout(new_Jinkela_wire_1678)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(new_Jinkela_wire_74),
        .b(new_Jinkela_wire_75),
        .c(new_Jinkela_wire_76)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(new_Jinkela_wire_1694),
        .dout(new_Jinkela_wire_1695)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1135),
        .dout(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(new_Jinkela_wire_1695),
        .dout(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_1710),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_109),
        .dout(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_1696),
        .dout(new_Jinkela_wire_1697)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_87),
        .b(new_Jinkela_wire_88),
        .c(new_Jinkela_wire_89)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_1080),
        .dout(new_Jinkela_wire_1081)
    );

    spl2 new_Jinkela_splitter_165 (
        .a(_068_),
        .b(new_Jinkela_wire_1720),
        .c(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    spl4L new_Jinkela_splitter_166 (
        .a(_013_),
        .b(new_Jinkela_wire_1722),
        .c(new_Jinkela_wire_1723),
        .d(new_Jinkela_wire_1724),
        .e(new_Jinkela_wire_1725)
    );

    spl3L new_Jinkela_splitter_131 (
        .a(_109_),
        .b(new_Jinkela_wire_1151),
        .c(new_Jinkela_wire_1152),
        .d(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(new_Jinkela_wire_1697),
        .dout(new_Jinkela_wire_1698)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(new_Jinkela_wire_107),
        .b(new_Jinkela_wire_108),
        .c(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1105),
        .dout(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_1711),
        .dout(new_Jinkela_wire_1712)
    );

    spl4L new_Jinkela_splitter_22 (
        .a(N195),
        .b(new_Jinkela_wire_135),
        .c(new_Jinkela_wire_136),
        .d(new_Jinkela_wire_137),
        .e(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_1698),
        .dout(new_Jinkela_wire_1699)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_net_524),
        .dout(new_Jinkela_wire_1154)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1136),
        .dout(new_Jinkela_wire_1137)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_Jinkela_wire_1699),
        .dout(new_Jinkela_wire_1700)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_1712),
        .dout(new_Jinkela_wire_1713)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_100),
        .dout(new_Jinkela_wire_101)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_1700),
        .dout(new_Jinkela_wire_1701)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_1084),
        .dout(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_101),
        .dout(new_Jinkela_wire_102)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1146),
        .dout(new_Jinkela_wire_1147)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(new_Jinkela_wire_1701),
        .dout(new_Jinkela_wire_1702)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    spl4L new_Jinkela_splitter_26 (
        .a(N59),
        .b(new_Jinkela_wire_163),
        .c(new_Jinkela_wire_164),
        .d(new_Jinkela_wire_165),
        .e(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_1085),
        .dout(new_Jinkela_wire_1086)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(new_Jinkela_wire_1713),
        .dout(new_Jinkela_wire_1714)
    );

    spl3L new_Jinkela_splitter_23 (
        .a(N171),
        .b(new_Jinkela_wire_146),
        .c(new_Jinkela_wire_147),
        .d(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_102),
        .dout(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(new_Jinkela_wire_1702),
        .dout(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1137),
        .dout(new_Jinkela_wire_1138)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(_246_),
        .b(new_Jinkela_wire_1726),
        .c(new_Jinkela_wire_1727)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(_211_),
        .dout(new_Jinkela_wire_1729)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(new_Jinkela_wire_1714),
        .dout(new_Jinkela_wire_1715)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(_010_),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_691),
        .dout(new_Jinkela_wire_692)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_692),
        .dout(new_Jinkela_wire_693)
    );

    spl2 new_Jinkela_splitter_104 (
        .a(_226_),
        .b(new_Jinkela_wire_764),
        .c(new_Jinkela_wire_765)
    );

    bfr new_Jinkela_buffer_502 (
        .din(_162_),
        .dout(new_Jinkela_wire_766)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_693),
        .dout(new_Jinkela_wire_694)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_721),
        .dout(new_Jinkela_wire_722)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_694),
        .dout(new_Jinkela_wire_695)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_695),
        .dout(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_722),
        .dout(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_696),
        .dout(new_Jinkela_wire_697)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_697),
        .dout(new_Jinkela_wire_698)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_698),
        .dout(new_Jinkela_wire_699)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_702),
        .dout(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_726),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_704),
        .dout(new_Jinkela_wire_705)
    );

    bfr new_Jinkela_buffer_508 (
        .din(_074_),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_705),
        .dout(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    spl2 new_Jinkela_splitter_105 (
        .a(_035_),
        .b(new_Jinkela_wire_778),
        .c(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(new_Jinkela_wire_729),
        .b(new_Jinkela_wire_730),
        .c(new_Jinkela_wire_731)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_520 (
        .din(_110_),
        .dout(new_Jinkela_wire_786)
    );

    spl2 new_Jinkela_splitter_173 (
        .a(new_Jinkela_wire_1947),
        .b(new_Jinkela_wire_1948),
        .c(new_Jinkela_wire_1950)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(new_Jinkela_wire_1920),
        .dout(new_Jinkela_wire_1921)
    );

    spl4L new_Jinkela_splitter_174 (
        .a(new_Jinkela_wire_1950),
        .b(new_Jinkela_wire_1951),
        .c(new_Jinkela_wire_1952),
        .d(new_Jinkela_wire_1953),
        .e(new_Jinkela_wire_1954)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_1921),
        .dout(new_Jinkela_wire_1922)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_1948),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_1922),
        .dout(new_Jinkela_wire_1923)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_1998),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(new_Jinkela_wire_1923),
        .dout(new_Jinkela_wire_1924)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    spl3L new_Jinkela_splitter_175 (
        .a(new_Jinkela_wire_1954),
        .b(new_Jinkela_wire_1955),
        .c(new_Jinkela_wire_1956),
        .d(new_Jinkela_wire_1957)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(new_Jinkela_wire_1924),
        .dout(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_1968),
        .dout(new_Jinkela_wire_1969)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(new_Jinkela_wire_1925),
        .dout(new_Jinkela_wire_1926)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_1926),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(new_Jinkela_wire_1969),
        .dout(new_Jinkela_wire_1970)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(new_Jinkela_wire_1928),
        .dout(new_Jinkela_wire_1929)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(_098_),
        .dout(new_Jinkela_wire_2022)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(new_Jinkela_wire_1929),
        .dout(new_Jinkela_wire_1930)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_1993),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(new_Jinkela_wire_1970),
        .dout(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(new_Jinkela_wire_1930),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_Jinkela_wire_1931),
        .dout(new_Jinkela_wire_1932)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(new_Jinkela_wire_1971),
        .dout(new_Jinkela_wire_1972)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_1932),
        .dout(new_Jinkela_wire_1933)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_1933),
        .dout(new_Jinkela_wire_1934)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(new_Jinkela_wire_1972),
        .dout(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_1934),
        .dout(new_Jinkela_wire_1935)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(_180_),
        .dout(new_Jinkela_wire_2029)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(new_Jinkela_wire_1973),
        .dout(new_Jinkela_wire_1974)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(new_Jinkela_wire_1974),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_1975),
        .dout(new_Jinkela_wire_1976)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_1976),
        .dout(new_Jinkela_wire_1977)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_2000),
        .dout(new_Jinkela_wire_2001)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_1977),
        .dout(new_Jinkela_wire_1978)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(_191_),
        .dout(new_Jinkela_wire_2028)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(new_Jinkela_wire_1978),
        .dout(new_Jinkela_wire_1979)
    );

    or_bi _442_ (
        .a(new_Jinkela_wire_616),
        .b(new_Jinkela_wire_1013),
        .c(_139_)
    );

    and_bi _443_ (
        .a(new_Jinkela_wire_614),
        .b(new_Jinkela_wire_1012),
        .c(_140_)
    );

    or_bb _444_ (
        .a(_140_),
        .b(new_Jinkela_wire_1445),
        .c(_141_)
    );

    and_bi _445_ (
        .a(new_Jinkela_wire_1936),
        .b(_141_),
        .c(_142_)
    );

    and_bb _446_ (
        .a(new_Jinkela_wire_997),
        .b(new_Jinkela_wire_388),
        .c(_143_)
    );

    and_bi _447_ (
        .a(new_Jinkela_wire_805),
        .b(new_Jinkela_wire_1952),
        .c(_144_)
    );

    and_bi _448_ (
        .a(new_Jinkela_wire_312),
        .b(new_Jinkela_wire_962),
        .c(_145_)
    );

    and_bb _449_ (
        .a(new_Jinkela_wire_441),
        .b(new_Jinkela_wire_197),
        .c(_146_)
    );

    and_bi _450_ (
        .a(new_Jinkela_wire_155),
        .b(new_Jinkela_wire_593),
        .c(_147_)
    );

    or_bb _451_ (
        .a(_147_),
        .b(new_Jinkela_wire_1482),
        .c(_148_)
    );

    or_bb _452_ (
        .a(new_Jinkela_wire_867),
        .b(_145_),
        .c(_149_)
    );

    or_bb _453_ (
        .a(new_Jinkela_wire_547),
        .b(_144_),
        .c(_150_)
    );

    or_bb _454_ (
        .a(new_Jinkela_wire_1049),
        .b(_143_),
        .c(_151_)
    );

    or_bb _455_ (
        .a(new_Jinkela_wire_979),
        .b(_142_),
        .c(new_net_532)
    );

    and_ii _456_ (
        .a(new_Jinkela_wire_1543),
        .b(new_Jinkela_wire_1639),
        .c(_152_)
    );

    and_bi _457_ (
        .a(new_Jinkela_wire_1768),
        .b(new_Jinkela_wire_1690),
        .c(_153_)
    );

    and_bi _458_ (
        .a(new_Jinkela_wire_1689),
        .b(new_Jinkela_wire_1766),
        .c(_154_)
    );

    or_bb _459_ (
        .a(_154_),
        .b(_153_),
        .c(_155_)
    );

    and_bi _460_ (
        .a(new_Jinkela_wire_368),
        .b(_155_),
        .c(_156_)
    );

    and_bb _461_ (
        .a(new_Jinkela_wire_1682),
        .b(new_Jinkela_wire_395),
        .c(_157_)
    );

    and_bi _462_ (
        .a(new_Jinkela_wire_1638),
        .b(new_Jinkela_wire_1958),
        .c(_158_)
    );

    and_bi _463_ (
        .a(new_Jinkela_wire_319),
        .b(new_Jinkela_wire_673),
        .c(_159_)
    );

    and_bi _464_ (
        .a(new_Jinkela_wire_67),
        .b(new_Jinkela_wire_589),
        .c(_160_)
    );

    and_bb _465_ (
        .a(new_Jinkela_wire_440),
        .b(new_Jinkela_wire_170),
        .c(_161_)
    );

    or_bb _466_ (
        .a(new_Jinkela_wire_584),
        .b(_160_),
        .c(_162_)
    );

    or_bb _467_ (
        .a(new_Jinkela_wire_771),
        .b(_159_),
        .c(_163_)
    );

    or_bb _468_ (
        .a(new_Jinkela_wire_1574),
        .b(_158_),
        .c(_164_)
    );

    or_bb _469_ (
        .a(new_Jinkela_wire_1893),
        .b(_157_),
        .c(_165_)
    );

    or_bb _470_ (
        .a(new_Jinkela_wire_578),
        .b(_156_),
        .c(new_net_564)
    );

    and_bi _471_ (
        .a(new_Jinkela_wire_778),
        .b(new_Jinkela_wire_982),
        .c(_166_)
    );

    and_bi _472_ (
        .a(new_Jinkela_wire_1575),
        .b(new_Jinkela_wire_1197),
        .c(_167_)
    );

    and_bi _473_ (
        .a(new_Jinkela_wire_1196),
        .b(new_Jinkela_wire_1577),
        .c(_168_)
    );

    or_bb _474_ (
        .a(_168_),
        .b(_167_),
        .c(_169_)
    );

    and_bi _475_ (
        .a(new_Jinkela_wire_364),
        .b(_169_),
        .c(_170_)
    );

    and_bb _476_ (
        .a(new_Jinkela_wire_1191),
        .b(new_Jinkela_wire_393),
        .c(_171_)
    );

    and_bi _477_ (
        .a(new_Jinkela_wire_983),
        .b(new_Jinkela_wire_1955),
        .c(_172_)
    );

    and_bi _478_ (
        .a(new_Jinkela_wire_316),
        .b(new_Jinkela_wire_1988),
        .c(_173_)
    );

    and_bi _479_ (
        .a(new_Jinkela_wire_329),
        .b(new_Jinkela_wire_587),
        .c(_174_)
    );

    and_bb _480_ (
        .a(new_Jinkela_wire_446),
        .b(new_Jinkela_wire_95),
        .c(_175_)
    );

    and_bb _481_ (
        .a(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_50),
        .c(_176_)
    );

    or_bb _482_ (
        .a(new_Jinkela_wire_738),
        .b(_175_),
        .c(_177_)
    );

    or_bb _483_ (
        .a(new_Jinkela_wire_837),
        .b(_174_),
        .c(_178_)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1109),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(_007_),
        .dout(new_Jinkela_wire_1492)
    );

    spl2 new_Jinkela_splitter_134 (
        .a(_271_),
        .b(new_Jinkela_wire_1198),
        .c(new_Jinkela_wire_1199)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1138),
        .dout(new_Jinkela_wire_1139)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1147),
        .dout(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_1483),
        .dout(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_Jinkela_wire_1479),
        .dout(new_Jinkela_wire_1480)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_1139),
        .dout(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_1426),
        .dout(new_Jinkela_wire_1427)
    );

    spl2 new_Jinkela_splitter_132 (
        .a(_166_),
        .b(new_Jinkela_wire_1191),
        .c(new_Jinkela_wire_1192)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1140),
        .dout(new_Jinkela_wire_1141)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_1428),
        .dout(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1154),
        .dout(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_1480),
        .dout(new_Jinkela_wire_1481)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1116),
        .dout(new_Jinkela_wire_1117)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_863 (
        .din(_193_),
        .dout(new_Jinkela_wire_1202)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(new_Jinkela_wire_1430),
        .b(new_Jinkela_wire_1431),
        .c(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1155),
        .dout(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_1488),
        .dout(new_Jinkela_wire_1489)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_1202),
        .dout(new_Jinkela_wire_1203)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1156),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_1484),
        .dout(new_Jinkela_wire_1485)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_1481),
        .dout(new_Jinkela_wire_1482)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1192),
        .dout(new_Jinkela_wire_1193)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_1465),
        .dout(new_Jinkela_wire_1466)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(_272_),
        .b(new_Jinkela_wire_1200),
        .c(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(new_Jinkela_wire_1435),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1122),
        .dout(new_Jinkela_wire_1123)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_1466),
        .dout(new_Jinkela_wire_1467)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1193),
        .dout(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_1123),
        .dout(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(_071_),
        .dout(new_Jinkela_wire_1499)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(new_Jinkela_wire_1438),
        .dout(new_Jinkela_wire_1439)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_1467),
        .dout(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_1439),
        .dout(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1159),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    spl2 new_Jinkela_splitter_144 (
        .a(new_Jinkela_wire_1485),
        .b(new_Jinkela_wire_1486),
        .c(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_1440),
        .dout(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1126),
        .dout(new_Jinkela_wire_1127)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(new_Jinkela_wire_1468),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1127),
        .dout(new_Jinkela_wire_1128)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(new_Jinkela_wire_1492),
        .dout(new_Jinkela_wire_1493)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(new_Jinkela_wire_1442),
        .dout(new_Jinkela_wire_1443)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1194),
        .dout(new_Jinkela_wire_1195)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1128),
        .dout(new_Jinkela_wire_1129)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_1469),
        .dout(new_Jinkela_wire_1470)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_1443),
        .dout(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_868 (
        .din(_194_),
        .dout(new_Jinkela_wire_1207)
    );

    spl2 new_Jinkela_splitter_141 (
        .a(new_Jinkela_wire_1444),
        .b(new_Jinkela_wire_1445),
        .c(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_112),
        .dout(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_779),
        .dout(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_773),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_770),
        .dout(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_126),
        .b(new_Jinkela_wire_127),
        .c(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    spl2 new_Jinkela_splitter_106 (
        .a(_103_),
        .b(new_Jinkela_wire_787),
        .c(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    spl2 new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_169),
        .b(new_Jinkela_wire_170),
        .c(new_Jinkela_wire_171)
    );

    spl3L new_Jinkela_splitter_107 (
        .a(_102_),
        .b(new_Jinkela_wire_805),
        .c(new_Jinkela_wire_806),
        .d(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_107 (
        .din(N126),
        .dout(new_Jinkela_wire_180)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_775),
        .dout(new_Jinkela_wire_776)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_142),
        .dout(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_776),
        .dout(new_Jinkela_wire_777)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(new_Jinkela_wire_132),
        .b(new_Jinkela_wire_133),
        .c(new_Jinkela_wire_134)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    spl2 new_Jinkela_splitter_30 (
        .a(N8),
        .b(new_Jinkela_wire_192),
        .c(new_Jinkela_wire_193)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    spl3L new_Jinkela_splitter_27 (
        .a(N106),
        .b(new_Jinkela_wire_167),
        .c(new_Jinkela_wire_168),
        .d(new_Jinkela_wire_169)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(_047_),
        .b(new_Jinkela_wire_825),
        .c(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_180),
        .dout(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    spl3L new_Jinkela_splitter_31 (
        .a(N96),
        .b(new_Jinkela_wire_194),
        .c(new_Jinkela_wire_195),
        .d(new_Jinkela_wire_196)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_172),
        .dout(new_Jinkela_wire_173)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(new_Jinkela_wire_154),
        .b(new_Jinkela_wire_155),
        .c(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    spl2 new_Jinkela_splitter_33 (
        .a(N17),
        .b(new_Jinkela_wire_207),
        .c(new_Jinkela_wire_211)
    );

    spl2 new_Jinkela_splitter_109 (
        .a(_252_),
        .b(new_Jinkela_wire_828),
        .c(new_Jinkela_wire_829)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_173),
        .dout(new_Jinkela_wire_174)
    );

    and_bi _333_ (
        .a(_030_),
        .b(_032_),
        .c(_033_)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_157),
        .dout(new_Jinkela_wire_158)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_791),
        .dout(new_Jinkela_wire_792)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_1715),
        .dout(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(_001_),
        .dout(new_Jinkela_wire_1730)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_1716),
        .dout(new_Jinkela_wire_1717)
    );

    spl3L new_Jinkela_splitter_168 (
        .a(_067_),
        .b(new_Jinkela_wire_1732),
        .c(new_Jinkela_wire_1733),
        .d(new_Jinkela_wire_1734)
    );

    spl2 new_Jinkela_splitter_169 (
        .a(_283_),
        .b(new_Jinkela_wire_1735),
        .c(new_Jinkela_wire_1736)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_1717),
        .dout(new_Jinkela_wire_1718)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_1730),
        .dout(new_Jinkela_wire_1731)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(_021_),
        .dout(new_Jinkela_wire_1737)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_1741),
        .dout(new_Jinkela_wire_1742)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(_136_),
        .dout(new_Jinkela_wire_1744)
    );

    spl4L new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_1737),
        .b(new_Jinkela_wire_1738),
        .c(new_Jinkela_wire_1739),
        .d(new_Jinkela_wire_1740),
        .e(new_Jinkela_wire_1741)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(_123_),
        .dout(new_Jinkela_wire_1745)
    );

    spl3L new_Jinkela_splitter_171 (
        .a(_055_),
        .b(new_Jinkela_wire_1766),
        .c(new_Jinkela_wire_1767),
        .d(new_Jinkela_wire_1768)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_net_536),
        .dout(new_Jinkela_wire_1769)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_1745),
        .dout(new_Jinkela_wire_1746)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_1742),
        .dout(new_Jinkela_wire_1743)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_net_560),
        .dout(new_Jinkela_wire_1804)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_1746),
        .dout(new_Jinkela_wire_1747)
    );

    and_bi _312_ (
        .a(new_Jinkela_wire_208),
        .b(new_Jinkela_wire_3),
        .c(_012_)
    );

    or_ii _290_ (
        .a(new_Jinkela_wire_540),
        .b(new_Jinkela_wire_223),
        .c(_277_)
    );

    and_bi _288_ (
        .a(new_Jinkela_wire_26),
        .b(new_Jinkela_wire_209),
        .c(_275_)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(new_Jinkela_wire_1747),
        .dout(new_Jinkela_wire_1748)
    );

    and_bi _289_ (
        .a(_274_),
        .b(_275_),
        .c(_276_)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_1769),
        .dout(new_Jinkela_wire_1770)
    );

    or_bi _287_ (
        .a(new_Jinkela_wire_27),
        .b(new_Jinkela_wire_213),
        .c(_274_)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_1748),
        .dout(new_Jinkela_wire_1749)
    );

    or_bi _291_ (
        .a(new_Jinkela_wire_994),
        .b(new_Jinkela_wire_422),
        .c(_278_)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_net_544),
        .dout(new_Jinkela_wire_1833)
    );

    inv _295_ (
        .din(new_Jinkela_wire_23),
        .dout(_282_)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(new_Jinkela_wire_1749),
        .dout(new_Jinkela_wire_1750)
    );

    or_bb _294_ (
        .a(_280_),
        .b(new_Jinkela_wire_884),
        .c(_281_)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_1770),
        .dout(new_Jinkela_wire_1771)
    );

    and_bb _292_ (
        .a(new_Jinkela_wire_417),
        .b(new_Jinkela_wire_166),
        .c(_279_)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_1750),
        .dout(new_Jinkela_wire_1751)
    );

    or_bb _304_ (
        .a(new_Jinkela_wire_545),
        .b(new_Jinkela_wire_878),
        .c(_004_)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_1804),
        .dout(new_Jinkela_wire_1805)
    );

    or_bi _293_ (
        .a(new_Jinkela_wire_880),
        .b(new_Jinkela_wire_546),
        .c(_280_)
    );

    or_ii _296_ (
        .a(new_Jinkela_wire_163),
        .b(new_Jinkela_wire_78),
        .c(_283_)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_1751),
        .dout(new_Jinkela_wire_1752)
    );

    or_bb _297_ (
        .a(new_Jinkela_wire_1736),
        .b(new_Jinkela_wire_1661),
        .c(_284_)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_1771),
        .dout(new_Jinkela_wire_1772)
    );

    or_ii _298_ (
        .a(new_Jinkela_wire_420),
        .b(new_Jinkela_wire_214),
        .c(_285_)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_1752),
        .dout(new_Jinkela_wire_1753)
    );

    or_ii _299_ (
        .a(new_Jinkela_wire_193),
        .b(new_Jinkela_wire_224),
        .c(_286_)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(new_net_562),
        .dout(new_Jinkela_wire_1852)
    );

    or_bb _300_ (
        .a(new_Jinkela_wire_627),
        .b(_285_),
        .c(_000_)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_1753),
        .dout(new_Jinkela_wire_1754)
    );

    and_bi _301_ (
        .a(_284_),
        .b(_000_),
        .c(_001_)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_1772),
        .dout(new_Jinkela_wire_1773)
    );

    and_bi _302_ (
        .a(_281_),
        .b(new_Jinkela_wire_1731),
        .c(_002_)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_1754),
        .dout(new_Jinkela_wire_1755)
    );

    or_bi _303_ (
        .a(new_Jinkela_wire_1659),
        .b(new_Jinkela_wire_179),
        .c(_003_)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_1805),
        .dout(new_Jinkela_wire_1806)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_1755),
        .dout(new_Jinkela_wire_1756)
    );

    or_bi _305_ (
        .a(new_Jinkela_wire_1632),
        .b(new_Jinkela_wire_522),
        .c(_005_)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(new_Jinkela_wire_1773),
        .dout(new_Jinkela_wire_1774)
    );

    and_bi _306_ (
        .a(new_Jinkela_wire_19),
        .b(new_Jinkela_wire_2021),
        .c(_006_)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    and_bb _307_ (
        .a(new_Jinkela_wire_409),
        .b(new_Jinkela_wire_438),
        .c(_007_)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_1833),
        .dout(new_Jinkela_wire_1834)
    );

    inv _308_ (
        .din(new_Jinkela_wire_486),
        .dout(_008_)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_1757),
        .dout(new_Jinkela_wire_1758)
    );

    or_ii _309_ (
        .a(new_Jinkela_wire_77),
        .b(new_Jinkela_wire_469),
        .c(_009_)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(new_Jinkela_wire_1774),
        .dout(new_Jinkela_wire_1775)
    );

    or_bb _310_ (
        .a(new_Jinkela_wire_625),
        .b(new_Jinkela_wire_1250),
        .c(_010_)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_Jinkela_wire_1758),
        .dout(new_Jinkela_wire_1759)
    );

    or_bb _311_ (
        .a(new_Jinkela_wire_1728),
        .b(new_Jinkela_wire_877),
        .c(_011_)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(new_Jinkela_wire_1806),
        .dout(new_Jinkela_wire_1807)
    );

endmodule
