module c5315(G124,G52,G48,G72,G100,G110,G53,G80,G132,G91,G55,G99,G134,G121,G61,G37,G165,G39,G157,G5,G62,G105,G117,G16,G44,G18,G96,G168,G36,G3,G43,G6,G78,G12,G42,G88,G57,G8,G137,G128,G153,G54,G118,G93,G169,G87,G73,G50,G174,G101,G67,G126,G103,G158,G161,G86,G138,G68,G113,G108,G140,G97,G135,G65,G92,G56,G66,G9,G112,G171,G64,G13,G142,G69,G14,G4,G150,G106,G109,G145,G139,G131,G160,G119,G159,G19,G11,G94,G120,G83,G123,G89,G152,G136,G46,G146,G32,G85,G47,G95,G114,G81,G45,G30,G111,G176,G148,G51,G162,G63,G149,G156,G155,G144,G1,G26,G102,G70,G17,G147,G129,G15,G24,G31,G141,G172,G49,G41,G84,G166,G20,G143,G107,G154,G122,G90,G77,G125,G82,G29,G74,G130,G164,G38,G10,G76,G116,G133,G35,G40,G7,G115,G177,G2,G104,G127,G27,G173,G60,G22,G21,G23,G170,G71,G98,G34,G33,G163,G59,G75,G167,G175,G28,G58,G79,G151,G178,G25);
    wire new_Jinkela_wire_3194;
    wire new_Jinkela_wire_3818;
    wire _0999_;
    wire new_Jinkela_wire_3971;
    wire new_Jinkela_wire_4255;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_3901;
    wire new_Jinkela_wire_3671;
    wire new_Jinkela_wire_6752;
    wire _0602_;
    wire new_Jinkela_wire_7513;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_2211;
    wire new_Jinkela_wire_2088;
    wire new_Jinkela_wire_4834;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_2406;
    wire new_Jinkela_wire_7288;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_3057;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_7843;
    wire new_Jinkela_wire_7161;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_5376;
    wire new_Jinkela_wire_2238;
    wire _1003_;
    wire new_Jinkela_wire_7324;
    wire _0102_;
    wire new_Jinkela_wire_3065;
    wire new_Jinkela_wire_4696;
    wire new_Jinkela_wire_6142;
    wire new_Jinkela_wire_7387;
    wire new_Jinkela_wire_4857;
    wire _0358_;
    wire _0910_;
    wire new_Jinkela_wire_4129;
    wire _0632_;
    wire new_Jinkela_wire_5959;
    wire new_Jinkela_wire_7954;
    wire new_Jinkela_wire_7703;
    wire _0963_;
    wire _1047_;
    wire new_Jinkela_wire_4161;
    wire _0330_;
    wire new_Jinkela_wire_3891;
    wire new_Jinkela_wire_7685;
    wire new_Jinkela_wire_4966;
    wire _1002_;
    wire new_Jinkela_wire_6740;
    wire new_Jinkela_wire_5421;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_2441;
    wire new_Jinkela_wire_7028;
    wire new_Jinkela_wire_2326;
    wire new_Jinkela_wire_5619;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_4796;
    wire new_Jinkela_wire_3529;
    wire _1182_;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_6681;
    wire new_Jinkela_wire_3134;
    wire new_Jinkela_wire_2150;
    wire _0085_;
    wire new_Jinkela_wire_3904;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_5414;
    wire new_Jinkela_wire_7791;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_2260;
    wire new_Jinkela_wire_5546;
    wire new_Jinkela_wire_6926;
    wire new_Jinkela_wire_6595;
    wire new_Jinkela_wire_5199;
    wire new_Jinkela_wire_1391;
    wire new_Jinkela_wire_5947;
    wire new_Jinkela_wire_2470;
    wire _0665_;
    wire _1108_;
    wire new_Jinkela_wire_3219;
    wire _0125_;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_1529;
    wire _0335_;
    wire new_Jinkela_wire_2420;
    wire new_Jinkela_wire_6490;
    wire new_Jinkela_wire_5768;
    wire _0553_;
    wire new_Jinkela_wire_5192;
    wire new_Jinkela_wire_5932;
    wire new_Jinkela_wire_5746;
    wire new_Jinkela_wire_7555;
    wire _1228_;
    wire _0930_;
    wire new_Jinkela_wire_6038;
    wire new_Jinkela_wire_4185;
    wire new_Jinkela_wire_3802;
    wire new_Jinkela_wire_1424;
    wire _0582_;
    wire new_Jinkela_wire_7020;
    wire new_Jinkela_wire_1135;
    wire _1097_;
    wire _0512_;
    wire new_Jinkela_wire_5057;
    wire new_Jinkela_wire_2722;
    wire new_Jinkela_wire_3200;
    wire new_Jinkela_wire_371;
    wire _0570_;
    wire new_Jinkela_wire_4150;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_5307;
    wire _0296_;
    wire new_Jinkela_wire_1719;
    wire new_Jinkela_wire_4401;
    wire new_Jinkela_wire_3147;
    wire _0497_;
    wire new_Jinkela_wire_6951;
    wire _0679_;
    wire new_Jinkela_wire_7955;
    wire new_Jinkela_wire_3613;
    wire new_Jinkela_wire_6512;
    wire new_Jinkela_wire_3854;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_7284;
    wire new_Jinkela_wire_6145;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_7330;
    wire new_Jinkela_wire_1975;
    wire new_Jinkela_wire_4659;
    wire new_Jinkela_wire_7167;
    wire _0710_;
    wire new_Jinkela_wire_5170;
    wire new_Jinkela_wire_3600;
    wire _0233_;
    wire new_Jinkela_wire_2098;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_1197;
    wire _0800_;
    wire new_Jinkela_wire_2807;
    wire new_Jinkela_wire_6665;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_5125;
    wire new_Jinkela_wire_5067;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_5339;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_1407;
    wire _0718_;
    wire new_Jinkela_wire_5061;
    wire new_Jinkela_wire_2997;
    wire new_Jinkela_wire_4557;
    wire new_Jinkela_wire_4866;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_5741;
    wire _0000_;
    wire new_Jinkela_wire_3846;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_5422;
    wire new_Jinkela_wire_2052;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_3329;
    wire new_Jinkela_wire_5457;
    wire new_Jinkela_wire_4041;
    wire new_Jinkela_wire_1138;
    wire _0547_;
    wire new_Jinkela_wire_2842;
    wire _0225_;
    wire new_Jinkela_wire_7612;
    wire new_Jinkela_wire_2382;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_6293;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_6498;
    wire new_Jinkela_wire_1063;
    wire _0707_;
    wire new_Jinkela_wire_5740;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_1684;
    wire _0871_;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_5017;
    wire new_Jinkela_wire_2730;
    wire new_Jinkela_wire_7663;
    wire _0896_;
    wire new_Jinkela_wire_4208;
    wire new_Jinkela_wire_6747;
    wire new_Jinkela_wire_2119;
    wire new_Jinkela_wire_6638;
    wire new_Jinkela_wire_4215;
    wire new_Jinkela_wire_4016;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_4535;
    wire new_Jinkela_wire_3425;
    wire new_Jinkela_wire_4621;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_4376;
    wire new_Jinkela_wire_3341;
    wire new_Jinkela_wire_3544;
    wire new_Jinkela_wire_2060;
    wire new_Jinkela_wire_5858;
    wire _1152_;
    wire _0897_;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_6278;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_4063;
    wire new_Jinkela_wire_3070;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_5528;
    wire new_Jinkela_wire_1688;
    wire new_Jinkela_wire_2284;
    wire new_Jinkela_wire_3589;
    wire _0969_;
    wire new_Jinkela_wire_2855;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_7952;
    wire new_Jinkela_wire_4229;
    wire new_Jinkela_wire_4598;
    wire new_Jinkela_wire_2237;
    wire _0484_;
    wire _0962_;
    wire new_Jinkela_wire_3718;
    wire new_Jinkela_wire_5925;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_6292;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_5163;
    wire new_Jinkela_wire_7373;
    wire new_Jinkela_wire_6499;
    wire new_Jinkela_wire_3397;
    wire new_Jinkela_wire_3936;
    wire _0086_;
    wire new_Jinkela_wire_6961;
    wire new_Jinkela_wire_6806;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_2801;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_5618;
    wire new_Jinkela_wire_3071;
    wire _1179_;
    wire new_Jinkela_wire_4868;
    wire new_Jinkela_wire_4685;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_2991;
    wire new_Jinkela_wire_7355;
    wire new_Jinkela_wire_7894;
    wire new_Jinkela_wire_4408;
    wire new_Jinkela_wire_4904;
    wire new_Jinkela_wire_4246;
    wire new_Jinkela_wire_634;
    wire _1160_;
    wire new_Jinkela_wire_3098;
    wire new_Jinkela_wire_4540;
    wire new_Jinkela_wire_4144;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_1223;
    wire _0244_;
    wire new_Jinkela_wire_3393;
    wire new_Jinkela_wire_7903;
    wire new_Jinkela_wire_7302;
    wire new_Jinkela_wire_1344;
    wire _0678_;
    wire new_Jinkela_wire_7047;
    wire new_Jinkela_wire_4056;
    wire new_Jinkela_wire_6291;
    wire new_Jinkela_wire_4649;
    wire _1017_;
    wire new_Jinkela_wire_3114;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_3842;
    wire new_Jinkela_wire_4234;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_7133;
    wire new_Jinkela_wire_6947;
    wire new_Jinkela_wire_2322;
    wire _0481_;
    wire new_Jinkela_wire_2469;
    wire new_Jinkela_wire_4681;
    wire _0739_;
    wire new_Jinkela_wire_2454;
    wire new_Jinkela_wire_7365;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_4320;
    wire new_Jinkela_wire_5312;
    wire _0077_;
    wire new_Jinkela_wire_5972;
    wire new_Jinkela_wire_3812;
    wire _0677_;
    wire new_Jinkela_wire_2396;
    wire new_Jinkela_wire_7262;
    wire new_Jinkela_wire_4998;
    wire new_Jinkela_wire_4459;
    wire new_Jinkela_wire_5101;
    wire new_Jinkela_wire_2825;
    wire new_Jinkela_wire_4521;
    wire new_Jinkela_wire_4570;
    wire new_Jinkela_wire_6267;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_5096;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_1066;
    wire new_Jinkela_wire_7958;
    wire new_Jinkela_wire_3451;
    wire new_Jinkela_wire_7606;
    wire new_Jinkela_wire_6779;
    wire new_Jinkela_wire_6721;
    wire new_Jinkela_wire_2712;
    wire new_Jinkela_wire_3701;
    wire new_Jinkela_wire_4140;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_4077;
    wire new_Jinkela_wire_7379;
    wire new_Jinkela_wire_6639;
    wire new_Jinkela_wire_546;
    wire _0367_;
    wire new_Jinkela_wire_4413;
    wire new_Jinkela_wire_2115;
    wire new_Jinkela_wire_6226;
    wire new_Jinkela_wire_5808;
    wire new_Jinkela_wire_3806;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_4292;
    wire new_Jinkela_wire_4672;
    wire new_Jinkela_wire_4261;
    wire new_Jinkela_wire_2571;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_3551;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_7548;
    wire new_Jinkela_wire_2191;
    wire new_Jinkela_wire_7928;
    wire new_Jinkela_wire_5789;
    wire _0067_;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_7421;
    wire _0538_;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_5543;
    wire _0138_;
    wire new_Jinkela_wire_1137;
    wire _0033_;
    wire new_Jinkela_wire_5420;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_5160;
    wire new_Jinkela_wire_5521;
    wire _1091_;
    wire new_Jinkela_wire_2848;
    wire new_Jinkela_wire_2346;
    wire new_Jinkela_wire_5031;
    wire new_Jinkela_wire_4135;
    wire _1122_;
    wire new_Jinkela_wire_2437;
    wire _0089_;
    wire new_Jinkela_wire_6044;
    wire new_Jinkela_wire_3950;
    wire new_Jinkela_wire_5319;
    wire _1055_;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_5169;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_2733;
    wire new_Jinkela_wire_3485;
    wire new_Jinkela_wire_3889;
    wire new_Jinkela_wire_5729;
    wire new_Jinkela_wire_6000;
    wire new_Jinkela_wire_4537;
    wire new_Jinkela_wire_3832;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_4004;
    wire _0514_;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_1543;
    wire _0082_;
    wire new_Jinkela_wire_4744;
    wire new_Jinkela_wire_2566;
    wire _0886_;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_5703;
    wire new_Jinkela_wire_4190;
    wire new_Jinkela_wire_2934;
    wire new_Jinkela_wire_5301;
    wire new_Jinkela_wire_4677;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_4624;
    wire new_Jinkela_wire_6801;
    wire new_Jinkela_wire_4117;
    wire new_Jinkela_wire_3512;
    wire new_Jinkela_wire_3312;
    wire new_Jinkela_wire_6256;
    wire new_Jinkela_wire_6616;
    wire new_Jinkela_wire_7801;
    wire new_Jinkela_wire_5187;
    wire _0157_;
    wire new_Jinkela_wire_4163;
    wire _0375_;
    wire new_Jinkela_wire_2085;
    wire new_Jinkela_wire_7580;
    wire new_Jinkela_wire_2367;
    wire new_Jinkela_wire_4584;
    wire new_Jinkela_wire_7214;
    wire new_Jinkela_wire_7804;
    wire _1070_;
    wire new_Jinkela_wire_4829;
    wire new_Jinkela_wire_2767;
    wire new_Jinkela_wire_6826;
    wire new_Jinkela_wire_1433;
    wire _0479_;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_2700;
    wire new_Jinkela_wire_6620;
    wire new_Jinkela_wire_6227;
    wire new_Jinkela_wire_2906;
    wire new_Jinkela_wire_6214;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_5527;
    wire new_Jinkela_wire_3256;
    wire new_Jinkela_wire_3669;
    wire new_Jinkela_wire_2553;
    wire new_Jinkela_wire_3882;
    wire new_Jinkela_wire_121;
    wire new_Jinkela_wire_7090;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_7834;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_2615;
    wire new_Jinkela_wire_2010;
    wire new_Jinkela_wire_6999;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_6010;
    wire new_Jinkela_wire_6184;
    wire new_Jinkela_wire_2698;
    wire _0377_;
    wire new_Jinkela_wire_5415;
    wire _0217_;
    wire new_Jinkela_wire_6982;
    wire _0573_;
    wire new_Jinkela_wire_7417;
    wire new_Jinkela_wire_2389;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_2465;
    wire _0539_;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_7235;
    wire new_Jinkela_wire_5398;
    wire new_Jinkela_wire_4491;
    wire new_Jinkela_wire_5616;
    wire new_Jinkela_wire_7113;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_6825;
    wire _0214_;
    wire new_Jinkela_wire_7873;
    wire _1107_;
    wire new_Jinkela_wire_5786;
    wire new_Jinkela_wire_5188;
    wire new_Jinkela_wire_7514;
    wire new_Jinkela_wire_6500;
    wire new_net_2445;
    wire new_Jinkela_wire_5000;
    wire new_Jinkela_wire_1816;
    wire new_Jinkela_wire_2575;
    wire new_net_2399;
    wire new_Jinkela_wire_2783;
    wire new_Jinkela_wire_3448;
    wire new_Jinkela_wire_2231;
    wire new_Jinkela_wire_3568;
    wire new_Jinkela_wire_4762;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_4010;
    wire new_Jinkela_wire_4417;
    wire _0549_;
    wire _0320_;
    wire new_Jinkela_wire_2266;
    wire _0590_;
    wire new_Jinkela_wire_3902;
    wire new_Jinkela_wire_3516;
    wire new_Jinkela_wire_2853;
    wire new_Jinkela_wire_5634;
    wire new_Jinkela_wire_5943;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_2797;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_2961;
    wire new_net_2447;
    wire _0882_;
    wire new_Jinkela_wire_7937;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_2256;
    wire new_Jinkela_wire_2585;
    wire new_net_6;
    wire _0879_;
    wire new_Jinkela_wire_3010;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_6091;
    wire new_Jinkela_wire_3655;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_3595;
    wire new_Jinkela_wire_6054;
    wire new_Jinkela_wire_5751;
    wire new_Jinkela_wire_4840;
    wire new_Jinkela_wire_6530;
    wire new_Jinkela_wire_3089;
    wire _0624_;
    wire new_Jinkela_wire_6344;
    wire new_Jinkela_wire_6406;
    wire _1151_;
    wire new_Jinkela_wire_5699;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_7504;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_4390;
    wire new_Jinkela_wire_621;
    wire _0420_;
    wire _1086_;
    wire new_Jinkela_wire_6992;
    wire new_Jinkela_wire_3355;
    wire new_Jinkela_wire_5919;
    wire new_Jinkela_wire_4506;
    wire _0183_;
    wire new_Jinkela_wire_5928;
    wire new_Jinkela_wire_5791;
    wire new_Jinkela_wire_3153;
    wire new_Jinkela_wire_5320;
    wire _0636_;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_7033;
    wire new_Jinkela_wire_6332;
    wire new_Jinkela_wire_6920;
    wire new_Jinkela_wire_7150;
    wire new_Jinkela_wire_2213;
    wire new_Jinkela_wire_4201;
    wire new_Jinkela_wire_3831;
    wire new_Jinkela_wire_1746;
    wire new_Jinkela_wire_4580;
    wire new_Jinkela_wire_6763;
    wire new_Jinkela_wire_3513;
    wire new_Jinkela_wire_2732;
    wire _0179_;
    wire _1062_;
    wire new_Jinkela_wire_5733;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_7016;
    wire new_Jinkela_wire_6549;
    wire new_Jinkela_wire_3502;
    wire new_Jinkela_wire_6407;
    wire new_Jinkela_wire_7303;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_4897;
    wire new_Jinkela_wire_149;
    wire _0419_;
    wire new_Jinkela_wire_5084;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_5735;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_5282;
    wire new_Jinkela_wire_4082;
    wire new_Jinkela_wire_2208;
    wire new_Jinkela_wire_2354;
    wire new_Jinkela_wire_2412;
    wire new_Jinkela_wire_3640;
    wire new_Jinkela_wire_6212;
    wire new_Jinkela_wire_6160;
    wire new_Jinkela_wire_3099;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_6334;
    wire _0083_;
    wire new_Jinkela_wire_7900;
    wire new_Jinkela_wire_962;
    wire _0502_;
    wire _0047_;
    wire new_Jinkela_wire_5284;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_2724;
    wire new_Jinkela_wire_5820;
    wire new_Jinkela_wire_6847;
    wire new_Jinkela_wire_5900;
    wire new_Jinkela_wire_2246;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_5370;
    wire _0396_;
    wire new_Jinkela_wire_5926;
    wire new_Jinkela_wire_3570;
    wire new_Jinkela_wire_5046;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_2480;
    wire _1112_;
    wire new_Jinkela_wire_4937;
    wire new_Jinkela_wire_4591;
    wire new_Jinkela_wire_3009;
    wire _1233_;
    wire new_Jinkela_wire_4489;
    wire new_Jinkela_wire_1553;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_1717;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_7240;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_6172;
    wire _0506_;
    wire new_Jinkela_wire_4926;
    wire new_Jinkela_wire_4250;
    wire _0297_;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_7024;
    wire new_Jinkela_wire_4574;
    wire new_Jinkela_wire_6247;
    wire new_Jinkela_wire_2756;
    wire _1095_;
    wire new_Jinkela_wire_5222;
    wire _1010_;
    wire new_Jinkela_wire_3770;
    wire _0595_;
    wire new_Jinkela_wire_16;
    wire _0469_;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_2075;
    wire new_Jinkela_wire_6892;
    wire new_Jinkela_wire_2004;
    wire new_Jinkela_wire_5128;
    wire new_Jinkela_wire_4976;
    wire new_Jinkela_wire_7500;
    wire new_Jinkela_wire_6325;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_2262;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_4346;
    wire new_Jinkela_wire_4361;
    wire new_Jinkela_wire_7925;
    wire new_Jinkela_wire_4472;
    wire new_Jinkela_wire_4406;
    wire new_Jinkela_wire_7883;
    wire new_Jinkela_wire_6520;
    wire new_Jinkela_wire_7265;
    wire new_Jinkela_wire_6663;
    wire new_Jinkela_wire_2775;
    wire new_Jinkela_wire_4699;
    wire new_Jinkela_wire_6524;
    wire new_Jinkela_wire_6389;
    wire new_Jinkela_wire_2443;
    wire new_Jinkela_wire_2236;
    wire _0977_;
    wire _0104_;
    wire new_Jinkela_wire_6359;
    wire _0192_;
    wire new_Jinkela_wire_5162;
    wire new_Jinkela_wire_3479;
    wire new_Jinkela_wire_6294;
    wire new_Jinkela_wire_4562;
    wire _0013_;
    wire new_Jinkela_wire_6137;
    wire new_net_2479;
    wire new_Jinkela_wire_3171;
    wire new_Jinkela_wire_5732;
    wire new_Jinkela_wire_4171;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_3441;
    wire new_Jinkela_wire_3539;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_6244;
    wire new_Jinkela_wire_4872;
    wire new_Jinkela_wire_1486;
    wire new_net_2495;
    wire new_Jinkela_wire_2380;
    wire new_Jinkela_wire_1724;
    wire new_Jinkela_wire_7468;
    wire new_Jinkela_wire_7129;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_1763;
    wire new_Jinkela_wire_4929;
    wire new_Jinkela_wire_4298;
    wire new_Jinkela_wire_6144;
    wire new_Jinkela_wire_1818;
    wire new_Jinkela_wire_6889;
    wire _0004_;
    wire new_Jinkela_wire_3838;
    wire new_Jinkela_wire_3628;
    wire new_Jinkela_wire_5906;
    wire new_Jinkela_wire_5835;
    wire new_Jinkela_wire_2784;
    wire new_Jinkela_wire_5574;
    wire new_Jinkela_wire_2777;
    wire new_Jinkela_wire_7710;
    wire new_Jinkela_wire_2157;
    wire new_Jinkela_wire_3795;
    wire new_Jinkela_wire_4893;
    wire _0744_;
    wire _0359_;
    wire new_Jinkela_wire_4869;
    wire _0322_;
    wire new_Jinkela_wire_3689;
    wire new_Jinkela_wire_5621;
    wire new_Jinkela_wire_4882;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_6174;
    wire new_Jinkela_wire_5438;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_4991;
    wire new_Jinkela_wire_1785;
    wire new_Jinkela_wire_3498;
    wire new_Jinkela_wire_5086;
    wire new_Jinkela_wire_4029;
    wire _0639_;
    wire new_Jinkela_wire_2563;
    wire new_Jinkela_wire_4365;
    wire new_Jinkela_wire_6822;
    wire _0018_;
    wire new_Jinkela_wire_7680;
    wire new_Jinkela_wire_3111;
    wire new_Jinkela_wire_2110;
    wire new_Jinkela_wire_7799;
    wire new_Jinkela_wire_4312;
    wire new_Jinkela_wire_3093;
    wire new_Jinkela_wire_3173;
    wire _1094_;
    wire new_Jinkela_wire_5709;
    wire new_Jinkela_wire_7847;
    wire new_Jinkela_wire_4090;
    wire new_Jinkela_wire_5579;
    wire new_Jinkela_wire_4735;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_7316;
    wire new_Jinkela_wire_4539;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_6434;
    wire _1225_;
    wire new_Jinkela_wire_4107;
    wire new_Jinkela_wire_4616;
    wire new_Jinkela_wire_4416;
    wire _0950_;
    wire _0486_;
    wire new_Jinkela_wire_5006;
    wire _0603_;
    wire new_Jinkela_wire_1704;
    wire _0968_;
    wire new_Jinkela_wire_1874;
    wire _1244_;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_3986;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_861;
    wire _0445_;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_1973;
    wire new_Jinkela_wire_5153;
    wire new_Jinkela_wire_4855;
    wire new_Jinkela_wire_6324;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_5043;
    wire new_Jinkela_wire_3365;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_780;
    wire _0835_;
    wire new_Jinkela_wire_2109;
    wire new_Jinkela_wire_2919;
    wire _0429_;
    wire new_Jinkela_wire_2081;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_7208;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_6328;
    wire new_Jinkela_wire_5738;
    wire new_Jinkela_wire_2694;
    wire new_net_2387;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_4597;
    wire new_Jinkela_wire_6109;
    wire new_Jinkela_wire_6372;
    wire new_Jinkela_wire_5164;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_2493;
    wire new_Jinkela_wire_4963;
    wire new_Jinkela_wire_2764;
    wire new_Jinkela_wire_2370;
    wire new_Jinkela_wire_7796;
    wire new_Jinkela_wire_7109;
    wire new_Jinkela_wire_7947;
    wire new_Jinkela_wire_3656;
    wire new_Jinkela_wire_7456;
    wire new_Jinkela_wire_2979;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_6350;
    wire new_Jinkela_wire_4484;
    wire _0491_;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_4345;
    wire new_Jinkela_wire_1506;
    wire new_Jinkela_wire_6249;
    wire new_Jinkela_wire_3712;
    wire new_Jinkela_wire_5366;
    wire new_Jinkela_wire_7931;
    wire new_Jinkela_wire_4799;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_1579;
    wire _0411_;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_7312;
    wire _1085_;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_7072;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_7872;
    wire new_Jinkela_wire_6983;
    wire new_Jinkela_wire_4726;
    wire new_Jinkela_wire_5981;
    wire new_Jinkela_wire_1870;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_7593;
    wire _0904_;
    wire new_Jinkela_wire_6331;
    wire new_Jinkela_wire_7359;
    wire new_Jinkela_wire_2083;
    wire new_Jinkela_wire_2632;
    wire new_Jinkela_wire_7413;
    wire new_Jinkela_wire_6546;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_3016;
    wire new_Jinkela_wire_4668;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_7082;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_3003;
    wire _0846_;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_79;
    wire _0574_;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_2856;
    wire new_Jinkela_wire_5558;
    wire new_Jinkela_wire_5220;
    wire new_Jinkela_wire_264;
    wire _0474_;
    wire new_Jinkela_wire_4614;
    wire new_Jinkela_wire_3972;
    wire new_Jinkela_wire_3104;
    wire new_Jinkela_wire_6139;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_5201;
    wire new_Jinkela_wire_3264;
    wire new_Jinkela_wire_3182;
    wire _0154_;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_1978;
    wire new_Jinkela_wire_5119;
    wire new_Jinkela_wire_3116;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_925;
    wire _1050_;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_4545;
    wire _0313_;
    wire new_Jinkela_wire_5394;
    wire new_Jinkela_wire_3992;
    wire _1117_;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_5922;
    wire _0412_;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_7876;
    wire new_Jinkela_wire_6573;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_4658;
    wire new_Jinkela_wire_6009;
    wire new_Jinkela_wire_3785;
    wire new_Jinkela_wire_5285;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_4674;
    wire new_Jinkela_wire_2725;
    wire new_Jinkela_wire_4881;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_2434;
    wire new_Jinkela_wire_6804;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_6705;
    wire new_Jinkela_wire_4262;
    wire new_Jinkela_wire_2495;
    wire new_Jinkela_wire_6251;
    wire new_Jinkela_wire_3186;
    wire new_Jinkela_wire_3119;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_2435;
    wire _0144_;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_4048;
    wire new_Jinkela_wire_6486;
    wire new_Jinkela_wire_7248;
    wire _0522_;
    wire new_Jinkela_wire_4723;
    wire new_Jinkela_wire_7358;
    wire new_Jinkela_wire_5765;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_1643;
    wire _0070_;
    wire new_Jinkela_wire_5409;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_7757;
    wire new_Jinkela_wire_1802;
    wire _1118_;
    wire _1029_;
    wire new_net_14;
    wire new_Jinkela_wire_3781;
    wire new_Jinkela_wire_3156;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_5123;
    wire new_Jinkela_wire_6361;
    wire new_Jinkela_wire_2537;
    wire new_Jinkela_wire_2520;
    wire new_Jinkela_wire_7228;
    wire _0966_;
    wire new_Jinkela_wire_2499;
    wire new_Jinkela_wire_5231;
    wire new_Jinkela_wire_4152;
    wire new_Jinkela_wire_7226;
    wire new_Jinkela_wire_4480;
    wire new_Jinkela_wire_5186;
    wire new_Jinkela_wire_1896;
    wire new_Jinkela_wire_5855;
    wire new_Jinkela_wire_3996;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_3927;
    wire new_Jinkela_wire_3653;
    wire new_Jinkela_wire_7636;
    wire new_Jinkela_wire_7348;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_7326;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_6141;
    wire new_Jinkela_wire_7467;
    wire new_Jinkela_wire_6572;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_7634;
    wire new_Jinkela_wire_2514;
    wire new_Jinkela_wire_1867;
    wire new_Jinkela_wire_2788;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_7671;
    wire _0232_;
    wire new_Jinkela_wire_6208;
    wire new_Jinkela_wire_5271;
    wire new_Jinkela_wire_5005;
    wire new_Jinkela_wire_4711;
    wire new_Jinkela_wire_3251;
    wire new_Jinkela_wire_6697;
    wire new_Jinkela_wire_6559;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_3768;
    wire new_Jinkela_wire_7192;
    wire new_Jinkela_wire_7157;
    wire new_Jinkela_wire_4751;
    wire _0374_;
    wire new_Jinkela_wire_7095;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_4617;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_6495;
    wire _0808_;
    wire _1172_;
    wire new_Jinkela_wire_4563;
    wire new_Jinkela_wire_6896;
    wire new_Jinkela_wire_3951;
    wire new_Jinkela_wire_3097;
    wire new_Jinkela_wire_5180;
    wire new_Jinkela_wire_2933;
    wire new_Jinkela_wire_2505;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_4436;
    wire _0610_;
    wire _0309_;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_3303;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_2820;
    wire new_Jinkela_wire_5931;
    wire _0720_;
    wire new_Jinkela_wire_7785;
    wire new_Jinkela_wire_3232;
    wire new_Jinkela_wire_2428;
    wire new_Jinkela_wire_5830;
    wire new_Jinkela_wire_7124;
    wire new_Jinkela_wire_4139;
    wire _1208_;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_3298;
    wire new_Jinkela_wire_5853;
    wire new_Jinkela_wire_4070;
    wire new_Jinkela_wire_3617;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_6772;
    wire new_Jinkela_wire_6408;
    wire new_Jinkela_wire_7592;
    wire new_Jinkela_wire_3541;
    wire new_Jinkela_wire_7516;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_5690;
    wire new_Jinkela_wire_6527;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_7048;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_2135;
    wire new_Jinkela_wire_52;
    wire _0141_;
    wire new_Jinkela_wire_4898;
    wire new_Jinkela_wire_3923;
    wire new_Jinkela_wire_4729;
    wire new_Jinkela_wire_7022;
    wire new_Jinkela_wire_5713;
    wire new_Jinkela_wire_2096;
    wire new_Jinkela_wire_6603;
    wire new_Jinkela_wire_5068;
    wire new_Jinkela_wire_3857;
    wire _0441_;
    wire new_Jinkela_wire_6412;
    wire _0177_;
    wire new_Jinkela_wire_3885;
    wire new_Jinkela_wire_5179;
    wire new_Jinkela_wire_6686;
    wire new_Jinkela_wire_2444;
    wire new_Jinkela_wire_2449;
    wire new_Jinkela_wire_8008;
    wire _0090_;
    wire new_Jinkela_wire_4803;
    wire new_Jinkela_wire_2929;
    wire new_Jinkela_wire_4172;
    wire new_Jinkela_wire_7988;
    wire new_Jinkela_wire_6410;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_3348;
    wire new_Jinkela_wire_5352;
    wire _0096_;
    wire new_Jinkela_wire_2630;
    wire new_Jinkela_wire_3405;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_7394;
    wire new_Jinkela_wire_7776;
    wire _0619_;
    wire new_Jinkela_wire_2393;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_5911;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_5514;
    wire _1101_;
    wire new_Jinkela_wire_4801;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_7408;
    wire new_Jinkela_wire_3732;
    wire new_Jinkela_wire_4941;
    wire new_Jinkela_wire_4817;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_5007;
    wire new_Jinkela_wire_3565;
    wire new_Jinkela_wire_7345;
    wire new_Jinkela_wire_7861;
    wire new_Jinkela_wire_2587;
    wire new_Jinkela_wire_5599;
    wire new_Jinkela_wire_4514;
    wire new_Jinkela_wire_6827;
    wire new_Jinkela_wire_5877;
    wire new_Jinkela_wire_3518;
    wire _1042_;
    wire new_Jinkela_wire_6924;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_6810;
    wire new_Jinkela_wire_2050;
    wire new_Jinkela_wire_7868;
    wire new_Jinkela_wire_2699;
    wire new_Jinkela_wire_5161;
    wire new_Jinkela_wire_3978;
    wire new_Jinkela_wire_6797;
    wire _0855_;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_7575;
    wire new_Jinkela_wire_4733;
    wire new_Jinkela_wire_6276;
    wire _0927_;
    wire _0294_;
    wire new_Jinkela_wire_6736;
    wire new_Jinkela_wire_161;
    wire _0695_;
    wire new_Jinkela_wire_1865;
    wire new_Jinkela_wire_5622;
    wire new_Jinkela_wire_4967;
    wire new_Jinkela_wire_5552;
    wire new_Jinkela_wire_2292;
    wire new_Jinkela_wire_4671;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_4605;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_4464;
    wire new_Jinkela_wire_4612;
    wire _0216_;
    wire _1212_;
    wire _0443_;
    wire new_Jinkela_wire_3500;
    wire new_Jinkela_wire_6948;
    wire new_Jinkela_wire_5433;
    wire new_Jinkela_wire_4774;
    wire new_Jinkela_wire_4510;
    wire new_net_11;
    wire _0028_;
    wire _0115_;
    wire _0751_;
    wire new_Jinkela_wire_2242;
    wire _0120_;
    wire new_Jinkela_wire_5263;
    wire new_Jinkela_wire_4323;
    wire new_Jinkela_wire_5615;
    wire new_Jinkela_wire_7173;
    wire new_Jinkela_wire_6202;
    wire new_Jinkela_wire_7684;
    wire new_Jinkela_wire_6734;
    wire _0593_;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_4211;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_4529;
    wire new_net_2441;
    wire new_Jinkela_wire_2198;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_2359;
    wire new_Jinkela_wire_7705;
    wire new_Jinkela_wire_6209;
    wire new_Jinkela_wire_5365;
    wire new_Jinkela_wire_7209;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_2810;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_6221;
    wire new_Jinkela_wire_2460;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_2492;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_597;
    wire _0865_;
    wire new_Jinkela_wire_6991;
    wire new_Jinkela_wire_3414;
    wire new_Jinkela_wire_4118;
    wire new_Jinkela_wire_4708;
    wire new_Jinkela_wire_6436;
    wire new_Jinkela_wire_5501;
    wire _0448_;
    wire new_Jinkela_wire_4372;
    wire new_Jinkela_wire_4609;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_178;
    wire new_Jinkela_wire_2545;
    wire new_Jinkela_wire_7012;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_4714;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_5261;
    wire new_Jinkela_wire_5467;
    wire new_Jinkela_wire_6477;
    wire new_Jinkela_wire_4531;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_4304;
    wire new_Jinkela_wire_2409;
    wire _0114_;
    wire _0392_;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_6450;
    wire new_Jinkela_wire_5435;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_86;
    wire _0622_;
    wire new_Jinkela_wire_3249;
    wire new_Jinkela_wire_1086;
    wire new_Jinkela_wire_3720;
    wire new_Jinkela_wire_7913;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_5568;
    wire _1032_;
    wire new_Jinkela_wire_3383;
    wire new_Jinkela_wire_2288;
    wire new_Jinkela_wire_7865;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_4600;
    wire new_Jinkela_wire_5566;
    wire new_Jinkela_wire_6316;
    wire _1153_;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_516;
    wire _0385_;
    wire new_Jinkela_wire_3404;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_6861;
    wire _0023_;
    wire new_Jinkela_wire_6015;
    wire _0031_;
    wire new_Jinkela_wire_6859;
    wire new_Jinkela_wire_3288;
    wire new_Jinkela_wire_4702;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_7026;
    wire new_Jinkela_wire_7013;
    wire _0750_;
    wire new_Jinkela_wire_1709;
    wire new_Jinkela_wire_5032;
    wire new_Jinkela_wire_2653;
    wire new_Jinkela_wire_7368;
    wire new_Jinkela_wire_2448;
    wire new_Jinkela_wire_5318;
    wire new_Jinkela_wire_3964;
    wire new_Jinkela_wire_7233;
    wire new_Jinkela_wire_7343;
    wire new_Jinkela_wire_2799;
    wire new_Jinkela_wire_3170;
    wire new_Jinkela_wire_4354;
    wire _0503_;
    wire new_Jinkela_wire_7731;
    wire new_Jinkela_wire_7598;
    wire new_Jinkela_wire_4994;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_6314;
    wire new_Jinkela_wire_6820;
    wire new_Jinkela_wire_7826;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_5098;
    wire new_Jinkela_wire_3687;
    wire new_Jinkela_wire_4653;
    wire new_Jinkela_wire_4914;
    wire _0719_;
    wire new_Jinkela_wire_5715;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_4209;
    wire new_Jinkela_wire_7156;
    wire new_Jinkela_wire_4394;
    wire new_Jinkela_wire_5002;
    wire _1103_;
    wire _0306_;
    wire new_Jinkela_wire_4017;
    wire new_Jinkela_wire_4179;
    wire new_Jinkela_wire_7537;
    wire new_Jinkela_wire_6733;
    wire new_Jinkela_wire_4264;
    wire new_Jinkela_wire_5913;
    wire new_Jinkela_wire_7542;
    wire new_Jinkela_wire_5630;
    wire new_Jinkela_wire_7075;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_6600;
    wire new_Jinkela_wire_2113;
    wire new_Jinkela_wire_5589;
    wire new_Jinkela_wire_5291;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_7439;
    wire new_Jinkela_wire_3033;
    wire _0243_;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_7329;
    wire new_Jinkela_wire_5204;
    wire new_Jinkela_wire_2962;
    wire new_Jinkela_wire_7031;
    wire _0137_;
    wire new_Jinkela_wire_5010;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_7061;
    wire new_Jinkela_wire_7247;
    wire _0528_;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_6452;
    wire new_Jinkela_wire_6248;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_5534;
    wire new_Jinkela_wire_6392;
    wire new_Jinkela_wire_2592;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_6739;
    wire new_Jinkela_wire_4148;
    wire new_Jinkela_wire_4724;
    wire _0838_;
    wire new_Jinkela_wire_2616;
    wire new_Jinkela_wire_1948;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_7647;
    wire new_Jinkela_wire_7682;
    wire _0253_;
    wire _0446_;
    wire new_Jinkela_wire_3252;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_2620;
    wire new_Jinkela_wire_2009;
    wire _0499_;
    wire new_Jinkela_wire_3989;
    wire new_Jinkela_wire_5238;
    wire new_Jinkela_wire_4820;
    wire new_Jinkela_wire_6238;
    wire new_Jinkela_wire_7519;
    wire new_Jinkela_wire_5345;
    wire new_Jinkela_wire_5549;
    wire new_Jinkela_wire_7916;
    wire new_Jinkela_wire_4776;
    wire new_Jinkela_wire_6431;
    wire new_Jinkela_wire_2928;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_2955;
    wire new_Jinkela_wire_7966;
    wire new_Jinkela_wire_6088;
    wire new_Jinkela_wire_2994;
    wire new_Jinkela_wire_8018;
    wire _0458_;
    wire new_Jinkela_wire_7653;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_6788;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_7820;
    wire new_Jinkela_wire_3637;
    wire _0063_;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_3711;
    wire new_Jinkela_wire_1844;
    wire new_Jinkela_wire_5001;
    wire new_Jinkela_wire_4560;
    wire new_Jinkela_wire_1906;
    wire _0276_;
    wire new_Jinkela_wire_1939;
    wire new_Jinkela_wire_5647;
    wire new_Jinkela_wire_2710;
    wire new_Jinkela_wire_6453;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_3221;
    wire new_Jinkela_wire_5812;
    wire new_Jinkela_wire_2385;
    wire new_Jinkela_wire_7964;
    wire new_Jinkela_wire_4722;
    wire new_Jinkela_wire_5127;
    wire new_Jinkela_wire_7767;
    wire new_Jinkela_wire_7666;
    wire new_Jinkela_wire_2582;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_2849;
    wire new_Jinkela_wire_3449;
    wire new_Jinkela_wire_6867;
    wire new_Jinkela_wire_4457;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_5103;
    wire new_Jinkela_wire_4080;
    wire new_Jinkela_wire_3468;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_5280;
    wire _1005_;
    wire _0874_;
    wire new_Jinkela_wire_7416;
    wire _0920_;
    wire new_Jinkela_wire_5447;
    wire new_Jinkela_wire_2605;
    wire new_net_2419;
    wire new_Jinkela_wire_4767;
    wire new_Jinkela_wire_5383;
    wire new_Jinkela_wire_6672;
    wire new_Jinkela_wire_7599;
    wire _0972_;
    wire new_Jinkela_wire_3642;
    wire _0416_;
    wire new_Jinkela_wire_7430;
    wire new_Jinkela_wire_2138;
    wire new_Jinkela_wire_7817;
    wire new_Jinkela_wire_5717;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_782;
    wire _0197_;
    wire new_Jinkela_wire_2297;
    wire new_Jinkela_wire_6478;
    wire new_Jinkela_wire_7108;
    wire new_Jinkela_wire_5175;
    wire new_Jinkela_wire_7623;
    wire new_Jinkela_wire_5026;
    wire _1201_;
    wire new_net_2407;
    wire new_Jinkela_wire_6834;
    wire new_Jinkela_wire_5785;
    wire _0298_;
    wire new_Jinkela_wire_794;
    wire _1216_;
    wire new_Jinkela_wire_7507;
    wire new_Jinkela_wire_6523;
    wire new_Jinkela_wire_7540;
    wire new_Jinkela_wire_5412;
    wire new_Jinkela_wire_6402;
    wire new_Jinkela_wire_2304;
    wire new_Jinkela_wire_1943;
    wire new_Jinkela_wire_1067;
    wire _0616_;
    wire _1130_;
    wire new_Jinkela_wire_4713;
    wire new_Jinkela_wire_4445;
    wire new_Jinkela_wire_5124;
    wire _0453_;
    wire _0789_;
    wire _0520_;
    wire new_Jinkela_wire_5905;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_3090;
    wire new_net_2465;
    wire new_Jinkela_wire_7193;
    wire new_Jinkela_wire_5639;
    wire _0255_;
    wire new_Jinkela_wire_6304;
    wire new_Jinkela_wire_7678;
    wire new_net_2463;
    wire new_Jinkela_wire_3179;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_2224;
    wire new_Jinkela_wire_6843;
    wire new_Jinkela_wire_3909;
    wire new_Jinkela_wire_2299;
    wire new_Jinkela_wire_5174;
    wire new_Jinkela_wire_80;
    wire _0038_;
    wire _0733_;
    wire new_Jinkela_wire_5677;
    wire _1014_;
    wire new_Jinkela_wire_4798;
    wire _0530_;
    wire new_Jinkela_wire_6076;
    wire new_Jinkela_wire_7904;
    wire new_Jinkela_wire_6060;
    wire new_Jinkela_wire_1549;
    wire new_Jinkela_wire_6528;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_5014;
    wire new_Jinkela_wire_6714;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_4061;
    wire new_Jinkela_wire_7552;
    wire new_Jinkela_wire_2711;
    wire new_Jinkela_wire_6691;
    wire new_Jinkela_wire_7102;
    wire new_Jinkela_wire_4692;
    wire new_Jinkela_wire_4875;
    wire _0827_;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_4912;
    wire _1021_;
    wire new_Jinkela_wire_5661;
    wire new_Jinkela_wire_2746;
    wire new_Jinkela_wire_3376;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_2151;
    wire new_Jinkela_wire_6519;
    wire new_Jinkela_wire_4536;
    wire _0580_;
    wire new_Jinkela_wire_7356;
    wire _0227_;
    wire new_Jinkela_wire_5696;
    wire new_Jinkela_wire_2331;
    wire new_Jinkela_wire_3012;
    wire new_Jinkela_wire_7880;
    wire new_Jinkela_wire_2422;
    wire new_Jinkela_wire_5773;
    wire new_Jinkela_wire_5684;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_4348;
    wire new_Jinkela_wire_5330;
    wire _0642_;
    wire new_Jinkela_wire_2720;
    wire new_Jinkela_wire_6701;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_5327;
    wire new_Jinkela_wire_7679;
    wire new_Jinkela_wire_4603;
    wire new_net_16;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_4961;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_6586;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_4551;
    wire _1131_;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_6950;
    wire new_Jinkela_wire_7625;
    wire new_Jinkela_wire_5651;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_7728;
    wire new_Jinkela_wire_7488;
    wire _0662_;
    wire new_Jinkela_wire_3839;
    wire new_Jinkela_wire_3060;
    wire new_Jinkela_wire_6710;
    wire new_Jinkela_wire_4895;
    wire new_Jinkela_wire_2378;
    wire new_Jinkela_wire_76;
    wire _0379_;
    wire new_Jinkela_wire_4703;
    wire _0584_;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_7716;
    wire new_Jinkela_wire_7251;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_2570;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_3704;
    wire _0738_;
    wire new_Jinkela_wire_4582;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_7318;
    wire new_Jinkela_wire_6759;
    wire new_Jinkela_wire_7017;
    wire new_Jinkela_wire_7870;
    wire new_Jinkela_wire_3649;
    wire new_Jinkela_wire_2487;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_6875;
    wire new_Jinkela_wire_4647;
    wire new_Jinkela_wire_154;
    wire _0937_;
    wire new_Jinkela_wire_5050;
    wire new_Jinkela_wire_3925;
    wire new_Jinkela_wire_3082;
    wire new_Jinkela_wire_4918;
    wire new_Jinkela_wire_5844;
    wire new_Jinkela_wire_281;
    wire _0060_;
    wire new_Jinkela_wire_7182;
    wire new_Jinkela_wire_2769;
    wire new_Jinkela_wire_1884;
    wire new_Jinkela_wire_3601;
    wire new_Jinkela_wire_6053;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_4814;
    wire new_Jinkela_wire_6110;
    wire new_Jinkela_wire_4239;
    wire new_Jinkela_wire_7676;
    wire new_Jinkela_wire_5837;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_6138;
    wire new_Jinkela_wire_1987;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_2159;
    wire new_Jinkela_wire_4717;
    wire new_Jinkela_wire_2229;
    wire new_Jinkela_wire_3816;
    wire new_Jinkela_wire_7215;
    wire _0478_;
    wire new_Jinkela_wire_7014;
    wire new_Jinkela_wire_7434;
    wire _1049_;
    wire new_Jinkela_wire_4960;
    wire new_Jinkela_wire_1754;
    wire new_Jinkela_wire_4253;
    wire new_Jinkela_wire_4256;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_3067;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_5308;
    wire new_Jinkela_wire_5625;
    wire new_Jinkela_wire_6677;
    wire new_Jinkela_wire_1979;
    wire new_Jinkela_wire_7274;
    wire new_Jinkela_wire_5513;
    wire new_Jinkela_wire_3775;
    wire new_Jinkela_wire_2932;
    wire new_Jinkela_wire_7652;
    wire _0383_;
    wire new_Jinkela_wire_3748;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_2687;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_3215;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_2925;
    wire new_Jinkela_wire_8006;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_6106;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_6296;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_3580;
    wire new_Jinkela_wire_1931;
    wire new_Jinkela_wire_2278;
    wire new_Jinkela_wire_4231;
    wire new_Jinkela_wire_3759;
    wire new_Jinkela_wire_6956;
    wire new_Jinkela_wire_3324;
    wire new_Jinkela_wire_4280;
    wire new_Jinkela_wire_4625;
    wire _0368_;
    wire new_Jinkela_wire_2280;
    wire new_Jinkela_wire_2813;
    wire new_Jinkela_wire_7735;
    wire new_Jinkela_wire_7159;
    wire new_Jinkela_wire_2511;
    wire new_Jinkela_wire_1043;
    wire _0256_;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_5845;
    wire new_Jinkela_wire_3632;
    wire new_Jinkela_wire_7581;
    wire new_Jinkela_wire_3911;
    wire _1197_;
    wire new_Jinkela_wire_7438;
    wire new_Jinkela_wire_7104;
    wire new_Jinkela_wire_6127;
    wire new_Jinkela_wire_4678;
    wire _0777_;
    wire new_Jinkela_wire_4368;
    wire _0166_;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_6360;
    wire new_Jinkela_wire_6988;
    wire new_Jinkela_wire_2895;
    wire new_Jinkela_wire_2744;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_3938;
    wire new_Jinkela_wire_6489;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_3788;
    wire new_Jinkela_wire_3993;
    wire new_Jinkela_wire_5693;
    wire new_Jinkela_wire_6848;
    wire _0844_;
    wire new_Jinkela_wire_5258;
    wire new_Jinkela_wire_3407;
    wire new_Jinkela_wire_3461;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_7457;
    wire _0321_;
    wire new_Jinkela_wire_4730;
    wire new_Jinkela_wire_6169;
    wire _0550_;
    wire new_Jinkela_wire_43;
    wire _0711_;
    wire _0543_;
    wire new_Jinkela_wire_3143;
    wire new_Jinkela_wire_6811;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_2148;
    wire new_Jinkela_wire_461;
    wire _0609_;
    wire new_Jinkela_wire_5861;
    wire new_Jinkela_wire_3274;
    wire new_Jinkela_wire_7732;
    wire new_Jinkela_wire_6502;
    wire new_Jinkela_wire_5708;
    wire new_Jinkela_wire_3761;
    wire new_Jinkela_wire_2364;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_3218;
    wire new_Jinkela_wire_568;
    wire _0995_;
    wire new_Jinkela_wire_6743;
    wire new_Jinkela_wire_7646;
    wire new_Jinkela_wire_7310;
    wire new_net_2453;
    wire new_Jinkela_wire_6460;
    wire new_Jinkela_wire_5875;
    wire new_Jinkela_wire_5085;
    wire new_Jinkela_wire_4449;
    wire new_Jinkela_wire_7409;
    wire new_Jinkela_wire_7501;
    wire new_Jinkela_wire_6488;
    wire _0035_;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_4885;
    wire new_Jinkela_wire_3954;
    wire new_Jinkela_wire_3744;
    wire new_Jinkela_wire_5091;
    wire _0988_;
    wire new_Jinkela_wire_3077;
    wire new_Jinkela_wire_5700;
    wire new_Jinkela_wire_2796;
    wire new_Jinkela_wire_4555;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_4072;
    wire new_Jinkela_wire_5914;
    wire new_Jinkela_wire_6483;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_1994;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_3666;
    wire new_Jinkela_wire_4845;
    wire new_Jinkela_wire_5737;
    wire new_Jinkela_wire_5512;
    wire new_Jinkela_wire_5961;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_7286;
    wire new_Jinkela_wire_4504;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_4736;
    wire new_Jinkela_wire_7813;
    wire new_Jinkela_wire_3006;
    wire new_Jinkela_wire_5819;
    wire new_Jinkela_wire_4880;
    wire new_Jinkela_wire_2886;
    wire new_Jinkela_wire_2619;
    wire new_Jinkela_wire_1659;
    wire _1189_;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_3610;
    wire new_Jinkela_wire_6545;
    wire _0053_;
    wire new_Jinkela_wire_1871;
    wire new_Jinkela_wire_7892;
    wire _0953_;
    wire new_Jinkela_wire_6510;
    wire new_Jinkela_wire_5824;
    wire new_Jinkela_wire_5024;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_7068;
    wire new_Jinkela_wire_5099;
    wire new_Jinkela_wire_4807;
    wire new_Jinkela_wire_3290;
    wire _0836_;
    wire new_Jinkela_wire_2281;
    wire new_Jinkela_wire_7268;
    wire new_Jinkela_wire_1949;
    wire new_Jinkela_wire_4136;
    wire new_Jinkela_wire_7448;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_4299;
    wire new_Jinkela_wire_3564;
    wire new_Jinkela_wire_3243;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_3638;
    wire new_Jinkela_wire_4973;
    wire new_Jinkela_wire_3206;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_5196;
    wire new_Jinkela_wire_4492;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_7272;
    wire new_Jinkela_wire_7441;
    wire new_Jinkela_wire_4120;
    wire new_Jinkela_wire_4878;
    wire new_Jinkela_wire_6986;
    wire new_Jinkela_wire_6648;
    wire new_Jinkela_wire_1862;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_4704;
    wire new_Jinkela_wire_6056;
    wire new_Jinkela_wire_6096;
    wire new_Jinkela_wire_6894;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_6794;
    wire _0637_;
    wire _0426_;
    wire new_Jinkela_wire_6560;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_3121;
    wire new_Jinkela_wire_5681;
    wire new_Jinkela_wire_2750;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_4106;
    wire new_Jinkela_wire_7695;
    wire new_Jinkela_wire_5294;
    wire new_Jinkela_wire_1985;
    wire new_Jinkela_wire_2066;
    wire _0365_;
    wire new_Jinkela_wire_6317;
    wire new_Jinkela_wire_1457;
    wire _0898_;
    wire new_Jinkela_wire_5910;
    wire new_Jinkela_wire_1750;
    wire new_Jinkela_wire_7035;
    wire new_Jinkela_wire_3998;
    wire new_Jinkela_wire_1649;
    wire _0036_;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_1815;
    wire _0628_;
    wire new_Jinkela_wire_7153;
    wire new_Jinkela_wire_3467;
    wire new_Jinkela_wire_2635;
    wire new_Jinkela_wire_4089;
    wire new_Jinkela_wire_5095;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_2323;
    wire new_Jinkela_wire_3408;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_7491;
    wire _1061_;
    wire new_Jinkela_wire_7543;
    wire new_Jinkela_wire_70;
    wire _1184_;
    wire new_Jinkela_wire_1503;
    wire new_Jinkela_wire_1857;
    wire new_Jinkela_wire_3723;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_5143;
    wire new_Jinkela_wire_4571;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_4268;
    wire new_Jinkela_wire_7484;
    wire _0199_;
    wire new_Jinkela_wire_1773;
    wire new_Jinkela_wire_6055;
    wire new_Jinkela_wire_3912;
    wire new_Jinkela_wire_5063;
    wire _0002_;
    wire new_Jinkela_wire_6445;
    wire _0203_;
    wire new_Jinkela_wire_7309;
    wire new_Jinkela_wire_5603;
    wire _1098_;
    wire new_Jinkela_wire_2812;
    wire new_net_2349;
    wire new_Jinkela_wire_5851;
    wire new_Jinkela_wire_4512;
    wire new_Jinkela_wire_2968;
    wire new_Jinkela_wire_1082;
    wire _1120_;
    wire _1031_;
    wire new_Jinkela_wire_6881;
    wire new_Jinkela_wire_5109;
    wire new_Jinkela_wire_3373;
    wire new_Jinkela_wire_3698;
    wire new_Jinkela_wire_3019;
    wire new_Jinkela_wire_4650;
    wire _0905_;
    wire new_Jinkela_wire_7829;
    wire new_Jinkela_wire_5660;
    wire _0325_;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_4938;
    wire _1194_;
    wire new_Jinkela_wire_5104;
    wire new_Jinkela_wire_6817;
    wire new_Jinkela_wire_3047;
    wire new_Jinkela_wire_3624;
    wire new_Jinkela_wire_3573;
    wire new_Jinkela_wire_4871;
    wire new_Jinkela_wire_3289;
    wire new_Jinkela_wire_3639;
    wire new_Jinkela_wire_2548;
    wire new_Jinkela_wire_7650;
    wire new_Jinkela_wire_6791;
    wire new_Jinkela_wire_7088;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_2249;
    wire new_Jinkela_wire_6394;
    wire _0526_;
    wire new_Jinkela_wire_1036;
    wire new_Jinkela_wire_7119;
    wire new_Jinkela_wire_3056;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_4576;
    wire new_Jinkela_wire_2667;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_7011;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_4483;
    wire new_Jinkela_wire_5874;
    wire new_Jinkela_wire_4113;
    wire new_Jinkela_wire_4527;
    wire new_Jinkela_wire_2178;
    wire new_Jinkela_wire_4216;
    wire new_Jinkela_wire_5479;
    wire new_Jinkela_wire_6658;
    wire new_Jinkela_wire_1561;
    wire _0548_;
    wire new_Jinkela_wire_1751;
    wire new_Jinkela_wire_3236;
    wire new_net_2379;
    wire new_Jinkela_wire_6666;
    wire new_Jinkela_wire_7833;
    wire new_Jinkela_wire_4012;
    wire new_Jinkela_wire_4732;
    wire _1150_;
    wire new_Jinkela_wire_5304;
    wire new_Jinkela_wire_6107;
    wire new_Jinkela_wire_2235;
    wire _0745_;
    wire new_Jinkela_wire_6253;
    wire new_Jinkela_wire_6158;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_5758;
    wire new_Jinkela_wire_931;
    wire _0803_;
    wire _1148_;
    wire new_net_2487;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_3633;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_5714;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_4414;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_2356;
    wire _0561_;
    wire _0757_;
    wire new_Jinkela_wire_7584;
    wire new_Jinkela_wire_6384;
    wire new_Jinkela_wire_6994;
    wire new_Jinkela_wire_6958;
    wire new_Jinkela_wire_3230;
    wire _0563_;
    wire new_Jinkela_wire_5234;
    wire new_Jinkela_wire_5456;
    wire new_Jinkela_wire_4932;
    wire new_Jinkela_wire_7125;
    wire new_Jinkela_wire_7196;
    wire new_Jinkela_wire_6590;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_2216;
    wire new_Jinkela_wire_5268;
    wire new_Jinkela_wire_7926;
    wire new_Jinkela_wire_4111;
    wire new_Jinkela_wire_3319;
    wire new_Jinkela_wire_8002;
    wire new_Jinkela_wire_2223;
    wire _0116_;
    wire new_Jinkela_wire_2139;
    wire new_Jinkela_wire_6451;
    wire new_Jinkela_wire_4212;
    wire new_Jinkela_wire_7600;
    wire _1011_;
    wire new_Jinkela_wire_7918;
    wire new_Jinkela_wire_2051;
    wire new_Jinkela_wire_7346;
    wire new_Jinkela_wire_5522;
    wire new_Jinkela_wire_3343;
    wire _1133_;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_6720;
    wire _1220_;
    wire new_Jinkela_wire_3674;
    wire new_Jinkela_wire_5803;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_4257;
    wire new_Jinkela_wire_4851;
    wire new_Jinkela_wire_4247;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_3172;
    wire new_Jinkela_wire_6140;
    wire new_Jinkela_wire_6352;
    wire new_Jinkela_wire_2417;
    wire new_Jinkela_wire_7962;
    wire new_Jinkela_wire_5117;
    wire _0936_;
    wire new_Jinkela_wire_7527;
    wire new_Jinkela_wire_6182;
    wire new_Jinkela_wire_2543;
    wire new_Jinkela_wire_7734;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_7295;
    wire new_Jinkela_wire_7465;
    wire _0417_;
    wire new_Jinkela_wire_3463;
    wire new_Jinkela_wire_3820;
    wire new_Jinkela_wire_7579;
    wire new_Jinkela_wire_7618;
    wire new_Jinkela_wire_3708;
    wire new_Jinkela_wire_5194;
    wire new_Jinkela_wire_4330;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_3803;
    wire _1083_;
    wire new_Jinkela_wire_2889;
    wire new_Jinkela_wire_3278;
    wire new_Jinkela_wire_7946;
    wire new_Jinkela_wire_7015;
    wire new_Jinkela_wire_4177;
    wire new_Jinkela_wire_1966;
    wire new_Jinkela_wire_5753;
    wire new_Jinkela_wire_5491;
    wire new_Jinkela_wire_3157;
    wire new_Jinkela_wire_2381;
    wire _0947_;
    wire new_Jinkela_wire_6872;
    wire new_Jinkela_wire_648;
    wire _0293_;
    wire new_Jinkela_wire_7874;
    wire new_Jinkela_wire_2193;
    wire new_Jinkela_wire_2885;
    wire new_Jinkela_wire_5033;
    wire new_Jinkela_wire_2153;
    wire _1198_;
    wire new_Jinkela_wire_7327;
    wire new_Jinkela_wire_2860;
    wire new_Jinkela_wire_4221;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_6821;
    wire new_Jinkela_wire_5520;
    wire new_Jinkela_wire_2782;
    wire _0251_;
    wire new_Jinkela_wire_3798;
    wire new_Jinkela_wire_5405;
    wire new_Jinkela_wire_5831;
    wire new_Jinkela_wire_5638;
    wire new_Jinkela_wire_4444;
    wire new_Jinkela_wire_3622;
    wire new_Jinkela_wire_5275;
    wire _1116_;
    wire new_Jinkela_wire_4426;
    wire new_Jinkela_wire_5218;
    wire new_Jinkela_wire_7336;
    wire new_Jinkela_wire_3224;
    wire new_Jinkela_wire_7505;
    wire new_Jinkela_wire_3763;
    wire _1238_;
    wire new_Jinkela_wire_1971;
    wire new_Jinkela_wire_3378;
    wire new_Jinkela_wire_5938;
    wire new_Jinkela_wire_5794;
    wire _0581_;
    wire new_Jinkela_wire_4860;
    wire new_Jinkela_wire_5039;
    wire _0376_;
    wire new_Jinkela_wire_2748;
    wire new_Jinkela_wire_6729;
    wire new_Jinkela_wire_481;
    wire _0455_;
    wire new_Jinkela_wire_5458;
    wire new_Jinkela_wire_7895;
    wire new_Jinkela_wire_3259;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_3526;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_4934;
    wire new_Jinkela_wire_6702;
    wire new_Jinkela_wire_4601;
    wire new_Jinkela_wire_3581;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_6882;
    wire new_Jinkela_wire_6241;
    wire new_Jinkela_wire_3920;
    wire new_Jinkela_wire_4594;
    wire new_Jinkela_wire_4005;
    wire new_Jinkela_wire_6675;
    wire new_Jinkela_wire_3962;
    wire new_Jinkela_wire_3095;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_6073;
    wire new_Jinkela_wire_7239;
    wire new_Jinkela_wire_7054;
    wire new_Jinkela_wire_5576;
    wire new_Jinkela_wire_5399;
    wire new_Jinkela_wire_4749;
    wire new_Jinkela_wire_3254;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_3729;
    wire new_Jinkela_wire_7630;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_6641;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_3548;
    wire new_Jinkela_wire_3054;
    wire new_Jinkela_wire_2641;
    wire new_Jinkela_wire_4547;
    wire new_Jinkela_wire_4956;
    wire _0363_;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_5776;
    wire new_Jinkela_wire_5941;
    wire _0763_;
    wire new_Jinkela_wire_7948;
    wire _0867_;
    wire new_Jinkela_wire_3668;
    wire new_Jinkela_wire_7969;
    wire new_Jinkela_wire_3945;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_2597;
    wire new_Jinkela_wire_2785;
    wire new_Jinkela_wire_6644;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_2800;
    wire new_Jinkela_wire_3472;
    wire new_Jinkela_wire_3080;
    wire new_Jinkela_wire_2774;
    wire new_Jinkela_wire_5952;
    wire new_Jinkela_wire_2680;
    wire new_Jinkela_wire_1832;
    wire new_Jinkela_wire_1481;
    wire _0132_;
    wire new_Jinkela_wire_5608;
    wire new_Jinkela_wire_6799;
    wire _1028_;
    wire new_Jinkela_wire_2416;
    wire new_Jinkela_wire_5159;
    wire new_Jinkela_wire_4957;
    wire _0791_;
    wire new_Jinkela_wire_5471;
    wire new_Jinkela_wire_3068;
    wire _0759_;
    wire _1068_;
    wire new_Jinkela_wire_1753;
    wire new_net_2431;
    wire new_Jinkela_wire_4626;
    wire _0817_;
    wire new_Jinkela_wire_4538;
    wire new_Jinkela_wire_5413;
    wire new_Jinkela_wire_4500;
    wire new_Jinkela_wire_193;
    wire _1026_;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_6418;
    wire new_Jinkela_wire_5767;
    wire new_Jinkela_wire_7269;
    wire _1193_;
    wire _0766_;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_5375;
    wire new_Jinkela_wire_3370;
    wire new_Jinkela_wire_2479;
    wire new_Jinkela_wire_7571;
    wire new_Jinkela_wire_2513;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_5205;
    wire new_Jinkela_wire_6007;
    wire new_Jinkela_wire_7908;
    wire new_Jinkela_wire_7832;
    wire new_Jinkela_wire_5624;
    wire new_Jinkela_wire_5937;
    wire new_Jinkela_wire_6943;
    wire new_Jinkela_wire_7968;
    wire _0598_;
    wire _0436_;
    wire _1072_;
    wire new_Jinkela_wire_4175;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_2591;
    wire new_Jinkela_wire_4181;
    wire new_Jinkela_wire_4731;
    wire new_Jinkela_wire_3749;
    wire new_Jinkela_wire_5825;
    wire new_Jinkela_wire_3605;
    wire new_Jinkela_wire_4183;
    wire new_Jinkela_wire_4768;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_2679;
    wire _1239_;
    wire new_Jinkela_wire_6783;
    wire _0095_;
    wire new_Jinkela_wire_542;
    wire _0760_;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_6592;
    wire new_Jinkela_wire_5016;
    wire new_Jinkela_wire_3159;
    wire new_Jinkela_wire_3429;
    wire _0993_;
    wire new_Jinkela_wire_6195;
    wire _0384_;
    wire new_net_2353;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_3509;
    wire new_Jinkela_wire_6310;
    wire new_Jinkela_wire_4321;
    wire new_Jinkela_wire_1989;
    wire new_Jinkela_wire_5920;
    wire new_Jinkela_wire_4350;
    wire _1200_;
    wire new_Jinkela_wire_4149;
    wire new_Jinkela_wire_5678;
    wire new_net_3;
    wire new_Jinkela_wire_7667;
    wire new_Jinkela_wire_3534;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_3535;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_3389;
    wire new_Jinkela_wire_4525;
    wire new_Jinkela_wire_6461;
    wire new_Jinkela_wire_5168;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_1697;
    wire new_Jinkela_wire_5669;
    wire new_Jinkela_wire_4125;
    wire new_Jinkela_wire_3673;
    wire new_Jinkela_wire_5597;
    wire new_Jinkela_wire_3559;
    wire new_Jinkela_wire_7658;
    wire new_Jinkela_wire_4290;
    wire new_Jinkela_wire_5667;
    wire new_Jinkela_wire_6373;
    wire new_Jinkela_wire_3222;
    wire new_Jinkela_wire_480;
    wire new_Jinkela_wire_2395;
    wire new_Jinkela_wire_3374;
    wire new_Jinkela_wire_5685;
    wire _1020_;
    wire new_Jinkela_wire_6035;
    wire new_net_2489;
    wire _1213_;
    wire new_Jinkela_wire_7073;
    wire new_Jinkela_wire_4336;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_3955;
    wire new_Jinkela_wire_6275;
    wire new_Jinkela_wire_3145;
    wire new_Jinkela_wire_2930;
    wire _0466_;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_5277;
    wire new_Jinkela_wire_5210;
    wire new_Jinkela_wire_7802;
    wire new_Jinkela_wire_4378;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_3594;
    wire new_Jinkela_wire_1583;
    wire _0876_;
    wire new_Jinkela_wire_979;
    wire _0331_;
    wire new_Jinkela_wire_3968;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_5229;
    wire new_Jinkela_wire_6636;
    wire new_Jinkela_wire_1538;
    wire _1138_;
    wire _0289_;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_4249;
    wire _0345_;
    wire new_Jinkela_wire_4592;
    wire new_Jinkela_wire_6540;
    wire new_Jinkela_wire_5224;
    wire new_Jinkela_wire_6588;
    wire new_Jinkela_wire_7464;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_7004;
    wire new_Jinkela_wire_4669;
    wire _0829_;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_2627;
    wire new_net_2507;
    wire new_Jinkela_wire_4981;
    wire new_Jinkela_wire_4828;
    wire new_Jinkela_wire_5890;
    wire new_Jinkela_wire_2484;
    wire new_Jinkela_wire_6447;
    wire new_Jinkela_wire_2649;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_5254;
    wire new_Jinkela_wire_4162;
    wire new_Jinkela_wire_5183;
    wire _0824_;
    wire _0567_;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_2232;
    wire new_Jinkela_wire_5028;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_6656;
    wire new_Jinkela_wire_2586;
    wire _0873_;
    wire new_Jinkela_wire_3907;
    wire new_Jinkela_wire_7480;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_765;
    wire _1039_;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_5829;
    wire new_Jinkela_wire_7112;
    wire new_Jinkela_wire_6741;
    wire _0558_;
    wire new_Jinkela_wire_3997;
    wire new_Jinkela_wire_5295;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_6189;
    wire new_Jinkela_wire_4642;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_4437;
    wire new_Jinkela_wire_6599;
    wire new_Jinkela_wire_3867;
    wire new_Jinkela_wire_3844;
    wire new_Jinkela_wire_3118;
    wire _0774_;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_6051;
    wire _0103_;
    wire new_Jinkela_wire_2989;
    wire new_Jinkela_wire_3786;
    wire _1025_;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_6777;
    wire _0123_;
    wire new_Jinkela_wire_6642;
    wire new_Jinkela_wire_3811;
    wire new_Jinkela_wire_1077;
    wire _1044_;
    wire new_Jinkela_wire_6432;
    wire _0611_;
    wire _1126_;
    wire new_Jinkela_wire_1628;
    wire _0500_;
    wire new_Jinkela_wire_7305;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_4160;
    wire new_Jinkela_wire_4146;
    wire _1166_;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_3828;
    wire new_Jinkela_wire_5832;
    wire new_Jinkela_wire_5893;
    wire new_Jinkela_wire_3458;
    wire _0081_;
    wire new_Jinkela_wire_3645;
    wire _0775_;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_4946;
    wire _0667_;
    wire _1226_;
    wire _0915_;
    wire new_Jinkela_wire_5426;
    wire new_Jinkela_wire_2475;
    wire new_Jinkela_wire_7249;
    wire _0250_;
    wire new_Jinkela_wire_2634;
    wire new_Jinkela_wire_3102;
    wire new_Jinkela_wire_7643;
    wire new_Jinkela_wire_6400;
    wire new_Jinkela_wire_1745;
    wire _0019_;
    wire new_Jinkela_wire_3108;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_4821;
    wire new_Jinkela_wire_7388;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_3515;
    wire new_Jinkela_wire_3417;
    wire new_Jinkela_wire_7528;
    wire new_Jinkela_wire_4453;
    wire _0207_;
    wire _0224_;
    wire new_Jinkela_wire_3758;
    wire new_Jinkela_wire_6175;
    wire new_Jinkela_wire_6492;
    wire new_net_2473;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_3799;
    wire new_Jinkela_wire_4151;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_7328;
    wire _0822_;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_6052;
    wire new_Jinkela_wire_6335;
    wire _0252_;
    wire new_Jinkela_wire_6273;
    wire new_Jinkela_wire_3574;
    wire new_Jinkela_wire_2951;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_7384;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_1617;
    wire new_Jinkela_wire_5640;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_2336;
    wire new_Jinkela_wire_3017;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_2399;
    wire new_Jinkela_wire_4430;
    wire new_Jinkela_wire_3064;
    wire _0507_;
    wire new_Jinkela_wire_2754;
    wire new_Jinkela_wire_7271;
    wire new_Jinkela_wire_5801;
    wire new_Jinkela_wire_6753;
    wire _0769_;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_1935;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_3894;
    wire new_Jinkela_wire_5653;
    wire new_Jinkela_wire_5698;
    wire new_Jinkela_wire_5775;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_6567;
    wire _1088_;
    wire new_Jinkela_wire_3824;
    wire new_Jinkela_wire_3177;
    wire new_Jinkela_wire_3641;
    wire new_Jinkela_wire_7536;
    wire _0958_;
    wire new_Jinkela_wire_7901;
    wire new_Jinkela_wire_5478;
    wire new_Jinkela_wire_2209;
    wire new_Jinkela_wire_3193;
    wire new_Jinkela_wire_1184;
    wire _1001_;
    wire new_Jinkela_wire_3113;
    wire _1242_;
    wire new_Jinkela_wire_3323;
    wire new_Jinkela_wire_3135;
    wire new_Jinkela_wire_6115;
    wire new_Jinkela_wire_3797;
    wire new_Jinkela_wire_5620;
    wire new_Jinkela_wire_1776;
    wire new_Jinkela_wire_4353;
    wire new_Jinkela_wire_3059;
    wire new_Jinkela_wire_6836;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_2661;
    wire _0351_;
    wire new_Jinkela_wire_5673;
    wire new_Jinkela_wire_3664;
    wire new_Jinkela_wire_7304;
    wire new_Jinkela_wire_5362;
    wire new_Jinkela_wire_7415;
    wire new_Jinkela_wire_7037;
    wire new_Jinkela_wire_6579;
    wire new_Jinkela_wire_2424;
    wire _0462_;
    wire new_Jinkela_wire_6050;
    wire _1089_;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_4636;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_6157;
    wire new_Jinkela_wire_7844;
    wire _0726_;
    wire new_Jinkela_wire_6049;
    wire new_Jinkela_wire_5526;
    wire new_Jinkela_wire_3959;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_4611;
    wire new_Jinkela_wire_7726;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_7270;
    wire new_Jinkela_wire_4054;
    wire _1096_;
    wire _0943_;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_3144;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_4990;
    wire new_Jinkela_wire_4174;
    wire new_Jinkela_wire_5652;
    wire new_Jinkela_wire_1723;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_5432;
    wire new_Jinkela_wire_6511;
    wire new_Jinkela_wire_5559;
    wire new_Jinkela_wire_65;
    wire _0287_;
    wire new_Jinkela_wire_7093;
    wire new_Jinkela_wire_4701;
    wire _1167_;
    wire _1100_;
    wire new_Jinkela_wire_5402;
    wire new_Jinkela_wire_1934;
    wire new_Jinkela_wire_2438;
    wire new_Jinkela_wire_2598;
    wire new_Jinkela_wire_5899;
    wire new_Jinkela_wire_3271;
    wire _0393_;
    wire new_Jinkela_wire_1224;
    wire new_Jinkela_wire_4786;
    wire new_Jinkela_wire_6605;
    wire new_Jinkela_wire_6935;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_7541;
    wire new_Jinkela_wire_6755;
    wire new_Jinkela_wire_2286;
    wire new_Jinkela_wire_6458;
    wire new_Jinkela_wire_2508;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_7722;
    wire new_Jinkela_wire_4337;
    wire new_Jinkela_wire_2881;
    wire new_Jinkela_wire_6306;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_7975;
    wire new_Jinkela_wire_7720;
    wire new_Jinkela_wire_3151;
    wire _0231_;
    wire new_Jinkela_wire_7835;
    wire new_Jinkela_wire_5492;
    wire new_Jinkela_wire_5221;
    wire new_Jinkela_wire_2847;
    wire _0806_;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_4230;
    wire new_Jinkela_wire_3614;
    wire new_Jinkela_wire_6883;
    wire new_Jinkela_wire_4936;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_1767;
    wire new_Jinkela_wire_7042;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_6773;
    wire new_Jinkela_wire_5090;
    wire new_Jinkela_wire_2415;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_3571;
    wire new_Jinkela_wire_3733;
    wire new_Jinkela_wire_4165;
    wire _1023_;
    wire new_Jinkela_wire_5269;
    wire new_Jinkela_wire_3937;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_5628;
    wire new_Jinkela_wire_2311;
    wire new_Jinkela_wire_2804;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_4380;
    wire new_Jinkela_wire_2911;
    wire new_Jinkela_wire_7282;
    wire new_Jinkela_wire_5604;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_4826;
    wire new_Jinkela_wire_5613;
    wire new_Jinkela_wire_2623;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_7702;
    wire new_Jinkela_wire_6809;
    wire new_Jinkela_wire_4447;
    wire new_Jinkela_wire_6374;
    wire new_Jinkela_wire_6152;
    wire _0440_;
    wire new_Jinkela_wire_2176;
    wire new_Jinkela_wire_4248;
    wire new_Jinkela_wire_3250;
    wire new_Jinkela_wire_4270;
    wire new_Jinkela_wire_3004;
    wire _0663_;
    wire new_Jinkela_wire_2099;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_7205;
    wire _1188_;
    wire new_Jinkela_wire_6724;
    wire new_Jinkela_wire_3181;
    wire new_Jinkela_wire_5148;
    wire _0020_;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_6888;
    wire new_Jinkela_wire_7224;
    wire new_Jinkela_wire_5131;
    wire new_Jinkela_wire_4235;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_6369;
    wire new_Jinkela_wire_4222;
    wire new_Jinkela_wire_4076;
    wire new_Jinkela_wire_3014;
    wire new_Jinkela_wire_4652;
    wire new_Jinkela_wire_7401;
    wire new_Jinkela_wire_6575;
    wire new_Jinkela_wire_3015;
    wire new_Jinkela_wire_3189;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_7779;
    wire new_Jinkela_wire_2963;
    wire _0194_;
    wire new_Jinkela_wire_1234;
    wire _0014_;
    wire new_Jinkela_wire_2590;
    wire new_Jinkela_wire_5705;
    wire new_Jinkela_wire_880;
    wire _0587_;
    wire _1135_;
    wire new_Jinkela_wire_6087;
    wire new_Jinkela_wire_3587;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_6839;
    wire new_Jinkela_wire_4157;
    wire new_Jinkela_wire_7189;
    wire new_Jinkela_wire_6662;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_3861;
    wire new_Jinkela_wire_6619;
    wire new_Jinkela_wire_304;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_2485;
    wire new_Jinkela_wire_2347;
    wire _0597_;
    wire _0218_;
    wire new_Jinkela_wire_4123;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_6853;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_4193;
    wire new_Jinkela_wire_5044;
    wire _0894_;
    wire new_Jinkela_wire_2270;
    wire new_Jinkela_wire_3020;
    wire new_Jinkela_wire_3899;
    wire new_Jinkela_wire_2197;
    wire new_Jinkela_wire_6505;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_7030;
    wire new_Jinkela_wire_7648;
    wire new_Jinkela_wire_3195;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_7452;
    wire new_Jinkela_wire_4720;
    wire new_Jinkela_wire_6842;
    wire new_Jinkela_wire_7923;
    wire new_Jinkela_wire_6946;
    wire new_Jinkela_wire_6046;
    wire new_Jinkela_wire_6798;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_4468;
    wire new_Jinkela_wire_1013;
    wire _0328_;
    wire _0736_;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_4969;
    wire new_Jinkela_wire_7531;
    wire new_Jinkela_wire_7206;
    wire new_Jinkela_wire_2043;
    wire new_Jinkela_wire_5967;
    wire new_Jinkela_wire_6838;
    wire new_Jinkela_wire_5689;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_2681;
    wire new_Jinkela_wire_3418;
    wire new_Jinkela_wire_3940;
    wire new_Jinkela_wire_3538;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_3066;
    wire new_Jinkela_wire_3626;
    wire new_Jinkela_wire_7563;
    wire new_net_17;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_3849;
    wire new_Jinkela_wire_5442;
    wire new_Jinkela_wire_3331;
    wire new_Jinkela_wire_6565;
    wire new_Jinkela_wire_5866;
    wire new_Jinkela_wire_3737;
    wire new_Jinkela_wire_6391;
    wire new_Jinkela_wire_3905;
    wire new_Jinkela_wire_1819;
    wire new_Jinkela_wire_5225;
    wire _1081_;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_6468;
    wire new_Jinkela_wire_1485;
    wire new_Jinkela_wire_7858;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_5115;
    wire new_Jinkela_wire_5642;
    wire new_Jinkela_wire_7756;
    wire new_Jinkela_wire_6229;
    wire new_Jinkela_wire_1455;
    wire _1074_;
    wire new_Jinkela_wire_3361;
    wire new_Jinkela_wire_2526;
    wire new_Jinkela_wire_4496;
    wire new_Jinkela_wire_6301;
    wire new_Jinkela_wire_7051;
    wire new_Jinkela_wire_7321;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_7243;
    wire new_Jinkela_wire_6254;
    wire _0312_;
    wire new_Jinkela_wire_4968;
    wire new_Jinkela_wire_1237;
    wire _0405_;
    wire new_Jinkela_wire_6617;
    wire new_Jinkela_wire_5547;
    wire _0230_;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_2455;
    wire new_Jinkela_wire_4513;
    wire _0560_;
    wire new_Jinkela_wire_6048;
    wire new_Jinkela_wire_4827;
    wire new_Jinkela_wire_4793;
    wire new_Jinkela_wire_7943;
    wire new_Jinkela_wire_4526;
    wire _0361_;
    wire new_Jinkela_wire_1921;
    wire new_Jinkela_wire_4327;
    wire _0724_;
    wire new_Jinkela_wire_4227;
    wire new_Jinkela_wire_6215;
    wire new_Jinkela_wire_7811;
    wire new_Jinkela_wire_4108;
    wire new_Jinkela_wire_2588;
    wire _0716_;
    wire new_Jinkela_wire_7521;
    wire new_Jinkela_wire_7115;
    wire new_Jinkela_wire_23;
    wire new_Jinkela_wire_6846;
    wire new_Jinkela_wire_3552;
    wire new_Jinkela_wire_7723;
    wire new_Jinkela_wire_1323;
    wire _0729_;
    wire new_Jinkela_wire_7529;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_4223;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_4779;
    wire _1158_;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_883;
    wire _0310_;
    wire _0781_;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_5631;
    wire new_Jinkela_wire_4395;
    wire new_net_2383;
    wire new_Jinkela_wire_2648;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_6409;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_5697;
    wire new_Jinkela_wire_4777;
    wire new_Jinkela_wire_2815;
    wire new_Jinkela_wire_2340;
    wire new_Jinkela_wire_7191;
    wire new_Jinkela_wire_7759;
    wire new_Jinkela_wire_5496;
    wire new_Jinkela_wire_7822;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_7098;
    wire new_Jinkela_wire_7428;
    wire new_Jinkela_wire_7963;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_4619;
    wire new_Jinkela_wire_2977;
    wire new_Jinkela_wire_3554;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_3562;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_7934;
    wire new_Jinkela_wire_3362;
    wire new_Jinkela_wire_3238;
    wire _0623_;
    wire new_Jinkela_wire_307;
    wire _0189_;
    wire _1035_;
    wire new_Jinkela_wire_6066;
    wire _0016_;
    wire new_Jinkela_wire_2617;
    wire new_Jinkela_wire_2742;
    wire new_Jinkela_wire_5594;
    wire new_Jinkela_wire_5011;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_8009;
    wire new_Jinkela_wire_993;
    wire new_net_2443;
    wire new_Jinkela_wire_4224;
    wire new_Jinkela_wire_7790;
    wire new_Jinkela_wire_4479;
    wire new_Jinkela_wire_4940;
    wire new_Jinkela_wire_5862;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_2998;
    wire _1057_;
    wire new_Jinkela_wire_7244;
    wire new_Jinkela_wire_6760;
    wire new_Jinkela_wire_4317;
    wire new_Jinkela_wire_6584;
    wire _0408_;
    wire _0261_;
    wire new_Jinkela_wire_5255;
    wire new_Jinkela_wire_4450;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_4775;
    wire _1051_;
    wire new_Jinkela_wire_2501;
    wire new_Jinkela_wire_4978;
    wire new_Jinkela_wire_5152;
    wire new_Jinkela_wire_5641;
    wire _0544_;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_3499;
    wire new_Jinkela_wire_2894;
    wire new_Jinkela_wire_5351;
    wire new_Jinkela_wire_5515;
    wire new_Jinkela_wire_1202;
    wire new_Jinkela_wire_2394;
    wire _1235_;
    wire _0650_;
    wire new_Jinkela_wire_6474;
    wire new_Jinkela_wire_3328;
    wire new_Jinkela_wire_6497;
    wire new_Jinkela_wire_3540;
    wire new_Jinkela_wire_2866;
    wire new_Jinkela_wire_6606;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_2803;
    wire new_Jinkela_wire_3207;
    wire new_Jinkela_wire_2303;
    wire _0160_;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_7597;
    wire new_Jinkela_wire_5894;
    wire new_Jinkela_wire_6776;
    wire new_Jinkela_wire_4800;
    wire new_Jinkela_wire_4196;
    wire new_Jinkela_wire_4996;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_7183;
    wire new_Jinkela_wire_7610;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_6655;
    wire new_Jinkela_wire_6645;
    wire new_Jinkela_wire_1439;
    wire new_Jinkela_wire_7717;
    wire _0945_;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_7715;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_5892;
    wire new_Jinkela_wire_3721;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_4315;
    wire new_Jinkela_wire_2554;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_5256;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_4274;
    wire _1186_;
    wire _0087_;
    wire _0430_;
    wire new_Jinkela_wire_4579;
    wire new_Jinkela_wire_2248;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_3809;
    wire _0832_;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_5828;
    wire new_Jinkela_wire_2121;
    wire new_Jinkela_wire_6556;
    wire new_Jinkela_wire_5997;
    wire new_Jinkela_wire_2741;
    wire new_Jinkela_wire_3465;
    wire _0201_;
    wire new_Jinkela_wire_2192;
    wire new_Jinkela_wire_3522;
    wire new_Jinkela_wire_6640;
    wire new_Jinkela_wire_1422;
    wire _0151_;
    wire new_Jinkela_wire_4403;
    wire new_Jinkela_wire_1403;
    wire new_Jinkela_wire_6851;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_7569;
    wire new_Jinkela_wire_2269;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_3593;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_2478;
    wire _0949_;
    wire new_Jinkela_wire_6927;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_1437;
    wire _0773_;
    wire new_Jinkela_wire_7983;
    wire new_Jinkela_wire_6646;
    wire new_Jinkela_wire_7172;
    wire new_Jinkela_wire_2291;
    wire new_Jinkela_wire_4105;
    wire _0178_;
    wire new_Jinkela_wire_4184;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_5879;
    wire _0163_;
    wire new_Jinkela_wire_3261;
    wire new_Jinkela_wire_7644;
    wire _0911_;
    wire new_Jinkela_wire_798;
    wire _0987_;
    wire new_Jinkela_wire_5092;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_4393;
    wire new_Jinkela_wire_4635;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_4170;
    wire new_Jinkela_wire_4695;
    wire _1060_;
    wire new_Jinkela_wire_2116;
    wire new_Jinkela_wire_2601;
    wire new_Jinkela_wire_5584;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_1139;
    wire _0661_;
    wire new_Jinkela_wire_3483;
    wire new_Jinkela_wire_4379;
    wire new_Jinkela_wire_2829;
    wire new_Jinkela_wire_3819;
    wire new_Jinkela_wire_5029;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_4756;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_2329;
    wire new_Jinkela_wire_3908;
    wire new_Jinkela_wire_3284;
    wire new_Jinkela_wire_2839;
    wire new_Jinkela_wire_5873;
    wire new_Jinkela_wire_5904;
    wire new_Jinkela_wire_2371;
    wire new_Jinkela_wire_6380;
    wire new_Jinkela_wire_5276;
    wire new_Jinkela_wire_1883;
    wire new_Jinkela_wire_4198;
    wire new_Jinkela_wire_2112;
    wire _1217_;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_6135;
    wire new_Jinkela_wire_6698;
    wire new_Jinkela_wire_4971;
    wire new_Jinkela_wire_1093;
    wire new_Jinkela_wire_7689;
    wire _0985_;
    wire new_Jinkela_wire_885;
    wire new_net_2403;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_7114;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_7202;
    wire _0957_;
    wire _0414_;
    wire new_Jinkela_wire_6841;
    wire new_Jinkela_wire_2683;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_5712;
    wire new_Jinkela_wire_3866;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_5305;
    wire new_Jinkela_wire_6576;
    wire new_Jinkela_wire_6218;
    wire new_Jinkela_wire_3858;
    wire new_Jinkela_wire_5477;
    wire new_Jinkela_wire_5876;
    wire new_Jinkela_wire_5887;
    wire _1127_;
    wire _1000_;
    wire _1030_;
    wire new_Jinkela_wire_3903;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_5971;
    wire _0279_;
    wire new_Jinkela_wire_7737;
    wire new_Jinkela_wire_2164;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_4924;
    wire new_Jinkela_wire_5570;
    wire new_Jinkela_wire_6070;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_3311;
    wire new_Jinkela_wire_2204;
    wire new_Jinkela_wire_6708;
    wire new_Jinkela_wire_3754;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_7669;
    wire new_Jinkela_wire_4933;
    wire new_Jinkela_wire_3707;
    wire new_Jinkela_wire_5816;
    wire new_Jinkela_wire_6025;
    wire new_Jinkela_wire_6034;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_4167;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_1743;
    wire new_Jinkela_wire_4244;
    wire new_Jinkela_wire_3291;
    wire new_Jinkela_wire_2902;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_3875;
    wire new_Jinkela_wire_6351;
    wire new_Jinkela_wire_5965;
    wire new_Jinkela_wire_6339;
    wire _0983_;
    wire new_Jinkela_wire_5583;
    wire _0146_;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_377;
    wire new_Jinkela_wire_3692;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_3257;
    wire new_Jinkela_wire_3625;
    wire new_Jinkela_wire_4665;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_5315;
    wire new_Jinkela_wire_3322;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_6111;
    wire new_Jinkela_wire_6746;
    wire new_Jinkela_wire_3310;
    wire new_Jinkela_wire_5400;
    wire new_Jinkela_wire_6198;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_4271;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_3340;
    wire new_Jinkela_wire_7664;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_5490;
    wire new_Jinkela_wire_6583;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_2880;
    wire new_Jinkela_wire_3514;
    wire new_Jinkela_wire_4002;
    wire new_Jinkela_wire_926;
    wire _0464_;
    wire new_Jinkela_wire_6235;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_7069;
    wire new_Jinkela_wire_2134;
    wire _0657_;
    wire _0319_;
    wire new_Jinkela_wire_4431;
    wire new_Jinkela_wire_6563;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_7360;
    wire new_Jinkela_wire_4419;
    wire _0494_;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_5966;
    wire new_Jinkela_wire_3354;
    wire new_Jinkela_wire_4541;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_1955;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_6309;
    wire new_Jinkela_wire_5744;
    wire new_Jinkela_wire_2988;
    wire new_Jinkela_wire_4958;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_2531;
    wire _0571_;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_3387;
    wire new_net_2481;
    wire new_Jinkela_wire_5948;
    wire new_Jinkela_wire_2002;
    wire new_Jinkela_wire_5133;
    wire new_Jinkela_wire_2646;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_3675;
    wire new_Jinkela_wire_2387;
    wire new_Jinkela_wire_7503;
    wire new_Jinkela_wire_3979;
    wire new_Jinkela_wire_6637;
    wire new_Jinkela_wire_2996;
    wire new_Jinkela_wire_3420;
    wire new_Jinkela_wire_2362;
    wire new_Jinkela_wire_7000;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_265;
    wire _0211_;
    wire new_Jinkela_wire_7067;
    wire new_Jinkela_wire_4187;
    wire new_Jinkela_wire_3356;
    wire new_Jinkela_wire_6197;
    wire new_Jinkela_wire_2368;
    wire new_net_2375;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_2671;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_2187;
    wire new_Jinkela_wire_5747;
    wire new_Jinkela_wire_614;
    wire _0814_;
    wire new_Jinkela_wire_5474;
    wire new_Jinkela_wire_6830;
    wire _0907_;
    wire _0354_;
    wire new_Jinkela_wire_7052;
    wire _0390_;
    wire new_Jinkela_wire_2662;
    wire new_Jinkela_wire_6913;
    wire new_Jinkela_wire_2672;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_5446;
    wire new_Jinkela_wire_3961;
    wire new_Jinkela_wire_7961;
    wire new_Jinkela_wire_3836;
    wire new_Jinkela_wire_6874;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_5782;
    wire new_Jinkela_wire_7974;
    wire new_Jinkela_wire_7838;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_2184;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_4951;
    wire new_Jinkela_wire_2790;
    wire _0542_;
    wire new_Jinkela_wire_7186;
    wire _0797_;
    wire new_Jinkela_wire_3349;
    wire new_Jinkela_wire_1436;
    wire _0699_;
    wire new_Jinkela_wire_6738;
    wire new_Jinkela_wire_6187;
    wire _0262_;
    wire new_Jinkela_wire_1646;
    wire _0161_;
    wire new_Jinkela_wire_2809;
    wire new_net_2459;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_7266;
    wire new_Jinkela_wire_6148;
    wire new_Jinkela_wire_2529;
    wire _0226_;
    wire _1078_;
    wire new_Jinkela_wire_4835;
    wire new_Jinkela_wire_4191;
    wire new_Jinkela_wire_6164;
    wire new_Jinkela_wire_2851;
    wire new_Jinkela_wire_6651;
    wire new_Jinkela_wire_4415;
    wire new_Jinkela_wire_3158;
    wire new_Jinkela_wire_7936;
    wire new_Jinkela_wire_6938;
    wire new_Jinkela_wire_2692;
    wire new_Jinkela_wire_3933;
    wire new_Jinkela_wire_4850;
    wire new_Jinkela_wire_4389;
    wire new_Jinkela_wire_7418;
    wire new_Jinkela_wire_2277;
    wire _1173_;
    wire new_Jinkela_wire_2766;
    wire new_Jinkela_wire_3358;
    wire new_Jinkela_wire_6028;
    wire new_Jinkela_wire_2941;
    wire new_Jinkela_wire_4456;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_6626;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_3873;
    wire new_Jinkela_wire_7929;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_6870;
    wire new_Jinkela_wire_2333;
    wire new_Jinkela_wire_4953;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_4085;
    wire _0105_;
    wire new_Jinkela_wire_2882;
    wire new_Jinkela_wire_652;
    wire _0702_;
    wire new_Jinkela_wire_6501;
    wire new_Jinkela_wire_4725;
    wire new_Jinkela_wire_7660;
    wire _0209_;
    wire new_Jinkela_wire_1705;
    wire new_Jinkela_wire_3480;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_7364;
    wire _1245_;
    wire new_Jinkela_wire_1470;
    wire new_net_8;
    wire new_Jinkela_wire_6245;
    wire new_Jinkela_wire_1938;
    wire _0802_;
    wire new_Jinkela_wire_5554;
    wire new_Jinkela_wire_6744;
    wire new_Jinkela_wire_5510;
    wire new_Jinkela_wire_5519;
    wire new_Jinkela_wire_3739;
    wire new_Jinkela_wire_3269;
    wire new_Jinkela_wire_2471;
    wire _0347_;
    wire new_Jinkela_wire_5723;
    wire new_Jinkela_wire_5403;
    wire new_Jinkela_wire_3939;
    wire new_Jinkela_wire_4269;
    wire new_Jinkela_wire_4281;
    wire new_Jinkela_wire_4301;
    wire _0939_;
    wire new_Jinkela_wire_1777;
    wire _1113_;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_4771;
    wire new_Jinkela_wire_3150;
    wire new_Jinkela_wire_3958;
    wire _1077_;
    wire new_Jinkela_wire_7888;
    wire new_Jinkela_wire_7616;
    wire new_Jinkela_wire_4400;
    wire new_Jinkela_wire_6855;
    wire new_Jinkela_wire_5670;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_5591;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_7366;
    wire new_net_2395;
    wire _0259_;
    wire new_Jinkela_wire_4091;
    wire new_Jinkela_wire_7372;
    wire new_Jinkela_wire_6008;
    wire new_Jinkela_wire_7558;
    wire new_Jinkela_wire_3442;
    wire _0174_;
    wire new_Jinkela_wire_3314;
    wire new_Jinkela_wire_3069;
    wire new_Jinkela_wire_6342;
    wire new_Jinkela_wire_7137;
    wire new_Jinkela_wire_1728;
    wire new_Jinkela_wire_4233;
    wire new_Jinkela_wire_7704;
    wire new_Jinkela_wire_3722;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_3476;
    wire new_Jinkela_wire_3532;
    wire new_Jinkela_wire_6832;
    wire new_Jinkela_wire_4823;
    wire new_Jinkela_wire_1954;
    wire new_Jinkela_wire_2106;
    wire new_Jinkela_wire_7499;
    wire new_Jinkela_wire_2263;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_7789;
    wire new_Jinkela_wire_906;
    wire _0236_;
    wire new_Jinkela_wire_5357;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_6367;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_4370;
    wire new_Jinkela_wire_4049;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_5518;
    wire _0525_;
    wire new_Jinkela_wire_3504;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_5995;
    wire new_Jinkela_wire_6580;
    wire new_Jinkela_wire_3599;
    wire new_Jinkela_wire_3084;
    wire new_Jinkela_wire_2556;
    wire new_Jinkela_wire_6193;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_5310;
    wire new_Jinkela_wire_2826;
    wire new_Jinkela_wire_6967;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_6987;
    wire _0110_;
    wire new_Jinkela_wire_452;
    wire new_net_15;
    wire new_Jinkela_wire_59;
    wire _0554_;
    wire new_Jinkela_wire_4867;
    wire new_Jinkela_wire_5214;
    wire new_Jinkela_wire_7615;
    wire _1161_;
    wire new_Jinkela_wire_6288;
    wire new_Jinkela_wire_3864;
    wire new_Jinkela_wire_7478;
    wire _1137_;
    wire new_Jinkela_wire_3270;
    wire new_Jinkela_wire_7446;
    wire new_Jinkela_wire_6613;
    wire new_Jinkela_wire_3092;
    wire new_Jinkela_wire_7221;
    wire new_Jinkela_wire_5121;
    wire new_Jinkela_wire_4446;
    wire _0149_;
    wire new_Jinkela_wire_4639;
    wire new_Jinkela_wire_1950;
    wire _0772_;
    wire new_Jinkela_wire_4099;
    wire new_Jinkela_wire_7217;
    wire new_Jinkela_wire_992;
    wire _0270_;
    wire new_Jinkela_wire_5377;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_5672;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_3714;
    wire new_Jinkela_wire_4454;
    wire new_Jinkela_wire_1089;
    wire new_Jinkela_wire_2844;
    wire new_Jinkela_wire_4307;
    wire new_Jinkela_wire_5909;
    wire new_Jinkela_wire_2515;
    wire new_Jinkela_wire_4602;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_5654;
    wire new_Jinkela_wire_5930;
    wire new_Jinkela_wire_2768;
    wire new_Jinkela_wire_5248;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_7232;
    wire new_Jinkela_wire_3385;
    wire new_Jinkela_wire_3892;
    wire _1008_;
    wire new_Jinkela_wire_3724;
    wire new_Jinkela_wire_4294;
    wire new_Jinkela_wire_2264;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_238;
    wire _0029_;
    wire _0686_;
    wire new_Jinkela_wire_6682;
    wire _0688_;
    wire new_Jinkela_wire_2414;
    wire new_net_2501;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_2576;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_4200;
    wire new_Jinkela_wire_7471;
    wire new_Jinkela_wire_6632;
    wire new_Jinkela_wire_6348;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_5886;
    wire new_Jinkela_wire_3464;
    wire _0557_;
    wire _0659_;
    wire new_Jinkela_wire_5582;
    wire new_Jinkela_wire_7560;
    wire new_Jinkela_wire_6277;
    wire _1191_;
    wire new_Jinkela_wire_5083;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_4746;
    wire new_Jinkela_wire_7296;
    wire _0787_;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_3833;
    wire new_Jinkela_wire_2573;
    wire new_Jinkela_wire_4025;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_6176;
    wire new_Jinkela_wire_3076;
    wire new_Jinkela_wire_4058;
    wire new_Jinkela_wire_4925;
    wire new_Jinkela_wire_4014;
    wire _0717_;
    wire new_Jinkela_wire_3489;
    wire new_Jinkela_wire_3335;
    wire new_Jinkela_wire_4423;
    wire new_Jinkela_wire_4645;
    wire new_Jinkela_wire_7577;
    wire new_Jinkela_wire_4266;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_4874;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_5316;
    wire new_Jinkela_wire_5381;
    wire new_Jinkela_wire_6354;
    wire new_Jinkela_wire_4719;
    wire new_Jinkela_wire_4710;
    wire new_Jinkela_wire_6340;
    wire new_Jinkela_wire_6042;
    wire new_Jinkela_wire_7570;
    wire new_Jinkela_wire_6845;
    wire new_Jinkela_wire_5111;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_5716;
    wire new_Jinkela_wire_4137;
    wire new_Jinkela_wire_2676;
    wire new_Jinkela_wire_7812;
    wire _0260_;
    wire new_Jinkela_wire_2686;
    wire new_Jinkela_wire_7941;
    wire new_Jinkela_wire_6623;
    wire new_Jinkela_wire_3350;
    wire new_Jinkela_wire_2654;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_7213;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_2391;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_3555;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_7473;
    wire new_Jinkela_wire_4288;
    wire new_Jinkela_wire_2076;
    wire new_Jinkela_wire_4052;
    wire new_Jinkela_wire_6426;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_6219;
    wire new_Jinkela_wire_7279;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_6090;
    wire new_Jinkela_wire_5889;
    wire new_Jinkela_wire_2201;
    wire new_Jinkela_wire_5682;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_7198;
    wire _0402_;
    wire new_Jinkela_wire_2690;
    wire _0372_;
    wire new_Jinkela_wire_7712;
    wire new_Jinkela_wire_6969;
    wire new_Jinkela_wire_3112;
    wire new_Jinkela_wire_2251;
    wire new_Jinkela_wire_6043;
    wire new_Jinkela_wire_3302;
    wire new_Jinkela_wire_6818;
    wire new_Jinkela_wire_6065;
    wire new_Jinkela_wire_6188;
    wire new_Jinkela_wire_7231;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_5430;
    wire new_Jinkela_wire_1408;
    wire _0410_;
    wire new_Jinkela_wire_2143;
    wire new_Jinkela_wire_4846;
    wire _1054_;
    wire new_net_2457;
    wire _0165_;
    wire new_Jinkela_wire_5138;
    wire new_Jinkela_wire_2194;
    wire new_Jinkela_wire_2656;
    wire new_Jinkela_wire_7898;
    wire _0888_;
    wire new_Jinkela_wire_763;
    wire _0755_;
    wire new_Jinkela_wire_2186;
    wire new_Jinkela_wire_6062;
    wire _0705_;
    wire new_Jinkela_wire_4631;
    wire new_Jinkela_wire_4947;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_3199;
    wire new_Jinkela_wire_7972;
    wire new_Jinkela_wire_5691;
    wire new_Jinkela_wire_3486;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_5444;
    wire new_Jinkela_wire_5354;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_2995;
    wire new_net_2475;
    wire new_Jinkela_wire_1526;
    wire new_net_2503;
    wire new_Jinkela_wire_7586;
    wire _1176_;
    wire new_Jinkela_wire_6762;
    wire new_Jinkela_wire_6585;
    wire new_Jinkela_wire_5774;
    wire new_Jinkela_wire_8001;
    wire _0150_;
    wire new_Jinkela_wire_6503;
    wire new_Jinkela_wire_6263;
    wire new_Jinkela_wire_5151;
    wire new_Jinkela_wire_4675;
    wire new_Jinkela_wire_6265;
    wire new_Jinkela_wire_6852;
    wire new_Jinkela_wire_6891;
    wire new_Jinkela_wire_6079;
    wire _0979_;
    wire new_Jinkela_wire_7564;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_2789;
    wire new_Jinkela_wire_5037;
    wire new_Jinkela_wire_6032;
    wire new_Jinkela_wire_5052;
    wire new_Jinkela_wire_4841;
    wire new_Jinkela_wire_6508;
    wire new_Jinkela_wire_3046;
    wire new_Jinkela_wire_5739;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_5166;
    wire _1222_;
    wire new_Jinkela_wire_7578;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_7341;
    wire new_Jinkela_wire_4853;
    wire new_Jinkela_wire_2095;
    wire new_Jinkela_wire_3146;
    wire new_Jinkela_wire_7203;
    wire new_Jinkela_wire_7062;
    wire new_Jinkela_wire_7163;
    wire new_Jinkela_wire_1514;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_5551;
    wire new_Jinkela_wire_4075;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_5469;
    wire new_Jinkela_wire_7385;
    wire new_Jinkela_wire_4917;
    wire new_Jinkela_wire_1801;
    wire new_Jinkela_wire_7332;
    wire new_Jinkela_wire_6531;
    wire new_Jinkela_wire_4794;
    wire new_net_2433;
    wire new_Jinkela_wire_4194;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_5390;
    wire new_Jinkela_wire_1627;
    wire new_Jinkela_wire_7825;
    wire new_Jinkela_wire_2170;
    wire new_Jinkela_wire_1847;
    wire _0088_;
    wire new_Jinkela_wire_7886;
    wire new_Jinkela_wire_5649;
    wire new_Jinkela_wire_6532;
    wire new_Jinkela_wire_2893;
    wire new_Jinkela_wire_2992;
    wire new_Jinkela_wire_6649;
    wire new_Jinkela_wire_3869;
    wire new_Jinkela_wire_4110;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_6466;
    wire new_Jinkela_wire_1833;
    wire new_Jinkela_wire_3437;
    wire new_Jinkela_wire_6191;
    wire new_Jinkela_wire_4098;
    wire new_Jinkela_wire_7977;
    wire _0559_;
    wire new_Jinkela_wire_6459;
    wire new_Jinkela_wire_4945;
    wire new_Jinkela_wire_6370;
    wire new_Jinkela_wire_5082;
    wire new_Jinkela_wire_7056;
    wire new_Jinkela_wire_6243;
    wire new_Jinkela_wire_7690;
    wire new_net_2377;
    wire new_Jinkela_wire_1804;
    wire new_Jinkela_wire_2657;
    wire new_Jinkela_wire_7122;
    wire new_Jinkela_wire_4050;
    wire new_Jinkela_wire_4112;
    wire new_Jinkela_wire_7375;
    wire new_Jinkela_wire_4641;
    wire new_Jinkela_wire_7741;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_6906;
    wire new_Jinkela_wire_6963;
    wire new_Jinkela_wire_3175;
    wire new_Jinkela_wire_6167;
    wire new_Jinkela_wire_5605;
    wire _1165_;
    wire new_Jinkela_wire_1866;
    wire new_Jinkela_wire_1727;
    wire new_Jinkela_wire_2160;
    wire new_Jinkela_wire_2579;
    wire new_Jinkela_wire_5976;
    wire _0737_;
    wire new_Jinkela_wire_2792;
    wire new_Jinkela_wire_5676;
    wire new_Jinkela_wire_6699;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_7081;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_1960;
    wire _0136_;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_3325;
    wire new_Jinkela_wire_5612;
    wire new_Jinkela_wire_5273;
    wire new_Jinkela_wire_5702;
    wire new_Jinkela_wire_7128;
    wire new_Jinkela_wire_5118;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_6481;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_2342;
    wire new_Jinkela_wire_2199;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_4515;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_3345;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_3210;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_1055;
    wire _0195_;
    wire new_Jinkela_wire_5251;
    wire new_Jinkela_wire_1757;
    wire new_Jinkela_wire_3444;
    wire new_net_2417;
    wire new_Jinkela_wire_5903;
    wire new_Jinkela_wire_4362;
    wire new_net_2437;
    wire new_Jinkela_wire_6005;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_3031;
    wire _0184_;
    wire new_Jinkela_wire_3817;
    wire _0885_;
    wire new_Jinkela_wire_3078;
    wire new_Jinkela_wire_4040;
    wire new_Jinkela_wire_2512;
    wire _0878_;
    wire new_Jinkela_wire_4388;
    wire _0693_;
    wire new_Jinkela_wire_5417;
    wire new_Jinkela_wire_3178;
    wire new_Jinkela_wire_3694;
    wire new_Jinkela_wire_7768;
    wire _1236_;
    wire new_Jinkela_wire_3148;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_2055;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_3371;
    wire new_Jinkela_wire_7397;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_7169;
    wire new_Jinkela_wire_5300;
    wire _0229_;
    wire new_Jinkela_wire_3657;
    wire _0799_;
    wire _0620_;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_5500;
    wire new_Jinkela_wire_3002;
    wire _1058_;
    wire new_Jinkela_wire_2971;
    wire _0845_;
    wire new_Jinkela_wire_7241;
    wire new_Jinkela_wire_6419;
    wire new_Jinkela_wire_2763;
    wire new_Jinkela_wire_2697;
    wire new_Jinkela_wire_5298;
    wire new_Jinkela_wire_7670;
    wire _0684_;
    wire new_Jinkela_wire_2535;
    wire new_Jinkela_wire_1779;
    wire new_Jinkela_wire_5611;
    wire new_Jinkela_wire_6252;
    wire new_Jinkela_wire_6470;
    wire new_Jinkela_wire_4983;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_4032;
    wire new_Jinkela_wire_2017;
    wire new_Jinkela_wire_3300;
    wire new_Jinkela_wire_2718;
    wire new_Jinkela_wire_3808;
    wire new_Jinkela_wire_3226;
    wire new_Jinkela_wire_6715;
    wire new_Jinkela_wire_7245;
    wire new_Jinkela_wire_6098;
    wire new_Jinkela_wire_968;
    wire _0487_;
    wire new_Jinkela_wire_5267;
    wire new_Jinkela_wire_5324;
    wire new_Jinkela_wire_4795;
    wire new_Jinkela_wire_4442;
    wire new_Jinkela_wire_5588;
    wire new_Jinkela_wire_7410;
    wire new_Jinkela_wire_2421;
    wire _0108_;
    wire new_Jinkela_wire_1661;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_4575;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_2685;
    wire new_Jinkela_wire_1942;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_4338;
    wire _0457_;
    wire _0039_;
    wire _0658_;
    wire new_Jinkela_wire_3209;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_2149;
    wire new_Jinkela_wire_4928;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_7639;
    wire new_Jinkela_wire_5242;
    wire new_Jinkela_wire_1655;
    wire new_Jinkela_wire_4142;
    wire new_Jinkela_wire_4782;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_2131;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_2125;
    wire new_Jinkela_wire_7875;
    wire new_Jinkela_wire_6929;
    wire new_Jinkela_wire_4530;
    wire new_Jinkela_wire_7141;
    wire new_Jinkela_wire_7135;
    wire new_Jinkela_wire_5374;
    wire new_Jinkela_wire_1156;
    wire _0037_;
    wire new_Jinkela_wire_7655;
    wire new_net_4;
    wire new_Jinkela_wire_2980;
    wire new_Jinkela_wire_5293;
    wire new_Jinkela_wire_6029;
    wire new_Jinkela_wire_4188;
    wire new_Jinkela_wire_2583;
    wire new_Jinkela_wire_7905;
    wire new_Jinkela_wire_1326;
    wire _0480_;
    wire new_Jinkela_wire_4364;
    wire _0994_;
    wire new_Jinkela_wire_5908;
    wire new_Jinkela_wire_6931;
    wire new_net_2413;
    wire new_Jinkela_wire_7701;
    wire new_Jinkela_wire_2290;
    wire _0752_;
    wire new_Jinkela_wire_4207;
    wire _0989_;
    wire new_Jinkela_wire_6180;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_7250;
    wire new_Jinkela_wire_5671;
    wire new_Jinkela_wire_2631;
    wire new_Jinkela_wire_7315;
    wire new_Jinkela_wire_3762;
    wire new_Jinkela_wire_7884;
    wire new_Jinkela_wire_7025;
    wire new_Jinkela_wire_7551;
    wire _0634_;
    wire _0465_;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_7476;
    wire new_Jinkela_wire_6303;
    wire new_Jinkela_wire_3975;
    wire new_Jinkela_wire_7788;
    wire _0698_;
    wire new_Jinkela_wire_3730;
    wire new_Jinkela_wire_3517;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_451;
    wire _0493_;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_4797;
    wire new_Jinkela_wire_5944;
    wire _0387_;
    wire new_Jinkela_wire_2990;
    wire new_Jinkela_wire_6312;
    wire new_Jinkela_wire_6547;
    wire new_Jinkela_wire_6414;
    wire new_Jinkela_wire_6749;
    wire new_Jinkela_wire_6727;
    wire new_Jinkela_wire_2510;
    wire new_Jinkela_wire_5675;
    wire _0459_;
    wire _1210_;
    wire new_Jinkela_wire_2220;
    wire new_Jinkela_wire_5322;
    wire new_Jinkela_wire_2817;
    wire _0676_;
    wire new_Jinkela_wire_4324;
    wire new_Jinkela_wire_3292;
    wire new_Jinkela_wire_3443;
    wire new_Jinkela_wire_67;
    wire _1175_;
    wire new_Jinkela_wire_6161;
    wire new_Jinkela_wire_1882;
    wire new_Jinkela_wire_4844;
    wire new_Jinkela_wire_6336;
    wire new_Jinkela_wire_1822;
    wire new_Jinkela_wire_5355;
    wire new_Jinkela_wire_2823;
    wire new_Jinkela_wire_7021;
    wire new_Jinkela_wire_3129;
    wire new_Jinkela_wire_3285;
    wire new_Jinkela_wire_6315;
    wire _0631_;
    wire new_Jinkela_wire_4883;
    wire _0516_;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_6258;
    wire new_Jinkela_wire_2123;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_3527;
    wire new_net_2427;
    wire new_Jinkela_wire_3608;
    wire new_Jinkela_wire_3163;
    wire new_Jinkela_wire_3629;
    wire new_Jinkela_wire_3883;
    wire _1006_;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_4030;
    wire new_Jinkela_wire_2226;
    wire new_Jinkela_wire_3212;
    wire new_Jinkela_wire_2490;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_7489;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_5053;
    wire _1162_;
    wire _0856_;
    wire _0780_;
    wire new_Jinkela_wire_7591;
    wire new_Jinkela_wire_5884;
    wire new_Jinkela_wire_2035;
    wire new_Jinkela_wire_6676;
    wire new_Jinkela_wire_2316;
    wire new_Jinkela_wire_5826;
    wire new_Jinkela_wire_908;
    wire _0140_;
    wire new_Jinkela_wire_5687;
    wire new_Jinkela_wire_6233;
    wire new_Jinkela_wire_6695;
    wire new_Jinkela_wire_7158;
    wire new_Jinkela_wire_1530;
    wire new_Jinkela_wire_6133;
    wire new_Jinkela_wire_6975;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_6349;
    wire new_Jinkela_wire_6186;
    wire new_Jinkela_wire_6101;
    wire new_Jinkela_wire_3375;
    wire new_Jinkela_wire_7848;
    wire new_Jinkela_wire_5694;
    wire new_Jinkela_wire_4094;
    wire new_Jinkela_wire_4053;
    wire new_Jinkela_wire_4325;
    wire new_Jinkela_wire_2016;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_4607;
    wire new_Jinkela_wire_2388;
    wire new_Jinkela_wire_7175;
    wire new_Jinkela_wire_3297;
    wire new_Jinkela_wire_2539;
    wire _0749_;
    wire new_Jinkela_wire_2869;
    wire new_Jinkela_wire_2884;
    wire new_Jinkela_wire_7437;
    wire new_Jinkela_wire_7700;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_3228;
    wire new_Jinkela_wire_6122;
    wire new_Jinkela_wire_5516;
    wire new_Jinkela_wire_7371;
    wire new_Jinkela_wire_1843;
    wire _0128_;
    wire new_Jinkela_wire_4955;
    wire new_Jinkela_wire_2871;
    wire new_Jinkela_wire_7445;
    wire new_Jinkela_wire_7794;
    wire new_Jinkela_wire_7176;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_2561;
    wire new_Jinkela_wire_6286;
    wire _0098_;
    wire _0240_;
    wire new_Jinkela_wire_6775;
    wire new_Jinkela_wire_4425;
    wire new_Jinkela_wire_2832;
    wire new_Jinkela_wire_2645;
    wire new_Jinkela_wire_3191;
    wire new_Jinkela_wire_3520;
    wire new_Jinkela_wire_7849;
    wire new_Jinkela_wire_2580;
    wire new_Jinkela_wire_4715;
    wire new_Jinkela_wire_7871;
    wire new_Jinkela_wire_4831;
    wire new_Jinkela_wire_1765;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_2907;
    wire new_Jinkela_wire_6513;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_1840;
    wire new_Jinkela_wire_3390;
    wire _0615_;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_7933;
    wire new_Jinkela_wire_2707;
    wire new_Jinkela_wire_6997;
    wire new_Jinkela_wire_7719;
    wire new_Jinkela_wire_7633;
    wire new_Jinkela_wire_5766;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_5023;
    wire _0119_;
    wire new_Jinkela_wire_4498;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_4959;
    wire new_Jinkela_wire_3887;
    wire new_Jinkela_wire_5475;
    wire new_Jinkela_wire_7253;
    wire new_Jinkela_wire_3402;
    wire new_Jinkela_wire_2852;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_2166;
    wire new_Jinkela_wire_1900;
    wire new_Jinkela_wire_6703;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_5240;
    wire _0449_;
    wire new_Jinkela_wire_7897;
    wire _1178_;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_3367;
    wire new_Jinkela_wire_288;
    wire _0352_;
    wire _0731_;
    wire new_Jinkela_wire_2867;
    wire new_Jinkela_wire_4122;
    wire _0468_;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_6071;
    wire _0049_;
    wire new_Jinkela_wire_2156;
    wire new_Jinkela_wire_3166;
    wire new_Jinkela_wire_5575;
    wire _0041_;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_5048;
    wire new_Jinkela_wire_7998;
    wire new_Jinkela_wire_6916;
    wire new_Jinkela_wire_5158;
    wire new_Jinkela_wire_6240;
    wire new_Jinkela_wire_3546;
    wire new_Jinkela_wire_4308;
    wire new_Jinkela_wire_3001;
    wire new_Jinkela_wire_7188;
    wire new_Jinkela_wire_5942;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_3731;
    wire new_Jinkela_wire_6713;
    wire new_Jinkela_wire_3872;
    wire new_Jinkela_wire_3203;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_3100;
    wire new_Jinkela_wire_7709;
    wire new_Jinkela_wire_4158;
    wire new_Jinkela_wire_2950;
    wire new_Jinkela_wire_7877;
    wire new_Jinkela_wire_7334;
    wire _0343_;
    wire new_Jinkela_wire_5495;
    wire _0812_;
    wire new_Jinkela_wire_4095;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_3507;
    wire new_Jinkela_wire_3360;
    wire new_Jinkela_wire_4523;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_7376;
    wire new_Jinkela_wire_2433;
    wire new_Jinkela_wire_2027;
    wire new_Jinkela_wire_2517;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_4291;
    wire new_Jinkela_wire_4101;
    wire new_Jinkela_wire_6255;
    wire new_Jinkela_wire_6404;
    wire _1207_;
    wire new_Jinkela_wire_1749;
    wire _0084_;
    wire new_Jinkela_wire_3929;
    wire new_Jinkela_wire_3351;
    wire _0672_;
    wire new_net_2423;
    wire new_Jinkela_wire_7472;
    wire new_Jinkela_wire_5250;
    wire _0861_;
    wire new_Jinkela_wire_4043;
    wire new_Jinkela_wire_5450;
    wire new_Jinkela_wire_3523;
    wire new_Jinkela_wire_3431;
    wire new_Jinkela_wire_7259;
    wire _0583_;
    wire new_Jinkela_wire_470;
    wire _0221_;
    wire new_Jinkela_wire_6873;
    wire new_Jinkela_wire_4086;
    wire new_Jinkela_wire_3494;
    wire new_Jinkela_wire_5659;
    wire new_Jinkela_wire_7454;
    wire new_Jinkela_wire_2128;
    wire _0043_;
    wire new_Jinkela_wire_4042;
    wire _0741_;
    wire new_Jinkela_wire_108;
    wire _0316_;
    wire new_Jinkela_wire_2082;
    wire new_Jinkela_wire_4475;
    wire new_Jinkela_wire_3648;
    wire new_Jinkela_wire_4632;
    wire _0756_;
    wire new_Jinkela_wire_4383;
    wire new_Jinkela_wire_2795;
    wire _0643_;
    wire new_Jinkela_wire_6622;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_7177;
    wire new_Jinkela_wire_6438;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_3436;
    wire _0485_;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_3283;
    wire new_Jinkela_wire_7718;
    wire new_Jinkela_wire_6905;
    wire new_Jinkela_wire_3931;
    wire new_Jinkela_wire_3086;
    wire new_Jinkela_wire_1913;
    wire new_Jinkela_wire_5927;
    wire new_Jinkela_wire_6968;
    wire new_Jinkela_wire_3801;
    wire new_Jinkela_wire_7254;
    wire new_Jinkela_wire_5679;
    wire new_Jinkela_wire_3487;
    wire new_Jinkela_wire_6429;
    wire new_Jinkela_wire_6700;
    wire new_Jinkela_wire_4608;
    wire new_Jinkela_wire_2179;
    wire new_Jinkela_wire_7453;
    wire new_Jinkela_wire_2061;
    wire new_Jinkela_wire_2059;
    wire new_Jinkela_wire_7980;
    wire new_Jinkela_wire_1930;
    wire new_Jinkela_wire_7179;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_5274;
    wire new_Jinkela_wire_7461;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_2488;
    wire new_Jinkela_wire_6401;
    wire new_Jinkela_wire_7490;
    wire new_Jinkela_wire_6850;
    wire _0748_;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_2949;
    wire new_Jinkela_wire_2152;
    wire new_Jinkela_wire_4003;
    wire new_Jinkela_wire_4461;
    wire new_Jinkela_wire_2172;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_8010;
    wire new_Jinkela_wire_6750;
    wire new_net_26;
    wire new_Jinkela_wire_5257;
    wire new_Jinkela_wire_2984;
    wire new_Jinkela_wire_3205;
    wire new_Jinkela_wire_6421;
    wire new_Jinkela_wire_6424;
    wire _0589_;
    wire new_Jinkela_wire_1781;
    wire new_Jinkela_wire_1083;
    wire _0467_;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_6981;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_4501;
    wire new_net_2461;
    wire new_Jinkela_wire_5391;
    wire new_Jinkela_wire_6484;
    wire new_Jinkela_wire_7117;
    wire new_Jinkela_wire_7781;
    wire new_Jinkela_wire_3946;
    wire new_Jinkela_wire_5757;
    wire new_Jinkela_wire_7775;
    wire _1163_;
    wire new_Jinkela_wire_5508;
    wire new_Jinkela_wire_5059;
    wire new_Jinkela_wire_2827;
    wire new_Jinkela_wire_1698;
    wire new_Jinkela_wire_6377;
    wire new_Jinkela_wire_152;
    wire new_net_2359;
    wire _0807_;
    wire new_Jinkela_wire_6555;
    wire new_Jinkela_wire_4673;
    wire new_Jinkela_wire_6977;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_6081;
    wire new_Jinkela_wire_263;
    wire _0170_;
    wire new_Jinkela_wire_6371;
    wire new_Jinkela_wire_2874;
    wire new_Jinkela_wire_5126;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_4554;
    wire new_Jinkela_wire_7010;
    wire new_Jinkela_wire_685;
    wire _0924_;
    wire new_Jinkela_wire_6627;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_5814;
    wire new_Jinkela_wire_4824;
    wire new_Jinkela_wire_5665;
    wire new_Jinkela_wire_4006;
    wire _0437_;
    wire new_Jinkela_wire_4305;
    wire _0339_;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_7755;
    wire new_Jinkela_wire_930;
    wire new_net_2391;
    wire _0788_;
    wire new_Jinkela_wire_3258;
    wire _0586_;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_2716;
    wire new_Jinkela_wire_2058;
    wire new_Jinkela_wire_6554;
    wire new_Jinkela_wire_6598;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_3041;
    wire new_Jinkela_wire_2120;
    wire new_Jinkela_wire_5581;
    wire new_Jinkela_wire_7778;
    wire new_Jinkela_wire_5356;
    wire new_Jinkela_wire_4458;
    wire new_Jinkela_wire_5592;
    wire new_Jinkela_wire_2240;
    wire new_Jinkela_wire_7058;
    wire new_Jinkela_wire_4300;
    wire new_Jinkela_wire_5895;
    wire new_Jinkela_wire_7809;
    wire new_Jinkela_wire_2307;
    wire new_Jinkela_wire_7736;
    wire new_Jinkela_wire_140;
    wire _1237_;
    wire _0668_;
    wire new_Jinkela_wire_7130;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_4556;
    wire new_Jinkela_wire_7494;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_5245;
    wire new_Jinkela_wire_2861;
    wire new_Jinkela_wire_5752;
    wire new_net_2393;
    wire new_Jinkela_wire_3967;
    wire new_Jinkela_wire_5289;
    wire new_Jinkela_wire_2923;
    wire new_Jinkela_wire_6690;
    wire new_Jinkela_wire_3481;
    wire new_Jinkela_wire_7487;
    wire new_Jinkela_wire_5815;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_2210;
    wire new_Jinkela_wire_7308;
    wire new_Jinkela_wire_5586;
    wire new_Jinkela_wire_184;
    wire _0626_;
    wire new_Jinkela_wire_5565;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_6517;
    wire new_Jinkela_wire_3728;
    wire new_Jinkela_wire_3447;
    wire new_Jinkela_wire_3738;
    wire new_Jinkela_wire_6006;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_6136;
    wire new_Jinkela_wire_6231;
    wire _0064_;
    wire new_Jinkela_wire_4812;
    wire new_Jinkela_wire_7107;
    wire new_Jinkela_wire_1908;
    wire _0656_;
    wire new_Jinkela_wire_3914;
    wire _0495_;
    wire new_net_2361;
    wire new_Jinkela_wire_3652;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_5455;
    wire new_Jinkela_wire_3296;
    wire new_Jinkela_wire_4114;
    wire new_Jinkela_wire_5533;
    wire new_Jinkela_wire_7990;
    wire new_Jinkela_wire_6069;
    wire new_Jinkela_wire_5139;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_1405;
    wire new_Jinkela_wire_7154;
    wire new_Jinkela_wire_3122;
    wire new_Jinkela_wire_5004;
    wire new_Jinkela_wire_3227;
    wire new_Jinkela_wire_5544;
    wire new_Jinkela_wire_7511;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_3293;
    wire new_Jinkela_wire_1742;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_4734;
    wire new_Jinkela_wire_5335;
    wire new_Jinkela_wire_5331;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_5859;
    wire new_Jinkela_wire_3477;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_4615;
    wire _0536_;
    wire new_Jinkela_wire_4578;
    wire _0982_;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_2734;
    wire new_Jinkela_wire_4451;
    wire new_Jinkela_wire_2811;
    wire new_Jinkela_wire_3852;
    wire new_Jinkela_wire_4739;
    wire new_Jinkela_wire_7649;
    wire new_Jinkela_wire_3043;
    wire new_Jinkela_wire_1475;
    wire new_Jinkela_wire_2688;
    wire new_Jinkela_wire_3678;
    wire _1169_;
    wire new_Jinkela_wire_2625;
    wire new_Jinkela_wire_2705;
    wire new_Jinkela_wire_2467;
    wire new_Jinkela_wire_5325;
    wire _1157_;
    wire new_Jinkela_wire_5799;
    wire new_Jinkela_wire_5598;
    wire new_Jinkela_wire_870;
    wire _1079_;
    wire new_Jinkela_wire_4102;
    wire new_Jinkela_wire_4982;
    wire new_Jinkela_wire_3034;
    wire new_Jinkela_wire_631;
    wire _0273_;
    wire new_Jinkela_wire_5635;
    wire new_Jinkela_wire_3471;
    wire new_Jinkela_wire_5657;
    wire new_Jinkela_wire_6479;
    wire new_Jinkela_wire_6902;
    wire new_Jinkela_wire_3886;
    wire new_Jinkela_wire_2392;
    wire new_Jinkela_wire_5393;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_5498;
    wire new_Jinkela_wire_6199;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_4024;
    wire new_Jinkela_wire_1782;
    wire _1009_;
    wire new_Jinkela_wire_6298;
    wire new_Jinkela_wire_6577;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_6748;
    wire new_Jinkela_wire_5333;
    wire new_Jinkela_wire_7168;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_5445;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_7760;
    wire new_Jinkela_wire_2607;
    wire new_Jinkela_wire_2898;
    wire new_Jinkela_wire_5838;
    wire new_Jinkela_wire_7984;
    wire new_Jinkela_wire_6915;
    wire new_Jinkela_wire_6117;
    wire _0534_;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_1880;
    wire new_Jinkela_wire_7242;
    wire _1230_;
    wire new_Jinkela_wire_2908;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_5145;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_5986;
    wire new_Jinkela_wire_2905;
    wire new_Jinkela_wire_5313;
    wire new_Jinkela_wire_7100;
    wire new_Jinkela_wire_6954;
    wire new_Jinkela_wire_5506;
    wire new_Jinkela_wire_4858;
    wire new_Jinkela_wire_2429;
    wire _0852_;
    wire new_Jinkela_wire_6611;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_4511;
    wire new_Jinkela_wire_6953;
    wire _0828_;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_4787;
    wire new_Jinkela_wire_3566;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_7657;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_5297;
    wire new_Jinkela_wire_6790;
    wire _1243_;
    wire _0299_;
    wire new_Jinkela_wire_5064;
    wire new_Jinkela_wire_5278;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_7353;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_6067;
    wire new_Jinkela_wire_6917;
    wire new_Jinkela_wire_2039;
    wire new_Jinkela_wire_6234;
    wire _0318_;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_7301;
    wire _0728_;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_5542;
    wire new_Jinkela_wire_2969;
    wire _0938_;
    wire _0601_;
    wire new_Jinkela_wire_4363;
    wire new_Jinkela_wire_2108;
    wire new_Jinkela_wire_6425;
    wire new_Jinkela_wire_5561;
    wire new_Jinkela_wire_3921;
    wire new_Jinkela_wire_7867;
    wire _0903_;
    wire new_Jinkela_wire_2319;
    wire new_Jinkela_wire_2970;
    wire new_Jinkela_wire_2611;
    wire new_Jinkela_wire_4237;
    wire new_Jinkela_wire_3306;
    wire new_Jinkela_wire_2145;
    wire _0428_;
    wire new_Jinkela_wire_7526;
    wire _0533_;
    wire new_Jinkela_wire_5078;
    wire new_Jinkela_wire_2695;
    wire new_Jinkela_wire_1888;
    wire new_Jinkela_wire_5577;
    wire new_Jinkela_wire_4173;
    wire new_Jinkela_wire_7275;
    wire new_Jinkela_wire_3890;
    wire new_Jinkela_wire_3621;
    wire new_Jinkela_wire_7349;
    wire new_Jinkela_wire_3459;
    wire new_Jinkela_wire_3848;
    wire new_Jinkela_wire_5580;
    wire new_Jinkela_wire_6093;
    wire new_Jinkela_wire_6290;
    wire _0646_;
    wire _0295_;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_3072;
    wire _0350_;
    wire new_Jinkela_wire_2477;
    wire new_Jinkela_wire_2808;
    wire _0167_;
    wire new_Jinkela_wire_3619;
    wire new_Jinkela_wire_2404;
    wire new_Jinkela_wire_4651;
    wire new_Jinkela_wire_7893;
    wire new_Jinkela_wire_3107;
    wire new_Jinkela_wire_6366;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_1823;
    wire new_Jinkela_wire_4154;
    wire new_Jinkela_wire_887;
    wire _0515_;
    wire new_Jinkela_wire_7944;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_5404;
    wire new_net_2397;
    wire new_Jinkela_wire_2431;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_3058;
    wire new_Jinkela_wire_2956;
    wire new_Jinkela_wire_5897;
    wire _0215_;
    wire new_Jinkela_wire_6264;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_4047;
    wire new_Jinkela_wire_6711;
    wire new_Jinkela_wire_2314;
    wire new_Jinkela_wire_3201;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_2509;
    wire new_Jinkela_wire_5134;
    wire new_Jinkela_wire_6940;
    wire new_Jinkela_wire_7545;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_7982;
    wire new_Jinkela_wire_3932;
    wire _0700_;
    wire new_Jinkela_wire_4630;
    wire new_Jinkela_wire_5497;
    wire new_Jinkela_wire_3963;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_2457;
    wire new_Jinkela_wire_2005;
    wire new_Jinkela_wire_6295;
    wire new_Jinkela_wire_6730;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_7283;
    wire new_Jinkela_wire_5364;
    wire new_Jinkela_wire_5314;
    wire new_Jinkela_wire_2013;
    wire _0284_;
    wire new_Jinkela_wire_6207;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_2318;
    wire _0926_;
    wire new_Jinkela_wire_6904;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_1151;
    wire new_Jinkela_wire_3746;
    wire _0840_;
    wire new_Jinkela_wire_5155;
    wire new_Jinkela_wire_1957;
    wire new_Jinkela_wire_7745;
    wire new_Jinkela_wire_2840;
    wire new_Jinkela_wire_3753;
    wire _0290_;
    wire _0612_;
    wire new_Jinkela_wire_2723;
    wire new_Jinkela_wire_3579;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_6165;
    wire new_Jinkela_wire_2738;
    wire _1139_;
    wire new_Jinkela_wire_6031;
    wire _0139_;
    wire new_Jinkela_wire_5030;
    wire new_Jinkela_wire_4577;
    wire new_Jinkela_wire_6311;
    wire _0032_;
    wire _0280_;
    wire new_Jinkela_wire_6844;
    wire new_Jinkela_wire_4289;
    wire new_Jinkela_wire_4493;
    wire new_Jinkela_wire_2859;
    wire new_Jinkela_wire_6064;
    wire new_Jinkela_wire_5763;
    wire new_Jinkela_wire_5140;
    wire new_Jinkela_wire_5593;
    wire new_Jinkela_wire_4275;
    wire new_Jinkela_wire_7525;
    wire new_Jinkela_wire_2343;
    wire new_Jinkela_wire_7390;
    wire _0510_;
    wire _1206_;
    wire new_Jinkela_wire_4481;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_5013;
    wire new_Jinkela_wire_5348;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_2976;
    wire new_Jinkela_wire_4773;
    wire new_Jinkela_wire_6669;
    wire new_Jinkela_wire_2247;
    wire new_Jinkela_wire_3679;
    wire new_Jinkela_wire_2677;
    wire new_Jinkela_wire_3382;
    wire new_Jinkela_wire_4808;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_7378;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_5136;
    wire new_net_2467;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_3877;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_6437;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_554;
    wire _0344_;
    wire new_Jinkela_wire_3482;
    wire new_Jinkela_wire_6482;
    wire new_Jinkela_wire_3898;
    wire new_Jinkela_wire_6395;
    wire new_net_2389;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_2500;
    wire _0156_;
    wire new_Jinkela_wire_7393;
    wire _0604_;
    wire new_Jinkela_wire_1567;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_5332;
    wire new_Jinkela_wire_2643;
    wire new_Jinkela_wire_3473;
    wire new_Jinkela_wire_2154;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_7398;
    wire _0685_;
    wire new_Jinkela_wire_4997;
    wire new_Jinkela_wire_3287;
    wire new_Jinkela_wire_5309;
    wire new_Jinkela_wire_6280;
    wire new_Jinkela_wire_6723;
    wire new_Jinkela_wire_6318;
    wire new_Jinkela_wire_2599;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_5342;
    wire new_Jinkela_wire_7306;
    wire _1146_;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_4232;
    wire _1209_;
    wire _0191_;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_5627;
    wire new_Jinkela_wire_5867;
    wire new_Jinkela_wire_5553;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_2759;
    wire new_Jinkela_wire_4036;
    wire new_Jinkela_wire_6083;
    wire _0068_;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_5975;
    wire new_Jinkela_wire_5846;
    wire new_Jinkela_wire_3469;
    wire new_Jinkela_wire_5731;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_7143;
    wire new_Jinkela_wire_4970;
    wire new_Jinkela_wire_6346;
    wire new_Jinkela_wire_2090;
    wire new_Jinkela_wire_6564;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_7019;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_4520;
    wire new_Jinkela_wire_1084;
    wire _1106_;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_2717;
    wire new_Jinkela_wire_7256;
    wire new_Jinkela_wire_7622;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_4533;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_7036;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_3235;
    wire new_Jinkela_wire_7171;
    wire new_Jinkela_wire_6353;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_4503;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_2983;
    wire _0746_;
    wire new_Jinkela_wire_7320;
    wire new_Jinkela_wire_5793;
    wire new_Jinkela_wire_4245;
    wire new_Jinkela_wire_4319;
    wire new_Jinkela_wire_3796;
    wire new_Jinkela_wire_4622;
    wire _0721_;
    wire new_Jinkela_wire_5076;
    wire new_Jinkela_wire_2419;
    wire _1192_;
    wire new_Jinkela_wire_3661;
    wire new_Jinkela_wire_4854;
    wire _0422_;
    wire _0112_;
    wire new_Jinkela_wire_1691;
    wire new_Jinkela_wire_6153;
    wire new_Jinkela_wire_6074;
    wire new_Jinkela_wire_2612;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_5704;
    wire new_Jinkela_wire_4402;
    wire new_net_18;
    wire new_Jinkela_wire_7694;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_5666;
    wire new_Jinkela_wire_5178;
    wire new_Jinkela_wire_2624;
    wire new_Jinkela_wire_6036;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_7762;
    wire new_Jinkela_wire_310;
    wire _0336_;
    wire new_Jinkela_wire_2271;
    wire _0569_;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_6803;
    wire _0556_;
    wire new_Jinkela_wire_1368;
    wire _0489_;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_4911;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_4643;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_6895;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_7562;
    wire new_Jinkela_wire_3879;
    wire _1059_;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_3363;
    wire _0674_;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_27;
    wire _1016_;
    wire new_Jinkela_wire_1689;
    wire new_Jinkela_wire_7479;
    wire new_Jinkela_wire_3550;
    wire new_Jinkela_wire_4217;
    wire new_Jinkela_wire_2532;
    wire new_Jinkela_wire_6119;
    wire new_Jinkela_wire_2965;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_5466;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_2669;
    wire new_Jinkela_wire_6570;
    wire new_Jinkela_wire_7749;
    wire _0940_;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_7110;
    wire _0706_;
    wire new_Jinkela_wire_2458;
    wire _0649_;
    wire new_Jinkela_wire_7132;
    wire new_Jinkela_wire_6417;
    wire _0809_;
    wire new_Jinkela_wire_3598;
    wire new_Jinkela_wire_2245;
    wire new_Jinkela_wire_5980;
    wire new_Jinkela_wire_626;
    wire _0471_;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_3162;
    wire new_Jinkela_wire_3406;
    wire _0532_;
    wire new_Jinkela_wire_6928;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_1918;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_3769;
    wire new_Jinkela_wire_4418;
    wire _1066_;
    wire new_Jinkela_wire_5493;
    wire new_Jinkela_wire_7740;
    wire new_Jinkela_wire_6568;
    wire _0785_;
    wire new_Jinkela_wire_5347;
    wire new_Jinkela_wire_6130;
    wire new_Jinkela_wire_2466;
    wire new_Jinkela_wire_3916;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_7105;
    wire new_Jinkela_wire_153;
    wire _0482_;
    wire new_Jinkela_wire_5120;
    wire new_Jinkela_wire_2144;
    wire new_Jinkela_wire_2077;
    wire new_Jinkela_wire_5065;
    wire new_Jinkela_wire_3780;
    wire new_Jinkela_wire_6061;
    wire new_Jinkela_wire_4903;
    wire new_Jinkela_wire_585;
    wire _0648_;
    wire new_Jinkela_wire_3683;
    wire new_Jinkela_wire_4369;
    wire new_Jinkela_wire_2105;
    wire new_Jinkela_wire_2430;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_7396;
    wire new_Jinkela_wire_5912;
    wire new_Jinkela_wire_2765;
    wire new_Jinkela_wire_2629;
    wire new_Jinkela_wire_6689;
    wire _1115_;
    wire new_Jinkela_wire_6692;
    wire new_Jinkela_wire_2401;
    wire new_Jinkela_wire_5762;
    wire new_Jinkela_wire_2857;
    wire new_Jinkela_wire_7828;
    wire new_Jinkela_wire_7573;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_2097;
    wire new_Jinkela_wire_7747;
    wire new_Jinkela_wire_4147;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_7662;
    wire new_Jinkela_wire_7481;
    wire _0050_;
    wire new_Jinkela_wire_4035;
    wire new_Jinkela_wire_4422;
    wire new_Jinkela_wire_5106;
    wire _0562_;
    wire new_Jinkela_wire_2057;
    wire new_Jinkela_wire_6768;
    wire new_Jinkela_wire_3139;
    wire new_Jinkela_wire_2541;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_4759;
    wire new_Jinkela_wire_7608;
    wire new_Jinkela_wire_7347;
    wire new_Jinkela_wire_6464;
    wire new_Jinkela_wire_5548;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_2063;
    wire new_Jinkela_wire_2324;
    wire new_Jinkela_wire_7227;
    wire new_Jinkela_wire_5529;
    wire new_Jinkela_wire_6732;
    wire new_Jinkela_wire_6396;
    wire new_Jinkela_wire_6472;
    wire new_Jinkela_wire_3432;
    wire new_Jinkela_wire_7780;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_7094;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_3771;
    wire new_Jinkela_wire_7620;
    wire new_Jinkela_wire_4396;
    wire new_Jinkela_wire_4168;
    wire new_Jinkela_wire_4145;
    wire new_Jinkela_wire_7631;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_4385;
    wire _0107_;
    wire _0764_;
    wire new_Jinkela_wire_4279;
    wire new_Jinkela_wire_4055;
    wire new_Jinkela_wire_5954;
    wire new_Jinkela_wire_2111;
    wire new_Jinkela_wire_6596;
    wire new_Jinkela_wire_6534;
    wire new_Jinkela_wire_5865;
    wire new_Jinkela_wire_3131;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_7854;
    wire _0566_;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_7166;
    wire new_Jinkela_wire_6712;
    wire _0275_;
    wire new_Jinkela_wire_4595;
    wire _0600_;
    wire new_Jinkela_wire_2727;
    wire new_Jinkela_wire_7951;
    wire new_Jinkela_wire_2883;
    wire _1121_;
    wire new_Jinkela_wire_5970;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_7230;
    wire new_Jinkela_wire_3805;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_2854;
    wire new_Jinkela_wire_5571;
    wire new_Jinkela_wire_6181;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_2954;
    wire new_Jinkela_wire_2254;
    wire new_Jinkela_wire_6574;
    wire new_Jinkela_wire_5441;
    wire new_Jinkela_wire_5451;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_3577;
    wire new_Jinkela_wire_6190;
    wire _0900_;
    wire new_Jinkela_wire_4428;
    wire new_Jinkela_wire_6393;
    wire new_Jinkela_wire_6506;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_3142;
    wire new_Jinkela_wire_7425;
    wire new_Jinkela_wire_1828;
    wire _0210_;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_3023;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_3777;
    wire new_Jinkela_wire_5462;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_6185;
    wire new_Jinkela_wire_5849;
    wire new_Jinkela_wire_2916;
    wire new_Jinkela_wire_6120;
    wire _0946_;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_6789;
    wire new_Jinkela_wire_5107;
    wire new_Jinkela_wire_7181;
    wire new_Jinkela_wire_4334;
    wire new_Jinkela_wire_5939;
    wire _0017_;
    wire _0269_;
    wire new_Jinkela_wire_1996;
    wire new_Jinkela_wire_5869;
    wire _1123_;
    wire _0159_;
    wire new_Jinkela_wire_5562;
    wire new_Jinkela_wire_6047;
    wire new_Jinkela_wire_2068;
    wire new_Jinkela_wire_5499;
    wire new_Jinkela_wire_3050;
    wire new_Jinkela_wire_5371;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_6907;
    wire new_Jinkela_wire_2345;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_4273;
    wire new_Jinkela_wire_7039;
    wire new_Jinkela_wire_3804;
    wire new_Jinkela_wire_3305;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_4789;
    wire new_Jinkela_wire_3190;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_6261;
    wire _0158_;
    wire new_Jinkela_wire_7395;
    wire new_Jinkela_wire_3800;
    wire new_Jinkela_wire_4921;
    wire new_Jinkela_wire_7460;
    wire _0022_;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_6462;
    wire new_Jinkela_wire_6465;
    wire new_Jinkela_wire_5633;
    wire new_Jinkela_wire_5358;
    wire _0860_;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_5336;
    wire new_Jinkela_wire_1729;
    wire new_Jinkela_wire_6974;
    wire new_Jinkela_wire_2426;
    wire new_Jinkela_wire_1333;
    wire _0404_;
    wire _0889_;
    wire new_Jinkela_wire_3860;
    wire new_Jinkela_wire_3394;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_5176;
    wire new_Jinkela_wire_1990;
    wire new_Jinkela_wire_5172;
    wire new_Jinkela_wire_6680;
    wire new_Jinkela_wire_2283;
    wire new_Jinkela_wire_7604;
    wire new_Jinkela_wire_3140;
    wire new_Jinkela_wire_2603;
    wire new_Jinkela_wire_5077;
    wire _0991_;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_2578;
    wire new_Jinkela_wire_4944;
    wire new_Jinkela_wire_3750;
    wire _0511_;
    wire new_Jinkela_wire_2704;
    wire new_Jinkela_wire_6569;
    wire new_Jinkela_wire_6876;
    wire new_net_2497;
    wire new_Jinkela_wire_7261;
    wire new_Jinkela_wire_1241;
    wire _1075_;
    wire new_Jinkela_wire_7136;
    wire _0431_;
    wire new_Jinkela_wire_5960;
    wire new_Jinkela_wire_5719;
    wire new_Jinkela_wire_5982;
    wire _0059_;
    wire _0024_;
    wire new_Jinkela_wire_2640;
    wire _0254_;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_6363;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_7455;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_4034;
    wire _1223_;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_4278;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_4008;
    wire new_Jinkela_wire_5617;
    wire new_Jinkela_wire_1897;
    wire new_Jinkela_wire_3725;
    wire new_Jinkela_wire_4411;
    wire new_Jinkela_wire_6657;
    wire new_Jinkela_wire_5239;
    wire new_Jinkela_wire_7589;
    wire new_Jinkela_wire_2296;
    wire _0271_;
    wire new_Jinkela_wire_3782;
    wire _1219_;
    wire new_Jinkela_wire_4022;
    wire _0627_;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_3399;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_6058;
    wire new_Jinkela_wire_7795;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_5079;
    wire new_Jinkela_wire_4287;
    wire new_Jinkela_wire_3557;
    wire _0285_;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_5988;
    wire new_Jinkela_wire_7959;
    wire new_Jinkela_wire_1951;
    wire new_Jinkela_wire_7891;
    wire new_Jinkela_wire_2405;
    wire _0078_;
    wire new_Jinkela_wire_2463;
    wire new_Jinkela_wire_1860;
    wire new_Jinkela_wire_5957;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_4202;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_2987;
    wire new_Jinkela_wire_7784;
    wire new_Jinkela_wire_3667;
    wire _0301_;
    wire _1181_;
    wire new_Jinkela_wire_6966;
    wire new_Jinkela_wire_4664;
    wire new_Jinkela_wire_7539;
    wire new_Jinkela_wire_2920;
    wire new_Jinkela_wire_1734;
    wire new_Jinkela_wire_4993;
    wire new_Jinkela_wire_3138;
    wire new_Jinkela_wire_7673;
    wire new_Jinkela_wire_3952;
    wire new_Jinkela_wire_4559;
    wire new_Jinkela_wire_4558;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_6683;
    wire new_Jinkela_wire_4258;
    wire new_Jinkela_wire_2234;
    wire new_Jinkela_wire_5215;
    wire new_Jinkela_wire_2794;
    wire new_Jinkela_wire_6129;
    wire new_Jinkela_wire_3160;
    wire _0629_;
    wire new_Jinkela_wire_3917;
    wire new_Jinkela_wire_2474;
    wire _0052_;
    wire new_Jinkela_wire_1676;
    wire _0034_;
    wire new_Jinkela_wire_3244;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_6934;
    wire new_Jinkela_wire_3415;
    wire new_Jinkela_wire_4066;
    wire new_Jinkela_wire_2305;
    wire new_Jinkela_wire_3511;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_2147;
    wire _0712_;
    wire new_Jinkela_wire_5247;
    wire new_Jinkela_wire_3681;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_3127;
    wire new_Jinkela_wire_4302;
    wire new_Jinkela_wire_4347;
    wire _0922_;
    wire new_Jinkela_wire_3578;
    wire new_Jinkela_wire_7278;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_4159;
    wire new_Jinkela_wire_2558;
    wire new_Jinkela_wire_6529;
    wire new_Jinkela_wire_7066;
    wire new_Jinkela_wire_1972;
    wire new_Jinkela_wire_2494;
    wire new_Jinkela_wire_6758;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_3491;
    wire new_Jinkela_wire_4667;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_4156;
    wire new_Jinkela_wire_7498;
    wire new_Jinkela_wire_2222;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_7841;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_7091;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_7483;
    wire new_Jinkela_wire_3321;
    wire _0381_;
    wire new_Jinkela_wire_2726;
    wire _1033_;
    wire new_Jinkela_wire_8017;
    wire new_Jinkela_wire_2527;
    wire new_Jinkela_wire_7469;
    wire new_Jinkela_wire_1984;
    wire _0219_;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_4687;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_5265;
    wire new_Jinkela_wire_6594;
    wire new_Jinkela_wire_5692;
    wire new_Jinkela_wire_2048;
    wire new_Jinkela_wire_6057;
    wire new_Jinkela_wire_7686;
    wire new_Jinkela_wire_3272;
    wire _0145_;
    wire _0776_;
    wire new_Jinkela_wire_6430;
    wire new_Jinkela_wire_4561;
    wire _0460_;
    wire _0881_;
    wire _0143_;
    wire new_Jinkela_wire_7609;
    wire new_Jinkela_wire_4740;
    wire new_Jinkela_wire_3253;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_2663;
    wire _0869_;
    wire new_Jinkela_wire_7675;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_4907;
    wire new_Jinkela_wire_1315;
    wire _0206_;
    wire new_Jinkela_wire_3435;
    wire new_Jinkela_wire_7497;
    wire _1215_;
    wire new_net_2449;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_1893;
    wire new_Jinkela_wire_3741;
    wire _0830_;
    wire _0892_;
    wire new_Jinkela_wire_2870;
    wire new_Jinkela_wire_2203;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_5993;
    wire new_Jinkela_wire_3934;
    wire new_Jinkela_wire_4785;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_4565;
    wire _1229_;
    wire new_Jinkela_wire_1953;
    wire new_Jinkela_wire_2130;
    wire new_Jinkela_wire_5058;
    wire new_Jinkela_wire_5427;
    wire new_Jinkela_wire_2306;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_3180;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_6909;
    wire new_Jinkela_wire_7576;
    wire new_Jinkela_wire_5343;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_4847;
    wire new_Jinkela_wire_1092;
    wire _0057_;
    wire new_Jinkela_wire_3957;
    wire new_Jinkela_wire_7086;
    wire new_Jinkela_wire_6516;
    wire new_Jinkela_wire_4509;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_3660;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_3154;
    wire new_Jinkela_wire_5730;
    wire new_Jinkela_wire_5113;
    wire new_Jinkela_wire_2729;
    wire new_Jinkela_wire_3152;
    wire new_Jinkela_wire_5852;
    wire new_Jinkela_wire_1748;
    wire _0967_;
    wire new_Jinkela_wire_6591;
    wire new_Jinkela_wire_3101;
    wire new_Jinkela_wire_2091;
    wire new_Jinkela_wire_5235;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_7839;
    wire new_Jinkela_wire_3558;
    wire new_Jinkela_wire_4276;
    wire new_Jinkela_wire_5607;
    wire new_Jinkela_wire_5464;
    wire new_Jinkela_wire_6345;
    wire new_Jinkela_wire_7707;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_3623;
    wire new_Jinkela_wire_2491;
    wire _0798_;
    wire new_Jinkela_wire_6593;
    wire new_Jinkela_wire_4286;
    wire new_Jinkela_wire_3995;
    wire new_Jinkela_wire_3970;
    wire new_Jinkela_wire_7981;
    wire new_Jinkela_wire_6877;
    wire new_Jinkela_wire_4694;
    wire new_Jinkela_wire_4398;
    wire new_Jinkela_wire_3620;
    wire new_Jinkela_wire_5449;
    wire _0997_;
    wire new_Jinkela_wire_6094;
    wire _0669_;
    wire new_Jinkela_wire_6539;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_3575;
    wire new_Jinkela_wire_4707;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_6962;
    wire _0434_;
    wire new_Jinkela_wire_3576;
    wire new_Jinkela_wire_2772;
    wire new_Jinkela_wire_2622;
    wire new_Jinkela_wire_6612;
    wire new_Jinkela_wire_2577;
    wire new_Jinkela_wire_3941;
    wire new_Jinkela_wire_4623;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_2310;
    wire _0585_;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_3778;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_5097;
    wire _0579_;
    wire _0608_;
    wire new_Jinkela_wire_3635;
    wire new_Jinkela_wire_2498;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_7005;
    wire new_Jinkela_wire_4084;
    wire new_Jinkela_wire_5636;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_2596;
    wire new_Jinkela_wire_6213;
    wire _0864_;
    wire new_Jinkela_wire_5360;
    wire new_Jinkela_wire_4067;
    wire new_Jinkela_wire_7906;
    wire new_Jinkela_wire_3506;
    wire new_Jinkela_wire_562;
    wire _1065_;
    wire new_Jinkela_wire_2584;
    wire new_Jinkela_wire_1737;
    wire new_Jinkela_wire_510;
    wire _0073_;
    wire new_Jinkela_wire_7890;
    wire new_Jinkela_wire_7583;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_1497;
    wire _0407_;
    wire new_Jinkela_wire_3337;
    wire new_Jinkela_wire_4026;
    wire new_Jinkela_wire_7596;
    wire new_Jinkela_wire_7683;
    wire new_Jinkela_wire_4943;
    wire new_Jinkela_wire_6722;
    wire _0913_;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_4984;
    wire new_Jinkela_wire_5395;
    wire new_Jinkela_wire_6504;
    wire new_Jinkela_wire_2129;
    wire new_Jinkela_wire_5863;
    wire _0998_;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_5945;
    wire _1071_;
    wire new_Jinkela_wire_7819;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_7851;
    wire new_Jinkela_wire_3391;
    wire new_Jinkela_wire_3919;
    wire new_Jinkela_wire_4440;
    wire new_Jinkela_wire_3214;
    wire _0875_;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_3336;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_2525;
    wire new_Jinkela_wire_6364;
    wire new_Jinkela_wire_7993;
    wire new_Jinkela_wire_7237;
    wire new_net_2471;
    wire new_Jinkela_wire_5821;
    wire _0877_;
    wire new_Jinkela_wire_2912;
    wire new_Jinkela_wire_4220;
    wire new_Jinkela_wire_7001;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_5108;
    wire new_Jinkela_wire_6020;
    wire new_Jinkela_wire_5834;
    wire new_Jinkela_wire_2706;
    wire new_Jinkela_wire_2294;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_2714;
    wire new_Jinkela_wire_3960;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_6223;
    wire new_Jinkela_wire_2014;
    wire _0714_;
    wire new_Jinkela_wire_3569;
    wire _0274_;
    wire new_Jinkela_wire_6201;
    wire new_Jinkela_wire_4889;
    wire new_Jinkela_wire_6260;
    wire new_Jinkela_wire_7882;
    wire _0341_;
    wire new_Jinkela_wire_6936;
    wire new_Jinkela_wire_1787;
    wire new_Jinkela_wire_4284;
    wire new_Jinkela_wire_6807;
    wire new_Jinkela_wire_5921;
    wire new_Jinkela_wire_7632;
    wire new_Jinkela_wire_6422;
    wire new_Jinkela_wire_4599;
    wire new_Jinkela_wire_7996;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_3332;
    wire new_Jinkela_wire_7403;
    wire new_Jinkela_wire_2506;
    wire new_Jinkela_wire_2255;
    wire _0288_;
    wire new_Jinkela_wire_6707;
    wire new_Jinkela_wire_5680;
    wire new_Jinkela_wire_2432;
    wire new_Jinkela_wire_3231;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_2865;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_5550;
    wire new_Jinkela_wire_1853;
    wire _0435_;
    wire _0307_;
    wire new_Jinkela_wire_6553;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_6897;
    wire new_Jinkela_wire_7187;
    wire new_Jinkela_wire_8012;
    wire new_Jinkela_wire_7956;
    wire new_Jinkela_wire_5870;
    wire new_Jinkela_wire_5181;
    wire new_Jinkela_wire_5424;
    wire new_Jinkela_wire_4727;
    wire new_Jinkela_wire_3133;
    wire new_net_21;
    wire new_Jinkela_wire_6196;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_7554;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_2935;
    wire new_Jinkela_wire_4587;
    wire new_Jinkela_wire_6173;
    wire new_Jinkela_wire_3790;
    wire new_Jinkela_wire_3631;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_3110;
    wire new_Jinkela_wire_7692;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_3693;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_3690;
    wire new_Jinkela_wire_3983;
    wire new_Jinkela_wire_5484;
    wire new_Jinkela_wire_4355;
    wire new_Jinkela_wire_2325;
    wire new_Jinkela_wire_7727;
    wire new_Jinkela_wire_6829;
    wire _1196_;
    wire new_Jinkela_wire_1800;
    wire _0450_;
    wire new_Jinkela_wire_4848;
    wire new_Jinkela_wire_6337;
    wire new_Jinkela_wire_3677;
    wire new_Jinkela_wire_2287;
    wire new_Jinkela_wire_150;
    wire _0042_;
    wire new_Jinkela_wire_6269;
    wire new_Jinkela_wire_6040;
    wire new_Jinkela_wire_5842;
    wire new_Jinkela_wire_6770;
    wire new_Jinkela_wire_4088;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_3853;
    wire new_Jinkela_wire_3045;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_6356;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_1899;
    wire _0045_;
    wire new_Jinkela_wire_7681;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_3366;
    wire new_Jinkela_wire_6236;
    wire new_Jinkela_wire_2747;
    wire _0805_;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_7991;
    wire new_Jinkela_wire_3213;
    wire new_Jinkela_wire_5868;
    wire _0572_;
    wire new_Jinkela_wire_5338;
    wire new_Jinkela_wire_7553;
    wire new_Jinkela_wire_4915;
    wire new_Jinkela_wire_3416;
    wire _0732_;
    wire new_Jinkela_wire_5648;
    wire new_Jinkela_wire_5724;
    wire new_Jinkela_wire_4879;
    wire new_Jinkela_wire_5100;
    wire _0106_;
    wire new_Jinkela_wire_4104;
    wire new_Jinkela_wire_4939;
    wire new_Jinkela_wire_2743;
    wire new_Jinkela_wire_7532;
    wire new_Jinkela_wire_6449;
    wire new_Jinkela_wire_4838;
    wire _0837_;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_6192;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_7382;
    wire new_Jinkela_wire_7713;
    wire new_Jinkela_wire_6522;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_3784;
    wire new_Jinkela_wire_4356;
    wire new_Jinkela_wire_5401;
    wire new_Jinkela_wire_5950;
    wire new_Jinkela_wire_4033;
    wire new_Jinkela_wire_7317;
    wire new_Jinkela_wire_2821;
    wire new_Jinkela_wire_5810;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_4128;
    wire new_Jinkela_wire_3308;
    wire new_Jinkela_wire_4589;
    wire new_Jinkela_wire_2459;
    wire new_Jinkela_wire_5999;
    wire new_Jinkela_wire_5209;
    wire _1007_;
    wire new_Jinkela_wire_2614;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_4646;
    wire new_Jinkela_wire_7613;
    wire new_Jinkela_wire_7383;
    wire new_Jinkela_wire_6793;
    wire new_Jinkela_wire_5093;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_6856;
    wire new_Jinkela_wire_2610;
    wire new_Jinkela_wire_4384;
    wire new_Jinkela_wire_2045;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_5259;
    wire new_Jinkela_wire_6728;
    wire new_Jinkela_wire_2173;
    wire new_Jinkela_wire_5141;
    wire _0400_;
    wire new_Jinkela_wire_7411;
    wire new_Jinkela_wire_5270;
    wire new_Jinkela_wire_1807;
    wire _0121_;
    wire new_Jinkela_wire_2781;
    wire new_Jinkela_wire_4770;
    wire new_Jinkela_wire_4435;
    wire new_Jinkela_wire_2675;
    wire new_Jinkela_wire_7985;
    wire new_Jinkela_wire_7637;
    wire new_Jinkela_wire_6163;
    wire new_Jinkela_wire_3549;
    wire new_Jinkela_wire_7185;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_6879;
    wire new_Jinkela_wire_7533;
    wire new_Jinkela_wire_4109;
    wire new_Jinkela_wire_2915;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_5989;
    wire new_Jinkela_wire_7149;
    wire new_Jinkela_wire_2850;
    wire new_Jinkela_wire_2070;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_4267;
    wire new_Jinkela_wire_4989;
    wire new_Jinkela_wire_3505;
    wire new_Jinkela_wire_6444;
    wire _1105_;
    wire new_Jinkela_wire_6476;
    wire new_Jinkela_wire_2946;
    wire _1214_;
    wire new_Jinkela_wire_1630;
    wire new_Jinkela_wire_3422;
    wire new_Jinkela_wire_6457;
    wire new_Jinkela_wire_4064;
    wire new_Jinkela_wire_2914;
    wire new_Jinkela_wire_1924;
    wire new_Jinkela_wire_5012;
    wire new_Jinkela_wire_3008;
    wire new_Jinkela_wire_5302;
    wire new_Jinkela_wire_7510;
    wire new_Jinkela_wire_3369;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_4297;
    wire new_Jinkela_wire_3688;
    wire new_Jinkela_wire_2639;
    wire new_Jinkela_wire_4116;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_7071;
    wire new_Jinkela_wire_2547;
    wire _0960_;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_1014;
    wire _1063_;
    wire _1177_;
    wire new_Jinkela_wire_3038;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_2461;
    wire new_Jinkela_wire_2814;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_1255;
    wire _0909_;
    wire new_Jinkela_wire_6866;
    wire _0901_;
    wire new_Jinkela_wire_6552;
    wire _0895_;
    wire new_Jinkela_wire_7106;
    wire new_Jinkela_wire_7126;
    wire _1064_;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_6964;
    wire new_Jinkela_wire_1626;
    wire new_Jinkela_wire_198;
    wire _0683_;
    wire new_Jinkela_wire_5777;
    wire new_Jinkela_wire_7792;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_4964;
    wire new_Jinkela_wire_2313;
    wire new_Jinkela_wire_6979;
    wire new_Jinkela_wire_7786;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_5779;
    wire new_Jinkela_wire_7758;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_3187;
    wire new_Jinkela_wire_7076;
    wire new_Jinkela_wire_5334;
    wire _0857_;
    wire new_Jinkela_wire_6696;
    wire new_Jinkela_wire_6589;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_2472;
    wire new_Jinkela_wire_7808;
    wire _0664_;
    wire new_Jinkela_wire_1619;
    wire _0394_;
    wire new_Jinkela_wire_2230;
    wire new_Jinkela_wire_5110;
    wire new_Jinkela_wire_2038;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_5984;
    wire _0186_;
    wire new_Jinkela_wire_7211;
    wire new_Jinkela_wire_6537;
    wire _0633_;
    wire _0425_;
    wire new_Jinkela_wire_7754;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_6725;
    wire _0066_;
    wire new_Jinkela_wire_5368;
    wire new_Jinkela_wire_5847;
    wire new_Jinkela_wire_2073;
    wire new_Jinkela_wire_6911;
    wire new_Jinkela_wire_3478;
    wire new_Jinkela_wire_6912;
    wire new_Jinkela_wire_2791;
    wire new_Jinkela_wire_6548;
    wire new_Jinkela_wire_5197;
    wire _0129_;
    wire new_Jinkela_wire_4314;
    wire new_Jinkela_wire_5601;
    wire new_Jinkela_wire_3241;
    wire new_net_2363;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_30;
    wire _0433_;
    wire new_Jinkela_wire_4712;
    wire new_Jinkela_wire_7354;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_5203;
    wire new_Jinkela_wire_7738;
    wire new_Jinkela_wire_7914;
    wire _0025_;
    wire new_Jinkela_wire_2887;
    wire new_Jinkela_wire_6761;
    wire _0238_;
    wire new_Jinkela_wire_2155;
    wire new_Jinkela_wire_5760;
    wire _0007_;
    wire new_Jinkela_wire_4670;
    wire new_Jinkela_wire_7549;
    wire new_Jinkela_wire_6858;
    wire _0919_;
    wire new_Jinkela_wire_2328;
    wire new_Jinkela_wire_3454;
    wire new_Jinkela_wire_5353;
    wire new_Jinkela_wire_1995;
    wire _0056_;
    wire new_Jinkela_wire_4153;
    wire _0292_;
    wire _0282_;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_4752;
    wire new_Jinkela_wire_3299;
    wire new_net_2511;
    wire new_net_2435;
    wire new_Jinkela_wire_3372;
    wire _1140_;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_4243;
    wire new_Jinkela_wire_2609;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_3128;
    wire new_Jinkela_wire_4618;
    wire new_Jinkela_wire_7236;
    wire new_Jinkela_wire_6910;
    wire new_Jinkela_wire_5749;
    wire new_Jinkela_wire_6828;
    wire new_Jinkela_wire_7121;
    wire new_Jinkela_wire_6716;
    wire new_Jinkela_wire_3895;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_7641;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_2446;
    wire new_Jinkela_wire_2064;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_5953;
    wire _0324_;
    wire new_Jinkela_wire_6671;
    wire new_Jinkela_wire_5200;
    wire new_Jinkela_wire_5856;
    wire new_Jinkela_wire_3834;
    wire new_Jinkela_wire_6128;
    wire _0051_;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_7561;
    wire new_Jinkela_wire_5216;
    wire new_Jinkela_wire_450;
    wire _0131_;
    wire new_Jinkela_wire_3386;
    wire new_Jinkela_wire_2921;
    wire new_Jinkela_wire_2334;
    wire new_Jinkela_wire_6284;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_7292;
    wire new_Jinkela_wire_2450;
    wire new_Jinkela_wire_2253;
    wire new_Jinkela_wire_7837;
    wire _0959_;
    wire new_Jinkela_wire_2227;
    wire new_Jinkela_wire_5840;
    wire new_Jinkela_wire_7325;
    wire new_Jinkela_wire_5923;
    wire new_Jinkela_wire_3615;
    wire new_Jinkela_wire_2348;
    wire new_Jinkela_wire_4062;
    wire new_Jinkela_wire_2837;
    wire _0072_;
    wire new_net_2491;
    wire new_Jinkela_wire_6442;
    wire new_Jinkela_wire_4604;
    wire new_Jinkela_wire_6024;
    wire new_Jinkela_wire_2289;
    wire new_Jinkela_wire_5397;
    wire new_net_2469;
    wire new_Jinkela_wire_6068;
    wire new_Jinkela_wire_3344;
    wire new_Jinkela_wire_3695;
    wire new_Jinkela_wire_4131;
    wire new_Jinkela_wire_5643;
    wire new_Jinkela_wire_1632;
    wire _0790_;
    wire new_Jinkela_wire_2749;
    wire new_Jinkela_wire_7442;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_4553;
    wire new_Jinkela_wire_2127;
    wire _0893_;
    wire _0854_;
    wire new_Jinkela_wire_1319;
    wire new_net_25;
    wire new_Jinkela_wire_7350;
    wire new_Jinkela_wire_5962;
    wire new_Jinkela_wire_5798;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_5940;
    wire new_Jinkela_wire_7436;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_3352;
    wire new_Jinkela_wire_4778;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_2757;
    wire _0329_;
    wire new_Jinkela_wire_5436;
    wire new_Jinkela_wire_2102;
    wire new_Jinkela_wire_5207;
    wire new_Jinkela_wire_7420;
    wire new_Jinkela_wire_4485;
    wire new_Jinkela_wire_3685;
    wire new_Jinkela_wire_5711;
    wire new_Jinkela_wire_1712;
    wire _0118_;
    wire new_Jinkela_wire_6849;
    wire new_Jinkela_wire_5361;
    wire _0884_;
    wire new_Jinkela_wire_6224;
    wire _0916_;
    wire new_Jinkela_wire_7063;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_1097;
    wire _1132_;
    wire _0099_;
    wire new_Jinkela_wire_2503;
    wire new_Jinkela_wire_7863;
    wire _0421_;
    wire new_Jinkela_wire_5184;
    wire new_Jinkela_wire_7920;
    wire new_Jinkela_wire_2771;
    wire _1041_;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_5587;
    wire new_Jinkela_wire_1755;
    wire new_Jinkela_wire_1771;
    wire _0825_;
    wire new_Jinkela_wire_4226;
    wire new_Jinkela_wire_7333;
    wire _1218_;
    wire _0291_;
    wire _0439_;
    wire new_Jinkela_wire_7431;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_3742;
    wire new_Jinkela_wire_5934;
    wire _0811_;
    wire new_Jinkela_wire_897;
    wire new_net_2401;
    wire new_Jinkela_wire_4815;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_2165;
    wire _0092_;
    wire _0868_;
    wire _0456_;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_4909;
    wire new_Jinkela_wire_4716;
    wire new_Jinkela_wire_2071;
    wire new_Jinkela_wire_6959;
    wire new_Jinkela_wire_3930;
    wire new_Jinkela_wire_7764;
    wire new_Jinkela_wire_6780;
    wire new_Jinkela_wire_7602;
    wire new_Jinkela_wire_6679;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_6823;
    wire new_Jinkela_wire_3245;
    wire new_Jinkela_wire_6742;
    wire _0722_;
    wire new_Jinkela_wire_3543;
    wire new_Jinkela_wire_4352;
    wire new_Jinkela_wire_4332;
    wire _0935_;
    wire new_Jinkela_wire_5811;
    wire new_Jinkela_wire_2660;
    wire new_Jinkela_wire_6416;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_4948;
    wire new_Jinkela_wire_4766;
    wire new_Jinkela_wire_7743;
    wire _0239_;
    wire new_Jinkela_wire_7294;
    wire _1022_;
    wire new_Jinkela_wire_2666;
    wire new_Jinkela_wire_4628;
    wire new_Jinkela_wire_3702;
    wire new_Jinkela_wire_4741;
    wire _0849_;
    wire new_Jinkela_wire_1878;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_3755;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_7857;
    wire new_Jinkela_wire_5062;
    wire _0496_;
    wire new_Jinkela_wire_1018;
    wire _0887_;
    wire new_Jinkela_wire_3137;
    wire new_Jinkela_wire_2824;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_2473;
    wire new_Jinkela_wire_2762;
    wire new_Jinkela_wire_2843;
    wire new_Jinkela_wire_7661;
    wire new_Jinkela_wire_3202;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_4386;
    wire new_Jinkela_wire_2689;
    wire new_Jinkela_wire_4358;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_7339;
    wire new_Jinkela_wire_6735;
    wire new_Jinkela_wire_2918;
    wire new_Jinkela_wire_6305;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_3044;
    wire new_Jinkela_wire_7797;
    wire new_Jinkela_wire_6814;
    wire new_Jinkela_wire_3596;
    wire _0213_;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_7628;
    wire new_Jinkela_wire_1941;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_4295;
    wire new_Jinkela_wire_2670;
    wire new_Jinkela_wire_5468;
    wire new_Jinkela_wire_3005;
    wire new_Jinkela_wire_3488;
    wire new_Jinkela_wire_5116;
    wire new_Jinkela_wire_1869;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_3125;
    wire new_Jinkela_wire_7582;
    wire _0670_;
    wire new_Jinkela_wire_2846;
    wire new_Jinkela_wire_2703;
    wire new_Jinkela_wire_4666;
    wire new_Jinkela_wire_3174;
    wire new_Jinkela_wire_3793;
    wire new_Jinkela_wire_2878;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_5955;
    wire new_Jinkela_wire_7338;
    wire new_Jinkela_wire_7611;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_2752;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_7524;
    wire new_Jinkela_wire_4199;
    wire new_Jinkela_wire_2993;
    wire new_Jinkela_wire_2174;
    wire new_Jinkela_wire_7412;
    wire new_Jinkela_wire_3117;
    wire _0190_;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_3609;
    wire new_Jinkela_wire_3922;
    wire new_Jinkela_wire_5536;
    wire new_Jinkela_wire_3825;
    wire new_Jinkela_wire_6156;
    wire _0635_;
    wire new_Jinkela_wire_3155;
    wire _0740_;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_5969;
    wire new_Jinkela_wire_6454;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_3026;
    wire new_Jinkela_wire_6271;
    wire new_Jinkela_wire_3843;
    wire new_Jinkela_wire_2056;
    wire new_Jinkela_wire_8007;
    wire new_Jinkela_wire_5623;
    wire new_Jinkela_wire_2279;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_5317;
    wire new_Jinkela_wire_1962;
    wire new_Jinkela_wire_5009;
    wire new_Jinkela_wire_4992;
    wire new_Jinkela_wire_5233;
    wire new_Jinkela_wire_6491;
    wire new_Jinkela_wire_7263;
    wire new_Jinkela_wire_7222;
    wire new_Jinkela_wire_4764;
    wire new_Jinkela_wire_4987;
    wire new_Jinkela_wire_6602;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_2836;
    wire new_Jinkela_wire_4843;
    wire new_Jinkela_wire_6125;
    wire new_Jinkela_wire_7423;
    wire _0588_;
    wire _0046_;
    wire new_net_2505;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_7287;
    wire _0418_;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_3327;
    wire _0117_;
    wire new_Jinkela_wire_7629;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_3103;
    wire new_Jinkela_wire_2608;
    wire new_Jinkela_wire_7725;
    wire new_Jinkela_wire_3495;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_7402;
    wire _0075_;
    wire new_Jinkela_wire_6200;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_7002;
    wire new_Jinkela_wire_6558;
    wire new_Jinkela_wire_7614;
    wire new_Jinkela_wire_4935;
    wire new_Jinkela_wire_4688;
    wire new_Jinkela_wire_2873;
    wire _0015_;
    wire new_Jinkela_wire_5833;
    wire new_Jinkela_wire_2400;
    wire new_net_2415;
    wire _0555_;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_6709;
    wire new_net_19;
    wire new_Jinkela_wire_4412;
    wire new_Jinkela_wire_6980;
    wire new_Jinkela_wire_6660;
    wire new_Jinkela_wire_3981;
    wire new_Jinkela_wire_6625;
    wire new_Jinkela_wire_5089;
    wire new_Jinkela_wire_4802;
    wire new_Jinkela_wire_7766;
    wire new_Jinkela_wire_4130;
    wire new_Jinkela_wire_7414;
    wire _0976_;
    wire new_Jinkela_wire_2522;
    wire new_Jinkela_wire_2375;
    wire _0923_;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_2451;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_4899;
    wire new_Jinkela_wire_7902;
    wire new_Jinkela_wire_2713;
    wire new_Jinkela_wire_1722;
    wire new_Jinkela_wire_7123;
    wire new_Jinkela_wire_4517;
    wire new_Jinkela_wire_6217;
    wire _0754_;
    wire _1136_;
    wire new_Jinkela_wire_279;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_3676;
    wire new_Jinkela_wire_7007;
    wire new_Jinkela_wire_7697;
    wire new_Jinkela_wire_6413;
    wire new_Jinkela_wire_4486;
    wire new_Jinkela_wire_4830;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_7477;
    wire new_Jinkela_wire_2309;
    wire _0266_;
    wire new_Jinkela_wire_3027;
    wire new_Jinkela_wire_7006;
    wire new_Jinkela_wire_7032;
    wire new_Jinkela_wire_4894;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_6018;
    wire new_Jinkela_wire_4502;
    wire new_Jinkela_wire_3474;
    wire new_Jinkela_wire_1016;
    wire new_Jinkela_wire_7180;
    wire _0673_;
    wire _1205_;
    wire new_Jinkela_wire_2739;
    wire new_Jinkela_wire_2952;
    wire new_Jinkela_wire_4508;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_7986;
    wire _1231_;
    wire new_Jinkela_wire_4381;
    wire new_Jinkela_wire_2162;
    wire new_Jinkela_wire_6805;
    wire new_Jinkela_wire_2702;
    wire new_Jinkela_wire_5208;
    wire new_Jinkela_wire_4985;
    wire new_Jinkela_wire_3665;
    wire new_Jinkela_wire_3659;
    wire new_Jinkela_wire_4610;
    wire new_Jinkela_wire_3682;
    wire _1142_;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_5535;
    wire _0727_;
    wire new_Jinkela_wire_2489;
    wire new_Jinkela_wire_7836;
    wire new_Jinkela_wire_7590;
    wire new_Jinkela_wire_5252;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_4700;
    wire new_Jinkela_wire_5041;
    wire _0929_;
    wire new_Jinkela_wire_4092;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_6230;
    wire new_Jinkela_wire_3582;
    wire new_Jinkela_wire_7976;
    wire new_Jinkela_wire_3295;
    wire new_Jinkela_wire_2550;
    wire new_Jinkela_wire_4443;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_4908;
    wire new_Jinkela_wire_1647;
    wire _0490_;
    wire new_Jinkela_wire_7218;
    wire new_Jinkela_wire_5511;
    wire new_Jinkela_wire_7899;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_1817;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_4452;
    wire new_Jinkela_wire_3705;
    wire new_Jinkela_wire_1693;
    wire new_Jinkela_wire_1963;
    wire new_Jinkela_wire_3395;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_3021;
    wire new_Jinkela_wire_2773;
    wire new_Jinkela_wire_2903;
    wire new_Jinkela_wire_2862;
    wire new_Jinkela_wire_5883;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_895;
    wire new_net_2409;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_3109;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_7367;
    wire new_Jinkela_wire_5772;
    wire new_Jinkela_wire_2241;
    wire new_Jinkela_wire_7077;
    wire new_Jinkela_wire_4132;
    wire new_Jinkela_wire_7084;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_4689;
    wire new_Jinkela_wire_6854;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_5418;
    wire _0770_;
    wire _0641_;
    wire new_Jinkela_wire_6358;
    wire new_Jinkela_wire_5722;
    wire new_Jinkela_wire_5538;
    wire _0546_;
    wire _1036_;
    wire new_Jinkela_wire_7043;
    wire _0730_;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_523;
    wire _0521_;
    wire new_Jinkela_wire_5189;
    wire new_Jinkela_wire_5411;
    wire new_Jinkela_wire_4683;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_4377;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_6387;
    wire new_Jinkela_wire_5363;
    wire new_Jinkela_wire_6228;
    wire new_Jinkela_wire_6785;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_357;
    wire _0541_;
    wire _0996_;
    wire new_Jinkela_wire_4311;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_3123;
    wire new_net_7;
    wire _0208_;
    wire new_Jinkela_wire_3484;
    wire _0617_;
    wire new_Jinkela_wire_4839;
    wire _0647_;
    wire new_Jinkela_wire_1852;
    wire new_Jinkela_wire_2533;
    wire new_Jinkela_wire_5459;
    wire new_Jinkela_wire_4890;
    wire new_Jinkela_wire_4494;
    wire new_Jinkela_wire_4096;
    wire new_Jinkela_wire_4322;
    wire new_Jinkela_wire_7134;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_7815;
    wire new_Jinkela_wire_2581;
    wire new_Jinkela_wire_4505;
    wire new_Jinkela_wire_3430;
    wire new_Jinkela_wire_6003;
    wire new_Jinkela_wire_6618;
    wire new_Jinkela_wire_3880;
    wire new_Jinkela_wire_3439;
    wire new_Jinkela_wire_6206;
    wire new_Jinkela_wire_5217;
    wire new_Jinkela_wire_5880;
    wire new_Jinkela_wire_3726;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_4071;
    wire _0618_;
    wire _0171_;
    wire new_Jinkela_wire_4037;
    wire new_Jinkela_wire_6784;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_6507;
    wire new_Jinkela_wire_4679;
    wire _1084_;
    wire new_Jinkela_wire_5202;
    wire new_Jinkela_wire_7087;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_6308;
    wire new_Jinkela_wire_3183;
    wire new_Jinkela_wire_5822;
    wire new_Jinkela_wire_3428;
    wire new_Jinkela_wire_2644;
    wire new_Jinkela_wire_3217;
    wire new_net_5;
    wire _0027_;
    wire new_Jinkela_wire_2200;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_6194;
    wire new_Jinkela_wire_7352;
    wire _0818_;
    wire new_Jinkela_wire_3510;
    wire new_Jinkela_wire_5481;
    wire new_Jinkela_wire_6166;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_4392;
    wire new_Jinkela_wire_8019;
    wire new_Jinkela_wire_7534;
    wire new_Jinkela_wire_2069;
    wire new_Jinkela_wire_5918;
    wire new_Jinkela_wire_5470;
    wire new_Jinkela_wire_3636;
    wire _0765_;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_5807;
    wire new_Jinkela_wire_4097;
    wire new_Jinkela_wire_4028;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_1656;
    wire _0300_;
    wire new_Jinkela_wire_6766;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_3452;
    wire new_Jinkela_wire_3814;
    wire _0524_;
    wire new_Jinkela_wire_5020;
    wire new_Jinkela_wire_5710;
    wire new_Jinkela_wire_6781;
    wire new_Jinkela_wire_7443;
    wire new_Jinkela_wire_7092;
    wire new_Jinkela_wire_5525;
    wire new_Jinkela_wire_5787;
    wire new_Jinkela_wire_3884;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_4856;
    wire new_Jinkela_wire_114;
    wire _0398_;
    wire new_Jinkela_wire_5329;
    wire new_Jinkela_wire_7850;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_4931;
    wire _0323_;
    wire new_Jinkela_wire_5983;
    wire new_Jinkela_wire_3810;
    wire _0523_;
    wire new_Jinkela_wire_147;
    wire new_net_2411;
    wire new_Jinkela_wire_6313;
    wire new_Jinkela_wire_6375;
    wire new_Jinkela_wire_5655;
    wire new_Jinkela_wire_6041;
    wire new_Jinkela_wire_4013;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_8013;
    wire new_Jinkela_wire_4809;
    wire _0477_;
    wire new_Jinkela_wire_4916;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_3533;
    wire new_Jinkela_wire_2183;
    wire new_Jinkela_wire_4421;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_5249;
    wire new_Jinkela_wire_6937;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_5557;
    wire _1185_;
    wire new_Jinkela_wire_5727;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_1040;
    wire new_Jinkela_wire_7823;
    wire new_Jinkela_wire_2080;
    wire new_Jinkela_wire_4263;
    wire new_Jinkela_wire_1309;
    wire new_Jinkela_wire_7322;
    wire new_Jinkela_wire_1278;
    wire _0843_;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_6737;
    wire new_Jinkela_wire_69;
    wire _0607_;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_1294;
    wire new_Jinkela_wire_4583;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_4852;
    wire new_Jinkela_wire_7721;
    wire new_Jinkela_wire_1713;
    wire new_Jinkela_wire_7285;
    wire _0564_;
    wire _1203_;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_6023;
    wire _0382_;
    wire new_net_2429;
    wire new_Jinkela_wire_2568;
    wire new_Jinkela_wire_6542;
    wire new_Jinkela_wire_6149;
    wire new_Jinkela_wire_5745;
    wire new_Jinkela_wire_6210;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_5898;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_2864;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_4876;
    wire new_Jinkela_wire_7638;
    wire new_Jinkela_wire_1258;
    wire _0030_;
    wire new_Jinkela_wire_5809;
    wire new_Jinkela_wire_4078;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_2755;
    wire new_Jinkela_wire_6667;
    wire new_Jinkela_wire_7800;
    wire new_Jinkela_wire_4892;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_2613;
    wire new_Jinkela_wire_3583;
    wire _0596_;
    wire new_Jinkela_wire_6299;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_2034;
    wire _1013_;
    wire new_Jinkela_wire_6272;
    wire new_Jinkela_wire_7040;
    wire new_Jinkela_wire_3276;
    wire new_Jinkela_wire_3686;
    wire new_Jinkela_wire_6944;
    wire new_Jinkela_wire_2897;
    wire _0831_;
    wire new_Jinkela_wire_2168;
    wire new_Jinkela_wire_5055;
    wire new_Jinkela_wire_3434;
    wire new_Jinkela_wire_2117;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_4434;
    wire new_Jinkela_wire_1911;
    wire new_Jinkela_wire_7246;
    wire new_Jinkela_wire_3030;
    wire new_Jinkela_wire_5578;
    wire new_Jinkela_wire_7405;
    wire new_Jinkela_wire_5211;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_5408;
    wire new_Jinkela_wire_4499;
    wire new_Jinkela_wire_3445;
    wire new_Jinkela_wire_3845;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_3906;
    wire new_Jinkela_wire_4986;
    wire new_Jinkela_wire_5564;
    wire new_Jinkela_wire_5728;
    wire new_Jinkela_wire_7971;
    wire _0540_;
    wire _0065_;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_3309;
    wire new_Jinkela_wire_4242;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_5964;
    wire new_Jinkela_wire_3973;
    wire _0380_;
    wire new_Jinkela_wire_4887;
    wire new_Jinkela_wire_6629;
    wire new_Jinkela_wire_5827;
    wire new_Jinkela_wire_2904;
    wire new_Jinkela_wire_4543;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_7544;
    wire new_Jinkela_wire_6802;
    wire new_Jinkela_wire_7621;
    wire new_Jinkela_wire_2618;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_2482;
    wire _0169_;
    wire new_Jinkela_wire_3736;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_3388;
    wire new_Jinkela_wire_6923;
    wire new_Jinkela_wire_3239;
    wire new_Jinkela_wire_6885;
    wire _0694_;
    wire new_Jinkela_wire_6089;
    wire new_Jinkela_wire_7881;
    wire _0964_;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_2376;
    wire new_Jinkela_wire_966;
    wire _0954_;
    wire _0021_;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_2981;
    wire new_Jinkela_wire_7927;
    wire new_Jinkela_wire_4634;
    wire new_net_2357;
    wire new_Jinkela_wire_3888;
    wire new_Jinkela_wire_7340;
    wire _0444_;
    wire _0697_;
    wire new_Jinkela_wire_7862;
    wire new_Jinkela_wire_4568;
    wire new_Jinkela_wire_3501;
    wire new_Jinkela_wire_2719;
    wire _0242_;
    wire _0399_;
    wire new_Jinkela_wire_5060;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_5193;
    wire _0133_;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_5406;
    wire _0715_;
    wire _0761_;
    wire new_Jinkela_wire_3603;
    wire new_Jinkela_wire_6257;
    wire new_Jinkela_wire_5299;
    wire new_Jinkela_wire_5328;
    wire new_Jinkela_wire_7407;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_7342;
    wire new_Jinkela_wire_6604;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_7856;
    wire _0955_;
    wire new_Jinkela_wire_4864;
    wire new_Jinkela_wire_3353;
    wire new_Jinkela_wire_4031;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_3751;
    wire _1024_;
    wire new_Jinkela_wire_6146;
    wire new_Jinkela_wire_3773;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_3630;
    wire new_Jinkela_wire_2668;
    wire new_Jinkela_wire_5963;
    wire new_Jinkela_wire_6587;
    wire new_Jinkela_wire_4127;
    wire new_Jinkela_wire_3561;
    wire _0061_;
    wire new_Jinkela_wire_7889;
    wire new_Jinkela_wire_5537;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_7879;
    wire new_Jinkela_wire_2678;
    wire new_Jinkela_wire_4126;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_3223;
    wire new_Jinkela_wire_4195;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_3976;
    wire new_Jinkela_wire_6322;
    wire new_Jinkela_wire_1780;
    wire new_Jinkela_wire_4805;
    wire _1048_;
    wire _0839_;
    wire new_Jinkela_wire_5349;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_2146;
    wire _0180_;
    wire new_Jinkela_wire_3783;
    wire _0026_;
    wire new_Jinkela_wire_6919;
    wire new_Jinkela_wire_2496;
    wire new_Jinkela_wire_6621;
    wire _0591_;
    wire new_Jinkela_wire_5384;
    wire new_Jinkela_wire_6397;
    wire new_Jinkela_wire_6080;
    wire new_Jinkela_wire_2308;
    wire new_Jinkela_wire_7111;
    wire _0093_;
    wire new_Jinkela_wire_3643;
    wire _0401_;
    wire _0614_;
    wire _1037_;
    wire new_Jinkela_wire_6901;
    wire new_Jinkela_wire_2302;
    wire _0277_;
    wire new_Jinkela_wire_4241;
    wire _0529_;
    wire new_net_2373;
    wire new_Jinkela_wire_5392;
    wire _0311_;
    wire new_Jinkela_wire_7502;
    wire new_Jinkela_wire_2142;
    wire new_Jinkela_wire_6659;
    wire new_Jinkela_wire_3984;
    wire new_Jinkela_wire_2107;
    wire new_Jinkela_wire_3542;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_2708;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_5346;
    wire new_Jinkela_wire_2985;
    wire new_Jinkela_wire_2701;
    wire new_Jinkela_wire_6535;
    wire _0451_;
    wire new_Jinkela_wire_3392;
    wire _1114_;
    wire new_Jinkela_wire_7530;
    wire new_Jinkela_wire_3757;
    wire new_Jinkela_wire_6411;
    wire new_Jinkela_wire_6684;
    wire new_Jinkela_wire_7699;
    wire _0645_;
    wire _0708_;
    wire new_Jinkela_wire_3756;
    wire new_Jinkela_wire_5102;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_6103;
    wire new_Jinkela_wire_2141;
    wire new_Jinkela_wire_2745;
    wire _0152_;
    wire _0986_;
    wire new_Jinkela_wire_492;
    wire _1149_;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_6480;
    wire new_Jinkela_wire_8011;
    wire new_Jinkela_wire_4228;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_2831;
    wire new_Jinkela_wire_5132;
    wire new_Jinkela_wire_7769;
    wire _0934_;
    wire new_Jinkela_wire_6386;
    wire new_Jinkela_wire_3556;
    wire new_Jinkela_wire_6704;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_3234;
    wire new_Jinkela_wire_2425;
    wire new_Jinkela_wire_3074;
    wire _0101_;
    wire new_net_2365;
    wire new_Jinkela_wire_6614;
    wire new_Jinkela_wire_5073;
    wire new_Jinkela_wire_2818;
    wire _0369_;
    wire new_Jinkela_wire_2779;
    wire new_Jinkela_wire_6485;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_5769;
    wire new_Jinkela_wire_5281;
    wire new_Jinkela_wire_6650;
    wire new_Jinkela_wire_4060;
    wire new_Jinkela_wire_3211;
    wire new_Jinkela_wire_2787;
    wire new_Jinkela_wire_3346;
    wire new_Jinkela_wire_4721;
    wire _0517_;
    wire new_Jinkela_wire_6685;
    wire new_Jinkela_wire_5157;
    wire new_Jinkela_wire_1157;
    wire _0870_;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_1252;
    wire _0599_;
    wire new_Jinkela_wire_4753;
    wire _0147_;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_4758;
    wire _0228_;
    wire new_Jinkela_wire_2078;
    wire new_Jinkela_wire_4340;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_4360;
    wire new_Jinkela_wire_4790;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_3497;
    wire new_Jinkela_wire_5936;
    wire _0452_;
    wire new_Jinkela_wire_7370;
    wire _0842_;
    wire new_Jinkela_wire_7493;
    wire _0109_;
    wire new_Jinkela_wire_5416;
    wire new_Jinkela_wire_3856;
    wire new_Jinkela_wire_6250;
    wire new_Jinkela_wire_2637;
    wire new_Jinkela_wire_7999;
    wire new_Jinkela_wire_1792;
    wire new_Jinkela_wire_7938;
    wire new_Jinkela_wire_7089;
    wire new_Jinkela_wire_2033;
    wire new_Jinkela_wire_3053;
    wire new_Jinkela_wire_2602;
    wire new_Jinkela_wire_2524;
    wire new_Jinkela_wire_5843;
    wire new_Jinkela_wire_2942;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_3347;
    wire new_Jinkela_wire_6835;
    wire new_Jinkela_wire_1450;
    wire _1099_;
    wire new_Jinkela_wire_1518;
    wire _0866_;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_3994;
    wire new_Jinkela_wire_2948;
    wire new_Jinkela_wire_7444;
    wire new_Jinkela_wire_7798;
    wire new_Jinkela_wire_4011;
    wire new_Jinkela_wire_5081;
    wire new_Jinkela_wire_1466;
    wire _0423_;
    wire new_Jinkela_wire_6045;
    wire _1053_;
    wire new_Jinkela_wire_4433;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_3881;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_7170;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_6526;
    wire new_Jinkela_wire_3185;
    wire new_Jinkela_wire_6932;
    wire new_Jinkela_wire_6957;
    wire new_Jinkela_wire_7207;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_2440;
    wire _1056_;
    wire new_Jinkela_wire_5042;
    wire new_Jinkela_wire_5483;
    wire new_Jinkela_wire_3999;
    wire new_Jinkela_wire_6865;
    wire _1040_;
    wire new_Jinkela_wire_4743;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_7746;
    wire new_Jinkela_wire_3204;
    wire new_Jinkela_wire_6237;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_6302;
    wire new_Jinkela_wire_7392;
    wire new_Jinkela_wire_6918;
    wire _0853_;
    wire _0011_;
    wire new_Jinkela_wire_6900;
    wire new_Jinkela_wire_5122;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_7212;
    wire new_Jinkela_wire_3216;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_2715;
    wire new_Jinkela_wire_6183;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_5946;
    wire _0990_;
    wire new_Jinkela_wire_2552;
    wire _0334_;
    wire new_Jinkela_wire_4138;
    wire new_Jinkela_wire_7997;
    wire new_Jinkela_wire_5243;
    wire new_Jinkela_wire_6279;
    wire new_Jinkela_wire_3169;
    wire _0941_;
    wire new_Jinkela_wire_4490;
    wire _0142_;
    wire _0973_;
    wire new_Jinkela_wire_5380;
    wire new_Jinkela_wire_4164;
    wire new_Jinkela_wire_6423;
    wire new_Jinkela_wire_4884;
    wire _1145_;
    wire new_Jinkela_wire_7466;
    wire new_Jinkela_wire_7049;
    wire new_Jinkela_wire_4471;
    wire new_Jinkela_wire_7474;
    wire new_Jinkela_wire_335;
    wire _0792_;
    wire new_Jinkela_wire_4569;
    wire new_Jinkela_wire_4405;
    wire new_Jinkela_wire_6338;
    wire new_Jinkela_wire_1300;
    wire _0793_;
    wire new_Jinkela_wire_5686;
    wire new_Jinkela_wire_5177;
    wire new_Jinkela_wire_4326;
    wire new_Jinkela_wire_641;
    wire _0317_;
    wire new_Jinkela_wire_2793;
    wire new_Jinkela_wire_2225;
    wire _0173_;
    wire new_Jinkela_wire_3410;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_6381;
    wire new_Jinkela_wire_6440;
    wire new_Jinkela_wire_4192;
    wire new_Jinkela_wire_2636;
    wire new_Jinkela_wire_4949;
    wire new_Jinkela_wire_7911;
    wire new_Jinkela_wire_7807;
    wire new_Jinkela_wire_2030;
    wire new_Jinkela_wire_6778;
    wire new_Jinkela_wire_3591;
    wire new_Jinkela_wire_4644;
    wire new_Jinkela_wire_3470;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_2761;
    wire new_Jinkela_wire_6973;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_6751;
    wire _1202_;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_5650;
    wire new_Jinkela_wire_4613;
    wire new_Jinkela_wire_3091;
    wire new_Jinkela_wire_7057;
    wire _0518_;
    wire new_Jinkela_wire_5668;
    wire _1015_;
    wire new_Jinkela_wire_7626;
    wire new_Jinkela_wire_5734;
    wire new_Jinkela_wire_5977;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_6022;
    wire new_Jinkela_wire_6955;
    wire new_Jinkela_wire_2664;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_2084;
    wire new_Jinkela_wire_3380;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_2124;
    wire new_Jinkela_wire_7930;
    wire new_Jinkela_wire_3791;
    wire new_Jinkela_wire_2486;
    wire new_Jinkela_wire_7714;
    wire _0779_;
    wire _0723_;
    wire new_Jinkela_wire_6647;
    wire new_Jinkela_wire_7921;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_5881;
    wire new_Jinkela_wire_4567;
    wire _0355_;
    wire new_Jinkela_wire_3301;
    wire new_Jinkela_wire_2798;
    wire new_Jinkela_wire_4709;
    wire new_Jinkela_wire_7827;
    wire new_Jinkela_wire_6694;
    wire new_Jinkela_wire_4283;
    wire new_Jinkela_wire_6118;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_7559;
    wire new_Jinkela_wire_1744;
    wire new_Jinkela_wire_5517;
    wire new_Jinkela_wire_4318;
    wire new_Jinkela_wire_3900;
    wire new_Jinkela_wire_2841;
    wire new_Jinkela_wire_3073;
    wire new_Jinkela_wire_2001;
    wire new_Jinkela_wire_7949;
    wire new_Jinkela_wire_5567;
    wire new_Jinkela_wire_2074;
    wire new_Jinkela_wire_2169;
    wire new_Jinkela_wire_3317;
    wire new_Jinkela_wire_3837;
    wire new_Jinkela_wire_6765;
    wire new_Jinkela_wire_5743;
    wire new_Jinkela_wire_4166;
    wire new_Jinkela_wire_2452;
    wire new_Jinkela_wire_2221;
    wire new_Jinkela_wire_4407;
    wire new_Jinkela_wire_4316;
    wire new_Jinkela_wire_2967;
    wire _0606_;
    wire new_Jinkela_wire_4769;
    wire _1183_;
    wire _1159_;
    wire _0786_;
    wire new_Jinkela_wire_3521;
    wire new_Jinkela_wire_3717;
    wire new_Jinkela_wire_4420;
    wire new_Jinkela_wire_6435;
    wire new_Jinkela_wire_3130;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_3096;
    wire new_Jinkela_wire_4833;
    wire new_Jinkela_wire_4818;
    wire new_Jinkela_wire_2317;
    wire new_Jinkela_wire_3384;
    wire _1045_;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_225;
    wire _0576_;
    wire new_Jinkela_wire_6343;
    wire new_Jinkela_wire_5764;
    wire _0200_;
    wire new_Jinkela_wire_7932;
    wire new_Jinkela_wire_3247;
    wire _0076_;
    wire new_Jinkela_wire_6321;
    wire _1076_;
    wire new_Jinkela_wire_2464;
    wire new_Jinkela_wire_4282;
    wire new_Jinkela_wire_6092;
    wire new_Jinkela_wire_5664;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_3268;
    wire new_Jinkela_wire_7363;
    wire new_Jinkela_wire_2674;
    wire new_Jinkela_wire_3650;
    wire new_Jinkela_wire_7556;
    wire _0008_;
    wire new_Jinkela_wire_5958;
    wire _0577_;
    wire new_Jinkela_wire_5385;
    wire new_Jinkela_wire_7451;
    wire new_Jinkela_wire_4115;
    wire new_Jinkela_wire_2557;
    wire new_Jinkela_wire_2872;
    wire new_Jinkela_wire_5725;
    wire new_Jinkela_wire_4548;
    wire new_Jinkela_wire_2212;
    wire _1190_;
    wire new_Jinkela_wire_2067;
    wire new_Jinkela_wire_5460;
    wire _0862_;
    wire new_Jinkela_wire_5262;
    wire new_Jinkela_wire_5796;
    wire new_Jinkela_wire_7142;
    wire new_Jinkela_wire_3611;
    wire new_Jinkela_wire_3248;
    wire new_Jinkela_wire_3088;
    wire new_Jinkela_wire_3807;
    wire new_Jinkela_wire_7044;
    wire new_Jinkela_wire_2072;
    wire new_Jinkela_wire_6026;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_4476;
    wire new_Jinkela_wire_4919;
    wire _0472_;
    wire new_Jinkela_wire_6390;
    wire new_Jinkela_wire_3196;
    wire new_Jinkela_wire_2758;
    wire _0182_;
    wire new_Jinkela_wire_7083;
    wire new_Jinkela_wire_7512;
    wire new_Jinkela_wire_4238;
    wire new_Jinkela_wire_7859;
    wire new_Jinkela_wire_7763;
    wire new_Jinkela_wire_4742;
    wire new_Jinkela_wire_4906;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_6030;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_5761;
    wire new_Jinkela_wire_7041;
    wire new_Jinkela_wire_7547;
    wire new_Jinkela_wire_3766;
    wire new_Jinkela_wire_5662;
    wire new_Jinkela_wire_3710;
    wire new_Jinkela_wire_4470;
    wire new_Jinkela_wire_2519;
    wire _0912_;
    wire new_Jinkela_wire_4691;
    wire new_net_2451;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_1022;
    wire _0778_;
    wire _0505_;
    wire new_Jinkela_wire_5088;
    wire new_Jinkela_wire_3049;
    wire new_Jinkela_wire_6515;
    wire new_Jinkela_wire_3493;
    wire new_Jinkela_wire_438;
    wire _0613_;
    wire _0176_;
    wire new_Jinkela_wire_3342;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_5018;
    wire new_Jinkela_wire_6002;
    wire new_Jinkela_wire_7234;
    wire new_Jinkela_wire_7038;
    wire _0241_;
    wire new_Jinkela_wire_5049;
    wire new_Jinkela_wire_3149;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_4409;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_7138;
    wire new_Jinkela_wire_3789;
    wire _1204_;
    wire new_Jinkela_wire_6323;
    wire new_Jinkela_wire_2218;
    wire new_Jinkela_wire_6719;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_2062;
    wire new_Jinkela_wire_2737;
    wire new_Jinkela_wire_4236;
    wire _0438_;
    wire new_Jinkela_wire_2523;
    wire _0833_;
    wire _0040_;
    wire new_Jinkela_wire_2628;
    wire new_Jinkela_wire_2092;
    wire new_Jinkela_wire_1238;
    wire _0134_;
    wire new_Jinkela_wire_3862;
    wire new_Jinkela_wire_6819;
    wire new_Jinkela_wire_3333;
    wire new_Jinkela_wire_7220;
    wire _0281_;
    wire new_Jinkela_wire_2806;
    wire new_Jinkela_wire_3607;
    wire new_Jinkela_wire_8005;
    wire _0651_;
    wire new_Jinkela_wire_6754;
    wire new_Jinkela_wire_1917;
    wire new_Jinkela_wire_4862;
    wire new_Jinkela_wire_4477;
    wire new_Jinkela_wire_6607;
    wire new_Jinkela_wire_5626;
    wire new_Jinkela_wire_5540;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_4462;
    wire new_Jinkela_wire_7155;
    wire new_Jinkela_wire_3466;
    wire new_Jinkela_wire_3051;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_2709;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_4564;
    wire new_Jinkela_wire_6469;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_6446;
    wire new_Jinkela_wire_2536;
    wire new_Jinkela_wire_349;
    wire _0630_;
    wire _0653_;
    wire new_Jinkela_wire_4474;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_4627;
    wire new_Jinkela_wire_6764;
    wire new_Jinkela_wire_5105;
    wire _0948_;
    wire new_Jinkela_wire_5034;
    wire _0925_;
    wire new_Jinkela_wire_5781;
    wire new_Jinkela_wire_2652;
    wire new_Jinkela_wire_5968;
    wire new_Jinkela_wire_2562;
    wire _1221_;
    wire new_Jinkela_wire_4519;
    wire new_Jinkela_wire_1747;
    wire new_Jinkela_wire_8000;
    wire new_Jinkela_wire_6815;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_3735;
    wire _0859_;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_2206;
    wire new_Jinkela_wire_4900;
    wire new_Jinkela_wire_6757;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_2958;
    wire new_Jinkela_wire_4974;
    wire _0804_;
    wire new_Jinkela_wire_7935;
    wire new_Jinkela_wire_3330;
    wire _0168_;
    wire new_Jinkela_wire_5695;
    wire new_Jinkela_wire_5688;
    wire new_Jinkela_wire_1786;
    wire new_Jinkela_wire_262;
    wire _0258_;
    wire new_Jinkela_wire_4680;
    wire new_Jinkela_wire_6756;
    wire _0235_;
    wire _0850_;
    wire new_Jinkela_wire_5530;
    wire new_net_2477;
    wire new_Jinkela_wire_4093;
    wire new_Jinkela_wire_7538;
    wire new_Jinkela_wire_5718;
    wire new_Jinkela_wire_7267;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_5223;
    wire _0447_;
    wire new_Jinkela_wire_7097;
    wire _0713_;
    wire new_Jinkela_wire_3987;
    wire new_Jinkela_wire_2476;
    wire new_Jinkela_wire_4902;
    wire _0671_;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_3105;
    wire new_Jinkela_wire_3368;
    wire new_Jinkela_wire_5595;
    wire new_Jinkela_wire_5074;
    wire new_Jinkela_wire_7293;
    wire _0743_;
    wire new_Jinkela_wire_7369;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_5340;
    wire new_Jinkela_wire_4524;
    wire new_Jinkela_wire_2944;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_7486;
    wire new_Jinkela_wire_3823;
    wire new_Jinkela_wire_2132;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_6661;
    wire new_Jinkela_wire_2780;
    wire new_Jinkela_wire_3563;
    wire new_Jinkela_wire_3876;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_4697;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_5916;
    wire new_Jinkela_wire_3262;
    wire new_Jinkela_wire_4837;
    wire _1174_;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_3545;
    wire new_Jinkela_wire_6131;
    wire new_Jinkela_wire_7299;
    wire _0353_;
    wire new_Jinkela_wire_6162;
    wire new_Jinkela_wire_5902;
    wire new_Jinkela_wire_7617;
    wire new_Jinkela_wire_5720;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_2901;
    wire new_Jinkela_wire_5848;
    wire new_Jinkela_wire_2534;
    wire _0395_;
    wire new_Jinkela_wire_5973;
    wire new_Jinkela_wire_7771;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_258;
    wire new_net_2381;
    wire _0537_;
    wire _0545_;
    wire _0931_;
    wire new_Jinkela_wire_4698;
    wire new_Jinkela_wire_7912;
    wire new_Jinkela_wire_7200;
    wire new_Jinkela_wire_2518;
    wire new_Jinkela_wire_3553;
    wire new_Jinkela_wire_7424;
    wire new_Jinkela_wire_1761;
    wire _1154_;
    wire new_net_0;
    wire new_Jinkela_wire_3840;
    wire _1143_;
    wire new_Jinkela_wire_3475;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_2945;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_1491;
    wire new_net_2493;
    wire new_Jinkela_wire_3663;
    wire _1019_;
    wire new_Jinkela_wire_2093;
    wire new_Jinkela_wire_3427;
    wire _0654_;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_7965;
    wire _0652_;
    wire _1195_;
    wire new_Jinkela_wire_2838;
    wire new_Jinkela_wire_4663;
    wire new_Jinkela_wire_1797;
    wire new_Jinkela_wire_4310;
    wire _0220_;
    wire new_Jinkela_wire_3094;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_4585;
    wire new_Jinkela_wire_2330;
    wire new_Jinkela_wire_5337;
    wire new_Jinkela_wire_5797;
    wire new_Jinkela_wire_4219;
    wire new_Jinkela_wire_7146;
    wire new_Jinkela_wire_7210;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_5378;
    wire new_Jinkela_wire_8015;
    wire _0185_;
    wire new_Jinkela_wire_7435;
    wire new_Jinkela_wire_1178;
    wire _0747_;
    wire _0193_;
    wire new_Jinkela_wire_7276;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_6155;
    wire new_Jinkela_wire_4180;
    wire new_Jinkela_wire_3969;
    wire new_Jinkela_wire_2053;
    wire new_Jinkela_wire_5494;
    wire new_Jinkela_wire_497;
    wire _1144_;
    wire new_Jinkela_wire_2320;
    wire new_Jinkela_wire_2504;
    wire new_Jinkela_wire_7178;
    wire _0005_;
    wire new_Jinkela_wire_5388;
    wire new_Jinkela_wire_1286;
    wire new_Jinkela_wire_5311;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_5770;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_3915;
    wire new_Jinkela_wire_3776;
    wire _1027_;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_3359;
    wire new_Jinkela_wire_1420;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_7195;
    wire new_Jinkela_wire_3697;
    wire new_Jinkela_wire_1886;
    wire new_Jinkela_wire_4810;
    wire new_Jinkela_wire_4473;
    wire _0001_;
    wire new_Jinkela_wire_5600;
    wire _0509_;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_2913;
    wire new_Jinkela_wire_3316;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_7064;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_2436;
    wire _0974_;
    wire new_Jinkela_wire_7957;
    wire new_Jinkela_wire_7831;
    wire new_Jinkela_wire_3433;
    wire _1180_;
    wire new_Jinkela_wire_7627;
    wire new_Jinkela_wire_4886;
    wire new_Jinkela_wire_7399;
    wire new_Jinkela_wire_2202;
    wire new_Jinkela_wire_6159;
    wire new_Jinkela_wire_6405;
    wire new_net_27;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_3313;
    wire new_Jinkela_wire_1114;
    wire new_Jinkela_wire_5817;
    wire new_Jinkela_wire_7806;
    wire new_Jinkela_wire_7672;
    wire new_Jinkela_wire_6220;
    wire new_Jinkela_wire_7458;
    wire new_Jinkela_wire_4737;
    wire _0263_;
    wire new_Jinkela_wire_4718;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_2665;
    wire new_Jinkela_wire_5129;
    wire new_Jinkela_wire_6448;
    wire new_Jinkela_wire_5230;
    wire _0508_;
    wire _0153_;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_2778;
    wire new_Jinkela_wire_1037;
    wire new_Jinkela_wire_4397;
    wire new_Jinkela_wire_6869;
    wire new_Jinkela_wire_5503;
    wire new_Jinkela_wire_4507;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_7979;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_2163;
    wire _0725_;
    wire new_Jinkela_wire_5606;
    wire new_Jinkela_wire_7223;
    wire new_Jinkela_wire_5341;
    wire new_Jinkela_wire_5167;
    wire new_Jinkela_wire_739;
    wire _1147_;
    wire new_Jinkela_wire_251;
    wire _1171_;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_5056;
    wire new_Jinkela_wire_4001;
    wire new_Jinkela_wire_3727;
    wire new_Jinkela_wire_3815;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_4204;
    wire new_Jinkela_wire_4206;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_7449;
    wire new_net_2371;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_5288;
    wire new_Jinkela_wire_3141;
    wire new_Jinkela_wire_4954;
    wire new_Jinkela_wire_4980;
    wire new_Jinkela_wire_2094;
    wire new_net_2421;
    wire new_Jinkela_wire_1651;
    wire _0127_;
    wire new_Jinkela_wire_4791;
    wire new_Jinkela_wire_7027;
    wire _0771_;
    wire new_Jinkela_wire_1338;
    wire _0592_;
    wire new_Jinkela_wire_2372;
    wire _0054_;
    wire new_Jinkela_wire_7688;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_4825;
    wire _0742_;
    wire new_Jinkela_wire_2301;
    wire new_Jinkela_wire_7496;
    wire new_Jinkela_wire_6320;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_5440;
    wire new_Jinkela_wire_5933;
    wire new_Jinkela_wire_7194;
    wire _0984_;
    wire new_Jinkela_wire_4073;
    wire new_Jinkela_wire_7814;
    wire new_Jinkela_wire_2369;
    wire new_Jinkela_wire_6077;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_7101;
    wire new_Jinkela_wire_6473;
    wire new_Jinkela_wire_7566;
    wire new_Jinkela_wire_3307;
    wire _0340_;
    wire new_Jinkela_wire_7060;
    wire new_Jinkela_wire_5373;
    wire new_Jinkela_wire_7197;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_4331;
    wire new_Jinkela_wire_5489;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_5045;
    wire new_Jinkela_wire_6121;
    wire new_Jinkela_wire_4792;
    wire new_Jinkela_wire_5147;
    wire new_Jinkela_wire_4861;
    wire new_Jinkela_wire_4832;
    wire new_Jinkela_wire_1848;
    wire _0245_;
    wire new_Jinkela_wire_8016;
    wire new_Jinkela_wire_2891;
    wire new_Jinkela_wire_4995;
    wire _0475_;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_6767;
    wire new_Jinkela_wire_4888;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_6925;
    wire new_Jinkela_wire_7023;
    wire new_Jinkela_wire_5386;
    wire new_Jinkela_wire_4923;
    wire _0823_;
    wire _0187_;
    wire new_Jinkela_wire_4690;
    wire _0278_;
    wire new_Jinkela_wire_6726;
    wire new_Jinkela_wire_7603;
    wire new_Jinkela_wire_6225;
    wire new_Jinkela_wire_4706;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_6774;
    wire new_Jinkela_wire_2344;
    wire new_Jinkela_wire_6428;
    wire new_Jinkela_wire_6787;
    wire new_Jinkela_wire_6300;
    wire new_Jinkela_wire_4573;
    wire new_Jinkela_wire_3743;
    wire new_Jinkela_wire_7148;
    wire new_Jinkela_wire_2642;
    wire new_Jinkela_wire_7595;
    wire new_Jinkela_wire_3745;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_7419;
    wire _0848_;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_6329;
    wire new_Jinkela_wire_4366;
    wire new_Jinkela_wire_2442;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_5488;
    wire new_Jinkela_wire_7400;
    wire new_Jinkela_wire_3868;
    wire new_Jinkela_wire_7782;
    wire new_Jinkela_wire_3326;
    wire new_Jinkela_wire_5502;
    wire new_Jinkela_wire_4662;
    wire new_Jinkela_wire_6171;
    wire new_Jinkela_wire_1421;
    wire new_Jinkela_wire_6123;
    wire new_Jinkela_wire_2938;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_5788;
    wire new_Jinkela_wire_3709;
    wire new_Jinkela_wire_3423;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_7433;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_7818;
    wire new_Jinkela_wire_6011;
    wire new_Jinkela_wire_7987;
    wire new_Jinkela_wire_5226;
    wire new_Jinkela_wire_2593;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_2383;
    wire new_Jinkela_wire_2357;
    wire new_Jinkela_wire_2398;
    wire new_Jinkela_wire_4103;
    wire new_Jinkela_wire_2339;
    wire new_Jinkela_wire_5326;
    wire new_Jinkela_wire_6433;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_4552;
    wire new_Jinkela_wire_3457;
    wire new_Jinkela_wire_6463;
    wire _0315_;
    wire new_Jinkela_wire_5555;
    wire new_Jinkela_wire_2161;
    wire new_Jinkela_wire_951;
    wire _0442_;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_4656;
    wire new_Jinkela_wire_4905;
    wire new_Jinkela_wire_3063;
    wire new_Jinkela_wire_5232;
    wire new_Jinkela_wire_7910;
    wire new_Jinkela_wire_2835;
    wire new_Jinkela_wire_6487;
    wire _0504_;
    wire new_Jinkela_wire_5951;
    wire new_Jinkela_wire_2802;
    wire new_Jinkela_wire_6813;
    wire new_Jinkela_wire_4432;
    wire new_Jinkela_wire_1892;
    wire _0346_;
    wire new_Jinkela_wire_1445;
    wire new_Jinkela_wire_3011;
    wire new_Jinkela_wire_3421;
    wire _1170_;
    wire new_Jinkela_wire_5429;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_5241;
    wire new_Jinkela_wire_3590;
    wire new_Jinkela_wire_5485;
    wire new_Jinkela_wire_4019;
    wire _0012_;
    wire new_Jinkela_wire_5560;
    wire new_Jinkela_wire_2252;
    wire _0980_;
    wire new_Jinkela_wire_7751;
    wire new_Jinkela_wire_4516;
    wire new_Jinkela_wire_7840;
    wire new_Jinkela_wire_3237;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_7654;
    wire new_Jinkela_wire_3286;
    wire new_Jinkela_wire_5610;
    wire _0918_;
    wire new_Jinkela_wire_7535;
    wire new_Jinkela_wire_5191;
    wire new_Jinkela_wire_2018;
    wire new_Jinkela_wire_5027;
    wire new_Jinkela_wire_2101;
    wire new_Jinkela_wire_6514;
    wire new_Jinkela_wire_4870;
    wire _0113_;
    wire new_Jinkela_wire_8020;
    wire new_Jinkela_wire_7866;
    wire new_Jinkela_wire_3670;
    wire new_Jinkela_wire_5915;
    wire new_Jinkela_wire_6004;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_3928;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_1015;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_7572;
    wire new_Jinkela_wire_3646;
    wire new_Jinkela_wire_5350;
    wire new_Jinkela_wire_5707;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_7574;
    wire new_Jinkela_wire_7103;
    wire _0734_;
    wire new_Jinkela_wire_6475;
    wire new_Jinkela_wire_4391;
    wire new_Jinkela_wire_4410;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_6287;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_5431;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_226;
    wire _0690_;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_5425;
    wire new_Jinkela_wire_4655;
    wire _0687_;
    wire new_Jinkela_wire_4920;
    wire new_Jinkela_wire_2103;
    wire new_Jinkela_wire_4210;
    wire new_Jinkela_wire_3124;
    wire new_Jinkela_wire_2312;
    wire new_Jinkela_wire_6441;
    wire new_Jinkela_wire_3339;
    wire new_Jinkela_wire_6654;
    wire new_Jinkela_wire_1398;
    wire new_Jinkela_wire_3826;
    wire new_Jinkela_wire_6995;
    wire new_Jinkela_wire_3338;
    wire new_Jinkela_wire_7739;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_5290;
    wire new_Jinkela_wire_2195;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_5070;
    wire new_Jinkela_wire_5112;
    wire new_Jinkela_wire_2751;
    wire new_Jinkela_wire_6985;
    wire new_Jinkela_wire_2468;
    wire new_Jinkela_wire_5080;
    wire new_Jinkela_wire_6782;
    wire new_Jinkela_wire_4252;
    wire new_Jinkela_wire_6628;
    wire new_Jinkela_wire_3267;
    wire new_Jinkela_wire_3255;
    wire new_Jinkela_wire_3083;
    wire new_Jinkela_wire_4455;
    wire new_Jinkela_wire_3411;
    wire _0338_;
    wire new_Jinkela_wire_3508;
    wire new_Jinkela_wire_7160;
    wire new_Jinkela_wire_7475;
    wire new_Jinkela_wire_4313;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_7258;
    wire _0492_;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_4550;
    wire new_Jinkela_wire_7139;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_5142;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_5287;
    wire _0933_;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_4863;
    wire new_Jinkela_wire_4755;
    wire new_Jinkela_wire_3850;
    wire new_Jinkela_wire_2638;
    wire new_Jinkela_wire_3450;
    wire new_Jinkela_wire_2567;
    wire _0863_;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_7440;
    wire _0205_;
    wire new_Jinkela_wire_3440;
    wire new_Jinkela_wire_2939;
    wire new_Jinkela_wire_7774;
    wire new_Jinkela_wire_5306;
    wire new_Jinkela_wire_6624;
    wire new_Jinkela_wire_2217;
    wire new_Jinkela_wire_1671;
    wire _0621_;
    wire new_Jinkela_wire_7922;
    wire new_Jinkela_wire_3953;
    wire new_Jinkela_wire_1907;
    wire _0079_;
    wire new_net_2509;
    wire new_Jinkela_wire_6837;
    wire new_Jinkela_wire_2574;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_6099;
    wire new_Jinkela_wire_5569;
    wire new_Jinkela_wire_5246;
    wire new_Jinkela_wire_7568;
    wire new_Jinkela_wire_7674;
    wire new_Jinkela_wire_718;
    wire _0704_;
    wire new_Jinkela_wire_6113;
    wire new_Jinkela_wire_2272;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_1788;
    wire new_Jinkela_wire_7506;
    wire new_Jinkela_wire_5286;
    wire _0097_;
    wire new_Jinkela_wire_6816;
    wire new_Jinkela_wire_3700;
    wire new_net_20;
    wire new_Jinkela_wire_3841;
    wire new_Jinkela_wire_2589;
    wire new_Jinkela_wire_7509;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_1284;
    wire new_Jinkela_wire_2244;
    wire new_Jinkela_wire_6016;
    wire new_net_2;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_3075;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_2828;
    wire new_Jinkela_wire_6108;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_2327;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_5428;
    wire new_Jinkela_wire_5644;
    wire new_Jinkela_wire_5857;
    wire new_Jinkela_wire_6205;
    wire new_Jinkela_wire_5805;
    wire new_Jinkela_wire_1721;
    wire new_Jinkela_wire_5917;
    wire new_Jinkela_wire_5173;
    wire new_Jinkela_wire_5541;
    wire new_Jinkela_wire_2909;
    wire new_Jinkela_wire_2940;
    wire new_Jinkela_wire_5885;
    wire new_Jinkela_wire_3266;
    wire new_Jinkela_wire_7824;
    wire new_Jinkela_wire_4371;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_2959;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_2373;
    wire new_Jinkela_wire_3280;
    wire new_Jinkela_wire_4399;
    wire new_Jinkela_wire_2408;
    wire new_Jinkela_wire_5924;
    wire new_Jinkela_wire_7742;
    wire new_Jinkela_wire_2258;
    wire new_Jinkela_wire_6899;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_1725;
    wire new_Jinkela_wire_4757;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_7659;
    wire new_Jinkela_wire_4633;
    wire new_Jinkela_wire_7651;
    wire new_Jinkela_wire_3455;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_8014;
    wire new_Jinkela_wire_3943;
    wire new_Jinkela_wire_2275;
    wire new_Jinkela_wire_7055;
    wire new_Jinkela_wire_4772;
    wire new_Jinkela_wire_6097;
    wire _0058_;
    wire _0247_;
    wire new_Jinkela_wire_2502;
    wire new_Jinkela_wire_6795;
    wire new_Jinkela_wire_3275;
    wire new_Jinkela_wire_2900;
    wire new_Jinkela_wire_2182;
    wire new_Jinkela_wire_7691;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_7300;
    wire new_Jinkela_wire_3715;
    wire new_Jinkela_wire_7588;
    wire _0055_;
    wire new_Jinkela_wire_3865;
    wire new_Jinkela_wire_7744;
    wire new_Jinkela_wire_1764;
    wire new_Jinkela_wire_7045;
    wire new_Jinkela_wire_4429;
    wire new_Jinkela_wire_3025;
    wire new_Jinkela_wire_4143;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_5149;
    wire new_Jinkela_wire_5171;
    wire new_Jinkela_wire_6674;
    wire new_Jinkela_wire_6283;
    wire new_Jinkela_wire_3240;
    wire new_Jinkela_wire_5726;
    wire new_Jinkela_wire_2402;
    wire new_Jinkela_wire_2974;
    wire new_Jinkela_wire_5448;
    wire new_Jinkela_wire_3942;
    wire new_Jinkela_wire_7816;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_4293;
    wire new_Jinkela_wire_5135;
    wire new_Jinkela_wire_6001;
    wire new_Jinkela_wire_5022;
    wire new_Jinkela_wire_6242;
    wire new_Jinkela_wire_4359;
    wire new_Jinkela_wire_5008;
    wire new_Jinkela_wire_2986;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_3977;
    wire new_Jinkela_wire_7459;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_4816;
    wire new_Jinkela_wire_2439;
    wire new_Jinkela_wire_2953;
    wire new_Jinkela_wire_2267;
    wire _0783_;
    wire new_Jinkela_wire_4804;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_3315;
    wire new_Jinkela_wire_6379;
    wire new_Jinkela_wire_3035;
    wire new_Jinkela_wire_5854;
    wire new_Jinkela_wire_3985;
    wire _0565_;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_7515;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_6796;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_6362;
    wire new_Jinkela_wire_3647;
    wire new_Jinkela_wire_6945;
    wire new_Jinkela_wire_3167;
    wire new_Jinkela_wire_5646;
    wire new_Jinkela_wire_7915;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_7645;
    wire new_Jinkela_wire_6439;
    wire new_Jinkela_wire_4765;
    wire new_Jinkela_wire_1715;
    wire new_Jinkela_wire_6893;
    wire new_Jinkela_wire_4972;
    wire new_Jinkela_wire_2104;
    wire new_Jinkela_wire_7677;
    wire new_Jinkela_wire_2118;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_6443;
    wire _0360_;
    wire new_Jinkela_wire_3855;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_5784;
    wire new_Jinkela_wire_2285;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_2560;
    wire new_Jinkela_wire_3612;
    wire new_Jinkela_wire_5025;
    wire new_Jinkela_wire_1967;
    wire new_Jinkela_wire_6706;
    wire new_Jinkela_wire_6415;
    wire new_Jinkela_wire_2274;
    wire new_Jinkela_wire_5974;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_7162;
    wire new_Jinkela_wire_5674;
    wire new_Jinkela_wire_7733;
    wire new_Jinkela_wire_3282;
    wire new_Jinkela_wire_3446;
    wire new_net_2483;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_4214;
    wire new_Jinkela_wire_3851;
    wire new_Jinkela_wire_5509;
    wire new_Jinkela_wire_5778;
    wire new_Jinkela_wire_7783;
    wire new_Jinkela_wire_4684;
    wire new_Jinkela_wire_2892;
    wire _0432_;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_6871;
    wire new_Jinkela_wire_1846;
    wire new_Jinkela_wire_7885;
    wire new_Jinkela_wire_3935;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_2999;
    wire _0692_;
    wire new_Jinkela_wire_3304;
    wire new_Jinkela_wire_4303;
    wire _0951_;
    wire _0899_;
    wire new_Jinkela_wire_7096;
    wire _0816_;
    wire new_Jinkela_wire_7070;
    wire new_Jinkela_wire_5452;
    wire _0701_;
    wire new_Jinkela_wire_5658;
    wire new_Jinkela_wire_40;
    wire new_net_22;
    wire new_Jinkela_wire_4342;
    wire new_Jinkela_wire_3536;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_6857;
    wire new_Jinkela_wire_2691;
    wire new_Jinkela_wire_3651;
    wire new_Jinkela_wire_6903;
    wire new_Jinkela_wire_7018;
    wire new_Jinkela_wire_5003;
    wire _0847_;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_4566;
    wire new_Jinkela_wire_5907;
    wire new_Jinkela_wire_1657;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_7099;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_3381;
    wire new_Jinkela_wire_5721;
    wire new_Jinkela_wire_4448;
    wire new_Jinkela_wire_3055;
    wire new_Jinkela_wire_2390;
    wire new_Jinkela_wire_3460;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_2133;
    wire _0682_;
    wire new_Jinkela_wire_4277;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_1726;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_7953;
    wire _1199_;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_5585;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_2753;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_4788;
    wire new_Jinkela_wire_3379;
    wire new_Jinkela_wire_2332;
    wire _0819_;
    wire new_Jinkela_wire_4079;
    wire new_Jinkela_wire_5237;
    wire new_Jinkela_wire_5683;
    wire new_Jinkela_wire_5434;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_4754;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_6941;
    wire _0267_;
    wire _0370_;
    wire new_Jinkela_wire_3878;
    wire new_Jinkela_wire_3822;
    wire new_Jinkela_wire_7351;
    wire new_Jinkela_wire_2003;
    wire new_Jinkela_wire_1575;
    wire _0094_;
    wire new_Jinkela_wire_7550;
    wire new_Jinkela_wire_2177;
    wire new_Jinkela_wire_3525;
    wire new_Jinkela_wire_7810;
    wire new_Jinkela_wire_6368;
    wire _0970_;
    wire new_Jinkela_wire_4606;
    wire _0181_;
    wire new_Jinkela_wire_3000;
    wire new_Jinkela_wire_3913;
    wire new_Jinkela_wire_7313;
    wire new_Jinkela_wire_2736;
    wire new_Jinkela_wire_3042;
    wire _1104_;
    wire new_Jinkela_wire_5754;
    wire _0971_;
    wire new_Jinkela_wire_6976;
    wire _0675_;
    wire new_Jinkela_wire_7750;
    wire _0568_;
    wire new_Jinkela_wire_3188;
    wire new_Jinkela_wire_2516;
    wire new_Jinkela_wire_7805;
    wire new_Jinkela_wire_5860;
    wire new_Jinkela_wire_7164;
    wire new_Jinkela_wire_4813;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_1269;
    wire _1227_;
    wire new_Jinkela_wire_7846;
    wire new_Jinkela_wire_6365;
    wire new_Jinkela_wire_6086;
    wire new_Jinkela_wire_5185;
    wire new_Jinkela_wire_3567;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_6014;
    wire new_Jinkela_wire_2564;
    wire new_Jinkela_wire_3294;
    wire new_Jinkela_wire_7144;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_4657;
    wire _0483_;
    wire new_Jinkela_wire_6134;
    wire new_Jinkela_wire_7950;
    wire new_Jinkela_wire_4877;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_3164;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_5054;
    wire new_Jinkela_wire_4039;
    wire new_Jinkela_wire_5590;
    wire new_Jinkela_wire_4965;
    wire new_Jinkela_wire_4693;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_5750;
    wire new_Jinkela_wire_3229;
    wire _0212_;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_5614;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_3242;
    wire new_Jinkela_wire_6687;
    wire new_Jinkela_wire_2521;
    wire new_Jinkela_wire_6533;
    wire new_Jinkela_wire_2456;
    wire new_Jinkela_wire_2181;
    wire new_Jinkela_wire_7520;
    wire _0357_;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_3774;
    wire _1092_;
    wire new_Jinkela_wire_4930;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_2315;
    wire new_Jinkela_wire_7656;
    wire new_Jinkela_wire_2366;
    wire new_Jinkela_wire_3767;
    wire new_Jinkela_wire_3699;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_2684;
    wire new_Jinkela_wire_3225;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_2595;
    wire _0551_;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_6427;
    wire new_Jinkela_wire_2158;
    wire new_Jinkela_wire_6536;
    wire new_Jinkela_wire_1997;
    wire new_Jinkela_wire_5094;
    wire new_net_23;
    wire new_Jinkela_wire_4021;
    wire _0386_;
    wire new_Jinkela_wire_6259;
    wire new_Jinkela_wire_2361;
    wire new_Jinkela_wire_5439;
    wire new_Jinkela_wire_6012;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_7127;
    wire new_Jinkela_wire_5190;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_6601;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_7635;
    wire new_Jinkela_wire_3760;
    wire new_Jinkela_wire_3847;
    wire _0327_;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_3752;
    wire new_Jinkela_wire_3863;
    wire new_Jinkela_wire_61;
    wire new_Jinkela_wire_2360;
    wire new_Jinkela_wire_5150;
    wire new_Jinkela_wire_2770;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_1675;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_5632;
    wire new_Jinkela_wire_7078;
    wire new_Jinkela_wire_2507;
    wire new_Jinkela_wire_2100;
    wire new_Jinkela_wire_7151;
    wire new_Jinkela_wire_4842;
    wire new_Jinkela_wire_6538;
    wire new_Jinkela_wire_4068;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_5038;
    wire new_Jinkela_wire_7034;
    wire new_Jinkela_wire_219;
    wire _0575_;
    wire new_Jinkela_wire_7696;
    wire new_Jinkela_wire_7059;
    wire new_Jinkela_wire_7711;
    wire new_Jinkela_wire_7601;
    wire _0100_;
    wire new_Jinkela_wire_6824;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_7290;
    wire new_Jinkela_wire_5292;
    wire new_Jinkela_wire_3874;
    wire new_Jinkela_wire_5748;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_7989;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_5507;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_7229;
    wire new_Jinkela_wire_6376;
    wire _0655_;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_5087;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_3400;
    wire new_Jinkela_wire_6786;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_6383;
    wire new_Jinkela_wire_1855;
    wire new_Jinkela_wire_5956;
    wire new_Jinkela_wire_2189;
    wire _1043_;
    wire new_Jinkela_wire_5531;
    wire _0044_;
    wire new_Jinkela_wire_2966;
    wire _1141_;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_4891;
    wire new_Jinkela_wire_3192;
    wire new_Jinkela_wire_4999;
    wire new_Jinkela_wire_4637;
    wire new_Jinkela_wire_196;
    wire _0625_;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_7864;
    wire new_Jinkela_wire_2910;
    wire new_Jinkela_wire_5253;
    wire _0902_;
    wire new_Jinkela_wire_2114;
    wire new_Jinkela_wire_3658;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_3032;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_5602;
    wire new_Jinkela_wire_4074;
    wire _0148_;
    wire new_Jinkela_wire_1856;
    wire _0880_;
    wire new_Jinkela_wire_3716;
    wire new_Jinkela_wire_25;
    wire _0821_;
    wire new_Jinkela_wire_2300;
    wire new_Jinkela_wire_2462;
    wire new_Jinkela_wire_4009;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_4705;
    wire new_Jinkela_wire_5891;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_1741;
    wire new_Jinkela_wire_2397;
    wire new_Jinkela_wire_3765;
    wire _0795_;
    wire new_Jinkela_wire_4522;
    wire new_Jinkela_wire_6378;
    wire new_Jinkela_wire_4660;
    wire new_Jinkela_wire_2259;
    wire _0388_;
    wire _0237_;
    wire new_Jinkela_wire_493;
    wire _0470_;
    wire _1234_;
    wire new_Jinkela_wire_2879;
    wire new_Jinkela_wire_3263;
    wire new_Jinkela_wire_6307;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_477;
    wire _0965_;
    wire new_Jinkela_wire_6143;
    wire new_Jinkela_wire_4488;
    wire new_Jinkela_wire_2447;
    wire new_Jinkela_wire_4087;
    wire new_Jinkela_wire_5539;
    wire new_Jinkela_wire_7277;
    wire new_Jinkela_wire_4901;
    wire new_Jinkela_wire_3503;
    wire new_Jinkela_wire_1859;
    wire new_Jinkela_wire_6668;
    wire new_Jinkela_wire_2876;
    wire new_Jinkela_wire_5387;
    wire new_Jinkela_wire_7264;
    wire new_Jinkela_wire_2233;
    wire new_Jinkela_wire_7752;
    wire new_Jinkela_wire_7273;
    wire new_Jinkela_wire_2122;
    wire new_Jinkela_wire_3980;
    wire new_Jinkela_wire_7377;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_5609;
    wire new_Jinkela_wire_5473;
    wire new_Jinkela_wire_1993;
    wire new_Jinkela_wire_256;
    wire _0638_;
    wire _0286_;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_5264;
    wire new_Jinkela_wire_7314;
    wire new_Jinkela_wire_3061;
    wire new_Jinkela_wire_5637;
    wire new_net_2499;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_4590;
    wire new_Jinkela_wire_4748;
    wire new_net_2439;
    wire new_Jinkela_wire_4169;
    wire new_Jinkela_wire_7485;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_3988;
    wire new_Jinkela_wire_4865;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_5;
    wire _0735_;
    wire _0681_;
    wire new_Jinkela_wire_2037;
    wire _0403_;
    wire new_Jinkela_wire_7406;
    wire new_Jinkela_wire_5994;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_2943;
    wire new_Jinkela_wire_6693;
    wire new_Jinkela_wire_3048;
    wire new_Jinkela_wire_3680;
    wire new_Jinkela_wire_6112;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_7311;
    wire new_Jinkela_wire_7426;
    wire new_Jinkela_wire_3136;
    wire new_Jinkela_wire_6930;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_5040;
    wire new_Jinkela_wire_3764;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_5524;
    wire new_Jinkela_wire_7462;
    wire new_Jinkela_wire_4463;
    wire new_Jinkela_wire_2219;
    wire _0975_;
    wire new_Jinkela_wire_5978;
    wire new_Jinkela_wire_5051;
    wire new_Jinkela_wire_6633;
    wire _0872_;
    wire new_Jinkela_wire_3438;
    wire new_Jinkela_wire_7184;
    wire new_Jinkela_wire_4544;
    wire new_Jinkela_wire_7773;
    wire new_Jinkela_wire_7724;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_3081;
    wire new_Jinkela_wire_7729;
    wire _0249_;
    wire new_Jinkela_wire_2171;
    wire new_Jinkela_wire_5736;
    wire new_Jinkela_wire_7803;
    wire new_Jinkela_wire_7907;
    wire new_Jinkela_wire_4686;
    wire _0424_;
    wire new_Jinkela_wire_7381;
    wire new_Jinkela_wire_2046;
    wire new_Jinkela_wire_5154;
    wire new_Jinkela_wire_7842;
    wire new_Jinkela_wire_104;
    wire _0768_;
    wire new_Jinkela_wire_7470;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_7116;
    wire new_Jinkela_wire_2413;
    wire new_Jinkela_wire_7432;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_4357;
    wire _0196_;
    wire new_Jinkela_wire_2927;
    wire new_Jinkela_wire_1775;
    wire _1067_;
    wire new_Jinkela_wire_6266;
    wire new_Jinkela_wire_6942;
    wire new_Jinkela_wire_2358;
    wire new_Jinkela_wire_3792;
    wire _0272_;
    wire _1110_;
    wire new_Jinkela_wire_6297;
    wire new_Jinkela_wire_7080;
    wire new_net_2355;
    wire new_Jinkela_wire_981;
    wire new_Jinkela_wire_5379;
    wire new_Jinkela_wire_6204;
    wire new_Jinkela_wire_2205;
    wire new_Jinkela_wire_1881;
    wire new_Jinkela_wire_1720;
    wire new_Jinkela_wire_1145;
    wire new_Jinkela_wire_4027;
    wire _0519_;
    wire new_Jinkela_wire_598;
    wire _0906_;
    wire new_Jinkela_wire_3859;
    wire _0961_;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_2731;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_4518;
    wire new_Jinkela_wire_6104;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_6960;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_4119;
    wire _0552_;
    wire new_Jinkela_wire_5563;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_2888;
    wire new_Jinkela_wire_4738;
    wire new_Jinkela_wire_7252;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_4059;
    wire new_Jinkela_wire_1672;
    wire new_Jinkela_wire_2257;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_1803;
    wire new_Jinkela_wire_5236;
    wire _0689_;
    wire new_Jinkela_wire_7687;
    wire new_Jinkela_wire_3835;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_7046;
    wire new_Jinkela_wire_4375;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_5663;
    wire _0111_;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_7665;
    wire new_Jinkela_wire_3456;
    wire new_Jinkela_wire_2947;
    wire new_Jinkela_wire_4197;
    wire new_Jinkela_wire_2868;
    wire new_Jinkela_wire_1929;
    wire new_Jinkela_wire_2659;
    wire new_Jinkela_wire_3197;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_2352;
    wire new_Jinkela_wire_4469;
    wire new_Jinkela_wire_6631;
    wire new_Jinkela_wire_3453;
    wire new_Jinkela_wire_2044;
    wire new_Jinkela_wire_4950;
    wire new_Jinkela_wire_3991;
    wire new_Jinkela_wire_5144;
    wire new_Jinkela_wire_2651;
    wire new_Jinkela_wire_7787;
    wire new_Jinkela_wire_2028;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_5901;
    wire new_Jinkela_wire_2975;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_4927;
    wire _1082_;
    wire _0155_;
    wire new_Jinkela_wire_6833;
    wire new_Jinkela_wire_6319;
    wire new_Jinkela_wire_6211;
    wire _0389_;
    wire new_Jinkela_wire_3926;
    wire new_Jinkela_wire_7323;
    wire new_Jinkela_wire_5871;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_7085;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_7522;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_4495;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_5303;
    wire new_Jinkela_wire_3734;
    wire new_Jinkela_wire_5545;
    wire new_Jinkela_wire_2355;
    wire new_Jinkela_wire_6615;
    wire new_Jinkela_wire_7855;
    wire new_Jinkela_wire_5573;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_6168;
    wire new_Jinkela_wire_2549;
    wire new_Jinkela_wire_6678;
    wire _1241_;
    wire new_Jinkela_wire_7174;
    wire new_Jinkela_wire_7140;
    wire new_Jinkela_wire_4441;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_5367;
    wire new_Jinkela_wire_2265;
    wire new_Jinkela_wire_5454;
    wire new_Jinkela_wire_5645;
    wire new_Jinkela_wire_5244;
    wire new_Jinkela_wire_6270;
    wire _1232_;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_4213;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_2453;
    wire new_Jinkela_wire_4182;
    wire new_Jinkela_wire_2196;
    wire new_Jinkela_wire_5227;
    wire _0463_;
    wire new_Jinkela_wire_2922;
    wire new_Jinkela_wire_6578;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_5800;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_3713;
    wire new_Jinkela_wire_4979;
    wire new_Jinkela_wire_5742;
    wire new_Jinkela_wire_6864;
    wire new_Jinkela_wire_6385;
    wire _1090_;
    wire new_Jinkela_wire_4784;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_6239;
    wire new_Jinkela_wire_7492;
    wire _0956_;
    wire new_Jinkela_wire_7291;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_5396;
    wire _0248_;
    wire new_Jinkela_wire_7852;
    wire new_Jinkela_wire_5841;
    wire _0303_;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_4285;
    wire new_Jinkela_wire_7255;
    wire new_Jinkela_wire_6100;
    wire _0640_;
    wire new_Jinkela_wire_2140;
    wire new_Jinkela_wire_4478;
    wire new_Jinkela_wire_3273;
    wire new_Jinkela_wire_5990;
    wire new_Jinkela_wire_5818;
    wire new_Jinkela_wire_3703;
    wire _1128_;
    wire new_Jinkela_wire_2696;
    wire new_Jinkela_wire_3208;
    wire _0342_;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_4349;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_4549;
    wire _0992_;
    wire new_Jinkela_wire_4155;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_3115;
    wire new_Jinkela_wire_2542;
    wire new_Jinkela_wire_6085;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_2214;
    wire new_Jinkela_wire_4640;
    wire new_Jinkela_wire_7447;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_2565;
    wire new_Jinkela_wire_3572;
    wire new_Jinkela_wire_6216;
    wire new_Jinkela_wire_3396;
    wire new_Jinkela_wire_5321;
    wire new_Jinkela_wire_7053;
    wire new_Jinkela_wire_6268;
    wire new_Jinkela_wire_6151;
    wire new_Jinkela_wire_4189;
    wire new_Jinkela_wire_3910;
    wire new_Jinkela_wire_3132;
    wire new_Jinkela_wire_4822;
    wire new_Jinkela_wire_5482;
    wire new_Jinkela_wire_1854;
    wire new_Jinkela_wire_2728;
    wire new_Jinkela_wire_2175;
    wire new_Jinkela_wire_2658;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_3990;
    wire new_Jinkela_wire_4596;
    wire new_Jinkela_wire_6562;
    wire _0703_;
    wire new_Jinkela_wire_3893;
    wire new_Jinkela_wire_1166;
    wire _1018_;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_6521;
    wire new_Jinkela_wire_5780;
    wire new_Jinkela_wire_7919;
    wire new_Jinkela_wire_7967;
    wire new_net_2455;
    wire new_Jinkela_wire_2964;
    wire new_Jinkela_wire_5146;
    wire new_Jinkela_wire_5114;
    wire new_Jinkela_wire_6178;
    wire new_Jinkela_wire_5156;
    wire new_Jinkela_wire_4203;
    wire new_Jinkela_wire_5198;
    wire new_Jinkela_wire_4747;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_5019;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_6922;
    wire _0364_;
    wire new_Jinkela_wire_6274;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_4045;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_7924;
    wire new_Jinkela_wire_2243;
    wire new_Jinkela_wire_4654;
    wire new_Jinkela_wire_2025;
    wire _0006_;
    wire new_Jinkela_wire_4581;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_6013;
    wire new_Jinkela_wire_1861;
    wire _0371_;
    wire new_Jinkela_wire_4750;
    wire new_Jinkela_wire_6179;
    wire new_Jinkela_wire_7939;
    wire new_Jinkela_wire_6971;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_6634;
    wire new_Jinkela_wire_7640;
    wire new_Jinkela_wire_3277;
    wire new_Jinkela_wire_3120;
    wire new_Jinkela_wire_7917;
    wire new_Jinkela_wire_3827;
    wire _0003_;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_430;
    wire _0349_;
    wire new_Jinkela_wire_3013;
    wire new_Jinkela_wire_3966;
    wire new_Jinkela_wire_6147;
    wire new_Jinkela_wire_4124;
    wire new_net_10;
    wire new_Jinkela_wire_4057;
    wire new_Jinkela_wire_2936;
    wire _0172_;
    wire new_Jinkela_wire_7668;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_3597;
    wire new_Jinkela_wire_3924;
    wire new_Jinkela_wire_4178;
    wire new_Jinkela_wire_4648;
    wire new_Jinkela_wire_6771;
    wire new_Jinkela_wire_7706;
    wire new_Jinkela_wire_4367;
    wire new_net_2351;
    wire _0978_;
    wire new_Jinkela_wire_5036;
    wire new_Jinkela_wire_4259;
    wire new_Jinkela_wire_7765;
    wire _0356_;
    wire _0202_;
    wire new_Jinkela_wire_5935;
    wire new_Jinkela_wire_6496;
    wire new_Jinkela_wire_6769;
    wire new_Jinkela_wire_7793;
    wire new_Jinkela_wire_3537;
    wire new_Jinkela_wire_7698;
    wire _0908_;
    wire new_Jinkela_wire_5260;
    wire new_Jinkela_wire_6670;
    wire new_Jinkela_wire_5165;
    wire new_Jinkela_wire_6084;
    wire new_Jinkela_wire_730;
    wire _0801_;
    wire new_Jinkela_wire_2298;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_2261;
    wire new_Jinkela_wire_3530;
    wire new_Jinkela_wire_6493;
    wire new_Jinkela_wire_6812;
    wire new_Jinkela_wire_1977;
    wire new_net_2367;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_1809;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_2295;
    wire new_Jinkela_wire_7753;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_6063;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_2528;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_4083;
    wire new_Jinkela_wire_6037;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_3870;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_6095;
    wire new_Jinkela_wire_7642;
    wire _0535_;
    wire new_Jinkela_wire_7624;
    wire new_Jinkela_wire_3087;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_7357;
    wire _0890_;
    wire new_Jinkela_wire_4272;
    wire new_Jinkela_wire_3364;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_2647;
    wire _0257_;
    wire new_Jinkela_wire_5523;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_6102;
    wire new_Jinkela_wire_6021;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_6949;
    wire new_Jinkela_wire_2822;
    wire new_Jinkela_wire_7973;
    wire new_Jinkela_wire_2682;
    wire new_Jinkela_wire_6996;
    wire new_Jinkela_wire_6610;
    wire new_Jinkela_wire_7587;
    wire new_Jinkela_wire_2926;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_6246;
    wire new_Jinkela_wire_4760;
    wire new_Jinkela_wire_6673;
    wire new_Jinkela_wire_7777;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_118;
    wire _0841_;
    wire _0917_;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_6420;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_2445;
    wire new_Jinkela_wire_2086;
    wire new_Jinkela_wire_2819;
    wire new_Jinkela_wire_1110;
    wire _1102_;
    wire new_Jinkela_wire_6965;
    wire new_Jinkela_wire_7845;
    wire new_Jinkela_wire_4439;
    wire new_Jinkela_wire_298;
    wire _0080_;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_6863;
    wire new_Jinkela_wire_1820;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_5130;
    wire new_Jinkela_wire_1279;
    wire _0164_;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_7147;
    wire new_Jinkela_wire_109;
    wire _0048_;
    wire new_Jinkela_wire_6831;
    wire new_Jinkela_wire_7380;
    wire new_Jinkela_wire_6027;
    wire _0326_;
    wire new_Jinkela_wire_3007;
    wire _0222_;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_7216;
    wire new_Jinkela_wire_7225;
    wire new_Jinkela_wire_3040;
    wire new_Jinkela_wire_42;
    wire new_net_12;
    wire new_Jinkela_wire_4588;
    wire new_Jinkela_wire_6984;
    wire new_Jinkela_wire_4333;
    wire new_Jinkela_wire_2268;
    wire _0454_;
    wire new_Jinkela_wire_6884;
    wire new_Jinkela_wire_5839;
    wire new_Jinkela_wire_3409;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_7145;
    wire new_Jinkela_wire_7050;
    wire new_Jinkela_wire_3492;
    wire new_Jinkela_wire_6840;
    wire new_Jinkela_wire_4781;
    wire new_Jinkela_wire_3085;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_4977;
    wire new_Jinkela_wire_6456;
    wire _0332_;
    wire _0680_;
    wire new_Jinkela_wire_2087;
    wire new_Jinkela_wire_5389;
    wire new_Jinkela_wire_1483;
    wire _0709_;
    wire new_Jinkela_wire_5759;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_2374;
    wire new_Jinkela_wire_6347;
    wire new_Jinkela_wire_6154;
    wire new_Jinkela_wire_4296;
    wire new_Jinkela_wire_5505;
    wire new_Jinkela_wire_4896;
    wire new_Jinkela_wire_4427;
    wire new_Jinkela_wire_1916;
    wire new_Jinkela_wire_5629;
    wire new_Jinkela_wire_2188;
    wire new_Jinkela_wire_7517;
    wire _0264_;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_5463;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_6635;
    wire new_Jinkela_wire_4467;
    wire _0858_;
    wire new_net_2405;
    wire new_Jinkela_wire_3320;
    wire new_Jinkela_wire_7374;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_2049;
    wire new_Jinkela_wire_3403;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_7772;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_3606;
    wire _0362_;
    wire _0397_;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_3279;
    wire _0921_;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_4046;
    wire new_Jinkela_wire_5802;
    wire _1038_;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_7508;
    wire new_Jinkela_wire_2559;
    wire new_Jinkela_wire_6039;
    wire new_Jinkela_wire_2483;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_1740;
    wire new_Jinkela_wire_3585;
    wire new_Jinkela_wire_4351;
    wire new_Jinkela_wire_4343;
    wire new_Jinkela_wire_5419;
    wire _0796_;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_7565;
    wire _0952_;
    wire new_Jinkela_wire_7821;
    wire new_Jinkela_wire_4466;
    wire new_Jinkela_wire_3524;
    wire new_Jinkela_wire_6403;
    wire new_Jinkela_wire_7463;
    wire new_Jinkela_wire_7619;
    wire new_Jinkela_wire_5850;
    wire new_Jinkela_wire_4205;
    wire new_Jinkela_wire_7945;
    wire new_Jinkela_wire_7281;
    wire new_Jinkela_wire_5878;
    wire new_Jinkela_wire_3547;
    wire _0476_;
    wire new_Jinkela_wire_2845;
    wire new_Jinkela_wire_8003;
    wire new_Jinkela_wire_7748;
    wire new_Jinkela_wire_795;
    wire _0932_;
    wire new_Jinkela_wire_5480;
    wire _0944_;
    wire new_Jinkela_wire_6745;
    wire new_Jinkela_wire_3787;
    wire new_Jinkela_wire_2089;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_5195;
    wire new_Jinkela_wire_5991;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_5813;
    wire new_Jinkela_wire_1141;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_5283;
    wire new_Jinkela_wire_3039;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_5219;
    wire new_Jinkela_wire_6868;
    wire new_Jinkela_wire_7238;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_2555;
    wire new_Jinkela_wire_4952;
    wire new_Jinkela_wire_6509;
    wire _0198_;
    wire new_Jinkela_wire_6718;
    wire new_Jinkela_wire_6800;
    wire new_Jinkela_wire_4225;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_6124;
    wire _0071_;
    wire new_Jinkela_wire_2293;
    wire new_Jinkela_wire_2875;
    wire new_Jinkela_wire_5372;
    wire new_Jinkela_wire_4811;
    wire new_Jinkela_wire_5792;
    wire new_Jinkela_wire_1599;
    wire _0074_;
    wire new_Jinkela_wire_3036;
    wire new_Jinkela_wire_5075;
    wire new_Jinkela_wire_6399;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_3401;
    wire new_Jinkela_wire_3584;
    wire new_Jinkela_wire_2877;
    wire new_Jinkela_wire_6978;
    wire new_Jinkela_wire_1969;
    wire _0501_;
    wire _1134_;
    wire new_Jinkela_wire_5212;
    wire new_Jinkela_wire_4382;
    wire new_Jinkela_wire_913;
    wire _0531_;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_6808;
    wire new_Jinkela_wire_6222;
    wire _0162_;
    wire new_Jinkela_wire_4728;
    wire new_Jinkela_wire_4424;
    wire new_Jinkela_wire_7940;
    wire new_Jinkela_wire_6289;
    wire new_Jinkela_wire_7853;
    wire new_Jinkela_wire_3062;
    wire new_Jinkela_wire_2407;
    wire new_Jinkela_wire_6880;
    wire new_Jinkela_wire_2776;
    wire new_Jinkela_wire_2538;
    wire new_Jinkela_wire_2410;
    wire _0302_;
    wire new_Jinkela_wire_7860;
    wire new_Jinkela_wire_4134;
    wire new_net_24;
    wire new_Jinkela_wire_2830;
    wire new_net_2425;
    wire new_Jinkela_wire_6970;
    wire new_Jinkela_wire_4942;
    wire new_Jinkela_wire_4176;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_6608;
    wire _1247_;
    wire new_Jinkela_wire_6341;
    wire new_Jinkela_wire_3947;
    wire _0942_;
    wire new_Jinkela_wire_3260;
    wire new_Jinkela_wire_7878;
    wire _1224_;
    wire new_Jinkela_wire_3398;
    wire _0810_;
    wire new_Jinkela_wire_3829;
    wire new_Jinkela_wire_2180;
    wire new_Jinkela_wire_7995;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_7482;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_2215;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_2250;
    wire new_Jinkela_wire_3684;
    wire new_Jinkela_wire_6116;
    wire new_Jinkela_wire_5504;
    wire new_Jinkela_wire_2377;
    wire new_Jinkela_wire_2540;
    wire new_Jinkela_wire_3198;
    wire _1046_;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_7567;
    wire new_Jinkela_wire_56;
    wire new_Jinkela_wire_5572;
    wire _1211_;
    wire new_Jinkela_wire_7523;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_2924;
    wire new_Jinkela_wire_7730;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_5790;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_4910;
    wire new_Jinkela_wire_5992;
    wire new_Jinkela_wire_2960;
    wire new_Jinkela_wire_5979;
    wire _0578_;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_4676;
    wire new_Jinkela_wire_6862;
    wire new_Jinkela_wire_3334;
    wire new_Jinkela_wire_6150;
    wire new_Jinkela_wire_6072;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_6398;
    wire new_Jinkela_wire_1266;
    wire new_Jinkela_wire_3281;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_1687;
    wire new_Jinkela_wire_3618;
    wire new_Jinkela_wire_1895;
    wire new_Jinkela_wire_2633;
    wire new_Jinkela_wire_7761;
    wire new_Jinkela_wire_3918;
    wire new_Jinkela_wire_2621;
    wire new_Jinkela_wire_7029;
    wire new_Jinkela_wire_4251;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_3948;
    wire new_Jinkela_wire_2273;
    wire new_Jinkela_wire_6285;
    wire new_Jinkela_wire_2338;
    wire _0605_;
    wire new_Jinkela_wire_5443;
    wire new_Jinkela_wire_5783;
    wire new_Jinkela_wire_6898;
    wire new_Jinkela_wire_4328;
    wire _0305_;
    wire new_Jinkela_wire_6333;
    wire new_Jinkela_wire_4922;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_1404;
    wire new_Jinkela_wire_5706;
    wire new_Jinkela_wire_701;
    wire _0660_;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_4546;
    wire new_Jinkela_wire_2012;
    wire new_Jinkela_wire_6717;
    wire new_Jinkela_wire_2136;
    wire new_Jinkela_wire_5929;
    wire new_Jinkela_wire_3644;
    wire new_Jinkela_wire_7830;
    wire new_Jinkela_wire_7970;
    wire new_Jinkela_wire_6203;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_3779;
    wire new_Jinkela_wire_6878;
    wire new_Jinkela_wire_6544;
    wire new_Jinkela_wire_4962;
    wire new_Jinkela_wire_1889;
    wire new_Jinkela_wire_7495;
    wire new_Jinkela_wire_4975;
    wire new_Jinkela_wire_6132;
    wire new_Jinkela_wire_7201;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_5137;
    wire new_Jinkela_wire_3424;
    wire new_Jinkela_wire_560;
    wire _0784_;
    wire new_Jinkela_wire_1806;
    wire new_Jinkela_wire_6105;
    wire new_Jinkela_wire_2760;
    wire new_Jinkela_wire_4344;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_2858;
    wire new_Jinkela_wire_3024;
    wire _0246_;
    wire new_Jinkela_wire_2546;
    wire _0691_;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_4528;
    wire _0124_;
    wire new_Jinkela_wire_4141;
    wire _0135_;
    wire new_Jinkela_wire_3233;
    wire _0337_;
    wire new_Jinkela_wire_5476;
    wire new_Jinkela_wire_3419;
    wire new_Jinkela_wire_7557;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_4387;
    wire _0391_;
    wire new_Jinkela_wire_5228;
    wire new_Jinkela_wire_2655;
    wire new_Jinkela_wire_6357;
    wire new_Jinkela_wire_3022;
    wire new_Jinkela_wire_7065;
    wire new_Jinkela_wire_6939;
    wire new_Jinkela_wire_5382;
    wire new_Jinkela_wire_7992;
    wire new_Jinkela_wire_3616;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_4065;
    wire new_Jinkela_wire_7219;
    wire new_Jinkela_wire_2786;
    wire new_Jinkela_wire_6494;
    wire new_Jinkela_wire_1245;
    wire new_Jinkela_wire_6653;
    wire new_Jinkela_wire_190;
    wire _0928_;
    wire new_Jinkela_wire_6581;
    wire _0851_;
    wire _1087_;
    wire new_Jinkela_wire_6664;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_6571;
    wire _0175_;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_6551;
    wire new_Jinkela_wire_5985;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_1591;
    wire new_Jinkela_wire_5072;
    wire new_Jinkela_wire_423;
    wire _0914_;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_5756;
    wire new_Jinkela_wire_7289;
    wire new_Jinkela_wire_2816;
    wire new_Jinkela_wire_2497;
    wire new_Jinkela_wire_4532;
    wire new_Jinkela_wire_4044;
    wire new_Jinkela_wire_365;
    wire _0373_;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_8004;
    wire new_net_2485;
    wire new_Jinkela_wire_4404;
    wire new_Jinkela_wire_6327;
    wire new_Jinkela_wire_6566;
    wire new_Jinkela_wire_4007;
    wire new_net_13;
    wire new_Jinkela_wire_2937;
    wire new_Jinkela_wire_2137;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_6471;
    wire new_Jinkela_wire_6993;
    wire new_Jinkela_wire_4015;
    wire new_Jinkela_wire_4572;
    wire new_Jinkela_wire_5206;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_5771;
    wire new_Jinkela_wire_4745;
    wire new_Jinkela_wire_2379;
    wire new_Jinkela_wire_5596;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_7518;
    wire new_Jinkela_wire_7199;
    wire _0304_;
    wire _0009_;
    wire new_Jinkela_wire_2673;
    wire new_Jinkela_wire_7152;
    wire new_Jinkela_wire_3490;
    wire new_Jinkela_wire_3126;
    wire new_Jinkela_wire_5213;
    wire new_Jinkela_wire_3772;
    wire _1012_;
    wire new_Jinkela_wire_6114;
    wire new_Jinkela_wire_6525;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_2572;
    wire new_Jinkela_wire_4329;
    wire new_Jinkela_wire_6355;
    wire new_Jinkela_wire_6017;
    wire new_Jinkela_wire_1262;
    wire new_Jinkela_wire_5461;
    wire new_Jinkela_wire_2423;
    wire new_Jinkela_wire_7008;
    wire new_Jinkela_wire_1612;
    wire new_Jinkela_wire_835;
    wire new_Jinkela_wire_3830;
    wire new_Jinkela_wire_1373;
    wire new_net_1;
    wire new_Jinkela_wire_7190;
    wire new_Jinkela_wire_6908;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_7389;
    wire new_Jinkela_wire_6890;
    wire new_Jinkela_wire_7307;
    wire new_Jinkela_wire_3588;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_3412;
    wire new_Jinkela_wire_2321;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_2604;
    wire _1109_;
    wire new_Jinkela_wire_7009;
    wire new_Jinkela_wire_1947;
    wire new_Jinkela_wire_4763;
    wire new_Jinkela_wire_5407;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_7337;
    wire new_Jinkela_wire_2899;
    wire _1129_;
    wire new_Jinkela_wire_4260;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_6282;
    wire _0782_;
    wire new_Jinkela_wire_3265;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_2403;
    wire new_Jinkela_wire_4254;
    wire new_Jinkela_wire_6019;
    wire new_Jinkela_wire_6597;
    wire new_Jinkela_wire_1829;
    wire new_Jinkela_wire_272;
    wire _0130_;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_4374;
    wire new_Jinkela_wire_3944;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_3176;
    wire new_Jinkela_wire_3634;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_6550;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_5882;
    wire _0696_;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_2353;
    wire new_Jinkela_wire_4629;
    wire new_Jinkela_wire_4306;
    wire new_Jinkela_wire_7909;
    wire new_Jinkela_wire_4836;
    wire new_Jinkela_wire_3028;
    wire new_Jinkela_wire_2350;
    wire new_Jinkela_wire_2411;
    wire new_Jinkela_wire_2239;
    wire new_Jinkela_wire_5369;
    wire new_Jinkela_wire_5453;
    wire new_Jinkela_wire_2079;
    wire _0834_;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_646;
    wire _0366_;
    wire new_Jinkela_wire_2917;
    wire new_Jinkela_wire_3896;
    wire new_Jinkela_wire_6989;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_4988;
    wire new_Jinkela_wire_4018;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_3604;
    wire new_Jinkela_wire_7204;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_5532;
    wire new_Jinkela_wire_3462;
    wire new_Jinkela_wire_4121;
    wire new_Jinkela_wire_2190;
    wire new_Jinkela_wire_7994;
    wire new_Jinkela_wire_5323;
    wire _0758_;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_6921;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_5465;
    wire new_Jinkela_wire_2569;
    wire new_Jinkela_wire_372;
    wire _0265_;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_6281;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_7450;
    wire new_Jinkela_wire_6688;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_7319;
    wire new_Jinkela_wire_2418;
    wire new_Jinkela_wire_7607;
    wire _1124_;
    wire new_Jinkela_wire_2982;
    wire new_Jinkela_wire_3949;
    wire new_Jinkela_wire_4240;
    wire new_Jinkela_wire_4069;
    wire new_Jinkela_wire_6643;
    wire new_Jinkela_wire_8021;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_1774;
    wire new_Jinkela_wire_7585;
    wire new_Jinkela_wire_2972;
    wire new_Jinkela_wire_4339;
    wire _0062_;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_5896;
    wire new_Jinkela_wire_2126;
    wire _1119_;
    wire new_Jinkela_wire_2735;
    wire _1004_;
    wire new_Jinkela_wire_1915;
    wire _0473_;
    wire new_Jinkela_wire_5272;
    wire new_Jinkela_wire_3672;
    wire new_Jinkela_wire_3184;
    wire new_Jinkela_wire_2065;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_3654;
    wire new_Jinkela_wire_7404;
    wire new_Jinkela_wire_5755;
    wire new_Jinkela_wire_2544;
    wire new_Jinkela_wire_1358;
    wire new_Jinkela_wire_3974;
    wire _0126_;
    wire new_Jinkela_wire_6557;
    wire new_Jinkela_wire_6082;
    wire new_Jinkela_wire_1991;
    wire new_Jinkela_wire_2931;
    wire new_Jinkela_wire_3377;
    wire new_Jinkela_wire_6326;
    wire new_Jinkela_wire_4806;
    wire new_Jinkela_wire_7546;
    wire new_Jinkela_wire_4534;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_5066;
    wire new_Jinkela_wire_7422;
    wire _0413_;
    wire new_Jinkela_wire_1140;
    wire _0415_;
    wire new_Jinkela_wire_2185;
    wire new_Jinkela_wire_3519;
    wire new_Jinkela_wire_3161;
    wire new_Jinkela_wire_6886;
    wire new_Jinkela_wire_6972;
    wire new_Jinkela_wire_4586;
    wire new_Jinkela_wire_7960;
    wire new_Jinkela_wire_6388;
    wire new_Jinkela_wire_7297;
    wire new_net_2369;
    wire new_Jinkela_wire_5656;
    wire new_Jinkela_wire_2650;
    wire new_Jinkela_wire_4783;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_5804;
    wire new_Jinkela_wire_3560;
    wire new_Jinkela_wire_5836;
    wire new_Jinkela_wire_7594;
    wire new_Jinkela_wire_4373;
    wire _0891_;
    wire new_Jinkela_wire_3413;
    wire new_Jinkela_wire_3052;
    wire new_Jinkela_wire_3956;
    wire new_Jinkela_wire_2351;
    wire new_Jinkela_wire_1759;
    wire new_Jinkela_wire_4620;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_7118;
    wire _0268_;
    wire new_Jinkela_wire_4000;
    wire _1034_;
    wire new_Jinkela_wire_3794;
    wire _0333_;
    wire new_Jinkela_wire_3871;
    wire new_Jinkela_wire_5069;
    wire new_Jinkela_wire_3220;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_3531;
    wire new_Jinkela_wire_7260;
    wire new_Jinkela_wire_3079;
    wire new_Jinkela_wire_7770;
    wire _1111_;
    wire new_Jinkela_wire_1073;
    wire new_Jinkela_wire_7605;
    wire _1069_;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_1500;
    wire _0762_;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_7887;
    wire new_Jinkela_wire_1702;
    wire _0283_;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_6860;
    wire new_Jinkela_wire_4100;
    wire new_Jinkela_wire_4682;
    wire new_Jinkela_wire_5047;
    wire new_Jinkela_wire_2833;
    wire new_Jinkela_wire_3165;
    wire new_Jinkela_wire_7978;
    wire new_Jinkela_wire_5701;
    wire new_Jinkela_wire_5359;
    wire new_Jinkela_wire_3168;
    wire new_Jinkela_wire_3528;
    wire new_Jinkela_wire_6990;
    wire new_Jinkela_wire_2721;
    wire new_Jinkela_wire_5035;
    wire new_Jinkela_wire_7429;
    wire _0666_;
    wire new_Jinkela_wire_7708;
    wire new_Jinkela_wire_5996;
    wire _0188_;
    wire new_Jinkela_wire_1739;
    wire new_Jinkela_wire_6582;
    wire new_Jinkela_wire_6731;
    wire new_Jinkela_wire_2349;
    wire new_Jinkela_wire_4133;
    wire _0813_;
    wire new_Jinkela_wire_7693;
    wire new_Jinkela_wire_7427;
    wire new_Jinkela_wire_2384;
    wire _1156_;
    wire new_Jinkela_wire_5344;
    wire new_Jinkela_wire_1126;
    wire _0594_;
    wire new_Jinkela_wire_2606;
    wire new_Jinkela_wire_4218;
    wire new_Jinkela_wire_5410;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_4497;
    wire new_Jinkela_wire_2054;
    wire new_Jinkela_wire_6914;
    wire _1246_;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_3037;
    wire _0794_;
    wire new_Jinkela_wire_3018;
    wire _0091_;
    wire new_Jinkela_wire_2740;
    wire _0767_;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_2626;
    wire _0204_;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_6232;
    wire _1080_;
    wire new_Jinkela_wire_2863;
    wire new_Jinkela_wire_7120;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_3602;
    wire new_Jinkela_wire_4593;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_6455;
    wire new_Jinkela_wire_3691;
    wire new_Jinkela_wire_6330;
    wire _0010_;
    wire new_net_9;
    wire new_Jinkela_wire_2015;
    wire new_Jinkela_wire_4859;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_4487;
    wire new_Jinkela_wire_3426;
    wire new_Jinkela_wire_5021;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_3965;
    wire new_Jinkela_wire_6952;
    wire new_Jinkela_wire_4023;
    wire new_Jinkela_wire_5888;
    wire new_Jinkela_wire_3627;
    wire new_Jinkela_wire_5949;
    wire new_Jinkela_wire_4542;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_5296;
    wire new_Jinkela_wire_5437;
    wire new_Jinkela_wire_7361;
    wire new_Jinkela_wire_1872;
    wire new_Jinkela_wire_3246;
    wire _1155_;
    wire new_Jinkela_wire_2481;
    wire _0427_;
    wire _0378_;
    wire new_Jinkela_wire_6467;
    wire new_Jinkela_wire_4438;
    wire new_Jinkela_wire_6933;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_6609;
    wire new_Jinkela_wire_5872;
    wire _0527_;
    wire _0644_;
    wire new_Jinkela_wire_1904;
    wire new_Jinkela_wire_2594;
    wire _0406_;
    wire new_Jinkela_wire_5472;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_6541;
    wire new_Jinkela_wire_2834;
    wire new_Jinkela_wire_4913;
    wire new_Jinkela_wire_2805;
    wire new_Jinkela_wire_3029;
    wire new_Jinkela_wire_2276;
    wire new_Jinkela_wire_6792;
    wire new_Jinkela_wire_1667;
    wire _0815_;
    wire new_Jinkela_wire_1945;
    wire _1240_;
    wire _0223_;
    wire _0234_;
    wire new_Jinkela_wire_5182;
    wire new_Jinkela_wire_3747;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_6887;
    wire _0753_;
    wire new_Jinkela_wire_5795;
    wire _0488_;
    wire new_Jinkela_wire_6543;
    wire _1093_;
    wire new_Jinkela_wire_2973;
    wire new_Jinkela_wire_7391;
    wire new_Jinkela_wire_4638;
    wire _0981_;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_7335;
    wire _0308_;
    wire new_Jinkela_wire_7079;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_7003;
    wire new_Jinkela_wire_7869;
    wire new_Jinkela_wire_3740;
    wire new_Jinkela_wire_6126;
    wire new_Jinkela_wire_2957;
    wire new_Jinkela_wire_6177;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_2551;
    wire new_Jinkela_wire_5266;
    wire new_Jinkela_wire_7896;
    wire new_Jinkela_wire_999;
    wire _1164_;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_3662;
    wire new_Jinkela_wire_3813;
    wire new_Jinkela_wire_6078;
    wire new_Jinkela_wire_7257;
    wire new_Jinkela_wire_7344;
    wire new_Jinkela_wire_6075;
    wire _0314_;
    wire new_Jinkela_wire_6561;
    wire new_Jinkela_wire_3106;
    wire new_Jinkela_wire_4265;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_5998;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_2896;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_6998;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_3696;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_2282;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_2978;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_6382;
    wire new_Jinkela_wire_2363;
    wire new_Jinkela_wire_3706;
    wire new_Jinkela_wire_6630;
    wire new_Jinkela_wire_4081;
    wire new_Jinkela_wire_7131;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_4051;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_7280;
    wire new_Jinkela_wire_6262;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_125;
    wire _0122_;
    wire new_Jinkela_wire_2335;
    wire new_Jinkela_wire_5987;
    wire _1187_;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_269;
    wire _0461_;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_6170;
    wire new_Jinkela_wire_6518;
    wire _1168_;
    wire new_Jinkela_wire_1463;
    wire _1073_;
    wire new_Jinkela_wire_66;
    wire _1125_;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_4873;
    wire new_Jinkela_wire_2341;
    wire new_Jinkela_wire_4335;
    wire new_Jinkela_wire_5864;
    wire new_Jinkela_wire_4341;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_4819;
    wire new_Jinkela_wire_7942;
    wire new_Jinkela_wire_241;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_2167;
    wire new_Jinkela_wire_6059;
    wire new_Jinkela_wire_3318;
    wire _0409_;
    wire new_Jinkela_wire_5556;
    wire new_Jinkela_wire_3982;
    wire new_Jinkela_wire_1347;
    wire _0498_;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_2427;
    wire new_Jinkela_wire_1308;
    wire _0826_;
    wire new_Jinkela_wire_2890;
    wire new_Jinkela_wire_2365;
    wire new_Jinkela_wire_850;
    wire _0883_;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_7165;
    wire new_Jinkela_wire_2386;
    wire new_Jinkela_wire_4020;
    wire new_Jinkela_wire_3592;
    wire new_Jinkela_wire_2207;
    wire new_Jinkela_wire_4465;
    wire _0513_;
    wire new_Jinkela_wire_2530;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_5487;
    wire new_Jinkela_wire_6652;
    wire new_Jinkela_wire_3897;
    wire _1052_;
    wire new_Jinkela_wire_2228;
    wire new_Jinkela_wire_4309;
    wire new_Jinkela_wire_4482;
    wire new_Jinkela_wire_4849;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_5071;
    wire new_Jinkela_wire_2337;
    wire _0820_;
    wire new_Jinkela_wire_4460;
    wire new_Jinkela_wire_3496;
    wire new_Jinkela_wire_7362;
    wire new_Jinkela_wire_3586;
    wire new_Jinkela_wire_5486;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_4780;
    wire new_Jinkela_wire_4761;
    wire new_Jinkela_wire_7331;
    wire _0069_;
    wire new_Jinkela_wire_3821;
    wire new_net_2385;
    wire new_Jinkela_wire_3719;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_5423;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_2693;
    wire new_Jinkela_wire_2600;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_1666;
    wire new_Jinkela_wire_6033;
    wire new_Jinkela_wire_4038;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_7386;
    wire new_Jinkela_wire_7298;
    wire new_Jinkela_wire_5279;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_4186;
    wire new_Jinkela_wire_4661;
    wire new_Jinkela_wire_7074;
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_5015;
    wire new_Jinkela_wire_1057;
    wire new_Jinkela_wire_3357;
    wire _0348_;
    wire new_Jinkela_wire_5806;
    wire new_Jinkela_wire_5823;
    input G124;
    input G52;
    input G48;
    input G72;
    input G100;
    input G110;
    input G53;
    input G80;
    input G132;
    input G91;
    input G55;
    input G99;
    input G134;
    input G121;
    input G61;
    input G37;
    input G165;
    input G39;
    input G157;
    input G5;
    input G62;
    input G105;
    input G117;
    input G16;
    input G44;
    input G18;
    input G96;
    input G168;
    input G36;
    input G3;
    input G43;
    input G6;
    input G78;
    input G12;
    input G42;
    input G88;
    input G57;
    input G8;
    input G137;
    input G128;
    input G153;
    input G54;
    input G118;
    input G93;
    input G169;
    input G87;
    input G73;
    input G50;
    input G174;
    input G101;
    input G67;
    input G126;
    input G103;
    input G158;
    input G161;
    input G86;
    input G138;
    input G68;
    input G113;
    input G108;
    input G140;
    input G97;
    input G135;
    input G65;
    input G92;
    input G56;
    input G66;
    input G9;
    input G112;
    input G171;
    input G64;
    input G13;
    input G142;
    input G69;
    input G14;
    input G4;
    input G150;
    input G106;
    input G109;
    input G145;
    input G139;
    input G131;
    input G160;
    input G119;
    input G159;
    input G19;
    input G11;
    input G94;
    input G120;
    input G83;
    input G123;
    input G89;
    input G152;
    input G136;
    input G46;
    input G146;
    input G32;
    input G85;
    input G47;
    input G95;
    input G114;
    input G81;
    input G45;
    input G30;
    input G111;
    input G176;
    input G148;
    input G51;
    input G162;
    input G63;
    input G149;
    input G156;
    input G155;
    input G144;
    input G1;
    input G26;
    input G102;
    input G70;
    input G17;
    input G147;
    input G129;
    input G15;
    input G24;
    input G31;
    input G141;
    input G172;
    input G49;
    input G41;
    input G84;
    input G166;
    input G20;
    input G143;
    input G107;
    input G154;
    input G122;
    input G90;
    input G77;
    input G125;
    input G82;
    input G29;
    input G74;
    input G130;
    input G164;
    input G38;
    input G10;
    input G76;
    input G116;
    input G133;
    input G35;
    input G40;
    input G7;
    input G115;
    input G177;
    input G2;
    input G104;
    input G127;
    input G27;
    input G173;
    input G60;
    input G22;
    input G21;
    input G23;
    input G170;
    input G71;
    input G98;
    input G34;
    input G33;
    input G163;
    input G59;
    input G75;
    input G167;
    input G175;
    input G28;
    input G58;
    input G79;
    input G151;
    input G178;
    input G25;
    output G5314;
    output G5252;
    output G5193;
    output G5196;
    output G5236;
    output G5269;
    output G5233;
    output G5223;
    output G5301;
    output G5231;
    output G5273;
    output G5279;
    output G5227;
    output G5262;
    output G5281;
    output G5234;
    output G5272;
    output G5228;
    output G5213;
    output G5244;
    output G5298;
    output G5240;
    output G5280;
    output G5232;
    output G5219;
    output G5218;
    output G5224;
    output G5241;
    output G5297;
    output G5274;
    output G5302;
    output G5289;
    output G5270;
    output G5290;
    output G5308;
    output G5215;
    output G5243;
    output G5287;
    output G5211;
    output G5249;
    output G5286;
    output G5205;
    output G5250;
    output G5299;
    output G5296;
    output G5230;
    output G5248;
    output G5292;
    output G5258;
    output G5263;
    output G5245;
    output G5197;
    output G5267;
    output G5275;
    output G5257;
    output G5271;
    output G5208;
    output G5210;
    output G5293;
    output G5204;
    output G5304;
    output G5239;
    output G5237;
    output G5261;
    output G5229;
    output G5238;
    output G5260;
    output G5266;
    output G5300;
    output G5303;
    output G5288;
    output G5311;
    output G5251;
    output G5313;
    output G5235;
    output G5246;
    output G5255;
    output G5291;
    output G5203;
    output G5195;
    output G5295;
    output G5264;
    output G5282;
    output G5259;
    output G5309;
    output G5256;
    output G5285;
    output G5194;
    output G5209;
    output G5242;
    output G5247;
    output G5207;
    output G5310;
    output G5226;
    output G5222;
    output G5315;
    output G5201;
    output G5220;
    output G5265;
    output G5225;
    output G5199;
    output G5278;
    output G5202;
    output G5206;
    output G5221;
    output G5307;
    output G5312;
    output G5294;
    output G5306;
    output G5253;
    output G5254;
    output G5284;
    output G5200;
    output G5214;
    output G5212;
    output G5217;
    output G5198;
    output G5216;
    output G5305;
    output G5276;
    output G5277;
    output G5268;
    output G5283;

    bfr new_Jinkela_buffer_4943 (
        .din(new_Jinkela_wire_6737),
        .dout(new_Jinkela_wire_6738)
    );

    bfr new_Jinkela_buffer_4964 (
        .din(new_Jinkela_wire_6771),
        .dout(new_Jinkela_wire_6772)
    );

    bfr new_Jinkela_buffer_4944 (
        .din(new_Jinkela_wire_6738),
        .dout(new_Jinkela_wire_6739)
    );

    spl2 new_Jinkela_splitter_702 (
        .a(new_Jinkela_wire_6848),
        .b(new_Jinkela_wire_6849),
        .c(new_Jinkela_wire_6850)
    );

    bfr new_Jinkela_buffer_4982 (
        .din(new_Jinkela_wire_6790),
        .dout(new_Jinkela_wire_6791)
    );

    bfr new_Jinkela_buffer_4945 (
        .din(new_Jinkela_wire_6739),
        .dout(new_Jinkela_wire_6740)
    );

    bfr new_Jinkela_buffer_4965 (
        .din(new_Jinkela_wire_6772),
        .dout(new_Jinkela_wire_6773)
    );

    bfr new_Jinkela_buffer_4946 (
        .din(new_Jinkela_wire_6740),
        .dout(new_Jinkela_wire_6741)
    );

    bfr new_Jinkela_buffer_5056 (
        .din(_0783_),
        .dout(new_Jinkela_wire_6892)
    );

    bfr new_Jinkela_buffer_4947 (
        .din(new_Jinkela_wire_6741),
        .dout(new_Jinkela_wire_6742)
    );

    bfr new_Jinkela_buffer_4966 (
        .din(new_Jinkela_wire_6773),
        .dout(new_Jinkela_wire_6774)
    );

    bfr new_Jinkela_buffer_4948 (
        .din(new_Jinkela_wire_6742),
        .dout(new_Jinkela_wire_6743)
    );

    bfr new_Jinkela_buffer_4983 (
        .din(new_Jinkela_wire_6796),
        .dout(new_Jinkela_wire_6797)
    );

    bfr new_Jinkela_buffer_4949 (
        .din(new_Jinkela_wire_6743),
        .dout(new_Jinkela_wire_6744)
    );

    bfr new_Jinkela_buffer_4967 (
        .din(new_Jinkela_wire_6774),
        .dout(new_Jinkela_wire_6775)
    );

    bfr new_Jinkela_buffer_4950 (
        .din(new_Jinkela_wire_6744),
        .dout(new_Jinkela_wire_6745)
    );

    spl4L new_Jinkela_splitter_693 (
        .a(new_Jinkela_wire_6792),
        .d(new_Jinkela_wire_6793),
        .e(new_Jinkela_wire_6794),
        .b(new_Jinkela_wire_6795),
        .c(new_Jinkela_wire_6796)
    );

    bfr new_Jinkela_buffer_4951 (
        .din(new_Jinkela_wire_6745),
        .dout(new_Jinkela_wire_6746)
    );

    bfr new_Jinkela_buffer_4968 (
        .din(new_Jinkela_wire_6775),
        .dout(new_Jinkela_wire_6776)
    );

    bfr new_Jinkela_buffer_4952 (
        .din(new_Jinkela_wire_6746),
        .dout(new_Jinkela_wire_6747)
    );

    bfr new_Jinkela_buffer_4953 (
        .din(new_Jinkela_wire_6747),
        .dout(new_Jinkela_wire_6748)
    );

    bfr new_Jinkela_buffer_4969 (
        .din(new_Jinkela_wire_6776),
        .dout(new_Jinkela_wire_6777)
    );

    bfr new_Jinkela_buffer_4954 (
        .din(new_Jinkela_wire_6748),
        .dout(new_Jinkela_wire_6749)
    );

    bfr new_Jinkela_buffer_4970 (
        .din(new_Jinkela_wire_6777),
        .dout(new_Jinkela_wire_6778)
    );

    bfr new_Jinkela_buffer_4984 (
        .din(new_Jinkela_wire_6797),
        .dout(new_Jinkela_wire_6798)
    );

    bfr new_Jinkela_buffer_4971 (
        .din(new_Jinkela_wire_6778),
        .dout(new_Jinkela_wire_6779)
    );

    spl2 new_Jinkela_splitter_704 (
        .a(_0055_),
        .b(new_Jinkela_wire_6890),
        .c(new_Jinkela_wire_6891)
    );

    bfr new_Jinkela_buffer_4972 (
        .din(new_Jinkela_wire_6779),
        .dout(new_Jinkela_wire_6780)
    );

    bfr new_Jinkela_buffer_4985 (
        .din(new_Jinkela_wire_6798),
        .dout(new_Jinkela_wire_6799)
    );

    bfr new_Jinkela_buffer_4973 (
        .din(new_Jinkela_wire_6780),
        .dout(new_Jinkela_wire_6781)
    );

    bfr new_Jinkela_buffer_5017 (
        .din(new_net_2),
        .dout(new_Jinkela_wire_6847)
    );

    spl2 new_Jinkela_splitter_703 (
        .a(_0247_),
        .b(new_Jinkela_wire_6888),
        .c(new_Jinkela_wire_6889)
    );

    bfr new_Jinkela_buffer_4974 (
        .din(new_Jinkela_wire_6781),
        .dout(new_Jinkela_wire_6782)
    );

    bfr new_Jinkela_buffer_4986 (
        .din(new_Jinkela_wire_6799),
        .dout(new_Jinkela_wire_6800)
    );

    bfr new_Jinkela_buffer_4975 (
        .din(new_Jinkela_wire_6782),
        .dout(new_Jinkela_wire_6783)
    );

    bfr new_Jinkela_buffer_4991 (
        .din(new_Jinkela_wire_6804),
        .dout(new_Jinkela_wire_6805)
    );

    bfr new_Jinkela_buffer_5019 (
        .din(new_Jinkela_wire_6850),
        .dout(new_Jinkela_wire_6851)
    );

    bfr new_Jinkela_buffer_4976 (
        .din(new_Jinkela_wire_6783),
        .dout(new_Jinkela_wire_6784)
    );

    bfr new_Jinkela_buffer_4987 (
        .din(new_Jinkela_wire_6800),
        .dout(new_Jinkela_wire_6801)
    );

    bfr new_Jinkela_buffer_4977 (
        .din(new_Jinkela_wire_6784),
        .dout(new_Jinkela_wire_6785)
    );

    bfr new_Jinkela_buffer_5018 (
        .din(new_Jinkela_wire_6847),
        .dout(new_Jinkela_wire_6848)
    );

    bfr new_Jinkela_buffer_4978 (
        .din(new_Jinkela_wire_6785),
        .dout(new_Jinkela_wire_6786)
    );

    bfr new_Jinkela_buffer_4988 (
        .din(new_Jinkela_wire_6801),
        .dout(new_Jinkela_wire_6802)
    );

    bfr new_Jinkela_buffer_2307 (
        .din(new_Jinkela_wire_3511),
        .dout(new_Jinkela_wire_3512)
    );

    spl2 new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_380),
        .b(new_Jinkela_wire_381),
        .c(new_Jinkela_wire_382)
    );

    bfr new_Jinkela_buffer_3687 (
        .din(new_Jinkela_wire_5159),
        .dout(new_Jinkela_wire_5160)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_2328 (
        .din(new_Jinkela_wire_3548),
        .dout(new_Jinkela_wire_3549)
    );

    bfr new_Jinkela_buffer_3644 (
        .din(new_Jinkela_wire_5102),
        .dout(new_Jinkela_wire_5103)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_3666 (
        .din(new_Jinkela_wire_5136),
        .dout(new_Jinkela_wire_5137)
    );

    bfr new_Jinkela_buffer_2308 (
        .din(new_Jinkela_wire_3512),
        .dout(new_Jinkela_wire_3513)
    );

    bfr new_Jinkela_buffer_3645 (
        .din(new_Jinkela_wire_5103),
        .dout(new_Jinkela_wire_5104)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    bfr new_Jinkela_buffer_2329 (
        .din(new_Jinkela_wire_3549),
        .dout(new_Jinkela_wire_3550)
    );

    bfr new_Jinkela_buffer_2309 (
        .din(new_Jinkela_wire_3513),
        .dout(new_Jinkela_wire_3514)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_3646 (
        .din(new_Jinkela_wire_5104),
        .dout(new_Jinkela_wire_5105)
    );

    bfr new_Jinkela_buffer_210 (
        .din(G97),
        .dout(new_Jinkela_wire_538)
    );

    bfr new_Jinkela_buffer_2358 (
        .din(new_Jinkela_wire_3581),
        .dout(new_Jinkela_wire_3582)
    );

    bfr new_Jinkela_buffer_3667 (
        .din(new_Jinkela_wire_5137),
        .dout(new_Jinkela_wire_5138)
    );

    bfr new_Jinkela_buffer_2310 (
        .din(new_Jinkela_wire_3514),
        .dout(new_Jinkela_wire_3515)
    );

    spl2 new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_384),
        .b(new_Jinkela_wire_385),
        .c(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_3647 (
        .din(new_Jinkela_wire_5105),
        .dout(new_Jinkela_wire_5106)
    );

    spl2 new_Jinkela_splitter_78 (
        .a(new_Jinkela_wire_386),
        .b(new_Jinkela_wire_387),
        .c(new_Jinkela_wire_388)
    );

    bfr new_Jinkela_buffer_2330 (
        .din(new_Jinkela_wire_3550),
        .dout(new_Jinkela_wire_3551)
    );

    bfr new_Jinkela_buffer_3688 (
        .din(new_Jinkela_wire_5160),
        .dout(new_Jinkela_wire_5161)
    );

    spl2 new_Jinkela_splitter_453 (
        .a(new_Jinkela_wire_3515),
        .b(new_Jinkela_wire_3516),
        .c(new_Jinkela_wire_3517)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    bfr new_Jinkela_buffer_3648 (
        .din(new_Jinkela_wire_5106),
        .dout(new_Jinkela_wire_5107)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    spl2 new_Jinkela_splitter_454 (
        .a(new_Jinkela_wire_3517),
        .b(new_Jinkela_wire_3518),
        .c(new_Jinkela_wire_3519)
    );

    spl2 new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_388),
        .b(new_Jinkela_wire_389),
        .c(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_3668 (
        .din(new_Jinkela_wire_5138),
        .dout(new_Jinkela_wire_5139)
    );

    spl4L new_Jinkela_splitter_461 (
        .a(new_Jinkela_wire_3583),
        .d(new_Jinkela_wire_3584),
        .e(new_Jinkela_wire_3585),
        .b(new_Jinkela_wire_3586),
        .c(new_Jinkela_wire_3587)
    );

    bfr new_Jinkela_buffer_3649 (
        .din(new_Jinkela_wire_5107),
        .dout(new_Jinkela_wire_5108)
    );

    bfr new_Jinkela_buffer_2311 (
        .din(new_Jinkela_wire_3519),
        .dout(new_Jinkela_wire_3520)
    );

    spl3L new_Jinkela_splitter_80 (
        .a(new_Jinkela_wire_390),
        .d(new_Jinkela_wire_391),
        .b(new_Jinkela_wire_392),
        .c(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_3726 (
        .din(_1223_),
        .dout(new_Jinkela_wire_5201)
    );

    bfr new_Jinkela_buffer_2362 (
        .din(new_Jinkela_wire_3591),
        .dout(new_Jinkela_wire_3592)
    );

    bfr new_Jinkela_buffer_3721 (
        .din(new_Jinkela_wire_5193),
        .dout(new_Jinkela_wire_5194)
    );

    bfr new_Jinkela_buffer_2331 (
        .din(new_Jinkela_wire_3551),
        .dout(new_Jinkela_wire_3552)
    );

    bfr new_Jinkela_buffer_3650 (
        .din(new_Jinkela_wire_5108),
        .dout(new_Jinkela_wire_5109)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    bfr new_Jinkela_buffer_3669 (
        .din(new_Jinkela_wire_5139),
        .dout(new_Jinkela_wire_5140)
    );

    spl2 new_Jinkela_splitter_455 (
        .a(new_Jinkela_wire_3520),
        .b(new_Jinkela_wire_3521),
        .c(new_Jinkela_wire_3522)
    );

    spl4L new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_393),
        .d(new_Jinkela_wire_394),
        .e(new_Jinkela_wire_395),
        .b(new_Jinkela_wire_396),
        .c(new_Jinkela_wire_397)
    );

    bfr new_Jinkela_buffer_3651 (
        .din(new_Jinkela_wire_5109),
        .dout(new_Jinkela_wire_5110)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    spl2 new_Jinkela_splitter_463 (
        .a(_0736_),
        .b(new_Jinkela_wire_3610),
        .c(new_Jinkela_wire_3611)
    );

    bfr new_Jinkela_buffer_3689 (
        .din(new_Jinkela_wire_5161),
        .dout(new_Jinkela_wire_5162)
    );

    spl2 new_Jinkela_splitter_464 (
        .a(new_net_17),
        .b(new_Jinkela_wire_3613),
        .c(new_Jinkela_wire_3615)
    );

    bfr new_Jinkela_buffer_2332 (
        .din(new_Jinkela_wire_3552),
        .dout(new_Jinkela_wire_3553)
    );

    bfr new_Jinkela_buffer_3652 (
        .din(new_Jinkela_wire_5110),
        .dout(new_Jinkela_wire_5111)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    bfr new_Jinkela_buffer_2360 (
        .din(new_Jinkela_wire_3587),
        .dout(new_Jinkela_wire_3588)
    );

    bfr new_Jinkela_buffer_2333 (
        .din(new_Jinkela_wire_3553),
        .dout(new_Jinkela_wire_3554)
    );

    bfr new_Jinkela_buffer_3670 (
        .din(new_Jinkela_wire_5140),
        .dout(new_Jinkela_wire_5141)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_3653 (
        .din(new_Jinkela_wire_5111),
        .dout(new_Jinkela_wire_5112)
    );

    bfr new_Jinkela_buffer_2334 (
        .din(new_Jinkela_wire_3554),
        .dout(new_Jinkela_wire_3555)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_2380 (
        .din(new_Jinkela_wire_3611),
        .dout(new_Jinkela_wire_3612)
    );

    bfr new_Jinkela_buffer_3654 (
        .din(new_Jinkela_wire_5112),
        .dout(new_Jinkela_wire_5113)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_2335 (
        .din(new_Jinkela_wire_3555),
        .dout(new_Jinkela_wire_3556)
    );

    bfr new_Jinkela_buffer_3671 (
        .din(new_Jinkela_wire_5141),
        .dout(new_Jinkela_wire_5142)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(new_Jinkela_wire_513),
        .b(new_Jinkela_wire_514),
        .c(new_Jinkela_wire_515)
    );

    spl4L new_Jinkela_splitter_110 (
        .a(new_Jinkela_wire_521),
        .d(new_Jinkela_wire_522),
        .e(new_Jinkela_wire_523),
        .b(new_Jinkela_wire_524),
        .c(new_Jinkela_wire_525)
    );

    spl2 new_Jinkela_splitter_462 (
        .a(new_Jinkela_wire_3588),
        .b(new_Jinkela_wire_3589),
        .c(new_Jinkela_wire_3590)
    );

    bfr new_Jinkela_buffer_3690 (
        .din(new_Jinkela_wire_5162),
        .dout(new_Jinkela_wire_5163)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    bfr new_Jinkela_buffer_2336 (
        .din(new_Jinkela_wire_3556),
        .dout(new_Jinkela_wire_3557)
    );

    bfr new_Jinkela_buffer_3672 (
        .din(new_Jinkela_wire_5142),
        .dout(new_Jinkela_wire_5143)
    );

    spl3L new_Jinkela_splitter_111 (
        .a(new_Jinkela_wire_525),
        .d(new_Jinkela_wire_526),
        .b(new_Jinkela_wire_527),
        .c(new_Jinkela_wire_528)
    );

    bfr new_Jinkela_buffer_3724 (
        .din(new_Jinkela_wire_5198),
        .dout(new_Jinkela_wire_5199)
    );

    bfr new_Jinkela_buffer_3722 (
        .din(new_Jinkela_wire_5194),
        .dout(new_Jinkela_wire_5195)
    );

    bfr new_Jinkela_buffer_2337 (
        .din(new_Jinkela_wire_3557),
        .dout(new_Jinkela_wire_3558)
    );

    bfr new_Jinkela_buffer_3673 (
        .din(new_Jinkela_wire_5143),
        .dout(new_Jinkela_wire_5144)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_468),
        .dout(new_Jinkela_wire_469)
    );

    bfr new_Jinkela_buffer_2363 (
        .din(new_Jinkela_wire_3592),
        .dout(new_Jinkela_wire_3593)
    );

    bfr new_Jinkela_buffer_3691 (
        .din(new_Jinkela_wire_5163),
        .dout(new_Jinkela_wire_5164)
    );

    spl2 new_Jinkela_splitter_109 (
        .a(new_Jinkela_wire_518),
        .b(new_Jinkela_wire_519),
        .c(new_Jinkela_wire_520)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    bfr new_Jinkela_buffer_2338 (
        .din(new_Jinkela_wire_3558),
        .dout(new_Jinkela_wire_3559)
    );

    bfr new_Jinkela_buffer_3674 (
        .din(new_Jinkela_wire_5144),
        .dout(new_Jinkela_wire_5145)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_469),
        .dout(new_Jinkela_wire_470)
    );

    bfr new_Jinkela_buffer_2364 (
        .din(new_Jinkela_wire_3593),
        .dout(new_Jinkela_wire_3594)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(G140),
        .b(new_Jinkela_wire_531),
        .c(new_Jinkela_wire_532)
    );

    bfr new_Jinkela_buffer_2339 (
        .din(new_Jinkela_wire_3559),
        .dout(new_Jinkela_wire_3560)
    );

    bfr new_Jinkela_buffer_3675 (
        .din(new_Jinkela_wire_5145),
        .dout(new_Jinkela_wire_5146)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_470),
        .dout(new_Jinkela_wire_471)
    );

    spl2 new_Jinkela_splitter_466 (
        .a(_1081_),
        .b(new_Jinkela_wire_3627),
        .c(new_Jinkela_wire_3628)
    );

    bfr new_Jinkela_buffer_3692 (
        .din(new_Jinkela_wire_5164),
        .dout(new_Jinkela_wire_5165)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_2340 (
        .din(new_Jinkela_wire_3560),
        .dout(new_Jinkela_wire_3561)
    );

    bfr new_Jinkela_buffer_3676 (
        .din(new_Jinkela_wire_5146),
        .dout(new_Jinkela_wire_5147)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_2365 (
        .din(new_Jinkela_wire_3594),
        .dout(new_Jinkela_wire_3595)
    );

    bfr new_Jinkela_buffer_3738 (
        .din(_0271_),
        .dout(new_Jinkela_wire_5213)
    );

    spl2 new_Jinkela_splitter_559 (
        .a(new_Jinkela_wire_5195),
        .b(new_Jinkela_wire_5196),
        .c(new_Jinkela_wire_5197)
    );

    bfr new_Jinkela_buffer_2341 (
        .din(new_Jinkela_wire_3561),
        .dout(new_Jinkela_wire_3562)
    );

    bfr new_Jinkela_buffer_3677 (
        .din(new_Jinkela_wire_5147),
        .dout(new_Jinkela_wire_5148)
    );

    spl2 new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_472),
        .b(new_Jinkela_wire_473),
        .c(new_Jinkela_wire_474)
    );

    bfr new_Jinkela_buffer_2381 (
        .din(new_Jinkela_wire_3613),
        .dout(new_Jinkela_wire_3614)
    );

    bfr new_Jinkela_buffer_3693 (
        .din(new_Jinkela_wire_5165),
        .dout(new_Jinkela_wire_5166)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_474),
        .dout(new_Jinkela_wire_475)
    );

    bfr new_Jinkela_buffer_2342 (
        .din(new_Jinkela_wire_3562),
        .dout(new_Jinkela_wire_3563)
    );

    bfr new_Jinkela_buffer_3678 (
        .din(new_Jinkela_wire_5148),
        .dout(new_Jinkela_wire_5149)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(G135),
        .b(new_Jinkela_wire_540),
        .c(new_Jinkela_wire_541)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_532),
        .dout(new_Jinkela_wire_533)
    );

    bfr new_Jinkela_buffer_2366 (
        .din(new_Jinkela_wire_3595),
        .dout(new_Jinkela_wire_3596)
    );

    bfr new_Jinkela_buffer_216 (
        .din(G65),
        .dout(new_Jinkela_wire_548)
    );

    bfr new_Jinkela_buffer_2343 (
        .din(new_Jinkela_wire_3563),
        .dout(new_Jinkela_wire_3564)
    );

    bfr new_Jinkela_buffer_3679 (
        .din(new_Jinkela_wire_5149),
        .dout(new_Jinkela_wire_5150)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_475),
        .dout(new_Jinkela_wire_476)
    );

    spl4L new_Jinkela_splitter_465 (
        .a(new_Jinkela_wire_3615),
        .d(new_Jinkela_wire_3616),
        .e(new_Jinkela_wire_3617),
        .b(new_Jinkela_wire_3618),
        .c(new_Jinkela_wire_3619)
    );

    bfr new_Jinkela_buffer_3694 (
        .din(new_Jinkela_wire_5166),
        .dout(new_Jinkela_wire_5167)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    bfr new_Jinkela_buffer_2344 (
        .din(new_Jinkela_wire_3564),
        .dout(new_Jinkela_wire_3565)
    );

    bfr new_Jinkela_buffer_3680 (
        .din(new_Jinkela_wire_5150),
        .dout(new_Jinkela_wire_5151)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_2367 (
        .din(new_Jinkela_wire_3596),
        .dout(new_Jinkela_wire_3597)
    );

    bfr new_Jinkela_buffer_3725 (
        .din(new_Jinkela_wire_5199),
        .dout(new_Jinkela_wire_5200)
    );

    spl3L new_Jinkela_splitter_424 (
        .a(new_Jinkela_wire_3308),
        .d(new_Jinkela_wire_3309),
        .b(new_Jinkela_wire_3310),
        .c(new_Jinkela_wire_3311)
    );

    bfr new_Jinkela_buffer_2131 (
        .din(new_Jinkela_wire_3247),
        .dout(new_Jinkela_wire_3248)
    );

    bfr new_Jinkela_buffer_338 (
        .din(G106),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    bfr new_Jinkela_buffer_2154 (
        .din(new_Jinkela_wire_3284),
        .dout(new_Jinkela_wire_3285)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_2132 (
        .din(new_Jinkela_wire_3248),
        .dout(new_Jinkela_wire_3249)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    bfr new_Jinkela_buffer_2178 (
        .din(new_Jinkela_wire_3317),
        .dout(new_Jinkela_wire_3318)
    );

    bfr new_Jinkela_buffer_2155 (
        .din(new_Jinkela_wire_3285),
        .dout(new_Jinkela_wire_3286)
    );

    spl2 new_Jinkela_splitter_137 (
        .a(new_Jinkela_wire_721),
        .b(new_Jinkela_wire_722),
        .c(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    bfr new_Jinkela_buffer_2156 (
        .din(new_Jinkela_wire_3286),
        .dout(new_Jinkela_wire_3287)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    spl4L new_Jinkela_splitter_425 (
        .a(new_Jinkela_wire_3312),
        .d(new_Jinkela_wire_3313),
        .e(new_Jinkela_wire_3314),
        .b(new_Jinkela_wire_3315),
        .c(new_Jinkela_wire_3316)
    );

    spl2 new_Jinkela_splitter_428 (
        .a(_0774_),
        .b(new_Jinkela_wire_3372),
        .c(new_Jinkela_wire_3373)
    );

    bfr new_Jinkela_buffer_2157 (
        .din(new_Jinkela_wire_3287),
        .dout(new_Jinkela_wire_3288)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    bfr new_Jinkela_buffer_2179 (
        .din(new_Jinkela_wire_3318),
        .dout(new_Jinkela_wire_3319)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_731),
        .dout(new_Jinkela_wire_732)
    );

    bfr new_Jinkela_buffer_2158 (
        .din(new_Jinkela_wire_3288),
        .dout(new_Jinkela_wire_3289)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    spl3L new_Jinkela_splitter_426 (
        .a(_0873_),
        .d(new_Jinkela_wire_3356),
        .b(new_Jinkela_wire_3357),
        .c(new_Jinkela_wire_3358)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_2159 (
        .din(new_Jinkela_wire_3289),
        .dout(new_Jinkela_wire_3290)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(new_Jinkela_wire_726),
        .b(new_Jinkela_wire_727),
        .c(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_660),
        .dout(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_2181 (
        .din(new_Jinkela_wire_3320),
        .dout(new_Jinkela_wire_3321)
    );

    bfr new_Jinkela_buffer_2160 (
        .din(new_Jinkela_wire_3290),
        .dout(new_Jinkela_wire_3291)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    spl2 new_Jinkela_splitter_434 (
        .a(_1025_),
        .b(new_Jinkela_wire_3390),
        .c(new_Jinkela_wire_3391)
    );

    spl3L new_Jinkela_splitter_430 (
        .a(_0103_),
        .d(new_Jinkela_wire_3377),
        .b(new_Jinkela_wire_3380),
        .c(new_Jinkela_wire_3385)
    );

    bfr new_Jinkela_buffer_2161 (
        .din(new_Jinkela_wire_3291),
        .dout(new_Jinkela_wire_3292)
    );

    spl3L new_Jinkela_splitter_125 (
        .a(new_Jinkela_wire_662),
        .d(new_Jinkela_wire_663),
        .b(new_Jinkela_wire_664),
        .c(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_2182 (
        .din(new_Jinkela_wire_3321),
        .dout(new_Jinkela_wire_3322)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_2162 (
        .din(new_Jinkela_wire_3292),
        .dout(new_Jinkela_wire_3293)
    );

    spl2 new_Jinkela_splitter_141 (
        .a(G109),
        .b(new_Jinkela_wire_740),
        .c(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_665),
        .dout(new_Jinkela_wire_666)
    );

    bfr new_Jinkela_buffer_2163 (
        .din(new_Jinkela_wire_3293),
        .dout(new_Jinkela_wire_3294)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_666),
        .dout(new_Jinkela_wire_667)
    );

    bfr new_Jinkela_buffer_2183 (
        .din(new_Jinkela_wire_3322),
        .dout(new_Jinkela_wire_3323)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_2164 (
        .din(new_Jinkela_wire_3294),
        .dout(new_Jinkela_wire_3295)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_667),
        .dout(new_Jinkela_wire_668)
    );

    bfr new_Jinkela_buffer_2216 (
        .din(new_Jinkela_wire_3358),
        .dout(new_Jinkela_wire_3359)
    );

    bfr new_Jinkela_buffer_2165 (
        .din(new_Jinkela_wire_3295),
        .dout(new_Jinkela_wire_3296)
    );

    spl3L new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_668),
        .d(new_Jinkela_wire_669),
        .b(new_Jinkela_wire_670),
        .c(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_2184 (
        .din(new_Jinkela_wire_3323),
        .dout(new_Jinkela_wire_3324)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(new_Jinkela_wire_733),
        .b(new_Jinkela_wire_734),
        .c(new_Jinkela_wire_735)
    );

    bfr new_Jinkela_buffer_2166 (
        .din(new_Jinkela_wire_3296),
        .dout(new_Jinkela_wire_3297)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    spl4L new_Jinkela_splitter_432 (
        .a(new_Jinkela_wire_3380),
        .d(new_Jinkela_wire_3381),
        .e(new_Jinkela_wire_3382),
        .b(new_Jinkela_wire_3383),
        .c(new_Jinkela_wire_3384)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    bfr new_Jinkela_buffer_2167 (
        .din(new_Jinkela_wire_3297),
        .dout(new_Jinkela_wire_3298)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_2185 (
        .din(new_Jinkela_wire_3324),
        .dout(new_Jinkela_wire_3325)
    );

    spl4L new_Jinkela_splitter_142 (
        .a(new_Jinkela_wire_742),
        .d(new_Jinkela_wire_743),
        .e(new_Jinkela_wire_744),
        .b(new_Jinkela_wire_746),
        .c(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_2168 (
        .din(new_Jinkela_wire_3298),
        .dout(new_Jinkela_wire_3299)
    );

    spl2 new_Jinkela_splitter_127 (
        .a(new_Jinkela_wire_673),
        .b(new_Jinkela_wire_674),
        .c(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_2217 (
        .din(new_Jinkela_wire_3359),
        .dout(new_Jinkela_wire_3360)
    );

    spl4L new_Jinkela_splitter_128 (
        .a(new_Jinkela_wire_676),
        .d(new_Jinkela_wire_677),
        .e(new_Jinkela_wire_678),
        .b(new_Jinkela_wire_679),
        .c(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_2169 (
        .din(new_Jinkela_wire_3299),
        .dout(new_Jinkela_wire_3300)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_2186 (
        .din(new_Jinkela_wire_3325),
        .dout(new_Jinkela_wire_3326)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(G145),
        .b(new_Jinkela_wire_756),
        .c(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_2170 (
        .din(new_Jinkela_wire_3300),
        .dout(new_Jinkela_wire_3301)
    );

    spl3L new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_680),
        .d(new_Jinkela_wire_681),
        .b(new_Jinkela_wire_682),
        .c(new_Jinkela_wire_683)
    );

    bfr new_Jinkela_buffer_2227 (
        .din(new_Jinkela_wire_3373),
        .dout(new_Jinkela_wire_3374)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_2171 (
        .din(new_Jinkela_wire_3301),
        .dout(new_Jinkela_wire_3302)
    );

    bfr new_Jinkela_buffer_2187 (
        .din(new_Jinkela_wire_3326),
        .dout(new_Jinkela_wire_3327)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(G139),
        .b(new_Jinkela_wire_765),
        .c(new_Jinkela_wire_766)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_2172 (
        .din(new_Jinkela_wire_3302),
        .dout(new_Jinkela_wire_3303)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_2218 (
        .din(new_Jinkela_wire_3360),
        .dout(new_Jinkela_wire_3361)
    );

    spl4L new_Jinkela_splitter_143 (
        .a(new_Jinkela_wire_746),
        .d(new_Jinkela_wire_747),
        .e(new_Jinkela_wire_748),
        .b(new_Jinkela_wire_749),
        .c(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_2173 (
        .din(new_Jinkela_wire_3303),
        .dout(new_Jinkela_wire_3304)
    );

    bfr new_Jinkela_buffer_2188 (
        .din(new_Jinkela_wire_3327),
        .dout(new_Jinkela_wire_3328)
    );

    bfr new_Jinkela_buffer_3143 (
        .din(new_Jinkela_wire_4500),
        .dout(new_Jinkela_wire_4501)
    );

    bfr new_Jinkela_buffer_3156 (
        .din(new_Jinkela_wire_4513),
        .dout(new_Jinkela_wire_4514)
    );

    bfr new_Jinkela_buffer_3144 (
        .din(new_Jinkela_wire_4501),
        .dout(new_Jinkela_wire_4502)
    );

    bfr new_Jinkela_buffer_3185 (
        .din(new_net_2423),
        .dout(new_Jinkela_wire_4547)
    );

    bfr new_Jinkela_buffer_3145 (
        .din(new_Jinkela_wire_4502),
        .dout(new_Jinkela_wire_4503)
    );

    bfr new_Jinkela_buffer_3157 (
        .din(new_Jinkela_wire_4514),
        .dout(new_Jinkela_wire_4515)
    );

    bfr new_Jinkela_buffer_3146 (
        .din(new_Jinkela_wire_4503),
        .dout(new_Jinkela_wire_4504)
    );

    bfr new_Jinkela_buffer_3176 (
        .din(new_Jinkela_wire_4537),
        .dout(new_Jinkela_wire_4538)
    );

    bfr new_Jinkela_buffer_3147 (
        .din(new_Jinkela_wire_4504),
        .dout(new_Jinkela_wire_4505)
    );

    bfr new_Jinkela_buffer_3158 (
        .din(new_Jinkela_wire_4515),
        .dout(new_Jinkela_wire_4516)
    );

    bfr new_Jinkela_buffer_3148 (
        .din(new_Jinkela_wire_4505),
        .dout(new_Jinkela_wire_4506)
    );

    spl3L new_Jinkela_splitter_518 (
        .a(_0672_),
        .d(new_Jinkela_wire_4568),
        .b(new_Jinkela_wire_4569),
        .c(new_Jinkela_wire_4570)
    );

    spl2 new_Jinkela_splitter_519 (
        .a(_0583_),
        .b(new_Jinkela_wire_4571),
        .c(new_Jinkela_wire_4575)
    );

    bfr new_Jinkela_buffer_3149 (
        .din(new_Jinkela_wire_4506),
        .dout(new_Jinkela_wire_4507)
    );

    bfr new_Jinkela_buffer_3159 (
        .din(new_Jinkela_wire_4516),
        .dout(new_Jinkela_wire_4517)
    );

    bfr new_Jinkela_buffer_3177 (
        .din(new_Jinkela_wire_4538),
        .dout(new_Jinkela_wire_4539)
    );

    bfr new_Jinkela_buffer_3160 (
        .din(new_Jinkela_wire_4517),
        .dout(new_Jinkela_wire_4518)
    );

    bfr new_Jinkela_buffer_3186 (
        .din(new_Jinkela_wire_4547),
        .dout(new_Jinkela_wire_4548)
    );

    bfr new_Jinkela_buffer_3161 (
        .din(new_Jinkela_wire_4518),
        .dout(new_Jinkela_wire_4519)
    );

    bfr new_Jinkela_buffer_3178 (
        .din(new_Jinkela_wire_4539),
        .dout(new_Jinkela_wire_4540)
    );

    bfr new_Jinkela_buffer_3162 (
        .din(new_Jinkela_wire_4519),
        .dout(new_Jinkela_wire_4520)
    );

    spl2 new_Jinkela_splitter_524 (
        .a(_0741_),
        .b(new_Jinkela_wire_4603),
        .c(new_Jinkela_wire_4604)
    );

    bfr new_Jinkela_buffer_3163 (
        .din(new_Jinkela_wire_4520),
        .dout(new_Jinkela_wire_4521)
    );

    bfr new_Jinkela_buffer_3179 (
        .din(new_Jinkela_wire_4540),
        .dout(new_Jinkela_wire_4541)
    );

    bfr new_Jinkela_buffer_3164 (
        .din(new_Jinkela_wire_4521),
        .dout(new_Jinkela_wire_4522)
    );

    bfr new_Jinkela_buffer_3187 (
        .din(new_Jinkela_wire_4548),
        .dout(new_Jinkela_wire_4549)
    );

    bfr new_Jinkela_buffer_3165 (
        .din(new_Jinkela_wire_4522),
        .dout(new_Jinkela_wire_4523)
    );

    bfr new_Jinkela_buffer_3180 (
        .din(new_Jinkela_wire_4541),
        .dout(new_Jinkela_wire_4542)
    );

    bfr new_Jinkela_buffer_3166 (
        .din(new_Jinkela_wire_4523),
        .dout(new_Jinkela_wire_4524)
    );

    bfr new_Jinkela_buffer_3224 (
        .din(_0221_),
        .dout(new_Jinkela_wire_4600)
    );

    bfr new_Jinkela_buffer_3167 (
        .din(new_Jinkela_wire_4524),
        .dout(new_Jinkela_wire_4525)
    );

    bfr new_Jinkela_buffer_3181 (
        .din(new_Jinkela_wire_4542),
        .dout(new_Jinkela_wire_4543)
    );

    bfr new_Jinkela_buffer_3168 (
        .din(new_Jinkela_wire_4525),
        .dout(new_Jinkela_wire_4526)
    );

    bfr new_Jinkela_buffer_3188 (
        .din(new_Jinkela_wire_4549),
        .dout(new_Jinkela_wire_4550)
    );

    bfr new_Jinkela_buffer_3169 (
        .din(new_Jinkela_wire_4526),
        .dout(new_Jinkela_wire_4527)
    );

    bfr new_Jinkela_buffer_3182 (
        .din(new_Jinkela_wire_4543),
        .dout(new_Jinkela_wire_4544)
    );

    bfr new_Jinkela_buffer_3170 (
        .din(new_Jinkela_wire_4527),
        .dout(new_Jinkela_wire_4528)
    );

    spl4L new_Jinkela_splitter_521 (
        .a(new_Jinkela_wire_4575),
        .d(new_Jinkela_wire_4576),
        .e(new_Jinkela_wire_4577),
        .b(new_Jinkela_wire_4578),
        .c(new_Jinkela_wire_4579)
    );

    bfr new_Jinkela_buffer_3183 (
        .din(new_Jinkela_wire_4544),
        .dout(new_Jinkela_wire_4545)
    );

    bfr new_Jinkela_buffer_3189 (
        .din(new_Jinkela_wire_4550),
        .dout(new_Jinkela_wire_4551)
    );

    bfr new_Jinkela_buffer_3184 (
        .din(new_Jinkela_wire_4545),
        .dout(new_Jinkela_wire_4546)
    );

    spl2 new_Jinkela_splitter_523 (
        .a(_0043_),
        .b(new_Jinkela_wire_4601),
        .c(new_Jinkela_wire_4602)
    );

    bfr new_Jinkela_buffer_3190 (
        .din(new_Jinkela_wire_4551),
        .dout(new_Jinkela_wire_4552)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    spl2 new_Jinkela_splitter_180 (
        .a(G114),
        .b(new_Jinkela_wire_970),
        .c(new_Jinkela_wire_971)
    );

    spl2 new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_960),
        .b(new_Jinkela_wire_961),
        .c(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_500 (
        .din(G81),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_503 (
        .din(G45),
        .dout(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(new_Jinkela_wire_972),
        .b(new_Jinkela_wire_973),
        .c(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    bfr new_Jinkela_buffer_508 (
        .din(G30),
        .dout(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_976),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    bfr new_Jinkela_buffer_3681 (
        .din(new_Jinkela_wire_5151),
        .dout(new_Jinkela_wire_5152)
    );

    bfr new_Jinkela_buffer_4979 (
        .din(new_Jinkela_wire_6786),
        .dout(new_Jinkela_wire_6787)
    );

    bfr new_Jinkela_buffer_3695 (
        .din(new_Jinkela_wire_5167),
        .dout(new_Jinkela_wire_5168)
    );

    bfr new_Jinkela_buffer_4992 (
        .din(new_Jinkela_wire_6805),
        .dout(new_Jinkela_wire_6806)
    );

    bfr new_Jinkela_buffer_3682 (
        .din(new_Jinkela_wire_5152),
        .dout(new_Jinkela_wire_5153)
    );

    bfr new_Jinkela_buffer_4980 (
        .din(new_Jinkela_wire_6787),
        .dout(new_Jinkela_wire_6788)
    );

    bfr new_Jinkela_buffer_3727 (
        .din(new_Jinkela_wire_5201),
        .dout(new_Jinkela_wire_5202)
    );

    bfr new_Jinkela_buffer_4989 (
        .din(new_Jinkela_wire_6802),
        .dout(new_Jinkela_wire_6803)
    );

    bfr new_Jinkela_buffer_3683 (
        .din(new_Jinkela_wire_5153),
        .dout(new_Jinkela_wire_5154)
    );

    bfr new_Jinkela_buffer_4981 (
        .din(new_Jinkela_wire_6788),
        .dout(new_Jinkela_wire_6789)
    );

    bfr new_Jinkela_buffer_3696 (
        .din(new_Jinkela_wire_5168),
        .dout(new_Jinkela_wire_5169)
    );

    bfr new_Jinkela_buffer_3684 (
        .din(new_Jinkela_wire_5154),
        .dout(new_Jinkela_wire_5155)
    );

    spl2 new_Jinkela_splitter_705 (
        .a(_0951_),
        .b(new_Jinkela_wire_6899),
        .c(new_Jinkela_wire_6900)
    );

    bfr new_Jinkela_buffer_3741 (
        .din(_1219_),
        .dout(new_Jinkela_wire_5216)
    );

    bfr new_Jinkela_buffer_4993 (
        .din(new_Jinkela_wire_6806),
        .dout(new_Jinkela_wire_6807)
    );

    bfr new_Jinkela_buffer_5057 (
        .din(new_net_2483),
        .dout(new_Jinkela_wire_6893)
    );

    bfr new_Jinkela_buffer_3697 (
        .din(new_Jinkela_wire_5169),
        .dout(new_Jinkela_wire_5170)
    );

    bfr new_Jinkela_buffer_4994 (
        .din(new_Jinkela_wire_6807),
        .dout(new_Jinkela_wire_6808)
    );

    bfr new_Jinkela_buffer_3728 (
        .din(new_Jinkela_wire_5202),
        .dout(new_Jinkela_wire_5203)
    );

    bfr new_Jinkela_buffer_4996 (
        .din(new_Jinkela_wire_6809),
        .dout(new_Jinkela_wire_6810)
    );

    bfr new_Jinkela_buffer_3698 (
        .din(new_Jinkela_wire_5170),
        .dout(new_Jinkela_wire_5171)
    );

    bfr new_Jinkela_buffer_4995 (
        .din(new_Jinkela_wire_6808),
        .dout(new_Jinkela_wire_6809)
    );

    bfr new_Jinkela_buffer_3739 (
        .din(new_Jinkela_wire_5213),
        .dout(new_Jinkela_wire_5214)
    );

    bfr new_Jinkela_buffer_5020 (
        .din(new_Jinkela_wire_6851),
        .dout(new_Jinkela_wire_6852)
    );

    bfr new_Jinkela_buffer_5058 (
        .din(new_Jinkela_wire_6893),
        .dout(new_Jinkela_wire_6894)
    );

    bfr new_Jinkela_buffer_3699 (
        .din(new_Jinkela_wire_5171),
        .dout(new_Jinkela_wire_5172)
    );

    bfr new_Jinkela_buffer_3729 (
        .din(new_Jinkela_wire_5203),
        .dout(new_Jinkela_wire_5204)
    );

    bfr new_Jinkela_buffer_4997 (
        .din(new_Jinkela_wire_6810),
        .dout(new_Jinkela_wire_6811)
    );

    spl2 new_Jinkela_splitter_710 (
        .a(_0819_),
        .b(new_Jinkela_wire_6934),
        .c(new_Jinkela_wire_6935)
    );

    bfr new_Jinkela_buffer_3700 (
        .din(new_Jinkela_wire_5172),
        .dout(new_Jinkela_wire_5173)
    );

    spl2 new_Jinkela_splitter_706 (
        .a(_0816_),
        .b(new_Jinkela_wire_6901),
        .c(new_Jinkela_wire_6902)
    );

    bfr new_Jinkela_buffer_5021 (
        .din(new_Jinkela_wire_6852),
        .dout(new_Jinkela_wire_6853)
    );

    spl2 new_Jinkela_splitter_560 (
        .a(_0034_),
        .b(new_Jinkela_wire_5217),
        .c(new_Jinkela_wire_5218)
    );

    bfr new_Jinkela_buffer_4998 (
        .din(new_Jinkela_wire_6811),
        .dout(new_Jinkela_wire_6812)
    );

    bfr new_Jinkela_buffer_3742 (
        .din(_0712_),
        .dout(new_Jinkela_wire_5219)
    );

    bfr new_Jinkela_buffer_3701 (
        .din(new_Jinkela_wire_5173),
        .dout(new_Jinkela_wire_5174)
    );

    bfr new_Jinkela_buffer_5022 (
        .din(new_Jinkela_wire_6853),
        .dout(new_Jinkela_wire_6854)
    );

    bfr new_Jinkela_buffer_3730 (
        .din(new_Jinkela_wire_5204),
        .dout(new_Jinkela_wire_5205)
    );

    bfr new_Jinkela_buffer_3702 (
        .din(new_Jinkela_wire_5174),
        .dout(new_Jinkela_wire_5175)
    );

    bfr new_Jinkela_buffer_4999 (
        .din(new_Jinkela_wire_6812),
        .dout(new_Jinkela_wire_6813)
    );

    bfr new_Jinkela_buffer_5059 (
        .din(new_Jinkela_wire_6894),
        .dout(new_Jinkela_wire_6895)
    );

    bfr new_Jinkela_buffer_3740 (
        .din(new_Jinkela_wire_5214),
        .dout(new_Jinkela_wire_5215)
    );

    bfr new_Jinkela_buffer_5000 (
        .din(new_Jinkela_wire_6813),
        .dout(new_Jinkela_wire_6814)
    );

    bfr new_Jinkela_buffer_3703 (
        .din(new_Jinkela_wire_5175),
        .dout(new_Jinkela_wire_5176)
    );

    bfr new_Jinkela_buffer_3731 (
        .din(new_Jinkela_wire_5205),
        .dout(new_Jinkela_wire_5206)
    );

    bfr new_Jinkela_buffer_5023 (
        .din(new_Jinkela_wire_6854),
        .dout(new_Jinkela_wire_6855)
    );

    bfr new_Jinkela_buffer_3704 (
        .din(new_Jinkela_wire_5176),
        .dout(new_Jinkela_wire_5177)
    );

    bfr new_Jinkela_buffer_5001 (
        .din(new_Jinkela_wire_6814),
        .dout(new_Jinkela_wire_6815)
    );

    spl2 new_Jinkela_splitter_562 (
        .a(_0881_),
        .b(new_Jinkela_wire_5236),
        .c(new_Jinkela_wire_5237)
    );

    bfr new_Jinkela_buffer_3743 (
        .din(new_Jinkela_wire_5219),
        .dout(new_Jinkela_wire_5220)
    );

    bfr new_Jinkela_buffer_3705 (
        .din(new_Jinkela_wire_5177),
        .dout(new_Jinkela_wire_5178)
    );

    spl2 new_Jinkela_splitter_694 (
        .a(new_Jinkela_wire_6815),
        .b(new_Jinkela_wire_6816),
        .c(new_Jinkela_wire_6817)
    );

    bfr new_Jinkela_buffer_3732 (
        .din(new_Jinkela_wire_5206),
        .dout(new_Jinkela_wire_5207)
    );

    bfr new_Jinkela_buffer_5002 (
        .din(new_Jinkela_wire_6817),
        .dout(new_Jinkela_wire_6818)
    );

    bfr new_Jinkela_buffer_3706 (
        .din(new_Jinkela_wire_5178),
        .dout(new_Jinkela_wire_5179)
    );

    bfr new_Jinkela_buffer_5024 (
        .din(new_Jinkela_wire_6855),
        .dout(new_Jinkela_wire_6856)
    );

    spl2 new_Jinkela_splitter_707 (
        .a(new_net_22),
        .b(new_Jinkela_wire_6903),
        .c(new_Jinkela_wire_6905)
    );

    bfr new_Jinkela_buffer_3707 (
        .din(new_Jinkela_wire_5179),
        .dout(new_Jinkela_wire_5180)
    );

    spl2 new_Jinkela_splitter_695 (
        .a(new_Jinkela_wire_6818),
        .b(new_Jinkela_wire_6819),
        .c(new_Jinkela_wire_6820)
    );

    bfr new_Jinkela_buffer_3733 (
        .din(new_Jinkela_wire_5207),
        .dout(new_Jinkela_wire_5208)
    );

    bfr new_Jinkela_buffer_5003 (
        .din(new_Jinkela_wire_6820),
        .dout(new_Jinkela_wire_6821)
    );

    bfr new_Jinkela_buffer_3708 (
        .din(new_Jinkela_wire_5180),
        .dout(new_Jinkela_wire_5181)
    );

    bfr new_Jinkela_buffer_5060 (
        .din(new_Jinkela_wire_6895),
        .dout(new_Jinkela_wire_6896)
    );

    bfr new_Jinkela_buffer_5025 (
        .din(new_Jinkela_wire_6856),
        .dout(new_Jinkela_wire_6857)
    );

    spl2 new_Jinkela_splitter_561 (
        .a(_0776_),
        .b(new_Jinkela_wire_5233),
        .c(new_Jinkela_wire_5234)
    );

    bfr new_Jinkela_buffer_3709 (
        .din(new_Jinkela_wire_5181),
        .dout(new_Jinkela_wire_5182)
    );

    bfr new_Jinkela_buffer_5004 (
        .din(new_Jinkela_wire_6821),
        .dout(new_Jinkela_wire_6822)
    );

    bfr new_Jinkela_buffer_3734 (
        .din(new_Jinkela_wire_5208),
        .dout(new_Jinkela_wire_5209)
    );

    bfr new_Jinkela_buffer_5026 (
        .din(new_Jinkela_wire_6857),
        .dout(new_Jinkela_wire_6858)
    );

    bfr new_Jinkela_buffer_3710 (
        .din(new_Jinkela_wire_5182),
        .dout(new_Jinkela_wire_5183)
    );

    spl2 new_Jinkela_splitter_696 (
        .a(new_Jinkela_wire_6822),
        .b(new_Jinkela_wire_6823),
        .c(new_Jinkela_wire_6824)
    );

    bfr new_Jinkela_buffer_3756 (
        .din(new_Jinkela_wire_5234),
        .dout(new_Jinkela_wire_5235)
    );

    bfr new_Jinkela_buffer_5005 (
        .din(new_Jinkela_wire_6824),
        .dout(new_Jinkela_wire_6825)
    );

    bfr new_Jinkela_buffer_3711 (
        .din(new_Jinkela_wire_5183),
        .dout(new_Jinkela_wire_5184)
    );

    spl2 new_Jinkela_splitter_709 (
        .a(_0682_),
        .b(new_Jinkela_wire_6921),
        .c(new_Jinkela_wire_6922)
    );

    bfr new_Jinkela_buffer_3735 (
        .din(new_Jinkela_wire_5209),
        .dout(new_Jinkela_wire_5210)
    );

    bfr new_Jinkela_buffer_5061 (
        .din(new_Jinkela_wire_6896),
        .dout(new_Jinkela_wire_6897)
    );

    bfr new_Jinkela_buffer_5027 (
        .din(new_Jinkela_wire_6858),
        .dout(new_Jinkela_wire_6859)
    );

    bfr new_Jinkela_buffer_3712 (
        .din(new_Jinkela_wire_5184),
        .dout(new_Jinkela_wire_5185)
    );

    bfr new_Jinkela_buffer_5006 (
        .din(new_Jinkela_wire_6825),
        .dout(new_Jinkela_wire_6826)
    );

    bfr new_Jinkela_buffer_3744 (
        .din(new_Jinkela_wire_5220),
        .dout(new_Jinkela_wire_5221)
    );

    bfr new_Jinkela_buffer_3713 (
        .din(new_Jinkela_wire_5185),
        .dout(new_Jinkela_wire_5186)
    );

    spl2 new_Jinkela_splitter_697 (
        .a(new_Jinkela_wire_6826),
        .b(new_Jinkela_wire_6827),
        .c(new_Jinkela_wire_6828)
    );

    bfr new_Jinkela_buffer_3736 (
        .din(new_Jinkela_wire_5210),
        .dout(new_Jinkela_wire_5211)
    );

    bfr new_Jinkela_buffer_5007 (
        .din(new_Jinkela_wire_6828),
        .dout(new_Jinkela_wire_6829)
    );

    and_bb _2327_ (
        .a(new_Jinkela_wire_4053),
        .b(new_Jinkela_wire_374),
        .c(_0337_)
    );

    or_bb _2328_ (
        .a(_0337_),
        .b(new_Jinkela_wire_3971),
        .c(_0338_)
    );

    and_bi _2329_ (
        .a(_0336_),
        .b(new_Jinkela_wire_6757),
        .c(_0339_)
    );

    and_bi _2330_ (
        .a(new_Jinkela_wire_1437),
        .b(new_Jinkela_wire_5813),
        .c(_0340_)
    );

    and_bi _2331_ (
        .a(new_Jinkela_wire_242),
        .b(new_Jinkela_wire_7876),
        .c(_0341_)
    );

    or_bb _2332_ (
        .a(_0341_),
        .b(_0340_),
        .c(_0342_)
    );

    or_bb _2333_ (
        .a(new_Jinkela_wire_7235),
        .b(_0339_),
        .c(new_net_2467)
    );

    or_bi _2334_ (
        .a(new_Jinkela_wire_377),
        .b(new_Jinkela_wire_7939),
        .c(_0343_)
    );

    and_bb _2335_ (
        .a(new_Jinkela_wire_7294),
        .b(new_Jinkela_wire_371),
        .c(_0344_)
    );

    or_bb _2336_ (
        .a(_0344_),
        .b(new_Jinkela_wire_3968),
        .c(_0345_)
    );

    and_bi _2337_ (
        .a(_0343_),
        .b(new_Jinkela_wire_3319),
        .c(_0346_)
    );

    and_bi _2338_ (
        .a(new_Jinkela_wire_151),
        .b(new_Jinkela_wire_7868),
        .c(_0347_)
    );

    and_bi _2339_ (
        .a(new_Jinkela_wire_1194),
        .b(new_Jinkela_wire_5806),
        .c(_0348_)
    );

    or_bb _2340_ (
        .a(_0348_),
        .b(_0347_),
        .c(_0349_)
    );

    or_bb _2341_ (
        .a(new_Jinkela_wire_7288),
        .b(_0346_),
        .c(new_net_2481)
    );

    or_bi _2342_ (
        .a(new_Jinkela_wire_370),
        .b(new_Jinkela_wire_2429),
        .c(_0350_)
    );

    and_bb _2343_ (
        .a(new_Jinkela_wire_7437),
        .b(new_Jinkela_wire_366),
        .c(_0351_)
    );

    or_bb _2344_ (
        .a(_0351_),
        .b(new_Jinkela_wire_3964),
        .c(_0352_)
    );

    and_bi _2345_ (
        .a(_0350_),
        .b(new_Jinkela_wire_4536),
        .c(_0353_)
    );

    and_bi _2346_ (
        .a(new_Jinkela_wire_1248),
        .b(new_Jinkela_wire_5814),
        .c(_0354_)
    );

    and_bi _2347_ (
        .a(new_Jinkela_wire_1611),
        .b(new_Jinkela_wire_7878),
        .c(_0355_)
    );

    or_bb _2348_ (
        .a(_0355_),
        .b(_0354_),
        .c(_0356_)
    );

    or_bb _2349_ (
        .a(new_Jinkela_wire_7370),
        .b(_0353_),
        .c(new_net_2365)
    );

    and_bi _2350_ (
        .a(new_Jinkela_wire_5909),
        .b(new_Jinkela_wire_486),
        .c(_0357_)
    );

    and_bi _2351_ (
        .a(new_Jinkela_wire_2067),
        .b(new_Jinkela_wire_1662),
        .c(_0358_)
    );

    or_bb _2352_ (
        .a(_0358_),
        .b(new_Jinkela_wire_1739),
        .c(_0359_)
    );

    or_bb _2353_ (
        .a(_0359_),
        .b(_0357_),
        .c(_0360_)
    );

    and_bi _2354_ (
        .a(new_Jinkela_wire_1375),
        .b(new_Jinkela_wire_7923),
        .c(_0361_)
    );

    and_bi _2355_ (
        .a(new_Jinkela_wire_506),
        .b(new_Jinkela_wire_6131),
        .c(_0362_)
    );

    or_bb _2356_ (
        .a(_0362_),
        .b(_0361_),
        .c(_0363_)
    );

    and_bi _2357_ (
        .a(_0360_),
        .b(new_Jinkela_wire_3159),
        .c(_0364_)
    );

    and_bi _2358_ (
        .a(new_Jinkela_wire_682),
        .b(_0364_),
        .c(new_net_2461)
    );

    and_bi _2359_ (
        .a(new_Jinkela_wire_2426),
        .b(new_Jinkela_wire_478),
        .c(_0365_)
    );

    and_bi _2360_ (
        .a(new_Jinkela_wire_7434),
        .b(new_Jinkela_wire_1652),
        .c(_0366_)
    );

    or_bb _2361_ (
        .a(_0366_),
        .b(new_Jinkela_wire_1729),
        .c(_0367_)
    );

    or_bb _2362_ (
        .a(new_Jinkela_wire_1968),
        .b(_0365_),
        .c(_0368_)
    );

    and_bi _2363_ (
        .a(new_Jinkela_wire_39),
        .b(new_Jinkela_wire_7918),
        .c(_0369_)
    );

    and_bi _2364_ (
        .a(new_Jinkela_wire_1352),
        .b(new_Jinkela_wire_6136),
        .c(_0370_)
    );

    or_bb _2365_ (
        .a(_0370_),
        .b(_0369_),
        .c(_0371_)
    );

    and_bi _2366_ (
        .a(_0368_),
        .b(new_Jinkela_wire_7265),
        .c(_0372_)
    );

    and_bi _2367_ (
        .a(new_Jinkela_wire_669),
        .b(_0372_),
        .c(new_net_2407)
    );

    and_bi _2368_ (
        .a(new_Jinkela_wire_7940),
        .b(new_Jinkela_wire_484),
        .c(_0373_)
    );

    or_bb _1613_ (
        .a(_0907_),
        .b(new_Jinkela_wire_4826),
        .c(_0908_)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    and_bi _1614_ (
        .a(_0896_),
        .b(new_Jinkela_wire_7391),
        .c(_0909_)
    );

    spl4L new_Jinkela_splitter_144 (
        .a(new_Jinkela_wire_751),
        .d(new_Jinkela_wire_752),
        .e(new_Jinkela_wire_753),
        .b(new_Jinkela_wire_754),
        .c(new_Jinkela_wire_755)
    );

    or_bb _1615_ (
        .a(_0909_),
        .b(new_Jinkela_wire_5155),
        .c(_0910_)
    );

    spl2 new_Jinkela_splitter_130 (
        .a(new_Jinkela_wire_686),
        .b(new_Jinkela_wire_687),
        .c(new_Jinkela_wire_688)
    );

    inv _1616_ (
        .din(new_Jinkela_wire_1616),
        .dout(new_net_2455)
    );

    spl2 new_Jinkela_splitter_131 (
        .a(new_Jinkela_wire_688),
        .b(new_Jinkela_wire_689),
        .c(new_Jinkela_wire_690)
    );

    and_bi _1617_ (
        .a(new_Jinkela_wire_237),
        .b(new_Jinkela_wire_6692),
        .c(_0911_)
    );

    spl2 new_Jinkela_splitter_148 (
        .a(G131),
        .b(new_Jinkela_wire_773),
        .c(new_Jinkela_wire_774)
    );

    and_bi _1618_ (
        .a(new_Jinkela_wire_3371),
        .b(new_Jinkela_wire_3311),
        .c(_0912_)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    or_bi _1619_ (
        .a(new_Jinkela_wire_3370),
        .b(new_Jinkela_wire_3315),
        .c(_0913_)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    and_bi _1620_ (
        .a(_0913_),
        .b(_0912_),
        .c(_0914_)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    or_bb _1621_ (
        .a(new_Jinkela_wire_7713),
        .b(new_Jinkela_wire_1088),
        .c(_0915_)
    );

    spl4L new_Jinkela_splitter_132 (
        .a(new_Jinkela_wire_691),
        .d(new_Jinkela_wire_692),
        .e(new_Jinkela_wire_693),
        .b(new_Jinkela_wire_694),
        .c(new_Jinkela_wire_695)
    );

    or_bb _1622_ (
        .a(new_Jinkela_wire_834),
        .b(new_Jinkela_wire_56),
        .c(_0916_)
    );

    spl4L new_Jinkela_splitter_133 (
        .a(new_Jinkela_wire_695),
        .d(new_Jinkela_wire_696),
        .e(new_Jinkela_wire_697),
        .b(new_Jinkela_wire_698),
        .c(new_Jinkela_wire_699)
    );

    and_bi _1623_ (
        .a(new_Jinkela_wire_831),
        .b(new_Jinkela_wire_413),
        .c(_0917_)
    );

    and_bi _1624_ (
        .a(_0916_),
        .b(_0917_),
        .c(_0918_)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    and_bi _1625_ (
        .a(new_Jinkela_wire_950),
        .b(_0918_),
        .c(_0919_)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    or_ii _1626_ (
        .a(new_Jinkela_wire_833),
        .b(new_Jinkela_wire_1203),
        .c(_0920_)
    );

    spl4L new_Jinkela_splitter_149 (
        .a(G160),
        .d(new_Jinkela_wire_777),
        .e(new_Jinkela_wire_778),
        .b(new_Jinkela_wire_779),
        .c(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    and_bi _1627_ (
        .a(new_Jinkela_wire_1535),
        .b(new_Jinkela_wire_829),
        .c(_0921_)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    and_bi _1628_ (
        .a(_0920_),
        .b(_0921_),
        .c(_0922_)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    or_bb _1629_ (
        .a(_0922_),
        .b(new_Jinkela_wire_949),
        .c(_0923_)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    and_bi _1630_ (
        .a(_0923_),
        .b(_0919_),
        .c(_0924_)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    and_bi _1631_ (
        .a(new_Jinkela_wire_1048),
        .b(new_Jinkela_wire_4707),
        .c(_0925_)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    or_bb _1632_ (
        .a(_0925_),
        .b(new_Jinkela_wire_4836),
        .c(_0926_)
    );

    bfr new_Jinkela_buffer_381 (
        .din(G119),
        .dout(new_Jinkela_wire_825)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    and_bi _1633_ (
        .a(_0915_),
        .b(new_Jinkela_wire_4916),
        .c(_0927_)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(new_Jinkela_wire_762),
        .b(new_Jinkela_wire_763),
        .c(new_Jinkela_wire_764)
    );

    and_ii _1634_ (
        .a(_0927_),
        .b(new_Jinkela_wire_3798),
        .c(new_net_22)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    and_bi _1635_ (
        .a(new_Jinkela_wire_944),
        .b(new_Jinkela_wire_6703),
        .c(_0928_)
    );

    spl4L new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_830),
        .d(new_Jinkela_wire_831),
        .e(new_Jinkela_wire_832),
        .b(new_Jinkela_wire_833),
        .c(new_Jinkela_wire_834)
    );

    or_ii _1636_ (
        .a(new_Jinkela_wire_263),
        .b(new_Jinkela_wire_18),
        .c(_0929_)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_775),
        .dout(new_Jinkela_wire_776)
    );

    and_bi _1637_ (
        .a(new_Jinkela_wire_895),
        .b(new_Jinkela_wire_2),
        .c(_0930_)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_770),
        .dout(new_Jinkela_wire_771)
    );

    and_bi _1638_ (
        .a(new_Jinkela_wire_5825),
        .b(new_Jinkela_wire_1753),
        .c(_0931_)
    );

    spl4L new_Jinkela_splitter_158 (
        .a(new_Jinkela_wire_825),
        .d(new_Jinkela_wire_826),
        .e(new_Jinkela_wire_827),
        .b(new_Jinkela_wire_828),
        .c(new_Jinkela_wire_830)
    );

    and_bi _1639_ (
        .a(new_Jinkela_wire_713),
        .b(new_Jinkela_wire_6498),
        .c(_0932_)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    inv _1640_ (
        .din(new_Jinkela_wire_705),
        .dout(_0933_)
    );

    or_bi _1641_ (
        .a(new_Jinkela_wire_1754),
        .b(new_Jinkela_wire_5826),
        .c(_0934_)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    and_bi _1642_ (
        .a(new_Jinkela_wire_6763),
        .b(new_Jinkela_wire_6191),
        .c(_0935_)
    );

    and_ii _1643_ (
        .a(new_Jinkela_wire_5654),
        .b(new_Jinkela_wire_7501),
        .c(_0936_)
    );

    spl3L new_Jinkela_splitter_160 (
        .a(G159),
        .d(new_Jinkela_wire_835),
        .b(new_Jinkela_wire_836),
        .c(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_838),
        .dout(new_Jinkela_wire_839)
    );

    inv _1644_ (
        .din(new_Jinkela_wire_1299),
        .dout(_0937_)
    );

    bfr new_Jinkela_buffer_388 (
        .din(G120),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    or_ii _1645_ (
        .a(new_Jinkela_wire_24),
        .b(new_Jinkela_wire_1339),
        .c(_0938_)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(G11),
        .b(new_Jinkela_wire_843),
        .c(new_Jinkela_wire_844)
    );

    and_bi _1646_ (
        .a(new_Jinkela_wire_82),
        .b(new_Jinkela_wire_12),
        .c(_0939_)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    and_bi _1647_ (
        .a(_0938_),
        .b(new_Jinkela_wire_4074),
        .c(_0940_)
    );

    or_bb _1648_ (
        .a(new_Jinkela_wire_5049),
        .b(new_Jinkela_wire_2860),
        .c(_0941_)
    );

    spl3L new_Jinkela_splitter_162 (
        .a(G94),
        .d(new_Jinkela_wire_845),
        .b(new_Jinkela_wire_849),
        .c(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    and_bi _1649_ (
        .a(new_Jinkela_wire_5048),
        .b(new_Jinkela_wire_1306),
        .c(_0942_)
    );

    inv _1650_ (
        .din(new_Jinkela_wire_1137),
        .dout(_0943_)
    );

    or_ii _1651_ (
        .a(new_Jinkela_wire_19),
        .b(new_Jinkela_wire_564),
        .c(_0944_)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    and_bi _1652_ (
        .a(new_Jinkela_wire_309),
        .b(new_Jinkela_wire_15),
        .c(_0945_)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    and_bi _1653_ (
        .a(_0944_),
        .b(new_Jinkela_wire_3749),
        .c(_0946_)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_785),
        .dout(new_Jinkela_wire_786)
    );

    or_bb _1654_ (
        .a(new_Jinkela_wire_5126),
        .b(new_Jinkela_wire_3576),
        .c(_0947_)
    );

    bfr new_Jinkela_buffer_383 (
        .din(G19),
        .dout(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_2174 (
        .din(new_Jinkela_wire_3304),
        .dout(new_Jinkela_wire_3305)
    );

    bfr new_Jinkela_buffer_2345 (
        .din(new_Jinkela_wire_3565),
        .dout(new_Jinkela_wire_3566)
    );

    bfr new_Jinkela_buffer_3093 (
        .din(new_Jinkela_wire_4448),
        .dout(new_Jinkela_wire_4449)
    );

    bfr new_Jinkela_buffer_3714 (
        .din(new_Jinkela_wire_5186),
        .dout(new_Jinkela_wire_5187)
    );

    spl2 new_Jinkela_splitter_467 (
        .a(_1074_),
        .b(new_Jinkela_wire_3629),
        .c(new_Jinkela_wire_3630)
    );

    bfr new_Jinkela_buffer_3113 (
        .din(new_Jinkela_wire_4470),
        .dout(new_Jinkela_wire_4471)
    );

    spl2 new_Jinkela_splitter_563 (
        .a(_1215_),
        .b(new_Jinkela_wire_5238),
        .c(new_Jinkela_wire_5239)
    );

    bfr new_Jinkela_buffer_2390 (
        .din(new_Jinkela_wire_3631),
        .dout(new_Jinkela_wire_3632)
    );

    bfr new_Jinkela_buffer_2189 (
        .din(new_Jinkela_wire_3328),
        .dout(new_Jinkela_wire_3329)
    );

    bfr new_Jinkela_buffer_2346 (
        .din(new_Jinkela_wire_3566),
        .dout(new_Jinkela_wire_3567)
    );

    bfr new_Jinkela_buffer_3094 (
        .din(new_Jinkela_wire_4449),
        .dout(new_Jinkela_wire_4450)
    );

    bfr new_Jinkela_buffer_3715 (
        .din(new_Jinkela_wire_5187),
        .dout(new_Jinkela_wire_5188)
    );

    bfr new_Jinkela_buffer_2219 (
        .din(new_Jinkela_wire_3361),
        .dout(new_Jinkela_wire_3362)
    );

    bfr new_Jinkela_buffer_2368 (
        .din(new_Jinkela_wire_3597),
        .dout(new_Jinkela_wire_3598)
    );

    bfr new_Jinkela_buffer_3151 (
        .din(new_Jinkela_wire_4508),
        .dout(new_Jinkela_wire_4509)
    );

    bfr new_Jinkela_buffer_3737 (
        .din(new_Jinkela_wire_5211),
        .dout(new_Jinkela_wire_5212)
    );

    bfr new_Jinkela_buffer_2190 (
        .din(new_Jinkela_wire_3329),
        .dout(new_Jinkela_wire_3330)
    );

    bfr new_Jinkela_buffer_2347 (
        .din(new_Jinkela_wire_3567),
        .dout(new_Jinkela_wire_3568)
    );

    bfr new_Jinkela_buffer_3095 (
        .din(new_Jinkela_wire_4450),
        .dout(new_Jinkela_wire_4451)
    );

    bfr new_Jinkela_buffer_3716 (
        .din(new_Jinkela_wire_5188),
        .dout(new_Jinkela_wire_5189)
    );

    spl2 new_Jinkela_splitter_429 (
        .a(new_Jinkela_wire_3374),
        .b(new_Jinkela_wire_3375),
        .c(new_Jinkela_wire_3376)
    );

    bfr new_Jinkela_buffer_2382 (
        .din(new_Jinkela_wire_3619),
        .dout(new_Jinkela_wire_3620)
    );

    bfr new_Jinkela_buffer_3114 (
        .din(new_Jinkela_wire_4471),
        .dout(new_Jinkela_wire_4472)
    );

    bfr new_Jinkela_buffer_3745 (
        .din(new_Jinkela_wire_5221),
        .dout(new_Jinkela_wire_5222)
    );

    bfr new_Jinkela_buffer_2191 (
        .din(new_Jinkela_wire_3330),
        .dout(new_Jinkela_wire_3331)
    );

    bfr new_Jinkela_buffer_2348 (
        .din(new_Jinkela_wire_3568),
        .dout(new_Jinkela_wire_3569)
    );

    bfr new_Jinkela_buffer_3096 (
        .din(new_Jinkela_wire_4451),
        .dout(new_Jinkela_wire_4452)
    );

    bfr new_Jinkela_buffer_3717 (
        .din(new_Jinkela_wire_5189),
        .dout(new_Jinkela_wire_5190)
    );

    bfr new_Jinkela_buffer_2220 (
        .din(new_Jinkela_wire_3362),
        .dout(new_Jinkela_wire_3363)
    );

    bfr new_Jinkela_buffer_2369 (
        .din(new_Jinkela_wire_3598),
        .dout(new_Jinkela_wire_3599)
    );

    bfr new_Jinkela_buffer_3134 (
        .din(new_Jinkela_wire_4491),
        .dout(new_Jinkela_wire_4492)
    );

    bfr new_Jinkela_buffer_3758 (
        .din(new_Jinkela_wire_5240),
        .dout(new_Jinkela_wire_5241)
    );

    bfr new_Jinkela_buffer_2192 (
        .din(new_Jinkela_wire_3331),
        .dout(new_Jinkela_wire_3332)
    );

    bfr new_Jinkela_buffer_2349 (
        .din(new_Jinkela_wire_3569),
        .dout(new_Jinkela_wire_3570)
    );

    bfr new_Jinkela_buffer_3097 (
        .din(new_Jinkela_wire_4452),
        .dout(new_Jinkela_wire_4453)
    );

    bfr new_Jinkela_buffer_3718 (
        .din(new_Jinkela_wire_5190),
        .dout(new_Jinkela_wire_5191)
    );

    bfr new_Jinkela_buffer_2229 (
        .din(new_Jinkela_wire_3392),
        .dout(new_Jinkela_wire_3393)
    );

    bfr new_Jinkela_buffer_3115 (
        .din(new_Jinkela_wire_4472),
        .dout(new_Jinkela_wire_4473)
    );

    bfr new_Jinkela_buffer_3746 (
        .din(new_Jinkela_wire_5222),
        .dout(new_Jinkela_wire_5223)
    );

    bfr new_Jinkela_buffer_2389 (
        .din(_0560_),
        .dout(new_Jinkela_wire_3631)
    );

    bfr new_Jinkela_buffer_2247 (
        .din(_0611_),
        .dout(new_Jinkela_wire_3411)
    );

    bfr new_Jinkela_buffer_2193 (
        .din(new_Jinkela_wire_3332),
        .dout(new_Jinkela_wire_3333)
    );

    bfr new_Jinkela_buffer_2370 (
        .din(new_Jinkela_wire_3599),
        .dout(new_Jinkela_wire_3600)
    );

    bfr new_Jinkela_buffer_3757 (
        .din(new_net_2449),
        .dout(new_Jinkela_wire_5240)
    );

    bfr new_Jinkela_buffer_3171 (
        .din(new_Jinkela_wire_4532),
        .dout(new_Jinkela_wire_4533)
    );

    bfr new_Jinkela_buffer_2221 (
        .din(new_Jinkela_wire_3363),
        .dout(new_Jinkela_wire_3364)
    );

    bfr new_Jinkela_buffer_3116 (
        .din(new_Jinkela_wire_4473),
        .dout(new_Jinkela_wire_4474)
    );

    bfr new_Jinkela_buffer_3747 (
        .din(new_Jinkela_wire_5223),
        .dout(new_Jinkela_wire_5224)
    );

    bfr new_Jinkela_buffer_2420 (
        .din(_0310_),
        .dout(new_Jinkela_wire_3664)
    );

    bfr new_Jinkela_buffer_2194 (
        .din(new_Jinkela_wire_3333),
        .dout(new_Jinkela_wire_3334)
    );

    bfr new_Jinkela_buffer_2371 (
        .din(new_Jinkela_wire_3600),
        .dout(new_Jinkela_wire_3601)
    );

    bfr new_Jinkela_buffer_3135 (
        .din(new_Jinkela_wire_4492),
        .dout(new_Jinkela_wire_4493)
    );

    spl2 new_Jinkela_splitter_565 (
        .a(_0892_),
        .b(new_Jinkela_wire_5245),
        .c(new_Jinkela_wire_5246)
    );

    spl4L new_Jinkela_splitter_433 (
        .a(new_Jinkela_wire_3385),
        .d(new_Jinkela_wire_3386),
        .e(new_Jinkela_wire_3387),
        .b(new_Jinkela_wire_3388),
        .c(new_Jinkela_wire_3389)
    );

    bfr new_Jinkela_buffer_2383 (
        .din(new_Jinkela_wire_3620),
        .dout(new_Jinkela_wire_3621)
    );

    bfr new_Jinkela_buffer_3117 (
        .din(new_Jinkela_wire_4474),
        .dout(new_Jinkela_wire_4475)
    );

    bfr new_Jinkela_buffer_3748 (
        .din(new_Jinkela_wire_5224),
        .dout(new_Jinkela_wire_5225)
    );

    bfr new_Jinkela_buffer_2195 (
        .din(new_Jinkela_wire_3334),
        .dout(new_Jinkela_wire_3335)
    );

    bfr new_Jinkela_buffer_2372 (
        .din(new_Jinkela_wire_3601),
        .dout(new_Jinkela_wire_3602)
    );

    bfr new_Jinkela_buffer_3152 (
        .din(new_Jinkela_wire_4509),
        .dout(new_Jinkela_wire_4510)
    );

    spl2 new_Jinkela_splitter_564 (
        .a(_0830_),
        .b(new_Jinkela_wire_5243),
        .c(new_Jinkela_wire_5244)
    );

    bfr new_Jinkela_buffer_2222 (
        .din(new_Jinkela_wire_3364),
        .dout(new_Jinkela_wire_3365)
    );

    spl2 new_Jinkela_splitter_468 (
        .a(_1158_),
        .b(new_Jinkela_wire_3662),
        .c(new_Jinkela_wire_3663)
    );

    bfr new_Jinkela_buffer_3118 (
        .din(new_Jinkela_wire_4475),
        .dout(new_Jinkela_wire_4476)
    );

    bfr new_Jinkela_buffer_3749 (
        .din(new_Jinkela_wire_5225),
        .dout(new_Jinkela_wire_5226)
    );

    bfr new_Jinkela_buffer_2196 (
        .din(new_Jinkela_wire_3335),
        .dout(new_Jinkela_wire_3336)
    );

    bfr new_Jinkela_buffer_2373 (
        .din(new_Jinkela_wire_3602),
        .dout(new_Jinkela_wire_3603)
    );

    bfr new_Jinkela_buffer_3136 (
        .din(new_Jinkela_wire_4493),
        .dout(new_Jinkela_wire_4494)
    );

    spl2 new_Jinkela_splitter_436 (
        .a(_0667_),
        .b(new_Jinkela_wire_3416),
        .c(new_Jinkela_wire_3417)
    );

    bfr new_Jinkela_buffer_2384 (
        .din(new_Jinkela_wire_3621),
        .dout(new_Jinkela_wire_3622)
    );

    bfr new_Jinkela_buffer_3119 (
        .din(new_Jinkela_wire_4476),
        .dout(new_Jinkela_wire_4477)
    );

    bfr new_Jinkela_buffer_3750 (
        .din(new_Jinkela_wire_5226),
        .dout(new_Jinkela_wire_5227)
    );

    bfr new_Jinkela_buffer_2197 (
        .din(new_Jinkela_wire_3336),
        .dout(new_Jinkela_wire_3337)
    );

    bfr new_Jinkela_buffer_2374 (
        .din(new_Jinkela_wire_3603),
        .dout(new_Jinkela_wire_3604)
    );

    bfr new_Jinkela_buffer_3759 (
        .din(new_Jinkela_wire_5241),
        .dout(new_Jinkela_wire_5242)
    );

    bfr new_Jinkela_buffer_2223 (
        .din(new_Jinkela_wire_3365),
        .dout(new_Jinkela_wire_3366)
    );

    bfr new_Jinkela_buffer_3120 (
        .din(new_Jinkela_wire_4477),
        .dout(new_Jinkela_wire_4478)
    );

    bfr new_Jinkela_buffer_3751 (
        .din(new_Jinkela_wire_5227),
        .dout(new_Jinkela_wire_5228)
    );

    bfr new_Jinkela_buffer_2433 (
        .din(_0189_),
        .dout(new_Jinkela_wire_3677)
    );

    bfr new_Jinkela_buffer_2198 (
        .din(new_Jinkela_wire_3337),
        .dout(new_Jinkela_wire_3338)
    );

    bfr new_Jinkela_buffer_2375 (
        .din(new_Jinkela_wire_3604),
        .dout(new_Jinkela_wire_3605)
    );

    bfr new_Jinkela_buffer_3137 (
        .din(new_Jinkela_wire_4494),
        .dout(new_Jinkela_wire_4495)
    );

    spl2 new_Jinkela_splitter_431 (
        .a(new_Jinkela_wire_3377),
        .b(new_Jinkela_wire_3378),
        .c(new_Jinkela_wire_3379)
    );

    bfr new_Jinkela_buffer_2385 (
        .din(new_Jinkela_wire_3622),
        .dout(new_Jinkela_wire_3623)
    );

    bfr new_Jinkela_buffer_3121 (
        .din(new_Jinkela_wire_4478),
        .dout(new_Jinkela_wire_4479)
    );

    bfr new_Jinkela_buffer_3752 (
        .din(new_Jinkela_wire_5228),
        .dout(new_Jinkela_wire_5229)
    );

    bfr new_Jinkela_buffer_2199 (
        .din(new_Jinkela_wire_3338),
        .dout(new_Jinkela_wire_3339)
    );

    bfr new_Jinkela_buffer_2376 (
        .din(new_Jinkela_wire_3605),
        .dout(new_Jinkela_wire_3606)
    );

    bfr new_Jinkela_buffer_3153 (
        .din(new_Jinkela_wire_4510),
        .dout(new_Jinkela_wire_4511)
    );

    spl2 new_Jinkela_splitter_566 (
        .a(_1229_),
        .b(new_Jinkela_wire_5247),
        .c(new_Jinkela_wire_5248)
    );

    bfr new_Jinkela_buffer_2224 (
        .din(new_Jinkela_wire_3366),
        .dout(new_Jinkela_wire_3367)
    );

    bfr new_Jinkela_buffer_2391 (
        .din(new_Jinkela_wire_3632),
        .dout(new_Jinkela_wire_3633)
    );

    bfr new_Jinkela_buffer_3122 (
        .din(new_Jinkela_wire_4479),
        .dout(new_Jinkela_wire_4480)
    );

    bfr new_Jinkela_buffer_3753 (
        .din(new_Jinkela_wire_5229),
        .dout(new_Jinkela_wire_5230)
    );

    bfr new_Jinkela_buffer_2200 (
        .din(new_Jinkela_wire_3339),
        .dout(new_Jinkela_wire_3340)
    );

    bfr new_Jinkela_buffer_2377 (
        .din(new_Jinkela_wire_3606),
        .dout(new_Jinkela_wire_3607)
    );

    bfr new_Jinkela_buffer_3138 (
        .din(new_Jinkela_wire_4495),
        .dout(new_Jinkela_wire_4496)
    );

    bfr new_Jinkela_buffer_3761 (
        .din(_0967_),
        .dout(new_Jinkela_wire_5250)
    );

    bfr new_Jinkela_buffer_3760 (
        .din(new_Jinkela_wire_5248),
        .dout(new_Jinkela_wire_5249)
    );

    bfr new_Jinkela_buffer_2386 (
        .din(new_Jinkela_wire_3623),
        .dout(new_Jinkela_wire_3624)
    );

    bfr new_Jinkela_buffer_3123 (
        .din(new_Jinkela_wire_4480),
        .dout(new_Jinkela_wire_4481)
    );

    bfr new_Jinkela_buffer_3754 (
        .din(new_Jinkela_wire_5230),
        .dout(new_Jinkela_wire_5231)
    );

    bfr new_Jinkela_buffer_2228 (
        .din(_1044_),
        .dout(new_Jinkela_wire_3392)
    );

    bfr new_Jinkela_buffer_2201 (
        .din(new_Jinkela_wire_3340),
        .dout(new_Jinkela_wire_3341)
    );

    bfr new_Jinkela_buffer_2378 (
        .din(new_Jinkela_wire_3607),
        .dout(new_Jinkela_wire_3608)
    );

    bfr new_Jinkela_buffer_3174 (
        .din(new_Jinkela_wire_4535),
        .dout(new_Jinkela_wire_4536)
    );

    spl2 new_Jinkela_splitter_570 (
        .a(_0669_),
        .b(new_Jinkela_wire_5273),
        .c(new_Jinkela_wire_5274)
    );

    bfr new_Jinkela_buffer_3175 (
        .din(_0084_),
        .dout(new_Jinkela_wire_4537)
    );

    bfr new_Jinkela_buffer_2225 (
        .din(new_Jinkela_wire_3367),
        .dout(new_Jinkela_wire_3368)
    );

    bfr new_Jinkela_buffer_3124 (
        .din(new_Jinkela_wire_4481),
        .dout(new_Jinkela_wire_4482)
    );

    bfr new_Jinkela_buffer_3755 (
        .din(new_Jinkela_wire_5231),
        .dout(new_Jinkela_wire_5232)
    );

    bfr new_Jinkela_buffer_2202 (
        .din(new_Jinkela_wire_3341),
        .dout(new_Jinkela_wire_3342)
    );

    bfr new_Jinkela_buffer_2379 (
        .din(new_Jinkela_wire_3608),
        .dout(new_Jinkela_wire_3609)
    );

    bfr new_Jinkela_buffer_3139 (
        .din(new_Jinkela_wire_4496),
        .dout(new_Jinkela_wire_4497)
    );

    bfr new_Jinkela_buffer_3778 (
        .din(new_Jinkela_wire_5275),
        .dout(new_Jinkela_wire_5276)
    );

    spl2 new_Jinkela_splitter_567 (
        .a(new_Jinkela_wire_5250),
        .b(new_Jinkela_wire_5251),
        .c(new_Jinkela_wire_5252)
    );

    bfr new_Jinkela_buffer_2387 (
        .din(new_Jinkela_wire_3624),
        .dout(new_Jinkela_wire_3625)
    );

    bfr new_Jinkela_buffer_3125 (
        .din(new_Jinkela_wire_4482),
        .dout(new_Jinkela_wire_4483)
    );

    bfr new_Jinkela_buffer_3762 (
        .din(new_Jinkela_wire_5252),
        .dout(new_Jinkela_wire_5253)
    );

    spl2 new_Jinkela_splitter_569 (
        .a(_0798_),
        .b(new_Jinkela_wire_5271),
        .c(new_Jinkela_wire_5272)
    );

    spl4L new_Jinkela_splitter_435 (
        .a(_1226_),
        .d(new_Jinkela_wire_3412),
        .e(new_Jinkela_wire_3413),
        .b(new_Jinkela_wire_3414),
        .c(new_Jinkela_wire_3415)
    );

    bfr new_Jinkela_buffer_2203 (
        .din(new_Jinkela_wire_3342),
        .dout(new_Jinkela_wire_3343)
    );

    bfr new_Jinkela_buffer_2392 (
        .din(new_Jinkela_wire_3633),
        .dout(new_Jinkela_wire_3634)
    );

    bfr new_Jinkela_buffer_3154 (
        .din(new_Jinkela_wire_4511),
        .dout(new_Jinkela_wire_4512)
    );

    bfr new_Jinkela_buffer_2226 (
        .din(new_Jinkela_wire_3368),
        .dout(new_Jinkela_wire_3369)
    );

    bfr new_Jinkela_buffer_2388 (
        .din(new_Jinkela_wire_3625),
        .dout(new_Jinkela_wire_3626)
    );

    bfr new_Jinkela_buffer_3126 (
        .din(new_Jinkela_wire_4483),
        .dout(new_Jinkela_wire_4484)
    );

    bfr new_Jinkela_buffer_3784 (
        .din(_0608_),
        .dout(new_Jinkela_wire_5285)
    );

    bfr new_Jinkela_buffer_3777 (
        .din(new_Jinkela_wire_5274),
        .dout(new_Jinkela_wire_5275)
    );

    bfr new_Jinkela_buffer_2204 (
        .din(new_Jinkela_wire_3343),
        .dout(new_Jinkela_wire_3344)
    );

    bfr new_Jinkela_buffer_2421 (
        .din(new_net_2383),
        .dout(new_Jinkela_wire_3665)
    );

    bfr new_Jinkela_buffer_3140 (
        .din(new_Jinkela_wire_4497),
        .dout(new_Jinkela_wire_4498)
    );

    bfr new_Jinkela_buffer_2434 (
        .din(new_net_2443),
        .dout(new_Jinkela_wire_3680)
    );

    bfr new_Jinkela_buffer_2230 (
        .din(new_Jinkela_wire_3393),
        .dout(new_Jinkela_wire_3394)
    );

    bfr new_Jinkela_buffer_2393 (
        .din(new_Jinkela_wire_3634),
        .dout(new_Jinkela_wire_3635)
    );

    bfr new_Jinkela_buffer_3127 (
        .din(new_Jinkela_wire_4484),
        .dout(new_Jinkela_wire_4485)
    );

    spl3L new_Jinkela_splitter_568 (
        .a(new_Jinkela_wire_5253),
        .d(new_Jinkela_wire_5254),
        .b(new_Jinkela_wire_5255),
        .c(new_Jinkela_wire_5256)
    );

    bfr new_Jinkela_buffer_2205 (
        .din(new_Jinkela_wire_3344),
        .dout(new_Jinkela_wire_3345)
    );

    bfr new_Jinkela_buffer_2422 (
        .din(new_Jinkela_wire_3665),
        .dout(new_Jinkela_wire_3666)
    );

    bfr new_Jinkela_buffer_3172 (
        .din(new_Jinkela_wire_4533),
        .dout(new_Jinkela_wire_4534)
    );

    spl2 new_Jinkela_splitter_427 (
        .a(new_Jinkela_wire_3369),
        .b(new_Jinkela_wire_3370),
        .c(new_Jinkela_wire_3371)
    );

    bfr new_Jinkela_buffer_2394 (
        .din(new_Jinkela_wire_3635),
        .dout(new_Jinkela_wire_3636)
    );

    bfr new_Jinkela_buffer_3128 (
        .din(new_Jinkela_wire_4485),
        .dout(new_Jinkela_wire_4486)
    );

    bfr new_Jinkela_buffer_3763 (
        .din(new_Jinkela_wire_5256),
        .dout(new_Jinkela_wire_5257)
    );

    bfr new_Jinkela_buffer_2206 (
        .din(new_Jinkela_wire_3345),
        .dout(new_Jinkela_wire_3346)
    );

    spl2 new_Jinkela_splitter_470 (
        .a(_1057_),
        .b(new_Jinkela_wire_3714),
        .c(new_Jinkela_wire_3715)
    );

    bfr new_Jinkela_buffer_3141 (
        .din(new_Jinkela_wire_4498),
        .dout(new_Jinkela_wire_4499)
    );

    spl3L new_Jinkela_splitter_572 (
        .a(_0864_),
        .d(new_Jinkela_wire_5296),
        .b(new_Jinkela_wire_5297),
        .c(new_Jinkela_wire_5298)
    );

    bfr new_Jinkela_buffer_3783 (
        .din(_0585_),
        .dout(new_Jinkela_wire_5284)
    );

    bfr new_Jinkela_buffer_2231 (
        .din(new_Jinkela_wire_3394),
        .dout(new_Jinkela_wire_3395)
    );

    bfr new_Jinkela_buffer_2395 (
        .din(new_Jinkela_wire_3636),
        .dout(new_Jinkela_wire_3637)
    );

    bfr new_Jinkela_buffer_3129 (
        .din(new_Jinkela_wire_4486),
        .dout(new_Jinkela_wire_4487)
    );

    bfr new_Jinkela_buffer_3764 (
        .din(new_Jinkela_wire_5257),
        .dout(new_Jinkela_wire_5258)
    );

    bfr new_Jinkela_buffer_2207 (
        .din(new_Jinkela_wire_3346),
        .dout(new_Jinkela_wire_3347)
    );

    bfr new_Jinkela_buffer_2423 (
        .din(new_Jinkela_wire_3666),
        .dout(new_Jinkela_wire_3667)
    );

    bfr new_Jinkela_buffer_3155 (
        .din(new_Jinkela_wire_4512),
        .dout(new_Jinkela_wire_4513)
    );

    spl2 new_Jinkela_splitter_573 (
        .a(_0073_),
        .b(new_Jinkela_wire_5300),
        .c(new_Jinkela_wire_5301)
    );

    bfr new_Jinkela_buffer_2396 (
        .din(new_Jinkela_wire_3637),
        .dout(new_Jinkela_wire_3638)
    );

    bfr new_Jinkela_buffer_3130 (
        .din(new_Jinkela_wire_4487),
        .dout(new_Jinkela_wire_4488)
    );

    bfr new_Jinkela_buffer_3765 (
        .din(new_Jinkela_wire_5258),
        .dout(new_Jinkela_wire_5259)
    );

    bfr new_Jinkela_buffer_2250 (
        .din(_0250_),
        .dout(new_Jinkela_wire_3420)
    );

    bfr new_Jinkela_buffer_2208 (
        .din(new_Jinkela_wire_3347),
        .dout(new_Jinkela_wire_3348)
    );

    spl2 new_Jinkela_splitter_469 (
        .a(new_Jinkela_wire_3677),
        .b(new_Jinkela_wire_3678),
        .c(new_Jinkela_wire_3679)
    );

    bfr new_Jinkela_buffer_3142 (
        .din(new_Jinkela_wire_4499),
        .dout(new_Jinkela_wire_4500)
    );

    bfr new_Jinkela_buffer_3785 (
        .din(new_Jinkela_wire_5285),
        .dout(new_Jinkela_wire_5286)
    );

    bfr new_Jinkela_buffer_2397 (
        .din(new_Jinkela_wire_3638),
        .dout(new_Jinkela_wire_3639)
    );

    bfr new_Jinkela_buffer_3766 (
        .din(new_Jinkela_wire_5259),
        .dout(new_Jinkela_wire_5260)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_2360),
        .dout(new_Jinkela_wire_2361)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(new_Jinkela_wire_2341),
        .dout(new_Jinkela_wire_2342)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(new_Jinkela_wire_2399),
        .dout(new_Jinkela_wire_2400)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(new_Jinkela_wire_2342),
        .dout(new_Jinkela_wire_2343)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_2361),
        .dout(new_Jinkela_wire_2362)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_2343),
        .dout(new_Jinkela_wire_2344)
    );

    spl2 new_Jinkela_splitter_368 (
        .a(_1042_),
        .b(new_Jinkela_wire_2413),
        .c(new_Jinkela_wire_2414)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(new_Jinkela_wire_2344),
        .dout(new_Jinkela_wire_2345)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_2362),
        .dout(new_Jinkela_wire_2363)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(new_Jinkela_wire_2345),
        .dout(new_Jinkela_wire_2346)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(new_Jinkela_wire_2400),
        .dout(new_Jinkela_wire_2401)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(new_Jinkela_wire_2346),
        .dout(new_Jinkela_wire_2347)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_2363),
        .dout(new_Jinkela_wire_2364)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_Jinkela_wire_2347),
        .dout(new_Jinkela_wire_2348)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(_1101_),
        .dout(new_Jinkela_wire_2409)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_2348),
        .dout(new_Jinkela_wire_2349)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_2364),
        .dout(new_Jinkela_wire_2365)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_2349),
        .dout(new_Jinkela_wire_2350)
    );

    spl2 new_Jinkela_splitter_364 (
        .a(new_Jinkela_wire_2401),
        .b(new_Jinkela_wire_2402),
        .c(new_Jinkela_wire_2403)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(new_Jinkela_wire_2350),
        .dout(new_Jinkela_wire_2351)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(new_Jinkela_wire_2365),
        .dout(new_Jinkela_wire_2366)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_2351),
        .dout(new_Jinkela_wire_2352)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_2352),
        .dout(new_Jinkela_wire_2353)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_2366),
        .dout(new_Jinkela_wire_2367)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_2353),
        .dout(new_Jinkela_wire_2354)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(new_Jinkela_wire_2409),
        .dout(new_Jinkela_wire_2410)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_2354),
        .dout(new_Jinkela_wire_2355)
    );

    spl4L new_Jinkela_splitter_369 (
        .a(_0855_),
        .d(new_Jinkela_wire_2417),
        .e(new_Jinkela_wire_2418),
        .b(new_Jinkela_wire_2419),
        .c(new_Jinkela_wire_2420)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_2367),
        .dout(new_Jinkela_wire_2368)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_2368),
        .dout(new_Jinkela_wire_2369)
    );

    spl2 new_Jinkela_splitter_367 (
        .a(new_Jinkela_wire_2410),
        .b(new_Jinkela_wire_2411),
        .c(new_Jinkela_wire_2412)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_2369),
        .dout(new_Jinkela_wire_2370)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_2421),
        .dout(new_Jinkela_wire_2422)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_2370),
        .dout(new_Jinkela_wire_2371)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(new_Jinkela_wire_2414),
        .dout(new_Jinkela_wire_2415)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(_0216_),
        .dout(new_Jinkela_wire_2421)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_2371),
        .dout(new_Jinkela_wire_2372)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_2415),
        .dout(new_Jinkela_wire_2416)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_2372),
        .dout(new_Jinkela_wire_2373)
    );

    spl2 new_Jinkela_splitter_371 (
        .a(new_net_11),
        .b(new_Jinkela_wire_2425),
        .c(new_Jinkela_wire_2427)
    );

    spl2 new_Jinkela_splitter_370 (
        .a(_1212_),
        .b(new_Jinkela_wire_2423),
        .c(new_Jinkela_wire_2424)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_2373),
        .dout(new_Jinkela_wire_2374)
    );

    bfr new_Jinkela_buffer_3052 (
        .din(new_Jinkela_wire_4403),
        .dout(new_Jinkela_wire_4404)
    );

    bfr new_Jinkela_buffer_3076 (
        .din(new_Jinkela_wire_4431),
        .dout(new_Jinkela_wire_4432)
    );

    bfr new_Jinkela_buffer_3053 (
        .din(new_Jinkela_wire_4404),
        .dout(new_Jinkela_wire_4405)
    );

    bfr new_Jinkela_buffer_3100 (
        .din(new_Jinkela_wire_4455),
        .dout(new_Jinkela_wire_4456)
    );

    bfr new_Jinkela_buffer_3054 (
        .din(new_Jinkela_wire_4405),
        .dout(new_Jinkela_wire_4406)
    );

    bfr new_Jinkela_buffer_3077 (
        .din(new_Jinkela_wire_4432),
        .dout(new_Jinkela_wire_4433)
    );

    bfr new_Jinkela_buffer_3055 (
        .din(new_Jinkela_wire_4406),
        .dout(new_Jinkela_wire_4407)
    );

    bfr new_Jinkela_buffer_3109 (
        .din(new_Jinkela_wire_4466),
        .dout(new_Jinkela_wire_4467)
    );

    bfr new_Jinkela_buffer_3056 (
        .din(new_Jinkela_wire_4407),
        .dout(new_Jinkela_wire_4408)
    );

    bfr new_Jinkela_buffer_3078 (
        .din(new_Jinkela_wire_4433),
        .dout(new_Jinkela_wire_4434)
    );

    bfr new_Jinkela_buffer_3057 (
        .din(new_Jinkela_wire_4408),
        .dout(new_Jinkela_wire_4409)
    );

    bfr new_Jinkela_buffer_3101 (
        .din(new_Jinkela_wire_4456),
        .dout(new_Jinkela_wire_4457)
    );

    bfr new_Jinkela_buffer_3058 (
        .din(new_Jinkela_wire_4409),
        .dout(new_Jinkela_wire_4410)
    );

    bfr new_Jinkela_buffer_3079 (
        .din(new_Jinkela_wire_4434),
        .dout(new_Jinkela_wire_4435)
    );

    bfr new_Jinkela_buffer_3131 (
        .din(new_net_2427),
        .dout(new_Jinkela_wire_4489)
    );

    bfr new_Jinkela_buffer_3080 (
        .din(new_Jinkela_wire_4435),
        .dout(new_Jinkela_wire_4436)
    );

    bfr new_Jinkela_buffer_3102 (
        .din(new_Jinkela_wire_4457),
        .dout(new_Jinkela_wire_4458)
    );

    bfr new_Jinkela_buffer_3081 (
        .din(new_Jinkela_wire_4436),
        .dout(new_Jinkela_wire_4437)
    );

    bfr new_Jinkela_buffer_3150 (
        .din(_1006_),
        .dout(new_Jinkela_wire_4508)
    );

    bfr new_Jinkela_buffer_3082 (
        .din(new_Jinkela_wire_4437),
        .dout(new_Jinkela_wire_4438)
    );

    bfr new_Jinkela_buffer_3103 (
        .din(new_Jinkela_wire_4458),
        .dout(new_Jinkela_wire_4459)
    );

    bfr new_Jinkela_buffer_3083 (
        .din(new_Jinkela_wire_4438),
        .dout(new_Jinkela_wire_4439)
    );

    bfr new_Jinkela_buffer_3110 (
        .din(new_Jinkela_wire_4467),
        .dout(new_Jinkela_wire_4468)
    );

    bfr new_Jinkela_buffer_3084 (
        .din(new_Jinkela_wire_4439),
        .dout(new_Jinkela_wire_4440)
    );

    bfr new_Jinkela_buffer_3104 (
        .din(new_Jinkela_wire_4459),
        .dout(new_Jinkela_wire_4460)
    );

    bfr new_Jinkela_buffer_3085 (
        .din(new_Jinkela_wire_4440),
        .dout(new_Jinkela_wire_4441)
    );

    bfr new_Jinkela_buffer_3132 (
        .din(new_Jinkela_wire_4489),
        .dout(new_Jinkela_wire_4490)
    );

    bfr new_Jinkela_buffer_3086 (
        .din(new_Jinkela_wire_4441),
        .dout(new_Jinkela_wire_4442)
    );

    bfr new_Jinkela_buffer_3105 (
        .din(new_Jinkela_wire_4460),
        .dout(new_Jinkela_wire_4461)
    );

    bfr new_Jinkela_buffer_3087 (
        .din(new_Jinkela_wire_4442),
        .dout(new_Jinkela_wire_4443)
    );

    bfr new_Jinkela_buffer_3111 (
        .din(new_Jinkela_wire_4468),
        .dout(new_Jinkela_wire_4469)
    );

    bfr new_Jinkela_buffer_3088 (
        .din(new_Jinkela_wire_4443),
        .dout(new_Jinkela_wire_4444)
    );

    bfr new_Jinkela_buffer_3106 (
        .din(new_Jinkela_wire_4461),
        .dout(new_Jinkela_wire_4462)
    );

    bfr new_Jinkela_buffer_3089 (
        .din(new_Jinkela_wire_4444),
        .dout(new_Jinkela_wire_4445)
    );

    spl4L new_Jinkela_splitter_517 (
        .a(_0615_),
        .d(new_Jinkela_wire_4529),
        .e(new_Jinkela_wire_4530),
        .b(new_Jinkela_wire_4531),
        .c(new_Jinkela_wire_4532)
    );

    bfr new_Jinkela_buffer_3173 (
        .din(_0352_),
        .dout(new_Jinkela_wire_4535)
    );

    bfr new_Jinkela_buffer_3090 (
        .din(new_Jinkela_wire_4445),
        .dout(new_Jinkela_wire_4446)
    );

    bfr new_Jinkela_buffer_3107 (
        .din(new_Jinkela_wire_4462),
        .dout(new_Jinkela_wire_4463)
    );

    bfr new_Jinkela_buffer_3091 (
        .din(new_Jinkela_wire_4446),
        .dout(new_Jinkela_wire_4447)
    );

    bfr new_Jinkela_buffer_3112 (
        .din(new_Jinkela_wire_4469),
        .dout(new_Jinkela_wire_4470)
    );

    bfr new_Jinkela_buffer_3092 (
        .din(new_Jinkela_wire_4447),
        .dout(new_Jinkela_wire_4448)
    );

    bfr new_Jinkela_buffer_3133 (
        .din(new_Jinkela_wire_4490),
        .dout(new_Jinkela_wire_4491)
    );

    and_bi _1655_ (
        .a(new_Jinkela_wire_5128),
        .b(new_Jinkela_wire_1145),
        .c(_0948_)
    );

    and_bi _2369_ (
        .a(new_Jinkela_wire_7290),
        .b(new_Jinkela_wire_1656),
        .c(_0374_)
    );

    bfr new_Jinkela_buffer_2424 (
        .din(new_Jinkela_wire_3667),
        .dout(new_Jinkela_wire_3668)
    );

    inv _1656_ (
        .din(new_Jinkela_wire_531),
        .dout(_0949_)
    );

    or_bb _2370_ (
        .a(_0374_),
        .b(new_Jinkela_wire_1733),
        .c(_0375_)
    );

    bfr new_Jinkela_buffer_2398 (
        .din(new_Jinkela_wire_3639),
        .dout(new_Jinkela_wire_3640)
    );

    or_ii _1657_ (
        .a(new_Jinkela_wire_14),
        .b(new_Jinkela_wire_848),
        .c(_0950_)
    );

    or_bb _2371_ (
        .a(new_Jinkela_wire_1982),
        .b(_0373_),
        .c(_0376_)
    );

    and_bi _1658_ (
        .a(new_Jinkela_wire_969),
        .b(new_Jinkela_wire_4),
        .c(_0951_)
    );

    and_bi _2372_ (
        .a(new_Jinkela_wire_1218),
        .b(new_Jinkela_wire_7924),
        .c(_0377_)
    );

    bfr new_Jinkela_buffer_2399 (
        .din(new_Jinkela_wire_3640),
        .dout(new_Jinkela_wire_3641)
    );

    and_bi _1659_ (
        .a(new_Jinkela_wire_2244),
        .b(new_Jinkela_wire_6899),
        .c(_0952_)
    );

    and_bi _2373_ (
        .a(new_Jinkela_wire_1525),
        .b(new_Jinkela_wire_6126),
        .c(_0378_)
    );

    bfr new_Jinkela_buffer_2425 (
        .din(new_Jinkela_wire_3668),
        .dout(new_Jinkela_wire_3669)
    );

    or_bb _1660_ (
        .a(new_Jinkela_wire_7470),
        .b(new_Jinkela_wire_3776),
        .c(_0953_)
    );

    or_bb _2374_ (
        .a(_0378_),
        .b(_0377_),
        .c(_0379_)
    );

    bfr new_Jinkela_buffer_2400 (
        .din(new_Jinkela_wire_3641),
        .dout(new_Jinkela_wire_3642)
    );

    and_ii _1661_ (
        .a(new_Jinkela_wire_2905),
        .b(new_Jinkela_wire_6380),
        .c(_0954_)
    );

    and_bi _2375_ (
        .a(_0376_),
        .b(new_Jinkela_wire_2840),
        .c(_0380_)
    );

    bfr new_Jinkela_buffer_2499 (
        .din(_0945_),
        .dout(new_Jinkela_wire_3749)
    );

    bfr new_Jinkela_buffer_2468 (
        .din(_0544_),
        .dout(new_Jinkela_wire_3716)
    );

    and_bi _1662_ (
        .a(new_Jinkela_wire_3093),
        .b(new_Jinkela_wire_6065),
        .c(_0955_)
    );

    and_bi _2376_ (
        .a(new_Jinkela_wire_675),
        .b(_0380_),
        .c(new_net_2413)
    );

    bfr new_Jinkela_buffer_2401 (
        .din(new_Jinkela_wire_3642),
        .dout(new_Jinkela_wire_3643)
    );

    and_ii _1663_ (
        .a(new_Jinkela_wire_6101),
        .b(new_Jinkela_wire_7600),
        .c(_0956_)
    );

    and_bi _2377_ (
        .a(new_Jinkela_wire_5882),
        .b(new_Jinkela_wire_483),
        .c(_0381_)
    );

    bfr new_Jinkela_buffer_2426 (
        .din(new_Jinkela_wire_3669),
        .dout(new_Jinkela_wire_3670)
    );

    and_bi _1664_ (
        .a(new_Jinkela_wire_6242),
        .b(new_Jinkela_wire_7204),
        .c(_0957_)
    );

    and_bi _2378_ (
        .a(new_Jinkela_wire_4055),
        .b(new_Jinkela_wire_1659),
        .c(_0382_)
    );

    bfr new_Jinkela_buffer_2402 (
        .din(new_Jinkela_wire_3643),
        .dout(new_Jinkela_wire_3644)
    );

    or_bb _1665_ (
        .a(new_Jinkela_wire_3251),
        .b(new_Jinkela_wire_2846),
        .c(_0958_)
    );

    or_bb _2379_ (
        .a(_0382_),
        .b(new_Jinkela_wire_1736),
        .c(_0383_)
    );

    bfr new_Jinkela_buffer_2435 (
        .din(new_Jinkela_wire_3680),
        .dout(new_Jinkela_wire_3681)
    );

    bfr new_Jinkela_buffer_2469 (
        .din(new_Jinkela_wire_3716),
        .dout(new_Jinkela_wire_3717)
    );

    and_ii _1666_ (
        .a(new_Jinkela_wire_3525),
        .b(new_Jinkela_wire_3538),
        .c(_0959_)
    );

    or_bb _2380_ (
        .a(new_Jinkela_wire_2862),
        .b(_0381_),
        .c(_0384_)
    );

    bfr new_Jinkela_buffer_2403 (
        .din(new_Jinkela_wire_3644),
        .dout(new_Jinkela_wire_3645)
    );

    and_bi _1667_ (
        .a(new_Jinkela_wire_3193),
        .b(new_Jinkela_wire_4309),
        .c(_0960_)
    );

    and_bi _2381_ (
        .a(new_Jinkela_wire_519),
        .b(new_Jinkela_wire_7919),
        .c(_0385_)
    );

    bfr new_Jinkela_buffer_2427 (
        .din(new_Jinkela_wire_3670),
        .dout(new_Jinkela_wire_3671)
    );

    or_bb _1668_ (
        .a(_0960_),
        .b(new_Jinkela_wire_3612),
        .c(_0961_)
    );

    and_bi _2382_ (
        .a(new_Jinkela_wire_717),
        .b(new_Jinkela_wire_6127),
        .c(_0386_)
    );

    bfr new_Jinkela_buffer_2404 (
        .din(new_Jinkela_wire_3645),
        .dout(new_Jinkela_wire_3646)
    );

    or_bb _1669_ (
        .a(new_Jinkela_wire_7151),
        .b(_0959_),
        .c(_0962_)
    );

    or_bb _2383_ (
        .a(_0386_),
        .b(_0385_),
        .c(_0387_)
    );

    bfr new_Jinkela_buffer_2436 (
        .din(new_Jinkela_wire_3681),
        .dout(new_Jinkela_wire_3682)
    );

    and_ii _1670_ (
        .a(new_Jinkela_wire_1911),
        .b(new_Jinkela_wire_5115),
        .c(_0963_)
    );

    and_bi _2384_ (
        .a(_0384_),
        .b(new_Jinkela_wire_4488),
        .c(_0388_)
    );

    bfr new_Jinkela_buffer_2405 (
        .din(new_Jinkela_wire_3646),
        .dout(new_Jinkela_wire_3647)
    );

    and_bi _1671_ (
        .a(new_Jinkela_wire_6234),
        .b(new_Jinkela_wire_7595),
        .c(_0964_)
    );

    and_bi _2385_ (
        .a(new_Jinkela_wire_679),
        .b(_0388_),
        .c(new_net_2387)
    );

    bfr new_Jinkela_buffer_2428 (
        .din(new_Jinkela_wire_3671),
        .dout(new_Jinkela_wire_3672)
    );

    and_bi _1672_ (
        .a(new_Jinkela_wire_3090),
        .b(new_Jinkela_wire_6381),
        .c(_0965_)
    );

    and_bi _2386_ (
        .a(new_Jinkela_wire_5912),
        .b(new_Jinkela_wire_811),
        .c(_0389_)
    );

    bfr new_Jinkela_buffer_2406 (
        .din(new_Jinkela_wire_3647),
        .dout(new_Jinkela_wire_3648)
    );

    or_bi _1673_ (
        .a(new_Jinkela_wire_6900),
        .b(new_Jinkela_wire_2245),
        .c(_0966_)
    );

    and_bi _2387_ (
        .a(new_Jinkela_wire_2069),
        .b(new_Jinkela_wire_6833),
        .c(_0390_)
    );

    or_bb _1674_ (
        .a(_0966_),
        .b(new_Jinkela_wire_537),
        .c(_0967_)
    );

    or_bb _2388_ (
        .a(_0390_),
        .b(new_Jinkela_wire_5584),
        .c(_0391_)
    );

    bfr new_Jinkela_buffer_2407 (
        .din(new_Jinkela_wire_3648),
        .dout(new_Jinkela_wire_3649)
    );

    or_ii _1675_ (
        .a(new_Jinkela_wire_5251),
        .b(new_Jinkela_wire_2904),
        .c(_0968_)
    );

    or_bb _2389_ (
        .a(_0391_),
        .b(_0389_),
        .c(_0392_)
    );

    bfr new_Jinkela_buffer_2429 (
        .din(new_Jinkela_wire_3672),
        .dout(new_Jinkela_wire_3673)
    );

    and_bi _1676_ (
        .a(new_Jinkela_wire_7016),
        .b(new_Jinkela_wire_2246),
        .c(_0969_)
    );

    and_bi _2390_ (
        .a(new_Jinkela_wire_1376),
        .b(new_Jinkela_wire_3387),
        .c(_0393_)
    );

    bfr new_Jinkela_buffer_2408 (
        .din(new_Jinkela_wire_3649),
        .dout(new_Jinkela_wire_3650)
    );

    or_ii _1677_ (
        .a(new_Jinkela_wire_1890),
        .b(new_Jinkela_wire_6047),
        .c(_0970_)
    );

    and_bi _2391_ (
        .a(new_Jinkela_wire_507),
        .b(new_Jinkela_wire_4031),
        .c(_0394_)
    );

    bfr new_Jinkela_buffer_2437 (
        .din(new_Jinkela_wire_3682),
        .dout(new_Jinkela_wire_3683)
    );

    and_ii _1678_ (
        .a(new_Jinkela_wire_6948),
        .b(new_Jinkela_wire_1630),
        .c(_0971_)
    );

    or_bb _2392_ (
        .a(_0394_),
        .b(_0393_),
        .c(_0395_)
    );

    bfr new_Jinkela_buffer_2409 (
        .din(new_Jinkela_wire_3650),
        .dout(new_Jinkela_wire_3651)
    );

    and_bi _1679_ (
        .a(new_Jinkela_wire_3887),
        .b(_0971_),
        .c(_0972_)
    );

    and_bi _2393_ (
        .a(_0392_),
        .b(new_Jinkela_wire_6495),
        .c(_0396_)
    );

    bfr new_Jinkela_buffer_2430 (
        .din(new_Jinkela_wire_3673),
        .dout(new_Jinkela_wire_3674)
    );

    and_bi _1680_ (
        .a(new_Jinkela_wire_2622),
        .b(new_Jinkela_wire_3083),
        .c(_0973_)
    );

    and_bi _2394_ (
        .a(new_Jinkela_wire_681),
        .b(_0396_),
        .c(new_net_2445)
    );

    bfr new_Jinkela_buffer_2410 (
        .din(new_Jinkela_wire_3651),
        .dout(new_Jinkela_wire_3652)
    );

    and_bi _1681_ (
        .a(new_Jinkela_wire_3082),
        .b(new_Jinkela_wire_2623),
        .c(_0974_)
    );

    and_bi _2395_ (
        .a(new_Jinkela_wire_2430),
        .b(new_Jinkela_wire_803),
        .c(_0397_)
    );

    spl2 new_Jinkela_splitter_471 (
        .a(_1235_),
        .b(new_Jinkela_wire_3747),
        .c(new_Jinkela_wire_3748)
    );

    and_ii _1682_ (
        .a(_0974_),
        .b(_0973_),
        .c(_0975_)
    );

    and_bi _2396_ (
        .a(new_Jinkela_wire_7436),
        .b(new_Jinkela_wire_6823),
        .c(_0398_)
    );

    bfr new_Jinkela_buffer_2411 (
        .din(new_Jinkela_wire_3652),
        .dout(new_Jinkela_wire_3653)
    );

    or_ii _1683_ (
        .a(new_Jinkela_wire_7105),
        .b(new_Jinkela_wire_7712),
        .c(_0976_)
    );

    or_bb _2397_ (
        .a(_0398_),
        .b(new_Jinkela_wire_5574),
        .c(_0399_)
    );

    bfr new_Jinkela_buffer_2431 (
        .din(new_Jinkela_wire_3674),
        .dout(new_Jinkela_wire_3675)
    );

    or_bb _1684_ (
        .a(new_Jinkela_wire_257),
        .b(new_Jinkela_wire_420),
        .c(_0977_)
    );

    or_bb _2398_ (
        .a(new_Jinkela_wire_6093),
        .b(_0397_),
        .c(_0400_)
    );

    bfr new_Jinkela_buffer_2412 (
        .din(new_Jinkela_wire_3653),
        .dout(new_Jinkela_wire_3654)
    );

    and_bi _1685_ (
        .a(new_Jinkela_wire_261),
        .b(new_Jinkela_wire_62),
        .c(_0978_)
    );

    and_bi _2399_ (
        .a(new_Jinkela_wire_40),
        .b(new_Jinkela_wire_3384),
        .c(_0401_)
    );

    bfr new_Jinkela_buffer_2438 (
        .din(new_Jinkela_wire_3683),
        .dout(new_Jinkela_wire_3684)
    );

    and_bi _1686_ (
        .a(_0977_),
        .b(_0978_),
        .c(_0979_)
    );

    and_bi _2400_ (
        .a(new_Jinkela_wire_1353),
        .b(new_Jinkela_wire_4028),
        .c(_0402_)
    );

    bfr new_Jinkela_buffer_2413 (
        .din(new_Jinkela_wire_3654),
        .dout(new_Jinkela_wire_3655)
    );

    and_bi _1687_ (
        .a(new_Jinkela_wire_710),
        .b(_0979_),
        .c(_0980_)
    );

    or_bb _2401_ (
        .a(_0402_),
        .b(_0401_),
        .c(_0403_)
    );

    bfr new_Jinkela_buffer_2432 (
        .din(new_Jinkela_wire_3675),
        .dout(new_Jinkela_wire_3676)
    );

    or_ii _1688_ (
        .a(new_Jinkela_wire_258),
        .b(new_Jinkela_wire_1540),
        .c(_0981_)
    );

    and_bi _2402_ (
        .a(_0400_),
        .b(new_Jinkela_wire_7104),
        .c(_0404_)
    );

    bfr new_Jinkela_buffer_2414 (
        .din(new_Jinkela_wire_3655),
        .dout(new_Jinkela_wire_3656)
    );

    and_bi _1689_ (
        .a(new_Jinkela_wire_1211),
        .b(new_Jinkela_wire_260),
        .c(_0982_)
    );

    and_bi _2403_ (
        .a(new_Jinkela_wire_670),
        .b(_0404_),
        .c(new_net_2475)
    );

    and_bi _1690_ (
        .a(_0981_),
        .b(_0982_),
        .c(_0983_)
    );

    and_bi _2404_ (
        .a(new_Jinkela_wire_7937),
        .b(new_Jinkela_wire_809),
        .c(_0405_)
    );

    bfr new_Jinkela_buffer_2415 (
        .din(new_Jinkela_wire_3656),
        .dout(new_Jinkela_wire_3657)
    );

    and_bi _1691_ (
        .a(new_Jinkela_wire_6760),
        .b(_0983_),
        .c(_0984_)
    );

    and_bi _2405_ (
        .a(new_Jinkela_wire_7292),
        .b(new_Jinkela_wire_6827),
        .c(_0406_)
    );

    bfr new_Jinkela_buffer_2439 (
        .din(new_Jinkela_wire_3684),
        .dout(new_Jinkela_wire_3685)
    );

    and_ii _1692_ (
        .a(_0984_),
        .b(_0980_),
        .c(_0985_)
    );

    or_bb _2406_ (
        .a(_0406_),
        .b(new_Jinkela_wire_5578),
        .c(_0407_)
    );

    bfr new_Jinkela_buffer_2416 (
        .din(new_Jinkela_wire_3657),
        .dout(new_Jinkela_wire_3658)
    );

    and_bi _1693_ (
        .a(new_Jinkela_wire_1052),
        .b(new_Jinkela_wire_3834),
        .c(_0986_)
    );

    or_bb _2407_ (
        .a(new_Jinkela_wire_5304),
        .b(_0405_),
        .c(_0408_)
    );

    bfr new_Jinkela_buffer_2470 (
        .din(new_Jinkela_wire_3717),
        .dout(new_Jinkela_wire_3718)
    );

    or_bb _1694_ (
        .a(_0986_),
        .b(new_Jinkela_wire_4834),
        .c(_0987_)
    );

    and_bi _2408_ (
        .a(new_Jinkela_wire_1219),
        .b(new_Jinkela_wire_3382),
        .c(_0409_)
    );

    bfr new_Jinkela_buffer_2417 (
        .din(new_Jinkela_wire_3658),
        .dout(new_Jinkela_wire_3659)
    );

    and_bi _1695_ (
        .a(_0976_),
        .b(new_Jinkela_wire_3819),
        .c(_0988_)
    );

    and_bi _2409_ (
        .a(new_Jinkela_wire_1526),
        .b(new_Jinkela_wire_4030),
        .c(_0410_)
    );

    bfr new_Jinkela_buffer_2440 (
        .din(new_Jinkela_wire_3685),
        .dout(new_Jinkela_wire_3686)
    );

    and_ii _1696_ (
        .a(_0988_),
        .b(new_Jinkela_wire_7681),
        .c(new_net_17)
    );

    or_bb _2410_ (
        .a(_0410_),
        .b(_0409_),
        .c(_0411_)
    );

    bfr new_Jinkela_buffer_2418 (
        .din(new_Jinkela_wire_3659),
        .dout(new_Jinkela_wire_3660)
    );

    spl2 new_Jinkela_splitter_457 (
        .a(new_Jinkela_wire_3526),
        .b(new_Jinkela_wire_3527),
        .c(new_Jinkela_wire_3528)
    );

    bfr new_Jinkela_buffer_2209 (
        .din(new_Jinkela_wire_3348),
        .dout(new_Jinkela_wire_3349)
    );

    bfr new_Jinkela_buffer_3779 (
        .din(new_Jinkela_wire_5276),
        .dout(new_Jinkela_wire_5277)
    );

    spl2 new_Jinkela_splitter_363 (
        .a(new_net_14),
        .b(new_Jinkela_wire_2356),
        .c(new_Jinkela_wire_2357)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_2291),
        .dout(new_Jinkela_wire_2292)
    );

    bfr new_Jinkela_buffer_2232 (
        .din(new_Jinkela_wire_3395),
        .dout(new_Jinkela_wire_3396)
    );

    bfr new_Jinkela_buffer_3767 (
        .din(new_Jinkela_wire_5260),
        .dout(new_Jinkela_wire_5261)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_2318),
        .dout(new_Jinkela_wire_2319)
    );

    bfr new_Jinkela_buffer_2210 (
        .din(new_Jinkela_wire_3349),
        .dout(new_Jinkela_wire_3350)
    );

    bfr new_Jinkela_buffer_3796 (
        .din(_0407_),
        .dout(new_Jinkela_wire_5302)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(_0232_),
        .dout(new_Jinkela_wire_2397)
    );

    bfr new_Jinkela_buffer_3795 (
        .din(new_Jinkela_wire_5298),
        .dout(new_Jinkela_wire_5299)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_Jinkela_wire_2292),
        .dout(new_Jinkela_wire_2293)
    );

    bfr new_Jinkela_buffer_3768 (
        .din(new_Jinkela_wire_5261),
        .dout(new_Jinkela_wire_5262)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(new_Jinkela_wire_2333),
        .dout(new_Jinkela_wire_2334)
    );

    bfr new_Jinkela_buffer_2211 (
        .din(new_Jinkela_wire_3350),
        .dout(new_Jinkela_wire_3351)
    );

    bfr new_Jinkela_buffer_3780 (
        .din(new_Jinkela_wire_5277),
        .dout(new_Jinkela_wire_5278)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_2319),
        .dout(new_Jinkela_wire_2320)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_2293),
        .dout(new_Jinkela_wire_2294)
    );

    bfr new_Jinkela_buffer_2233 (
        .din(new_Jinkela_wire_3396),
        .dout(new_Jinkela_wire_3397)
    );

    bfr new_Jinkela_buffer_3769 (
        .din(new_Jinkela_wire_5262),
        .dout(new_Jinkela_wire_5263)
    );

    bfr new_Jinkela_buffer_2212 (
        .din(new_Jinkela_wire_3351),
        .dout(new_Jinkela_wire_3352)
    );

    bfr new_Jinkela_buffer_3786 (
        .din(new_Jinkela_wire_5286),
        .dout(new_Jinkela_wire_5287)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_2294),
        .dout(new_Jinkela_wire_2295)
    );

    bfr new_Jinkela_buffer_2248 (
        .din(new_Jinkela_wire_3417),
        .dout(new_Jinkela_wire_3418)
    );

    bfr new_Jinkela_buffer_3770 (
        .din(new_Jinkela_wire_5263),
        .dout(new_Jinkela_wire_5264)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_2357),
        .dout(new_Jinkela_wire_2358)
    );

    bfr new_Jinkela_buffer_2213 (
        .din(new_Jinkela_wire_3352),
        .dout(new_Jinkela_wire_3353)
    );

    spl3L new_Jinkela_splitter_571 (
        .a(new_Jinkela_wire_5278),
        .d(new_Jinkela_wire_5279),
        .b(new_Jinkela_wire_5280),
        .c(new_Jinkela_wire_5281)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(new_Jinkela_wire_2320),
        .dout(new_Jinkela_wire_2321)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_2295),
        .dout(new_Jinkela_wire_2296)
    );

    bfr new_Jinkela_buffer_2234 (
        .din(new_Jinkela_wire_3397),
        .dout(new_Jinkela_wire_3398)
    );

    bfr new_Jinkela_buffer_3771 (
        .din(new_Jinkela_wire_5264),
        .dout(new_Jinkela_wire_5265)
    );

    bfr new_Jinkela_buffer_2214 (
        .din(new_Jinkela_wire_3353),
        .dout(new_Jinkela_wire_3354)
    );

    bfr new_Jinkela_buffer_3799 (
        .din(new_net_2471),
        .dout(new_Jinkela_wire_5307)
    );

    bfr new_Jinkela_buffer_3797 (
        .din(new_Jinkela_wire_5302),
        .dout(new_Jinkela_wire_5303)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_2296),
        .dout(new_Jinkela_wire_2297)
    );

    bfr new_Jinkela_buffer_3772 (
        .din(new_Jinkela_wire_5265),
        .dout(new_Jinkela_wire_5266)
    );

    bfr new_Jinkela_buffer_2249 (
        .din(new_Jinkela_wire_3418),
        .dout(new_Jinkela_wire_3419)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_2334),
        .dout(new_Jinkela_wire_2335)
    );

    bfr new_Jinkela_buffer_2215 (
        .din(new_Jinkela_wire_3354),
        .dout(new_Jinkela_wire_3355)
    );

    bfr new_Jinkela_buffer_3781 (
        .din(new_Jinkela_wire_5281),
        .dout(new_Jinkela_wire_5282)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_2321),
        .dout(new_Jinkela_wire_2322)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_2297),
        .dout(new_Jinkela_wire_2298)
    );

    bfr new_Jinkela_buffer_2235 (
        .din(new_Jinkela_wire_3398),
        .dout(new_Jinkela_wire_3399)
    );

    bfr new_Jinkela_buffer_3773 (
        .din(new_Jinkela_wire_5266),
        .dout(new_Jinkela_wire_5267)
    );

    bfr new_Jinkela_buffer_3787 (
        .din(new_Jinkela_wire_5287),
        .dout(new_Jinkela_wire_5288)
    );

    bfr new_Jinkela_buffer_2275 (
        .din(new_Jinkela_wire_3467),
        .dout(new_Jinkela_wire_3468)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_2298),
        .dout(new_Jinkela_wire_2299)
    );

    bfr new_Jinkela_buffer_2236 (
        .din(new_Jinkela_wire_3399),
        .dout(new_Jinkela_wire_3400)
    );

    bfr new_Jinkela_buffer_3774 (
        .din(new_Jinkela_wire_5267),
        .dout(new_Jinkela_wire_5268)
    );

    bfr new_Jinkela_buffer_3782 (
        .din(new_Jinkela_wire_5282),
        .dout(new_Jinkela_wire_5283)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_2322),
        .dout(new_Jinkela_wire_2323)
    );

    bfr new_Jinkela_buffer_2274 (
        .din(_0224_),
        .dout(new_Jinkela_wire_3467)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_Jinkela_wire_2299),
        .dout(new_Jinkela_wire_2300)
    );

    bfr new_Jinkela_buffer_2237 (
        .din(new_Jinkela_wire_3400),
        .dout(new_Jinkela_wire_3401)
    );

    bfr new_Jinkela_buffer_3775 (
        .din(new_Jinkela_wire_5268),
        .dout(new_Jinkela_wire_5269)
    );

    spl2 new_Jinkela_splitter_446 (
        .a(_0207_),
        .b(new_Jinkela_wire_3465),
        .c(new_Jinkela_wire_3466)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_2300),
        .dout(new_Jinkela_wire_2301)
    );

    bfr new_Jinkela_buffer_2238 (
        .din(new_Jinkela_wire_3401),
        .dout(new_Jinkela_wire_3402)
    );

    bfr new_Jinkela_buffer_3776 (
        .din(new_Jinkela_wire_5269),
        .dout(new_Jinkela_wire_5270)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_2335),
        .dout(new_Jinkela_wire_2336)
    );

    bfr new_Jinkela_buffer_3788 (
        .din(new_Jinkela_wire_5288),
        .dout(new_Jinkela_wire_5289)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_2323),
        .dout(new_Jinkela_wire_2324)
    );

    bfr new_Jinkela_buffer_2277 (
        .din(new_Jinkela_wire_3469),
        .dout(new_Jinkela_wire_3470)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_2301),
        .dout(new_Jinkela_wire_2302)
    );

    bfr new_Jinkela_buffer_2239 (
        .din(new_Jinkela_wire_3402),
        .dout(new_Jinkela_wire_3403)
    );

    bfr new_Jinkela_buffer_2251 (
        .din(new_Jinkela_wire_3420),
        .dout(new_Jinkela_wire_3421)
    );

    bfr new_Jinkela_buffer_3789 (
        .din(new_Jinkela_wire_5289),
        .dout(new_Jinkela_wire_5290)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_2302),
        .dout(new_Jinkela_wire_2303)
    );

    bfr new_Jinkela_buffer_2240 (
        .din(new_Jinkela_wire_3403),
        .dout(new_Jinkela_wire_3404)
    );

    spl2 new_Jinkela_splitter_574 (
        .a(_1071_),
        .b(new_Jinkela_wire_5305),
        .c(new_Jinkela_wire_5306)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(_0141_),
        .dout(new_Jinkela_wire_2399)
    );

    bfr new_Jinkela_buffer_3790 (
        .din(new_Jinkela_wire_5290),
        .dout(new_Jinkela_wire_5291)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_2324),
        .dout(new_Jinkela_wire_2325)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_2303),
        .dout(new_Jinkela_wire_2304)
    );

    bfr new_Jinkela_buffer_2241 (
        .din(new_Jinkela_wire_3404),
        .dout(new_Jinkela_wire_3405)
    );

    bfr new_Jinkela_buffer_3800 (
        .din(new_Jinkela_wire_5307),
        .dout(new_Jinkela_wire_5308)
    );

    bfr new_Jinkela_buffer_2276 (
        .din(new_net_2473),
        .dout(new_Jinkela_wire_3469)
    );

    bfr new_Jinkela_buffer_3791 (
        .din(new_Jinkela_wire_5291),
        .dout(new_Jinkela_wire_5292)
    );

    spl2 new_Jinkela_splitter_365 (
        .a(_0177_),
        .b(new_Jinkela_wire_2404),
        .c(new_Jinkela_wire_2405)
    );

    bfr new_Jinkela_buffer_2278 (
        .din(new_Jinkela_wire_3470),
        .dout(new_Jinkela_wire_3471)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_2336),
        .dout(new_Jinkela_wire_2337)
    );

    bfr new_Jinkela_buffer_2242 (
        .din(new_Jinkela_wire_3405),
        .dout(new_Jinkela_wire_3406)
    );

    bfr new_Jinkela_buffer_3798 (
        .din(new_Jinkela_wire_5303),
        .dout(new_Jinkela_wire_5304)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_2325),
        .dout(new_Jinkela_wire_2326)
    );

    bfr new_Jinkela_buffer_3792 (
        .din(new_Jinkela_wire_5292),
        .dout(new_Jinkela_wire_5293)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(new_Jinkela_wire_2397),
        .dout(new_Jinkela_wire_2398)
    );

    bfr new_Jinkela_buffer_2243 (
        .din(new_Jinkela_wire_3406),
        .dout(new_Jinkela_wire_3407)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_2326),
        .dout(new_Jinkela_wire_2327)
    );

    bfr new_Jinkela_buffer_2287 (
        .din(_0252_),
        .dout(new_Jinkela_wire_3480)
    );

    bfr new_Jinkela_buffer_3793 (
        .din(new_Jinkela_wire_5293),
        .dout(new_Jinkela_wire_5294)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_2358),
        .dout(new_Jinkela_wire_2359)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(new_Jinkela_wire_2337),
        .dout(new_Jinkela_wire_2338)
    );

    bfr new_Jinkela_buffer_2244 (
        .din(new_Jinkela_wire_3407),
        .dout(new_Jinkela_wire_3408)
    );

    bfr new_Jinkela_buffer_3810 (
        .din(_0714_),
        .dout(new_Jinkela_wire_5318)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(new_Jinkela_wire_2327),
        .dout(new_Jinkela_wire_2328)
    );

    bfr new_Jinkela_buffer_3794 (
        .din(new_Jinkela_wire_5294),
        .dout(new_Jinkela_wire_5295)
    );

    spl4L new_Jinkela_splitter_456 (
        .a(_0769_),
        .d(new_Jinkela_wire_3523),
        .e(new_Jinkela_wire_3524),
        .b(new_Jinkela_wire_3525),
        .c(new_Jinkela_wire_3526)
    );

    bfr new_Jinkela_buffer_2245 (
        .din(new_Jinkela_wire_3408),
        .dout(new_Jinkela_wire_3409)
    );

    bfr new_Jinkela_buffer_3824 (
        .din(_0274_),
        .dout(new_Jinkela_wire_5332)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_2328),
        .dout(new_Jinkela_wire_2329)
    );

    spl2 new_Jinkela_splitter_459 (
        .a(_1088_),
        .b(new_Jinkela_wire_3534),
        .c(new_Jinkela_wire_3535)
    );

    bfr new_Jinkela_buffer_3801 (
        .din(new_Jinkela_wire_5308),
        .dout(new_Jinkela_wire_5309)
    );

    bfr new_Jinkela_buffer_2254 (
        .din(new_Jinkela_wire_3423),
        .dout(new_Jinkela_wire_3424)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(new_Jinkela_wire_2338),
        .dout(new_Jinkela_wire_2339)
    );

    bfr new_Jinkela_buffer_2246 (
        .din(new_Jinkela_wire_3409),
        .dout(new_Jinkela_wire_3410)
    );

    bfr new_Jinkela_buffer_3811 (
        .din(new_Jinkela_wire_5318),
        .dout(new_Jinkela_wire_5319)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_2329),
        .dout(new_Jinkela_wire_2330)
    );

    bfr new_Jinkela_buffer_2252 (
        .din(new_Jinkela_wire_3421),
        .dout(new_Jinkela_wire_3422)
    );

    bfr new_Jinkela_buffer_3802 (
        .din(new_Jinkela_wire_5309),
        .dout(new_Jinkela_wire_5310)
    );

    bfr new_Jinkela_buffer_2279 (
        .din(new_Jinkela_wire_3471),
        .dout(new_Jinkela_wire_3472)
    );

    bfr new_Jinkela_buffer_2255 (
        .din(new_Jinkela_wire_3424),
        .dout(new_Jinkela_wire_3425)
    );

    bfr new_Jinkela_buffer_3826 (
        .din(_0307_),
        .dout(new_Jinkela_wire_5334)
    );

    spl2 new_Jinkela_splitter_362 (
        .a(new_Jinkela_wire_2330),
        .b(new_Jinkela_wire_2331),
        .c(new_Jinkela_wire_2332)
    );

    bfr new_Jinkela_buffer_2253 (
        .din(new_Jinkela_wire_3422),
        .dout(new_Jinkela_wire_3423)
    );

    bfr new_Jinkela_buffer_2256 (
        .din(new_Jinkela_wire_3425),
        .dout(new_Jinkela_wire_3426)
    );

    bfr new_Jinkela_buffer_3803 (
        .din(new_Jinkela_wire_5310),
        .dout(new_Jinkela_wire_5311)
    );

    bfr new_Jinkela_buffer_2315 (
        .din(_0958_),
        .dout(new_Jinkela_wire_3536)
    );

    bfr new_Jinkela_buffer_2280 (
        .din(new_Jinkela_wire_3472),
        .dout(new_Jinkela_wire_3473)
    );

    bfr new_Jinkela_buffer_3812 (
        .din(new_Jinkela_wire_5319),
        .dout(new_Jinkela_wire_5320)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_2359),
        .dout(new_Jinkela_wire_2360)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_2339),
        .dout(new_Jinkela_wire_2340)
    );

    bfr new_Jinkela_buffer_3804 (
        .din(new_Jinkela_wire_5311),
        .dout(new_Jinkela_wire_5312)
    );

    spl3L new_Jinkela_splitter_366 (
        .a(_0619_),
        .d(new_Jinkela_wire_2406),
        .b(new_Jinkela_wire_2407),
        .c(new_Jinkela_wire_2408)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(new_Jinkela_wire_2340),
        .dout(new_Jinkela_wire_2341)
    );

    bfr new_Jinkela_buffer_3825 (
        .din(new_Jinkela_wire_5332),
        .dout(new_Jinkela_wire_5333)
    );

    bfr new_Jinkela_buffer_3034 (
        .din(new_Jinkela_wire_4385),
        .dout(new_Jinkela_wire_4386)
    );

    bfr new_Jinkela_buffer_3024 (
        .din(new_Jinkela_wire_4369),
        .dout(new_Jinkela_wire_4370)
    );

    bfr new_Jinkela_buffer_3061 (
        .din(new_Jinkela_wire_4414),
        .dout(new_Jinkela_wire_4415)
    );

    bfr new_Jinkela_buffer_3025 (
        .din(new_Jinkela_wire_4370),
        .dout(new_Jinkela_wire_4371)
    );

    bfr new_Jinkela_buffer_3035 (
        .din(new_Jinkela_wire_4386),
        .dout(new_Jinkela_wire_4387)
    );

    bfr new_Jinkela_buffer_3026 (
        .din(new_Jinkela_wire_4371),
        .dout(new_Jinkela_wire_4372)
    );

    bfr new_Jinkela_buffer_3027 (
        .din(new_Jinkela_wire_4372),
        .dout(new_Jinkela_wire_4373)
    );

    bfr new_Jinkela_buffer_3036 (
        .din(new_Jinkela_wire_4387),
        .dout(new_Jinkela_wire_4388)
    );

    bfr new_Jinkela_buffer_3028 (
        .din(new_Jinkela_wire_4373),
        .dout(new_Jinkela_wire_4374)
    );

    bfr new_Jinkela_buffer_3062 (
        .din(new_Jinkela_wire_4415),
        .dout(new_Jinkela_wire_4416)
    );

    bfr new_Jinkela_buffer_3029 (
        .din(new_Jinkela_wire_4374),
        .dout(new_Jinkela_wire_4375)
    );

    bfr new_Jinkela_buffer_3037 (
        .din(new_Jinkela_wire_4388),
        .dout(new_Jinkela_wire_4389)
    );

    bfr new_Jinkela_buffer_3030 (
        .din(new_Jinkela_wire_4375),
        .dout(new_Jinkela_wire_4376)
    );

    bfr new_Jinkela_buffer_3098 (
        .din(_0634_),
        .dout(new_Jinkela_wire_4454)
    );

    bfr new_Jinkela_buffer_3038 (
        .din(new_Jinkela_wire_4389),
        .dout(new_Jinkela_wire_4390)
    );

    bfr new_Jinkela_buffer_3063 (
        .din(new_Jinkela_wire_4416),
        .dout(new_Jinkela_wire_4417)
    );

    bfr new_Jinkela_buffer_3039 (
        .din(new_Jinkela_wire_4390),
        .dout(new_Jinkela_wire_4391)
    );

    bfr new_Jinkela_buffer_3073 (
        .din(new_Jinkela_wire_4428),
        .dout(new_Jinkela_wire_4429)
    );

    bfr new_Jinkela_buffer_3071 (
        .din(new_Jinkela_wire_4426),
        .dout(new_Jinkela_wire_4427)
    );

    bfr new_Jinkela_buffer_3040 (
        .din(new_Jinkela_wire_4391),
        .dout(new_Jinkela_wire_4392)
    );

    bfr new_Jinkela_buffer_3064 (
        .din(new_Jinkela_wire_4417),
        .dout(new_Jinkela_wire_4418)
    );

    bfr new_Jinkela_buffer_3041 (
        .din(new_Jinkela_wire_4392),
        .dout(new_Jinkela_wire_4393)
    );

    bfr new_Jinkela_buffer_3042 (
        .din(new_Jinkela_wire_4393),
        .dout(new_Jinkela_wire_4394)
    );

    bfr new_Jinkela_buffer_3065 (
        .din(new_Jinkela_wire_4418),
        .dout(new_Jinkela_wire_4419)
    );

    bfr new_Jinkela_buffer_3043 (
        .din(new_Jinkela_wire_4394),
        .dout(new_Jinkela_wire_4395)
    );

    spl2 new_Jinkela_splitter_516 (
        .a(_0698_),
        .b(new_Jinkela_wire_4464),
        .c(new_Jinkela_wire_4465)
    );

    bfr new_Jinkela_buffer_3108 (
        .din(_0387_),
        .dout(new_Jinkela_wire_4466)
    );

    bfr new_Jinkela_buffer_3044 (
        .din(new_Jinkela_wire_4395),
        .dout(new_Jinkela_wire_4396)
    );

    bfr new_Jinkela_buffer_3066 (
        .din(new_Jinkela_wire_4419),
        .dout(new_Jinkela_wire_4420)
    );

    bfr new_Jinkela_buffer_3045 (
        .din(new_Jinkela_wire_4396),
        .dout(new_Jinkela_wire_4397)
    );

    bfr new_Jinkela_buffer_3074 (
        .din(new_Jinkela_wire_4429),
        .dout(new_Jinkela_wire_4430)
    );

    bfr new_Jinkela_buffer_3046 (
        .din(new_Jinkela_wire_4397),
        .dout(new_Jinkela_wire_4398)
    );

    bfr new_Jinkela_buffer_3067 (
        .din(new_Jinkela_wire_4420),
        .dout(new_Jinkela_wire_4421)
    );

    bfr new_Jinkela_buffer_3047 (
        .din(new_Jinkela_wire_4398),
        .dout(new_Jinkela_wire_4399)
    );

    bfr new_Jinkela_buffer_3099 (
        .din(new_Jinkela_wire_4454),
        .dout(new_Jinkela_wire_4455)
    );

    bfr new_Jinkela_buffer_3048 (
        .din(new_Jinkela_wire_4399),
        .dout(new_Jinkela_wire_4400)
    );

    bfr new_Jinkela_buffer_3068 (
        .din(new_Jinkela_wire_4421),
        .dout(new_Jinkela_wire_4422)
    );

    bfr new_Jinkela_buffer_3049 (
        .din(new_Jinkela_wire_4400),
        .dout(new_Jinkela_wire_4401)
    );

    bfr new_Jinkela_buffer_3075 (
        .din(new_Jinkela_wire_4430),
        .dout(new_Jinkela_wire_4431)
    );

    bfr new_Jinkela_buffer_3050 (
        .din(new_Jinkela_wire_4401),
        .dout(new_Jinkela_wire_4402)
    );

    bfr new_Jinkela_buffer_3069 (
        .din(new_Jinkela_wire_4422),
        .dout(new_Jinkela_wire_4423)
    );

    bfr new_Jinkela_buffer_3051 (
        .din(new_Jinkela_wire_4402),
        .dout(new_Jinkela_wire_4403)
    );

    bfr new_Jinkela_buffer_2514 (
        .din(_0949_),
        .dout(new_Jinkela_wire_3770)
    );

    bfr new_Jinkela_buffer_3805 (
        .din(new_Jinkela_wire_5312),
        .dout(new_Jinkela_wire_5313)
    );

    spl4L new_Jinkela_splitter_472 (
        .a(_0087_),
        .d(new_Jinkela_wire_3750),
        .e(new_Jinkela_wire_3751),
        .b(new_Jinkela_wire_3752),
        .c(new_Jinkela_wire_3753)
    );

    bfr new_Jinkela_buffer_2419 (
        .din(new_Jinkela_wire_3660),
        .dout(new_Jinkela_wire_3661)
    );

    bfr new_Jinkela_buffer_3813 (
        .din(new_Jinkela_wire_5320),
        .dout(new_Jinkela_wire_5321)
    );

    bfr new_Jinkela_buffer_2441 (
        .din(new_Jinkela_wire_3686),
        .dout(new_Jinkela_wire_3687)
    );

    bfr new_Jinkela_buffer_3806 (
        .din(new_Jinkela_wire_5313),
        .dout(new_Jinkela_wire_5314)
    );

    bfr new_Jinkela_buffer_2471 (
        .din(new_Jinkela_wire_3718),
        .dout(new_Jinkela_wire_3719)
    );

    spl2 new_Jinkela_splitter_575 (
        .a(new_net_21),
        .b(new_Jinkela_wire_5358),
        .c(new_Jinkela_wire_5360)
    );

    bfr new_Jinkela_buffer_3858 (
        .din(_0732_),
        .dout(new_Jinkela_wire_5372)
    );

    bfr new_Jinkela_buffer_2442 (
        .din(new_Jinkela_wire_3687),
        .dout(new_Jinkela_wire_3688)
    );

    bfr new_Jinkela_buffer_3807 (
        .din(new_Jinkela_wire_5314),
        .dout(new_Jinkela_wire_5315)
    );

    bfr new_Jinkela_buffer_2500 (
        .din(_0832_),
        .dout(new_Jinkela_wire_3754)
    );

    bfr new_Jinkela_buffer_3814 (
        .din(new_Jinkela_wire_5321),
        .dout(new_Jinkela_wire_5322)
    );

    bfr new_Jinkela_buffer_2443 (
        .din(new_Jinkela_wire_3688),
        .dout(new_Jinkela_wire_3689)
    );

    bfr new_Jinkela_buffer_3808 (
        .din(new_Jinkela_wire_5315),
        .dout(new_Jinkela_wire_5316)
    );

    bfr new_Jinkela_buffer_2472 (
        .din(new_Jinkela_wire_3719),
        .dout(new_Jinkela_wire_3720)
    );

    bfr new_Jinkela_buffer_3827 (
        .din(new_Jinkela_wire_5334),
        .dout(new_Jinkela_wire_5335)
    );

    bfr new_Jinkela_buffer_2444 (
        .din(new_Jinkela_wire_3689),
        .dout(new_Jinkela_wire_3690)
    );

    bfr new_Jinkela_buffer_3809 (
        .din(new_Jinkela_wire_5316),
        .dout(new_Jinkela_wire_5317)
    );

    bfr new_Jinkela_buffer_2539 (
        .din(_0987_),
        .dout(new_Jinkela_wire_3799)
    );

    bfr new_Jinkela_buffer_3815 (
        .din(new_Jinkela_wire_5322),
        .dout(new_Jinkela_wire_5323)
    );

    bfr new_Jinkela_buffer_2501 (
        .din(new_Jinkela_wire_3754),
        .dout(new_Jinkela_wire_3755)
    );

    bfr new_Jinkela_buffer_2445 (
        .din(new_Jinkela_wire_3690),
        .dout(new_Jinkela_wire_3691)
    );

    bfr new_Jinkela_buffer_3878 (
        .din(_1105_),
        .dout(new_Jinkela_wire_5394)
    );

    bfr new_Jinkela_buffer_3851 (
        .din(new_Jinkela_wire_5364),
        .dout(new_Jinkela_wire_5365)
    );

    bfr new_Jinkela_buffer_2473 (
        .din(new_Jinkela_wire_3720),
        .dout(new_Jinkela_wire_3721)
    );

    bfr new_Jinkela_buffer_3816 (
        .din(new_Jinkela_wire_5323),
        .dout(new_Jinkela_wire_5324)
    );

    bfr new_Jinkela_buffer_2446 (
        .din(new_Jinkela_wire_3691),
        .dout(new_Jinkela_wire_3692)
    );

    bfr new_Jinkela_buffer_3828 (
        .din(new_Jinkela_wire_5335),
        .dout(new_Jinkela_wire_5336)
    );

    bfr new_Jinkela_buffer_3817 (
        .din(new_Jinkela_wire_5324),
        .dout(new_Jinkela_wire_5325)
    );

    bfr new_Jinkela_buffer_2513 (
        .din(_0201_),
        .dout(new_Jinkela_wire_3767)
    );

    bfr new_Jinkela_buffer_2447 (
        .din(new_Jinkela_wire_3692),
        .dout(new_Jinkela_wire_3693)
    );

    bfr new_Jinkela_buffer_3850 (
        .din(new_Jinkela_wire_5358),
        .dout(new_Jinkela_wire_5359)
    );

    spl4L new_Jinkela_splitter_576 (
        .a(new_Jinkela_wire_5360),
        .d(new_Jinkela_wire_5361),
        .e(new_Jinkela_wire_5362),
        .b(new_Jinkela_wire_5363),
        .c(new_Jinkela_wire_5364)
    );

    bfr new_Jinkela_buffer_2474 (
        .din(new_Jinkela_wire_3721),
        .dout(new_Jinkela_wire_3722)
    );

    bfr new_Jinkela_buffer_3818 (
        .din(new_Jinkela_wire_5325),
        .dout(new_Jinkela_wire_5326)
    );

    bfr new_Jinkela_buffer_2448 (
        .din(new_Jinkela_wire_3693),
        .dout(new_Jinkela_wire_3694)
    );

    bfr new_Jinkela_buffer_3829 (
        .din(new_Jinkela_wire_5336),
        .dout(new_Jinkela_wire_5337)
    );

    bfr new_Jinkela_buffer_3819 (
        .din(new_Jinkela_wire_5326),
        .dout(new_Jinkela_wire_5327)
    );

    bfr new_Jinkela_buffer_2517 (
        .din(_0911_),
        .dout(new_Jinkela_wire_3777)
    );

    bfr new_Jinkela_buffer_2449 (
        .din(new_Jinkela_wire_3694),
        .dout(new_Jinkela_wire_3695)
    );

    bfr new_Jinkela_buffer_3877 (
        .din(_0121_),
        .dout(new_Jinkela_wire_5391)
    );

    bfr new_Jinkela_buffer_2475 (
        .din(new_Jinkela_wire_3722),
        .dout(new_Jinkela_wire_3723)
    );

    bfr new_Jinkela_buffer_3820 (
        .din(new_Jinkela_wire_5327),
        .dout(new_Jinkela_wire_5328)
    );

    bfr new_Jinkela_buffer_2450 (
        .din(new_Jinkela_wire_3695),
        .dout(new_Jinkela_wire_3696)
    );

    bfr new_Jinkela_buffer_3830 (
        .din(new_Jinkela_wire_5337),
        .dout(new_Jinkela_wire_5338)
    );

    bfr new_Jinkela_buffer_2502 (
        .din(new_Jinkela_wire_3755),
        .dout(new_Jinkela_wire_3756)
    );

    bfr new_Jinkela_buffer_3821 (
        .din(new_Jinkela_wire_5328),
        .dout(new_Jinkela_wire_5329)
    );

    bfr new_Jinkela_buffer_2451 (
        .din(new_Jinkela_wire_3696),
        .dout(new_Jinkela_wire_3697)
    );

    bfr new_Jinkela_buffer_2476 (
        .din(new_Jinkela_wire_3723),
        .dout(new_Jinkela_wire_3724)
    );

    bfr new_Jinkela_buffer_3822 (
        .din(new_Jinkela_wire_5329),
        .dout(new_Jinkela_wire_5330)
    );

    bfr new_Jinkela_buffer_2452 (
        .din(new_Jinkela_wire_3697),
        .dout(new_Jinkela_wire_3698)
    );

    bfr new_Jinkela_buffer_3831 (
        .din(new_Jinkela_wire_5338),
        .dout(new_Jinkela_wire_5339)
    );

    spl2 new_Jinkela_splitter_473 (
        .a(new_Jinkela_wire_3767),
        .b(new_Jinkela_wire_3768),
        .c(new_Jinkela_wire_3769)
    );

    bfr new_Jinkela_buffer_3823 (
        .din(new_Jinkela_wire_5330),
        .dout(new_Jinkela_wire_5331)
    );

    bfr new_Jinkela_buffer_2453 (
        .din(new_Jinkela_wire_3698),
        .dout(new_Jinkela_wire_3699)
    );

    bfr new_Jinkela_buffer_2477 (
        .din(new_Jinkela_wire_3724),
        .dout(new_Jinkela_wire_3725)
    );

    bfr new_Jinkela_buffer_3832 (
        .din(new_Jinkela_wire_5339),
        .dout(new_Jinkela_wire_5340)
    );

    bfr new_Jinkela_buffer_2454 (
        .din(new_Jinkela_wire_3699),
        .dout(new_Jinkela_wire_3700)
    );

    bfr new_Jinkela_buffer_3859 (
        .din(new_Jinkela_wire_5372),
        .dout(new_Jinkela_wire_5373)
    );

    bfr new_Jinkela_buffer_2503 (
        .din(new_Jinkela_wire_3756),
        .dout(new_Jinkela_wire_3757)
    );

    bfr new_Jinkela_buffer_3833 (
        .din(new_Jinkela_wire_5340),
        .dout(new_Jinkela_wire_5341)
    );

    bfr new_Jinkela_buffer_2455 (
        .din(new_Jinkela_wire_3700),
        .dout(new_Jinkela_wire_3701)
    );

    spl2 new_Jinkela_splitter_578 (
        .a(_0895_),
        .b(new_Jinkela_wire_5395),
        .c(new_Jinkela_wire_5396)
    );

    bfr new_Jinkela_buffer_2478 (
        .din(new_Jinkela_wire_3725),
        .dout(new_Jinkela_wire_3726)
    );

    bfr new_Jinkela_buffer_3834 (
        .din(new_Jinkela_wire_5341),
        .dout(new_Jinkela_wire_5342)
    );

    bfr new_Jinkela_buffer_2456 (
        .din(new_Jinkela_wire_3701),
        .dout(new_Jinkela_wire_3702)
    );

    bfr new_Jinkela_buffer_3852 (
        .din(new_Jinkela_wire_5365),
        .dout(new_Jinkela_wire_5366)
    );

    bfr new_Jinkela_buffer_3835 (
        .din(new_Jinkela_wire_5342),
        .dout(new_Jinkela_wire_5343)
    );

    bfr new_Jinkela_buffer_2457 (
        .din(new_Jinkela_wire_3702),
        .dout(new_Jinkela_wire_3703)
    );

    bfr new_Jinkela_buffer_3860 (
        .din(new_Jinkela_wire_5373),
        .dout(new_Jinkela_wire_5374)
    );

    bfr new_Jinkela_buffer_2479 (
        .din(new_Jinkela_wire_3726),
        .dout(new_Jinkela_wire_3727)
    );

    bfr new_Jinkela_buffer_3836 (
        .din(new_Jinkela_wire_5343),
        .dout(new_Jinkela_wire_5344)
    );

    bfr new_Jinkela_buffer_2458 (
        .din(new_Jinkela_wire_3703),
        .dout(new_Jinkela_wire_3704)
    );

    bfr new_Jinkela_buffer_3853 (
        .din(new_Jinkela_wire_5366),
        .dout(new_Jinkela_wire_5367)
    );

    bfr new_Jinkela_buffer_2504 (
        .din(new_Jinkela_wire_3757),
        .dout(new_Jinkela_wire_3758)
    );

    bfr new_Jinkela_buffer_3837 (
        .din(new_Jinkela_wire_5344),
        .dout(new_Jinkela_wire_5345)
    );

    bfr new_Jinkela_buffer_2459 (
        .din(new_Jinkela_wire_3704),
        .dout(new_Jinkela_wire_3705)
    );

    spl2 new_Jinkela_splitter_577 (
        .a(new_Jinkela_wire_5391),
        .b(new_Jinkela_wire_5392),
        .c(new_Jinkela_wire_5393)
    );

    bfr new_Jinkela_buffer_2480 (
        .din(new_Jinkela_wire_3727),
        .dout(new_Jinkela_wire_3728)
    );

    bfr new_Jinkela_buffer_3838 (
        .din(new_Jinkela_wire_5345),
        .dout(new_Jinkela_wire_5346)
    );

    bfr new_Jinkela_buffer_2460 (
        .din(new_Jinkela_wire_3705),
        .dout(new_Jinkela_wire_3706)
    );

    bfr new_Jinkela_buffer_3854 (
        .din(new_Jinkela_wire_5367),
        .dout(new_Jinkela_wire_5368)
    );

    bfr new_Jinkela_buffer_3839 (
        .din(new_Jinkela_wire_5346),
        .dout(new_Jinkela_wire_5347)
    );

    bfr new_Jinkela_buffer_2257 (
        .din(new_Jinkela_wire_3426),
        .dout(new_Jinkela_wire_3427)
    );

    bfr new_Jinkela_buffer_2318 (
        .din(_0462_),
        .dout(new_Jinkela_wire_3539)
    );

    bfr new_Jinkela_buffer_2258 (
        .din(new_Jinkela_wire_3427),
        .dout(new_Jinkela_wire_3428)
    );

    bfr new_Jinkela_buffer_2312 (
        .din(new_Jinkela_wire_3528),
        .dout(new_Jinkela_wire_3529)
    );

    bfr new_Jinkela_buffer_2281 (
        .din(new_Jinkela_wire_3473),
        .dout(new_Jinkela_wire_3474)
    );

    bfr new_Jinkela_buffer_2259 (
        .din(new_Jinkela_wire_3428),
        .dout(new_Jinkela_wire_3429)
    );

    bfr new_Jinkela_buffer_2260 (
        .din(new_Jinkela_wire_3429),
        .dout(new_Jinkela_wire_3430)
    );

    bfr new_Jinkela_buffer_2282 (
        .din(new_Jinkela_wire_3474),
        .dout(new_Jinkela_wire_3475)
    );

    bfr new_Jinkela_buffer_2261 (
        .din(new_Jinkela_wire_3430),
        .dout(new_Jinkela_wire_3431)
    );

    bfr new_Jinkela_buffer_2316 (
        .din(new_Jinkela_wire_3536),
        .dout(new_Jinkela_wire_3537)
    );

    spl2 new_Jinkela_splitter_437 (
        .a(new_Jinkela_wire_3431),
        .b(new_Jinkela_wire_3432),
        .c(new_Jinkela_wire_3433)
    );

    bfr new_Jinkela_buffer_2262 (
        .din(new_Jinkela_wire_3433),
        .dout(new_Jinkela_wire_3434)
    );

    bfr new_Jinkela_buffer_2288 (
        .din(new_Jinkela_wire_3480),
        .dout(new_Jinkela_wire_3481)
    );

    bfr new_Jinkela_buffer_2283 (
        .din(new_Jinkela_wire_3475),
        .dout(new_Jinkela_wire_3476)
    );

    spl2 new_Jinkela_splitter_438 (
        .a(new_Jinkela_wire_3434),
        .b(new_Jinkela_wire_3435),
        .c(new_Jinkela_wire_3436)
    );

    bfr new_Jinkela_buffer_2263 (
        .din(new_Jinkela_wire_3436),
        .dout(new_Jinkela_wire_3437)
    );

    bfr new_Jinkela_buffer_2284 (
        .din(new_Jinkela_wire_3476),
        .dout(new_Jinkela_wire_3477)
    );

    bfr new_Jinkela_buffer_2289 (
        .din(new_Jinkela_wire_3481),
        .dout(new_Jinkela_wire_3482)
    );

    spl2 new_Jinkela_splitter_439 (
        .a(new_Jinkela_wire_3437),
        .b(new_Jinkela_wire_3438),
        .c(new_Jinkela_wire_3439)
    );

    spl2 new_Jinkela_splitter_440 (
        .a(new_Jinkela_wire_3439),
        .b(new_Jinkela_wire_3440),
        .c(new_Jinkela_wire_3441)
    );

    bfr new_Jinkela_buffer_2313 (
        .din(new_Jinkela_wire_3529),
        .dout(new_Jinkela_wire_3530)
    );

    bfr new_Jinkela_buffer_2285 (
        .din(new_Jinkela_wire_3477),
        .dout(new_Jinkela_wire_3478)
    );

    bfr new_Jinkela_buffer_2264 (
        .din(new_Jinkela_wire_3441),
        .dout(new_Jinkela_wire_3442)
    );

    bfr new_Jinkela_buffer_2286 (
        .din(new_Jinkela_wire_3478),
        .dout(new_Jinkela_wire_3479)
    );

    bfr new_Jinkela_buffer_2265 (
        .din(new_Jinkela_wire_3442),
        .dout(new_Jinkela_wire_3443)
    );

    bfr new_Jinkela_buffer_2353 (
        .din(_0287_),
        .dout(new_Jinkela_wire_3577)
    );

    spl3L new_Jinkela_splitter_441 (
        .a(new_Jinkela_wire_3443),
        .d(new_Jinkela_wire_3444),
        .b(new_Jinkela_wire_3445),
        .c(new_Jinkela_wire_3446)
    );

    bfr new_Jinkela_buffer_2290 (
        .din(new_Jinkela_wire_3482),
        .dout(new_Jinkela_wire_3483)
    );

    bfr new_Jinkela_buffer_2266 (
        .din(new_Jinkela_wire_3446),
        .dout(new_Jinkela_wire_3447)
    );

    bfr new_Jinkela_buffer_2350 (
        .din(_0943_),
        .dout(new_Jinkela_wire_3571)
    );

    spl2 new_Jinkela_splitter_442 (
        .a(new_Jinkela_wire_3447),
        .b(new_Jinkela_wire_3448),
        .c(new_Jinkela_wire_3449)
    );

    bfr new_Jinkela_buffer_2267 (
        .din(new_Jinkela_wire_3449),
        .dout(new_Jinkela_wire_3450)
    );

    bfr new_Jinkela_buffer_2291 (
        .din(new_Jinkela_wire_3483),
        .dout(new_Jinkela_wire_3484)
    );

    bfr new_Jinkela_buffer_2317 (
        .din(new_Jinkela_wire_3537),
        .dout(new_Jinkela_wire_3538)
    );

    spl4L new_Jinkela_splitter_443 (
        .a(new_Jinkela_wire_3450),
        .d(new_Jinkela_wire_3451),
        .e(new_Jinkela_wire_3452),
        .b(new_Jinkela_wire_3453),
        .c(new_Jinkela_wire_3454)
    );

    spl2 new_Jinkela_splitter_444 (
        .a(new_Jinkela_wire_3454),
        .b(new_Jinkela_wire_3455),
        .c(new_Jinkela_wire_3456)
    );

    bfr new_Jinkela_buffer_2292 (
        .din(new_Jinkela_wire_3484),
        .dout(new_Jinkela_wire_3485)
    );

    bfr new_Jinkela_buffer_2314 (
        .din(new_Jinkela_wire_3530),
        .dout(new_Jinkela_wire_3531)
    );

    bfr new_Jinkela_buffer_2268 (
        .din(new_Jinkela_wire_3456),
        .dout(new_Jinkela_wire_3457)
    );

    bfr new_Jinkela_buffer_2293 (
        .din(new_Jinkela_wire_3485),
        .dout(new_Jinkela_wire_3486)
    );

    bfr new_Jinkela_buffer_2319 (
        .din(new_Jinkela_wire_3539),
        .dout(new_Jinkela_wire_3540)
    );

    bfr new_Jinkela_buffer_2269 (
        .din(new_Jinkela_wire_3457),
        .dout(new_Jinkela_wire_3458)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_2232),
        .dout(new_Jinkela_wire_2233)
    );

    bfr new_Jinkela_buffer_2976 (
        .din(new_Jinkela_wire_4303),
        .dout(new_Jinkela_wire_4304)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_Jinkela_wire_2256),
        .dout(new_Jinkela_wire_2257)
    );

    bfr new_Jinkela_buffer_3005 (
        .din(_1058_),
        .dout(new_Jinkela_wire_4345)
    );

    bfr new_Jinkela_buffer_3006 (
        .din(new_Jinkela_wire_4349),
        .dout(new_Jinkela_wire_4350)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_2233),
        .dout(new_Jinkela_wire_2234)
    );

    bfr new_Jinkela_buffer_2977 (
        .din(new_Jinkela_wire_4304),
        .dout(new_Jinkela_wire_4305)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(new_Jinkela_wire_2272),
        .dout(new_Jinkela_wire_2273)
    );

    bfr new_Jinkela_buffer_2998 (
        .din(new_Jinkela_wire_4329),
        .dout(new_Jinkela_wire_4330)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(new_Jinkela_wire_2234),
        .dout(new_Jinkela_wire_2235)
    );

    bfr new_Jinkela_buffer_2978 (
        .din(new_Jinkela_wire_4305),
        .dout(new_Jinkela_wire_4306)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_2257),
        .dout(new_Jinkela_wire_2258)
    );

    bfr new_Jinkela_buffer_3013 (
        .din(_0658_),
        .dout(new_Jinkela_wire_4359)
    );

    spl2 new_Jinkela_splitter_509 (
        .a(_0620_),
        .b(new_Jinkela_wire_4343),
        .c(new_Jinkela_wire_4344)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(new_Jinkela_wire_2235),
        .dout(new_Jinkela_wire_2236)
    );

    bfr new_Jinkela_buffer_2979 (
        .din(new_Jinkela_wire_4306),
        .dout(new_Jinkela_wire_4307)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_2282),
        .dout(new_Jinkela_wire_2283)
    );

    bfr new_Jinkela_buffer_2999 (
        .din(new_Jinkela_wire_4330),
        .dout(new_Jinkela_wire_4331)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_2236),
        .dout(new_Jinkela_wire_2237)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_2258),
        .dout(new_Jinkela_wire_2259)
    );

    bfr new_Jinkela_buffer_3000 (
        .din(new_Jinkela_wire_4331),
        .dout(new_Jinkela_wire_4332)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(new_Jinkela_wire_2237),
        .dout(new_Jinkela_wire_2238)
    );

    spl4L new_Jinkela_splitter_510 (
        .a(_0684_),
        .d(new_Jinkela_wire_4346),
        .e(new_Jinkela_wire_4347),
        .b(new_Jinkela_wire_4348),
        .c(new_Jinkela_wire_4349)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_2273),
        .dout(new_Jinkela_wire_2274)
    );

    bfr new_Jinkela_buffer_3001 (
        .din(new_Jinkela_wire_4332),
        .dout(new_Jinkela_wire_4333)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(new_Jinkela_wire_2238),
        .dout(new_Jinkela_wire_2239)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_2259),
        .dout(new_Jinkela_wire_2260)
    );

    bfr new_Jinkela_buffer_3002 (
        .din(new_Jinkela_wire_4333),
        .dout(new_Jinkela_wire_4334)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(new_Jinkela_wire_2239),
        .dout(new_Jinkela_wire_2240)
    );

    spl2 new_Jinkela_splitter_512 (
        .a(new_net_4),
        .b(new_Jinkela_wire_4377),
        .c(new_Jinkela_wire_4379)
    );

    bfr new_Jinkela_buffer_3008 (
        .din(new_Jinkela_wire_4351),
        .dout(new_Jinkela_wire_4352)
    );

    bfr new_Jinkela_buffer_3003 (
        .din(new_Jinkela_wire_4334),
        .dout(new_Jinkela_wire_4335)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(_0070_),
        .dout(new_Jinkela_wire_2315)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(new_Jinkela_wire_2240),
        .dout(new_Jinkela_wire_2241)
    );

    spl2 new_Jinkela_splitter_514 (
        .a(_0994_),
        .b(new_Jinkela_wire_4411),
        .c(new_Jinkela_wire_4412)
    );

    spl2 new_Jinkela_splitter_355 (
        .a(new_Jinkela_wire_2260),
        .b(new_Jinkela_wire_2261),
        .c(new_Jinkela_wire_2262)
    );

    bfr new_Jinkela_buffer_3007 (
        .din(new_Jinkela_wire_4350),
        .dout(new_Jinkela_wire_4351)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(new_Jinkela_wire_2241),
        .dout(new_Jinkela_wire_2242)
    );

    bfr new_Jinkela_buffer_3060 (
        .din(new_Jinkela_wire_4413),
        .dout(new_Jinkela_wire_4414)
    );

    bfr new_Jinkela_buffer_3032 (
        .din(new_Jinkela_wire_4383),
        .dout(new_Jinkela_wire_4384)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(new_Jinkela_wire_2283),
        .dout(new_Jinkela_wire_2284)
    );

    bfr new_Jinkela_buffer_3014 (
        .din(new_Jinkela_wire_4359),
        .dout(new_Jinkela_wire_4360)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(new_Jinkela_wire_2242),
        .dout(new_Jinkela_wire_2243)
    );

    bfr new_Jinkela_buffer_3015 (
        .din(new_Jinkela_wire_4360),
        .dout(new_Jinkela_wire_4361)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(new_Jinkela_wire_2274),
        .dout(new_Jinkela_wire_2275)
    );

    bfr new_Jinkela_buffer_3009 (
        .din(new_Jinkela_wire_4352),
        .dout(new_Jinkela_wire_4353)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_2275),
        .dout(new_Jinkela_wire_2276)
    );

    bfr new_Jinkela_buffer_3031 (
        .din(new_Jinkela_wire_4377),
        .dout(new_Jinkela_wire_4378)
    );

    spl4L new_Jinkela_splitter_513 (
        .a(new_Jinkela_wire_4379),
        .d(new_Jinkela_wire_4380),
        .e(new_Jinkela_wire_4381),
        .b(new_Jinkela_wire_4382),
        .c(new_Jinkela_wire_4383)
    );

    bfr new_Jinkela_buffer_3010 (
        .din(new_Jinkela_wire_4353),
        .dout(new_Jinkela_wire_4354)
    );

    spl3L new_Jinkela_splitter_359 (
        .a(_1050_),
        .d(new_Jinkela_wire_2309),
        .b(new_Jinkela_wire_2310),
        .c(new_Jinkela_wire_2311)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_2276),
        .dout(new_Jinkela_wire_2277)
    );

    bfr new_Jinkela_buffer_3016 (
        .din(new_Jinkela_wire_4361),
        .dout(new_Jinkela_wire_4362)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_2284),
        .dout(new_Jinkela_wire_2285)
    );

    bfr new_Jinkela_buffer_3011 (
        .din(new_Jinkela_wire_4354),
        .dout(new_Jinkela_wire_4355)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(new_Jinkela_wire_2277),
        .dout(new_Jinkela_wire_2278)
    );

    bfr new_Jinkela_buffer_3072 (
        .din(_0989_),
        .dout(new_Jinkela_wire_4428)
    );

    spl2 new_Jinkela_splitter_360 (
        .a(_0144_),
        .b(new_Jinkela_wire_2313),
        .c(new_Jinkela_wire_2314)
    );

    bfr new_Jinkela_buffer_3012 (
        .din(new_Jinkela_wire_4355),
        .dout(new_Jinkela_wire_4356)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(_1117_),
        .dout(new_Jinkela_wire_2312)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(new_Jinkela_wire_2278),
        .dout(new_Jinkela_wire_2279)
    );

    bfr new_Jinkela_buffer_3017 (
        .din(new_Jinkela_wire_4362),
        .dout(new_Jinkela_wire_4363)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_2285),
        .dout(new_Jinkela_wire_2286)
    );

    spl2 new_Jinkela_splitter_511 (
        .a(new_Jinkela_wire_4356),
        .b(new_Jinkela_wire_4357),
        .c(new_Jinkela_wire_4358)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_2279),
        .dout(new_Jinkela_wire_2280)
    );

    bfr new_Jinkela_buffer_3018 (
        .din(new_Jinkela_wire_4363),
        .dout(new_Jinkela_wire_4364)
    );

    bfr new_Jinkela_buffer_3059 (
        .din(new_net_2413),
        .dout(new_Jinkela_wire_4413)
    );

    spl2 new_Jinkela_splitter_361 (
        .a(new_Jinkela_wire_2315),
        .b(new_Jinkela_wire_2316),
        .c(new_Jinkela_wire_2317)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_2280),
        .dout(new_Jinkela_wire_2281)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_2286),
        .dout(new_Jinkela_wire_2287)
    );

    bfr new_Jinkela_buffer_3019 (
        .din(new_Jinkela_wire_4364),
        .dout(new_Jinkela_wire_4365)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_2287),
        .dout(new_Jinkela_wire_2288)
    );

    bfr new_Jinkela_buffer_3020 (
        .din(new_Jinkela_wire_4365),
        .dout(new_Jinkela_wire_4366)
    );

    spl2 new_Jinkela_splitter_515 (
        .a(_0752_),
        .b(new_Jinkela_wire_4424),
        .c(new_Jinkela_wire_4425)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(_1118_),
        .dout(new_Jinkela_wire_2318)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_2288),
        .dout(new_Jinkela_wire_2289)
    );

    bfr new_Jinkela_buffer_3021 (
        .din(new_Jinkela_wire_4366),
        .dout(new_Jinkela_wire_4367)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(_1029_),
        .dout(new_Jinkela_wire_2333)
    );

    bfr new_Jinkela_buffer_3033 (
        .din(new_Jinkela_wire_4384),
        .dout(new_Jinkela_wire_4385)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_2289),
        .dout(new_Jinkela_wire_2290)
    );

    bfr new_Jinkela_buffer_3022 (
        .din(new_Jinkela_wire_4367),
        .dout(new_Jinkela_wire_4368)
    );

    bfr new_Jinkela_buffer_3070 (
        .din(new_Jinkela_wire_4425),
        .dout(new_Jinkela_wire_4426)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_2290),
        .dout(new_Jinkela_wire_2291)
    );

    bfr new_Jinkela_buffer_3023 (
        .din(new_Jinkela_wire_4368),
        .dout(new_Jinkela_wire_4369)
    );

    bfr new_Jinkela_buffer_3861 (
        .din(new_Jinkela_wire_5374),
        .dout(new_Jinkela_wire_5375)
    );

    bfr new_Jinkela_buffer_3840 (
        .din(new_Jinkela_wire_5347),
        .dout(new_Jinkela_wire_5348)
    );

    bfr new_Jinkela_buffer_3855 (
        .din(new_Jinkela_wire_5368),
        .dout(new_Jinkela_wire_5369)
    );

    bfr new_Jinkela_buffer_3841 (
        .din(new_Jinkela_wire_5348),
        .dout(new_Jinkela_wire_5349)
    );

    bfr new_Jinkela_buffer_3842 (
        .din(new_Jinkela_wire_5349),
        .dout(new_Jinkela_wire_5350)
    );

    bfr new_Jinkela_buffer_3856 (
        .din(new_Jinkela_wire_5369),
        .dout(new_Jinkela_wire_5370)
    );

    bfr new_Jinkela_buffer_3843 (
        .din(new_Jinkela_wire_5350),
        .dout(new_Jinkela_wire_5351)
    );

    bfr new_Jinkela_buffer_3862 (
        .din(new_Jinkela_wire_5375),
        .dout(new_Jinkela_wire_5376)
    );

    bfr new_Jinkela_buffer_3844 (
        .din(new_Jinkela_wire_5351),
        .dout(new_Jinkela_wire_5352)
    );

    bfr new_Jinkela_buffer_3857 (
        .din(new_Jinkela_wire_5370),
        .dout(new_Jinkela_wire_5371)
    );

    bfr new_Jinkela_buffer_3845 (
        .din(new_Jinkela_wire_5352),
        .dout(new_Jinkela_wire_5353)
    );

    bfr new_Jinkela_buffer_3880 (
        .din(_1064_),
        .dout(new_Jinkela_wire_5398)
    );

    bfr new_Jinkela_buffer_3846 (
        .din(new_Jinkela_wire_5353),
        .dout(new_Jinkela_wire_5354)
    );

    bfr new_Jinkela_buffer_3863 (
        .din(new_Jinkela_wire_5376),
        .dout(new_Jinkela_wire_5377)
    );

    bfr new_Jinkela_buffer_3847 (
        .din(new_Jinkela_wire_5354),
        .dout(new_Jinkela_wire_5355)
    );

    bfr new_Jinkela_buffer_3879 (
        .din(new_Jinkela_wire_5396),
        .dout(new_Jinkela_wire_5397)
    );

    bfr new_Jinkela_buffer_3848 (
        .din(new_Jinkela_wire_5355),
        .dout(new_Jinkela_wire_5356)
    );

    bfr new_Jinkela_buffer_3864 (
        .din(new_Jinkela_wire_5377),
        .dout(new_Jinkela_wire_5378)
    );

    bfr new_Jinkela_buffer_3849 (
        .din(new_Jinkela_wire_5356),
        .dout(new_Jinkela_wire_5357)
    );

    spl2 new_Jinkela_splitter_580 (
        .a(_0683_),
        .b(new_Jinkela_wire_5404),
        .c(new_Jinkela_wire_5405)
    );

    bfr new_Jinkela_buffer_3865 (
        .din(new_Jinkela_wire_5378),
        .dout(new_Jinkela_wire_5379)
    );

    bfr new_Jinkela_buffer_3894 (
        .din(_0857_),
        .dout(new_Jinkela_wire_5416)
    );

    bfr new_Jinkela_buffer_3881 (
        .din(new_Jinkela_wire_5398),
        .dout(new_Jinkela_wire_5399)
    );

    bfr new_Jinkela_buffer_3866 (
        .din(new_Jinkela_wire_5379),
        .dout(new_Jinkela_wire_5380)
    );

    bfr new_Jinkela_buffer_3867 (
        .din(new_Jinkela_wire_5380),
        .dout(new_Jinkela_wire_5381)
    );

    bfr new_Jinkela_buffer_3882 (
        .din(new_Jinkela_wire_5399),
        .dout(new_Jinkela_wire_5400)
    );

    bfr new_Jinkela_buffer_3868 (
        .din(new_Jinkela_wire_5381),
        .dout(new_Jinkela_wire_5382)
    );

    bfr new_Jinkela_buffer_3884 (
        .din(new_Jinkela_wire_5405),
        .dout(new_Jinkela_wire_5406)
    );

    bfr new_Jinkela_buffer_3869 (
        .din(new_Jinkela_wire_5382),
        .dout(new_Jinkela_wire_5383)
    );

    spl2 new_Jinkela_splitter_581 (
        .a(_0186_),
        .b(new_Jinkela_wire_5421),
        .c(new_Jinkela_wire_5422)
    );

    bfr new_Jinkela_buffer_3883 (
        .din(new_Jinkela_wire_5400),
        .dout(new_Jinkela_wire_5401)
    );

    bfr new_Jinkela_buffer_3870 (
        .din(new_Jinkela_wire_5383),
        .dout(new_Jinkela_wire_5384)
    );

    bfr new_Jinkela_buffer_3899 (
        .din(_0425_),
        .dout(new_Jinkela_wire_5423)
    );

    bfr new_Jinkela_buffer_3871 (
        .din(new_Jinkela_wire_5384),
        .dout(new_Jinkela_wire_5385)
    );

    bfr new_Jinkela_buffer_3895 (
        .din(new_Jinkela_wire_5416),
        .dout(new_Jinkela_wire_5417)
    );

    spl2 new_Jinkela_splitter_579 (
        .a(new_Jinkela_wire_5401),
        .b(new_Jinkela_wire_5402),
        .c(new_Jinkela_wire_5403)
    );

    bfr new_Jinkela_buffer_3872 (
        .din(new_Jinkela_wire_5385),
        .dout(new_Jinkela_wire_5386)
    );

    bfr new_Jinkela_buffer_3873 (
        .din(new_Jinkela_wire_5386),
        .dout(new_Jinkela_wire_5387)
    );

    bfr new_Jinkela_buffer_3885 (
        .din(new_Jinkela_wire_5406),
        .dout(new_Jinkela_wire_5407)
    );

    bfr new_Jinkela_buffer_3874 (
        .din(new_Jinkela_wire_5387),
        .dout(new_Jinkela_wire_5388)
    );

    bfr new_Jinkela_buffer_3886 (
        .din(new_Jinkela_wire_5407),
        .dout(new_Jinkela_wire_5408)
    );

    bfr new_Jinkela_buffer_3875 (
        .din(new_Jinkela_wire_5388),
        .dout(new_Jinkela_wire_5389)
    );

    and_bi _1697_ (
        .a(new_Jinkela_wire_1023),
        .b(new_Jinkela_wire_6694),
        .c(_0989_)
    );

    and_bi _2411_ (
        .a(_0408_),
        .b(new_Jinkela_wire_2304),
        .c(_0412_)
    );

    and_bi _1698_ (
        .a(new_Jinkela_wire_1903),
        .b(new_Jinkela_wire_1632),
        .c(_0990_)
    );

    and_bi _2412_ (
        .a(new_Jinkela_wire_677),
        .b(_0412_),
        .c(new_net_2431)
    );

    and_bi _1699_ (
        .a(new_Jinkela_wire_6116),
        .b(_0990_),
        .c(_0991_)
    );

    and_bi _2413_ (
        .a(new_Jinkela_wire_5881),
        .b(new_Jinkela_wire_808),
        .c(_0413_)
    );

    or_bb _1700_ (
        .a(new_Jinkela_wire_5156),
        .b(new_Jinkela_wire_6064),
        .c(_0992_)
    );

    and_bi _2414_ (
        .a(new_Jinkela_wire_4051),
        .b(new_Jinkela_wire_6830),
        .c(_0414_)
    );

    and_bb _1701_ (
        .a(new_Jinkela_wire_5157),
        .b(new_Jinkela_wire_6063),
        .c(_0993_)
    );

    or_bb _2415_ (
        .a(_0414_),
        .b(new_Jinkela_wire_5581),
        .c(_0415_)
    );

    and_bi _1702_ (
        .a(_0992_),
        .b(_0993_),
        .c(_0994_)
    );

    or_bb _2416_ (
        .a(new_Jinkela_wire_7850),
        .b(_0413_),
        .c(_0416_)
    );

    or_bb _1703_ (
        .a(new_Jinkela_wire_4411),
        .b(new_Jinkela_wire_1097),
        .c(_0995_)
    );

    and_bi _2417_ (
        .a(new_Jinkela_wire_520),
        .b(new_Jinkela_wire_3378),
        .c(_0417_)
    );

    or_bb _1704_ (
        .a(new_Jinkela_wire_1334),
        .b(new_Jinkela_wire_323),
        .c(_0996_)
    );

    and_bi _2418_ (
        .a(new_Jinkela_wire_718),
        .b(new_Jinkela_wire_4027),
        .c(_0418_)
    );

    and_bi _1705_ (
        .a(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_216),
        .c(_0997_)
    );

    or_bb _2419_ (
        .a(_0418_),
        .b(_0417_),
        .c(_0419_)
    );

    and_bi _1706_ (
        .a(_0996_),
        .b(_0997_),
        .c(_0998_)
    );

    and_bi _2420_ (
        .a(_0416_),
        .b(new_Jinkela_wire_2117),
        .c(_0420_)
    );

    or_bb _1707_ (
        .a(_0998_),
        .b(new_Jinkela_wire_2856),
        .c(_0999_)
    );

    and_bi _2421_ (
        .a(new_Jinkela_wire_678),
        .b(_0420_),
        .c(new_net_2471)
    );

    or_ii _1708_ (
        .a(new_Jinkela_wire_1591),
        .b(new_Jinkela_wire_1336),
        .c(_1000_)
    );

    or_ii _2422_ (
        .a(new_Jinkela_wire_7790),
        .b(new_Jinkela_wire_1521),
        .c(_0421_)
    );

    and_bi _1709_ (
        .a(new_Jinkela_wire_1286),
        .b(new_Jinkela_wire_1328),
        .c(_1001_)
    );

    and_ii _2423_ (
        .a(new_Jinkela_wire_2766),
        .b(new_Jinkela_wire_113),
        .c(_0422_)
    );

    and_bi _1710_ (
        .a(_1000_),
        .b(_1001_),
        .c(_1002_)
    );

    and_bb _2424_ (
        .a(new_Jinkela_wire_2765),
        .b(new_Jinkela_wire_114),
        .c(_0423_)
    );

    and_bi _1711_ (
        .a(new_Jinkela_wire_2857),
        .b(_1002_),
        .c(_1003_)
    );

    and_ii _2425_ (
        .a(_0423_),
        .b(_0422_),
        .c(_0424_)
    );

    and_bi _1712_ (
        .a(_0999_),
        .b(_1003_),
        .c(_1004_)
    );

    and_bi _2426_ (
        .a(new_Jinkela_wire_7130),
        .b(new_Jinkela_wire_1517),
        .c(_0425_)
    );

    and_bi _1713_ (
        .a(new_Jinkela_wire_1047),
        .b(new_Jinkela_wire_7848),
        .c(_1005_)
    );

    and_bi _2427_ (
        .a(_0421_),
        .b(new_Jinkela_wire_5425),
        .c(_0426_)
    );

    or_bb _1714_ (
        .a(_1005_),
        .b(new_Jinkela_wire_4843),
        .c(_1006_)
    );

    and_bi _2428_ (
        .a(new_Jinkela_wire_640),
        .b(_0426_),
        .c(_0427_)
    );

    and_bi _1715_ (
        .a(_0995_),
        .b(new_Jinkela_wire_4528),
        .c(_1007_)
    );

    or_ii _2429_ (
        .a(G178),
        .b(G62),
        .c(_0428_)
    );

    and_ii _1716_ (
        .a(_1007_),
        .b(new_Jinkela_wire_4453),
        .c(new_net_20)
    );

    or_bi _2430_ (
        .a(new_Jinkela_wire_299),
        .b(new_Jinkela_wire_1507),
        .c(_0429_)
    );

    and_bi _1717_ (
        .a(new_Jinkela_wire_1298),
        .b(new_Jinkela_wire_6689),
        .c(_1008_)
    );

    and_ii _2431_ (
        .a(new_Jinkela_wire_2420),
        .b(new_Jinkela_wire_1513),
        .c(_0430_)
    );

    and_bi _1718_ (
        .a(new_Jinkela_wire_5270),
        .b(new_Jinkela_wire_1626),
        .c(_1009_)
    );

    and_bi _2432_ (
        .a(new_Jinkela_wire_2270),
        .b(_0430_),
        .c(_0431_)
    );

    and_bb _1719_ (
        .a(new_Jinkela_wire_1629),
        .b(new_Jinkela_wire_2923),
        .c(_1010_)
    );

    or_bb _2433_ (
        .a(_0431_),
        .b(new_Jinkela_wire_633),
        .c(_0432_)
    );

    and_ii _1720_ (
        .a(_1010_),
        .b(_1009_),
        .c(_1011_)
    );

    or_ii _2434_ (
        .a(_0432_),
        .b(new_Jinkela_wire_4864),
        .c(_0433_)
    );

    or_bb _1721_ (
        .a(new_Jinkela_wire_3061),
        .b(new_Jinkela_wire_7035),
        .c(_1012_)
    );

    and_ii _2435_ (
        .a(new_Jinkela_wire_5432),
        .b(_0427_),
        .c(new_net_2485)
    );

    or_bi _1722_ (
        .a(new_Jinkela_wire_6379),
        .b(new_Jinkela_wire_3089),
        .c(_1013_)
    );

    and_bi _2436_ (
        .a(new_Jinkela_wire_7789),
        .b(new_Jinkela_wire_7135),
        .c(_0434_)
    );

    and_bi _1723_ (
        .a(new_Jinkela_wire_3062),
        .b(new_Jinkela_wire_6042),
        .c(_1014_)
    );

    and_bi _2437_ (
        .a(new_Jinkela_wire_7134),
        .b(new_Jinkela_wire_7787),
        .c(_0435_)
    );

    and_bi _1724_ (
        .a(_1012_),
        .b(_1014_),
        .c(_1015_)
    );

    or_bb _2438_ (
        .a(_0435_),
        .b(_0434_),
        .c(new_net_2377)
    );

    or_bb _1725_ (
        .a(new_Jinkela_wire_6250),
        .b(new_Jinkela_wire_1098),
        .c(_1016_)
    );

    or_ii _2439_ (
        .a(new_Jinkela_wire_1136),
        .b(new_Jinkela_wire_89),
        .c(_0436_)
    );

    or_bb _1726_ (
        .a(new_Jinkela_wire_567),
        .b(new_Jinkela_wire_324),
        .c(_1017_)
    );

    and_ii _2440_ (
        .a(_0436_),
        .b(new_Jinkela_wire_7741),
        .c(_0437_)
    );

    and_bi _1727_ (
        .a(new_Jinkela_wire_562),
        .b(new_Jinkela_wire_212),
        .c(_1018_)
    );

    and_bb _2441_ (
        .a(_0437_),
        .b(new_Jinkela_wire_2356),
        .c(_0438_)
    );

    and_bi _1728_ (
        .a(_1017_),
        .b(_1018_),
        .c(_1019_)
    );

    or_ii _2442_ (
        .a(new_Jinkela_wire_6374),
        .b(new_Jinkela_wire_4079),
        .c(_0439_)
    );

    and_bi _1729_ (
        .a(new_Jinkela_wire_1143),
        .b(_1019_),
        .c(_1020_)
    );

    or_bb _2443_ (
        .a(_0439_),
        .b(new_Jinkela_wire_5130),
        .c(_0440_)
    );

    or_ii _1730_ (
        .a(new_Jinkela_wire_1589),
        .b(new_Jinkela_wire_559),
        .c(_1021_)
    );

    or_bb _2444_ (
        .a(new_Jinkela_wire_3582),
        .b(new_Jinkela_wire_5422),
        .c(_0441_)
    );

    and_bi _1731_ (
        .a(new_Jinkela_wire_1287),
        .b(new_Jinkela_wire_560),
        .c(_1022_)
    );

    and_bi _2445_ (
        .a(new_Jinkela_wire_2781),
        .b(_0441_),
        .c(new_net_2423)
    );

    and_bi _1732_ (
        .a(_1021_),
        .b(_1022_),
        .c(_1023_)
    );

    or_bi _2446_ (
        .a(new_Jinkela_wire_396),
        .b(new_Jinkela_wire_3616),
        .c(_0442_)
    );

    and_bi _1733_ (
        .a(new_Jinkela_wire_3573),
        .b(_1023_),
        .c(_1024_)
    );

    and_bb _2447_ (
        .a(new_Jinkela_wire_5000),
        .b(new_Jinkela_wire_361),
        .c(_0443_)
    );

    and_ii _1734_ (
        .a(_1024_),
        .b(_1020_),
        .c(_1025_)
    );

    or_bb _2448_ (
        .a(_0443_),
        .b(new_Jinkela_wire_3960),
        .c(_0444_)
    );

    and_bi _1735_ (
        .a(new_Jinkela_wire_1050),
        .b(new_Jinkela_wire_3390),
        .c(_1026_)
    );

    and_bi _2449_ (
        .a(_0442_),
        .b(new_Jinkela_wire_6091),
        .c(_0445_)
    );

    or_bb _1736_ (
        .a(_1026_),
        .b(new_Jinkela_wire_4837),
        .c(_1027_)
    );

    and_bi _2450_ (
        .a(new_Jinkela_wire_1270),
        .b(new_Jinkela_wire_7872),
        .c(_0446_)
    );

    and_bi _1737_ (
        .a(_1016_),
        .b(new_Jinkela_wire_6584),
        .c(_1028_)
    );

    and_bi _2451_ (
        .a(new_Jinkela_wire_252),
        .b(new_Jinkela_wire_5803),
        .c(_0447_)
    );

    and_ii _1738_ (
        .a(_1028_),
        .b(new_Jinkela_wire_4154),
        .c(new_net_21)
    );

    or_bb _2452_ (
        .a(_0447_),
        .b(_0446_),
        .c(_0448_)
    );

    bfr new_Jinkela_buffer_5244 (
        .din(new_Jinkela_wire_7150),
        .dout(new_Jinkela_wire_7151)
    );

    bfr new_Jinkela_buffer_5247 (
        .din(new_Jinkela_wire_7153),
        .dout(new_Jinkela_wire_7154)
    );

    bfr new_Jinkela_buffer_5279 (
        .din(_1241_),
        .dout(new_Jinkela_wire_7191)
    );

    bfr new_Jinkela_buffer_5248 (
        .din(new_Jinkela_wire_7154),
        .dout(new_Jinkela_wire_7155)
    );

    bfr new_Jinkela_buffer_5280 (
        .din(new_Jinkela_wire_7191),
        .dout(new_Jinkela_wire_7192)
    );

    spl3L new_Jinkela_splitter_735 (
        .a(new_Jinkela_wire_7185),
        .d(new_Jinkela_wire_7186),
        .b(new_Jinkela_wire_7187),
        .c(new_Jinkela_wire_7188)
    );

    bfr new_Jinkela_buffer_5249 (
        .din(new_Jinkela_wire_7155),
        .dout(new_Jinkela_wire_7156)
    );

    bfr new_Jinkela_buffer_5278 (
        .din(new_Jinkela_wire_7184),
        .dout(new_Jinkela_wire_7185)
    );

    bfr new_Jinkela_buffer_5250 (
        .din(new_Jinkela_wire_7156),
        .dout(new_Jinkela_wire_7157)
    );

    bfr new_Jinkela_buffer_5251 (
        .din(new_Jinkela_wire_7157),
        .dout(new_Jinkela_wire_7158)
    );

    bfr new_Jinkela_buffer_5285 (
        .din(_1232_),
        .dout(new_Jinkela_wire_7197)
    );

    bfr new_Jinkela_buffer_5252 (
        .din(new_Jinkela_wire_7158),
        .dout(new_Jinkela_wire_7159)
    );

    bfr new_Jinkela_buffer_5286 (
        .din(_0463_),
        .dout(new_Jinkela_wire_7198)
    );

    bfr new_Jinkela_buffer_5253 (
        .din(new_Jinkela_wire_7159),
        .dout(new_Jinkela_wire_7160)
    );

    bfr new_Jinkela_buffer_5281 (
        .din(new_Jinkela_wire_7192),
        .dout(new_Jinkela_wire_7193)
    );

    bfr new_Jinkela_buffer_5254 (
        .din(new_Jinkela_wire_7160),
        .dout(new_Jinkela_wire_7161)
    );

    spl2 new_Jinkela_splitter_737 (
        .a(_1090_),
        .b(new_Jinkela_wire_7200),
        .c(new_Jinkela_wire_7201)
    );

    spl2 new_Jinkela_splitter_738 (
        .a(_0956_),
        .b(new_Jinkela_wire_7204),
        .c(new_Jinkela_wire_7205)
    );

    bfr new_Jinkela_buffer_5255 (
        .din(new_Jinkela_wire_7161),
        .dout(new_Jinkela_wire_7162)
    );

    bfr new_Jinkela_buffer_5282 (
        .din(new_Jinkela_wire_7193),
        .dout(new_Jinkela_wire_7194)
    );

    bfr new_Jinkela_buffer_5256 (
        .din(new_Jinkela_wire_7162),
        .dout(new_Jinkela_wire_7163)
    );

    bfr new_Jinkela_buffer_5287 (
        .din(new_Jinkela_wire_7198),
        .dout(new_Jinkela_wire_7199)
    );

    bfr new_Jinkela_buffer_5257 (
        .din(new_Jinkela_wire_7163),
        .dout(new_Jinkela_wire_7164)
    );

    bfr new_Jinkela_buffer_5283 (
        .din(new_Jinkela_wire_7194),
        .dout(new_Jinkela_wire_7195)
    );

    bfr new_Jinkela_buffer_5258 (
        .din(new_Jinkela_wire_7164),
        .dout(new_Jinkela_wire_7165)
    );

    bfr new_Jinkela_buffer_5288 (
        .din(new_Jinkela_wire_7201),
        .dout(new_Jinkela_wire_7202)
    );

    bfr new_Jinkela_buffer_5259 (
        .din(new_Jinkela_wire_7165),
        .dout(new_Jinkela_wire_7166)
    );

    bfr new_Jinkela_buffer_5284 (
        .din(new_Jinkela_wire_7195),
        .dout(new_Jinkela_wire_7196)
    );

    bfr new_Jinkela_buffer_5260 (
        .din(new_Jinkela_wire_7166),
        .dout(new_Jinkela_wire_7167)
    );

    bfr new_Jinkela_buffer_5261 (
        .din(new_Jinkela_wire_7167),
        .dout(new_Jinkela_wire_7168)
    );

    spl3L new_Jinkela_splitter_739 (
        .a(_0640_),
        .d(new_Jinkela_wire_7206),
        .b(new_Jinkela_wire_7207),
        .c(new_Jinkela_wire_7208)
    );

    bfr new_Jinkela_buffer_5262 (
        .din(new_Jinkela_wire_7168),
        .dout(new_Jinkela_wire_7169)
    );

    bfr new_Jinkela_buffer_5290 (
        .din(_0342_),
        .dout(new_Jinkela_wire_7213)
    );

    bfr new_Jinkela_buffer_5289 (
        .din(new_Jinkela_wire_7202),
        .dout(new_Jinkela_wire_7203)
    );

    bfr new_Jinkela_buffer_5263 (
        .din(new_Jinkela_wire_7169),
        .dout(new_Jinkela_wire_7170)
    );

    bfr new_Jinkela_buffer_5291 (
        .din(new_Jinkela_wire_7213),
        .dout(new_Jinkela_wire_7214)
    );

    bfr new_Jinkela_buffer_5264 (
        .din(new_Jinkela_wire_7170),
        .dout(new_Jinkela_wire_7171)
    );

    bfr new_Jinkela_buffer_5313 (
        .din(new_net_2455),
        .dout(new_Jinkela_wire_7240)
    );

    bfr new_Jinkela_buffer_5265 (
        .din(new_Jinkela_wire_7171),
        .dout(new_Jinkela_wire_7172)
    );

    spl2 new_Jinkela_splitter_740 (
        .a(new_Jinkela_wire_7208),
        .b(new_Jinkela_wire_7209),
        .c(new_Jinkela_wire_7210)
    );

    spl4L new_Jinkela_splitter_742 (
        .a(_0703_),
        .d(new_Jinkela_wire_7236),
        .e(new_Jinkela_wire_7237),
        .b(new_Jinkela_wire_7238),
        .c(new_Jinkela_wire_7239)
    );

    bfr new_Jinkela_buffer_5266 (
        .din(new_Jinkela_wire_7172),
        .dout(new_Jinkela_wire_7173)
    );

    bfr new_Jinkela_buffer_2270 (
        .din(new_Jinkela_wire_3458),
        .dout(new_Jinkela_wire_3459)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(new_net_2387),
        .dout(new_Jinkela_wire_2271)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(new_Jinkela_wire_2183),
        .dout(new_Jinkela_wire_2184)
    );

    bfr new_Jinkela_buffer_2271 (
        .din(new_Jinkela_wire_3459),
        .dout(new_Jinkela_wire_3460)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_2218),
        .dout(new_Jinkela_wire_2219)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_2184),
        .dout(new_Jinkela_wire_2185)
    );

    spl2 new_Jinkela_splitter_458 (
        .a(new_Jinkela_wire_3531),
        .b(new_Jinkela_wire_3532),
        .c(new_Jinkela_wire_3533)
    );

    bfr new_Jinkela_buffer_2272 (
        .din(new_Jinkela_wire_3460),
        .dout(new_Jinkela_wire_3461)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_2249),
        .dout(new_Jinkela_wire_2250)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(new_Jinkela_wire_2185),
        .dout(new_Jinkela_wire_2186)
    );

    bfr new_Jinkela_buffer_2320 (
        .din(new_Jinkela_wire_3540),
        .dout(new_Jinkela_wire_3541)
    );

    spl2 new_Jinkela_splitter_445 (
        .a(new_Jinkela_wire_3461),
        .b(new_Jinkela_wire_3462),
        .c(new_Jinkela_wire_3463)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(new_Jinkela_wire_2219),
        .dout(new_Jinkela_wire_2220)
    );

    bfr new_Jinkela_buffer_2273 (
        .din(new_Jinkela_wire_3463),
        .dout(new_Jinkela_wire_3464)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_2186),
        .dout(new_Jinkela_wire_2187)
    );

    bfr new_Jinkela_buffer_2296 (
        .din(new_Jinkela_wire_3488),
        .dout(new_Jinkela_wire_3489)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_2266),
        .dout(new_Jinkela_wire_2267)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_2187),
        .dout(new_Jinkela_wire_2188)
    );

    bfr new_Jinkela_buffer_2295 (
        .din(new_Jinkela_wire_3487),
        .dout(new_Jinkela_wire_3488)
    );

    bfr new_Jinkela_buffer_2297 (
        .din(new_Jinkela_wire_3489),
        .dout(new_Jinkela_wire_3490)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_2220),
        .dout(new_Jinkela_wire_2221)
    );

    bfr new_Jinkela_buffer_2356 (
        .din(_0440_),
        .dout(new_Jinkela_wire_3580)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_2188),
        .dout(new_Jinkela_wire_2189)
    );

    bfr new_Jinkela_buffer_2294 (
        .din(new_Jinkela_wire_3486),
        .dout(new_Jinkela_wire_3487)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(new_Jinkela_wire_2250),
        .dout(new_Jinkela_wire_2251)
    );

    bfr new_Jinkela_buffer_2298 (
        .din(new_Jinkela_wire_3490),
        .dout(new_Jinkela_wire_3491)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(new_Jinkela_wire_2189),
        .dout(new_Jinkela_wire_2190)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_2221),
        .dout(new_Jinkela_wire_2222)
    );

    bfr new_Jinkela_buffer_2321 (
        .din(new_Jinkela_wire_3541),
        .dout(new_Jinkela_wire_3542)
    );

    bfr new_Jinkela_buffer_2299 (
        .din(new_Jinkela_wire_3491),
        .dout(new_Jinkela_wire_3492)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_2190),
        .dout(new_Jinkela_wire_2191)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(_0411_),
        .dout(new_Jinkela_wire_2282)
    );

    spl2 new_Jinkela_splitter_447 (
        .a(new_Jinkela_wire_3492),
        .b(new_Jinkela_wire_3493),
        .c(new_Jinkela_wire_3494)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(new_Jinkela_wire_2191),
        .dout(new_Jinkela_wire_2192)
    );

    bfr new_Jinkela_buffer_2300 (
        .din(new_Jinkela_wire_3494),
        .dout(new_Jinkela_wire_3495)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(new_Jinkela_wire_2222),
        .dout(new_Jinkela_wire_2223)
    );

    spl3L new_Jinkela_splitter_460 (
        .a(new_Jinkela_wire_3572),
        .d(new_Jinkela_wire_3573),
        .b(new_Jinkela_wire_3574),
        .c(new_Jinkela_wire_3575)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_2192),
        .dout(new_Jinkela_wire_2193)
    );

    bfr new_Jinkela_buffer_2322 (
        .din(new_Jinkela_wire_3542),
        .dout(new_Jinkela_wire_3543)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_2251),
        .dout(new_Jinkela_wire_2252)
    );

    bfr new_Jinkela_buffer_2354 (
        .din(new_Jinkela_wire_3577),
        .dout(new_Jinkela_wire_3578)
    );

    spl2 new_Jinkela_splitter_448 (
        .a(new_Jinkela_wire_3495),
        .b(new_Jinkela_wire_3496),
        .c(new_Jinkela_wire_3497)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_2193),
        .dout(new_Jinkela_wire_2194)
    );

    bfr new_Jinkela_buffer_2301 (
        .din(new_Jinkela_wire_3497),
        .dout(new_Jinkela_wire_3498)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_2223),
        .dout(new_Jinkela_wire_2224)
    );

    bfr new_Jinkela_buffer_2351 (
        .din(new_Jinkela_wire_3571),
        .dout(new_Jinkela_wire_3572)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_2194),
        .dout(new_Jinkela_wire_2195)
    );

    bfr new_Jinkela_buffer_2323 (
        .din(new_Jinkela_wire_3543),
        .dout(new_Jinkela_wire_3544)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_2267),
        .dout(new_Jinkela_wire_2268)
    );

    bfr new_Jinkela_buffer_2302 (
        .din(new_Jinkela_wire_3498),
        .dout(new_Jinkela_wire_3499)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_2195),
        .dout(new_Jinkela_wire_2196)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_2224),
        .dout(new_Jinkela_wire_2225)
    );

    bfr new_Jinkela_buffer_2324 (
        .din(new_Jinkela_wire_3544),
        .dout(new_Jinkela_wire_3545)
    );

    spl2 new_Jinkela_splitter_449 (
        .a(new_Jinkela_wire_3499),
        .b(new_Jinkela_wire_3500),
        .c(new_Jinkela_wire_3501)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_Jinkela_wire_2252),
        .dout(new_Jinkela_wire_2253)
    );

    bfr new_Jinkela_buffer_2303 (
        .din(new_Jinkela_wire_3501),
        .dout(new_Jinkela_wire_3502)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_2225),
        .dout(new_Jinkela_wire_2226)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(new_Jinkela_wire_2271),
        .dout(new_Jinkela_wire_2272)
    );

    bfr new_Jinkela_buffer_2359 (
        .din(_0663_),
        .dout(new_Jinkela_wire_3583)
    );

    bfr new_Jinkela_buffer_2352 (
        .din(new_Jinkela_wire_3575),
        .dout(new_Jinkela_wire_3576)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_2226),
        .dout(new_Jinkela_wire_2227)
    );

    bfr new_Jinkela_buffer_2325 (
        .din(new_Jinkela_wire_3545),
        .dout(new_Jinkela_wire_3546)
    );

    bfr new_Jinkela_buffer_2304 (
        .din(new_Jinkela_wire_3502),
        .dout(new_Jinkela_wire_3503)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_2253),
        .dout(new_Jinkela_wire_2254)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(new_Jinkela_wire_2227),
        .dout(new_Jinkela_wire_2228)
    );

    spl2 new_Jinkela_splitter_450 (
        .a(new_Jinkela_wire_3503),
        .b(new_Jinkela_wire_3504),
        .c(new_Jinkela_wire_3505)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_2268),
        .dout(new_Jinkela_wire_2269)
    );

    bfr new_Jinkela_buffer_2305 (
        .din(new_Jinkela_wire_3505),
        .dout(new_Jinkela_wire_3506)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(new_Jinkela_wire_2228),
        .dout(new_Jinkela_wire_2229)
    );

    bfr new_Jinkela_buffer_2361 (
        .din(_0328_),
        .dout(new_Jinkela_wire_3591)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(new_Jinkela_wire_2254),
        .dout(new_Jinkela_wire_2255)
    );

    bfr new_Jinkela_buffer_2326 (
        .din(new_Jinkela_wire_3546),
        .dout(new_Jinkela_wire_3547)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_2229),
        .dout(new_Jinkela_wire_2230)
    );

    bfr new_Jinkela_buffer_2355 (
        .din(new_Jinkela_wire_3578),
        .dout(new_Jinkela_wire_3579)
    );

    spl2 new_Jinkela_splitter_451 (
        .a(new_Jinkela_wire_3506),
        .b(new_Jinkela_wire_3507),
        .c(new_Jinkela_wire_3508)
    );

    spl2 new_Jinkela_splitter_357 (
        .a(_1085_),
        .b(new_Jinkela_wire_2305),
        .c(new_Jinkela_wire_2306)
    );

    spl2 new_Jinkela_splitter_358 (
        .a(_0846_),
        .b(new_Jinkela_wire_2307),
        .c(new_Jinkela_wire_2308)
    );

    bfr new_Jinkela_buffer_2306 (
        .din(new_Jinkela_wire_3508),
        .dout(new_Jinkela_wire_3509)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_2230),
        .dout(new_Jinkela_wire_2231)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(new_Jinkela_wire_2255),
        .dout(new_Jinkela_wire_2256)
    );

    bfr new_Jinkela_buffer_2327 (
        .din(new_Jinkela_wire_3547),
        .dout(new_Jinkela_wire_3548)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(new_Jinkela_wire_2231),
        .dout(new_Jinkela_wire_2232)
    );

    bfr new_Jinkela_buffer_2357 (
        .din(new_Jinkela_wire_3580),
        .dout(new_Jinkela_wire_3581)
    );

    spl2 new_Jinkela_splitter_452 (
        .a(new_Jinkela_wire_3509),
        .b(new_Jinkela_wire_3510),
        .c(new_Jinkela_wire_3511)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(new_Jinkela_wire_2269),
        .dout(new_Jinkela_wire_2270)
    );

    spl2 new_Jinkela_splitter_505 (
        .a(new_Jinkela_wire_4312),
        .b(new_Jinkela_wire_4313),
        .c(new_Jinkela_wire_4314)
    );

    bfr new_Jinkela_buffer_2926 (
        .din(new_Jinkela_wire_4251),
        .dout(new_Jinkela_wire_4252)
    );

    bfr new_Jinkela_buffer_2944 (
        .din(new_Jinkela_wire_4271),
        .dout(new_Jinkela_wire_4272)
    );

    bfr new_Jinkela_buffer_3876 (
        .din(new_Jinkela_wire_5389),
        .dout(new_Jinkela_wire_5390)
    );

    bfr new_Jinkela_buffer_2927 (
        .din(new_Jinkela_wire_4252),
        .dout(new_Jinkela_wire_4253)
    );

    bfr new_Jinkela_buffer_3896 (
        .din(new_Jinkela_wire_5417),
        .dout(new_Jinkela_wire_5418)
    );

    bfr new_Jinkela_buffer_3887 (
        .din(new_Jinkela_wire_5408),
        .dout(new_Jinkela_wire_5409)
    );

    bfr new_Jinkela_buffer_2960 (
        .din(new_Jinkela_wire_4287),
        .dout(new_Jinkela_wire_4288)
    );

    bfr new_Jinkela_buffer_2945 (
        .din(new_Jinkela_wire_4272),
        .dout(new_Jinkela_wire_4273)
    );

    bfr new_Jinkela_buffer_3900 (
        .din(new_Jinkela_wire_5423),
        .dout(new_Jinkela_wire_5424)
    );

    bfr new_Jinkela_buffer_3888 (
        .din(new_Jinkela_wire_5409),
        .dout(new_Jinkela_wire_5410)
    );

    bfr new_Jinkela_buffer_2946 (
        .din(new_Jinkela_wire_4273),
        .dout(new_Jinkela_wire_4274)
    );

    bfr new_Jinkela_buffer_3897 (
        .din(new_Jinkela_wire_5418),
        .dout(new_Jinkela_wire_5419)
    );

    bfr new_Jinkela_buffer_3889 (
        .din(new_Jinkela_wire_5410),
        .dout(new_Jinkela_wire_5411)
    );

    bfr new_Jinkela_buffer_2961 (
        .din(new_Jinkela_wire_4288),
        .dout(new_Jinkela_wire_4289)
    );

    bfr new_Jinkela_buffer_2947 (
        .din(new_Jinkela_wire_4274),
        .dout(new_Jinkela_wire_4275)
    );

    bfr new_Jinkela_buffer_3902 (
        .din(new_net_2363),
        .dout(new_Jinkela_wire_5426)
    );

    bfr new_Jinkela_buffer_3890 (
        .din(new_Jinkela_wire_5411),
        .dout(new_Jinkela_wire_5412)
    );

    bfr new_Jinkela_buffer_2994 (
        .din(new_Jinkela_wire_4325),
        .dout(new_Jinkela_wire_4326)
    );

    spl2 new_Jinkela_splitter_508 (
        .a(_0878_),
        .b(new_Jinkela_wire_4340),
        .c(new_Jinkela_wire_4341)
    );

    bfr new_Jinkela_buffer_2948 (
        .din(new_Jinkela_wire_4275),
        .dout(new_Jinkela_wire_4276)
    );

    bfr new_Jinkela_buffer_3898 (
        .din(new_Jinkela_wire_5419),
        .dout(new_Jinkela_wire_5420)
    );

    bfr new_Jinkela_buffer_3891 (
        .din(new_Jinkela_wire_5412),
        .dout(new_Jinkela_wire_5413)
    );

    bfr new_Jinkela_buffer_2962 (
        .din(new_Jinkela_wire_4289),
        .dout(new_Jinkela_wire_4290)
    );

    bfr new_Jinkela_buffer_2949 (
        .din(new_Jinkela_wire_4276),
        .dout(new_Jinkela_wire_4277)
    );

    bfr new_Jinkela_buffer_3904 (
        .din(_0433_),
        .dout(new_Jinkela_wire_5428)
    );

    bfr new_Jinkela_buffer_3892 (
        .din(new_Jinkela_wire_5413),
        .dout(new_Jinkela_wire_5414)
    );

    bfr new_Jinkela_buffer_2985 (
        .din(new_Jinkela_wire_4316),
        .dout(new_Jinkela_wire_4317)
    );

    bfr new_Jinkela_buffer_2950 (
        .din(new_Jinkela_wire_4277),
        .dout(new_Jinkela_wire_4278)
    );

    bfr new_Jinkela_buffer_3901 (
        .din(new_Jinkela_wire_5424),
        .dout(new_Jinkela_wire_5425)
    );

    bfr new_Jinkela_buffer_3893 (
        .din(new_Jinkela_wire_5414),
        .dout(new_Jinkela_wire_5415)
    );

    bfr new_Jinkela_buffer_2963 (
        .din(new_Jinkela_wire_4290),
        .dout(new_Jinkela_wire_4291)
    );

    bfr new_Jinkela_buffer_2951 (
        .din(new_Jinkela_wire_4278),
        .dout(new_Jinkela_wire_4279)
    );

    bfr new_Jinkela_buffer_3903 (
        .din(new_Jinkela_wire_5426),
        .dout(new_Jinkela_wire_5427)
    );

    bfr new_Jinkela_buffer_2986 (
        .din(new_Jinkela_wire_4317),
        .dout(new_Jinkela_wire_4318)
    );

    bfr new_Jinkela_buffer_3909 (
        .din(_0025_),
        .dout(new_Jinkela_wire_5433)
    );

    bfr new_Jinkela_buffer_2964 (
        .din(new_Jinkela_wire_4291),
        .dout(new_Jinkela_wire_4292)
    );

    bfr new_Jinkela_buffer_3905 (
        .din(new_Jinkela_wire_5428),
        .dout(new_Jinkela_wire_5429)
    );

    bfr new_Jinkela_buffer_3910 (
        .din(_0238_),
        .dout(new_Jinkela_wire_5434)
    );

    spl2 new_Jinkela_splitter_507 (
        .a(new_Jinkela_wire_4337),
        .b(new_Jinkela_wire_4338),
        .c(new_Jinkela_wire_4339)
    );

    bfr new_Jinkela_buffer_2965 (
        .din(new_Jinkela_wire_4292),
        .dout(new_Jinkela_wire_4293)
    );

    bfr new_Jinkela_buffer_3906 (
        .din(new_Jinkela_wire_5429),
        .dout(new_Jinkela_wire_5430)
    );

    bfr new_Jinkela_buffer_2987 (
        .din(new_Jinkela_wire_4318),
        .dout(new_Jinkela_wire_4319)
    );

    spl2 new_Jinkela_splitter_582 (
        .a(_0007_),
        .b(new_Jinkela_wire_5435),
        .c(new_Jinkela_wire_5436)
    );

    bfr new_Jinkela_buffer_3911 (
        .din(_0282_),
        .dout(new_Jinkela_wire_5437)
    );

    bfr new_Jinkela_buffer_2966 (
        .din(new_Jinkela_wire_4293),
        .dout(new_Jinkela_wire_4294)
    );

    bfr new_Jinkela_buffer_3907 (
        .din(new_Jinkela_wire_5430),
        .dout(new_Jinkela_wire_5431)
    );

    bfr new_Jinkela_buffer_2995 (
        .din(new_Jinkela_wire_4326),
        .dout(new_Jinkela_wire_4327)
    );

    bfr new_Jinkela_buffer_3912 (
        .din(new_Jinkela_wire_5437),
        .dout(new_Jinkela_wire_5438)
    );

    bfr new_Jinkela_buffer_2967 (
        .din(new_Jinkela_wire_4294),
        .dout(new_Jinkela_wire_4295)
    );

    bfr new_Jinkela_buffer_3908 (
        .din(new_Jinkela_wire_5431),
        .dout(new_Jinkela_wire_5432)
    );

    bfr new_Jinkela_buffer_2988 (
        .din(new_Jinkela_wire_4319),
        .dout(new_Jinkela_wire_4320)
    );

    bfr new_Jinkela_buffer_2968 (
        .din(new_Jinkela_wire_4295),
        .dout(new_Jinkela_wire_4296)
    );

    bfr new_Jinkela_buffer_3914 (
        .din(new_net_2511),
        .dout(new_Jinkela_wire_5440)
    );

    bfr new_Jinkela_buffer_3921 (
        .din(new_net_2435),
        .dout(new_Jinkela_wire_5447)
    );

    bfr new_Jinkela_buffer_2969 (
        .din(new_Jinkela_wire_4296),
        .dout(new_Jinkela_wire_4297)
    );

    bfr new_Jinkela_buffer_3913 (
        .din(new_Jinkela_wire_5438),
        .dout(new_Jinkela_wire_5439)
    );

    bfr new_Jinkela_buffer_2989 (
        .din(new_Jinkela_wire_4320),
        .dout(new_Jinkela_wire_4321)
    );

    bfr new_Jinkela_buffer_3915 (
        .din(new_Jinkela_wire_5440),
        .dout(new_Jinkela_wire_5441)
    );

    bfr new_Jinkela_buffer_2970 (
        .din(new_Jinkela_wire_4297),
        .dout(new_Jinkela_wire_4298)
    );

    bfr new_Jinkela_buffer_3961 (
        .din(_0324_),
        .dout(new_Jinkela_wire_5487)
    );

    bfr new_Jinkela_buffer_2996 (
        .din(new_Jinkela_wire_4327),
        .dout(new_Jinkela_wire_4328)
    );

    bfr new_Jinkela_buffer_3916 (
        .din(new_Jinkela_wire_5441),
        .dout(new_Jinkela_wire_5442)
    );

    bfr new_Jinkela_buffer_2971 (
        .din(new_Jinkela_wire_4298),
        .dout(new_Jinkela_wire_4299)
    );

    bfr new_Jinkela_buffer_3922 (
        .din(new_Jinkela_wire_5447),
        .dout(new_Jinkela_wire_5448)
    );

    bfr new_Jinkela_buffer_2990 (
        .din(new_Jinkela_wire_4321),
        .dout(new_Jinkela_wire_4322)
    );

    bfr new_Jinkela_buffer_3917 (
        .din(new_Jinkela_wire_5442),
        .dout(new_Jinkela_wire_5443)
    );

    bfr new_Jinkela_buffer_2972 (
        .din(new_Jinkela_wire_4299),
        .dout(new_Jinkela_wire_4300)
    );

    bfr new_Jinkela_buffer_3963 (
        .din(_0072_),
        .dout(new_Jinkela_wire_5489)
    );

    bfr new_Jinkela_buffer_3004 (
        .din(_0229_),
        .dout(new_Jinkela_wire_4342)
    );

    bfr new_Jinkela_buffer_3918 (
        .din(new_Jinkela_wire_5443),
        .dout(new_Jinkela_wire_5444)
    );

    bfr new_Jinkela_buffer_2973 (
        .din(new_Jinkela_wire_4300),
        .dout(new_Jinkela_wire_4301)
    );

    bfr new_Jinkela_buffer_3923 (
        .din(new_Jinkela_wire_5448),
        .dout(new_Jinkela_wire_5449)
    );

    bfr new_Jinkela_buffer_2991 (
        .din(new_Jinkela_wire_4322),
        .dout(new_Jinkela_wire_4323)
    );

    bfr new_Jinkela_buffer_3919 (
        .din(new_Jinkela_wire_5444),
        .dout(new_Jinkela_wire_5445)
    );

    bfr new_Jinkela_buffer_2974 (
        .din(new_Jinkela_wire_4301),
        .dout(new_Jinkela_wire_4302)
    );

    bfr new_Jinkela_buffer_3962 (
        .din(new_Jinkela_wire_5487),
        .dout(new_Jinkela_wire_5488)
    );

    bfr new_Jinkela_buffer_2997 (
        .din(new_Jinkela_wire_4328),
        .dout(new_Jinkela_wire_4329)
    );

    bfr new_Jinkela_buffer_3920 (
        .din(new_Jinkela_wire_5445),
        .dout(new_Jinkela_wire_5446)
    );

    bfr new_Jinkela_buffer_2975 (
        .din(new_Jinkela_wire_4302),
        .dout(new_Jinkela_wire_4303)
    );

    bfr new_Jinkela_buffer_3924 (
        .din(new_Jinkela_wire_5449),
        .dout(new_Jinkela_wire_5450)
    );

    bfr new_Jinkela_buffer_2992 (
        .din(new_Jinkela_wire_4323),
        .dout(new_Jinkela_wire_4324)
    );

    bfr new_Jinkela_buffer_3964 (
        .din(new_net_2491),
        .dout(new_Jinkela_wire_5490)
    );

    spl2 new_Jinkela_splitter_354 (
        .a(_0968_),
        .b(new_Jinkela_wire_2246),
        .c(new_Jinkela_wire_2247)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(new_Jinkela_wire_2142),
        .dout(new_Jinkela_wire_2143)
    );

    bfr new_Jinkela_buffer_2617 (
        .din(new_Jinkela_wire_3886),
        .dout(new_Jinkela_wire_3887)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(new_Jinkela_wire_2167),
        .dout(new_Jinkela_wire_2168)
    );

    bfr new_Jinkela_buffer_2588 (
        .din(new_Jinkela_wire_3855),
        .dout(new_Jinkela_wire_3856)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_2143),
        .dout(new_Jinkela_wire_2144)
    );

    bfr new_Jinkela_buffer_2697 (
        .din(new_Jinkela_wire_3986),
        .dout(new_Jinkela_wire_3987)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_2211),
        .dout(new_Jinkela_wire_2212)
    );

    bfr new_Jinkela_buffer_2589 (
        .din(new_Jinkela_wire_3856),
        .dout(new_Jinkela_wire_3857)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_2207),
        .dout(new_Jinkela_wire_2208)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(new_Jinkela_wire_2144),
        .dout(new_Jinkela_wire_2145)
    );

    bfr new_Jinkela_buffer_2624 (
        .din(new_Jinkela_wire_3893),
        .dout(new_Jinkela_wire_3894)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(new_Jinkela_wire_2168),
        .dout(new_Jinkela_wire_2169)
    );

    bfr new_Jinkela_buffer_2590 (
        .din(new_Jinkela_wire_3857),
        .dout(new_Jinkela_wire_3858)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_2145),
        .dout(new_Jinkela_wire_2146)
    );

    bfr new_Jinkela_buffer_2634 (
        .din(new_Jinkela_wire_3903),
        .dout(new_Jinkela_wire_3904)
    );

    bfr new_Jinkela_buffer_2591 (
        .din(new_Jinkela_wire_3858),
        .dout(new_Jinkela_wire_3859)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(new_Jinkela_wire_2146),
        .dout(new_Jinkela_wire_2147)
    );

    bfr new_Jinkela_buffer_2625 (
        .din(new_Jinkela_wire_3894),
        .dout(new_Jinkela_wire_3895)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(new_Jinkela_wire_2169),
        .dout(new_Jinkela_wire_2170)
    );

    bfr new_Jinkela_buffer_2592 (
        .din(new_Jinkela_wire_3859),
        .dout(new_Jinkela_wire_3860)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_Jinkela_wire_2147),
        .dout(new_Jinkela_wire_2148)
    );

    bfr new_Jinkela_buffer_2698 (
        .din(new_Jinkela_wire_3987),
        .dout(new_Jinkela_wire_3988)
    );

    spl2 new_Jinkela_splitter_353 (
        .a(_0950_),
        .b(new_Jinkela_wire_2244),
        .c(new_Jinkela_wire_2245)
    );

    bfr new_Jinkela_buffer_2593 (
        .din(new_Jinkela_wire_3860),
        .dout(new_Jinkela_wire_3861)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_2148),
        .dout(new_Jinkela_wire_2149)
    );

    bfr new_Jinkela_buffer_2626 (
        .din(new_Jinkela_wire_3895),
        .dout(new_Jinkela_wire_3896)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(new_Jinkela_wire_2170),
        .dout(new_Jinkela_wire_2171)
    );

    bfr new_Jinkela_buffer_2594 (
        .din(new_Jinkela_wire_3861),
        .dout(new_Jinkela_wire_3862)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_2149),
        .dout(new_Jinkela_wire_2150)
    );

    bfr new_Jinkela_buffer_2635 (
        .din(new_Jinkela_wire_3904),
        .dout(new_Jinkela_wire_3905)
    );

    bfr new_Jinkela_buffer_2595 (
        .din(new_Jinkela_wire_3862),
        .dout(new_Jinkela_wire_3863)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_2150),
        .dout(new_Jinkela_wire_2151)
    );

    bfr new_Jinkela_buffer_2627 (
        .din(new_Jinkela_wire_3896),
        .dout(new_Jinkela_wire_3897)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(new_Jinkela_wire_2171),
        .dout(new_Jinkela_wire_2172)
    );

    bfr new_Jinkela_buffer_2596 (
        .din(new_Jinkela_wire_3863),
        .dout(new_Jinkela_wire_3864)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_2151),
        .dout(new_Jinkela_wire_2152)
    );

    spl2 new_Jinkela_splitter_493 (
        .a(new_net_8),
        .b(new_Jinkela_wire_4050),
        .c(new_Jinkela_wire_4052)
    );

    spl3L new_Jinkela_splitter_489 (
        .a(_0105_),
        .d(new_Jinkela_wire_4021),
        .b(new_Jinkela_wire_4024),
        .c(new_Jinkela_wire_4029)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_2212),
        .dout(new_Jinkela_wire_2213)
    );

    bfr new_Jinkela_buffer_2597 (
        .din(new_Jinkela_wire_3864),
        .dout(new_Jinkela_wire_3865)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(new_Jinkela_wire_2152),
        .dout(new_Jinkela_wire_2153)
    );

    bfr new_Jinkela_buffer_2628 (
        .din(new_Jinkela_wire_3897),
        .dout(new_Jinkela_wire_3898)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_2172),
        .dout(new_Jinkela_wire_2173)
    );

    bfr new_Jinkela_buffer_2598 (
        .din(new_Jinkela_wire_3865),
        .dout(new_Jinkela_wire_3866)
    );

    bfr new_Jinkela_buffer_2636 (
        .din(new_Jinkela_wire_3905),
        .dout(new_Jinkela_wire_3906)
    );

    spl2 new_Jinkela_splitter_356 (
        .a(_1244_),
        .b(new_Jinkela_wire_2263),
        .c(new_Jinkela_wire_2264)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_2173),
        .dout(new_Jinkela_wire_2174)
    );

    bfr new_Jinkela_buffer_2599 (
        .din(new_Jinkela_wire_3866),
        .dout(new_Jinkela_wire_3867)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(new_Jinkela_wire_2213),
        .dout(new_Jinkela_wire_2214)
    );

    bfr new_Jinkela_buffer_2629 (
        .din(new_Jinkela_wire_3898),
        .dout(new_Jinkela_wire_3899)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_2174),
        .dout(new_Jinkela_wire_2175)
    );

    bfr new_Jinkela_buffer_2600 (
        .din(new_Jinkela_wire_3867),
        .dout(new_Jinkela_wire_3868)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(_0429_),
        .dout(new_Jinkela_wire_2266)
    );

    bfr new_Jinkela_buffer_2696 (
        .din(new_net_2459),
        .dout(new_Jinkela_wire_3986)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(new_Jinkela_wire_2175),
        .dout(new_Jinkela_wire_2176)
    );

    bfr new_Jinkela_buffer_2601 (
        .din(new_Jinkela_wire_3868),
        .dout(new_Jinkela_wire_3869)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(new_Jinkela_wire_2214),
        .dout(new_Jinkela_wire_2215)
    );

    bfr new_Jinkela_buffer_2630 (
        .din(new_Jinkela_wire_3899),
        .dout(new_Jinkela_wire_3900)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_2176),
        .dout(new_Jinkela_wire_2177)
    );

    bfr new_Jinkela_buffer_2602 (
        .din(new_Jinkela_wire_3869),
        .dout(new_Jinkela_wire_3870)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(new_Jinkela_wire_2247),
        .dout(new_Jinkela_wire_2248)
    );

    bfr new_Jinkela_buffer_2637 (
        .din(new_Jinkela_wire_3906),
        .dout(new_Jinkela_wire_3907)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(_0835_),
        .dout(new_Jinkela_wire_2265)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_2177),
        .dout(new_Jinkela_wire_2178)
    );

    bfr new_Jinkela_buffer_2603 (
        .din(new_Jinkela_wire_3870),
        .dout(new_Jinkela_wire_3871)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(new_Jinkela_wire_2215),
        .dout(new_Jinkela_wire_2216)
    );

    bfr new_Jinkela_buffer_2631 (
        .din(new_Jinkela_wire_3900),
        .dout(new_Jinkela_wire_3901)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_2178),
        .dout(new_Jinkela_wire_2179)
    );

    bfr new_Jinkela_buffer_2604 (
        .din(new_Jinkela_wire_3871),
        .dout(new_Jinkela_wire_3872)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(new_Jinkela_wire_2179),
        .dout(new_Jinkela_wire_2180)
    );

    bfr new_Jinkela_buffer_2605 (
        .din(new_Jinkela_wire_3872),
        .dout(new_Jinkela_wire_3873)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_2216),
        .dout(new_Jinkela_wire_2217)
    );

    bfr new_Jinkela_buffer_2638 (
        .din(new_Jinkela_wire_3907),
        .dout(new_Jinkela_wire_3908)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_2180),
        .dout(new_Jinkela_wire_2181)
    );

    bfr new_Jinkela_buffer_2606 (
        .din(new_Jinkela_wire_3873),
        .dout(new_Jinkela_wire_3874)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(new_Jinkela_wire_2248),
        .dout(new_Jinkela_wire_2249)
    );

    bfr new_Jinkela_buffer_2731 (
        .din(_0702_),
        .dout(new_Jinkela_wire_4034)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(new_Jinkela_wire_2181),
        .dout(new_Jinkela_wire_2182)
    );

    bfr new_Jinkela_buffer_2607 (
        .din(new_Jinkela_wire_3874),
        .dout(new_Jinkela_wire_3875)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_2217),
        .dout(new_Jinkela_wire_2218)
    );

    bfr new_Jinkela_buffer_2639 (
        .din(new_Jinkela_wire_3908),
        .dout(new_Jinkela_wire_3909)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(new_Jinkela_wire_2182),
        .dout(new_Jinkela_wire_2183)
    );

    bfr new_Jinkela_buffer_2608 (
        .din(new_Jinkela_wire_3875),
        .dout(new_Jinkela_wire_3876)
    );

    bfr new_Jinkela_buffer_2905 (
        .din(new_Jinkela_wire_4230),
        .dout(new_Jinkela_wire_4231)
    );

    bfr new_Jinkela_buffer_5191 (
        .din(new_Jinkela_wire_7069),
        .dout(new_Jinkela_wire_7070)
    );

    bfr new_Jinkela_buffer_2993 (
        .din(new_net_2437),
        .dout(new_Jinkela_wire_4325)
    );

    bfr new_Jinkela_buffer_5220 (
        .din(new_Jinkela_wire_7114),
        .dout(new_Jinkela_wire_7115)
    );

    bfr new_Jinkela_buffer_2906 (
        .din(new_Jinkela_wire_4231),
        .dout(new_Jinkela_wire_4232)
    );

    bfr new_Jinkela_buffer_5192 (
        .din(new_Jinkela_wire_7070),
        .dout(new_Jinkela_wire_7071)
    );

    bfr new_Jinkela_buffer_2934 (
        .din(new_Jinkela_wire_4261),
        .dout(new_Jinkela_wire_4262)
    );

    bfr new_Jinkela_buffer_5209 (
        .din(new_Jinkela_wire_7095),
        .dout(new_Jinkela_wire_7096)
    );

    bfr new_Jinkela_buffer_2907 (
        .din(new_Jinkela_wire_4232),
        .dout(new_Jinkela_wire_4233)
    );

    bfr new_Jinkela_buffer_5193 (
        .din(new_Jinkela_wire_7071),
        .dout(new_Jinkela_wire_7072)
    );

    bfr new_Jinkela_buffer_2955 (
        .din(new_Jinkela_wire_4282),
        .dout(new_Jinkela_wire_4283)
    );

    bfr new_Jinkela_buffer_2908 (
        .din(new_Jinkela_wire_4233),
        .dout(new_Jinkela_wire_4234)
    );

    bfr new_Jinkela_buffer_5194 (
        .din(new_Jinkela_wire_7072),
        .dout(new_Jinkela_wire_7073)
    );

    bfr new_Jinkela_buffer_2935 (
        .din(new_Jinkela_wire_4262),
        .dout(new_Jinkela_wire_4263)
    );

    bfr new_Jinkela_buffer_5210 (
        .din(new_Jinkela_wire_7096),
        .dout(new_Jinkela_wire_7097)
    );

    bfr new_Jinkela_buffer_2909 (
        .din(new_Jinkela_wire_4234),
        .dout(new_Jinkela_wire_4235)
    );

    bfr new_Jinkela_buffer_5221 (
        .din(new_Jinkela_wire_7115),
        .dout(new_Jinkela_wire_7116)
    );

    bfr new_Jinkela_buffer_5211 (
        .din(new_Jinkela_wire_7097),
        .dout(new_Jinkela_wire_7098)
    );

    bfr new_Jinkela_buffer_2981 (
        .din(new_Jinkela_wire_4310),
        .dout(new_Jinkela_wire_4311)
    );

    bfr new_Jinkela_buffer_2910 (
        .din(new_Jinkela_wire_4235),
        .dout(new_Jinkela_wire_4236)
    );

    spl2 new_Jinkela_splitter_733 (
        .a(_0906_),
        .b(new_Jinkela_wire_7143),
        .c(new_Jinkela_wire_7144)
    );

    bfr new_Jinkela_buffer_5236 (
        .din(new_Jinkela_wire_7136),
        .dout(new_Jinkela_wire_7137)
    );

    bfr new_Jinkela_buffer_2936 (
        .din(new_Jinkela_wire_4263),
        .dout(new_Jinkela_wire_4264)
    );

    bfr new_Jinkela_buffer_5212 (
        .din(new_Jinkela_wire_7098),
        .dout(new_Jinkela_wire_7099)
    );

    bfr new_Jinkela_buffer_2911 (
        .din(new_Jinkela_wire_4236),
        .dout(new_Jinkela_wire_4237)
    );

    bfr new_Jinkela_buffer_5222 (
        .din(new_Jinkela_wire_7116),
        .dout(new_Jinkela_wire_7117)
    );

    bfr new_Jinkela_buffer_2956 (
        .din(new_Jinkela_wire_4283),
        .dout(new_Jinkela_wire_4284)
    );

    bfr new_Jinkela_buffer_5213 (
        .din(new_Jinkela_wire_7099),
        .dout(new_Jinkela_wire_7100)
    );

    bfr new_Jinkela_buffer_2912 (
        .din(new_Jinkela_wire_4237),
        .dout(new_Jinkela_wire_4238)
    );

    bfr new_Jinkela_buffer_5234 (
        .din(new_Jinkela_wire_7132),
        .dout(new_Jinkela_wire_7133)
    );

    bfr new_Jinkela_buffer_2937 (
        .din(new_Jinkela_wire_4264),
        .dout(new_Jinkela_wire_4265)
    );

    bfr new_Jinkela_buffer_5214 (
        .din(new_Jinkela_wire_7100),
        .dout(new_Jinkela_wire_7101)
    );

    bfr new_Jinkela_buffer_2913 (
        .din(new_Jinkela_wire_4238),
        .dout(new_Jinkela_wire_4239)
    );

    bfr new_Jinkela_buffer_5223 (
        .din(new_Jinkela_wire_7117),
        .dout(new_Jinkela_wire_7118)
    );

    bfr new_Jinkela_buffer_5215 (
        .din(new_Jinkela_wire_7101),
        .dout(new_Jinkela_wire_7102)
    );

    bfr new_Jinkela_buffer_2914 (
        .din(new_Jinkela_wire_4239),
        .dout(new_Jinkela_wire_4240)
    );

    bfr new_Jinkela_buffer_5240 (
        .din(_0961_),
        .dout(new_Jinkela_wire_7147)
    );

    bfr new_Jinkela_buffer_2938 (
        .din(new_Jinkela_wire_4265),
        .dout(new_Jinkela_wire_4266)
    );

    bfr new_Jinkela_buffer_5216 (
        .din(new_Jinkela_wire_7102),
        .dout(new_Jinkela_wire_7103)
    );

    bfr new_Jinkela_buffer_2915 (
        .din(new_Jinkela_wire_4240),
        .dout(new_Jinkela_wire_4241)
    );

    bfr new_Jinkela_buffer_5224 (
        .din(new_Jinkela_wire_7118),
        .dout(new_Jinkela_wire_7119)
    );

    bfr new_Jinkela_buffer_2957 (
        .din(new_Jinkela_wire_4284),
        .dout(new_Jinkela_wire_4285)
    );

    bfr new_Jinkela_buffer_5217 (
        .din(new_Jinkela_wire_7103),
        .dout(new_Jinkela_wire_7104)
    );

    bfr new_Jinkela_buffer_2916 (
        .din(new_Jinkela_wire_4241),
        .dout(new_Jinkela_wire_4242)
    );

    spl2 new_Jinkela_splitter_731 (
        .a(new_Jinkela_wire_7133),
        .b(new_Jinkela_wire_7134),
        .c(new_Jinkela_wire_7135)
    );

    bfr new_Jinkela_buffer_2939 (
        .din(new_Jinkela_wire_4266),
        .dout(new_Jinkela_wire_4267)
    );

    bfr new_Jinkela_buffer_5225 (
        .din(new_Jinkela_wire_7119),
        .dout(new_Jinkela_wire_7120)
    );

    bfr new_Jinkela_buffer_2917 (
        .din(new_Jinkela_wire_4242),
        .dout(new_Jinkela_wire_4243)
    );

    spl2 new_Jinkela_splitter_734 (
        .a(new_Jinkela_wire_7144),
        .b(new_Jinkela_wire_7145),
        .c(new_Jinkela_wire_7146)
    );

    bfr new_Jinkela_buffer_2984 (
        .din(new_Jinkela_wire_4315),
        .dout(new_Jinkela_wire_4316)
    );

    bfr new_Jinkela_buffer_5226 (
        .din(new_Jinkela_wire_7120),
        .dout(new_Jinkela_wire_7121)
    );

    bfr new_Jinkela_buffer_2982 (
        .din(new_Jinkela_wire_4311),
        .dout(new_Jinkela_wire_4312)
    );

    bfr new_Jinkela_buffer_2918 (
        .din(new_Jinkela_wire_4243),
        .dout(new_Jinkela_wire_4244)
    );

    bfr new_Jinkela_buffer_5238 (
        .din(new_Jinkela_wire_7140),
        .dout(new_Jinkela_wire_7141)
    );

    spl2 new_Jinkela_splitter_732 (
        .a(new_Jinkela_wire_7137),
        .b(new_Jinkela_wire_7138),
        .c(new_Jinkela_wire_7139)
    );

    bfr new_Jinkela_buffer_2940 (
        .din(new_Jinkela_wire_4267),
        .dout(new_Jinkela_wire_4268)
    );

    bfr new_Jinkela_buffer_5227 (
        .din(new_Jinkela_wire_7121),
        .dout(new_Jinkela_wire_7122)
    );

    bfr new_Jinkela_buffer_2919 (
        .din(new_Jinkela_wire_4244),
        .dout(new_Jinkela_wire_4245)
    );

    bfr new_Jinkela_buffer_5239 (
        .din(new_Jinkela_wire_7141),
        .dout(new_Jinkela_wire_7142)
    );

    bfr new_Jinkela_buffer_2958 (
        .din(new_Jinkela_wire_4285),
        .dout(new_Jinkela_wire_4286)
    );

    bfr new_Jinkela_buffer_5228 (
        .din(new_Jinkela_wire_7122),
        .dout(new_Jinkela_wire_7123)
    );

    bfr new_Jinkela_buffer_2920 (
        .din(new_Jinkela_wire_4245),
        .dout(new_Jinkela_wire_4246)
    );

    bfr new_Jinkela_buffer_2941 (
        .din(new_Jinkela_wire_4268),
        .dout(new_Jinkela_wire_4269)
    );

    bfr new_Jinkela_buffer_5229 (
        .din(new_Jinkela_wire_7123),
        .dout(new_Jinkela_wire_7124)
    );

    bfr new_Jinkela_buffer_2921 (
        .din(new_Jinkela_wire_4246),
        .dout(new_Jinkela_wire_4247)
    );

    bfr new_Jinkela_buffer_5245 (
        .din(_0552_),
        .dout(new_Jinkela_wire_7152)
    );

    bfr new_Jinkela_buffer_5230 (
        .din(new_Jinkela_wire_7124),
        .dout(new_Jinkela_wire_7125)
    );

    bfr new_Jinkela_buffer_2922 (
        .din(new_Jinkela_wire_4247),
        .dout(new_Jinkela_wire_4248)
    );

    bfr new_Jinkela_buffer_2942 (
        .din(new_Jinkela_wire_4269),
        .dout(new_Jinkela_wire_4270)
    );

    bfr new_Jinkela_buffer_5231 (
        .din(new_Jinkela_wire_7125),
        .dout(new_Jinkela_wire_7126)
    );

    bfr new_Jinkela_buffer_2923 (
        .din(new_Jinkela_wire_4248),
        .dout(new_Jinkela_wire_4249)
    );

    bfr new_Jinkela_buffer_5277 (
        .din(_0689_),
        .dout(new_Jinkela_wire_7184)
    );

    spl2 new_Jinkela_splitter_736 (
        .a(_0111_),
        .b(new_Jinkela_wire_7189),
        .c(new_Jinkela_wire_7190)
    );

    bfr new_Jinkela_buffer_2959 (
        .din(new_Jinkela_wire_4286),
        .dout(new_Jinkela_wire_4287)
    );

    bfr new_Jinkela_buffer_5232 (
        .din(new_Jinkela_wire_7126),
        .dout(new_Jinkela_wire_7127)
    );

    bfr new_Jinkela_buffer_2924 (
        .din(new_Jinkela_wire_4249),
        .dout(new_Jinkela_wire_4250)
    );

    bfr new_Jinkela_buffer_5241 (
        .din(new_Jinkela_wire_7147),
        .dout(new_Jinkela_wire_7148)
    );

    bfr new_Jinkela_buffer_2943 (
        .din(new_Jinkela_wire_4270),
        .dout(new_Jinkela_wire_4271)
    );

    bfr new_Jinkela_buffer_5242 (
        .din(new_Jinkela_wire_7148),
        .dout(new_Jinkela_wire_7149)
    );

    bfr new_Jinkela_buffer_2925 (
        .din(new_Jinkela_wire_4250),
        .dout(new_Jinkela_wire_4251)
    );

    bfr new_Jinkela_buffer_5246 (
        .din(new_Jinkela_wire_7152),
        .dout(new_Jinkela_wire_7153)
    );

    spl2 new_Jinkela_splitter_506 (
        .a(_0885_),
        .b(new_Jinkela_wire_4336),
        .c(new_Jinkela_wire_4337)
    );

    bfr new_Jinkela_buffer_5243 (
        .din(new_Jinkela_wire_7149),
        .dout(new_Jinkela_wire_7150)
    );

    or_bb _2453_ (
        .a(new_Jinkela_wire_2531),
        .b(_0445_),
        .c(new_net_2439)
    );

    or_ii _2454_ (
        .a(new_Jinkela_wire_3617),
        .b(new_Jinkela_wire_3464),
        .c(_0449_)
    );

    and_bi _2455_ (
        .a(new_Jinkela_wire_5002),
        .b(new_Jinkela_wire_3435),
        .c(_0450_)
    );

    or_bb _2456_ (
        .a(_0450_),
        .b(new_Jinkela_wire_3496),
        .c(_0451_)
    );

    and_bi _2457_ (
        .a(_0449_),
        .b(new_Jinkela_wire_6184),
        .c(_0452_)
    );

    and_bi _2458_ (
        .a(new_Jinkela_wire_1271),
        .b(new_Jinkela_wire_6414),
        .c(_0453_)
    );

    and_bi _2459_ (
        .a(new_Jinkela_wire_253),
        .b(new_Jinkela_wire_2870),
        .c(_0454_)
    );

    or_bb _2460_ (
        .a(_0454_),
        .b(_0453_),
        .c(_0455_)
    );

    or_bb _2461_ (
        .a(new_Jinkela_wire_3135),
        .b(_0452_),
        .c(new_net_2401)
    );

    and_bi _2466_ (
        .a(new_Jinkela_wire_1223),
        .b(new_Jinkela_wire_2865),
        .c(_0460_)
    );

    and_bi _2467_ (
        .a(new_Jinkela_wire_190),
        .b(new_Jinkela_wire_6424),
        .c(_0461_)
    );

    or_bb _2468_ (
        .a(_0461_),
        .b(_0460_),
        .c(_0462_)
    );

    or_bb _2469_ (
        .a(new_Jinkela_wire_3570),
        .b(_0459_),
        .c(new_net_2355)
    );

    or_bb _2470_ (
        .a(new_Jinkela_wire_1615),
        .b(new_Jinkela_wire_3462),
        .c(_0463_)
    );

    and_bi _2471_ (
        .a(new_Jinkela_wire_5359),
        .b(new_Jinkela_wire_1480),
        .c(_0464_)
    );

    or_bb _2472_ (
        .a(_0464_),
        .b(new_Jinkela_wire_3522),
        .c(_0465_)
    );

    and_bi _2473_ (
        .a(new_Jinkela_wire_7199),
        .b(_0465_),
        .c(_0466_)
    );

    and_bi _2474_ (
        .a(new_Jinkela_wire_121),
        .b(new_Jinkela_wire_2868),
        .c(_0467_)
    );

    and_bi _2475_ (
        .a(new_Jinkela_wire_1388),
        .b(new_Jinkela_wire_6419),
        .c(_0468_)
    );

    or_bb _2476_ (
        .a(_0468_),
        .b(_0467_),
        .c(_0469_)
    );

    or_bb _2477_ (
        .a(new_Jinkela_wire_2153),
        .b(_0466_),
        .c(new_net_2457)
    );

    or_ii _2478_ (
        .a(new_Jinkela_wire_6908),
        .b(new_Jinkela_wire_1471),
        .c(_0470_)
    );

    and_bi _2479_ (
        .a(new_Jinkela_wire_6990),
        .b(new_Jinkela_wire_1473),
        .c(_0471_)
    );

    or_bb _2480_ (
        .a(_0471_),
        .b(new_Jinkela_wire_3516),
        .c(_0472_)
    );

    and_bi _2481_ (
        .a(new_Jinkela_wire_7015),
        .b(_0472_),
        .c(_0473_)
    );

    and_bi _2482_ (
        .a(new_Jinkela_wire_226),
        .b(new_Jinkela_wire_2864),
        .c(_0474_)
    );

    and_bi _2483_ (
        .a(new_Jinkela_wire_1242),
        .b(new_Jinkela_wire_6420),
        .c(_0475_)
    );

    or_bb _2484_ (
        .a(_0475_),
        .b(_0474_),
        .c(_0476_)
    );

    or_bb _2485_ (
        .a(new_Jinkela_wire_7500),
        .b(_0473_),
        .c(new_net_2483)
    );

    or_bi _2486_ (
        .a(new_Jinkela_wire_395),
        .b(new_Jinkela_wire_6791),
        .c(_0477_)
    );

    and_bb _2487_ (
        .a(new_Jinkela_wire_5774),
        .b(new_Jinkela_wire_392),
        .c(_0478_)
    );

    or_bb _2488_ (
        .a(_0478_),
        .b(new_Jinkela_wire_3984),
        .c(_0479_)
    );

    and_bi _2489_ (
        .a(_0477_),
        .b(_0479_),
        .c(_0480_)
    );

    and_bi _2490_ (
        .a(new_Jinkela_wire_1224),
        .b(new_Jinkela_wire_5811),
        .c(_0481_)
    );

    and_bi _2491_ (
        .a(new_Jinkela_wire_191),
        .b(new_Jinkela_wire_7879),
        .c(_0482_)
    );

    or_bb _2492_ (
        .a(_0482_),
        .b(_0481_),
        .c(_0483_)
    );

    or_bb _2493_ (
        .a(new_Jinkela_wire_6986),
        .b(_0480_),
        .c(new_net_2479)
    );

    or_bi _2494_ (
        .a(new_Jinkela_wire_394),
        .b(new_Jinkela_wire_5363),
        .c(_0484_)
    );

    and_bi _2495_ (
        .a(new_Jinkela_wire_391),
        .b(new_Jinkela_wire_1618),
        .c(_0485_)
    );

    or_bb _2496_ (
        .a(_0485_),
        .b(new_Jinkela_wire_3985),
        .c(_0486_)
    );

    and_bi _2497_ (
        .a(_0484_),
        .b(_0486_),
        .c(_0487_)
    );

    and_bi _1739_ (
        .a(new_Jinkela_wire_186),
        .b(new_Jinkela_wire_6693),
        .c(_1029_)
    );

    bfr new_Jinkela_buffer_2765 (
        .din(_0939_),
        .dout(new_Jinkela_wire_4074)
    );

    bfr new_Jinkela_buffer_3925 (
        .din(new_Jinkela_wire_5450),
        .dout(new_Jinkela_wire_5451)
    );

    bfr new_Jinkela_buffer_2673 (
        .din(new_Jinkela_wire_3944),
        .dout(new_Jinkela_wire_3945)
    );

    or_ii _1740_ (
        .a(new_Jinkela_wire_2262),
        .b(new_Jinkela_wire_1631),
        .c(_1030_)
    );

    bfr new_Jinkela_buffer_2640 (
        .din(new_Jinkela_wire_3909),
        .dout(new_Jinkela_wire_3910)
    );

    bfr new_Jinkela_buffer_3970 (
        .din(new_net_2469),
        .dout(new_Jinkela_wire_5496)
    );

    and_ii _1741_ (
        .a(new_Jinkela_wire_2261),
        .b(new_Jinkela_wire_1627),
        .c(_1031_)
    );

    bfr new_Jinkela_buffer_3926 (
        .din(new_Jinkela_wire_5451),
        .dout(new_Jinkela_wire_5452)
    );

    and_bi _1742_ (
        .a(_1030_),
        .b(_1031_),
        .c(_1032_)
    );

    bfr new_Jinkela_buffer_2641 (
        .din(new_Jinkela_wire_3910),
        .dout(new_Jinkela_wire_3911)
    );

    bfr new_Jinkela_buffer_3965 (
        .din(new_Jinkela_wire_5490),
        .dout(new_Jinkela_wire_5491)
    );

    or_bb _1743_ (
        .a(new_Jinkela_wire_2534),
        .b(new_Jinkela_wire_1091),
        .c(_1033_)
    );

    bfr new_Jinkela_buffer_2674 (
        .din(new_Jinkela_wire_3945),
        .dout(new_Jinkela_wire_3946)
    );

    bfr new_Jinkela_buffer_3927 (
        .din(new_Jinkela_wire_5452),
        .dout(new_Jinkela_wire_5453)
    );

    or_bb _1744_ (
        .a(new_Jinkela_wire_851),
        .b(new_Jinkela_wire_312),
        .c(_1034_)
    );

    bfr new_Jinkela_buffer_2642 (
        .din(new_Jinkela_wire_3911),
        .dout(new_Jinkela_wire_3912)
    );

    bfr new_Jinkela_buffer_3981 (
        .din(new_net_25),
        .dout(new_Jinkela_wire_5507)
    );

    bfr new_Jinkela_buffer_4020 (
        .din(_0118_),
        .dout(new_Jinkela_wire_5550)
    );

    and_bi _1745_ (
        .a(new_Jinkela_wire_855),
        .b(new_Jinkela_wire_210),
        .c(_1035_)
    );

    spl4L new_Jinkela_splitter_491 (
        .a(new_Jinkela_wire_4024),
        .d(new_Jinkela_wire_4025),
        .e(new_Jinkela_wire_4026),
        .b(new_Jinkela_wire_4027),
        .c(new_Jinkela_wire_4028)
    );

    bfr new_Jinkela_buffer_3928 (
        .din(new_Jinkela_wire_5453),
        .dout(new_Jinkela_wire_5454)
    );

    bfr new_Jinkela_buffer_2699 (
        .din(new_Jinkela_wire_3988),
        .dout(new_Jinkela_wire_3989)
    );

    and_bi _1746_ (
        .a(_1034_),
        .b(_1035_),
        .c(_1036_)
    );

    bfr new_Jinkela_buffer_2643 (
        .din(new_Jinkela_wire_3912),
        .dout(new_Jinkela_wire_3913)
    );

    bfr new_Jinkela_buffer_3966 (
        .din(new_Jinkela_wire_5491),
        .dout(new_Jinkela_wire_5492)
    );

    or_bb _1747_ (
        .a(_1036_),
        .b(new_Jinkela_wire_3771),
        .c(_1037_)
    );

    bfr new_Jinkela_buffer_3929 (
        .din(new_Jinkela_wire_5454),
        .dout(new_Jinkela_wire_5455)
    );

    or_ii _1748_ (
        .a(new_Jinkela_wire_1582),
        .b(new_Jinkela_wire_850),
        .c(_1038_)
    );

    bfr new_Jinkela_buffer_2644 (
        .din(new_Jinkela_wire_3913),
        .dout(new_Jinkela_wire_3914)
    );

    bfr new_Jinkela_buffer_3971 (
        .din(new_Jinkela_wire_5496),
        .dout(new_Jinkela_wire_5497)
    );

    and_bi _1749_ (
        .a(new_Jinkela_wire_1279),
        .b(new_Jinkela_wire_852),
        .c(_1039_)
    );

    bfr new_Jinkela_buffer_2675 (
        .din(new_Jinkela_wire_3946),
        .dout(new_Jinkela_wire_3947)
    );

    bfr new_Jinkela_buffer_3930 (
        .din(new_Jinkela_wire_5455),
        .dout(new_Jinkela_wire_5456)
    );

    bfr new_Jinkela_buffer_2700 (
        .din(new_Jinkela_wire_3989),
        .dout(new_Jinkela_wire_3990)
    );

    and_bi _1750_ (
        .a(_1038_),
        .b(_1039_),
        .c(_1040_)
    );

    bfr new_Jinkela_buffer_2645 (
        .din(new_Jinkela_wire_3914),
        .dout(new_Jinkela_wire_3915)
    );

    bfr new_Jinkela_buffer_3967 (
        .din(new_Jinkela_wire_5492),
        .dout(new_Jinkela_wire_5493)
    );

    and_bi _1751_ (
        .a(new_Jinkela_wire_3773),
        .b(_1040_),
        .c(_1041_)
    );

    bfr new_Jinkela_buffer_3931 (
        .din(new_Jinkela_wire_5456),
        .dout(new_Jinkela_wire_5457)
    );

    bfr new_Jinkela_buffer_2676 (
        .din(new_Jinkela_wire_3947),
        .dout(new_Jinkela_wire_3948)
    );

    and_bi _1752_ (
        .a(_1037_),
        .b(_1041_),
        .c(_1042_)
    );

    bfr new_Jinkela_buffer_2646 (
        .din(new_Jinkela_wire_3915),
        .dout(new_Jinkela_wire_3916)
    );

    bfr new_Jinkela_buffer_3982 (
        .din(new_Jinkela_wire_5507),
        .dout(new_Jinkela_wire_5508)
    );

    and_bi _1753_ (
        .a(new_Jinkela_wire_1042),
        .b(new_Jinkela_wire_2413),
        .c(_1043_)
    );

    bfr new_Jinkela_buffer_3932 (
        .din(new_Jinkela_wire_5457),
        .dout(new_Jinkela_wire_5458)
    );

    or_bb _1754_ (
        .a(_1043_),
        .b(new_Jinkela_wire_4827),
        .c(_1044_)
    );

    bfr new_Jinkela_buffer_2647 (
        .din(new_Jinkela_wire_3916),
        .dout(new_Jinkela_wire_3917)
    );

    bfr new_Jinkela_buffer_3968 (
        .din(new_Jinkela_wire_5493),
        .dout(new_Jinkela_wire_5494)
    );

    and_bi _1755_ (
        .a(_1033_),
        .b(new_Jinkela_wire_3410),
        .c(_1045_)
    );

    bfr new_Jinkela_buffer_3933 (
        .din(new_Jinkela_wire_5458),
        .dout(new_Jinkela_wire_5459)
    );

    bfr new_Jinkela_buffer_2677 (
        .din(new_Jinkela_wire_3948),
        .dout(new_Jinkela_wire_3949)
    );

    and_ii _1756_ (
        .a(_1045_),
        .b(new_Jinkela_wire_2355),
        .c(new_net_23)
    );

    bfr new_Jinkela_buffer_2648 (
        .din(new_Jinkela_wire_3917),
        .dout(new_Jinkela_wire_3918)
    );

    bfr new_Jinkela_buffer_3972 (
        .din(new_Jinkela_wire_5497),
        .dout(new_Jinkela_wire_5498)
    );

    inv _1757_ (
        .din(new_Jinkela_wire_641),
        .dout(_1046_)
    );

    bfr new_Jinkela_buffer_3934 (
        .din(new_Jinkela_wire_5459),
        .dout(new_Jinkela_wire_5460)
    );

    inv _1758_ (
        .din(new_Jinkela_wire_452),
        .dout(_1047_)
    );

    bfr new_Jinkela_buffer_2649 (
        .din(new_Jinkela_wire_3918),
        .dout(new_Jinkela_wire_3919)
    );

    bfr new_Jinkela_buffer_3969 (
        .din(new_Jinkela_wire_5494),
        .dout(new_Jinkela_wire_5495)
    );

    and_bi _1759_ (
        .a(new_Jinkela_wire_4991),
        .b(new_Jinkela_wire_7209),
        .c(_1048_)
    );

    bfr new_Jinkela_buffer_2678 (
        .din(new_Jinkela_wire_3949),
        .dout(new_Jinkela_wire_3950)
    );

    bfr new_Jinkela_buffer_3935 (
        .din(new_Jinkela_wire_5460),
        .dout(new_Jinkela_wire_5461)
    );

    bfr new_Jinkela_buffer_2701 (
        .din(new_Jinkela_wire_3990),
        .dout(new_Jinkela_wire_3991)
    );

    and_bi _1760_ (
        .a(new_Jinkela_wire_7212),
        .b(new_Jinkela_wire_6559),
        .c(_1049_)
    );

    bfr new_Jinkela_buffer_2650 (
        .din(new_Jinkela_wire_3919),
        .dout(new_Jinkela_wire_3920)
    );

    bfr new_Jinkela_buffer_4047 (
        .din(_0291_),
        .dout(new_Jinkela_wire_5599)
    );

    and_bi _1761_ (
        .a(new_Jinkela_wire_4614),
        .b(new_Jinkela_wire_2861),
        .c(_1050_)
    );

    bfr new_Jinkela_buffer_2679 (
        .din(new_Jinkela_wire_3950),
        .dout(new_Jinkela_wire_3951)
    );

    bfr new_Jinkela_buffer_3936 (
        .din(new_Jinkela_wire_5461),
        .dout(new_Jinkela_wire_5462)
    );

    or_bb _1762_ (
        .a(new_Jinkela_wire_4988),
        .b(new_Jinkela_wire_7040),
        .c(_1051_)
    );

    bfr new_Jinkela_buffer_2651 (
        .din(new_Jinkela_wire_3920),
        .dout(new_Jinkela_wire_3921)
    );

    bfr new_Jinkela_buffer_3973 (
        .din(new_Jinkela_wire_5498),
        .dout(new_Jinkela_wire_5499)
    );

    or_bi _1763_ (
        .a(new_Jinkela_wire_3216),
        .b(_1051_),
        .c(_1052_)
    );

    bfr new_Jinkela_buffer_3937 (
        .din(new_Jinkela_wire_5462),
        .dout(new_Jinkela_wire_5463)
    );

    spl2 new_Jinkela_splitter_490 (
        .a(new_Jinkela_wire_4021),
        .b(new_Jinkela_wire_4022),
        .c(new_Jinkela_wire_4023)
    );

    and_bi _1764_ (
        .a(new_Jinkela_wire_7999),
        .b(new_Jinkela_wire_2310),
        .c(_1053_)
    );

    bfr new_Jinkela_buffer_2652 (
        .din(new_Jinkela_wire_3921),
        .dout(new_Jinkela_wire_3922)
    );

    spl2 new_Jinkela_splitter_594 (
        .a(_1218_),
        .b(new_Jinkela_wire_5597),
        .c(new_Jinkela_wire_5598)
    );

    bfr new_Jinkela_buffer_3983 (
        .din(new_Jinkela_wire_5508),
        .dout(new_Jinkela_wire_5509)
    );

    or_bb _1765_ (
        .a(_1053_),
        .b(new_Jinkela_wire_6121),
        .c(_1054_)
    );

    bfr new_Jinkela_buffer_3938 (
        .din(new_Jinkela_wire_5463),
        .dout(new_Jinkela_wire_5464)
    );

    and_bi _1766_ (
        .a(new_Jinkela_wire_4194),
        .b(new_Jinkela_wire_3532),
        .c(_1055_)
    );

    bfr new_Jinkela_buffer_2653 (
        .din(new_Jinkela_wire_3922),
        .dout(new_Jinkela_wire_3923)
    );

    bfr new_Jinkela_buffer_3974 (
        .din(new_Jinkela_wire_5499),
        .dout(new_Jinkela_wire_5500)
    );

    and_bi _1767_ (
        .a(new_Jinkela_wire_3533),
        .b(new_Jinkela_wire_4195),
        .c(_1056_)
    );

    bfr new_Jinkela_buffer_3939 (
        .din(new_Jinkela_wire_5464),
        .dout(new_Jinkela_wire_5465)
    );

    or_bb _1768_ (
        .a(_1056_),
        .b(_1055_),
        .c(_1057_)
    );

    bfr new_Jinkela_buffer_2654 (
        .din(new_Jinkela_wire_3923),
        .dout(new_Jinkela_wire_3924)
    );

    or_bb _1769_ (
        .a(new_Jinkela_wire_3714),
        .b(new_Jinkela_wire_3376),
        .c(_1058_)
    );

    spl4L new_Jinkela_splitter_492 (
        .a(new_Jinkela_wire_4029),
        .d(new_Jinkela_wire_4030),
        .e(new_Jinkela_wire_4031),
        .b(new_Jinkela_wire_4032),
        .c(new_Jinkela_wire_4033)
    );

    bfr new_Jinkela_buffer_3940 (
        .din(new_Jinkela_wire_5465),
        .dout(new_Jinkela_wire_5466)
    );

    bfr new_Jinkela_buffer_2681 (
        .din(new_Jinkela_wire_3952),
        .dout(new_Jinkela_wire_3953)
    );

    and_bb _1770_ (
        .a(new_Jinkela_wire_3715),
        .b(new_Jinkela_wire_3375),
        .c(_1059_)
    );

    bfr new_Jinkela_buffer_2655 (
        .din(new_Jinkela_wire_3924),
        .dout(new_Jinkela_wire_3925)
    );

    bfr new_Jinkela_buffer_3975 (
        .din(new_Jinkela_wire_5500),
        .dout(new_Jinkela_wire_5501)
    );

    or_bb _1771_ (
        .a(_1059_),
        .b(new_Jinkela_wire_146),
        .c(_1060_)
    );

    bfr new_Jinkela_buffer_3941 (
        .din(new_Jinkela_wire_5466),
        .dout(new_Jinkela_wire_5467)
    );

    bfr new_Jinkela_buffer_2680 (
        .din(new_Jinkela_wire_3951),
        .dout(new_Jinkela_wire_3952)
    );

    and_bi _1772_ (
        .a(new_Jinkela_wire_4345),
        .b(_1060_),
        .c(_1061_)
    );

    bfr new_Jinkela_buffer_2656 (
        .din(new_Jinkela_wire_3925),
        .dout(new_Jinkela_wire_3926)
    );

    bfr new_Jinkela_buffer_3984 (
        .din(new_Jinkela_wire_5509),
        .dout(new_Jinkela_wire_5510)
    );

    and_ii _1773_ (
        .a(new_Jinkela_wire_2199),
        .b(new_Jinkela_wire_2205),
        .c(_1062_)
    );

    bfr new_Jinkela_buffer_2703 (
        .din(new_Jinkela_wire_3992),
        .dout(new_Jinkela_wire_3993)
    );

    bfr new_Jinkela_buffer_3942 (
        .din(new_Jinkela_wire_5467),
        .dout(new_Jinkela_wire_5468)
    );

    and_bi _1774_ (
        .a(new_Jinkela_wire_2208),
        .b(new_Jinkela_wire_4987),
        .c(_1063_)
    );

    bfr new_Jinkela_buffer_2657 (
        .din(new_Jinkela_wire_3926),
        .dout(new_Jinkela_wire_3927)
    );

    bfr new_Jinkela_buffer_3976 (
        .din(new_Jinkela_wire_5501),
        .dout(new_Jinkela_wire_5502)
    );

    and_ii _1775_ (
        .a(_1063_),
        .b(new_Jinkela_wire_2094),
        .c(_1064_)
    );

    bfr new_Jinkela_buffer_2702 (
        .din(new_Jinkela_wire_3991),
        .dout(new_Jinkela_wire_3992)
    );

    bfr new_Jinkela_buffer_3943 (
        .din(new_Jinkela_wire_5468),
        .dout(new_Jinkela_wire_5469)
    );

    bfr new_Jinkela_buffer_2682 (
        .din(new_Jinkela_wire_3953),
        .dout(new_Jinkela_wire_3954)
    );

    or_bb _1776_ (
        .a(new_Jinkela_wire_5402),
        .b(new_Jinkela_wire_6246),
        .c(_1065_)
    );

    bfr new_Jinkela_buffer_2658 (
        .din(new_Jinkela_wire_3927),
        .dout(new_Jinkela_wire_3928)
    );

    bfr new_Jinkela_buffer_4021 (
        .din(new_Jinkela_wire_5550),
        .dout(new_Jinkela_wire_5551)
    );

    bfr new_Jinkela_buffer_4022 (
        .din(_0099_),
        .dout(new_Jinkela_wire_5554)
    );

    and_bb _1777_ (
        .a(new_Jinkela_wire_5403),
        .b(new_Jinkela_wire_6244),
        .c(_1066_)
    );

    bfr new_Jinkela_buffer_3944 (
        .din(new_Jinkela_wire_5469),
        .dout(new_Jinkela_wire_5470)
    );

    bfr new_Jinkela_buffer_2732 (
        .din(new_Jinkela_wire_4034),
        .dout(new_Jinkela_wire_4035)
    );

    and_bi _1778_ (
        .a(_1065_),
        .b(_1066_),
        .c(_1067_)
    );

    bfr new_Jinkela_buffer_2659 (
        .din(new_Jinkela_wire_3928),
        .dout(new_Jinkela_wire_3929)
    );

    bfr new_Jinkela_buffer_3977 (
        .din(new_Jinkela_wire_5502),
        .dout(new_Jinkela_wire_5503)
    );

    or_bb _1779_ (
        .a(new_Jinkela_wire_2309),
        .b(new_Jinkela_wire_1960),
        .c(_1068_)
    );

    bfr new_Jinkela_buffer_3945 (
        .din(new_Jinkela_wire_5470),
        .dout(new_Jinkela_wire_5471)
    );

    bfr new_Jinkela_buffer_2683 (
        .din(new_Jinkela_wire_3954),
        .dout(new_Jinkela_wire_3955)
    );

    and_bi _1780_ (
        .a(new_Jinkela_wire_2311),
        .b(new_Jinkela_wire_2853),
        .c(_1069_)
    );

    bfr new_Jinkela_buffer_2660 (
        .din(new_Jinkela_wire_3929),
        .dout(new_Jinkela_wire_3930)
    );

    spl3L new_Jinkela_splitter_350 (
        .a(_0744_),
        .d(new_Jinkela_wire_2199),
        .b(new_Jinkela_wire_2200),
        .c(new_Jinkela_wire_2201)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(new_Jinkela_wire_2107),
        .dout(new_Jinkela_wire_2108)
    );

    bfr new_Jinkela_buffer_2867 (
        .din(new_Jinkela_wire_4188),
        .dout(new_Jinkela_wire_4189)
    );

    bfr new_Jinkela_buffer_5160 (
        .din(new_Jinkela_wire_7033),
        .dout(new_Jinkela_wire_7034)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_2126),
        .dout(new_Jinkela_wire_2127)
    );

    spl2 new_Jinkela_splitter_503 (
        .a(_0150_),
        .b(new_Jinkela_wire_4254),
        .c(new_Jinkela_wire_4255)
    );

    bfr new_Jinkela_buffer_5171 (
        .din(new_Jinkela_wire_7049),
        .dout(new_Jinkela_wire_7050)
    );

    spl2 new_Jinkela_splitter_502 (
        .a(new_Jinkela_wire_4201),
        .b(new_Jinkela_wire_4202),
        .c(new_Jinkela_wire_4203)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_2108),
        .dout(new_Jinkela_wire_2109)
    );

    bfr new_Jinkela_buffer_2868 (
        .din(new_Jinkela_wire_4189),
        .dout(new_Jinkela_wire_4190)
    );

    bfr new_Jinkela_buffer_5161 (
        .din(new_Jinkela_wire_7034),
        .dout(new_Jinkela_wire_7035)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(new_Jinkela_wire_2157),
        .dout(new_Jinkela_wire_2158)
    );

    bfr new_Jinkela_buffer_5198 (
        .din(new_Jinkela_wire_7076),
        .dout(new_Jinkela_wire_7077)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(new_Jinkela_wire_2109),
        .dout(new_Jinkela_wire_2110)
    );

    bfr new_Jinkela_buffer_2869 (
        .din(new_Jinkela_wire_4190),
        .dout(new_Jinkela_wire_4191)
    );

    bfr new_Jinkela_buffer_5172 (
        .din(new_Jinkela_wire_7050),
        .dout(new_Jinkela_wire_7051)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_2127),
        .dout(new_Jinkela_wire_2128)
    );

    bfr new_Jinkela_buffer_2894 (
        .din(new_Jinkela_wire_4219),
        .dout(new_Jinkela_wire_4220)
    );

    spl2 new_Jinkela_splitter_724 (
        .a(new_Jinkela_wire_7080),
        .b(new_Jinkela_wire_7081),
        .c(new_Jinkela_wire_7082)
    );

    bfr new_Jinkela_buffer_2928 (
        .din(new_net_2433),
        .dout(new_Jinkela_wire_4256)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_2110),
        .dout(new_Jinkela_wire_2111)
    );

    bfr new_Jinkela_buffer_2870 (
        .din(new_Jinkela_wire_4191),
        .dout(new_Jinkela_wire_4192)
    );

    bfr new_Jinkela_buffer_5173 (
        .din(new_Jinkela_wire_7051),
        .dout(new_Jinkela_wire_7052)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_2160),
        .dout(new_Jinkela_wire_2161)
    );

    bfr new_Jinkela_buffer_2880 (
        .din(new_Jinkela_wire_4205),
        .dout(new_Jinkela_wire_4206)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_Jinkela_wire_2111),
        .dout(new_Jinkela_wire_2112)
    );

    bfr new_Jinkela_buffer_2871 (
        .din(new_Jinkela_wire_4192),
        .dout(new_Jinkela_wire_4193)
    );

    bfr new_Jinkela_buffer_5174 (
        .din(new_Jinkela_wire_7052),
        .dout(new_Jinkela_wire_7053)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(new_Jinkela_wire_2128),
        .dout(new_Jinkela_wire_2129)
    );

    bfr new_Jinkela_buffer_2881 (
        .din(new_Jinkela_wire_4206),
        .dout(new_Jinkela_wire_4207)
    );

    spl2 new_Jinkela_splitter_727 (
        .a(_0872_),
        .b(new_Jinkela_wire_7107),
        .c(new_Jinkela_wire_7109)
    );

    bfr new_Jinkela_buffer_5200 (
        .din(new_Jinkela_wire_7086),
        .dout(new_Jinkela_wire_7087)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_2112),
        .dout(new_Jinkela_wire_2113)
    );

    bfr new_Jinkela_buffer_5175 (
        .din(new_Jinkela_wire_7053),
        .dout(new_Jinkela_wire_7054)
    );

    bfr new_Jinkela_buffer_2929 (
        .din(new_Jinkela_wire_4256),
        .dout(new_Jinkela_wire_4257)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(new_Jinkela_wire_2158),
        .dout(new_Jinkela_wire_2159)
    );

    bfr new_Jinkela_buffer_2882 (
        .din(new_Jinkela_wire_4207),
        .dout(new_Jinkela_wire_4208)
    );

    bfr new_Jinkela_buffer_5219 (
        .din(new_Jinkela_wire_7113),
        .dout(new_Jinkela_wire_7114)
    );

    spl2 new_Jinkela_splitter_726 (
        .a(_0975_),
        .b(new_Jinkela_wire_7105),
        .c(new_Jinkela_wire_7106)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_2113),
        .dout(new_Jinkela_wire_2114)
    );

    bfr new_Jinkela_buffer_2895 (
        .din(new_Jinkela_wire_4220),
        .dout(new_Jinkela_wire_4221)
    );

    bfr new_Jinkela_buffer_5176 (
        .din(new_Jinkela_wire_7054),
        .dout(new_Jinkela_wire_7055)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(new_Jinkela_wire_2129),
        .dout(new_Jinkela_wire_2130)
    );

    bfr new_Jinkela_buffer_2883 (
        .din(new_Jinkela_wire_4208),
        .dout(new_Jinkela_wire_4209)
    );

    bfr new_Jinkela_buffer_5201 (
        .din(new_Jinkela_wire_7087),
        .dout(new_Jinkela_wire_7088)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_2114),
        .dout(new_Jinkela_wire_2115)
    );

    bfr new_Jinkela_buffer_5177 (
        .din(new_Jinkela_wire_7055),
        .dout(new_Jinkela_wire_7056)
    );

    bfr new_Jinkela_buffer_2884 (
        .din(new_Jinkela_wire_4209),
        .dout(new_Jinkela_wire_4210)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_2201),
        .dout(new_Jinkela_wire_2202)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(new_Jinkela_wire_2115),
        .dout(new_Jinkela_wire_2116)
    );

    bfr new_Jinkela_buffer_2896 (
        .din(new_Jinkela_wire_4221),
        .dout(new_Jinkela_wire_4222)
    );

    bfr new_Jinkela_buffer_5178 (
        .din(new_Jinkela_wire_7056),
        .dout(new_Jinkela_wire_7057)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(new_Jinkela_wire_2130),
        .dout(new_Jinkela_wire_2131)
    );

    bfr new_Jinkela_buffer_2885 (
        .din(new_Jinkela_wire_4210),
        .dout(new_Jinkela_wire_4211)
    );

    bfr new_Jinkela_buffer_5202 (
        .din(new_Jinkela_wire_7088),
        .dout(new_Jinkela_wire_7089)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_2116),
        .dout(new_Jinkela_wire_2117)
    );

    bfr new_Jinkela_buffer_2952 (
        .din(new_net_2377),
        .dout(new_Jinkela_wire_4280)
    );

    bfr new_Jinkela_buffer_5179 (
        .din(new_Jinkela_wire_7057),
        .dout(new_Jinkela_wire_7058)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_2161),
        .dout(new_Jinkela_wire_2162)
    );

    bfr new_Jinkela_buffer_2886 (
        .din(new_Jinkela_wire_4211),
        .dout(new_Jinkela_wire_4212)
    );

    spl2 new_Jinkela_splitter_729 (
        .a(_0249_),
        .b(new_Jinkela_wire_7128),
        .c(new_Jinkela_wire_7129)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_2131),
        .dout(new_Jinkela_wire_2132)
    );

    bfr new_Jinkela_buffer_2897 (
        .din(new_Jinkela_wire_4222),
        .dout(new_Jinkela_wire_4223)
    );

    bfr new_Jinkela_buffer_5180 (
        .din(new_Jinkela_wire_7058),
        .dout(new_Jinkela_wire_7059)
    );

    bfr new_Jinkela_buffer_2887 (
        .din(new_Jinkela_wire_4212),
        .dout(new_Jinkela_wire_4213)
    );

    bfr new_Jinkela_buffer_5203 (
        .din(new_Jinkela_wire_7089),
        .dout(new_Jinkela_wire_7090)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_2132),
        .dout(new_Jinkela_wire_2133)
    );

    spl2 new_Jinkela_splitter_504 (
        .a(_0737_),
        .b(new_Jinkela_wire_4308),
        .c(new_Jinkela_wire_4309)
    );

    bfr new_Jinkela_buffer_5181 (
        .din(new_Jinkela_wire_7059),
        .dout(new_Jinkela_wire_7060)
    );

    bfr new_Jinkela_buffer_2980 (
        .din(_0195_),
        .dout(new_Jinkela_wire_4310)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_Jinkela_wire_2162),
        .dout(new_Jinkela_wire_2163)
    );

    bfr new_Jinkela_buffer_2888 (
        .din(new_Jinkela_wire_4213),
        .dout(new_Jinkela_wire_4214)
    );

    spl2 new_Jinkela_splitter_730 (
        .a(_0424_),
        .b(new_Jinkela_wire_7130),
        .c(new_Jinkela_wire_7131)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(new_Jinkela_wire_2133),
        .dout(new_Jinkela_wire_2134)
    );

    bfr new_Jinkela_buffer_2898 (
        .din(new_Jinkela_wire_4223),
        .dout(new_Jinkela_wire_4224)
    );

    bfr new_Jinkela_buffer_5182 (
        .din(new_Jinkela_wire_7060),
        .dout(new_Jinkela_wire_7061)
    );

    spl3L new_Jinkela_splitter_351 (
        .a(_0639_),
        .d(new_Jinkela_wire_2204),
        .b(new_Jinkela_wire_2205),
        .c(new_Jinkela_wire_2206)
    );

    bfr new_Jinkela_buffer_2889 (
        .din(new_Jinkela_wire_4214),
        .dout(new_Jinkela_wire_4215)
    );

    bfr new_Jinkela_buffer_5204 (
        .din(new_Jinkela_wire_7090),
        .dout(new_Jinkela_wire_7091)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_2134),
        .dout(new_Jinkela_wire_2135)
    );

    bfr new_Jinkela_buffer_2930 (
        .din(new_Jinkela_wire_4257),
        .dout(new_Jinkela_wire_4258)
    );

    bfr new_Jinkela_buffer_5183 (
        .din(new_Jinkela_wire_7061),
        .dout(new_Jinkela_wire_7062)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_2163),
        .dout(new_Jinkela_wire_2164)
    );

    bfr new_Jinkela_buffer_2890 (
        .din(new_Jinkela_wire_4215),
        .dout(new_Jinkela_wire_4216)
    );

    spl4L new_Jinkela_splitter_728 (
        .a(new_Jinkela_wire_7109),
        .d(new_Jinkela_wire_7110),
        .e(new_Jinkela_wire_7111),
        .b(new_Jinkela_wire_7112),
        .c(new_Jinkela_wire_7113)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_2135),
        .dout(new_Jinkela_wire_2136)
    );

    bfr new_Jinkela_buffer_2899 (
        .din(new_Jinkela_wire_4224),
        .dout(new_Jinkela_wire_4225)
    );

    bfr new_Jinkela_buffer_5184 (
        .din(new_Jinkela_wire_7062),
        .dout(new_Jinkela_wire_7063)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_2206),
        .dout(new_Jinkela_wire_2207)
    );

    bfr new_Jinkela_buffer_2891 (
        .din(new_Jinkela_wire_4216),
        .dout(new_Jinkela_wire_4217)
    );

    bfr new_Jinkela_buffer_5205 (
        .din(new_Jinkela_wire_7091),
        .dout(new_Jinkela_wire_7092)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_2136),
        .dout(new_Jinkela_wire_2137)
    );

    bfr new_Jinkela_buffer_2953 (
        .din(new_Jinkela_wire_4280),
        .dout(new_Jinkela_wire_4281)
    );

    bfr new_Jinkela_buffer_5185 (
        .din(new_Jinkela_wire_7063),
        .dout(new_Jinkela_wire_7064)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_2164),
        .dout(new_Jinkela_wire_2165)
    );

    bfr new_Jinkela_buffer_2892 (
        .din(new_Jinkela_wire_4217),
        .dout(new_Jinkela_wire_4218)
    );

    bfr new_Jinkela_buffer_5237 (
        .din(new_net_2355),
        .dout(new_Jinkela_wire_7140)
    );

    bfr new_Jinkela_buffer_5218 (
        .din(new_Jinkela_wire_7107),
        .dout(new_Jinkela_wire_7108)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_2137),
        .dout(new_Jinkela_wire_2138)
    );

    bfr new_Jinkela_buffer_2900 (
        .din(new_Jinkela_wire_4225),
        .dout(new_Jinkela_wire_4226)
    );

    bfr new_Jinkela_buffer_5186 (
        .din(new_Jinkela_wire_7064),
        .dout(new_Jinkela_wire_7065)
    );

    spl2 new_Jinkela_splitter_352 (
        .a(_0018_),
        .b(new_Jinkela_wire_2209),
        .c(new_Jinkela_wire_2210)
    );

    bfr new_Jinkela_buffer_2931 (
        .din(new_Jinkela_wire_4258),
        .dout(new_Jinkela_wire_4259)
    );

    bfr new_Jinkela_buffer_5206 (
        .din(new_Jinkela_wire_7092),
        .dout(new_Jinkela_wire_7093)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(new_Jinkela_wire_2202),
        .dout(new_Jinkela_wire_2203)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(new_Jinkela_wire_2138),
        .dout(new_Jinkela_wire_2139)
    );

    bfr new_Jinkela_buffer_2901 (
        .din(new_Jinkela_wire_4226),
        .dout(new_Jinkela_wire_4227)
    );

    bfr new_Jinkela_buffer_5187 (
        .din(new_Jinkela_wire_7065),
        .dout(new_Jinkela_wire_7066)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_2165),
        .dout(new_Jinkela_wire_2166)
    );

    bfr new_Jinkela_buffer_2983 (
        .din(new_net_2417),
        .dout(new_Jinkela_wire_4315)
    );

    bfr new_Jinkela_buffer_5235 (
        .din(_1067_),
        .dout(new_Jinkela_wire_7136)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(new_Jinkela_wire_2139),
        .dout(new_Jinkela_wire_2140)
    );

    bfr new_Jinkela_buffer_2902 (
        .din(new_Jinkela_wire_4227),
        .dout(new_Jinkela_wire_4228)
    );

    bfr new_Jinkela_buffer_5188 (
        .din(new_Jinkela_wire_7066),
        .dout(new_Jinkela_wire_7067)
    );

    bfr new_Jinkela_buffer_2932 (
        .din(new_Jinkela_wire_4259),
        .dout(new_Jinkela_wire_4260)
    );

    bfr new_Jinkela_buffer_5207 (
        .din(new_Jinkela_wire_7093),
        .dout(new_Jinkela_wire_7094)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(_1225_),
        .dout(new_Jinkela_wire_2211)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_2140),
        .dout(new_Jinkela_wire_2141)
    );

    bfr new_Jinkela_buffer_2903 (
        .din(new_Jinkela_wire_4228),
        .dout(new_Jinkela_wire_4229)
    );

    bfr new_Jinkela_buffer_5189 (
        .din(new_Jinkela_wire_7067),
        .dout(new_Jinkela_wire_7068)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_2166),
        .dout(new_Jinkela_wire_2167)
    );

    bfr new_Jinkela_buffer_2954 (
        .din(new_Jinkela_wire_4281),
        .dout(new_Jinkela_wire_4282)
    );

    bfr new_Jinkela_buffer_5233 (
        .din(new_Jinkela_wire_7131),
        .dout(new_Jinkela_wire_7132)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_2141),
        .dout(new_Jinkela_wire_2142)
    );

    bfr new_Jinkela_buffer_2904 (
        .din(new_Jinkela_wire_4229),
        .dout(new_Jinkela_wire_4230)
    );

    bfr new_Jinkela_buffer_5190 (
        .din(new_Jinkela_wire_7068),
        .dout(new_Jinkela_wire_7069)
    );

    bfr new_Jinkela_buffer_2933 (
        .din(new_Jinkela_wire_4260),
        .dout(new_Jinkela_wire_4261)
    );

    bfr new_Jinkela_buffer_5208 (
        .din(new_Jinkela_wire_7094),
        .dout(new_Jinkela_wire_7095)
    );

    bfr new_Jinkela_buffer_4075 (
        .din(new_net_2401),
        .dout(new_Jinkela_wire_5627)
    );

    bfr new_Jinkela_buffer_3946 (
        .din(new_Jinkela_wire_5471),
        .dout(new_Jinkela_wire_5472)
    );

    bfr new_Jinkela_buffer_3978 (
        .din(new_Jinkela_wire_5503),
        .dout(new_Jinkela_wire_5504)
    );

    bfr new_Jinkela_buffer_3947 (
        .din(new_Jinkela_wire_5472),
        .dout(new_Jinkela_wire_5473)
    );

    bfr new_Jinkela_buffer_3985 (
        .din(new_Jinkela_wire_5510),
        .dout(new_Jinkela_wire_5511)
    );

    bfr new_Jinkela_buffer_3948 (
        .din(new_Jinkela_wire_5473),
        .dout(new_Jinkela_wire_5474)
    );

    bfr new_Jinkela_buffer_3979 (
        .din(new_Jinkela_wire_5504),
        .dout(new_Jinkela_wire_5505)
    );

    bfr new_Jinkela_buffer_3949 (
        .din(new_Jinkela_wire_5474),
        .dout(new_Jinkela_wire_5475)
    );

    spl2 new_Jinkela_splitter_584 (
        .a(new_Jinkela_wire_5551),
        .b(new_Jinkela_wire_5552),
        .c(new_Jinkela_wire_5553)
    );

    bfr new_Jinkela_buffer_3950 (
        .din(new_Jinkela_wire_5475),
        .dout(new_Jinkela_wire_5476)
    );

    bfr new_Jinkela_buffer_3980 (
        .din(new_Jinkela_wire_5505),
        .dout(new_Jinkela_wire_5506)
    );

    bfr new_Jinkela_buffer_3951 (
        .din(new_Jinkela_wire_5476),
        .dout(new_Jinkela_wire_5477)
    );

    bfr new_Jinkela_buffer_3986 (
        .din(new_Jinkela_wire_5511),
        .dout(new_Jinkela_wire_5512)
    );

    bfr new_Jinkela_buffer_3952 (
        .din(new_Jinkela_wire_5477),
        .dout(new_Jinkela_wire_5478)
    );

    bfr new_Jinkela_buffer_4048 (
        .din(new_Jinkela_wire_5599),
        .dout(new_Jinkela_wire_5600)
    );

    bfr new_Jinkela_buffer_3953 (
        .din(new_Jinkela_wire_5478),
        .dout(new_Jinkela_wire_5479)
    );

    bfr new_Jinkela_buffer_3987 (
        .din(new_Jinkela_wire_5512),
        .dout(new_Jinkela_wire_5513)
    );

    bfr new_Jinkela_buffer_3954 (
        .din(new_Jinkela_wire_5479),
        .dout(new_Jinkela_wire_5480)
    );

    bfr new_Jinkela_buffer_4062 (
        .din(_0811_),
        .dout(new_Jinkela_wire_5614)
    );

    bfr new_Jinkela_buffer_3955 (
        .din(new_Jinkela_wire_5480),
        .dout(new_Jinkela_wire_5481)
    );

    bfr new_Jinkela_buffer_3988 (
        .din(new_Jinkela_wire_5513),
        .dout(new_Jinkela_wire_5514)
    );

    bfr new_Jinkela_buffer_3956 (
        .din(new_Jinkela_wire_5481),
        .dout(new_Jinkela_wire_5482)
    );

    bfr new_Jinkela_buffer_3957 (
        .din(new_Jinkela_wire_5482),
        .dout(new_Jinkela_wire_5483)
    );

    bfr new_Jinkela_buffer_3989 (
        .din(new_Jinkela_wire_5514),
        .dout(new_Jinkela_wire_5515)
    );

    bfr new_Jinkela_buffer_3958 (
        .din(new_Jinkela_wire_5483),
        .dout(new_Jinkela_wire_5484)
    );

    bfr new_Jinkela_buffer_3959 (
        .din(new_Jinkela_wire_5484),
        .dout(new_Jinkela_wire_5485)
    );

    bfr new_Jinkela_buffer_4049 (
        .din(new_Jinkela_wire_5600),
        .dout(new_Jinkela_wire_5601)
    );

    bfr new_Jinkela_buffer_3990 (
        .din(new_Jinkela_wire_5515),
        .dout(new_Jinkela_wire_5516)
    );

    bfr new_Jinkela_buffer_3960 (
        .din(new_Jinkela_wire_5485),
        .dout(new_Jinkela_wire_5486)
    );

    bfr new_Jinkela_buffer_4023 (
        .din(new_Jinkela_wire_5554),
        .dout(new_Jinkela_wire_5555)
    );

    bfr new_Jinkela_buffer_3991 (
        .din(new_Jinkela_wire_5516),
        .dout(new_Jinkela_wire_5517)
    );

    bfr new_Jinkela_buffer_3992 (
        .din(new_Jinkela_wire_5517),
        .dout(new_Jinkela_wire_5518)
    );

    bfr new_Jinkela_buffer_4024 (
        .din(new_Jinkela_wire_5555),
        .dout(new_Jinkela_wire_5556)
    );

    bfr new_Jinkela_buffer_4050 (
        .din(new_Jinkela_wire_5601),
        .dout(new_Jinkela_wire_5602)
    );

    bfr new_Jinkela_buffer_3993 (
        .din(new_Jinkela_wire_5518),
        .dout(new_Jinkela_wire_5519)
    );

    bfr new_Jinkela_buffer_4063 (
        .din(new_Jinkela_wire_5614),
        .dout(new_Jinkela_wire_5615)
    );

    bfr new_Jinkela_buffer_3994 (
        .din(new_Jinkela_wire_5519),
        .dout(new_Jinkela_wire_5520)
    );

    bfr new_Jinkela_buffer_4025 (
        .din(new_Jinkela_wire_5556),
        .dout(new_Jinkela_wire_5557)
    );

    bfr new_Jinkela_buffer_3995 (
        .din(new_Jinkela_wire_5520),
        .dout(new_Jinkela_wire_5521)
    );

    spl2 new_Jinkela_splitter_595 (
        .a(_0868_),
        .b(new_Jinkela_wire_5631),
        .c(new_Jinkela_wire_5633)
    );

    bfr new_Jinkela_buffer_3996 (
        .din(new_Jinkela_wire_5521),
        .dout(new_Jinkela_wire_5522)
    );

    bfr new_Jinkela_buffer_5121 (
        .din(new_Jinkela_wire_6976),
        .dout(new_Jinkela_wire_6977)
    );

    bfr new_Jinkela_buffer_2661 (
        .din(new_Jinkela_wire_3930),
        .dout(new_Jinkela_wire_3931)
    );

    bfr new_Jinkela_buffer_5139 (
        .din(new_Jinkela_wire_7002),
        .dout(new_Jinkela_wire_7003)
    );

    bfr new_Jinkela_buffer_2704 (
        .din(new_Jinkela_wire_3993),
        .dout(new_Jinkela_wire_3994)
    );

    bfr new_Jinkela_buffer_5122 (
        .din(new_Jinkela_wire_6977),
        .dout(new_Jinkela_wire_6978)
    );

    bfr new_Jinkela_buffer_2684 (
        .din(new_Jinkela_wire_3955),
        .dout(new_Jinkela_wire_3956)
    );

    bfr new_Jinkela_buffer_2662 (
        .din(new_Jinkela_wire_3931),
        .dout(new_Jinkela_wire_3932)
    );

    bfr new_Jinkela_buffer_5146 (
        .din(new_Jinkela_wire_7019),
        .dout(new_Jinkela_wire_7020)
    );

    bfr new_Jinkela_buffer_5123 (
        .din(new_Jinkela_wire_6978),
        .dout(new_Jinkela_wire_6979)
    );

    bfr new_Jinkela_buffer_2663 (
        .din(new_Jinkela_wire_3932),
        .dout(new_Jinkela_wire_3933)
    );

    bfr new_Jinkela_buffer_5140 (
        .din(new_Jinkela_wire_7003),
        .dout(new_Jinkela_wire_7004)
    );

    bfr new_Jinkela_buffer_5124 (
        .din(new_Jinkela_wire_6979),
        .dout(new_Jinkela_wire_6980)
    );

    spl2 new_Jinkela_splitter_480 (
        .a(new_Jinkela_wire_3956),
        .b(new_Jinkela_wire_3957),
        .c(new_Jinkela_wire_3958)
    );

    bfr new_Jinkela_buffer_2664 (
        .din(new_Jinkela_wire_3933),
        .dout(new_Jinkela_wire_3934)
    );

    bfr new_Jinkela_buffer_5195 (
        .din(new_net_2439),
        .dout(new_Jinkela_wire_7074)
    );

    bfr new_Jinkela_buffer_5125 (
        .din(new_Jinkela_wire_6980),
        .dout(new_Jinkela_wire_6981)
    );

    bfr new_Jinkela_buffer_2685 (
        .din(new_Jinkela_wire_3958),
        .dout(new_Jinkela_wire_3959)
    );

    bfr new_Jinkela_buffer_2665 (
        .din(new_Jinkela_wire_3934),
        .dout(new_Jinkela_wire_3935)
    );

    bfr new_Jinkela_buffer_5141 (
        .din(new_Jinkela_wire_7004),
        .dout(new_Jinkela_wire_7005)
    );

    bfr new_Jinkela_buffer_5126 (
        .din(new_Jinkela_wire_6981),
        .dout(new_Jinkela_wire_6982)
    );

    bfr new_Jinkela_buffer_2733 (
        .din(new_Jinkela_wire_4035),
        .dout(new_Jinkela_wire_4036)
    );

    bfr new_Jinkela_buffer_2666 (
        .din(new_Jinkela_wire_3935),
        .dout(new_Jinkela_wire_3936)
    );

    bfr new_Jinkela_buffer_5162 (
        .din(new_Jinkela_wire_7038),
        .dout(new_Jinkela_wire_7039)
    );

    bfr new_Jinkela_buffer_2705 (
        .din(new_Jinkela_wire_3994),
        .dout(new_Jinkela_wire_3995)
    );

    bfr new_Jinkela_buffer_5127 (
        .din(new_Jinkela_wire_6982),
        .dout(new_Jinkela_wire_6983)
    );

    bfr new_Jinkela_buffer_2667 (
        .din(new_Jinkela_wire_3936),
        .dout(new_Jinkela_wire_3937)
    );

    bfr new_Jinkela_buffer_5147 (
        .din(new_Jinkela_wire_7020),
        .dout(new_Jinkela_wire_7021)
    );

    bfr new_Jinkela_buffer_5128 (
        .din(new_Jinkela_wire_6983),
        .dout(new_Jinkela_wire_6984)
    );

    spl2 new_Jinkela_splitter_481 (
        .a(new_Jinkela_wire_3959),
        .b(new_Jinkela_wire_3960),
        .c(new_Jinkela_wire_3961)
    );

    bfr new_Jinkela_buffer_2668 (
        .din(new_Jinkela_wire_3937),
        .dout(new_Jinkela_wire_3938)
    );

    bfr new_Jinkela_buffer_5166 (
        .din(new_Jinkela_wire_7044),
        .dout(new_Jinkela_wire_7045)
    );

    spl2 new_Jinkela_splitter_722 (
        .a(new_Jinkela_wire_7039),
        .b(new_Jinkela_wire_7040),
        .c(new_Jinkela_wire_7041)
    );

    bfr new_Jinkela_buffer_5129 (
        .din(new_Jinkela_wire_6984),
        .dout(new_Jinkela_wire_6985)
    );

    bfr new_Jinkela_buffer_2686 (
        .din(new_Jinkela_wire_3961),
        .dout(new_Jinkela_wire_3962)
    );

    bfr new_Jinkela_buffer_2669 (
        .din(new_Jinkela_wire_3938),
        .dout(new_Jinkela_wire_3939)
    );

    bfr new_Jinkela_buffer_5148 (
        .din(new_Jinkela_wire_7021),
        .dout(new_Jinkela_wire_7022)
    );

    bfr new_Jinkela_buffer_5130 (
        .din(new_Jinkela_wire_6985),
        .dout(new_Jinkela_wire_6986)
    );

    bfr new_Jinkela_buffer_2670 (
        .din(new_Jinkela_wire_3939),
        .dout(new_Jinkela_wire_3940)
    );

    bfr new_Jinkela_buffer_2706 (
        .din(new_Jinkela_wire_3995),
        .dout(new_Jinkela_wire_3996)
    );

    bfr new_Jinkela_buffer_5149 (
        .din(new_Jinkela_wire_7022),
        .dout(new_Jinkela_wire_7023)
    );

    bfr new_Jinkela_buffer_2671 (
        .din(new_Jinkela_wire_3940),
        .dout(new_Jinkela_wire_3941)
    );

    bfr new_Jinkela_buffer_5163 (
        .din(new_Jinkela_wire_7041),
        .dout(new_Jinkela_wire_7042)
    );

    bfr new_Jinkela_buffer_2734 (
        .din(new_Jinkela_wire_4036),
        .dout(new_Jinkela_wire_4037)
    );

    bfr new_Jinkela_buffer_5150 (
        .din(new_Jinkela_wire_7023),
        .dout(new_Jinkela_wire_7024)
    );

    bfr new_Jinkela_buffer_2687 (
        .din(new_Jinkela_wire_3962),
        .dout(new_Jinkela_wire_3963)
    );

    spl3L new_Jinkela_splitter_723 (
        .a(_0735_),
        .d(new_Jinkela_wire_7078),
        .b(new_Jinkela_wire_7079),
        .c(new_Jinkela_wire_7080)
    );

    spl3L new_Jinkela_splitter_725 (
        .a(_0681_),
        .d(new_Jinkela_wire_7083),
        .b(new_Jinkela_wire_7084),
        .c(new_Jinkela_wire_7085)
    );

    bfr new_Jinkela_buffer_2707 (
        .din(new_Jinkela_wire_3996),
        .dout(new_Jinkela_wire_3997)
    );

    bfr new_Jinkela_buffer_5151 (
        .din(new_Jinkela_wire_7024),
        .dout(new_Jinkela_wire_7025)
    );

    spl2 new_Jinkela_splitter_482 (
        .a(new_Jinkela_wire_3963),
        .b(new_Jinkela_wire_3964),
        .c(new_Jinkela_wire_3965)
    );

    bfr new_Jinkela_buffer_5167 (
        .din(new_Jinkela_wire_7045),
        .dout(new_Jinkela_wire_7046)
    );

    bfr new_Jinkela_buffer_2688 (
        .din(new_Jinkela_wire_3965),
        .dout(new_Jinkela_wire_3966)
    );

    bfr new_Jinkela_buffer_5152 (
        .din(new_Jinkela_wire_7025),
        .dout(new_Jinkela_wire_7026)
    );

    bfr new_Jinkela_buffer_2766 (
        .din(new_net_2395),
        .dout(new_Jinkela_wire_4075)
    );

    bfr new_Jinkela_buffer_5164 (
        .din(new_Jinkela_wire_7042),
        .dout(new_Jinkela_wire_7043)
    );

    spl4L new_Jinkela_splitter_494 (
        .a(new_Jinkela_wire_4052),
        .d(new_Jinkela_wire_4053),
        .e(new_Jinkela_wire_4054),
        .b(new_Jinkela_wire_4055),
        .c(new_Jinkela_wire_4056)
    );

    bfr new_Jinkela_buffer_2708 (
        .din(new_Jinkela_wire_3997),
        .dout(new_Jinkela_wire_3998)
    );

    bfr new_Jinkela_buffer_5153 (
        .din(new_Jinkela_wire_7026),
        .dout(new_Jinkela_wire_7027)
    );

    bfr new_Jinkela_buffer_2689 (
        .din(new_Jinkela_wire_3966),
        .dout(new_Jinkela_wire_3967)
    );

    bfr new_Jinkela_buffer_5196 (
        .din(new_Jinkela_wire_7074),
        .dout(new_Jinkela_wire_7075)
    );

    bfr new_Jinkela_buffer_2735 (
        .din(new_Jinkela_wire_4037),
        .dout(new_Jinkela_wire_4038)
    );

    bfr new_Jinkela_buffer_5154 (
        .din(new_Jinkela_wire_7027),
        .dout(new_Jinkela_wire_7028)
    );

    spl2 new_Jinkela_splitter_483 (
        .a(new_Jinkela_wire_3967),
        .b(new_Jinkela_wire_3968),
        .c(new_Jinkela_wire_3969)
    );

    bfr new_Jinkela_buffer_5168 (
        .din(new_Jinkela_wire_7046),
        .dout(new_Jinkela_wire_7047)
    );

    bfr new_Jinkela_buffer_2690 (
        .din(new_Jinkela_wire_3969),
        .dout(new_Jinkela_wire_3970)
    );

    bfr new_Jinkela_buffer_5155 (
        .din(new_Jinkela_wire_7028),
        .dout(new_Jinkela_wire_7029)
    );

    bfr new_Jinkela_buffer_2709 (
        .din(new_Jinkela_wire_3998),
        .dout(new_Jinkela_wire_3999)
    );

    bfr new_Jinkela_buffer_5199 (
        .din(_0403_),
        .dout(new_Jinkela_wire_7086)
    );

    bfr new_Jinkela_buffer_5156 (
        .din(new_Jinkela_wire_7029),
        .dout(new_Jinkela_wire_7030)
    );

    spl2 new_Jinkela_splitter_484 (
        .a(new_Jinkela_wire_3970),
        .b(new_Jinkela_wire_3971),
        .c(new_Jinkela_wire_3972)
    );

    bfr new_Jinkela_buffer_5169 (
        .din(new_Jinkela_wire_7047),
        .dout(new_Jinkela_wire_7048)
    );

    bfr new_Jinkela_buffer_2691 (
        .din(new_Jinkela_wire_3972),
        .dout(new_Jinkela_wire_3973)
    );

    bfr new_Jinkela_buffer_5157 (
        .din(new_Jinkela_wire_7030),
        .dout(new_Jinkela_wire_7031)
    );

    bfr new_Jinkela_buffer_2747 (
        .din(new_Jinkela_wire_4050),
        .dout(new_Jinkela_wire_4051)
    );

    bfr new_Jinkela_buffer_2710 (
        .din(new_Jinkela_wire_3999),
        .dout(new_Jinkela_wire_4000)
    );

    bfr new_Jinkela_buffer_5197 (
        .din(new_Jinkela_wire_7075),
        .dout(new_Jinkela_wire_7076)
    );

    bfr new_Jinkela_buffer_2736 (
        .din(new_Jinkela_wire_4038),
        .dout(new_Jinkela_wire_4039)
    );

    bfr new_Jinkela_buffer_5158 (
        .din(new_Jinkela_wire_7031),
        .dout(new_Jinkela_wire_7032)
    );

    spl2 new_Jinkela_splitter_485 (
        .a(new_Jinkela_wire_3973),
        .b(new_Jinkela_wire_3974),
        .c(new_Jinkela_wire_3975)
    );

    bfr new_Jinkela_buffer_5170 (
        .din(new_Jinkela_wire_7048),
        .dout(new_Jinkela_wire_7049)
    );

    bfr new_Jinkela_buffer_2692 (
        .din(new_Jinkela_wire_3975),
        .dout(new_Jinkela_wire_3976)
    );

    bfr new_Jinkela_buffer_5159 (
        .din(new_Jinkela_wire_7032),
        .dout(new_Jinkela_wire_7033)
    );

    bfr new_Jinkela_buffer_2711 (
        .din(new_Jinkela_wire_4000),
        .dout(new_Jinkela_wire_4001)
    );

    bfr new_Jinkela_buffer_2855 (
        .din(new_Jinkela_wire_4172),
        .dout(new_Jinkela_wire_4173)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_2095),
        .dout(new_Jinkela_wire_2096)
    );

    bfr new_Jinkela_buffer_2826 (
        .din(new_Jinkela_wire_4140),
        .dout(new_Jinkela_wire_4141)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(new_Jinkela_wire_2053),
        .dout(new_Jinkela_wire_2054)
    );

    bfr new_Jinkela_buffer_2846 (
        .din(new_Jinkela_wire_4160),
        .dout(new_Jinkela_wire_4161)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_2077),
        .dout(new_Jinkela_wire_2078)
    );

    bfr new_Jinkela_buffer_2827 (
        .din(new_Jinkela_wire_4141),
        .dout(new_Jinkela_wire_4142)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_2054),
        .dout(new_Jinkela_wire_2055)
    );

    bfr new_Jinkela_buffer_2872 (
        .din(new_net_2457),
        .dout(new_Jinkela_wire_4196)
    );

    spl2 new_Jinkela_splitter_347 (
        .a(_1095_),
        .b(new_Jinkela_wire_2120),
        .c(new_Jinkela_wire_2121)
    );

    bfr new_Jinkela_buffer_2828 (
        .din(new_Jinkela_wire_4142),
        .dout(new_Jinkela_wire_4143)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(_0469_),
        .dout(new_Jinkela_wire_2122)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_2055),
        .dout(new_Jinkela_wire_2056)
    );

    bfr new_Jinkela_buffer_2847 (
        .din(new_Jinkela_wire_4161),
        .dout(new_Jinkela_wire_4162)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(new_Jinkela_wire_2078),
        .dout(new_Jinkela_wire_2079)
    );

    bfr new_Jinkela_buffer_2829 (
        .din(new_Jinkela_wire_4143),
        .dout(new_Jinkela_wire_4144)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(new_Jinkela_wire_2056),
        .dout(new_Jinkela_wire_2057)
    );

    bfr new_Jinkela_buffer_2858 (
        .din(new_Jinkela_wire_4179),
        .dout(new_Jinkela_wire_4180)
    );

    bfr new_Jinkela_buffer_2856 (
        .din(new_Jinkela_wire_4173),
        .dout(new_Jinkela_wire_4174)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_2096),
        .dout(new_Jinkela_wire_2097)
    );

    bfr new_Jinkela_buffer_2830 (
        .din(new_Jinkela_wire_4144),
        .dout(new_Jinkela_wire_4145)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_2057),
        .dout(new_Jinkela_wire_2058)
    );

    bfr new_Jinkela_buffer_2848 (
        .din(new_Jinkela_wire_4162),
        .dout(new_Jinkela_wire_4163)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(new_Jinkela_wire_2079),
        .dout(new_Jinkela_wire_2080)
    );

    bfr new_Jinkela_buffer_2831 (
        .din(new_Jinkela_wire_4145),
        .dout(new_Jinkela_wire_4146)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_2058),
        .dout(new_Jinkela_wire_2059)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_2118),
        .dout(new_Jinkela_wire_2119)
    );

    bfr new_Jinkela_buffer_2832 (
        .din(new_Jinkela_wire_4146),
        .dout(new_Jinkela_wire_4147)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_2059),
        .dout(new_Jinkela_wire_2060)
    );

    bfr new_Jinkela_buffer_2849 (
        .din(new_Jinkela_wire_4163),
        .dout(new_Jinkela_wire_4164)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_2080),
        .dout(new_Jinkela_wire_2081)
    );

    bfr new_Jinkela_buffer_2833 (
        .din(new_Jinkela_wire_4147),
        .dout(new_Jinkela_wire_4148)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(new_Jinkela_wire_2060),
        .dout(new_Jinkela_wire_2061)
    );

    spl2 new_Jinkela_splitter_501 (
        .a(_1054_),
        .b(new_Jinkela_wire_4194),
        .c(new_Jinkela_wire_4195)
    );

    spl2 new_Jinkela_splitter_499 (
        .a(new_Jinkela_wire_4174),
        .b(new_Jinkela_wire_4175),
        .c(new_Jinkela_wire_4176)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(new_Jinkela_wire_2097),
        .dout(new_Jinkela_wire_2098)
    );

    bfr new_Jinkela_buffer_2834 (
        .din(new_Jinkela_wire_4148),
        .dout(new_Jinkela_wire_4149)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(new_Jinkela_wire_2061),
        .dout(new_Jinkela_wire_2062)
    );

    bfr new_Jinkela_buffer_2850 (
        .din(new_Jinkela_wire_4164),
        .dout(new_Jinkela_wire_4165)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_2081),
        .dout(new_Jinkela_wire_2082)
    );

    bfr new_Jinkela_buffer_2835 (
        .din(new_Jinkela_wire_4149),
        .dout(new_Jinkela_wire_4150)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(new_Jinkela_wire_2062),
        .dout(new_Jinkela_wire_2063)
    );

    bfr new_Jinkela_buffer_2873 (
        .din(new_Jinkela_wire_4196),
        .dout(new_Jinkela_wire_4197)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_net_2479),
        .dout(new_Jinkela_wire_2156)
    );

    bfr new_Jinkela_buffer_2836 (
        .din(new_Jinkela_wire_4150),
        .dout(new_Jinkela_wire_4151)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_2122),
        .dout(new_Jinkela_wire_2123)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_2082),
        .dout(new_Jinkela_wire_2083)
    );

    bfr new_Jinkela_buffer_2851 (
        .din(new_Jinkela_wire_4165),
        .dout(new_Jinkela_wire_4166)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_2098),
        .dout(new_Jinkela_wire_2099)
    );

    bfr new_Jinkela_buffer_2837 (
        .din(new_Jinkela_wire_4151),
        .dout(new_Jinkela_wire_4152)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(new_Jinkela_wire_2083),
        .dout(new_Jinkela_wire_2084)
    );

    bfr new_Jinkela_buffer_2859 (
        .din(new_Jinkela_wire_4180),
        .dout(new_Jinkela_wire_4181)
    );

    bfr new_Jinkela_buffer_2838 (
        .din(new_Jinkela_wire_4152),
        .dout(new_Jinkela_wire_4153)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_2084),
        .dout(new_Jinkela_wire_2085)
    );

    bfr new_Jinkela_buffer_2878 (
        .din(new_net_2475),
        .dout(new_Jinkela_wire_4204)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(new_Jinkela_wire_2099),
        .dout(new_Jinkela_wire_2100)
    );

    bfr new_Jinkela_buffer_2839 (
        .din(new_Jinkela_wire_4153),
        .dout(new_Jinkela_wire_4154)
    );

    spl2 new_Jinkela_splitter_348 (
        .a(_0192_),
        .b(new_Jinkela_wire_2154),
        .c(new_Jinkela_wire_2155)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_2100),
        .dout(new_Jinkela_wire_2101)
    );

    bfr new_Jinkela_buffer_2860 (
        .din(new_Jinkela_wire_4181),
        .dout(new_Jinkela_wire_4182)
    );

    bfr new_Jinkela_buffer_2875 (
        .din(_0165_),
        .dout(new_Jinkela_wire_4199)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(new_Jinkela_wire_2156),
        .dout(new_Jinkela_wire_2157)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_2101),
        .dout(new_Jinkela_wire_2102)
    );

    bfr new_Jinkela_buffer_2861 (
        .din(new_Jinkela_wire_4182),
        .dout(new_Jinkela_wire_4183)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_2123),
        .dout(new_Jinkela_wire_2124)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_2102),
        .dout(new_Jinkela_wire_2103)
    );

    bfr new_Jinkela_buffer_2862 (
        .din(new_Jinkela_wire_4183),
        .dout(new_Jinkela_wire_4184)
    );

    bfr new_Jinkela_buffer_2874 (
        .din(new_Jinkela_wire_4197),
        .dout(new_Jinkela_wire_4198)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_2103),
        .dout(new_Jinkela_wire_2104)
    );

    bfr new_Jinkela_buffer_2863 (
        .din(new_Jinkela_wire_4184),
        .dout(new_Jinkela_wire_4185)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_2124),
        .dout(new_Jinkela_wire_2125)
    );

    bfr new_Jinkela_buffer_2893 (
        .din(new_net_2503),
        .dout(new_Jinkela_wire_4219)
    );

    bfr new_Jinkela_buffer_2876 (
        .din(new_Jinkela_wire_4199),
        .dout(new_Jinkela_wire_4200)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(new_Jinkela_wire_2104),
        .dout(new_Jinkela_wire_2105)
    );

    bfr new_Jinkela_buffer_2864 (
        .din(new_Jinkela_wire_4185),
        .dout(new_Jinkela_wire_4186)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_net_2495),
        .dout(new_Jinkela_wire_2160)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(new_Jinkela_wire_2105),
        .dout(new_Jinkela_wire_2106)
    );

    bfr new_Jinkela_buffer_2865 (
        .din(new_Jinkela_wire_4186),
        .dout(new_Jinkela_wire_4187)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_2125),
        .dout(new_Jinkela_wire_2126)
    );

    bfr new_Jinkela_buffer_2879 (
        .din(new_Jinkela_wire_4204),
        .dout(new_Jinkela_wire_4205)
    );

    bfr new_Jinkela_buffer_2877 (
        .din(new_Jinkela_wire_4200),
        .dout(new_Jinkela_wire_4201)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_2106),
        .dout(new_Jinkela_wire_2107)
    );

    bfr new_Jinkela_buffer_2866 (
        .din(new_Jinkela_wire_4187),
        .dout(new_Jinkela_wire_4188)
    );

    spl2 new_Jinkela_splitter_349 (
        .a(_0004_),
        .b(new_Jinkela_wire_2197),
        .c(new_Jinkela_wire_2198)
    );

    and_bi _2498_ (
        .a(new_Jinkela_wire_122),
        .b(new_Jinkela_wire_5807),
        .c(_0488_)
    );

    bfr new_Jinkela_buffer_4027 (
        .din(new_Jinkela_wire_5558),
        .dout(new_Jinkela_wire_5559)
    );

    or_bi _1781_ (
        .a(_1069_),
        .b(_1068_),
        .c(_1070_)
    );

    and_bi _2499_ (
        .a(new_Jinkela_wire_1389),
        .b(new_Jinkela_wire_7873),
        .c(_0489_)
    );

    bfr new_Jinkela_buffer_3997 (
        .din(new_Jinkela_wire_5522),
        .dout(new_Jinkela_wire_5523)
    );

    and_bi _1782_ (
        .a(new_Jinkela_wire_7886),
        .b(new_Jinkela_wire_6676),
        .c(_1071_)
    );

    or_bb _2500_ (
        .a(_0489_),
        .b(_0488_),
        .c(_0490_)
    );

    or_bi _1783_ (
        .a(new_Jinkela_wire_1983),
        .b(new_Jinkela_wire_5305),
        .c(_1072_)
    );

    bfr new_Jinkela_buffer_4094 (
        .din(_0456_),
        .dout(new_Jinkela_wire_5652)
    );

    or_bb _2501_ (
        .a(new_Jinkela_wire_5857),
        .b(_0487_),
        .c(new_net_2405)
    );

    bfr new_Jinkela_buffer_3998 (
        .din(new_Jinkela_wire_5523),
        .dout(new_Jinkela_wire_5524)
    );

    and_bi _1784_ (
        .a(new_Jinkela_wire_1984),
        .b(new_Jinkela_wire_5306),
        .c(_1073_)
    );

    or_bi _2502_ (
        .a(new_Jinkela_wire_387),
        .b(new_Jinkela_wire_6994),
        .c(_0491_)
    );

    bfr new_Jinkela_buffer_4051 (
        .din(new_Jinkela_wire_5602),
        .dout(new_Jinkela_wire_5603)
    );

    or_bi _1785_ (
        .a(_1073_),
        .b(_1072_),
        .c(_1074_)
    );

    and_bb _2503_ (
        .a(new_Jinkela_wire_6907),
        .b(new_Jinkela_wire_385),
        .c(_0492_)
    );

    bfr new_Jinkela_buffer_3999 (
        .din(new_Jinkela_wire_5524),
        .dout(new_Jinkela_wire_5525)
    );

    or_bi _1786_ (
        .a(new_Jinkela_wire_7138),
        .b(new_Jinkela_wire_3629),
        .c(_1075_)
    );

    or_bb _2504_ (
        .a(_0492_),
        .b(new_Jinkela_wire_3979),
        .c(_0493_)
    );

    bfr new_Jinkela_buffer_4026 (
        .din(new_Jinkela_wire_5557),
        .dout(new_Jinkela_wire_5558)
    );

    inv _1787_ (
        .din(new_Jinkela_wire_123),
        .dout(_1076_)
    );

    bfr new_Jinkela_buffer_4028 (
        .din(new_Jinkela_wire_5559),
        .dout(new_Jinkela_wire_5560)
    );

    and_bi _2505_ (
        .a(_0491_),
        .b(_0493_),
        .c(_0494_)
    );

    bfr new_Jinkela_buffer_4000 (
        .din(new_Jinkela_wire_5525),
        .dout(new_Jinkela_wire_5526)
    );

    and_bi _1788_ (
        .a(new_Jinkela_wire_7139),
        .b(new_Jinkela_wire_3630),
        .c(_1077_)
    );

    and_bi _2506_ (
        .a(new_Jinkela_wire_227),
        .b(new_Jinkela_wire_5808),
        .c(_0495_)
    );

    bfr new_Jinkela_buffer_4064 (
        .din(new_Jinkela_wire_5615),
        .dout(new_Jinkela_wire_5616)
    );

    or_bb _1789_ (
        .a(_1077_),
        .b(new_Jinkela_wire_6282),
        .c(_1078_)
    );

    bfr new_Jinkela_buffer_4029 (
        .din(new_Jinkela_wire_5560),
        .dout(new_Jinkela_wire_5561)
    );

    and_bi _2507_ (
        .a(new_Jinkela_wire_1243),
        .b(new_Jinkela_wire_7874),
        .c(_0496_)
    );

    bfr new_Jinkela_buffer_4001 (
        .din(new_Jinkela_wire_5526),
        .dout(new_Jinkela_wire_5527)
    );

    and_bi _1790_ (
        .a(new_Jinkela_wire_5192),
        .b(_1078_),
        .c(_1079_)
    );

    or_bb _2508_ (
        .a(_0496_),
        .b(_0495_),
        .c(_0497_)
    );

    or_bb _1791_ (
        .a(_1079_),
        .b(_1061_),
        .c(_1080_)
    );

    bfr new_Jinkela_buffer_4052 (
        .din(new_Jinkela_wire_5603),
        .dout(new_Jinkela_wire_5604)
    );

    or_bb _2509_ (
        .a(new_Jinkela_wire_1848),
        .b(_0494_),
        .c(new_net_2511)
    );

    bfr new_Jinkela_buffer_4002 (
        .din(new_Jinkela_wire_5527),
        .dout(new_Jinkela_wire_5528)
    );

    or_bi _1792_ (
        .a(new_Jinkela_wire_1889),
        .b(new_Jinkela_wire_6100),
        .c(_1081_)
    );

    and_bi _2510_ (
        .a(new_Jinkela_wire_6906),
        .b(new_Jinkela_wire_1667),
        .c(_0498_)
    );

    and_bb _1793_ (
        .a(new_Jinkela_wire_3627),
        .b(new_Jinkela_wire_6243),
        .c(_1082_)
    );

    and_bi _2511_ (
        .a(new_Jinkela_wire_6993),
        .b(new_Jinkela_wire_491),
        .c(_0499_)
    );

    bfr new_Jinkela_buffer_4003 (
        .din(new_Jinkela_wire_5528),
        .dout(new_Jinkela_wire_5529)
    );

    or_bb _1794_ (
        .a(_1082_),
        .b(new_Jinkela_wire_7604),
        .c(_1083_)
    );

    or_bb _2512_ (
        .a(_0499_),
        .b(new_Jinkela_wire_1745),
        .c(_0500_)
    );

    or_bb _1795_ (
        .a(new_Jinkela_wire_7018),
        .b(new_Jinkela_wire_3064),
        .c(_1084_)
    );

    or_bb _2513_ (
        .a(_0500_),
        .b(new_Jinkela_wire_7994),
        .c(_0501_)
    );

    bfr new_Jinkela_buffer_4004 (
        .din(new_Jinkela_wire_5529),
        .dout(new_Jinkela_wire_5530)
    );

    and_bi _1796_ (
        .a(new_Jinkela_wire_3063),
        .b(new_Jinkela_wire_6025),
        .c(_1085_)
    );

    and_bi _2514_ (
        .a(new_Jinkela_wire_1343),
        .b(new_Jinkela_wire_7916),
        .c(_0502_)
    );

    or_bi _1797_ (
        .a(new_Jinkela_wire_2305),
        .b(new_Jinkela_wire_5906),
        .c(_1086_)
    );

    bfr new_Jinkela_buffer_4053 (
        .din(new_Jinkela_wire_5604),
        .dout(new_Jinkela_wire_5605)
    );

    and_bi _2515_ (
        .a(new_Jinkela_wire_330),
        .b(new_Jinkela_wire_6132),
        .c(_0503_)
    );

    bfr new_Jinkela_buffer_4005 (
        .din(new_Jinkela_wire_5530),
        .dout(new_Jinkela_wire_5531)
    );

    and_bi _1798_ (
        .a(new_Jinkela_wire_2912),
        .b(new_Jinkela_wire_3628),
        .c(_1087_)
    );

    or_bb _2516_ (
        .a(_0503_),
        .b(_0502_),
        .c(_0504_)
    );

    bfr new_Jinkela_buffer_4031 (
        .din(new_Jinkela_wire_5562),
        .dout(new_Jinkela_wire_5563)
    );

    or_bb _1799_ (
        .a(_1087_),
        .b(new_Jinkela_wire_6071),
        .c(_1088_)
    );

    and_bi _2517_ (
        .a(_0501_),
        .b(new_Jinkela_wire_6749),
        .c(_0505_)
    );

    bfr new_Jinkela_buffer_4006 (
        .din(new_Jinkela_wire_5531),
        .dout(new_Jinkela_wire_5532)
    );

    or_bb _1800_ (
        .a(new_Jinkela_wire_3534),
        .b(new_Jinkela_wire_2089),
        .c(_1089_)
    );

    and_bi _2518_ (
        .a(new_Jinkela_wire_689),
        .b(_0505_),
        .c(new_net_2361)
    );

    bfr new_Jinkela_buffer_4030 (
        .din(new_Jinkela_wire_5561),
        .dout(new_Jinkela_wire_5562)
    );

    and_bi _1801_ (
        .a(new_Jinkela_wire_5907),
        .b(new_Jinkela_wire_2306),
        .c(_1090_)
    );

    bfr new_Jinkela_buffer_4065 (
        .din(new_Jinkela_wire_5616),
        .dout(new_Jinkela_wire_5617)
    );

    and_bi _2519_ (
        .a(new_Jinkela_wire_495),
        .b(new_Jinkela_wire_1617),
        .c(_0506_)
    );

    bfr new_Jinkela_buffer_4007 (
        .din(new_Jinkela_wire_5532),
        .dout(new_Jinkela_wire_5533)
    );

    and_bi _1802_ (
        .a(new_Jinkela_wire_3535),
        .b(new_Jinkela_wire_7203),
        .c(_1091_)
    );

    and_bi _2520_ (
        .a(new_Jinkela_wire_5362),
        .b(new_Jinkela_wire_497),
        .c(_0507_)
    );

    and_bi _1803_ (
        .a(_1089_),
        .b(_1091_),
        .c(_1092_)
    );

    bfr new_Jinkela_buffer_4076 (
        .din(new_Jinkela_wire_5627),
        .dout(new_Jinkela_wire_5628)
    );

    or_bb _2521_ (
        .a(_0507_),
        .b(new_Jinkela_wire_1751),
        .c(_0508_)
    );

    bfr new_Jinkela_buffer_4008 (
        .din(new_Jinkela_wire_5533),
        .dout(new_Jinkela_wire_5534)
    );

    and_bi _1804_ (
        .a(new_Jinkela_wire_6987),
        .b(new_Jinkela_wire_3087),
        .c(_1093_)
    );

    or_bb _2522_ (
        .a(_0508_),
        .b(new_Jinkela_wire_2119),
        .c(_0509_)
    );

    bfr new_Jinkela_buffer_4032 (
        .din(new_Jinkela_wire_5563),
        .dout(new_Jinkela_wire_5564)
    );

    and_bi _1805_ (
        .a(new_Jinkela_wire_3088),
        .b(new_Jinkela_wire_6988),
        .c(_1094_)
    );

    and_bi _2523_ (
        .a(new_Jinkela_wire_1575),
        .b(new_Jinkela_wire_7915),
        .c(_0510_)
    );

    bfr new_Jinkela_buffer_4009 (
        .din(new_Jinkela_wire_5534),
        .dout(new_Jinkela_wire_5535)
    );

    or_bb _1806_ (
        .a(_1094_),
        .b(_1093_),
        .c(_1095_)
    );

    and_bi _2524_ (
        .a(new_Jinkela_wire_961),
        .b(new_Jinkela_wire_6137),
        .c(_0511_)
    );

    bfr new_Jinkela_buffer_4054 (
        .din(new_Jinkela_wire_5605),
        .dout(new_Jinkela_wire_5606)
    );

    or_bi _1807_ (
        .a(new_Jinkela_wire_2120),
        .b(new_Jinkela_wire_1914),
        .c(_1096_)
    );

    or_bb _2525_ (
        .a(_0511_),
        .b(_0510_),
        .c(_0512_)
    );

    bfr new_Jinkela_buffer_4010 (
        .din(new_Jinkela_wire_5535),
        .dout(new_Jinkela_wire_5536)
    );

    and_bb _1808_ (
        .a(new_Jinkela_wire_6102),
        .b(new_Jinkela_wire_6239),
        .c(_1097_)
    );

    and_bi _2526_ (
        .a(_0509_),
        .b(new_Jinkela_wire_1787),
        .c(_0513_)
    );

    bfr new_Jinkela_buffer_4033 (
        .din(new_Jinkela_wire_5564),
        .dout(new_Jinkela_wire_5565)
    );

    and_ii _1809_ (
        .a(new_Jinkela_wire_1755),
        .b(new_Jinkela_wire_7205),
        .c(_1098_)
    );

    and_bi _2527_ (
        .a(new_Jinkela_wire_696),
        .b(_0513_),
        .c(new_net_2381)
    );

    bfr new_Jinkela_buffer_4011 (
        .din(new_Jinkela_wire_5536),
        .dout(new_Jinkela_wire_5537)
    );

    or_bi _1810_ (
        .a(new_Jinkela_wire_6043),
        .b(new_Jinkela_wire_5254),
        .c(_1099_)
    );

    and_bi _2528_ (
        .a(new_Jinkela_wire_5777),
        .b(new_Jinkela_wire_1671),
        .c(_0514_)
    );

    and_bi _1811_ (
        .a(new_Jinkela_wire_6044),
        .b(new_Jinkela_wire_5255),
        .c(_1100_)
    );

    and_bi _2529_ (
        .a(new_Jinkela_wire_6793),
        .b(new_Jinkela_wire_498),
        .c(_0515_)
    );

    bfr new_Jinkela_buffer_4012 (
        .din(new_Jinkela_wire_5537),
        .dout(new_Jinkela_wire_5538)
    );

    or_bi _1812_ (
        .a(_1100_),
        .b(_1099_),
        .c(_1101_)
    );

    or_bb _2530_ (
        .a(_0515_),
        .b(new_Jinkela_wire_1750),
        .c(_0516_)
    );

    bfr new_Jinkela_buffer_4034 (
        .din(new_Jinkela_wire_5565),
        .dout(new_Jinkela_wire_5566)
    );

    or_bb _1813_ (
        .a(new_Jinkela_wire_2411),
        .b(new_Jinkela_wire_2086),
        .c(_1102_)
    );

    or_bb _2531_ (
        .a(_0516_),
        .b(new_Jinkela_wire_1979),
        .c(_0517_)
    );

    bfr new_Jinkela_buffer_4013 (
        .din(new_Jinkela_wire_5538),
        .dout(new_Jinkela_wire_5539)
    );

    and_bi _1814_ (
        .a(new_Jinkela_wire_2412),
        .b(new_Jinkela_wire_7200),
        .c(_1103_)
    );

    and_bi _2532_ (
        .a(new_Jinkela_wire_1275),
        .b(new_Jinkela_wire_6134),
        .c(_0518_)
    );

    and_bi _1815_ (
        .a(_1102_),
        .b(_1103_),
        .c(_1104_)
    );

    bfr new_Jinkela_buffer_4055 (
        .din(new_Jinkela_wire_5606),
        .dout(new_Jinkela_wire_5607)
    );

    and_bi _2533_ (
        .a(new_Jinkela_wire_1359),
        .b(new_Jinkela_wire_7925),
        .c(_0519_)
    );

    bfr new_Jinkela_buffer_4014 (
        .din(new_Jinkela_wire_5539),
        .dout(new_Jinkela_wire_5540)
    );

    or_bi _1816_ (
        .a(new_Jinkela_wire_2942),
        .b(new_Jinkela_wire_6949),
        .c(_1105_)
    );

    or_bb _2534_ (
        .a(_0519_),
        .b(_0518_),
        .c(_0520_)
    );

    spl2 new_Jinkela_splitter_585 (
        .a(new_Jinkela_wire_5566),
        .b(new_Jinkela_wire_5567),
        .c(new_Jinkela_wire_5568)
    );

    and_bi _1817_ (
        .a(new_Jinkela_wire_2943),
        .b(new_Jinkela_wire_6950),
        .c(_1106_)
    );

    and_bi _2535_ (
        .a(_0517_),
        .b(new_Jinkela_wire_2684),
        .c(_0521_)
    );

    bfr new_Jinkela_buffer_4015 (
        .din(new_Jinkela_wire_5540),
        .dout(new_Jinkela_wire_5541)
    );

    or_bb _1818_ (
        .a(_1106_),
        .b(new_Jinkela_wire_1908),
        .c(_1107_)
    );

    and_bi _2536_ (
        .a(new_Jinkela_wire_698),
        .b(_0521_),
        .c(new_net_2395)
    );

    bfr new_Jinkela_buffer_4035 (
        .din(new_Jinkela_wire_5568),
        .dout(new_Jinkela_wire_5569)
    );

    or_bi _1819_ (
        .a(_1107_),
        .b(new_Jinkela_wire_5394),
        .c(_1108_)
    );

    and_bi _2537_ (
        .a(new_Jinkela_wire_3618),
        .b(new_Jinkela_wire_499),
        .c(_0522_)
    );

    bfr new_Jinkela_buffer_4016 (
        .din(new_Jinkela_wire_5541),
        .dout(new_Jinkela_wire_5542)
    );

    or_ii _1820_ (
        .a(new_Jinkela_wire_1683),
        .b(new_Jinkela_wire_6279),
        .c(_1109_)
    );

    and_bi _2538_ (
        .a(new_Jinkela_wire_5004),
        .b(new_Jinkela_wire_1648),
        .c(_0523_)
    );

    and_bi _1821_ (
        .a(_1096_),
        .b(new_Jinkela_wire_7823),
        .c(_1110_)
    );

    bfr new_Jinkela_buffer_4066 (
        .din(new_Jinkela_wire_5617),
        .dout(new_Jinkela_wire_5618)
    );

    or_bb _2539_ (
        .a(_0523_),
        .b(new_Jinkela_wire_1725),
        .c(_0524_)
    );

    bfr new_Jinkela_buffer_4017 (
        .din(new_Jinkela_wire_5542),
        .dout(new_Jinkela_wire_5543)
    );

    and_bi _1822_ (
        .a(new_Jinkela_wire_3161),
        .b(new_Jinkela_wire_1907),
        .c(_1111_)
    );

    bfr new_Jinkela_buffer_5099 (
        .din(new_Jinkela_wire_6954),
        .dout(new_Jinkela_wire_6955)
    );

    bfr new_Jinkela_buffer_5094 (
        .din(new_Jinkela_wire_6945),
        .dout(new_Jinkela_wire_6946)
    );

    bfr new_Jinkela_buffer_5132 (
        .din(new_Jinkela_wire_6995),
        .dout(new_Jinkela_wire_6996)
    );

    bfr new_Jinkela_buffer_5102 (
        .din(new_Jinkela_wire_6957),
        .dout(new_Jinkela_wire_6958)
    );

    bfr new_Jinkela_buffer_5095 (
        .din(new_Jinkela_wire_6946),
        .dout(new_Jinkela_wire_6947)
    );

    bfr new_Jinkela_buffer_5131 (
        .din(new_Jinkela_wire_6989),
        .dout(new_Jinkela_wire_6990)
    );

    bfr new_Jinkela_buffer_5096 (
        .din(new_Jinkela_wire_6947),
        .dout(new_Jinkela_wire_6948)
    );

    bfr new_Jinkela_buffer_5142 (
        .din(_0821_),
        .dout(new_Jinkela_wire_7006)
    );

    bfr new_Jinkela_buffer_5103 (
        .din(new_Jinkela_wire_6958),
        .dout(new_Jinkela_wire_6959)
    );

    bfr new_Jinkela_buffer_5143 (
        .din(new_Jinkela_wire_7006),
        .dout(new_Jinkela_wire_7007)
    );

    spl4L new_Jinkela_splitter_716 (
        .a(new_Jinkela_wire_6991),
        .d(new_Jinkela_wire_6992),
        .e(new_Jinkela_wire_6993),
        .b(new_Jinkela_wire_6994),
        .c(new_Jinkela_wire_6995)
    );

    bfr new_Jinkela_buffer_5104 (
        .din(new_Jinkela_wire_6959),
        .dout(new_Jinkela_wire_6960)
    );

    bfr new_Jinkela_buffer_5105 (
        .din(new_Jinkela_wire_6960),
        .dout(new_Jinkela_wire_6961)
    );

    spl2 new_Jinkela_splitter_718 (
        .a(_0795_),
        .b(new_Jinkela_wire_7012),
        .c(new_Jinkela_wire_7013)
    );

    bfr new_Jinkela_buffer_5106 (
        .din(new_Jinkela_wire_6961),
        .dout(new_Jinkela_wire_6962)
    );

    bfr new_Jinkela_buffer_5107 (
        .din(new_Jinkela_wire_6962),
        .dout(new_Jinkela_wire_6963)
    );

    bfr new_Jinkela_buffer_5108 (
        .din(new_Jinkela_wire_6963),
        .dout(new_Jinkela_wire_6964)
    );

    spl4L new_Jinkela_splitter_717 (
        .a(new_Jinkela_wire_7007),
        .d(new_Jinkela_wire_7008),
        .e(new_Jinkela_wire_7009),
        .b(new_Jinkela_wire_7010),
        .c(new_Jinkela_wire_7011)
    );

    bfr new_Jinkela_buffer_5109 (
        .din(new_Jinkela_wire_6964),
        .dout(new_Jinkela_wire_6965)
    );

    bfr new_Jinkela_buffer_5133 (
        .din(new_Jinkela_wire_6996),
        .dout(new_Jinkela_wire_6997)
    );

    bfr new_Jinkela_buffer_5110 (
        .din(new_Jinkela_wire_6965),
        .dout(new_Jinkela_wire_6966)
    );

    bfr new_Jinkela_buffer_5145 (
        .din(new_Jinkela_wire_7014),
        .dout(new_Jinkela_wire_7015)
    );

    bfr new_Jinkela_buffer_5111 (
        .din(new_Jinkela_wire_6966),
        .dout(new_Jinkela_wire_6967)
    );

    bfr new_Jinkela_buffer_5134 (
        .din(new_Jinkela_wire_6997),
        .dout(new_Jinkela_wire_6998)
    );

    bfr new_Jinkela_buffer_5112 (
        .din(new_Jinkela_wire_6967),
        .dout(new_Jinkela_wire_6968)
    );

    bfr new_Jinkela_buffer_5144 (
        .din(_0470_),
        .dout(new_Jinkela_wire_7014)
    );

    bfr new_Jinkela_buffer_5113 (
        .din(new_Jinkela_wire_6968),
        .dout(new_Jinkela_wire_6969)
    );

    bfr new_Jinkela_buffer_5135 (
        .din(new_Jinkela_wire_6998),
        .dout(new_Jinkela_wire_6999)
    );

    bfr new_Jinkela_buffer_5114 (
        .din(new_Jinkela_wire_6969),
        .dout(new_Jinkela_wire_6970)
    );

    spl3L new_Jinkela_splitter_721 (
        .a(_0638_),
        .d(new_Jinkela_wire_7036),
        .b(new_Jinkela_wire_7037),
        .c(new_Jinkela_wire_7038)
    );

    bfr new_Jinkela_buffer_5115 (
        .din(new_Jinkela_wire_6970),
        .dout(new_Jinkela_wire_6971)
    );

    bfr new_Jinkela_buffer_5136 (
        .din(new_Jinkela_wire_6999),
        .dout(new_Jinkela_wire_7000)
    );

    bfr new_Jinkela_buffer_5116 (
        .din(new_Jinkela_wire_6971),
        .dout(new_Jinkela_wire_6972)
    );

    spl2 new_Jinkela_splitter_719 (
        .a(_0965_),
        .b(new_Jinkela_wire_7016),
        .c(new_Jinkela_wire_7017)
    );

    spl2 new_Jinkela_splitter_720 (
        .a(new_Jinkela_wire_7017),
        .b(new_Jinkela_wire_7018),
        .c(new_Jinkela_wire_7019)
    );

    bfr new_Jinkela_buffer_5117 (
        .din(new_Jinkela_wire_6972),
        .dout(new_Jinkela_wire_6973)
    );

    bfr new_Jinkela_buffer_5137 (
        .din(new_Jinkela_wire_7000),
        .dout(new_Jinkela_wire_7001)
    );

    bfr new_Jinkela_buffer_5118 (
        .din(new_Jinkela_wire_6973),
        .dout(new_Jinkela_wire_6974)
    );

    bfr new_Jinkela_buffer_5165 (
        .din(new_net_2499),
        .dout(new_Jinkela_wire_7044)
    );

    bfr new_Jinkela_buffer_5119 (
        .din(new_Jinkela_wire_6974),
        .dout(new_Jinkela_wire_6975)
    );

    bfr new_Jinkela_buffer_5138 (
        .din(new_Jinkela_wire_7001),
        .dout(new_Jinkela_wire_7002)
    );

    bfr new_Jinkela_buffer_5120 (
        .din(new_Jinkela_wire_6975),
        .dout(new_Jinkela_wire_6976)
    );

    spl4L new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_405),
        .d(new_Jinkela_wire_406),
        .e(new_Jinkela_wire_407),
        .b(new_Jinkela_wire_411),
        .c(new_Jinkela_wire_416)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    bfr new_Jinkela_buffer_2841 (
        .din(new_Jinkela_wire_4155),
        .dout(new_Jinkela_wire_4156)
    );

    bfr new_Jinkela_buffer_4056 (
        .din(new_Jinkela_wire_5607),
        .dout(new_Jinkela_wire_5608)
    );

    bfr new_Jinkela_buffer_2782 (
        .din(new_Jinkela_wire_4094),
        .dout(new_Jinkela_wire_4095)
    );

    bfr new_Jinkela_buffer_4018 (
        .din(new_Jinkela_wire_5543),
        .dout(new_Jinkela_wire_5544)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_32),
        .dout(new_Jinkela_wire_33)
    );

    spl2 new_Jinkela_splitter_586 (
        .a(new_Jinkela_wire_5569),
        .b(new_Jinkela_wire_5570),
        .c(new_Jinkela_wire_5571)
    );

    bfr new_Jinkela_buffer_14 (
        .din(G110),
        .dout(new_Jinkela_wire_64)
    );

    bfr new_Jinkela_buffer_2805 (
        .din(new_Jinkela_wire_4119),
        .dout(new_Jinkela_wire_4120)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_36),
        .dout(new_Jinkela_wire_37)
    );

    bfr new_Jinkela_buffer_2783 (
        .din(new_Jinkela_wire_4095),
        .dout(new_Jinkela_wire_4096)
    );

    bfr new_Jinkela_buffer_4019 (
        .din(new_Jinkela_wire_5544),
        .dout(new_Jinkela_wire_5545)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_33),
        .dout(new_Jinkela_wire_34)
    );

    bfr new_Jinkela_buffer_4036 (
        .din(new_Jinkela_wire_5571),
        .dout(new_Jinkela_wire_5572)
    );

    bfr new_Jinkela_buffer_2817 (
        .din(new_Jinkela_wire_4131),
        .dout(new_Jinkela_wire_4132)
    );

    bfr new_Jinkela_buffer_2784 (
        .din(new_Jinkela_wire_4096),
        .dout(new_Jinkela_wire_4097)
    );

    spl4L new_Jinkela_splitter_583 (
        .a(new_Jinkela_wire_5545),
        .d(new_Jinkela_wire_5546),
        .e(new_Jinkela_wire_5547),
        .b(new_Jinkela_wire_5548),
        .c(new_Jinkela_wire_5549)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    spl4L new_Jinkela_splitter_9 (
        .a(new_Jinkela_wire_43),
        .d(new_Jinkela_wire_44),
        .e(new_Jinkela_wire_45),
        .b(new_Jinkela_wire_46),
        .c(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_2806 (
        .din(new_Jinkela_wire_4120),
        .dout(new_Jinkela_wire_4121)
    );

    bfr new_Jinkela_buffer_4057 (
        .din(new_Jinkela_wire_5608),
        .dout(new_Jinkela_wire_5609)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_37),
        .dout(new_Jinkela_wire_38)
    );

    bfr new_Jinkela_buffer_2785 (
        .din(new_Jinkela_wire_4097),
        .dout(new_Jinkela_wire_4098)
    );

    bfr new_Jinkela_buffer_4077 (
        .din(new_Jinkela_wire_5628),
        .dout(new_Jinkela_wire_5629)
    );

    bfr new_Jinkela_buffer_4037 (
        .din(new_Jinkela_wire_5572),
        .dout(new_Jinkela_wire_5573)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    spl2 new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_39),
        .c(new_Jinkela_wire_40)
    );

    bfr new_Jinkela_buffer_2786 (
        .din(new_Jinkela_wire_4098),
        .dout(new_Jinkela_wire_4099)
    );

    bfr new_Jinkela_buffer_4067 (
        .din(new_Jinkela_wire_5618),
        .dout(new_Jinkela_wire_5619)
    );

    bfr new_Jinkela_buffer_2852 (
        .din(new_Jinkela_wire_4169),
        .dout(new_Jinkela_wire_4170)
    );

    spl2 new_Jinkela_splitter_587 (
        .a(new_Jinkela_wire_5573),
        .b(new_Jinkela_wire_5574),
        .c(new_Jinkela_wire_5575)
    );

    bfr new_Jinkela_buffer_2807 (
        .din(new_Jinkela_wire_4121),
        .dout(new_Jinkela_wire_4122)
    );

    spl4L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_48),
        .d(new_Jinkela_wire_49),
        .e(new_Jinkela_wire_50),
        .b(new_Jinkela_wire_54),
        .c(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_2787 (
        .din(new_Jinkela_wire_4099),
        .dout(new_Jinkela_wire_4100)
    );

    bfr new_Jinkela_buffer_4038 (
        .din(new_Jinkela_wire_5575),
        .dout(new_Jinkela_wire_5576)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_41),
        .dout(new_Jinkela_wire_42)
    );

    spl3L new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_50),
        .d(new_Jinkela_wire_51),
        .b(new_Jinkela_wire_52),
        .c(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_2818 (
        .din(new_Jinkela_wire_4132),
        .dout(new_Jinkela_wire_4133)
    );

    bfr new_Jinkela_buffer_4058 (
        .din(new_Jinkela_wire_5609),
        .dout(new_Jinkela_wire_5610)
    );

    bfr new_Jinkela_buffer_2788 (
        .din(new_Jinkela_wire_4100),
        .dout(new_Jinkela_wire_4101)
    );

    bfr new_Jinkela_buffer_16 (
        .din(G53),
        .dout(new_Jinkela_wire_66)
    );

    spl2 new_Jinkela_splitter_597 (
        .a(_0935_),
        .b(new_Jinkela_wire_5654),
        .c(new_Jinkela_wire_5655)
    );

    bfr new_Jinkela_buffer_4039 (
        .din(new_Jinkela_wire_5576),
        .dout(new_Jinkela_wire_5577)
    );

    bfr new_Jinkela_buffer_21 (
        .din(G80),
        .dout(new_Jinkela_wire_71)
    );

    bfr new_Jinkela_buffer_2808 (
        .din(new_Jinkela_wire_4122),
        .dout(new_Jinkela_wire_4123)
    );

    spl3L new_Jinkela_splitter_15 (
        .a(G132),
        .d(new_Jinkela_wire_76),
        .b(new_Jinkela_wire_77),
        .c(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_2789 (
        .din(new_Jinkela_wire_4101),
        .dout(new_Jinkela_wire_4102)
    );

    bfr new_Jinkela_buffer_4079 (
        .din(new_Jinkela_wire_5631),
        .dout(new_Jinkela_wire_5632)
    );

    spl4L new_Jinkela_splitter_12 (
        .a(new_Jinkela_wire_54),
        .d(new_Jinkela_wire_55),
        .e(new_Jinkela_wire_56),
        .b(new_Jinkela_wire_57),
        .c(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_4059 (
        .din(new_Jinkela_wire_5610),
        .dout(new_Jinkela_wire_5611)
    );

    spl2 new_Jinkela_splitter_588 (
        .a(new_Jinkela_wire_5577),
        .b(new_Jinkela_wire_5578),
        .c(new_Jinkela_wire_5579)
    );

    spl4L new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_59),
        .d(new_Jinkela_wire_60),
        .e(new_Jinkela_wire_61),
        .b(new_Jinkela_wire_62),
        .c(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_2842 (
        .din(new_Jinkela_wire_4156),
        .dout(new_Jinkela_wire_4157)
    );

    bfr new_Jinkela_buffer_2790 (
        .din(new_Jinkela_wire_4102),
        .dout(new_Jinkela_wire_4103)
    );

    bfr new_Jinkela_buffer_4040 (
        .din(new_Jinkela_wire_5579),
        .dout(new_Jinkela_wire_5580)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_67),
        .dout(new_Jinkela_wire_68)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_66),
        .dout(new_Jinkela_wire_67)
    );

    bfr new_Jinkela_buffer_2809 (
        .din(new_Jinkela_wire_4123),
        .dout(new_Jinkela_wire_4124)
    );

    bfr new_Jinkela_buffer_4068 (
        .din(new_Jinkela_wire_5619),
        .dout(new_Jinkela_wire_5620)
    );

    bfr new_Jinkela_buffer_2791 (
        .din(new_Jinkela_wire_4103),
        .dout(new_Jinkela_wire_4104)
    );

    bfr new_Jinkela_buffer_4060 (
        .din(new_Jinkela_wire_5611),
        .dout(new_Jinkela_wire_5612)
    );

    spl2 new_Jinkela_splitter_589 (
        .a(new_Jinkela_wire_5580),
        .b(new_Jinkela_wire_5581),
        .c(new_Jinkela_wire_5582)
    );

    bfr new_Jinkela_buffer_26 (
        .din(G91),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_2819 (
        .din(new_Jinkela_wire_4133),
        .dout(new_Jinkela_wire_4134)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_71),
        .dout(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_2792 (
        .din(new_Jinkela_wire_4104),
        .dout(new_Jinkela_wire_4105)
    );

    bfr new_Jinkela_buffer_4041 (
        .din(new_Jinkela_wire_5582),
        .dout(new_Jinkela_wire_5583)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_28 (
        .din(G55),
        .dout(new_Jinkela_wire_83)
    );

    bfr new_Jinkela_buffer_2810 (
        .din(new_Jinkela_wire_4124),
        .dout(new_Jinkela_wire_4125)
    );

    bfr new_Jinkela_buffer_4078 (
        .din(new_Jinkela_wire_5629),
        .dout(new_Jinkela_wire_5630)
    );

    bfr new_Jinkela_buffer_2793 (
        .din(new_Jinkela_wire_4105),
        .dout(new_Jinkela_wire_4106)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_4061 (
        .din(new_Jinkela_wire_5612),
        .dout(new_Jinkela_wire_5613)
    );

    spl2 new_Jinkela_splitter_590 (
        .a(new_Jinkela_wire_5583),
        .b(new_Jinkela_wire_5584),
        .c(new_Jinkela_wire_5585)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    spl2 new_Jinkela_splitter_500 (
        .a(_0787_),
        .b(new_Jinkela_wire_4177),
        .c(new_Jinkela_wire_4178)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_2794 (
        .din(new_Jinkela_wire_4106),
        .dout(new_Jinkela_wire_4107)
    );

    bfr new_Jinkela_buffer_4042 (
        .din(new_Jinkela_wire_5585),
        .dout(new_Jinkela_wire_5586)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_2811 (
        .din(new_Jinkela_wire_4125),
        .dout(new_Jinkela_wire_4126)
    );

    bfr new_Jinkela_buffer_4069 (
        .din(new_Jinkela_wire_5620),
        .dout(new_Jinkela_wire_5621)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_73),
        .b(new_Jinkela_wire_74),
        .c(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_2795 (
        .din(new_Jinkela_wire_4107),
        .dout(new_Jinkela_wire_4108)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_79),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_4043 (
        .din(new_Jinkela_wire_5586),
        .dout(new_Jinkela_wire_5587)
    );

    bfr new_Jinkela_buffer_2820 (
        .din(new_Jinkela_wire_4134),
        .dout(new_Jinkela_wire_4135)
    );

    bfr new_Jinkela_buffer_2812 (
        .din(new_Jinkela_wire_4126),
        .dout(new_Jinkela_wire_4127)
    );

    bfr new_Jinkela_buffer_4070 (
        .din(new_Jinkela_wire_5621),
        .dout(new_Jinkela_wire_5622)
    );

    bfr new_Jinkela_buffer_4044 (
        .din(new_Jinkela_wire_5587),
        .dout(new_Jinkela_wire_5588)
    );

    spl2 new_Jinkela_splitter_16 (
        .a(G99),
        .b(new_Jinkela_wire_88),
        .c(new_Jinkela_wire_89)
    );

    bfr new_Jinkela_buffer_2843 (
        .din(new_Jinkela_wire_4157),
        .dout(new_Jinkela_wire_4158)
    );

    bfr new_Jinkela_buffer_33 (
        .din(G134),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_2813 (
        .din(new_Jinkela_wire_4127),
        .dout(new_Jinkela_wire_4128)
    );

    bfr new_Jinkela_buffer_4103 (
        .din(_0239_),
        .dout(new_Jinkela_wire_5663)
    );

    spl2 new_Jinkela_splitter_591 (
        .a(new_Jinkela_wire_5588),
        .b(new_Jinkela_wire_5589),
        .c(new_Jinkela_wire_5590)
    );

    bfr new_Jinkela_buffer_36 (
        .din(G61),
        .dout(new_Jinkela_wire_108)
    );

    bfr new_Jinkela_buffer_2821 (
        .din(new_Jinkela_wire_4135),
        .dout(new_Jinkela_wire_4136)
    );

    spl3L new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_91),
        .d(new_Jinkela_wire_92),
        .b(new_Jinkela_wire_94),
        .c(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_4045 (
        .din(new_Jinkela_wire_5590),
        .dout(new_Jinkela_wire_5591)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    spl4L new_Jinkela_splitter_596 (
        .a(new_Jinkela_wire_5633),
        .d(new_Jinkela_wire_5634),
        .e(new_Jinkela_wire_5635),
        .b(new_Jinkela_wire_5636),
        .c(new_Jinkela_wire_5637)
    );

    bfr new_Jinkela_buffer_2822 (
        .din(new_Jinkela_wire_4136),
        .dout(new_Jinkela_wire_4137)
    );

    bfr new_Jinkela_buffer_4071 (
        .din(new_Jinkela_wire_5622),
        .dout(new_Jinkela_wire_5623)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_2844 (
        .din(new_Jinkela_wire_4158),
        .dout(new_Jinkela_wire_4159)
    );

    bfr new_Jinkela_buffer_4080 (
        .din(new_Jinkela_wire_5637),
        .dout(new_Jinkela_wire_5638)
    );

    spl2 new_Jinkela_splitter_592 (
        .a(new_Jinkela_wire_5591),
        .b(new_Jinkela_wire_5592),
        .c(new_Jinkela_wire_5593)
    );

    bfr new_Jinkela_buffer_34 (
        .din(G121),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_2823 (
        .din(new_Jinkela_wire_4137),
        .dout(new_Jinkela_wire_4138)
    );

    spl2 new_Jinkela_splitter_593 (
        .a(new_Jinkela_wire_5593),
        .b(new_Jinkela_wire_5594),
        .c(new_Jinkela_wire_5595)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_2857 (
        .din(_0260_),
        .dout(new_Jinkela_wire_4179)
    );

    bfr new_Jinkela_buffer_2853 (
        .din(new_Jinkela_wire_4170),
        .dout(new_Jinkela_wire_4171)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_108),
        .dout(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_2824 (
        .din(new_Jinkela_wire_4138),
        .dout(new_Jinkela_wire_4139)
    );

    bfr new_Jinkela_buffer_4072 (
        .din(new_Jinkela_wire_5623),
        .dout(new_Jinkela_wire_5624)
    );

    bfr new_Jinkela_buffer_41 (
        .din(G37),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_4046 (
        .din(new_Jinkela_wire_5595),
        .dout(new_Jinkela_wire_5596)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(G165),
        .b(new_Jinkela_wire_116),
        .c(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_2845 (
        .din(new_Jinkela_wire_4159),
        .dout(new_Jinkela_wire_4160)
    );

    bfr new_Jinkela_buffer_2825 (
        .din(new_Jinkela_wire_4139),
        .dout(new_Jinkela_wire_4140)
    );

    bfr new_Jinkela_buffer_4095 (
        .din(new_Jinkela_wire_5652),
        .dout(new_Jinkela_wire_5653)
    );

    bfr new_Jinkela_buffer_4073 (
        .din(new_Jinkela_wire_5624),
        .dout(new_Jinkela_wire_5625)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1763),
        .dout(new_Jinkela_wire_1764)
    );

    spl2 new_Jinkela_splitter_313 (
        .a(new_Jinkela_wire_1724),
        .b(new_Jinkela_wire_1725),
        .c(new_Jinkela_wire_1726)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1726),
        .dout(new_Jinkela_wire_1727)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1791),
        .dout(new_Jinkela_wire_1792)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1764),
        .dout(new_Jinkela_wire_1765)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_1727),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1822),
        .dout(new_Jinkela_wire_1823)
    );

    spl2 new_Jinkela_splitter_314 (
        .a(new_Jinkela_wire_1728),
        .b(new_Jinkela_wire_1729),
        .c(new_Jinkela_wire_1730)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1730),
        .dout(new_Jinkela_wire_1731)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1765),
        .dout(new_Jinkela_wire_1766)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1792),
        .dout(new_Jinkela_wire_1793)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1731),
        .dout(new_Jinkela_wire_1732)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1766),
        .dout(new_Jinkela_wire_1767)
    );

    spl2 new_Jinkela_splitter_315 (
        .a(new_Jinkela_wire_1732),
        .b(new_Jinkela_wire_1733),
        .c(new_Jinkela_wire_1734)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1734),
        .dout(new_Jinkela_wire_1735)
    );

    spl2 new_Jinkela_splitter_325 (
        .a(_0718_),
        .b(new_Jinkela_wire_1858),
        .c(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1767),
        .dout(new_Jinkela_wire_1768)
    );

    spl2 new_Jinkela_splitter_316 (
        .a(new_Jinkela_wire_1735),
        .b(new_Jinkela_wire_1736),
        .c(new_Jinkela_wire_1737)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1737),
        .dout(new_Jinkela_wire_1738)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_1768),
        .dout(new_Jinkela_wire_1769)
    );

    spl2 new_Jinkela_splitter_317 (
        .a(new_Jinkela_wire_1738),
        .b(new_Jinkela_wire_1739),
        .c(new_Jinkela_wire_1740)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1740),
        .dout(new_Jinkela_wire_1741)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1823),
        .dout(new_Jinkela_wire_1824)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1769),
        .dout(new_Jinkela_wire_1770)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1741),
        .dout(new_Jinkela_wire_1742)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1794),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1742),
        .dout(new_Jinkela_wire_1743)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1770),
        .dout(new_Jinkela_wire_1771)
    );

    bfr new_Jinkela_buffer_872 (
        .din(new_Jinkela_wire_1743),
        .dout(new_Jinkela_wire_1744)
    );

    bfr new_Jinkela_buffer_969 (
        .din(_0800_),
        .dout(new_Jinkela_wire_1853)
    );

    spl2 new_Jinkela_splitter_318 (
        .a(new_Jinkela_wire_1744),
        .b(new_Jinkela_wire_1745),
        .c(new_Jinkela_wire_1746)
    );

    spl2 new_Jinkela_splitter_319 (
        .a(new_Jinkela_wire_1746),
        .b(new_Jinkela_wire_1747),
        .c(new_Jinkela_wire_1748)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1771),
        .dout(new_Jinkela_wire_1772)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_1748),
        .dout(new_Jinkela_wire_1749)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1795),
        .dout(new_Jinkela_wire_1796)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1772),
        .dout(new_Jinkela_wire_1773)
    );

    spl2 new_Jinkela_splitter_320 (
        .a(new_Jinkela_wire_1749),
        .b(new_Jinkela_wire_1750),
        .c(new_Jinkela_wire_1751)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1773),
        .dout(new_Jinkela_wire_1774)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1824),
        .dout(new_Jinkela_wire_1825)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1796),
        .dout(new_Jinkela_wire_1797)
    );

    bfr new_Jinkela_buffer_5042 (
        .din(new_Jinkela_wire_6873),
        .dout(new_Jinkela_wire_6874)
    );

    bfr new_Jinkela_buffer_5087 (
        .din(new_Jinkela_wire_6938),
        .dout(new_Jinkela_wire_6939)
    );

    bfr new_Jinkela_buffer_5069 (
        .din(new_Jinkela_wire_6914),
        .dout(new_Jinkela_wire_6915)
    );

    bfr new_Jinkela_buffer_5043 (
        .din(new_Jinkela_wire_6874),
        .dout(new_Jinkela_wire_6875)
    );

    bfr new_Jinkela_buffer_5044 (
        .din(new_Jinkela_wire_6875),
        .dout(new_Jinkela_wire_6876)
    );

    bfr new_Jinkela_buffer_5078 (
        .din(new_Jinkela_wire_6925),
        .dout(new_Jinkela_wire_6926)
    );

    bfr new_Jinkela_buffer_5070 (
        .din(new_Jinkela_wire_6915),
        .dout(new_Jinkela_wire_6916)
    );

    bfr new_Jinkela_buffer_5045 (
        .din(new_Jinkela_wire_6876),
        .dout(new_Jinkela_wire_6877)
    );

    bfr new_Jinkela_buffer_5046 (
        .din(new_Jinkela_wire_6877),
        .dout(new_Jinkela_wire_6878)
    );

    spl2 new_Jinkela_splitter_713 (
        .a(_0675_),
        .b(new_Jinkela_wire_6951),
        .c(new_Jinkela_wire_6952)
    );

    bfr new_Jinkela_buffer_5071 (
        .din(new_Jinkela_wire_6916),
        .dout(new_Jinkela_wire_6917)
    );

    bfr new_Jinkela_buffer_5047 (
        .din(new_Jinkela_wire_6878),
        .dout(new_Jinkela_wire_6879)
    );

    bfr new_Jinkela_buffer_5048 (
        .din(new_Jinkela_wire_6879),
        .dout(new_Jinkela_wire_6880)
    );

    bfr new_Jinkela_buffer_5079 (
        .din(new_Jinkela_wire_6926),
        .dout(new_Jinkela_wire_6927)
    );

    bfr new_Jinkela_buffer_5072 (
        .din(new_Jinkela_wire_6917),
        .dout(new_Jinkela_wire_6918)
    );

    bfr new_Jinkela_buffer_5049 (
        .din(new_Jinkela_wire_6880),
        .dout(new_Jinkela_wire_6881)
    );

    bfr new_Jinkela_buffer_5050 (
        .din(new_Jinkela_wire_6881),
        .dout(new_Jinkela_wire_6882)
    );

    bfr new_Jinkela_buffer_5073 (
        .din(new_Jinkela_wire_6918),
        .dout(new_Jinkela_wire_6919)
    );

    bfr new_Jinkela_buffer_5051 (
        .din(new_Jinkela_wire_6882),
        .dout(new_Jinkela_wire_6883)
    );

    bfr new_Jinkela_buffer_5052 (
        .din(new_Jinkela_wire_6883),
        .dout(new_Jinkela_wire_6884)
    );

    bfr new_Jinkela_buffer_5080 (
        .din(new_Jinkela_wire_6927),
        .dout(new_Jinkela_wire_6928)
    );

    bfr new_Jinkela_buffer_5074 (
        .din(new_Jinkela_wire_6919),
        .dout(new_Jinkela_wire_6920)
    );

    bfr new_Jinkela_buffer_5053 (
        .din(new_Jinkela_wire_6884),
        .dout(new_Jinkela_wire_6885)
    );

    bfr new_Jinkela_buffer_5054 (
        .din(new_Jinkela_wire_6885),
        .dout(new_Jinkela_wire_6886)
    );

    bfr new_Jinkela_buffer_5088 (
        .din(new_Jinkela_wire_6939),
        .dout(new_Jinkela_wire_6940)
    );

    bfr new_Jinkela_buffer_5055 (
        .din(new_Jinkela_wire_6886),
        .dout(new_Jinkela_wire_6887)
    );

    bfr new_Jinkela_buffer_5081 (
        .din(new_Jinkela_wire_6928),
        .dout(new_Jinkela_wire_6929)
    );

    bfr new_Jinkela_buffer_5100 (
        .din(_0483_),
        .dout(new_Jinkela_wire_6956)
    );

    bfr new_Jinkela_buffer_5097 (
        .din(new_Jinkela_wire_6952),
        .dout(new_Jinkela_wire_6953)
    );

    bfr new_Jinkela_buffer_5082 (
        .din(new_Jinkela_wire_6929),
        .dout(new_Jinkela_wire_6930)
    );

    bfr new_Jinkela_buffer_5089 (
        .din(new_Jinkela_wire_6940),
        .dout(new_Jinkela_wire_6941)
    );

    bfr new_Jinkela_buffer_5083 (
        .din(new_Jinkela_wire_6930),
        .dout(new_Jinkela_wire_6931)
    );

    spl2 new_Jinkela_splitter_714 (
        .a(_1092_),
        .b(new_Jinkela_wire_6987),
        .c(new_Jinkela_wire_6988)
    );

    bfr new_Jinkela_buffer_5084 (
        .din(new_Jinkela_wire_6931),
        .dout(new_Jinkela_wire_6932)
    );

    bfr new_Jinkela_buffer_5090 (
        .din(new_Jinkela_wire_6941),
        .dout(new_Jinkela_wire_6942)
    );

    bfr new_Jinkela_buffer_5085 (
        .din(new_Jinkela_wire_6932),
        .dout(new_Jinkela_wire_6933)
    );

    spl2 new_Jinkela_splitter_715 (
        .a(new_net_23),
        .b(new_Jinkela_wire_6989),
        .c(new_Jinkela_wire_6991)
    );

    bfr new_Jinkela_buffer_5101 (
        .din(new_Jinkela_wire_6956),
        .dout(new_Jinkela_wire_6957)
    );

    bfr new_Jinkela_buffer_5091 (
        .din(new_Jinkela_wire_6942),
        .dout(new_Jinkela_wire_6943)
    );

    bfr new_Jinkela_buffer_5098 (
        .din(new_Jinkela_wire_6953),
        .dout(new_Jinkela_wire_6954)
    );

    bfr new_Jinkela_buffer_5092 (
        .din(new_Jinkela_wire_6943),
        .dout(new_Jinkela_wire_6944)
    );

    bfr new_Jinkela_buffer_5093 (
        .din(new_Jinkela_wire_6944),
        .dout(new_Jinkela_wire_6945)
    );

    spl4L new_Jinkela_splitter_18 (
        .a(new_Jinkela_wire_94),
        .d(new_Jinkela_wire_95),
        .e(new_Jinkela_wire_96),
        .b(new_Jinkela_wire_97),
        .c(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    spl4L new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_99),
        .d(new_Jinkela_wire_100),
        .e(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_102),
        .c(new_Jinkela_wire_103)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_103),
        .b(new_Jinkela_wire_104),
        .c(new_Jinkela_wire_105)
    );

    bfr new_Jinkela_buffer_42 (
        .din(G39),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_109),
        .dout(new_Jinkela_wire_110)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(new_Jinkela_wire_105),
        .b(new_Jinkela_wire_106),
        .c(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_67 (
        .din(G5),
        .dout(new_Jinkela_wire_147)
    );

    spl2 new_Jinkela_splitter_25 (
        .a(G157),
        .b(new_Jinkela_wire_123),
        .c(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    spl2 new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_112),
        .b(new_Jinkela_wire_113),
        .c(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_70 (
        .din(G105),
        .dout(new_Jinkela_wire_152)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(new_Jinkela_wire_120),
        .b(new_Jinkela_wire_121),
        .c(new_Jinkela_wire_122)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_147),
        .dout(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    spl3L new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_167),
        .d(new_Jinkela_wire_168),
        .b(new_Jinkela_wire_169),
        .c(new_Jinkela_wire_170)
    );

    spl2 new_Jinkela_splitter_31 (
        .a(G117),
        .b(new_Jinkela_wire_167),
        .c(new_Jinkela_wire_171)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    spl4L new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_157),
        .d(new_Jinkela_wire_158),
        .e(new_Jinkela_wire_159),
        .b(new_Jinkela_wire_160),
        .c(new_Jinkela_wire_161)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    spl2 new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_149),
        .b(new_Jinkela_wire_150),
        .c(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    spl4L new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_152),
        .d(new_Jinkela_wire_153),
        .e(new_Jinkela_wire_154),
        .b(new_Jinkela_wire_157),
        .c(new_Jinkela_wire_162)
    );

    spl4L new_Jinkela_splitter_33 (
        .a(new_Jinkela_wire_171),
        .d(new_Jinkela_wire_172),
        .e(new_Jinkela_wire_173),
        .b(new_Jinkela_wire_174),
        .c(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    spl2 new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_154),
        .b(new_Jinkela_wire_155),
        .c(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_72 (
        .din(G16),
        .dout(new_Jinkela_wire_177)
    );

    spl4L new_Jinkela_splitter_30 (
        .a(new_Jinkela_wire_162),
        .d(new_Jinkela_wire_163),
        .e(new_Jinkela_wire_164),
        .b(new_Jinkela_wire_165),
        .c(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    bfr new_Jinkela_buffer_80 (
        .din(G18),
        .dout(new_Jinkela_wire_187)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_136),
        .dout(new_Jinkela_wire_137)
    );

    bfr new_Jinkela_buffer_75 (
        .din(G44),
        .dout(new_Jinkela_wire_182)
    );

    or_bb _2540_ (
        .a(new_Jinkela_wire_5948),
        .b(_0522_),
        .c(_0525_)
    );

    or_bb _1823_ (
        .a(new_Jinkela_wire_7882),
        .b(new_Jinkela_wire_2121),
        .c(_1112_)
    );

    bfr new_Jinkela_buffer_2752 (
        .din(new_Jinkela_wire_4060),
        .dout(new_Jinkela_wire_4061)
    );

    and_bi _2541_ (
        .a(new_Jinkela_wire_335),
        .b(new_Jinkela_wire_7926),
        .c(_0526_)
    );

    and_bi _1824_ (
        .a(new_Jinkela_wire_3169),
        .b(new_Jinkela_wire_1684),
        .c(_1113_)
    );

    bfr new_Jinkela_buffer_2730 (
        .din(new_Jinkela_wire_4019),
        .dout(new_Jinkela_wire_4020)
    );

    and_bi _2542_ (
        .a(new_Jinkela_wire_865),
        .b(new_Jinkela_wire_6129),
        .c(_0527_)
    );

    or_bb _1825_ (
        .a(_1113_),
        .b(new_Jinkela_wire_6281),
        .c(_1114_)
    );

    bfr new_Jinkela_buffer_2746 (
        .din(new_Jinkela_wire_4048),
        .dout(new_Jinkela_wire_4049)
    );

    or_bb _2543_ (
        .a(_0527_),
        .b(_0526_),
        .c(_0528_)
    );

    and_bi _1826_ (
        .a(_1112_),
        .b(_1114_),
        .c(_1115_)
    );

    and_bi _2544_ (
        .a(_0525_),
        .b(new_Jinkela_wire_2569),
        .c(_0529_)
    );

    or_bb _1827_ (
        .a(_1115_),
        .b(_1110_),
        .c(_1116_)
    );

    bfr new_Jinkela_buffer_2753 (
        .din(new_Jinkela_wire_4061),
        .dout(new_Jinkela_wire_4062)
    );

    and_bi _2545_ (
        .a(new_Jinkela_wire_693),
        .b(_0529_),
        .c(new_net_2449)
    );

    and_bb _1828_ (
        .a(new_Jinkela_wire_3252),
        .b(new_Jinkela_wire_5789),
        .c(_1117_)
    );

    bfr new_Jinkela_buffer_2814 (
        .din(_1008_),
        .dout(new_Jinkela_wire_4129)
    );

    and_bi _2546_ (
        .a(new_Jinkela_wire_6992),
        .b(new_Jinkela_wire_816),
        .c(_0530_)
    );

    bfr new_Jinkela_buffer_2769 (
        .din(new_Jinkela_wire_4081),
        .dout(new_Jinkela_wire_4082)
    );

    and_bi _1829_ (
        .a(new_Jinkela_wire_6096),
        .b(new_Jinkela_wire_2312),
        .c(_1118_)
    );

    bfr new_Jinkela_buffer_2754 (
        .din(new_Jinkela_wire_4062),
        .dout(new_Jinkela_wire_4063)
    );

    and_bi _2547_ (
        .a(new_Jinkela_wire_6904),
        .b(new_Jinkela_wire_6838),
        .c(_0531_)
    );

    or_bb _1830_ (
        .a(new_Jinkela_wire_2331),
        .b(new_Jinkela_wire_3094),
        .c(_1119_)
    );

    or_bb _2548_ (
        .a(_0531_),
        .b(new_Jinkela_wire_5589),
        .c(_0532_)
    );

    bfr new_Jinkela_buffer_2797 (
        .din(new_Jinkela_wire_4109),
        .dout(new_Jinkela_wire_4110)
    );

    and_bb _1831_ (
        .a(new_Jinkela_wire_2332),
        .b(new_Jinkela_wire_3095),
        .c(_1120_)
    );

    bfr new_Jinkela_buffer_2755 (
        .din(new_Jinkela_wire_4063),
        .dout(new_Jinkela_wire_4064)
    );

    or_bb _2549_ (
        .a(_0532_),
        .b(_0530_),
        .c(_0533_)
    );

    and_bi _1832_ (
        .a(_1119_),
        .b(_1120_),
        .c(_1121_)
    );

    and_bi _2550_ (
        .a(new_Jinkela_wire_1344),
        .b(new_Jinkela_wire_3386),
        .c(_0534_)
    );

    bfr new_Jinkela_buffer_2770 (
        .din(new_Jinkela_wire_4082),
        .dout(new_Jinkela_wire_4083)
    );

    and_ii _1833_ (
        .a(new_Jinkela_wire_5121),
        .b(new_Jinkela_wire_7933),
        .c(_1122_)
    );

    bfr new_Jinkela_buffer_2756 (
        .din(new_Jinkela_wire_4064),
        .dout(new_Jinkela_wire_4065)
    );

    and_bi _2551_ (
        .a(new_Jinkela_wire_331),
        .b(new_Jinkela_wire_4032),
        .c(_0535_)
    );

    and_bb _1834_ (
        .a(new_Jinkela_wire_5122),
        .b(new_Jinkela_wire_7934),
        .c(_1123_)
    );

    or_bb _2552_ (
        .a(_0535_),
        .b(_0534_),
        .c(_0536_)
    );

    or_bb _1835_ (
        .a(_1123_),
        .b(new_Jinkela_wire_1100),
        .c(_1124_)
    );

    bfr new_Jinkela_buffer_2757 (
        .din(new_Jinkela_wire_4065),
        .dout(new_Jinkela_wire_4066)
    );

    and_bi _2553_ (
        .a(_0533_),
        .b(new_Jinkela_wire_4795),
        .c(_0537_)
    );

    or_bb _1836_ (
        .a(_1124_),
        .b(new_Jinkela_wire_1974),
        .c(_1125_)
    );

    bfr new_Jinkela_buffer_2800 (
        .din(new_Jinkela_wire_4114),
        .dout(new_Jinkela_wire_4115)
    );

    and_bi _2554_ (
        .a(new_Jinkela_wire_687),
        .b(_0537_),
        .c(new_net_2491)
    );

    bfr new_Jinkela_buffer_2771 (
        .din(new_Jinkela_wire_4083),
        .dout(new_Jinkela_wire_4084)
    );

    or_bb _1837_ (
        .a(new_Jinkela_wire_1332),
        .b(new_Jinkela_wire_57),
        .c(_1126_)
    );

    bfr new_Jinkela_buffer_2758 (
        .din(new_Jinkela_wire_4066),
        .dout(new_Jinkela_wire_4067)
    );

    and_bi _2555_ (
        .a(new_Jinkela_wire_5361),
        .b(new_Jinkela_wire_824),
        .c(_0538_)
    );

    and_bi _1838_ (
        .a(new_Jinkela_wire_1329),
        .b(new_Jinkela_wire_409),
        .c(_1127_)
    );

    and_bi _2556_ (
        .a(new_Jinkela_wire_820),
        .b(new_Jinkela_wire_1613),
        .c(_0539_)
    );

    bfr new_Jinkela_buffer_2798 (
        .din(new_Jinkela_wire_4110),
        .dout(new_Jinkela_wire_4111)
    );

    and_bi _1839_ (
        .a(_1126_),
        .b(_1127_),
        .c(_1128_)
    );

    bfr new_Jinkela_buffer_2759 (
        .din(new_Jinkela_wire_4067),
        .dout(new_Jinkela_wire_4068)
    );

    or_bb _2557_ (
        .a(_0539_),
        .b(new_Jinkela_wire_5594),
        .c(_0540_)
    );

    and_bi _1840_ (
        .a(new_Jinkela_wire_1304),
        .b(_1128_),
        .c(_1129_)
    );

    or_bb _2558_ (
        .a(_0540_),
        .b(_0538_),
        .c(_0541_)
    );

    bfr new_Jinkela_buffer_2772 (
        .din(new_Jinkela_wire_4084),
        .dout(new_Jinkela_wire_4085)
    );

    or_ii _1841_ (
        .a(new_Jinkela_wire_1338),
        .b(new_Jinkela_wire_1212),
        .c(_1130_)
    );

    bfr new_Jinkela_buffer_2760 (
        .din(new_Jinkela_wire_4068),
        .dout(new_Jinkela_wire_4069)
    );

    and_bi _2559_ (
        .a(new_Jinkela_wire_962),
        .b(new_Jinkela_wire_4033),
        .c(_0542_)
    );

    and_bi _1842_ (
        .a(new_Jinkela_wire_1536),
        .b(new_Jinkela_wire_1327),
        .c(_1131_)
    );

    and_bi _2560_ (
        .a(new_Jinkela_wire_1576),
        .b(new_Jinkela_wire_3389),
        .c(_0543_)
    );

    and_bi _1843_ (
        .a(_1130_),
        .b(_1131_),
        .c(_1132_)
    );

    bfr new_Jinkela_buffer_2761 (
        .din(new_Jinkela_wire_4069),
        .dout(new_Jinkela_wire_4070)
    );

    or_bb _2561_ (
        .a(_0543_),
        .b(_0542_),
        .c(_0544_)
    );

    and_bi _1844_ (
        .a(new_Jinkela_wire_2858),
        .b(_1132_),
        .c(_1133_)
    );

    bfr new_Jinkela_buffer_2840 (
        .din(new_net_2501),
        .dout(new_Jinkela_wire_4155)
    );

    and_bi _2562_ (
        .a(_0541_),
        .b(new_Jinkela_wire_3746),
        .c(_0545_)
    );

    bfr new_Jinkela_buffer_2773 (
        .din(new_Jinkela_wire_4085),
        .dout(new_Jinkela_wire_4086)
    );

    and_ii _1845_ (
        .a(_1133_),
        .b(_1129_),
        .c(_1134_)
    );

    bfr new_Jinkela_buffer_2762 (
        .din(new_Jinkela_wire_4070),
        .dout(new_Jinkela_wire_4071)
    );

    and_bi _2563_ (
        .a(new_Jinkela_wire_692),
        .b(_0545_),
        .c(new_net_2493)
    );

    or_bb _1846_ (
        .a(new_Jinkela_wire_565),
        .b(new_Jinkela_wire_61),
        .c(_1135_)
    );

    and_bi _2564_ (
        .a(new_Jinkela_wire_5776),
        .b(new_Jinkela_wire_6842),
        .c(_0546_)
    );

    spl2 new_Jinkela_splitter_497 (
        .a(new_Jinkela_wire_4111),
        .b(new_Jinkela_wire_4112),
        .c(new_Jinkela_wire_4113)
    );

    and_bi _1847_ (
        .a(new_Jinkela_wire_557),
        .b(new_Jinkela_wire_418),
        .c(_1136_)
    );

    bfr new_Jinkela_buffer_2763 (
        .din(new_Jinkela_wire_4071),
        .dout(new_Jinkela_wire_4072)
    );

    and_bi _2565_ (
        .a(new_Jinkela_wire_6795),
        .b(new_Jinkela_wire_822),
        .c(_0547_)
    );

    and_bi _1848_ (
        .a(_1135_),
        .b(_1136_),
        .c(_1137_)
    );

    or_bb _2566_ (
        .a(_0547_),
        .b(new_Jinkela_wire_5596),
        .c(_0548_)
    );

    bfr new_Jinkela_buffer_2774 (
        .din(new_Jinkela_wire_4086),
        .dout(new_Jinkela_wire_4087)
    );

    and_bi _1849_ (
        .a(new_Jinkela_wire_1142),
        .b(_1137_),
        .c(_1138_)
    );

    bfr new_Jinkela_buffer_2764 (
        .din(new_Jinkela_wire_4072),
        .dout(new_Jinkela_wire_4073)
    );

    or_bb _2567_ (
        .a(_0548_),
        .b(new_Jinkela_wire_5867),
        .c(_0549_)
    );

    or_ii _1850_ (
        .a(new_Jinkela_wire_561),
        .b(new_Jinkela_wire_1208),
        .c(_1139_)
    );

    and_bi _2568_ (
        .a(new_Jinkela_wire_1360),
        .b(new_Jinkela_wire_3388),
        .c(_0550_)
    );

    and_bi _1851_ (
        .a(new_Jinkela_wire_1546),
        .b(new_Jinkela_wire_566),
        .c(_1140_)
    );

    bfr new_Jinkela_buffer_2815 (
        .din(new_Jinkela_wire_4129),
        .dout(new_Jinkela_wire_4130)
    );

    and_bi _2569_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_4023),
        .c(_0551_)
    );

    bfr new_Jinkela_buffer_2775 (
        .din(new_Jinkela_wire_4087),
        .dout(new_Jinkela_wire_4088)
    );

    and_bi _1852_ (
        .a(_1139_),
        .b(_1140_),
        .c(_1141_)
    );

    or_bb _2570_ (
        .a(_0551_),
        .b(_0550_),
        .c(_0552_)
    );

    and_bi _1853_ (
        .a(new_Jinkela_wire_3574),
        .b(_1141_),
        .c(_1142_)
    );

    bfr new_Jinkela_buffer_2801 (
        .din(new_Jinkela_wire_4115),
        .dout(new_Jinkela_wire_4116)
    );

    and_bi _2571_ (
        .a(_0549_),
        .b(new_Jinkela_wire_7183),
        .c(_0553_)
    );

    bfr new_Jinkela_buffer_2776 (
        .din(new_Jinkela_wire_4088),
        .dout(new_Jinkela_wire_4089)
    );

    and_ii _1854_ (
        .a(_1142_),
        .b(_1138_),
        .c(_1143_)
    );

    and_bi _2572_ (
        .a(new_Jinkela_wire_697),
        .b(_0553_),
        .c(new_net_2363)
    );

    and_bi _1855_ (
        .a(new_Jinkela_wire_6549),
        .b(new_Jinkela_wire_7522),
        .c(_1144_)
    );

    bfr new_Jinkela_buffer_2802 (
        .din(new_Jinkela_wire_4116),
        .dout(new_Jinkela_wire_4117)
    );

    and_bi _2573_ (
        .a(new_Jinkela_wire_3614),
        .b(new_Jinkela_wire_823),
        .c(_0554_)
    );

    bfr new_Jinkela_buffer_2777 (
        .din(new_Jinkela_wire_4089),
        .dout(new_Jinkela_wire_4090)
    );

    and_bi _1856_ (
        .a(new_Jinkela_wire_7523),
        .b(new_Jinkela_wire_6550),
        .c(_1145_)
    );

    and_bi _2574_ (
        .a(new_Jinkela_wire_5003),
        .b(new_Jinkela_wire_6819),
        .c(_0555_)
    );

    and_ii _1857_ (
        .a(_1145_),
        .b(_1144_),
        .c(_1146_)
    );

    spl3L new_Jinkela_splitter_498 (
        .a(_0659_),
        .d(new_Jinkela_wire_4167),
        .b(new_Jinkela_wire_4168),
        .c(new_Jinkela_wire_4169)
    );

    or_bb _2575_ (
        .a(_0555_),
        .b(new_Jinkela_wire_5570),
        .c(_0556_)
    );

    bfr new_Jinkela_buffer_2778 (
        .din(new_Jinkela_wire_4090),
        .dout(new_Jinkela_wire_4091)
    );

    or_bb _1858_ (
        .a(new_Jinkela_wire_846),
        .b(new_Jinkela_wire_46),
        .c(_1147_)
    );

    or_bb _2576_ (
        .a(new_Jinkela_wire_5047),
        .b(_0554_),
        .c(_0557_)
    );

    bfr new_Jinkela_buffer_2854 (
        .din(_1191_),
        .dout(new_Jinkela_wire_4172)
    );

    and_bi _1859_ (
        .a(new_Jinkela_wire_856),
        .b(new_Jinkela_wire_406),
        .c(_1148_)
    );

    bfr new_Jinkela_buffer_2803 (
        .din(new_Jinkela_wire_4117),
        .dout(new_Jinkela_wire_4118)
    );

    and_bi _2577_ (
        .a(new_Jinkela_wire_336),
        .b(new_Jinkela_wire_3379),
        .c(_0558_)
    );

    bfr new_Jinkela_buffer_2779 (
        .din(new_Jinkela_wire_4091),
        .dout(new_Jinkela_wire_4092)
    );

    and_bi _1860_ (
        .a(_1147_),
        .b(_1148_),
        .c(_1149_)
    );

    and_bi _2578_ (
        .a(new_Jinkela_wire_866),
        .b(new_Jinkela_wire_4022),
        .c(_0559_)
    );

    and_bi _1861_ (
        .a(new_Jinkela_wire_535),
        .b(_1149_),
        .c(_1150_)
    );

    bfr new_Jinkela_buffer_2816 (
        .din(new_Jinkela_wire_4130),
        .dout(new_Jinkela_wire_4131)
    );

    or_bb _2579_ (
        .a(_0559_),
        .b(_0558_),
        .c(_0560_)
    );

    bfr new_Jinkela_buffer_2780 (
        .din(new_Jinkela_wire_4092),
        .dout(new_Jinkela_wire_4093)
    );

    or_ii _1862_ (
        .a(new_Jinkela_wire_857),
        .b(new_Jinkela_wire_1197),
        .c(_1151_)
    );

    and_bi _2580_ (
        .a(_0557_),
        .b(new_Jinkela_wire_3661),
        .c(_0561_)
    );

    and_bi _1863_ (
        .a(new_Jinkela_wire_1530),
        .b(new_Jinkela_wire_853),
        .c(_1152_)
    );

    bfr new_Jinkela_buffer_2804 (
        .din(new_Jinkela_wire_4118),
        .dout(new_Jinkela_wire_4119)
    );

    and_bi _2581_ (
        .a(new_Jinkela_wire_694),
        .b(_0561_),
        .c(new_net_2391)
    );

    bfr new_Jinkela_buffer_2781 (
        .din(new_Jinkela_wire_4093),
        .dout(new_Jinkela_wire_4094)
    );

    and_bi _1864_ (
        .a(_1151_),
        .b(_1152_),
        .c(_1153_)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_137),
        .dout(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_2545),
        .dout(new_Jinkela_wire_2546)
    );

    bfr new_Jinkela_buffer_83 (
        .din(G96),
        .dout(new_Jinkela_wire_192)
    );

    bfr new_Jinkela_buffer_5028 (
        .din(new_Jinkela_wire_6859),
        .dout(new_Jinkela_wire_6860)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_2498),
        .dout(new_Jinkela_wire_2499)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    bfr new_Jinkela_buffer_5063 (
        .din(new_Jinkela_wire_6903),
        .dout(new_Jinkela_wire_6904)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_2519),
        .dout(new_Jinkela_wire_2520)
    );

    spl2 new_Jinkela_splitter_698 (
        .a(new_Jinkela_wire_6829),
        .b(new_Jinkela_wire_6830),
        .c(new_Jinkela_wire_6831)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(new_Jinkela_wire_2499),
        .dout(new_Jinkela_wire_2500)
    );

    bfr new_Jinkela_buffer_5008 (
        .din(new_Jinkela_wire_6831),
        .dout(new_Jinkela_wire_6832)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_5062 (
        .din(new_Jinkela_wire_6897),
        .dout(new_Jinkela_wire_6898)
    );

    bfr new_Jinkela_buffer_5029 (
        .din(new_Jinkela_wire_6860),
        .dout(new_Jinkela_wire_6861)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(new_Jinkela_wire_2520),
        .dout(new_Jinkela_wire_2521)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(new_Jinkela_wire_2546),
        .dout(new_Jinkela_wire_2547)
    );

    spl2 new_Jinkela_splitter_699 (
        .a(new_Jinkela_wire_6832),
        .b(new_Jinkela_wire_6833),
        .c(new_Jinkela_wire_6834)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_178),
        .dout(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_2521),
        .dout(new_Jinkela_wire_2522)
    );

    bfr new_Jinkela_buffer_5009 (
        .din(new_Jinkela_wire_6834),
        .dout(new_Jinkela_wire_6835)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(new_Jinkela_wire_2583),
        .dout(new_Jinkela_wire_2584)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_2574),
        .dout(new_Jinkela_wire_2575)
    );

    bfr new_Jinkela_buffer_5030 (
        .din(new_Jinkela_wire_6861),
        .dout(new_Jinkela_wire_6862)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_2522),
        .dout(new_Jinkela_wire_2523)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_142),
        .dout(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(new_Jinkela_wire_2547),
        .dout(new_Jinkela_wire_2548)
    );

    bfr new_Jinkela_buffer_5010 (
        .din(new_Jinkela_wire_6835),
        .dout(new_Jinkela_wire_6836)
    );

    spl2 new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_180),
        .c(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_2523),
        .dout(new_Jinkela_wire_2524)
    );

    bfr new_Jinkela_buffer_5075 (
        .din(new_Jinkela_wire_6922),
        .dout(new_Jinkela_wire_6923)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    bfr new_Jinkela_buffer_5031 (
        .din(new_Jinkela_wire_6862),
        .dout(new_Jinkela_wire_6863)
    );

    bfr new_Jinkela_buffer_5011 (
        .din(new_Jinkela_wire_6836),
        .dout(new_Jinkela_wire_6837)
    );

    spl2 new_Jinkela_splitter_40 (
        .a(G168),
        .b(new_Jinkela_wire_207),
        .c(new_Jinkela_wire_209)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_2524),
        .dout(new_Jinkela_wire_2525)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    spl4L new_Jinkela_splitter_708 (
        .a(new_Jinkela_wire_6905),
        .d(new_Jinkela_wire_6906),
        .e(new_Jinkela_wire_6907),
        .b(new_Jinkela_wire_6908),
        .c(new_Jinkela_wire_6909)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(new_Jinkela_wire_2548),
        .dout(new_Jinkela_wire_2549)
    );

    spl2 new_Jinkela_splitter_700 (
        .a(new_Jinkela_wire_6837),
        .b(new_Jinkela_wire_6838),
        .c(new_Jinkela_wire_6839)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_2525),
        .dout(new_Jinkela_wire_2526)
    );

    bfr new_Jinkela_buffer_5012 (
        .din(new_Jinkela_wire_6839),
        .dout(new_Jinkela_wire_6840)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_145),
        .dout(new_Jinkela_wire_146)
    );

    bfr new_Jinkela_buffer_1613 (
        .din(new_Jinkela_wire_2624),
        .dout(new_Jinkela_wire_2625)
    );

    bfr new_Jinkela_buffer_5064 (
        .din(new_Jinkela_wire_6909),
        .dout(new_Jinkela_wire_6910)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(new_Jinkela_wire_2575),
        .dout(new_Jinkela_wire_2576)
    );

    bfr new_Jinkela_buffer_5032 (
        .din(new_Jinkela_wire_6863),
        .dout(new_Jinkela_wire_6864)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_2526),
        .dout(new_Jinkela_wire_2527)
    );

    spl4L new_Jinkela_splitter_36 (
        .a(new_Jinkela_wire_192),
        .d(new_Jinkela_wire_193),
        .e(new_Jinkela_wire_194),
        .b(new_Jinkela_wire_197),
        .c(new_Jinkela_wire_202)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(new_Jinkela_wire_2549),
        .dout(new_Jinkela_wire_2550)
    );

    bfr new_Jinkela_buffer_5013 (
        .din(new_Jinkela_wire_6840),
        .dout(new_Jinkela_wire_6841)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_2527),
        .dout(new_Jinkela_wire_2528)
    );

    bfr new_Jinkela_buffer_5033 (
        .din(new_Jinkela_wire_6864),
        .dout(new_Jinkela_wire_6865)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_207),
        .dout(new_Jinkela_wire_208)
    );

    spl2 new_Jinkela_splitter_701 (
        .a(new_Jinkela_wire_6841),
        .b(new_Jinkela_wire_6842),
        .c(new_Jinkela_wire_6843)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(new_Jinkela_wire_2528),
        .dout(new_Jinkela_wire_2529)
    );

    bfr new_Jinkela_buffer_5014 (
        .din(new_Jinkela_wire_6843),
        .dout(new_Jinkela_wire_6844)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_2550),
        .dout(new_Jinkela_wire_2551)
    );

    spl2 new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_189),
        .b(new_Jinkela_wire_190),
        .c(new_Jinkela_wire_191)
    );

    spl2 new_Jinkela_splitter_711 (
        .a(_0970_),
        .b(new_Jinkela_wire_6937),
        .c(new_Jinkela_wire_6938)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(new_Jinkela_wire_2529),
        .dout(new_Jinkela_wire_2530)
    );

    bfr new_Jinkela_buffer_5086 (
        .din(new_Jinkela_wire_6935),
        .dout(new_Jinkela_wire_6936)
    );

    spl4L new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_209),
        .d(new_Jinkela_wire_210),
        .e(new_Jinkela_wire_211),
        .b(new_Jinkela_wire_213),
        .c(new_Jinkela_wire_218)
    );

    bfr new_Jinkela_buffer_5034 (
        .din(new_Jinkela_wire_6865),
        .dout(new_Jinkela_wire_6866)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(new_Jinkela_wire_2584),
        .dout(new_Jinkela_wire_2585)
    );

    bfr new_Jinkela_buffer_5015 (
        .din(new_Jinkela_wire_6844),
        .dout(new_Jinkela_wire_6845)
    );

    spl4L new_Jinkela_splitter_38 (
        .a(new_Jinkela_wire_197),
        .d(new_Jinkela_wire_198),
        .e(new_Jinkela_wire_199),
        .b(new_Jinkela_wire_200),
        .c(new_Jinkela_wire_201)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_2576),
        .dout(new_Jinkela_wire_2577)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(new_Jinkela_wire_2530),
        .dout(new_Jinkela_wire_2531)
    );

    spl2 new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_194),
        .b(new_Jinkela_wire_195),
        .c(new_Jinkela_wire_196)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_Jinkela_wire_2551),
        .dout(new_Jinkela_wire_2552)
    );

    bfr new_Jinkela_buffer_5016 (
        .din(new_Jinkela_wire_6845),
        .dout(new_Jinkela_wire_6846)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    bfr new_Jinkela_buffer_5065 (
        .din(new_Jinkela_wire_6910),
        .dout(new_Jinkela_wire_6911)
    );

    bfr new_Jinkela_buffer_5035 (
        .din(new_Jinkela_wire_6866),
        .dout(new_Jinkela_wire_6867)
    );

    spl4L new_Jinkela_splitter_39 (
        .a(new_Jinkela_wire_202),
        .d(new_Jinkela_wire_203),
        .e(new_Jinkela_wire_204),
        .b(new_Jinkela_wire_205),
        .c(new_Jinkela_wire_206)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(new_Jinkela_wire_2552),
        .dout(new_Jinkela_wire_2553)
    );

    bfr new_Jinkela_buffer_1627 (
        .din(_0789_),
        .dout(new_Jinkela_wire_2639)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_211),
        .dout(new_Jinkela_wire_212)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(new_Jinkela_wire_2577),
        .dout(new_Jinkela_wire_2578)
    );

    bfr new_Jinkela_buffer_5036 (
        .din(new_Jinkela_wire_6867),
        .dout(new_Jinkela_wire_6868)
    );

    bfr new_Jinkela_buffer_89 (
        .din(G3),
        .dout(new_Jinkela_wire_228)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_2553),
        .dout(new_Jinkela_wire_2554)
    );

    spl4L new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_213),
        .d(new_Jinkela_wire_214),
        .e(new_Jinkela_wire_215),
        .b(new_Jinkela_wire_216),
        .c(new_Jinkela_wire_217)
    );

    bfr new_Jinkela_buffer_5076 (
        .din(new_Jinkela_wire_6923),
        .dout(new_Jinkela_wire_6924)
    );

    bfr new_Jinkela_buffer_86 (
        .din(G36),
        .dout(new_Jinkela_wire_223)
    );

    bfr new_Jinkela_buffer_5066 (
        .din(new_Jinkela_wire_6911),
        .dout(new_Jinkela_wire_6912)
    );

    bfr new_Jinkela_buffer_92 (
        .din(G43),
        .dout(new_Jinkela_wire_233)
    );

    bfr new_Jinkela_buffer_5037 (
        .din(new_Jinkela_wire_6868),
        .dout(new_Jinkela_wire_6869)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_2554),
        .dout(new_Jinkela_wire_2555)
    );

    spl4L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_218),
        .d(new_Jinkela_wire_219),
        .e(new_Jinkela_wire_220),
        .b(new_Jinkela_wire_221),
        .c(new_Jinkela_wire_222)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(new_Jinkela_wire_2585),
        .dout(new_Jinkela_wire_2586)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_2578),
        .dout(new_Jinkela_wire_2579)
    );

    bfr new_Jinkela_buffer_5038 (
        .din(new_Jinkela_wire_6869),
        .dout(new_Jinkela_wire_6870)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_2555),
        .dout(new_Jinkela_wire_2556)
    );

    spl2 new_Jinkela_splitter_712 (
        .a(_1104_),
        .b(new_Jinkela_wire_6949),
        .c(new_Jinkela_wire_6950)
    );

    bfr new_Jinkela_buffer_5067 (
        .din(new_Jinkela_wire_6912),
        .dout(new_Jinkela_wire_6913)
    );

    bfr new_Jinkela_buffer_100 (
        .din(G78),
        .dout(new_Jinkela_wire_243)
    );

    bfr new_Jinkela_buffer_5039 (
        .din(new_Jinkela_wire_6870),
        .dout(new_Jinkela_wire_6871)
    );

    bfr new_Jinkela_buffer_97 (
        .din(G6),
        .dout(new_Jinkela_wire_238)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_2556),
        .dout(new_Jinkela_wire_2557)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    bfr new_Jinkela_buffer_1641 (
        .din(_0520_),
        .dout(new_Jinkela_wire_2653)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_225),
        .b(new_Jinkela_wire_226),
        .c(new_Jinkela_wire_227)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(new_Jinkela_wire_2579),
        .dout(new_Jinkela_wire_2580)
    );

    bfr new_Jinkela_buffer_5040 (
        .din(new_Jinkela_wire_6871),
        .dout(new_Jinkela_wire_6872)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_2557),
        .dout(new_Jinkela_wire_2558)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    bfr new_Jinkela_buffer_5077 (
        .din(new_Jinkela_wire_6924),
        .dout(new_Jinkela_wire_6925)
    );

    bfr new_Jinkela_buffer_5068 (
        .din(new_Jinkela_wire_6913),
        .dout(new_Jinkela_wire_6914)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_233),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_5041 (
        .din(new_Jinkela_wire_6872),
        .dout(new_Jinkela_wire_6873)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_2558),
        .dout(new_Jinkela_wire_2559)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(new_Jinkela_wire_2586),
        .dout(new_Jinkela_wire_2587)
    );

    bfr new_Jinkela_buffer_3373 (
        .din(new_Jinkela_wire_4766),
        .dout(new_Jinkela_wire_4767)
    );

    bfr new_Jinkela_buffer_3317 (
        .din(new_Jinkela_wire_4703),
        .dout(new_Jinkela_wire_4704)
    );

    bfr new_Jinkela_buffer_5866 (
        .din(new_Jinkela_wire_7864),
        .dout(new_Jinkela_wire_7865)
    );

    bfr new_Jinkela_buffer_3339 (
        .din(new_Jinkela_wire_4730),
        .dout(new_Jinkela_wire_4731)
    );

    spl3L new_Jinkela_splitter_782 (
        .a(_0091_),
        .d(new_Jinkela_wire_7914),
        .b(new_Jinkela_wire_7917),
        .c(new_Jinkela_wire_7922)
    );

    spl2 new_Jinkela_splitter_781 (
        .a(new_Jinkela_wire_7891),
        .b(new_Jinkela_wire_7892),
        .c(new_Jinkela_wire_7893)
    );

    bfr new_Jinkela_buffer_3318 (
        .din(new_Jinkela_wire_4704),
        .dout(new_Jinkela_wire_4705)
    );

    bfr new_Jinkela_buffer_5867 (
        .din(new_Jinkela_wire_7865),
        .dout(new_Jinkela_wire_7866)
    );

    bfr new_Jinkela_buffer_3376 (
        .din(new_Jinkela_wire_4769),
        .dout(new_Jinkela_wire_4770)
    );

    bfr new_Jinkela_buffer_5892 (
        .din(_0794_),
        .dout(new_Jinkela_wire_7912)
    );

    bfr new_Jinkela_buffer_5895 (
        .din(_1080_),
        .dout(new_Jinkela_wire_7930)
    );

    bfr new_Jinkela_buffer_3340 (
        .din(new_Jinkela_wire_4731),
        .dout(new_Jinkela_wire_4732)
    );

    bfr new_Jinkela_buffer_5875 (
        .din(new_Jinkela_wire_7894),
        .dout(new_Jinkela_wire_7895)
    );

    bfr new_Jinkela_buffer_3403 (
        .din(new_Jinkela_wire_4796),
        .dout(new_Jinkela_wire_4797)
    );

    bfr new_Jinkela_buffer_5876 (
        .din(new_Jinkela_wire_7895),
        .dout(new_Jinkela_wire_7896)
    );

    bfr new_Jinkela_buffer_3341 (
        .din(new_Jinkela_wire_4732),
        .dout(new_Jinkela_wire_4733)
    );

    bfr new_Jinkela_buffer_5893 (
        .din(new_Jinkela_wire_7912),
        .dout(new_Jinkela_wire_7913)
    );

    bfr new_Jinkela_buffer_3377 (
        .din(new_Jinkela_wire_4770),
        .dout(new_Jinkela_wire_4771)
    );

    bfr new_Jinkela_buffer_5877 (
        .din(new_Jinkela_wire_7896),
        .dout(new_Jinkela_wire_7897)
    );

    bfr new_Jinkela_buffer_3342 (
        .din(new_Jinkela_wire_4733),
        .dout(new_Jinkela_wire_4734)
    );

    spl2 new_Jinkela_splitter_531 (
        .a(_0728_),
        .b(new_Jinkela_wire_4814),
        .c(new_Jinkela_wire_4815)
    );

    bfr new_Jinkela_buffer_5878 (
        .din(new_Jinkela_wire_7897),
        .dout(new_Jinkela_wire_7898)
    );

    bfr new_Jinkela_buffer_3421 (
        .din(_0601_),
        .dout(new_Jinkela_wire_4817)
    );

    bfr new_Jinkela_buffer_3343 (
        .din(new_Jinkela_wire_4734),
        .dout(new_Jinkela_wire_4735)
    );

    bfr new_Jinkela_buffer_5894 (
        .din(_0204_),
        .dout(new_Jinkela_wire_7927)
    );

    bfr new_Jinkela_buffer_3378 (
        .din(new_Jinkela_wire_4771),
        .dout(new_Jinkela_wire_4772)
    );

    bfr new_Jinkela_buffer_5879 (
        .din(new_Jinkela_wire_7898),
        .dout(new_Jinkela_wire_7899)
    );

    bfr new_Jinkela_buffer_3344 (
        .din(new_Jinkela_wire_4735),
        .dout(new_Jinkela_wire_4736)
    );

    bfr new_Jinkela_buffer_5898 (
        .din(_0010_),
        .dout(new_Jinkela_wire_7935)
    );

    bfr new_Jinkela_buffer_3404 (
        .din(new_Jinkela_wire_4797),
        .dout(new_Jinkela_wire_4798)
    );

    bfr new_Jinkela_buffer_5880 (
        .din(new_Jinkela_wire_7899),
        .dout(new_Jinkela_wire_7900)
    );

    bfr new_Jinkela_buffer_3345 (
        .din(new_Jinkela_wire_4736),
        .dout(new_Jinkela_wire_4737)
    );

    spl2 new_Jinkela_splitter_783 (
        .a(new_Jinkela_wire_7914),
        .b(new_Jinkela_wire_7915),
        .c(new_Jinkela_wire_7916)
    );

    bfr new_Jinkela_buffer_3379 (
        .din(new_Jinkela_wire_4772),
        .dout(new_Jinkela_wire_4773)
    );

    bfr new_Jinkela_buffer_5881 (
        .din(new_Jinkela_wire_7900),
        .dout(new_Jinkela_wire_7901)
    );

    bfr new_Jinkela_buffer_3346 (
        .din(new_Jinkela_wire_4737),
        .dout(new_Jinkela_wire_4738)
    );

    spl4L new_Jinkela_splitter_784 (
        .a(new_Jinkela_wire_7917),
        .d(new_Jinkela_wire_7918),
        .e(new_Jinkela_wire_7919),
        .b(new_Jinkela_wire_7920),
        .c(new_Jinkela_wire_7921)
    );

    bfr new_Jinkela_buffer_5915 (
        .din(_1155_),
        .dout(new_Jinkela_wire_7958)
    );

    bfr new_Jinkela_buffer_3406 (
        .din(new_Jinkela_wire_4799),
        .dout(new_Jinkela_wire_4800)
    );

    bfr new_Jinkela_buffer_5882 (
        .din(new_Jinkela_wire_7901),
        .dout(new_Jinkela_wire_7902)
    );

    bfr new_Jinkela_buffer_3347 (
        .din(new_Jinkela_wire_4738),
        .dout(new_Jinkela_wire_4739)
    );

    spl4L new_Jinkela_splitter_785 (
        .a(new_Jinkela_wire_7922),
        .d(new_Jinkela_wire_7923),
        .e(new_Jinkela_wire_7924),
        .b(new_Jinkela_wire_7925),
        .c(new_Jinkela_wire_7926)
    );

    bfr new_Jinkela_buffer_3380 (
        .din(new_Jinkela_wire_4773),
        .dout(new_Jinkela_wire_4774)
    );

    bfr new_Jinkela_buffer_5883 (
        .din(new_Jinkela_wire_7902),
        .dout(new_Jinkela_wire_7903)
    );

    bfr new_Jinkela_buffer_3348 (
        .din(new_Jinkela_wire_4739),
        .dout(new_Jinkela_wire_4740)
    );

    spl2 new_Jinkela_splitter_786 (
        .a(new_Jinkela_wire_7927),
        .b(new_Jinkela_wire_7928),
        .c(new_Jinkela_wire_7929)
    );

    bfr new_Jinkela_buffer_3420 (
        .din(new_Jinkela_wire_4815),
        .dout(new_Jinkela_wire_4816)
    );

    bfr new_Jinkela_buffer_5884 (
        .din(new_Jinkela_wire_7903),
        .dout(new_Jinkela_wire_7904)
    );

    bfr new_Jinkela_buffer_3349 (
        .din(new_Jinkela_wire_4740),
        .dout(new_Jinkela_wire_4741)
    );

    bfr new_Jinkela_buffer_5896 (
        .din(new_Jinkela_wire_7930),
        .dout(new_Jinkela_wire_7931)
    );

    bfr new_Jinkela_buffer_3381 (
        .din(new_Jinkela_wire_4774),
        .dout(new_Jinkela_wire_4775)
    );

    bfr new_Jinkela_buffer_5885 (
        .din(new_Jinkela_wire_7904),
        .dout(new_Jinkela_wire_7905)
    );

    bfr new_Jinkela_buffer_3350 (
        .din(new_Jinkela_wire_4741),
        .dout(new_Jinkela_wire_4742)
    );

    spl2 new_Jinkela_splitter_788 (
        .a(new_net_9),
        .b(new_Jinkela_wire_7936),
        .c(new_Jinkela_wire_7938)
    );

    spl2 new_Jinkela_splitter_791 (
        .a(_0815_),
        .b(new_Jinkela_wire_7961),
        .c(new_Jinkela_wire_7962)
    );

    bfr new_Jinkela_buffer_3407 (
        .din(new_Jinkela_wire_4800),
        .dout(new_Jinkela_wire_4801)
    );

    bfr new_Jinkela_buffer_5886 (
        .din(new_Jinkela_wire_7905),
        .dout(new_Jinkela_wire_7906)
    );

    bfr new_Jinkela_buffer_3351 (
        .din(new_Jinkela_wire_4742),
        .dout(new_Jinkela_wire_4743)
    );

    bfr new_Jinkela_buffer_5897 (
        .din(new_Jinkela_wire_7931),
        .dout(new_Jinkela_wire_7932)
    );

    bfr new_Jinkela_buffer_3382 (
        .din(new_Jinkela_wire_4775),
        .dout(new_Jinkela_wire_4776)
    );

    bfr new_Jinkela_buffer_5887 (
        .din(new_Jinkela_wire_7906),
        .dout(new_Jinkela_wire_7907)
    );

    bfr new_Jinkela_buffer_3352 (
        .din(new_Jinkela_wire_4743),
        .dout(new_Jinkela_wire_4744)
    );

    bfr new_Jinkela_buffer_5900 (
        .din(new_Jinkela_wire_7942),
        .dout(new_Jinkela_wire_7943)
    );

    bfr new_Jinkela_buffer_5888 (
        .din(new_Jinkela_wire_7907),
        .dout(new_Jinkela_wire_7908)
    );

    bfr new_Jinkela_buffer_3434 (
        .din(_0428_),
        .dout(new_Jinkela_wire_4857)
    );

    bfr new_Jinkela_buffer_3353 (
        .din(new_Jinkela_wire_4744),
        .dout(new_Jinkela_wire_4745)
    );

    bfr new_Jinkela_buffer_5899 (
        .din(new_Jinkela_wire_7936),
        .dout(new_Jinkela_wire_7937)
    );

    spl2 new_Jinkela_splitter_787 (
        .a(new_Jinkela_wire_7932),
        .b(new_Jinkela_wire_7933),
        .c(new_Jinkela_wire_7934)
    );

    bfr new_Jinkela_buffer_3383 (
        .din(new_Jinkela_wire_4776),
        .dout(new_Jinkela_wire_4777)
    );

    bfr new_Jinkela_buffer_5889 (
        .din(new_Jinkela_wire_7908),
        .dout(new_Jinkela_wire_7909)
    );

    bfr new_Jinkela_buffer_3354 (
        .din(new_Jinkela_wire_4745),
        .dout(new_Jinkela_wire_4746)
    );

    bfr new_Jinkela_buffer_3408 (
        .din(new_Jinkela_wire_4801),
        .dout(new_Jinkela_wire_4802)
    );

    bfr new_Jinkela_buffer_5890 (
        .din(new_Jinkela_wire_7909),
        .dout(new_Jinkela_wire_7910)
    );

    bfr new_Jinkela_buffer_3355 (
        .din(new_Jinkela_wire_4746),
        .dout(new_Jinkela_wire_4747)
    );

    spl4L new_Jinkela_splitter_789 (
        .a(new_Jinkela_wire_7938),
        .d(new_Jinkela_wire_7939),
        .e(new_Jinkela_wire_7940),
        .b(new_Jinkela_wire_7941),
        .c(new_Jinkela_wire_7942)
    );

    bfr new_Jinkela_buffer_3384 (
        .din(new_Jinkela_wire_4777),
        .dout(new_Jinkela_wire_4778)
    );

    bfr new_Jinkela_buffer_5891 (
        .din(new_Jinkela_wire_7910),
        .dout(new_Jinkela_wire_7911)
    );

    bfr new_Jinkela_buffer_3356 (
        .din(new_Jinkela_wire_4747),
        .dout(new_Jinkela_wire_4748)
    );

    spl2 new_Jinkela_splitter_792 (
        .a(_0753_),
        .b(new_Jinkela_wire_7964),
        .c(new_Jinkela_wire_7965)
    );

    bfr new_Jinkela_buffer_3442 (
        .din(_0295_),
        .dout(new_Jinkela_wire_4865)
    );

    bfr new_Jinkela_buffer_3357 (
        .din(new_Jinkela_wire_4748),
        .dout(new_Jinkela_wire_4749)
    );

    spl2 new_Jinkela_splitter_790 (
        .a(new_Jinkela_wire_7958),
        .b(new_Jinkela_wire_7959),
        .c(new_Jinkela_wire_7960)
    );

    bfr new_Jinkela_buffer_3385 (
        .din(new_Jinkela_wire_4778),
        .dout(new_Jinkela_wire_4779)
    );

    bfr new_Jinkela_buffer_5916 (
        .din(new_Jinkela_wire_7962),
        .dout(new_Jinkela_wire_7963)
    );

    bfr new_Jinkela_buffer_3358 (
        .din(new_Jinkela_wire_4749),
        .dout(new_Jinkela_wire_4750)
    );

    bfr new_Jinkela_buffer_5901 (
        .din(new_Jinkela_wire_7943),
        .dout(new_Jinkela_wire_7944)
    );

    spl2 new_Jinkela_splitter_385 (
        .a(new_Jinkela_wire_2812),
        .b(new_Jinkela_wire_2813),
        .c(new_Jinkela_wire_2814)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_1468),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_1747 (
        .din(new_Jinkela_wire_2758),
        .dout(new_Jinkela_wire_2759)
    );

    spl2 new_Jinkela_splitter_274 (
        .a(new_Jinkela_wire_1512),
        .b(new_Jinkela_wire_1513),
        .c(new_Jinkela_wire_1514)
    );

    bfr new_Jinkela_buffer_1768 (
        .din(new_Jinkela_wire_2794),
        .dout(new_Jinkela_wire_2795)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_1469),
        .dout(new_Jinkela_wire_1470)
    );

    bfr new_Jinkela_buffer_1748 (
        .din(new_Jinkela_wire_2759),
        .dout(new_Jinkela_wire_2760)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_1514),
        .dout(new_Jinkela_wire_1515)
    );

    bfr new_Jinkela_buffer_1783 (
        .din(new_Jinkela_wire_2814),
        .dout(new_Jinkela_wire_2815)
    );

    spl2 new_Jinkela_splitter_265 (
        .a(new_Jinkela_wire_1470),
        .b(new_Jinkela_wire_1471),
        .c(new_Jinkela_wire_1472)
    );

    bfr new_Jinkela_buffer_1749 (
        .din(new_Jinkela_wire_2760),
        .dout(new_Jinkela_wire_2761)
    );

    spl2 new_Jinkela_splitter_266 (
        .a(new_Jinkela_wire_1472),
        .b(new_Jinkela_wire_1473),
        .c(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_1769 (
        .din(new_Jinkela_wire_2795),
        .dout(new_Jinkela_wire_2796)
    );

    bfr new_Jinkela_buffer_1750 (
        .din(new_Jinkela_wire_2761),
        .dout(new_Jinkela_wire_2762)
    );

    spl2 new_Jinkela_splitter_276 (
        .a(new_Jinkela_wire_1524),
        .b(new_Jinkela_wire_1525),
        .c(new_Jinkela_wire_1526)
    );

    spl2 new_Jinkela_splitter_267 (
        .a(new_Jinkela_wire_1474),
        .b(new_Jinkela_wire_1475),
        .c(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_1818 (
        .din(_1049_),
        .dout(new_Jinkela_wire_2861)
    );

    bfr new_Jinkela_buffer_1751 (
        .din(new_Jinkela_wire_2762),
        .dout(new_Jinkela_wire_2763)
    );

    spl2 new_Jinkela_splitter_268 (
        .a(new_Jinkela_wire_1476),
        .b(new_Jinkela_wire_1477),
        .c(new_Jinkela_wire_1478)
    );

    bfr new_Jinkela_buffer_1788 (
        .din(new_Jinkela_wire_2821),
        .dout(new_Jinkela_wire_2822)
    );

    bfr new_Jinkela_buffer_1770 (
        .din(new_Jinkela_wire_2796),
        .dout(new_Jinkela_wire_2797)
    );

    bfr new_Jinkela_buffer_1752 (
        .din(new_Jinkela_wire_2763),
        .dout(new_Jinkela_wire_2764)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_1515),
        .dout(new_Jinkela_wire_1516)
    );

    spl3L new_Jinkela_splitter_269 (
        .a(new_Jinkela_wire_1478),
        .d(new_Jinkela_wire_1479),
        .b(new_Jinkela_wire_1480),
        .c(new_Jinkela_wire_1481)
    );

    spl4L new_Jinkela_splitter_280 (
        .a(new_Jinkela_wire_1533),
        .d(new_Jinkela_wire_1534),
        .e(new_Jinkela_wire_1535),
        .b(new_Jinkela_wire_1536),
        .c(new_Jinkela_wire_1537)
    );

    bfr new_Jinkela_buffer_1771 (
        .din(new_Jinkela_wire_2797),
        .dout(new_Jinkela_wire_2798)
    );

    spl2 new_Jinkela_splitter_275 (
        .a(new_Jinkela_wire_1516),
        .b(new_Jinkela_wire_1517),
        .c(new_Jinkela_wire_1518)
    );

    spl2 new_Jinkela_splitter_386 (
        .a(new_Jinkela_wire_2815),
        .b(new_Jinkela_wire_2816),
        .c(new_Jinkela_wire_2817)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_1481),
        .dout(new_Jinkela_wire_1482)
    );

    bfr new_Jinkela_buffer_1772 (
        .din(new_Jinkela_wire_2798),
        .dout(new_Jinkela_wire_2799)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_1518),
        .dout(new_Jinkela_wire_1519)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_1482),
        .dout(new_Jinkela_wire_1483)
    );

    bfr new_Jinkela_buffer_1773 (
        .din(new_Jinkela_wire_2799),
        .dout(new_Jinkela_wire_2800)
    );

    spl4L new_Jinkela_splitter_279 (
        .a(new_Jinkela_wire_1531),
        .d(new_Jinkela_wire_1532),
        .e(new_Jinkela_wire_1533),
        .b(new_Jinkela_wire_1538),
        .c(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_1808 (
        .din(new_Jinkela_wire_2843),
        .dout(new_Jinkela_wire_2844)
    );

    bfr new_Jinkela_buffer_1789 (
        .din(new_Jinkela_wire_2822),
        .dout(new_Jinkela_wire_2823)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_1774 (
        .din(new_Jinkela_wire_2800),
        .dout(new_Jinkela_wire_2801)
    );

    spl3L new_Jinkela_splitter_278 (
        .a(new_Jinkela_wire_1527),
        .d(new_Jinkela_wire_1528),
        .b(new_Jinkela_wire_1529),
        .c(new_Jinkela_wire_1530)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_1519),
        .dout(new_Jinkela_wire_1520)
    );

    bfr new_Jinkela_buffer_1809 (
        .din(new_Jinkela_wire_2847),
        .dout(new_Jinkela_wire_2848)
    );

    bfr new_Jinkela_buffer_1790 (
        .din(new_Jinkela_wire_2823),
        .dout(new_Jinkela_wire_2824)
    );

    spl3L new_Jinkela_splitter_283 (
        .a(G163),
        .d(new_Jinkela_wire_1552),
        .b(new_Jinkela_wire_1557),
        .c(new_Jinkela_wire_1562)
    );

    bfr new_Jinkela_buffer_1775 (
        .din(new_Jinkela_wire_2801),
        .dout(new_Jinkela_wire_2802)
    );

    spl4L new_Jinkela_splitter_281 (
        .a(new_Jinkela_wire_1538),
        .d(new_Jinkela_wire_1539),
        .e(new_Jinkela_wire_1540),
        .b(new_Jinkela_wire_1541),
        .c(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_1520),
        .dout(new_Jinkela_wire_1521)
    );

    bfr new_Jinkela_buffer_1776 (
        .din(new_Jinkela_wire_2802),
        .dout(new_Jinkela_wire_2803)
    );

    spl4L new_Jinkela_splitter_285 (
        .a(new_Jinkela_wire_1557),
        .d(new_Jinkela_wire_1558),
        .e(new_Jinkela_wire_1559),
        .b(new_Jinkela_wire_1560),
        .c(new_Jinkela_wire_1561)
    );

    spl4L new_Jinkela_splitter_282 (
        .a(new_Jinkela_wire_1543),
        .d(new_Jinkela_wire_1544),
        .e(new_Jinkela_wire_1545),
        .b(new_Jinkela_wire_1546),
        .c(new_Jinkela_wire_1547)
    );

    bfr new_Jinkela_buffer_1791 (
        .din(new_Jinkela_wire_2824),
        .dout(new_Jinkela_wire_2825)
    );

    bfr new_Jinkela_buffer_1777 (
        .din(new_Jinkela_wire_2803),
        .dout(new_Jinkela_wire_2804)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_1568),
        .dout(new_Jinkela_wire_1569)
    );

    bfr new_Jinkela_buffer_767 (
        .din(G59),
        .dout(new_Jinkela_wire_1567)
    );

    bfr new_Jinkela_buffer_1810 (
        .din(new_Jinkela_wire_2848),
        .dout(new_Jinkela_wire_2849)
    );

    bfr new_Jinkela_buffer_1792 (
        .din(new_Jinkela_wire_2825),
        .dout(new_Jinkela_wire_2826)
    );

    bfr new_Jinkela_buffer_772 (
        .din(G75),
        .dout(new_Jinkela_wire_1572)
    );

    spl4L new_Jinkela_splitter_284 (
        .a(new_Jinkela_wire_1552),
        .d(new_Jinkela_wire_1553),
        .e(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_1555),
        .c(new_Jinkela_wire_1556)
    );

    spl4L new_Jinkela_splitter_389 (
        .a(new_Jinkela_wire_2855),
        .d(new_Jinkela_wire_2856),
        .e(new_Jinkela_wire_2857),
        .b(new_Jinkela_wire_2858),
        .c(new_Jinkela_wire_2859)
    );

    spl2 new_Jinkela_splitter_288 (
        .a(G167),
        .b(new_Jinkela_wire_1577),
        .c(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_1793 (
        .din(new_Jinkela_wire_2826),
        .dout(new_Jinkela_wire_2827)
    );

    spl4L new_Jinkela_splitter_286 (
        .a(new_Jinkela_wire_1562),
        .d(new_Jinkela_wire_1563),
        .e(new_Jinkela_wire_1564),
        .b(new_Jinkela_wire_1565),
        .c(new_Jinkela_wire_1566)
    );

    bfr new_Jinkela_buffer_1819 (
        .din(_0383_),
        .dout(new_Jinkela_wire_2862)
    );

    bfr new_Jinkela_buffer_1811 (
        .din(new_Jinkela_wire_2849),
        .dout(new_Jinkela_wire_2850)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_1567),
        .dout(new_Jinkela_wire_1568)
    );

    bfr new_Jinkela_buffer_1794 (
        .din(new_Jinkela_wire_2827),
        .dout(new_Jinkela_wire_2828)
    );

    bfr new_Jinkela_buffer_1817 (
        .din(new_Jinkela_wire_2859),
        .dout(new_Jinkela_wire_2860)
    );

    bfr new_Jinkela_buffer_1795 (
        .din(new_Jinkela_wire_2828),
        .dout(new_Jinkela_wire_2829)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1572),
        .dout(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_1569),
        .dout(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_1812 (
        .din(new_Jinkela_wire_2850),
        .dout(new_Jinkela_wire_2851)
    );

    spl4L new_Jinkela_splitter_290 (
        .a(new_Jinkela_wire_1580),
        .d(new_Jinkela_wire_1581),
        .e(new_Jinkela_wire_1582),
        .b(new_Jinkela_wire_1583),
        .c(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_1796 (
        .din(new_Jinkela_wire_2829),
        .dout(new_Jinkela_wire_2830)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_1797 (
        .din(new_Jinkela_wire_2830),
        .dout(new_Jinkela_wire_2831)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1573),
        .dout(new_Jinkela_wire_1574)
    );

    spl3L new_Jinkela_splitter_390 (
        .a(_0256_),
        .d(new_Jinkela_wire_2863),
        .b(new_Jinkela_wire_2866),
        .c(new_Jinkela_wire_2871)
    );

    bfr new_Jinkela_buffer_1813 (
        .din(new_Jinkela_wire_2851),
        .dout(new_Jinkela_wire_2852)
    );

    spl3L new_Jinkela_splitter_293 (
        .a(G175),
        .d(new_Jinkela_wire_1592),
        .b(new_Jinkela_wire_1593),
        .c(new_Jinkela_wire_1594)
    );

    bfr new_Jinkela_buffer_1798 (
        .din(new_Jinkela_wire_2831),
        .dout(new_Jinkela_wire_2832)
    );

    spl2 new_Jinkela_splitter_287 (
        .a(new_Jinkela_wire_1574),
        .b(new_Jinkela_wire_1575),
        .c(new_Jinkela_wire_1576)
    );

    bfr new_Jinkela_buffer_775 (
        .din(G28),
        .dout(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_1816 (
        .din(new_Jinkela_wire_2854),
        .dout(new_Jinkela_wire_2855)
    );

    bfr new_Jinkela_buffer_777 (
        .din(G58),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_1799 (
        .din(new_Jinkela_wire_2832),
        .dout(new_Jinkela_wire_2833)
    );

    or_bb _2582_ (
        .a(new_Jinkela_wire_6699),
        .b(new_Jinkela_wire_1116),
        .c(_0562_)
    );

    bfr new_Jinkela_buffer_3328 (
        .din(new_Jinkela_wire_4719),
        .dout(new_Jinkela_wire_4720)
    );

    bfr new_Jinkela_buffer_5267 (
        .din(new_Jinkela_wire_7173),
        .dout(new_Jinkela_wire_7174)
    );

    and_bi _2583_ (
        .a(new_Jinkela_wire_5080),
        .b(new_Jinkela_wire_1682),
        .c(new_net_2353)
    );

    bfr new_Jinkela_buffer_4663 (
        .din(new_Jinkela_wire_6377),
        .dout(new_Jinkela_wire_6378)
    );

    bfr new_Jinkela_buffer_3296 (
        .din(new_Jinkela_wire_4682),
        .dout(new_Jinkela_wire_4683)
    );

    bfr new_Jinkela_buffer_4640 (
        .din(new_Jinkela_wire_6344),
        .dout(new_Jinkela_wire_6345)
    );

    spl2 new_Jinkela_splitter_741 (
        .a(new_Jinkela_wire_7210),
        .b(new_Jinkela_wire_7211),
        .c(new_Jinkela_wire_7212)
    );

    and_ii _2584_ (
        .a(new_Jinkela_wire_6682),
        .b(new_Jinkela_wire_1266),
        .c(_0563_)
    );

    bfr new_Jinkela_buffer_3374 (
        .din(_0536_),
        .dout(new_Jinkela_wire_4768)
    );

    bfr new_Jinkela_buffer_4655 (
        .din(new_Jinkela_wire_6367),
        .dout(new_Jinkela_wire_6368)
    );

    bfr new_Jinkela_buffer_5268 (
        .din(new_Jinkela_wire_7174),
        .dout(new_Jinkela_wire_7175)
    );

    and_bi _2585_ (
        .a(new_Jinkela_wire_7606),
        .b(new_Jinkela_wire_3060),
        .c(new_net_2409)
    );

    bfr new_Jinkela_buffer_3297 (
        .din(new_Jinkela_wire_4683),
        .dout(new_Jinkela_wire_4684)
    );

    bfr new_Jinkela_buffer_4641 (
        .din(new_Jinkela_wire_6345),
        .dout(new_Jinkela_wire_6346)
    );

    or_bb _2586_ (
        .a(new_Jinkela_wire_3415),
        .b(new_Jinkela_wire_1483),
        .c(_0564_)
    );

    bfr new_Jinkela_buffer_3329 (
        .din(new_Jinkela_wire_4720),
        .dout(new_Jinkela_wire_4721)
    );

    bfr new_Jinkela_buffer_5269 (
        .din(new_Jinkela_wire_7175),
        .dout(new_Jinkela_wire_7176)
    );

    and_bi _2587_ (
        .a(new_Jinkela_wire_1475),
        .b(new_Jinkela_wire_3753),
        .c(_0565_)
    );

    bfr new_Jinkela_buffer_4664 (
        .din(_0859_),
        .dout(new_Jinkela_wire_6382)
    );

    bfr new_Jinkela_buffer_3298 (
        .din(new_Jinkela_wire_4684),
        .dout(new_Jinkela_wire_4685)
    );

    bfr new_Jinkela_buffer_4642 (
        .din(new_Jinkela_wire_6346),
        .dout(new_Jinkela_wire_6347)
    );

    or_bb _2588_ (
        .a(_0565_),
        .b(new_Jinkela_wire_3518),
        .c(_0566_)
    );

    bfr new_Jinkela_buffer_3366 (
        .din(new_Jinkela_wire_4759),
        .dout(new_Jinkela_wire_4760)
    );

    bfr new_Jinkela_buffer_4656 (
        .din(new_Jinkela_wire_6368),
        .dout(new_Jinkela_wire_6369)
    );

    bfr new_Jinkela_buffer_5270 (
        .din(new_Jinkela_wire_7176),
        .dout(new_Jinkela_wire_7177)
    );

    and_bi _2589_ (
        .a(_0564_),
        .b(new_Jinkela_wire_5118),
        .c(_0567_)
    );

    bfr new_Jinkela_buffer_3299 (
        .din(new_Jinkela_wire_4685),
        .dout(new_Jinkela_wire_4686)
    );

    bfr new_Jinkela_buffer_4643 (
        .din(new_Jinkela_wire_6347),
        .dout(new_Jinkela_wire_6348)
    );

    bfr new_Jinkela_buffer_5292 (
        .din(new_Jinkela_wire_7214),
        .dout(new_Jinkela_wire_7215)
    );

    and_bi _2590_ (
        .a(new_Jinkela_wire_1505),
        .b(new_Jinkela_wire_6417),
        .c(_0568_)
    );

    bfr new_Jinkela_buffer_3330 (
        .din(new_Jinkela_wire_4721),
        .dout(new_Jinkela_wire_4722)
    );

    bfr new_Jinkela_buffer_5271 (
        .din(new_Jinkela_wire_7177),
        .dout(new_Jinkela_wire_7178)
    );

    and_bi _2591_ (
        .a(new_Jinkela_wire_727),
        .b(new_Jinkela_wire_2873),
        .c(_0569_)
    );

    bfr new_Jinkela_buffer_4689 (
        .din(_0168_),
        .dout(new_Jinkela_wire_6407)
    );

    bfr new_Jinkela_buffer_3300 (
        .din(new_Jinkela_wire_4686),
        .dout(new_Jinkela_wire_4687)
    );

    bfr new_Jinkela_buffer_4657 (
        .din(new_Jinkela_wire_6369),
        .dout(new_Jinkela_wire_6370)
    );

    bfr new_Jinkela_buffer_5293 (
        .din(new_Jinkela_wire_7215),
        .dout(new_Jinkela_wire_7216)
    );

    or_bb _2592_ (
        .a(_0569_),
        .b(_0568_),
        .c(_0570_)
    );

    bfr new_Jinkela_buffer_3370 (
        .din(new_Jinkela_wire_4763),
        .dout(new_Jinkela_wire_4764)
    );

    spl3L new_Jinkela_splitter_660 (
        .a(_0258_),
        .d(new_Jinkela_wire_6413),
        .b(new_Jinkela_wire_6416),
        .c(new_Jinkela_wire_6421)
    );

    bfr new_Jinkela_buffer_5272 (
        .din(new_Jinkela_wire_7178),
        .dout(new_Jinkela_wire_7179)
    );

    or_bb _2593_ (
        .a(new_Jinkela_wire_1820),
        .b(_0567_),
        .c(new_net_2489)
    );

    bfr new_Jinkela_buffer_3301 (
        .din(new_Jinkela_wire_4687),
        .dout(new_Jinkela_wire_4688)
    );

    bfr new_Jinkela_buffer_4658 (
        .din(new_Jinkela_wire_6370),
        .dout(new_Jinkela_wire_6371)
    );

    bfr new_Jinkela_buffer_5339 (
        .din(_0349_),
        .dout(new_Jinkela_wire_7266)
    );

    or_bb _2594_ (
        .a(new_Jinkela_wire_3412),
        .b(new_Jinkela_wire_399),
        .c(_0571_)
    );

    bfr new_Jinkela_buffer_5320 (
        .din(_0371_),
        .dout(new_Jinkela_wire_7247)
    );

    bfr new_Jinkela_buffer_3331 (
        .din(new_Jinkela_wire_4722),
        .dout(new_Jinkela_wire_4723)
    );

    bfr new_Jinkela_buffer_4665 (
        .din(new_Jinkela_wire_6382),
        .dout(new_Jinkela_wire_6383)
    );

    bfr new_Jinkela_buffer_5273 (
        .din(new_Jinkela_wire_7179),
        .dout(new_Jinkela_wire_7180)
    );

    and_bi _2595_ (
        .a(new_Jinkela_wire_389),
        .b(new_Jinkela_wire_3750),
        .c(_0572_)
    );

    bfr new_Jinkela_buffer_3302 (
        .din(new_Jinkela_wire_4688),
        .dout(new_Jinkela_wire_4689)
    );

    bfr new_Jinkela_buffer_4659 (
        .din(new_Jinkela_wire_6371),
        .dout(new_Jinkela_wire_6372)
    );

    bfr new_Jinkela_buffer_5294 (
        .din(new_Jinkela_wire_7216),
        .dout(new_Jinkela_wire_7217)
    );

    or_bb _2596_ (
        .a(_0572_),
        .b(new_Jinkela_wire_3982),
        .c(_0573_)
    );

    bfr new_Jinkela_buffer_3367 (
        .din(new_Jinkela_wire_4760),
        .dout(new_Jinkela_wire_4761)
    );

    bfr new_Jinkela_buffer_4737 (
        .din(_0395_),
        .dout(new_Jinkela_wire_6472)
    );

    bfr new_Jinkela_buffer_5274 (
        .din(new_Jinkela_wire_7180),
        .dout(new_Jinkela_wire_7181)
    );

    and_bi _2597_ (
        .a(_0571_),
        .b(new_Jinkela_wire_1988),
        .c(_0574_)
    );

    bfr new_Jinkela_buffer_3303 (
        .din(new_Jinkela_wire_4689),
        .dout(new_Jinkela_wire_4690)
    );

    bfr new_Jinkela_buffer_4660 (
        .din(new_Jinkela_wire_6372),
        .dout(new_Jinkela_wire_6373)
    );

    bfr new_Jinkela_buffer_5314 (
        .din(new_Jinkela_wire_7240),
        .dout(new_Jinkela_wire_7241)
    );

    and_bi _2598_ (
        .a(new_Jinkela_wire_1506),
        .b(new_Jinkela_wire_7877),
        .c(_0575_)
    );

    bfr new_Jinkela_buffer_3332 (
        .din(new_Jinkela_wire_4723),
        .dout(new_Jinkela_wire_4724)
    );

    bfr new_Jinkela_buffer_4666 (
        .din(new_Jinkela_wire_6383),
        .dout(new_Jinkela_wire_6384)
    );

    bfr new_Jinkela_buffer_5275 (
        .din(new_Jinkela_wire_7181),
        .dout(new_Jinkela_wire_7182)
    );

    and_bi _2599_ (
        .a(new_Jinkela_wire_728),
        .b(new_Jinkela_wire_5804),
        .c(_0576_)
    );

    bfr new_Jinkela_buffer_3304 (
        .din(new_Jinkela_wire_4690),
        .dout(new_Jinkela_wire_4691)
    );

    bfr new_Jinkela_buffer_4661 (
        .din(new_Jinkela_wire_6373),
        .dout(new_Jinkela_wire_6374)
    );

    bfr new_Jinkela_buffer_5295 (
        .din(new_Jinkela_wire_7217),
        .dout(new_Jinkela_wire_7218)
    );

    or_bb _2600_ (
        .a(_0576_),
        .b(_0575_),
        .c(_0577_)
    );

    bfr new_Jinkela_buffer_3402 (
        .din(_1230_),
        .dout(new_Jinkela_wire_4796)
    );

    bfr new_Jinkela_buffer_5276 (
        .din(new_Jinkela_wire_7182),
        .dout(new_Jinkela_wire_7183)
    );

    or_bb _2601_ (
        .a(new_Jinkela_wire_6316),
        .b(_0574_),
        .c(new_net_2349)
    );

    bfr new_Jinkela_buffer_4690 (
        .din(new_Jinkela_wire_6407),
        .dout(new_Jinkela_wire_6408)
    );

    bfr new_Jinkela_buffer_3305 (
        .din(new_Jinkela_wire_4691),
        .dout(new_Jinkela_wire_4692)
    );

    bfr new_Jinkela_buffer_4667 (
        .din(new_Jinkela_wire_6384),
        .dout(new_Jinkela_wire_6385)
    );

    bfr new_Jinkela_buffer_5315 (
        .din(new_Jinkela_wire_7241),
        .dout(new_Jinkela_wire_7242)
    );

    and_bi _2602_ (
        .a(new_Jinkela_wire_4570),
        .b(new_Jinkela_wire_7651),
        .c(new_net_2433)
    );

    bfr new_Jinkela_buffer_3333 (
        .din(new_Jinkela_wire_4724),
        .dout(new_Jinkela_wire_4725)
    );

    bfr new_Jinkela_buffer_5296 (
        .din(new_Jinkela_wire_7218),
        .dout(new_Jinkela_wire_7219)
    );

    and_ii _2603_ (
        .a(new_Jinkela_wire_1951),
        .b(new_Jinkela_wire_3165),
        .c(new_net_2421)
    );

    bfr new_Jinkela_buffer_3306 (
        .din(new_Jinkela_wire_4692),
        .dout(new_Jinkela_wire_4693)
    );

    bfr new_Jinkela_buffer_4668 (
        .din(new_Jinkela_wire_6385),
        .dout(new_Jinkela_wire_6386)
    );

    bfr new_Jinkela_buffer_5321 (
        .din(new_Jinkela_wire_7247),
        .dout(new_Jinkela_wire_7248)
    );

    or_bb _2604_ (
        .a(new_Jinkela_wire_7129),
        .b(new_Jinkela_wire_6889),
        .c(new_net_2385)
    );

    bfr new_Jinkela_buffer_3368 (
        .din(new_Jinkela_wire_4761),
        .dout(new_Jinkela_wire_4762)
    );

    bfr new_Jinkela_buffer_5297 (
        .din(new_Jinkela_wire_7219),
        .dout(new_Jinkela_wire_7220)
    );

    or_bi _2605_ (
        .a(new_Jinkela_wire_4573),
        .b(new_Jinkela_wire_2769),
        .c(new_net_2497)
    );

    bfr new_Jinkela_buffer_4691 (
        .din(new_Jinkela_wire_6408),
        .dout(new_Jinkela_wire_6409)
    );

    bfr new_Jinkela_buffer_3307 (
        .din(new_Jinkela_wire_4693),
        .dout(new_Jinkela_wire_4694)
    );

    bfr new_Jinkela_buffer_4669 (
        .din(new_Jinkela_wire_6386),
        .dout(new_Jinkela_wire_6387)
    );

    bfr new_Jinkela_buffer_5316 (
        .din(new_Jinkela_wire_7242),
        .dout(new_Jinkela_wire_7243)
    );

    bfr new_Jinkela_buffer_3334 (
        .din(new_Jinkela_wire_4725),
        .dout(new_Jinkela_wire_4726)
    );

    bfr new_Jinkela_buffer_5298 (
        .din(new_Jinkela_wire_7220),
        .dout(new_Jinkela_wire_7221)
    );

    bfr new_Jinkela_buffer_4693 (
        .din(_0235_),
        .dout(new_Jinkela_wire_6426)
    );

    bfr new_Jinkela_buffer_3308 (
        .din(new_Jinkela_wire_4694),
        .dout(new_Jinkela_wire_4695)
    );

    bfr new_Jinkela_buffer_4670 (
        .din(new_Jinkela_wire_6387),
        .dout(new_Jinkela_wire_6388)
    );

    spl2 new_Jinkela_splitter_743 (
        .a(new_net_10),
        .b(new_Jinkela_wire_7289),
        .c(new_Jinkela_wire_7291)
    );

    bfr new_Jinkela_buffer_5382 (
        .din(new_net_2351),
        .dout(new_Jinkela_wire_7315)
    );

    bfr new_Jinkela_buffer_3371 (
        .din(new_Jinkela_wire_4764),
        .dout(new_Jinkela_wire_4765)
    );

    spl2 new_Jinkela_splitter_664 (
        .a(_0671_),
        .b(new_Jinkela_wire_6470),
        .c(new_Jinkela_wire_6471)
    );

    bfr new_Jinkela_buffer_5299 (
        .din(new_Jinkela_wire_7221),
        .dout(new_Jinkela_wire_7222)
    );

    bfr new_Jinkela_buffer_4692 (
        .din(new_Jinkela_wire_6409),
        .dout(new_Jinkela_wire_6410)
    );

    bfr new_Jinkela_buffer_3309 (
        .din(new_Jinkela_wire_4695),
        .dout(new_Jinkela_wire_4696)
    );

    bfr new_Jinkela_buffer_4671 (
        .din(new_Jinkela_wire_6388),
        .dout(new_Jinkela_wire_6389)
    );

    bfr new_Jinkela_buffer_5317 (
        .din(new_Jinkela_wire_7243),
        .dout(new_Jinkela_wire_7244)
    );

    bfr new_Jinkela_buffer_3335 (
        .din(new_Jinkela_wire_4726),
        .dout(new_Jinkela_wire_4727)
    );

    bfr new_Jinkela_buffer_5300 (
        .din(new_Jinkela_wire_7222),
        .dout(new_Jinkela_wire_7223)
    );

    spl4L new_Jinkela_splitter_662 (
        .a(new_Jinkela_wire_6416),
        .d(new_Jinkela_wire_6417),
        .e(new_Jinkela_wire_6418),
        .b(new_Jinkela_wire_6419),
        .c(new_Jinkela_wire_6420)
    );

    bfr new_Jinkela_buffer_3310 (
        .din(new_Jinkela_wire_4696),
        .dout(new_Jinkela_wire_4697)
    );

    bfr new_Jinkela_buffer_4672 (
        .din(new_Jinkela_wire_6389),
        .dout(new_Jinkela_wire_6390)
    );

    bfr new_Jinkela_buffer_5322 (
        .din(new_Jinkela_wire_7248),
        .dout(new_Jinkela_wire_7249)
    );

    bfr new_Jinkela_buffer_3375 (
        .din(new_Jinkela_wire_4768),
        .dout(new_Jinkela_wire_4769)
    );

    bfr new_Jinkela_buffer_4694 (
        .din(_0850_),
        .dout(new_Jinkela_wire_6427)
    );

    bfr new_Jinkela_buffer_5301 (
        .din(new_Jinkela_wire_7223),
        .dout(new_Jinkela_wire_7224)
    );

    spl2 new_Jinkela_splitter_659 (
        .a(new_Jinkela_wire_6410),
        .b(new_Jinkela_wire_6411),
        .c(new_Jinkela_wire_6412)
    );

    bfr new_Jinkela_buffer_3311 (
        .din(new_Jinkela_wire_4697),
        .dout(new_Jinkela_wire_4698)
    );

    bfr new_Jinkela_buffer_4673 (
        .din(new_Jinkela_wire_6390),
        .dout(new_Jinkela_wire_6391)
    );

    bfr new_Jinkela_buffer_5318 (
        .din(new_Jinkela_wire_7244),
        .dout(new_Jinkela_wire_7245)
    );

    bfr new_Jinkela_buffer_3336 (
        .din(new_Jinkela_wire_4727),
        .dout(new_Jinkela_wire_4728)
    );

    bfr new_Jinkela_buffer_5302 (
        .din(new_Jinkela_wire_7224),
        .dout(new_Jinkela_wire_7225)
    );

    bfr new_Jinkela_buffer_3312 (
        .din(new_Jinkela_wire_4698),
        .dout(new_Jinkela_wire_4699)
    );

    bfr new_Jinkela_buffer_4674 (
        .din(new_Jinkela_wire_6391),
        .dout(new_Jinkela_wire_6392)
    );

    bfr new_Jinkela_buffer_5340 (
        .din(new_Jinkela_wire_7266),
        .dout(new_Jinkela_wire_7267)
    );

    bfr new_Jinkela_buffer_3372 (
        .din(new_Jinkela_wire_4765),
        .dout(new_Jinkela_wire_4766)
    );

    spl4L new_Jinkela_splitter_663 (
        .a(new_Jinkela_wire_6421),
        .d(new_Jinkela_wire_6422),
        .e(new_Jinkela_wire_6423),
        .b(new_Jinkela_wire_6424),
        .c(new_Jinkela_wire_6425)
    );

    bfr new_Jinkela_buffer_5303 (
        .din(new_Jinkela_wire_7225),
        .dout(new_Jinkela_wire_7226)
    );

    bfr new_Jinkela_buffer_3313 (
        .din(new_Jinkela_wire_4699),
        .dout(new_Jinkela_wire_4700)
    );

    bfr new_Jinkela_buffer_4675 (
        .din(new_Jinkela_wire_6392),
        .dout(new_Jinkela_wire_6393)
    );

    bfr new_Jinkela_buffer_5319 (
        .din(new_Jinkela_wire_7245),
        .dout(new_Jinkela_wire_7246)
    );

    bfr new_Jinkela_buffer_3337 (
        .din(new_Jinkela_wire_4728),
        .dout(new_Jinkela_wire_4729)
    );

    spl2 new_Jinkela_splitter_661 (
        .a(new_Jinkela_wire_6413),
        .b(new_Jinkela_wire_6414),
        .c(new_Jinkela_wire_6415)
    );

    bfr new_Jinkela_buffer_5304 (
        .din(new_Jinkela_wire_7226),
        .dout(new_Jinkela_wire_7227)
    );

    bfr new_Jinkela_buffer_3314 (
        .din(new_Jinkela_wire_4700),
        .dout(new_Jinkela_wire_4701)
    );

    bfr new_Jinkela_buffer_4676 (
        .din(new_Jinkela_wire_6393),
        .dout(new_Jinkela_wire_6394)
    );

    bfr new_Jinkela_buffer_5323 (
        .din(new_Jinkela_wire_7249),
        .dout(new_Jinkela_wire_7250)
    );

    bfr new_Jinkela_buffer_3405 (
        .din(_0299_),
        .dout(new_Jinkela_wire_4799)
    );

    bfr new_Jinkela_buffer_4702 (
        .din(new_net_2477),
        .dout(new_Jinkela_wire_6435)
    );

    bfr new_Jinkela_buffer_5305 (
        .din(new_Jinkela_wire_7227),
        .dout(new_Jinkela_wire_7228)
    );

    bfr new_Jinkela_buffer_3315 (
        .din(new_Jinkela_wire_4701),
        .dout(new_Jinkela_wire_4702)
    );

    bfr new_Jinkela_buffer_4677 (
        .din(new_Jinkela_wire_6394),
        .dout(new_Jinkela_wire_6395)
    );

    bfr new_Jinkela_buffer_3338 (
        .din(new_Jinkela_wire_4729),
        .dout(new_Jinkela_wire_4730)
    );

    bfr new_Jinkela_buffer_4695 (
        .din(new_Jinkela_wire_6427),
        .dout(new_Jinkela_wire_6428)
    );

    bfr new_Jinkela_buffer_5306 (
        .din(new_Jinkela_wire_7228),
        .dout(new_Jinkela_wire_7229)
    );

    bfr new_Jinkela_buffer_3316 (
        .din(new_Jinkela_wire_4702),
        .dout(new_Jinkela_wire_4703)
    );

    bfr new_Jinkela_buffer_4678 (
        .din(new_Jinkela_wire_6395),
        .dout(new_Jinkela_wire_6396)
    );

    bfr new_Jinkela_buffer_5324 (
        .din(new_Jinkela_wire_7250),
        .dout(new_Jinkela_wire_7251)
    );

    and_bi _1865_ (
        .a(new_Jinkela_wire_3772),
        .b(_1153_),
        .c(_1154_)
    );

    and_ii _1866_ (
        .a(_1154_),
        .b(_1150_),
        .c(_1155_)
    );

    and_ii _1867_ (
        .a(new_Jinkela_wire_7959),
        .b(new_Jinkela_wire_3833),
        .c(_1156_)
    );

    and_bb _1868_ (
        .a(new_Jinkela_wire_7960),
        .b(new_Jinkela_wire_3835),
        .c(_1157_)
    );

    and_ii _1869_ (
        .a(_1157_),
        .b(_1156_),
        .c(_1158_)
    );

    and_bb _1870_ (
        .a(new_Jinkela_wire_3662),
        .b(new_Jinkela_wire_4980),
        .c(_1159_)
    );

    and_ii _1871_ (
        .a(new_Jinkela_wire_3663),
        .b(new_Jinkela_wire_4981),
        .c(_1160_)
    );

    or_bb _1872_ (
        .a(_1160_),
        .b(_1159_),
        .c(_1161_)
    );

    or_bb _1873_ (
        .a(new_Jinkela_wire_1314),
        .b(new_Jinkela_wire_51),
        .c(_1162_)
    );

    and_bi _1874_ (
        .a(new_Jinkela_wire_1313),
        .b(new_Jinkela_wire_415),
        .c(_1163_)
    );

    and_bi _1875_ (
        .a(_1162_),
        .b(_1163_),
        .c(_1164_)
    );

    or_bb _1876_ (
        .a(_1164_),
        .b(new_Jinkela_wire_5702),
        .c(_1165_)
    );

    or_ii _1877_ (
        .a(new_Jinkela_wire_1315),
        .b(new_Jinkela_wire_1209),
        .c(_1166_)
    );

    and_bi _1878_ (
        .a(new_Jinkela_wire_1544),
        .b(new_Jinkela_wire_1310),
        .c(_1167_)
    );

    and_bi _1879_ (
        .a(_1166_),
        .b(_1167_),
        .c(_1168_)
    );

    and_bi _1880_ (
        .a(new_Jinkela_wire_5700),
        .b(_1168_),
        .c(_1169_)
    );

    and_bi _1881_ (
        .a(_1165_),
        .b(_1169_),
        .c(_1170_)
    );

    or_bb _1882_ (
        .a(new_Jinkela_wire_166),
        .b(new_Jinkela_wire_53),
        .c(_1171_)
    );

    and_bi _1883_ (
        .a(new_Jinkela_wire_159),
        .b(new_Jinkela_wire_410),
        .c(_1172_)
    );

    and_bi _1884_ (
        .a(_1171_),
        .b(_1172_),
        .c(_1173_)
    );

    or_bb _1885_ (
        .a(_1173_),
        .b(new_Jinkela_wire_7008),
        .c(_1174_)
    );

    or_ii _1886_ (
        .a(new_Jinkela_wire_164),
        .b(new_Jinkela_wire_1207),
        .c(_1175_)
    );

    and_bi _1887_ (
        .a(new_Jinkela_wire_1542),
        .b(new_Jinkela_wire_158),
        .c(_1176_)
    );

    and_bi _1888_ (
        .a(_1175_),
        .b(_1176_),
        .c(_1177_)
    );

    and_bi _1889_ (
        .a(new_Jinkela_wire_7011),
        .b(_1177_),
        .c(_1178_)
    );

    and_bi _1890_ (
        .a(_1174_),
        .b(_1178_),
        .c(_1179_)
    );

    and_ii _1891_ (
        .a(new_Jinkela_wire_1944),
        .b(new_Jinkela_wire_6750),
        .c(_1180_)
    );

    and_bb _1892_ (
        .a(new_Jinkela_wire_1945),
        .b(new_Jinkela_wire_6751),
        .c(_1181_)
    );

    and_ii _1893_ (
        .a(_1181_),
        .b(_1180_),
        .c(_1182_)
    );

    or_bb _1894_ (
        .a(new_Jinkela_wire_196),
        .b(new_Jinkela_wire_55),
        .c(_1183_)
    );

    and_bi _1895_ (
        .a(new_Jinkela_wire_199),
        .b(new_Jinkela_wire_414),
        .c(_1184_)
    );

    and_bi _1896_ (
        .a(_1183_),
        .b(_1184_),
        .c(_1185_)
    );

    or_bb _1897_ (
        .a(_1185_),
        .b(new_Jinkela_wire_6353),
        .c(_1186_)
    );

    or_ii _1898_ (
        .a(new_Jinkela_wire_198),
        .b(new_Jinkela_wire_1202),
        .c(_1187_)
    );

    and_bi _1899_ (
        .a(new_Jinkela_wire_1547),
        .b(new_Jinkela_wire_206),
        .c(_1188_)
    );

    and_bi _1900_ (
        .a(_1187_),
        .b(_1188_),
        .c(_1189_)
    );

    and_bi _1901_ (
        .a(new_Jinkela_wire_6354),
        .b(_1189_),
        .c(_1190_)
    );

    and_bi _1902_ (
        .a(_1186_),
        .b(_1190_),
        .c(_1191_)
    );

    or_bb _1903_ (
        .a(new_Jinkela_wire_749),
        .b(new_Jinkela_wire_52),
        .c(_1192_)
    );

    and_bi _1904_ (
        .a(new_Jinkela_wire_747),
        .b(new_Jinkela_wire_419),
        .c(_1193_)
    );

    and_bi _1905_ (
        .a(_1192_),
        .b(_1193_),
        .c(_1194_)
    );

    or_bb _1906_ (
        .a(_1194_),
        .b(new_Jinkela_wire_6187),
        .c(_1195_)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(new_Jinkela_wire_230),
        .b(new_Jinkela_wire_231),
        .c(new_Jinkela_wire_232)
    );

    bfr new_Jinkela_buffer_5917 (
        .din(new_Jinkela_wire_7965),
        .dout(new_Jinkela_wire_7966)
    );

    bfr new_Jinkela_buffer_103 (
        .din(G12),
        .dout(new_Jinkela_wire_248)
    );

    bfr new_Jinkela_buffer_5902 (
        .din(new_Jinkela_wire_7944),
        .dout(new_Jinkela_wire_7945)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    bfr new_Jinkela_buffer_5921 (
        .din(_0314_),
        .dout(new_Jinkela_wire_7970)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_238),
        .dout(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    bfr new_Jinkela_buffer_5903 (
        .din(new_Jinkela_wire_7945),
        .dout(new_Jinkela_wire_7946)
    );

    bfr new_Jinkela_buffer_107 (
        .din(G88),
        .dout(new_Jinkela_wire_254)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    bfr new_Jinkela_buffer_5904 (
        .din(new_Jinkela_wire_7946),
        .dout(new_Jinkela_wire_7947)
    );

    bfr new_Jinkela_buffer_104 (
        .din(G42),
        .dout(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_5944 (
        .din(_0498_),
        .dout(new_Jinkela_wire_7993)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_5905 (
        .din(new_Jinkela_wire_7947),
        .dout(new_Jinkela_wire_7948)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    bfr new_Jinkela_buffer_5922 (
        .din(new_Jinkela_wire_7970),
        .dout(new_Jinkela_wire_7971)
    );

    spl2 new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_240),
        .b(new_Jinkela_wire_241),
        .c(new_Jinkela_wire_242)
    );

    bfr new_Jinkela_buffer_5918 (
        .din(new_Jinkela_wire_7966),
        .dout(new_Jinkela_wire_7967)
    );

    bfr new_Jinkela_buffer_5906 (
        .din(new_Jinkela_wire_7948),
        .dout(new_Jinkela_wire_7949)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_244),
        .dout(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_5907 (
        .din(new_Jinkela_wire_7949),
        .dout(new_Jinkela_wire_7950)
    );

    bfr new_Jinkela_buffer_5946 (
        .din(_0826_),
        .dout(new_Jinkela_wire_7995)
    );

    spl2 new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_245),
        .b(new_Jinkela_wire_246),
        .c(new_Jinkela_wire_247)
    );

    bfr new_Jinkela_buffer_5919 (
        .din(new_Jinkela_wire_7967),
        .dout(new_Jinkela_wire_7968)
    );

    bfr new_Jinkela_buffer_5908 (
        .din(new_Jinkela_wire_7950),
        .dout(new_Jinkela_wire_7951)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    bfr new_Jinkela_buffer_5909 (
        .din(new_Jinkela_wire_7951),
        .dout(new_Jinkela_wire_7952)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    bfr new_Jinkela_buffer_5923 (
        .din(new_Jinkela_wire_7971),
        .dout(new_Jinkela_wire_7972)
    );

    spl3L new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_255),
        .d(new_Jinkela_wire_256),
        .b(new_Jinkela_wire_257),
        .c(new_Jinkela_wire_258)
    );

    bfr new_Jinkela_buffer_5920 (
        .din(new_Jinkela_wire_7968),
        .dout(new_Jinkela_wire_7969)
    );

    bfr new_Jinkela_buffer_5910 (
        .din(new_Jinkela_wire_7952),
        .dout(new_Jinkela_wire_7953)
    );

    spl2 new_Jinkela_splitter_48 (
        .a(new_Jinkela_wire_251),
        .b(new_Jinkela_wire_252),
        .c(new_Jinkela_wire_253)
    );

    spl2 new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_254),
        .b(new_Jinkela_wire_255),
        .c(new_Jinkela_wire_259)
    );

    bfr new_Jinkela_buffer_5911 (
        .din(new_Jinkela_wire_7953),
        .dout(new_Jinkela_wire_7954)
    );

    bfr new_Jinkela_buffer_113 (
        .din(G8),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_5945 (
        .din(new_Jinkela_wire_7993),
        .dout(new_Jinkela_wire_7994)
    );

    spl4L new_Jinkela_splitter_51 (
        .a(new_Jinkela_wire_259),
        .d(new_Jinkela_wire_260),
        .e(new_Jinkela_wire_261),
        .b(new_Jinkela_wire_262),
        .c(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_5912 (
        .din(new_Jinkela_wire_7954),
        .dout(new_Jinkela_wire_7955)
    );

    bfr new_Jinkela_buffer_108 (
        .din(G57),
        .dout(new_Jinkela_wire_264)
    );

    spl2 new_Jinkela_splitter_52 (
        .a(G137),
        .b(new_Jinkela_wire_271),
        .c(new_Jinkela_wire_272)
    );

    bfr new_Jinkela_buffer_5924 (
        .din(new_Jinkela_wire_7972),
        .dout(new_Jinkela_wire_7973)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    bfr new_Jinkela_buffer_5913 (
        .din(new_Jinkela_wire_7955),
        .dout(new_Jinkela_wire_7956)
    );

    spl4L new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_282),
        .d(new_Jinkela_wire_283),
        .e(new_Jinkela_wire_284),
        .b(new_Jinkela_wire_286),
        .c(new_Jinkela_wire_291)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    bfr new_Jinkela_buffer_5947 (
        .din(_1052_),
        .dout(new_Jinkela_wire_7996)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_266),
        .dout(new_Jinkela_wire_267)
    );

    bfr new_Jinkela_buffer_5914 (
        .din(new_Jinkela_wire_7956),
        .dout(new_Jinkela_wire_7957)
    );

    bfr new_Jinkela_buffer_5925 (
        .din(new_Jinkela_wire_7973),
        .dout(new_Jinkela_wire_7974)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_267),
        .dout(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_5951 (
        .din(new_net_2385),
        .dout(new_Jinkela_wire_8000)
    );

    bfr new_Jinkela_buffer_5926 (
        .din(new_Jinkela_wire_7974),
        .dout(new_Jinkela_wire_7975)
    );

    bfr new_Jinkela_buffer_5948 (
        .din(new_Jinkela_wire_7996),
        .dout(new_Jinkela_wire_7997)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_5927 (
        .din(new_Jinkela_wire_7975),
        .dout(new_Jinkela_wire_7976)
    );

    spl2 new_Jinkela_splitter_55 (
        .a(G128),
        .b(new_Jinkela_wire_280),
        .c(new_Jinkela_wire_282)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(G54),
        .b(new_Jinkela_wire_299),
        .c(new_Jinkela_wire_300)
    );

    bfr new_Jinkela_buffer_5928 (
        .din(new_Jinkela_wire_7976),
        .dout(new_Jinkela_wire_7977)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_273),
        .dout(new_Jinkela_wire_274)
    );

    bfr new_Jinkela_buffer_5949 (
        .din(new_Jinkela_wire_7997),
        .dout(new_Jinkela_wire_7998)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_274),
        .dout(new_Jinkela_wire_275)
    );

    bfr new_Jinkela_buffer_5929 (
        .din(new_Jinkela_wire_7977),
        .dout(new_Jinkela_wire_7978)
    );

    bfr new_Jinkela_buffer_5952 (
        .din(new_Jinkela_wire_8000),
        .dout(new_Jinkela_wire_8001)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_275),
        .b(new_Jinkela_wire_276),
        .c(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_5930 (
        .din(new_Jinkela_wire_7978),
        .dout(new_Jinkela_wire_7979)
    );

    spl2 new_Jinkela_splitter_54 (
        .a(new_Jinkela_wire_277),
        .b(new_Jinkela_wire_278),
        .c(new_Jinkela_wire_279)
    );

    bfr new_Jinkela_buffer_5950 (
        .din(new_Jinkela_wire_7998),
        .dout(new_Jinkela_wire_7999)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(G153),
        .b(new_Jinkela_wire_297),
        .c(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_5931 (
        .din(new_Jinkela_wire_7979),
        .dout(new_Jinkela_wire_7980)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_280),
        .dout(new_Jinkela_wire_281)
    );

    spl4L new_Jinkela_splitter_57 (
        .a(new_Jinkela_wire_286),
        .d(new_Jinkela_wire_287),
        .e(new_Jinkela_wire_288),
        .b(new_Jinkela_wire_289),
        .c(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_5932 (
        .din(new_Jinkela_wire_7980),
        .dout(new_Jinkela_wire_7981)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_291),
        .d(new_Jinkela_wire_292),
        .e(new_Jinkela_wire_293),
        .b(new_Jinkela_wire_294),
        .c(new_Jinkela_wire_295)
    );

    bfr new_Jinkela_buffer_125 (
        .din(G118),
        .dout(new_Jinkela_wire_305)
    );

    bfr new_Jinkela_buffer_5953 (
        .din(new_Jinkela_wire_8001),
        .dout(new_Jinkela_wire_8002)
    );

    bfr new_Jinkela_buffer_1706 (
        .din(new_Jinkela_wire_2717),
        .dout(new_Jinkela_wire_2718)
    );

    spl4L new_Jinkela_splitter_655 (
        .a(new_Jinkela_wire_6350),
        .d(new_Jinkela_wire_6351),
        .e(new_Jinkela_wire_6352),
        .b(new_Jinkela_wire_6353),
        .c(new_Jinkela_wire_6354)
    );

    bfr new_Jinkela_buffer_4602 (
        .din(new_Jinkela_wire_6298),
        .dout(new_Jinkela_wire_6299)
    );

    bfr new_Jinkela_buffer_1759 (
        .din(new_Jinkela_wire_2785),
        .dout(new_Jinkela_wire_2786)
    );

    bfr new_Jinkela_buffer_1707 (
        .din(new_Jinkela_wire_2718),
        .dout(new_Jinkela_wire_2719)
    );

    bfr new_Jinkela_buffer_4628 (
        .din(new_Jinkela_wire_6332),
        .dout(new_Jinkela_wire_6333)
    );

    bfr new_Jinkela_buffer_1730 (
        .din(new_Jinkela_wire_2741),
        .dout(new_Jinkela_wire_2742)
    );

    bfr new_Jinkela_buffer_4603 (
        .din(new_Jinkela_wire_6299),
        .dout(new_Jinkela_wire_6300)
    );

    bfr new_Jinkela_buffer_1708 (
        .din(new_Jinkela_wire_2719),
        .dout(new_Jinkela_wire_2720)
    );

    bfr new_Jinkela_buffer_4646 (
        .din(new_Jinkela_wire_6358),
        .dout(new_Jinkela_wire_6359)
    );

    bfr new_Jinkela_buffer_4604 (
        .din(new_Jinkela_wire_6300),
        .dout(new_Jinkela_wire_6301)
    );

    spl3L new_Jinkela_splitter_384 (
        .a(new_Jinkela_wire_2806),
        .d(new_Jinkela_wire_2807),
        .b(new_Jinkela_wire_2808),
        .c(new_Jinkela_wire_2809)
    );

    bfr new_Jinkela_buffer_1709 (
        .din(new_Jinkela_wire_2720),
        .dout(new_Jinkela_wire_2721)
    );

    bfr new_Jinkela_buffer_4629 (
        .din(new_Jinkela_wire_6333),
        .dout(new_Jinkela_wire_6334)
    );

    bfr new_Jinkela_buffer_1731 (
        .din(new_Jinkela_wire_2742),
        .dout(new_Jinkela_wire_2743)
    );

    bfr new_Jinkela_buffer_4605 (
        .din(new_Jinkela_wire_6301),
        .dout(new_Jinkela_wire_6302)
    );

    bfr new_Jinkela_buffer_1710 (
        .din(new_Jinkela_wire_2721),
        .dout(new_Jinkela_wire_2722)
    );

    bfr new_Jinkela_buffer_4652 (
        .din(_0438_),
        .dout(new_Jinkela_wire_6365)
    );

    bfr new_Jinkela_buffer_1807 (
        .din(new_Jinkela_wire_2842),
        .dout(new_Jinkela_wire_2843)
    );

    bfr new_Jinkela_buffer_4606 (
        .din(new_Jinkela_wire_6302),
        .dout(new_Jinkela_wire_6303)
    );

    bfr new_Jinkela_buffer_1760 (
        .din(new_Jinkela_wire_2786),
        .dout(new_Jinkela_wire_2787)
    );

    bfr new_Jinkela_buffer_1711 (
        .din(new_Jinkela_wire_2722),
        .dout(new_Jinkela_wire_2723)
    );

    bfr new_Jinkela_buffer_4630 (
        .din(new_Jinkela_wire_6334),
        .dout(new_Jinkela_wire_6335)
    );

    bfr new_Jinkela_buffer_1732 (
        .din(new_Jinkela_wire_2743),
        .dout(new_Jinkela_wire_2744)
    );

    bfr new_Jinkela_buffer_4607 (
        .din(new_Jinkela_wire_6303),
        .dout(new_Jinkela_wire_6304)
    );

    bfr new_Jinkela_buffer_1712 (
        .din(new_Jinkela_wire_2723),
        .dout(new_Jinkela_wire_2724)
    );

    bfr new_Jinkela_buffer_4608 (
        .din(new_Jinkela_wire_6304),
        .dout(new_Jinkela_wire_6305)
    );

    bfr new_Jinkela_buffer_1733 (
        .din(new_Jinkela_wire_2744),
        .dout(new_Jinkela_wire_2745)
    );

    bfr new_Jinkela_buffer_4631 (
        .din(new_Jinkela_wire_6335),
        .dout(new_Jinkela_wire_6336)
    );

    bfr new_Jinkela_buffer_1780 (
        .din(new_Jinkela_wire_2809),
        .dout(new_Jinkela_wire_2810)
    );

    bfr new_Jinkela_buffer_4609 (
        .din(new_Jinkela_wire_6305),
        .dout(new_Jinkela_wire_6306)
    );

    bfr new_Jinkela_buffer_1761 (
        .din(new_Jinkela_wire_2787),
        .dout(new_Jinkela_wire_2788)
    );

    bfr new_Jinkela_buffer_1734 (
        .din(new_Jinkela_wire_2745),
        .dout(new_Jinkela_wire_2746)
    );

    bfr new_Jinkela_buffer_4651 (
        .din(new_Jinkela_wire_6363),
        .dout(new_Jinkela_wire_6364)
    );

    bfr new_Jinkela_buffer_4647 (
        .din(new_Jinkela_wire_6359),
        .dout(new_Jinkela_wire_6360)
    );

    bfr new_Jinkela_buffer_4610 (
        .din(new_Jinkela_wire_6306),
        .dout(new_Jinkela_wire_6307)
    );

    bfr new_Jinkela_buffer_1735 (
        .din(new_Jinkela_wire_2746),
        .dout(new_Jinkela_wire_2747)
    );

    bfr new_Jinkela_buffer_4632 (
        .din(new_Jinkela_wire_6336),
        .dout(new_Jinkela_wire_6337)
    );

    bfr new_Jinkela_buffer_4611 (
        .din(new_Jinkela_wire_6307),
        .dout(new_Jinkela_wire_6308)
    );

    bfr new_Jinkela_buffer_1762 (
        .din(new_Jinkela_wire_2788),
        .dout(new_Jinkela_wire_2789)
    );

    bfr new_Jinkela_buffer_1736 (
        .din(new_Jinkela_wire_2747),
        .dout(new_Jinkela_wire_2748)
    );

    bfr new_Jinkela_buffer_4612 (
        .din(new_Jinkela_wire_6308),
        .dout(new_Jinkela_wire_6309)
    );

    bfr new_Jinkela_buffer_1786 (
        .din(new_Jinkela_wire_2819),
        .dout(new_Jinkela_wire_2820)
    );

    bfr new_Jinkela_buffer_1737 (
        .din(new_Jinkela_wire_2748),
        .dout(new_Jinkela_wire_2749)
    );

    bfr new_Jinkela_buffer_4633 (
        .din(new_Jinkela_wire_6337),
        .dout(new_Jinkela_wire_6338)
    );

    bfr new_Jinkela_buffer_4613 (
        .din(new_Jinkela_wire_6309),
        .dout(new_Jinkela_wire_6310)
    );

    bfr new_Jinkela_buffer_1763 (
        .din(new_Jinkela_wire_2789),
        .dout(new_Jinkela_wire_2790)
    );

    bfr new_Jinkela_buffer_1738 (
        .din(new_Jinkela_wire_2749),
        .dout(new_Jinkela_wire_2750)
    );

    bfr new_Jinkela_buffer_4662 (
        .din(_0281_),
        .dout(new_Jinkela_wire_6375)
    );

    bfr new_Jinkela_buffer_4648 (
        .din(new_Jinkela_wire_6360),
        .dout(new_Jinkela_wire_6361)
    );

    bfr new_Jinkela_buffer_4614 (
        .din(new_Jinkela_wire_6310),
        .dout(new_Jinkela_wire_6311)
    );

    bfr new_Jinkela_buffer_1781 (
        .din(new_Jinkela_wire_2810),
        .dout(new_Jinkela_wire_2811)
    );

    bfr new_Jinkela_buffer_1739 (
        .din(new_Jinkela_wire_2750),
        .dout(new_Jinkela_wire_2751)
    );

    bfr new_Jinkela_buffer_4634 (
        .din(new_Jinkela_wire_6338),
        .dout(new_Jinkela_wire_6339)
    );

    bfr new_Jinkela_buffer_4615 (
        .din(new_Jinkela_wire_6311),
        .dout(new_Jinkela_wire_6312)
    );

    bfr new_Jinkela_buffer_1764 (
        .din(new_Jinkela_wire_2790),
        .dout(new_Jinkela_wire_2791)
    );

    bfr new_Jinkela_buffer_1740 (
        .din(new_Jinkela_wire_2751),
        .dout(new_Jinkela_wire_2752)
    );

    bfr new_Jinkela_buffer_4616 (
        .din(new_Jinkela_wire_6312),
        .dout(new_Jinkela_wire_6313)
    );

    bfr new_Jinkela_buffer_1741 (
        .din(new_Jinkela_wire_2752),
        .dout(new_Jinkela_wire_2753)
    );

    bfr new_Jinkela_buffer_4635 (
        .din(new_Jinkela_wire_6339),
        .dout(new_Jinkela_wire_6340)
    );

    bfr new_Jinkela_buffer_1787 (
        .din(new_Jinkela_wire_2820),
        .dout(new_Jinkela_wire_2821)
    );

    bfr new_Jinkela_buffer_4617 (
        .din(new_Jinkela_wire_6313),
        .dout(new_Jinkela_wire_6314)
    );

    bfr new_Jinkela_buffer_1765 (
        .din(new_Jinkela_wire_2791),
        .dout(new_Jinkela_wire_2792)
    );

    bfr new_Jinkela_buffer_1742 (
        .din(new_Jinkela_wire_2753),
        .dout(new_Jinkela_wire_2754)
    );

    bfr new_Jinkela_buffer_4653 (
        .din(new_Jinkela_wire_6365),
        .dout(new_Jinkela_wire_6366)
    );

    bfr new_Jinkela_buffer_4649 (
        .din(new_Jinkela_wire_6361),
        .dout(new_Jinkela_wire_6362)
    );

    bfr new_Jinkela_buffer_4618 (
        .din(new_Jinkela_wire_6314),
        .dout(new_Jinkela_wire_6315)
    );

    bfr new_Jinkela_buffer_1782 (
        .din(new_Jinkela_wire_2811),
        .dout(new_Jinkela_wire_2812)
    );

    bfr new_Jinkela_buffer_1743 (
        .din(new_Jinkela_wire_2754),
        .dout(new_Jinkela_wire_2755)
    );

    bfr new_Jinkela_buffer_4636 (
        .din(new_Jinkela_wire_6340),
        .dout(new_Jinkela_wire_6341)
    );

    bfr new_Jinkela_buffer_4619 (
        .din(new_Jinkela_wire_6315),
        .dout(new_Jinkela_wire_6316)
    );

    bfr new_Jinkela_buffer_1766 (
        .din(new_Jinkela_wire_2792),
        .dout(new_Jinkela_wire_2793)
    );

    bfr new_Jinkela_buffer_1744 (
        .din(new_Jinkela_wire_2755),
        .dout(new_Jinkela_wire_2756)
    );

    bfr new_Jinkela_buffer_4637 (
        .din(new_Jinkela_wire_6341),
        .dout(new_Jinkela_wire_6342)
    );

    bfr new_Jinkela_buffer_1745 (
        .din(new_Jinkela_wire_2756),
        .dout(new_Jinkela_wire_2757)
    );

    spl2 new_Jinkela_splitter_657 (
        .a(_0630_),
        .b(new_Jinkela_wire_6376),
        .c(new_Jinkela_wire_6377)
    );

    spl3L new_Jinkela_splitter_658 (
        .a(_0948_),
        .d(new_Jinkela_wire_6379),
        .b(new_Jinkela_wire_6380),
        .c(new_Jinkela_wire_6381)
    );

    bfr new_Jinkela_buffer_1815 (
        .din(_0937_),
        .dout(new_Jinkela_wire_2854)
    );

    bfr new_Jinkela_buffer_4638 (
        .din(new_Jinkela_wire_6342),
        .dout(new_Jinkela_wire_6343)
    );

    bfr new_Jinkela_buffer_1767 (
        .din(new_Jinkela_wire_2793),
        .dout(new_Jinkela_wire_2794)
    );

    bfr new_Jinkela_buffer_1746 (
        .din(new_Jinkela_wire_2757),
        .dout(new_Jinkela_wire_2758)
    );

    bfr new_Jinkela_buffer_4654 (
        .din(new_Jinkela_wire_6366),
        .dout(new_Jinkela_wire_6367)
    );

    bfr new_Jinkela_buffer_4639 (
        .din(new_Jinkela_wire_6343),
        .dout(new_Jinkela_wire_6344)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(new_Jinkela_wire_2014),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_5307 (
        .din(new_Jinkela_wire_7229),
        .dout(new_Jinkela_wire_7230)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_2041),
        .dout(new_Jinkela_wire_2042)
    );

    bfr new_Jinkela_buffer_5341 (
        .din(new_Jinkela_wire_7267),
        .dout(new_Jinkela_wire_7268)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(new_Jinkela_wire_2015),
        .dout(new_Jinkela_wire_2016)
    );

    bfr new_Jinkela_buffer_5308 (
        .din(new_Jinkela_wire_7230),
        .dout(new_Jinkela_wire_7231)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(new_Jinkela_wire_2071),
        .dout(new_Jinkela_wire_2072)
    );

    bfr new_Jinkela_buffer_5325 (
        .din(new_Jinkela_wire_7251),
        .dout(new_Jinkela_wire_7252)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(new_Jinkela_wire_2016),
        .dout(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_5309 (
        .din(new_Jinkela_wire_7231),
        .dout(new_Jinkela_wire_7232)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_2042),
        .dout(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_5419 (
        .din(_0356_),
        .dout(new_Jinkela_wire_7352)
    );

    bfr new_Jinkela_buffer_5362 (
        .din(new_Jinkela_wire_7289),
        .dout(new_Jinkela_wire_7290)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_2017),
        .dout(new_Jinkela_wire_2018)
    );

    bfr new_Jinkela_buffer_5310 (
        .din(new_Jinkela_wire_7232),
        .dout(new_Jinkela_wire_7233)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(_0419_),
        .dout(new_Jinkela_wire_2095)
    );

    bfr new_Jinkela_buffer_5326 (
        .din(new_Jinkela_wire_7252),
        .dout(new_Jinkela_wire_7253)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_2088),
        .dout(new_Jinkela_wire_2089)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_2018),
        .dout(new_Jinkela_wire_2019)
    );

    bfr new_Jinkela_buffer_5311 (
        .din(new_Jinkela_wire_7233),
        .dout(new_Jinkela_wire_7234)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    bfr new_Jinkela_buffer_5342 (
        .din(new_Jinkela_wire_7268),
        .dout(new_Jinkela_wire_7269)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(new_Jinkela_wire_2019),
        .dout(new_Jinkela_wire_2020)
    );

    bfr new_Jinkela_buffer_5312 (
        .din(new_Jinkela_wire_7234),
        .dout(new_Jinkela_wire_7235)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_Jinkela_wire_2072),
        .dout(new_Jinkela_wire_2073)
    );

    bfr new_Jinkela_buffer_5327 (
        .din(new_Jinkela_wire_7253),
        .dout(new_Jinkela_wire_7254)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(new_Jinkela_wire_2020),
        .dout(new_Jinkela_wire_2021)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_2044),
        .dout(new_Jinkela_wire_2045)
    );

    bfr new_Jinkela_buffer_5328 (
        .din(new_Jinkela_wire_7254),
        .dout(new_Jinkela_wire_7255)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_2021),
        .dout(new_Jinkela_wire_2022)
    );

    bfr new_Jinkela_buffer_5343 (
        .din(new_Jinkela_wire_7269),
        .dout(new_Jinkela_wire_7270)
    );

    bfr new_Jinkela_buffer_5329 (
        .din(new_Jinkela_wire_7255),
        .dout(new_Jinkela_wire_7256)
    );

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    spl4L new_Jinkela_splitter_744 (
        .a(new_Jinkela_wire_7291),
        .d(new_Jinkela_wire_7292),
        .e(new_Jinkela_wire_7293),
        .b(new_Jinkela_wire_7294),
        .c(new_Jinkela_wire_7295)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_5330 (
        .din(new_Jinkela_wire_7256),
        .dout(new_Jinkela_wire_7257)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(new_Jinkela_wire_2023),
        .dout(new_Jinkela_wire_2024)
    );

    bfr new_Jinkela_buffer_5344 (
        .din(new_Jinkela_wire_7270),
        .dout(new_Jinkela_wire_7271)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(new_Jinkela_wire_2073),
        .dout(new_Jinkela_wire_2074)
    );

    bfr new_Jinkela_buffer_5331 (
        .din(new_Jinkela_wire_7257),
        .dout(new_Jinkela_wire_7258)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_2024),
        .dout(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_5363 (
        .din(new_Jinkela_wire_7295),
        .dout(new_Jinkela_wire_7296)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_2046),
        .dout(new_Jinkela_wire_2047)
    );

    bfr new_Jinkela_buffer_5332 (
        .din(new_Jinkela_wire_7258),
        .dout(new_Jinkela_wire_7259)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_2025),
        .dout(new_Jinkela_wire_2026)
    );

    bfr new_Jinkela_buffer_5345 (
        .din(new_Jinkela_wire_7271),
        .dout(new_Jinkela_wire_7272)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(_1062_),
        .dout(new_Jinkela_wire_2093)
    );

    bfr new_Jinkela_buffer_5333 (
        .din(new_Jinkela_wire_7259),
        .dout(new_Jinkela_wire_7260)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_5383 (
        .din(new_Jinkela_wire_7315),
        .dout(new_Jinkela_wire_7316)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(new_Jinkela_wire_2047),
        .dout(new_Jinkela_wire_2048)
    );

    bfr new_Jinkela_buffer_5334 (
        .din(new_Jinkela_wire_7260),
        .dout(new_Jinkela_wire_7261)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_2027),
        .dout(new_Jinkela_wire_2028)
    );

    bfr new_Jinkela_buffer_5346 (
        .din(new_Jinkela_wire_7272),
        .dout(new_Jinkela_wire_7273)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(new_Jinkela_wire_2074),
        .dout(new_Jinkela_wire_2075)
    );

    bfr new_Jinkela_buffer_5335 (
        .din(new_Jinkela_wire_7261),
        .dout(new_Jinkela_wire_7262)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_2028),
        .dout(new_Jinkela_wire_2029)
    );

    bfr new_Jinkela_buffer_5438 (
        .din(_0908_),
        .dout(new_Jinkela_wire_7371)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(new_Jinkela_wire_2048),
        .dout(new_Jinkela_wire_2049)
    );

    bfr new_Jinkela_buffer_5336 (
        .din(new_Jinkela_wire_7262),
        .dout(new_Jinkela_wire_7263)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_2029),
        .dout(new_Jinkela_wire_2030)
    );

    bfr new_Jinkela_buffer_5347 (
        .din(new_Jinkela_wire_7273),
        .dout(new_Jinkela_wire_7274)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_2093),
        .dout(new_Jinkela_wire_2094)
    );

    bfr new_Jinkela_buffer_5337 (
        .din(new_Jinkela_wire_7263),
        .dout(new_Jinkela_wire_7264)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_2030),
        .dout(new_Jinkela_wire_2031)
    );

    bfr new_Jinkela_buffer_5364 (
        .din(new_Jinkela_wire_7296),
        .dout(new_Jinkela_wire_7297)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(new_Jinkela_wire_2049),
        .dout(new_Jinkela_wire_2050)
    );

    bfr new_Jinkela_buffer_5338 (
        .din(new_Jinkela_wire_7264),
        .dout(new_Jinkela_wire_7265)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_2031),
        .dout(new_Jinkela_wire_2032)
    );

    bfr new_Jinkela_buffer_5348 (
        .din(new_Jinkela_wire_7274),
        .dout(new_Jinkela_wire_7275)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_2075),
        .dout(new_Jinkela_wire_2076)
    );

    bfr new_Jinkela_buffer_5384 (
        .din(new_Jinkela_wire_7316),
        .dout(new_Jinkela_wire_7317)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_2032),
        .dout(new_Jinkela_wire_2033)
    );

    bfr new_Jinkela_buffer_5349 (
        .din(new_Jinkela_wire_7275),
        .dout(new_Jinkela_wire_7276)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_Jinkela_wire_2050),
        .dout(new_Jinkela_wire_2051)
    );

    bfr new_Jinkela_buffer_5365 (
        .din(new_Jinkela_wire_7297),
        .dout(new_Jinkela_wire_7298)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(_0506_),
        .dout(new_Jinkela_wire_2118)
    );

    bfr new_Jinkela_buffer_5350 (
        .din(new_Jinkela_wire_7276),
        .dout(new_Jinkela_wire_7277)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_2051),
        .dout(new_Jinkela_wire_2052)
    );

    bfr new_Jinkela_buffer_5420 (
        .din(new_Jinkela_wire_7352),
        .dout(new_Jinkela_wire_7353)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_2076),
        .dout(new_Jinkela_wire_2077)
    );

    bfr new_Jinkela_buffer_5351 (
        .din(new_Jinkela_wire_7277),
        .dout(new_Jinkela_wire_7278)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_2052),
        .dout(new_Jinkela_wire_2053)
    );

    bfr new_Jinkela_buffer_5366 (
        .din(new_Jinkela_wire_7298),
        .dout(new_Jinkela_wire_7299)
    );

    bfr new_Jinkela_buffer_3250 (
        .din(new_Jinkela_wire_4634),
        .dout(new_Jinkela_wire_4635)
    );

    bfr new_Jinkela_buffer_3321 (
        .din(new_Jinkela_wire_4710),
        .dout(new_Jinkela_wire_4711)
    );

    bfr new_Jinkela_buffer_3251 (
        .din(new_Jinkela_wire_4635),
        .dout(new_Jinkela_wire_4636)
    );

    bfr new_Jinkela_buffer_3285 (
        .din(new_Jinkela_wire_4671),
        .dout(new_Jinkela_wire_4672)
    );

    bfr new_Jinkela_buffer_3252 (
        .din(new_Jinkela_wire_4636),
        .dout(new_Jinkela_wire_4637)
    );

    bfr new_Jinkela_buffer_3253 (
        .din(new_Jinkela_wire_4637),
        .dout(new_Jinkela_wire_4638)
    );

    bfr new_Jinkela_buffer_3286 (
        .din(new_Jinkela_wire_4672),
        .dout(new_Jinkela_wire_4673)
    );

    bfr new_Jinkela_buffer_3254 (
        .din(new_Jinkela_wire_4638),
        .dout(new_Jinkela_wire_4639)
    );

    bfr new_Jinkela_buffer_3363 (
        .din(_0064_),
        .dout(new_Jinkela_wire_4755)
    );

    bfr new_Jinkela_buffer_3255 (
        .din(new_Jinkela_wire_4639),
        .dout(new_Jinkela_wire_4640)
    );

    bfr new_Jinkela_buffer_3364 (
        .din(_0656_),
        .dout(new_Jinkela_wire_4758)
    );

    bfr new_Jinkela_buffer_3287 (
        .din(new_Jinkela_wire_4673),
        .dout(new_Jinkela_wire_4674)
    );

    bfr new_Jinkela_buffer_3256 (
        .din(new_Jinkela_wire_4640),
        .dout(new_Jinkela_wire_4641)
    );

    bfr new_Jinkela_buffer_3324 (
        .din(new_Jinkela_wire_4715),
        .dout(new_Jinkela_wire_4716)
    );

    bfr new_Jinkela_buffer_3257 (
        .din(new_Jinkela_wire_4641),
        .dout(new_Jinkela_wire_4642)
    );

    bfr new_Jinkela_buffer_3288 (
        .din(new_Jinkela_wire_4674),
        .dout(new_Jinkela_wire_4675)
    );

    bfr new_Jinkela_buffer_3258 (
        .din(new_Jinkela_wire_4642),
        .dout(new_Jinkela_wire_4643)
    );

    bfr new_Jinkela_buffer_3369 (
        .din(new_net_2361),
        .dout(new_Jinkela_wire_4763)
    );

    bfr new_Jinkela_buffer_3259 (
        .din(new_Jinkela_wire_4643),
        .dout(new_Jinkela_wire_4644)
    );

    bfr new_Jinkela_buffer_3289 (
        .din(new_Jinkela_wire_4675),
        .dout(new_Jinkela_wire_4676)
    );

    bfr new_Jinkela_buffer_3260 (
        .din(new_Jinkela_wire_4644),
        .dout(new_Jinkela_wire_4645)
    );

    bfr new_Jinkela_buffer_3325 (
        .din(new_Jinkela_wire_4716),
        .dout(new_Jinkela_wire_4717)
    );

    bfr new_Jinkela_buffer_3261 (
        .din(new_Jinkela_wire_4645),
        .dout(new_Jinkela_wire_4646)
    );

    bfr new_Jinkela_buffer_3290 (
        .din(new_Jinkela_wire_4676),
        .dout(new_Jinkela_wire_4677)
    );

    bfr new_Jinkela_buffer_3262 (
        .din(new_Jinkela_wire_4646),
        .dout(new_Jinkela_wire_4647)
    );

    spl2 new_Jinkela_splitter_530 (
        .a(new_Jinkela_wire_4755),
        .b(new_Jinkela_wire_4756),
        .c(new_Jinkela_wire_4757)
    );

    bfr new_Jinkela_buffer_3263 (
        .din(new_Jinkela_wire_4647),
        .dout(new_Jinkela_wire_4648)
    );

    bfr new_Jinkela_buffer_3291 (
        .din(new_Jinkela_wire_4677),
        .dout(new_Jinkela_wire_4678)
    );

    bfr new_Jinkela_buffer_3264 (
        .din(new_Jinkela_wire_4648),
        .dout(new_Jinkela_wire_4649)
    );

    bfr new_Jinkela_buffer_3326 (
        .din(new_Jinkela_wire_4717),
        .dout(new_Jinkela_wire_4718)
    );

    bfr new_Jinkela_buffer_3265 (
        .din(new_Jinkela_wire_4649),
        .dout(new_Jinkela_wire_4650)
    );

    bfr new_Jinkela_buffer_3292 (
        .din(new_Jinkela_wire_4678),
        .dout(new_Jinkela_wire_4679)
    );

    bfr new_Jinkela_buffer_3266 (
        .din(new_Jinkela_wire_4650),
        .dout(new_Jinkela_wire_4651)
    );

    bfr new_Jinkela_buffer_3267 (
        .din(new_Jinkela_wire_4651),
        .dout(new_Jinkela_wire_4652)
    );

    bfr new_Jinkela_buffer_3365 (
        .din(new_Jinkela_wire_4758),
        .dout(new_Jinkela_wire_4759)
    );

    bfr new_Jinkela_buffer_3293 (
        .din(new_Jinkela_wire_4679),
        .dout(new_Jinkela_wire_4680)
    );

    bfr new_Jinkela_buffer_3268 (
        .din(new_Jinkela_wire_4652),
        .dout(new_Jinkela_wire_4653)
    );

    bfr new_Jinkela_buffer_3327 (
        .din(new_Jinkela_wire_4718),
        .dout(new_Jinkela_wire_4719)
    );

    spl2 new_Jinkela_splitter_527 (
        .a(new_Jinkela_wire_4653),
        .b(new_Jinkela_wire_4654),
        .c(new_Jinkela_wire_4655)
    );

    bfr new_Jinkela_buffer_3294 (
        .din(new_Jinkela_wire_4680),
        .dout(new_Jinkela_wire_4681)
    );

    bfr new_Jinkela_buffer_3295 (
        .din(new_Jinkela_wire_4681),
        .dout(new_Jinkela_wire_4682)
    );

    or_ii _1907_ (
        .a(new_Jinkela_wire_755),
        .b(new_Jinkela_wire_1213),
        .c(_1196_)
    );

    bfr new_Jinkela_buffer_4571 (
        .din(new_Jinkela_wire_6263),
        .dout(new_Jinkela_wire_6264)
    );

    bfr new_Jinkela_buffer_5933 (
        .din(new_Jinkela_wire_7981),
        .dout(new_Jinkela_wire_7982)
    );

    and_bi _1908_ (
        .a(new_Jinkela_wire_1541),
        .b(new_Jinkela_wire_745),
        .c(_1197_)
    );

    bfr new_Jinkela_buffer_4589 (
        .din(new_Jinkela_wire_6285),
        .dout(new_Jinkela_wire_6286)
    );

    and_bi _1909_ (
        .a(_1196_),
        .b(_1197_),
        .c(_1198_)
    );

    bfr new_Jinkela_buffer_4572 (
        .din(new_Jinkela_wire_6264),
        .dout(new_Jinkela_wire_6265)
    );

    bfr new_Jinkela_buffer_5934 (
        .din(new_Jinkela_wire_7982),
        .dout(new_Jinkela_wire_7983)
    );

    and_bi _1910_ (
        .a(new_Jinkela_wire_6189),
        .b(_1198_),
        .c(_1199_)
    );

    bfr new_Jinkela_buffer_5954 (
        .din(new_Jinkela_wire_8002),
        .dout(new_Jinkela_wire_8003)
    );

    spl4L new_Jinkela_splitter_656 (
        .a(_0613_),
        .d(new_Jinkela_wire_6355),
        .e(new_Jinkela_wire_6356),
        .b(new_Jinkela_wire_6357),
        .c(new_Jinkela_wire_6358)
    );

    and_bi _1911_ (
        .a(_1195_),
        .b(_1199_),
        .c(_1200_)
    );

    bfr new_Jinkela_buffer_4573 (
        .din(new_Jinkela_wire_6265),
        .dout(new_Jinkela_wire_6266)
    );

    bfr new_Jinkela_buffer_5935 (
        .din(new_Jinkela_wire_7983),
        .dout(new_Jinkela_wire_7984)
    );

    or_bb _1912_ (
        .a(new_Jinkela_wire_448),
        .b(new_Jinkela_wire_60),
        .c(_1201_)
    );

    bfr new_Jinkela_buffer_4590 (
        .din(new_Jinkela_wire_6286),
        .dout(new_Jinkela_wire_6287)
    );

    and_bi _1913_ (
        .a(new_Jinkela_wire_440),
        .b(new_Jinkela_wire_408),
        .c(_1202_)
    );

    bfr new_Jinkela_buffer_4574 (
        .din(new_Jinkela_wire_6266),
        .dout(new_Jinkela_wire_6267)
    );

    bfr new_Jinkela_buffer_5936 (
        .din(new_Jinkela_wire_7984),
        .dout(new_Jinkela_wire_7985)
    );

    and_bi _1914_ (
        .a(_1201_),
        .b(_1202_),
        .c(_1203_)
    );

    bfr new_Jinkela_buffer_5955 (
        .din(new_Jinkela_wire_8003),
        .dout(new_Jinkela_wire_8004)
    );

    bfr new_Jinkela_buffer_4644 (
        .din(_0778_),
        .dout(new_Jinkela_wire_6349)
    );

    and_bi _1915_ (
        .a(new_Jinkela_wire_276),
        .b(_1203_),
        .c(_1204_)
    );

    bfr new_Jinkela_buffer_4575 (
        .din(new_Jinkela_wire_6267),
        .dout(new_Jinkela_wire_6268)
    );

    bfr new_Jinkela_buffer_5937 (
        .din(new_Jinkela_wire_7985),
        .dout(new_Jinkela_wire_7986)
    );

    or_ii _1916_ (
        .a(new_Jinkela_wire_449),
        .b(new_Jinkela_wire_1204),
        .c(_1205_)
    );

    bfr new_Jinkela_buffer_4591 (
        .din(new_Jinkela_wire_6287),
        .dout(new_Jinkela_wire_6288)
    );

    and_bi _1917_ (
        .a(new_Jinkela_wire_1545),
        .b(new_Jinkela_wire_450),
        .c(_1206_)
    );

    bfr new_Jinkela_buffer_4576 (
        .din(new_Jinkela_wire_6268),
        .dout(new_Jinkela_wire_6269)
    );

    bfr new_Jinkela_buffer_5938 (
        .din(new_Jinkela_wire_7986),
        .dout(new_Jinkela_wire_7987)
    );

    and_bi _1918_ (
        .a(_1205_),
        .b(_1206_),
        .c(_1207_)
    );

    spl2 new_Jinkela_splitter_653 (
        .a(new_Jinkela_wire_6317),
        .b(new_Jinkela_wire_6318),
        .c(new_Jinkela_wire_6319)
    );

    bfr new_Jinkela_buffer_5956 (
        .din(new_Jinkela_wire_8004),
        .dout(new_Jinkela_wire_8005)
    );

    and_bi _1919_ (
        .a(new_Jinkela_wire_1857),
        .b(_1207_),
        .c(_1208_)
    );

    bfr new_Jinkela_buffer_4577 (
        .din(new_Jinkela_wire_6269),
        .dout(new_Jinkela_wire_6270)
    );

    bfr new_Jinkela_buffer_5939 (
        .din(new_Jinkela_wire_7987),
        .dout(new_Jinkela_wire_7988)
    );

    and_ii _1920_ (
        .a(_1208_),
        .b(_1204_),
        .c(_1209_)
    );

    bfr new_Jinkela_buffer_4592 (
        .din(new_Jinkela_wire_6288),
        .dout(new_Jinkela_wire_6289)
    );

    or_bb _1921_ (
        .a(new_Jinkela_wire_4982),
        .b(new_Jinkela_wire_3274),
        .c(_1210_)
    );

    bfr new_Jinkela_buffer_4578 (
        .din(new_Jinkela_wire_6270),
        .dout(new_Jinkela_wire_6271)
    );

    bfr new_Jinkela_buffer_5940 (
        .din(new_Jinkela_wire_7988),
        .dout(new_Jinkela_wire_7989)
    );

    and_bb _1922_ (
        .a(new_Jinkela_wire_4983),
        .b(new_Jinkela_wire_3275),
        .c(_1211_)
    );

    spl4L new_Jinkela_splitter_654 (
        .a(new_Jinkela_wire_6320),
        .d(new_Jinkela_wire_6321),
        .e(new_Jinkela_wire_6322),
        .b(new_Jinkela_wire_6323),
        .c(new_Jinkela_wire_6324)
    );

    bfr new_Jinkela_buffer_5957 (
        .din(new_Jinkela_wire_8005),
        .dout(new_Jinkela_wire_8006)
    );

    bfr new_Jinkela_buffer_4620 (
        .din(new_Jinkela_wire_6324),
        .dout(new_Jinkela_wire_6325)
    );

    and_bi _1923_ (
        .a(_1210_),
        .b(_1211_),
        .c(_1212_)
    );

    bfr new_Jinkela_buffer_4579 (
        .din(new_Jinkela_wire_6271),
        .dout(new_Jinkela_wire_6272)
    );

    bfr new_Jinkela_buffer_5941 (
        .din(new_Jinkela_wire_7989),
        .dout(new_Jinkela_wire_7990)
    );

    and_ii _1924_ (
        .a(new_Jinkela_wire_2423),
        .b(new_Jinkela_wire_4175),
        .c(_1213_)
    );

    bfr new_Jinkela_buffer_4593 (
        .din(new_Jinkela_wire_6289),
        .dout(new_Jinkela_wire_6290)
    );

    and_bb _1925_ (
        .a(new_Jinkela_wire_2424),
        .b(new_Jinkela_wire_4176),
        .c(_1214_)
    );

    bfr new_Jinkela_buffer_4580 (
        .din(new_Jinkela_wire_6272),
        .dout(new_Jinkela_wire_6273)
    );

    bfr new_Jinkela_buffer_5942 (
        .din(new_Jinkela_wire_7990),
        .dout(new_Jinkela_wire_7991)
    );

    and_ii _1926_ (
        .a(_1214_),
        .b(_1213_),
        .c(_1215_)
    );

    bfr new_Jinkela_buffer_4625 (
        .din(new_Jinkela_wire_6329),
        .dout(new_Jinkela_wire_6330)
    );

    bfr new_Jinkela_buffer_5958 (
        .din(new_Jinkela_wire_8006),
        .dout(new_Jinkela_wire_8007)
    );

    and_ii _1927_ (
        .a(new_Jinkela_wire_5238),
        .b(new_Jinkela_wire_1679),
        .c(_1216_)
    );

    bfr new_Jinkela_buffer_4581 (
        .din(new_Jinkela_wire_6273),
        .dout(new_Jinkela_wire_6274)
    );

    bfr new_Jinkela_buffer_5943 (
        .din(new_Jinkela_wire_7991),
        .dout(new_Jinkela_wire_7992)
    );

    and_bb _1928_ (
        .a(new_Jinkela_wire_5239),
        .b(new_Jinkela_wire_1680),
        .c(_1217_)
    );

    bfr new_Jinkela_buffer_4594 (
        .din(new_Jinkela_wire_6290),
        .dout(new_Jinkela_wire_6291)
    );

    or_bb _1929_ (
        .a(_1217_),
        .b(_1216_),
        .c(_1218_)
    );

    bfr new_Jinkela_buffer_4582 (
        .din(new_Jinkela_wire_6274),
        .dout(new_Jinkela_wire_6275)
    );

    bfr new_Jinkela_buffer_5959 (
        .din(new_Jinkela_wire_8007),
        .dout(new_Jinkela_wire_8008)
    );

    or_bi _1930_ (
        .a(new_Jinkela_wire_4112),
        .b(new_Jinkela_wire_5597),
        .c(_1219_)
    );

    bfr new_Jinkela_buffer_4645 (
        .din(new_Jinkela_wire_6349),
        .dout(new_Jinkela_wire_6350)
    );

    and_bi _1931_ (
        .a(new_Jinkela_wire_4113),
        .b(new_Jinkela_wire_5598),
        .c(_1220_)
    );

    bfr new_Jinkela_buffer_4583 (
        .din(new_Jinkela_wire_6275),
        .dout(new_Jinkela_wire_6276)
    );

    bfr new_Jinkela_buffer_5960 (
        .din(new_Jinkela_wire_8008),
        .dout(new_Jinkela_wire_8009)
    );

    or_bb _1932_ (
        .a(_1220_),
        .b(new_Jinkela_wire_7699),
        .c(_1221_)
    );

    bfr new_Jinkela_buffer_4595 (
        .din(new_Jinkela_wire_6291),
        .dout(new_Jinkela_wire_6292)
    );

    and_bi _1933_ (
        .a(new_Jinkela_wire_5216),
        .b(_1221_),
        .c(_1222_)
    );

    bfr new_Jinkela_buffer_4584 (
        .din(new_Jinkela_wire_6276),
        .dout(new_Jinkela_wire_6277)
    );

    bfr new_Jinkela_buffer_5961 (
        .din(new_Jinkela_wire_8009),
        .dout(new_Jinkela_wire_8010)
    );

    or_bb _1934_ (
        .a(_1222_),
        .b(new_Jinkela_wire_4856),
        .c(_1223_)
    );

    bfr new_Jinkela_buffer_4626 (
        .din(new_Jinkela_wire_6330),
        .dout(new_Jinkela_wire_6331)
    );

    bfr new_Jinkela_buffer_4621 (
        .din(new_Jinkela_wire_6325),
        .dout(new_Jinkela_wire_6326)
    );

    or_bi _1935_ (
        .a(new_Jinkela_wire_5212),
        .b(_1125_),
        .c(_1224_)
    );

    bfr new_Jinkela_buffer_4585 (
        .din(new_Jinkela_wire_6277),
        .dout(new_Jinkela_wire_6278)
    );

    bfr new_Jinkela_buffer_5962 (
        .din(new_Jinkela_wire_8010),
        .dout(new_Jinkela_wire_8011)
    );

    or_bi _1936_ (
        .a(new_Jinkela_wire_1400),
        .b(new_Jinkela_wire_1369),
        .c(_1225_)
    );

    bfr new_Jinkela_buffer_4596 (
        .din(new_Jinkela_wire_6292),
        .dout(new_Jinkela_wire_6293)
    );

    or_ii _1937_ (
        .a(new_Jinkela_wire_2243),
        .b(new_Jinkela_wire_7605),
        .c(_1226_)
    );

    spl2 new_Jinkela_splitter_650 (
        .a(new_Jinkela_wire_6278),
        .b(new_Jinkela_wire_6279),
        .c(new_Jinkela_wire_6280)
    );

    bfr new_Jinkela_buffer_5963 (
        .din(new_Jinkela_wire_8011),
        .dout(new_Jinkela_wire_8012)
    );

    and_bi _1938_ (
        .a(new_Jinkela_wire_1675),
        .b(new_Jinkela_wire_3413),
        .c(_1227_)
    );

    spl2 new_Jinkela_splitter_651 (
        .a(new_Jinkela_wire_6280),
        .b(new_Jinkela_wire_6281),
        .c(new_Jinkela_wire_6282)
    );

    inv _1939_ (
        .din(new_Jinkela_wire_836),
        .dout(_1228_)
    );

    bfr new_Jinkela_buffer_5964 (
        .din(new_Jinkela_wire_8012),
        .dout(new_Jinkela_wire_8013)
    );

    and_bi _1940_ (
        .a(new_Jinkela_wire_1885),
        .b(new_Jinkela_wire_6318),
        .c(_1229_)
    );

    bfr new_Jinkela_buffer_4650 (
        .din(_0176_),
        .dout(new_Jinkela_wire_6363)
    );

    bfr new_Jinkela_buffer_4622 (
        .din(new_Jinkela_wire_6326),
        .dout(new_Jinkela_wire_6327)
    );

    or_bi _1941_ (
        .a(new_Jinkela_wire_5247),
        .b(new_Jinkela_wire_5636),
        .c(_1230_)
    );

    bfr new_Jinkela_buffer_4597 (
        .din(new_Jinkela_wire_6293),
        .dout(new_Jinkela_wire_6294)
    );

    bfr new_Jinkela_buffer_5965 (
        .din(new_Jinkela_wire_8013),
        .dout(new_Jinkela_wire_8014)
    );

    and_bi _1942_ (
        .a(new_Jinkela_wire_7112),
        .b(new_Jinkela_wire_1888),
        .c(_1231_)
    );

    bfr new_Jinkela_buffer_4598 (
        .din(new_Jinkela_wire_6294),
        .dout(new_Jinkela_wire_6295)
    );

    or_bb _1943_ (
        .a(_1231_),
        .b(new_Jinkela_wire_5249),
        .c(_1232_)
    );

    bfr new_Jinkela_buffer_5966 (
        .din(new_Jinkela_wire_8014),
        .dout(new_Jinkela_wire_8015)
    );

    and_ii _1944_ (
        .a(new_Jinkela_wire_3357),
        .b(new_Jinkela_wire_6328),
        .c(_1233_)
    );

    bfr new_Jinkela_buffer_4599 (
        .din(new_Jinkela_wire_6295),
        .dout(new_Jinkela_wire_6296)
    );

    and_bi _1945_ (
        .a(new_Jinkela_wire_7197),
        .b(_1233_),
        .c(_1234_)
    );

    bfr new_Jinkela_buffer_4627 (
        .din(new_Jinkela_wire_6331),
        .dout(new_Jinkela_wire_6332)
    );

    bfr new_Jinkela_buffer_5967 (
        .din(new_Jinkela_wire_8015),
        .dout(new_Jinkela_wire_8016)
    );

    bfr new_Jinkela_buffer_4623 (
        .din(new_Jinkela_wire_6327),
        .dout(new_Jinkela_wire_6328)
    );

    and_bi _1946_ (
        .a(new_Jinkela_wire_4798),
        .b(_1234_),
        .c(_1235_)
    );

    bfr new_Jinkela_buffer_4600 (
        .din(new_Jinkela_wire_6296),
        .dout(new_Jinkela_wire_6297)
    );

    and_ii _1947_ (
        .a(new_Jinkela_wire_6323),
        .b(new_Jinkela_wire_2770),
        .c(_1236_)
    );

    bfr new_Jinkela_buffer_5968 (
        .din(new_Jinkela_wire_8016),
        .dout(new_Jinkela_wire_8017)
    );

    and_bb _1948_ (
        .a(new_Jinkela_wire_6321),
        .b(new_Jinkela_wire_2774),
        .c(_1237_)
    );

    bfr new_Jinkela_buffer_4601 (
        .din(new_Jinkela_wire_6297),
        .dout(new_Jinkela_wire_6298)
    );

    bfr new_Jinkela_buffer_1669 (
        .din(new_Jinkela_wire_2680),
        .dout(new_Jinkela_wire_2681)
    );

    bfr new_Jinkela_buffer_5352 (
        .din(new_Jinkela_wire_7278),
        .dout(new_Jinkela_wire_7279)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    bfr new_Jinkela_buffer_128 (
        .din(G93),
        .dout(new_Jinkela_wire_308)
    );

    bfr new_Jinkela_buffer_1687 (
        .din(new_Jinkela_wire_2698),
        .dout(new_Jinkela_wire_2699)
    );

    bfr new_Jinkela_buffer_5385 (
        .din(new_Jinkela_wire_7317),
        .dout(new_Jinkela_wire_7318)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_305),
        .dout(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_1670 (
        .din(new_Jinkela_wire_2681),
        .dout(new_Jinkela_wire_2682)
    );

    bfr new_Jinkela_buffer_5353 (
        .din(new_Jinkela_wire_7279),
        .dout(new_Jinkela_wire_7280)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_1720 (
        .din(new_Jinkela_wire_2731),
        .dout(new_Jinkela_wire_2732)
    );

    bfr new_Jinkela_buffer_5367 (
        .din(new_Jinkela_wire_7299),
        .dout(new_Jinkela_wire_7300)
    );

    spl2 new_Jinkela_splitter_61 (
        .a(G169),
        .b(new_Jinkela_wire_310),
        .c(new_Jinkela_wire_313)
    );

    bfr new_Jinkela_buffer_1671 (
        .din(new_Jinkela_wire_2682),
        .dout(new_Jinkela_wire_2683)
    );

    bfr new_Jinkela_buffer_5354 (
        .din(new_Jinkela_wire_7280),
        .dout(new_Jinkela_wire_7281)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_1688 (
        .din(new_Jinkela_wire_2699),
        .dout(new_Jinkela_wire_2700)
    );

    bfr new_Jinkela_buffer_5459 (
        .din(new_net_2367),
        .dout(new_Jinkela_wire_7392)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_1672 (
        .din(new_Jinkela_wire_2683),
        .dout(new_Jinkela_wire_2684)
    );

    bfr new_Jinkela_buffer_5355 (
        .din(new_Jinkela_wire_7281),
        .dout(new_Jinkela_wire_7282)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_5368 (
        .din(new_Jinkela_wire_7300),
        .dout(new_Jinkela_wire_7301)
    );

    spl2 new_Jinkela_splitter_383 (
        .a(new_Jinkela_wire_2780),
        .b(new_Jinkela_wire_2781),
        .c(new_Jinkela_wire_2782)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_1689 (
        .din(new_Jinkela_wire_2700),
        .dout(new_Jinkela_wire_2701)
    );

    bfr new_Jinkela_buffer_5356 (
        .din(new_Jinkela_wire_7282),
        .dout(new_Jinkela_wire_7283)
    );

    bfr new_Jinkela_buffer_1721 (
        .din(new_Jinkela_wire_2732),
        .dout(new_Jinkela_wire_2733)
    );

    bfr new_Jinkela_buffer_5386 (
        .din(new_Jinkela_wire_7318),
        .dout(new_Jinkela_wire_7319)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_315),
        .dout(new_Jinkela_wire_316)
    );

    bfr new_Jinkela_buffer_131 (
        .din(G87),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_1690 (
        .din(new_Jinkela_wire_2701),
        .dout(new_Jinkela_wire_2702)
    );

    bfr new_Jinkela_buffer_5357 (
        .din(new_Jinkela_wire_7283),
        .dout(new_Jinkela_wire_7284)
    );

    bfr new_Jinkela_buffer_137 (
        .din(G50),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_5369 (
        .din(new_Jinkela_wire_7301),
        .dout(new_Jinkela_wire_7302)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    bfr new_Jinkela_buffer_1756 (
        .din(new_Jinkela_wire_2782),
        .dout(new_Jinkela_wire_2783)
    );

    bfr new_Jinkela_buffer_1691 (
        .din(new_Jinkela_wire_2702),
        .dout(new_Jinkela_wire_2703)
    );

    bfr new_Jinkela_buffer_5358 (
        .din(new_Jinkela_wire_7284),
        .dout(new_Jinkela_wire_7285)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_311),
        .c(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_1722 (
        .din(new_Jinkela_wire_2733),
        .dout(new_Jinkela_wire_2734)
    );

    bfr new_Jinkela_buffer_5421 (
        .din(new_Jinkela_wire_7353),
        .dout(new_Jinkela_wire_7354)
    );

    spl4L new_Jinkela_splitter_63 (
        .a(new_Jinkela_wire_313),
        .d(new_Jinkela_wire_314),
        .e(new_Jinkela_wire_315),
        .b(new_Jinkela_wire_317),
        .c(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_1692 (
        .din(new_Jinkela_wire_2703),
        .dout(new_Jinkela_wire_2704)
    );

    bfr new_Jinkela_buffer_5359 (
        .din(new_Jinkela_wire_7285),
        .dout(new_Jinkela_wire_7286)
    );

    bfr new_Jinkela_buffer_134 (
        .din(G73),
        .dout(new_Jinkela_wire_332)
    );

    spl2 new_Jinkela_splitter_382 (
        .a(new_Jinkela_wire_2776),
        .b(new_Jinkela_wire_2777),
        .c(new_Jinkela_wire_2778)
    );

    bfr new_Jinkela_buffer_5370 (
        .din(new_Jinkela_wire_7302),
        .dout(new_Jinkela_wire_7303)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_317),
        .d(new_Jinkela_wire_318),
        .e(new_Jinkela_wire_319),
        .b(new_Jinkela_wire_320),
        .c(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_1693 (
        .din(new_Jinkela_wire_2704),
        .dout(new_Jinkela_wire_2705)
    );

    bfr new_Jinkela_buffer_5360 (
        .din(new_Jinkela_wire_7286),
        .dout(new_Jinkela_wire_7287)
    );

    spl4L new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_322),
        .d(new_Jinkela_wire_323),
        .e(new_Jinkela_wire_324),
        .b(new_Jinkela_wire_325),
        .c(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_1723 (
        .din(new_Jinkela_wire_2734),
        .dout(new_Jinkela_wire_2735)
    );

    bfr new_Jinkela_buffer_5387 (
        .din(new_Jinkela_wire_7319),
        .dout(new_Jinkela_wire_7320)
    );

    bfr new_Jinkela_buffer_1694 (
        .din(new_Jinkela_wire_2705),
        .dout(new_Jinkela_wire_2706)
    );

    bfr new_Jinkela_buffer_5361 (
        .din(new_Jinkela_wire_7287),
        .dout(new_Jinkela_wire_7288)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    spl3L new_Jinkela_splitter_68 (
        .a(G174),
        .d(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_343),
        .c(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_5371 (
        .din(new_Jinkela_wire_7303),
        .dout(new_Jinkela_wire_7304)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    bfr new_Jinkela_buffer_1779 (
        .din(new_Jinkela_wire_2805),
        .dout(new_Jinkela_wire_2806)
    );

    bfr new_Jinkela_buffer_1695 (
        .din(new_Jinkela_wire_2706),
        .dout(new_Jinkela_wire_2707)
    );

    bfr new_Jinkela_buffer_5439 (
        .din(new_Jinkela_wire_7371),
        .dout(new_Jinkela_wire_7372)
    );

    spl2 new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_329),
        .b(new_Jinkela_wire_330),
        .c(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_1724 (
        .din(new_Jinkela_wire_2735),
        .dout(new_Jinkela_wire_2736)
    );

    bfr new_Jinkela_buffer_5372 (
        .din(new_Jinkela_wire_7304),
        .dout(new_Jinkela_wire_7305)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_1696 (
        .din(new_Jinkela_wire_2707),
        .dout(new_Jinkela_wire_2708)
    );

    bfr new_Jinkela_buffer_5388 (
        .din(new_Jinkela_wire_7320),
        .dout(new_Jinkela_wire_7321)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_337),
        .dout(new_Jinkela_wire_338)
    );

    bfr new_Jinkela_buffer_5373 (
        .din(new_Jinkela_wire_7305),
        .dout(new_Jinkela_wire_7306)
    );

    spl2 new_Jinkela_splitter_387 (
        .a(_0584_),
        .b(new_Jinkela_wire_2841),
        .c(new_Jinkela_wire_2842)
    );

    bfr new_Jinkela_buffer_1697 (
        .din(new_Jinkela_wire_2708),
        .dout(new_Jinkela_wire_2709)
    );

    bfr new_Jinkela_buffer_5422 (
        .din(new_Jinkela_wire_7354),
        .dout(new_Jinkela_wire_7355)
    );

    spl2 new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_334),
        .b(new_Jinkela_wire_335),
        .c(new_Jinkela_wire_336)
    );

    bfr new_Jinkela_buffer_1725 (
        .din(new_Jinkela_wire_2736),
        .dout(new_Jinkela_wire_2737)
    );

    bfr new_Jinkela_buffer_5374 (
        .din(new_Jinkela_wire_7306),
        .dout(new_Jinkela_wire_7307)
    );

    spl4L new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_416),
        .d(new_Jinkela_wire_417),
        .e(new_Jinkela_wire_418),
        .b(new_Jinkela_wire_419),
        .c(new_Jinkela_wire_420)
    );

    bfr new_Jinkela_buffer_1698 (
        .din(new_Jinkela_wire_2709),
        .dout(new_Jinkela_wire_2710)
    );

    bfr new_Jinkela_buffer_5389 (
        .din(new_Jinkela_wire_7321),
        .dout(new_Jinkela_wire_7322)
    );

    spl4L new_Jinkela_splitter_96 (
        .a(G158),
        .d(new_Jinkela_wire_452),
        .e(new_Jinkela_wire_453),
        .b(new_Jinkela_wire_454),
        .c(new_Jinkela_wire_455)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_338),
        .dout(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_1785 (
        .din(new_Jinkela_wire_2818),
        .dout(new_Jinkela_wire_2819)
    );

    bfr new_Jinkela_buffer_5375 (
        .din(new_Jinkela_wire_7307),
        .dout(new_Jinkela_wire_7308)
    );

    spl3L new_Jinkela_splitter_105 (
        .a(G161),
        .d(new_Jinkela_wire_500),
        .b(new_Jinkela_wire_501),
        .c(new_Jinkela_wire_502)
    );

    bfr new_Jinkela_buffer_1757 (
        .din(new_Jinkela_wire_2783),
        .dout(new_Jinkela_wire_2784)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_1699 (
        .din(new_Jinkela_wire_2710),
        .dout(new_Jinkela_wire_2711)
    );

    bfr new_Jinkela_buffer_5499 (
        .din(_0080_),
        .dout(new_Jinkela_wire_7432)
    );

    spl4L new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_411),
        .d(new_Jinkela_wire_412),
        .e(new_Jinkela_wire_413),
        .b(new_Jinkela_wire_414),
        .c(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_1726 (
        .din(new_Jinkela_wire_2737),
        .dout(new_Jinkela_wire_2738)
    );

    bfr new_Jinkela_buffer_5376 (
        .din(new_Jinkela_wire_7308),
        .dout(new_Jinkela_wire_7309)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_340),
        .dout(new_Jinkela_wire_341)
    );

    bfr new_Jinkela_buffer_1700 (
        .din(new_Jinkela_wire_2711),
        .dout(new_Jinkela_wire_2712)
    );

    bfr new_Jinkela_buffer_5390 (
        .din(new_Jinkela_wire_7322),
        .dout(new_Jinkela_wire_7323)
    );

    bfr new_Jinkela_buffer_5377 (
        .din(new_Jinkela_wire_7309),
        .dout(new_Jinkela_wire_7310)
    );

    spl3L new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_407),
        .d(new_Jinkela_wire_408),
        .b(new_Jinkela_wire_409),
        .c(new_Jinkela_wire_410)
    );

    spl3L new_Jinkela_splitter_388 (
        .a(_0738_),
        .d(new_Jinkela_wire_2845),
        .b(new_Jinkela_wire_2846),
        .c(new_Jinkela_wire_2847)
    );

    bfr new_Jinkela_buffer_1701 (
        .din(new_Jinkela_wire_2712),
        .dout(new_Jinkela_wire_2713)
    );

    bfr new_Jinkela_buffer_5423 (
        .din(new_Jinkela_wire_7355),
        .dout(new_Jinkela_wire_7356)
    );

    bfr new_Jinkela_buffer_1727 (
        .din(new_Jinkela_wire_2738),
        .dout(new_Jinkela_wire_2739)
    );

    bfr new_Jinkela_buffer_5378 (
        .din(new_Jinkela_wire_7310),
        .dout(new_Jinkela_wire_7311)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_1702 (
        .din(new_Jinkela_wire_2713),
        .dout(new_Jinkela_wire_2714)
    );

    bfr new_Jinkela_buffer_5391 (
        .din(new_Jinkela_wire_7323),
        .dout(new_Jinkela_wire_7324)
    );

    bfr new_Jinkela_buffer_167 (
        .din(G103),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_5379 (
        .din(new_Jinkela_wire_7311),
        .dout(new_Jinkela_wire_7312)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_1758 (
        .din(new_Jinkela_wire_2784),
        .dout(new_Jinkela_wire_2785)
    );

    bfr new_Jinkela_buffer_1703 (
        .din(new_Jinkela_wire_2714),
        .dout(new_Jinkela_wire_2715)
    );

    bfr new_Jinkela_buffer_5440 (
        .din(new_Jinkela_wire_7372),
        .dout(new_Jinkela_wire_7373)
    );

    spl3L new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_422),
        .d(new_Jinkela_wire_423),
        .b(new_Jinkela_wire_424),
        .c(new_Jinkela_wire_425)
    );

    bfr new_Jinkela_buffer_1728 (
        .din(new_Jinkela_wire_2739),
        .dout(new_Jinkela_wire_2740)
    );

    bfr new_Jinkela_buffer_5380 (
        .din(new_Jinkela_wire_7312),
        .dout(new_Jinkela_wire_7313)
    );

    bfr new_Jinkela_buffer_165 (
        .din(G67),
        .dout(new_Jinkela_wire_421)
    );

    bfr new_Jinkela_buffer_1704 (
        .din(new_Jinkela_wire_2715),
        .dout(new_Jinkela_wire_2716)
    );

    bfr new_Jinkela_buffer_5392 (
        .din(new_Jinkela_wire_7324),
        .dout(new_Jinkela_wire_7325)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    spl4L new_Jinkela_splitter_90 (
        .a(new_Jinkela_wire_426),
        .d(new_Jinkela_wire_427),
        .e(new_Jinkela_wire_428),
        .b(new_Jinkela_wire_429),
        .c(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_5381 (
        .din(new_Jinkela_wire_7313),
        .dout(new_Jinkela_wire_7314)
    );

    bfr new_Jinkela_buffer_1705 (
        .din(new_Jinkela_wire_2716),
        .dout(new_Jinkela_wire_2717)
    );

    bfr new_Jinkela_buffer_5424 (
        .din(new_Jinkela_wire_7356),
        .dout(new_Jinkela_wire_7357)
    );

    spl3L new_Jinkela_splitter_88 (
        .a(G126),
        .d(new_Jinkela_wire_422),
        .b(new_Jinkela_wire_426),
        .c(new_Jinkela_wire_431)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_348),
        .dout(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_1729 (
        .din(new_Jinkela_wire_2740),
        .dout(new_Jinkela_wire_2741)
    );

    bfr new_Jinkela_buffer_5393 (
        .din(new_Jinkela_wire_7325),
        .dout(new_Jinkela_wire_7326)
    );

    bfr new_Jinkela_buffer_3218 (
        .din(new_Jinkela_wire_4591),
        .dout(new_Jinkela_wire_4592)
    );

    spl3L new_Jinkela_splitter_528 (
        .a(_0924_),
        .d(new_Jinkela_wire_4706),
        .b(new_Jinkela_wire_4707),
        .c(new_Jinkela_wire_4708)
    );

    bfr new_Jinkela_buffer_3233 (
        .din(new_Jinkela_wire_4617),
        .dout(new_Jinkela_wire_4618)
    );

    bfr new_Jinkela_buffer_3219 (
        .din(new_Jinkela_wire_4592),
        .dout(new_Jinkela_wire_4593)
    );

    bfr new_Jinkela_buffer_3319 (
        .din(new_net_2391),
        .dout(new_Jinkela_wire_4709)
    );

    bfr new_Jinkela_buffer_3220 (
        .din(new_Jinkela_wire_4593),
        .dout(new_Jinkela_wire_4594)
    );

    bfr new_Jinkela_buffer_3271 (
        .din(new_Jinkela_wire_4657),
        .dout(new_Jinkela_wire_4658)
    );

    bfr new_Jinkela_buffer_3234 (
        .din(new_Jinkela_wire_4618),
        .dout(new_Jinkela_wire_4619)
    );

    bfr new_Jinkela_buffer_3221 (
        .din(new_Jinkela_wire_4594),
        .dout(new_Jinkela_wire_4595)
    );

    bfr new_Jinkela_buffer_3222 (
        .din(new_Jinkela_wire_4595),
        .dout(new_Jinkela_wire_4596)
    );

    bfr new_Jinkela_buffer_3280 (
        .din(new_Jinkela_wire_4666),
        .dout(new_Jinkela_wire_4667)
    );

    bfr new_Jinkela_buffer_3235 (
        .din(new_Jinkela_wire_4619),
        .dout(new_Jinkela_wire_4620)
    );

    bfr new_Jinkela_buffer_3223 (
        .din(new_Jinkela_wire_4596),
        .dout(new_Jinkela_wire_4597)
    );

    spl2 new_Jinkela_splitter_522 (
        .a(new_Jinkela_wire_4597),
        .b(new_Jinkela_wire_4598),
        .c(new_Jinkela_wire_4599)
    );

    bfr new_Jinkela_buffer_3272 (
        .din(new_Jinkela_wire_4658),
        .dout(new_Jinkela_wire_4659)
    );

    bfr new_Jinkela_buffer_3236 (
        .din(new_Jinkela_wire_4620),
        .dout(new_Jinkela_wire_4621)
    );

    bfr new_Jinkela_buffer_3237 (
        .din(new_Jinkela_wire_4621),
        .dout(new_Jinkela_wire_4622)
    );

    spl2 new_Jinkela_splitter_529 (
        .a(_0668_),
        .b(new_Jinkela_wire_4712),
        .c(new_Jinkela_wire_4713)
    );

    bfr new_Jinkela_buffer_3273 (
        .din(new_Jinkela_wire_4659),
        .dout(new_Jinkela_wire_4660)
    );

    bfr new_Jinkela_buffer_3238 (
        .din(new_Jinkela_wire_4622),
        .dout(new_Jinkela_wire_4623)
    );

    bfr new_Jinkela_buffer_3281 (
        .din(new_Jinkela_wire_4667),
        .dout(new_Jinkela_wire_4668)
    );

    bfr new_Jinkela_buffer_3239 (
        .din(new_Jinkela_wire_4623),
        .dout(new_Jinkela_wire_4624)
    );

    bfr new_Jinkela_buffer_3274 (
        .din(new_Jinkela_wire_4660),
        .dout(new_Jinkela_wire_4661)
    );

    bfr new_Jinkela_buffer_3240 (
        .din(new_Jinkela_wire_4624),
        .dout(new_Jinkela_wire_4625)
    );

    bfr new_Jinkela_buffer_3323 (
        .din(new_net_2393),
        .dout(new_Jinkela_wire_4715)
    );

    bfr new_Jinkela_buffer_3241 (
        .din(new_Jinkela_wire_4625),
        .dout(new_Jinkela_wire_4626)
    );

    bfr new_Jinkela_buffer_3275 (
        .din(new_Jinkela_wire_4661),
        .dout(new_Jinkela_wire_4662)
    );

    bfr new_Jinkela_buffer_3242 (
        .din(new_Jinkela_wire_4626),
        .dout(new_Jinkela_wire_4627)
    );

    bfr new_Jinkela_buffer_3282 (
        .din(new_Jinkela_wire_4668),
        .dout(new_Jinkela_wire_4669)
    );

    bfr new_Jinkela_buffer_3243 (
        .din(new_Jinkela_wire_4627),
        .dout(new_Jinkela_wire_4628)
    );

    bfr new_Jinkela_buffer_3276 (
        .din(new_Jinkela_wire_4662),
        .dout(new_Jinkela_wire_4663)
    );

    bfr new_Jinkela_buffer_3244 (
        .din(new_Jinkela_wire_4628),
        .dout(new_Jinkela_wire_4629)
    );

    bfr new_Jinkela_buffer_3320 (
        .din(new_Jinkela_wire_4709),
        .dout(new_Jinkela_wire_4710)
    );

    bfr new_Jinkela_buffer_3245 (
        .din(new_Jinkela_wire_4629),
        .dout(new_Jinkela_wire_4630)
    );

    bfr new_Jinkela_buffer_3277 (
        .din(new_Jinkela_wire_4663),
        .dout(new_Jinkela_wire_4664)
    );

    bfr new_Jinkela_buffer_3246 (
        .din(new_Jinkela_wire_4630),
        .dout(new_Jinkela_wire_4631)
    );

    bfr new_Jinkela_buffer_3283 (
        .din(new_Jinkela_wire_4669),
        .dout(new_Jinkela_wire_4670)
    );

    bfr new_Jinkela_buffer_3247 (
        .din(new_Jinkela_wire_4631),
        .dout(new_Jinkela_wire_4632)
    );

    bfr new_Jinkela_buffer_3278 (
        .din(new_Jinkela_wire_4664),
        .dout(new_Jinkela_wire_4665)
    );

    bfr new_Jinkela_buffer_3248 (
        .din(new_Jinkela_wire_4632),
        .dout(new_Jinkela_wire_4633)
    );

    bfr new_Jinkela_buffer_3322 (
        .din(new_Jinkela_wire_4713),
        .dout(new_Jinkela_wire_4714)
    );

    bfr new_Jinkela_buffer_3249 (
        .din(new_Jinkela_wire_4633),
        .dout(new_Jinkela_wire_4634)
    );

    bfr new_Jinkela_buffer_3284 (
        .din(new_Jinkela_wire_4670),
        .dout(new_Jinkela_wire_4671)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1637),
        .dout(new_Jinkela_wire_1638)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1638),
        .dout(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1686),
        .dout(new_Jinkela_wire_1687)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1639),
        .dout(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1640),
        .dout(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1687),
        .dout(new_Jinkela_wire_1688)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1641),
        .dout(new_Jinkela_wire_1642)
    );

    spl2 new_Jinkela_splitter_321 (
        .a(new_Jinkela_wire_1752),
        .b(new_Jinkela_wire_1753),
        .c(new_Jinkela_wire_1754)
    );

    bfr new_Jinkela_buffer_876 (
        .din(_0512_),
        .dout(new_Jinkela_wire_1756)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1642),
        .dout(new_Jinkela_wire_1643)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1688),
        .dout(new_Jinkela_wire_1689)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    spl2 new_Jinkela_splitter_301 (
        .a(new_Jinkela_wire_1644),
        .b(new_Jinkela_wire_1645),
        .c(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1689),
        .dout(new_Jinkela_wire_1690)
    );

    bfr new_Jinkela_buffer_908 (
        .din(_0570_),
        .dout(new_Jinkela_wire_1788)
    );

    spl2 new_Jinkela_splitter_302 (
        .a(new_Jinkela_wire_1647),
        .b(new_Jinkela_wire_1648),
        .c(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1690),
        .dout(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_875 (
        .din(_1097_),
        .dout(new_Jinkela_wire_1755)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1709),
        .dout(new_Jinkela_wire_1710)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1650),
        .dout(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1691),
        .dout(new_Jinkela_wire_1692)
    );

    spl2 new_Jinkela_splitter_303 (
        .a(new_Jinkela_wire_1651),
        .b(new_Jinkela_wire_1652),
        .c(new_Jinkela_wire_1653)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1653),
        .dout(new_Jinkela_wire_1654)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1692),
        .dout(new_Jinkela_wire_1693)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1654),
        .dout(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1710),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1711),
        .dout(new_Jinkela_wire_1712)
    );

    spl2 new_Jinkela_splitter_304 (
        .a(new_Jinkela_wire_1655),
        .b(new_Jinkela_wire_1656),
        .c(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1657),
        .dout(new_Jinkela_wire_1658)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1693),
        .dout(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_941 (
        .din(_0497_),
        .dout(new_Jinkela_wire_1821)
    );

    spl2 new_Jinkela_splitter_305 (
        .a(new_Jinkela_wire_1658),
        .b(new_Jinkela_wire_1659),
        .c(new_Jinkela_wire_1660)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1660),
        .dout(new_Jinkela_wire_1661)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1694),
        .dout(new_Jinkela_wire_1695)
    );

    spl2 new_Jinkela_splitter_306 (
        .a(new_Jinkela_wire_1661),
        .b(new_Jinkela_wire_1662),
        .c(new_Jinkela_wire_1663)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_1663),
        .dout(new_Jinkela_wire_1664)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_1695),
        .dout(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1757),
        .dout(new_Jinkela_wire_1758)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_840),
        .dout(new_Jinkela_wire_841)
    );

    bfr new_Jinkela_buffer_1648 (
        .din(new_Jinkela_wire_2659),
        .dout(new_Jinkela_wire_2660)
    );

    bfr new_Jinkela_buffer_4531 (
        .din(new_Jinkela_wire_6206),
        .dout(new_Jinkela_wire_6207)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_5969 (
        .din(new_Jinkela_wire_8017),
        .dout(new_Jinkela_wire_8018)
    );

    bfr new_Jinkela_buffer_1755 (
        .din(new_net_16),
        .dout(new_Jinkela_wire_2780)
    );

    spl2 new_Jinkela_splitter_643 (
        .a(new_Jinkela_wire_6229),
        .b(new_Jinkela_wire_6230),
        .c(new_Jinkela_wire_6231)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(G123),
        .b(new_Jinkela_wire_867),
        .c(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_1649 (
        .din(new_Jinkela_wire_2660),
        .dout(new_Jinkela_wire_2661)
    );

    bfr new_Jinkela_buffer_4532 (
        .din(new_Jinkela_wire_6207),
        .dout(new_Jinkela_wire_6208)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_787),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_5970 (
        .din(new_Jinkela_wire_8018),
        .dout(new_Jinkela_wire_8019)
    );

    bfr new_Jinkela_buffer_1677 (
        .din(new_Jinkela_wire_2688),
        .dout(new_Jinkela_wire_2689)
    );

    bfr new_Jinkela_buffer_4542 (
        .din(new_Jinkela_wire_6217),
        .dout(new_Jinkela_wire_6218)
    );

    spl4L new_Jinkela_splitter_164 (
        .a(new_Jinkela_wire_849),
        .d(new_Jinkela_wire_850),
        .e(new_Jinkela_wire_851),
        .b(new_Jinkela_wire_852),
        .c(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_841),
        .dout(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_1650 (
        .din(new_Jinkela_wire_2661),
        .dout(new_Jinkela_wire_2662)
    );

    bfr new_Jinkela_buffer_4533 (
        .din(new_Jinkela_wire_6208),
        .dout(new_Jinkela_wire_6209)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_5971 (
        .din(new_Jinkela_wire_8019),
        .dout(new_Jinkela_wire_8020)
    );

    bfr new_Jinkela_buffer_1715 (
        .din(new_Jinkela_wire_2726),
        .dout(new_Jinkela_wire_2727)
    );

    bfr new_Jinkela_buffer_391 (
        .din(G83),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_1651 (
        .din(new_Jinkela_wire_2662),
        .dout(new_Jinkela_wire_2663)
    );

    bfr new_Jinkela_buffer_4534 (
        .din(new_Jinkela_wire_6209),
        .dout(new_Jinkela_wire_6210)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_5972 (
        .din(new_Jinkela_wire_8020),
        .dout(new_Jinkela_wire_8021)
    );

    bfr new_Jinkela_buffer_1678 (
        .din(new_Jinkela_wire_2689),
        .dout(new_Jinkela_wire_2690)
    );

    bfr new_Jinkela_buffer_4543 (
        .din(new_Jinkela_wire_6218),
        .dout(new_Jinkela_wire_6219)
    );

    spl3L new_Jinkela_splitter_163 (
        .a(new_Jinkela_wire_845),
        .d(new_Jinkela_wire_846),
        .b(new_Jinkela_wire_847),
        .c(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_1652 (
        .din(new_Jinkela_wire_2663),
        .dout(new_Jinkela_wire_2664)
    );

    bfr new_Jinkela_buffer_4535 (
        .din(new_Jinkela_wire_6210),
        .dout(new_Jinkela_wire_6211)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    spl3L new_Jinkela_splitter_380 (
        .a(new_Jinkela_wire_2767),
        .d(new_Jinkela_wire_2768),
        .b(new_Jinkela_wire_2769),
        .c(new_Jinkela_wire_2770)
    );

    spl4L new_Jinkela_splitter_381 (
        .a(new_Jinkela_wire_2771),
        .d(new_Jinkela_wire_2772),
        .e(new_Jinkela_wire_2773),
        .b(new_Jinkela_wire_2774),
        .c(new_Jinkela_wire_2775)
    );

    bfr new_Jinkela_buffer_1653 (
        .din(new_Jinkela_wire_2664),
        .dout(new_Jinkela_wire_2665)
    );

    bfr new_Jinkela_buffer_4544 (
        .din(new_Jinkela_wire_6219),
        .dout(new_Jinkela_wire_6220)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_791),
        .dout(new_Jinkela_wire_792)
    );

    bfr new_Jinkela_buffer_1679 (
        .din(new_Jinkela_wire_2690),
        .dout(new_Jinkela_wire_2691)
    );

    bfr new_Jinkela_buffer_4553 (
        .din(new_Jinkela_wire_6232),
        .dout(new_Jinkela_wire_6233)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    spl4L new_Jinkela_splitter_165 (
        .a(new_Jinkela_wire_854),
        .d(new_Jinkela_wire_855),
        .e(new_Jinkela_wire_856),
        .b(new_Jinkela_wire_857),
        .c(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_1654 (
        .din(new_Jinkela_wire_2665),
        .dout(new_Jinkela_wire_2666)
    );

    bfr new_Jinkela_buffer_4545 (
        .din(new_Jinkela_wire_6220),
        .dout(new_Jinkela_wire_6221)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    bfr new_Jinkela_buffer_1716 (
        .din(new_Jinkela_wire_2727),
        .dout(new_Jinkela_wire_2728)
    );

    spl2 new_Jinkela_splitter_648 (
        .a(_1015_),
        .b(new_Jinkela_wire_6250),
        .c(new_Jinkela_wire_6251)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_1655 (
        .din(new_Jinkela_wire_2666),
        .dout(new_Jinkela_wire_2667)
    );

    bfr new_Jinkela_buffer_4546 (
        .din(new_Jinkela_wire_6221),
        .dout(new_Jinkela_wire_6222)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_1680 (
        .din(new_Jinkela_wire_2691),
        .dout(new_Jinkela_wire_2692)
    );

    bfr new_Jinkela_buffer_4558 (
        .din(_0317_),
        .dout(new_Jinkela_wire_6247)
    );

    bfr new_Jinkela_buffer_4554 (
        .din(new_Jinkela_wire_6235),
        .dout(new_Jinkela_wire_6236)
    );

    bfr new_Jinkela_buffer_1656 (
        .din(new_Jinkela_wire_2667),
        .dout(new_Jinkela_wire_2668)
    );

    bfr new_Jinkela_buffer_4547 (
        .din(new_Jinkela_wire_6222),
        .dout(new_Jinkela_wire_6223)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    bfr new_Jinkela_buffer_4561 (
        .din(_0606_),
        .dout(new_Jinkela_wire_6252)
    );

    bfr new_Jinkela_buffer_1778 (
        .din(_0662_),
        .dout(new_Jinkela_wire_2805)
    );

    bfr new_Jinkela_buffer_1657 (
        .din(new_Jinkela_wire_2668),
        .dout(new_Jinkela_wire_2669)
    );

    bfr new_Jinkela_buffer_4548 (
        .din(new_Jinkela_wire_6223),
        .dout(new_Jinkela_wire_6224)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    bfr new_Jinkela_buffer_1681 (
        .din(new_Jinkela_wire_2692),
        .dout(new_Jinkela_wire_2693)
    );

    bfr new_Jinkela_buffer_4559 (
        .din(new_Jinkela_wire_6247),
        .dout(new_Jinkela_wire_6248)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_1658 (
        .din(new_Jinkela_wire_2669),
        .dout(new_Jinkela_wire_2670)
    );

    spl3L new_Jinkela_splitter_647 (
        .a(_0793_),
        .d(new_Jinkela_wire_6244),
        .b(new_Jinkela_wire_6245),
        .c(new_Jinkela_wire_6246)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_4567 (
        .din(_1076_),
        .dout(new_Jinkela_wire_6260)
    );

    bfr new_Jinkela_buffer_1717 (
        .din(new_Jinkela_wire_2728),
        .dout(new_Jinkela_wire_2729)
    );

    bfr new_Jinkela_buffer_4555 (
        .din(new_Jinkela_wire_6236),
        .dout(new_Jinkela_wire_6237)
    );

    bfr new_Jinkela_buffer_4556 (
        .din(new_Jinkela_wire_6237),
        .dout(new_Jinkela_wire_6238)
    );

    spl4L new_Jinkela_splitter_169 (
        .a(new_Jinkela_wire_871),
        .d(new_Jinkela_wire_872),
        .e(new_Jinkela_wire_877),
        .b(new_Jinkela_wire_882),
        .c(new_Jinkela_wire_887)
    );

    bfr new_Jinkela_buffer_1659 (
        .din(new_Jinkela_wire_2670),
        .dout(new_Jinkela_wire_2671)
    );

    spl2 new_Jinkela_splitter_150 (
        .a(new_Jinkela_wire_797),
        .b(new_Jinkela_wire_798),
        .c(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_4562 (
        .din(new_Jinkela_wire_6252),
        .dout(new_Jinkela_wire_6253)
    );

    bfr new_Jinkela_buffer_1682 (
        .din(new_Jinkela_wire_2693),
        .dout(new_Jinkela_wire_2694)
    );

    bfr new_Jinkela_buffer_4560 (
        .din(new_Jinkela_wire_6248),
        .dout(new_Jinkela_wire_6249)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    spl2 new_Jinkela_splitter_645 (
        .a(new_Jinkela_wire_6238),
        .b(new_Jinkela_wire_6239),
        .c(new_Jinkela_wire_6240)
    );

    bfr new_Jinkela_buffer_1660 (
        .din(new_Jinkela_wire_2671),
        .dout(new_Jinkela_wire_2672)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_4557 (
        .din(new_Jinkela_wire_6240),
        .dout(new_Jinkela_wire_6241)
    );

    bfr new_Jinkela_buffer_1784 (
        .din(_0379_),
        .dout(new_Jinkela_wire_2818)
    );

    bfr new_Jinkela_buffer_437 (
        .din(G46),
        .dout(new_Jinkela_wire_940)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_1661 (
        .din(new_Jinkela_wire_2672),
        .dout(new_Jinkela_wire_2673)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_1683 (
        .din(new_Jinkela_wire_2694),
        .dout(new_Jinkela_wire_2695)
    );

    bfr new_Jinkela_buffer_4565 (
        .din(_0076_),
        .dout(new_Jinkela_wire_6256)
    );

    spl2 new_Jinkela_splitter_166 (
        .a(new_Jinkela_wire_864),
        .b(new_Jinkela_wire_865),
        .c(new_Jinkela_wire_866)
    );

    spl2 new_Jinkela_splitter_646 (
        .a(new_Jinkela_wire_6241),
        .b(new_Jinkela_wire_6242),
        .c(new_Jinkela_wire_6243)
    );

    bfr new_Jinkela_buffer_1662 (
        .din(new_Jinkela_wire_2673),
        .dout(new_Jinkela_wire_2674)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    bfr new_Jinkela_buffer_1718 (
        .din(new_Jinkela_wire_2729),
        .dout(new_Jinkela_wire_2730)
    );

    bfr new_Jinkela_buffer_4563 (
        .din(new_Jinkela_wire_6253),
        .dout(new_Jinkela_wire_6254)
    );

    bfr new_Jinkela_buffer_395 (
        .din(G89),
        .dout(new_Jinkela_wire_894)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(G152),
        .b(new_Jinkela_wire_896),
        .c(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_1663 (
        .din(new_Jinkela_wire_2674),
        .dout(new_Jinkela_wire_2675)
    );

    bfr new_Jinkela_buffer_4566 (
        .din(new_Jinkela_wire_6256),
        .dout(new_Jinkela_wire_6257)
    );

    spl2 new_Jinkela_splitter_151 (
        .a(new_Jinkela_wire_802),
        .b(new_Jinkela_wire_803),
        .c(new_Jinkela_wire_804)
    );

    bfr new_Jinkela_buffer_1684 (
        .din(new_Jinkela_wire_2695),
        .dout(new_Jinkela_wire_2696)
    );

    bfr new_Jinkela_buffer_4586 (
        .din(_0008_),
        .dout(new_Jinkela_wire_6283)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_804),
        .dout(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_1664 (
        .din(new_Jinkela_wire_2675),
        .dout(new_Jinkela_wire_2676)
    );

    bfr new_Jinkela_buffer_4564 (
        .din(new_Jinkela_wire_6254),
        .dout(new_Jinkela_wire_6255)
    );

    bfr new_Jinkela_buffer_1753 (
        .din(new_Jinkela_wire_2775),
        .dout(new_Jinkela_wire_2776)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_1665 (
        .din(new_Jinkela_wire_2676),
        .dout(new_Jinkela_wire_2677)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    spl2 new_Jinkela_splitter_649 (
        .a(new_Jinkela_wire_6257),
        .b(new_Jinkela_wire_6258),
        .c(new_Jinkela_wire_6259)
    );

    bfr new_Jinkela_buffer_1685 (
        .din(new_Jinkela_wire_2696),
        .dout(new_Jinkela_wire_2697)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_1666 (
        .din(new_Jinkela_wire_2677),
        .dout(new_Jinkela_wire_2678)
    );

    spl2 new_Jinkela_splitter_652 (
        .a(_0862_),
        .b(new_Jinkela_wire_6317),
        .c(new_Jinkela_wire_6320)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_4587 (
        .din(_0577_),
        .dout(new_Jinkela_wire_6284)
    );

    bfr new_Jinkela_buffer_1719 (
        .din(new_Jinkela_wire_2730),
        .dout(new_Jinkela_wire_2731)
    );

    bfr new_Jinkela_buffer_4568 (
        .din(new_Jinkela_wire_6260),
        .dout(new_Jinkela_wire_6261)
    );

    bfr new_Jinkela_buffer_4624 (
        .din(new_net_2451),
        .dout(new_Jinkela_wire_6329)
    );

    spl2 new_Jinkela_splitter_168 (
        .a(new_Jinkela_wire_868),
        .b(new_Jinkela_wire_869),
        .c(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_1667 (
        .din(new_Jinkela_wire_2678),
        .dout(new_Jinkela_wire_2679)
    );

    bfr new_Jinkela_buffer_4569 (
        .din(new_Jinkela_wire_6261),
        .dout(new_Jinkela_wire_6262)
    );

    spl3L new_Jinkela_splitter_152 (
        .a(new_Jinkela_wire_807),
        .d(new_Jinkela_wire_808),
        .b(new_Jinkela_wire_809),
        .c(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_1686 (
        .din(new_Jinkela_wire_2697),
        .dout(new_Jinkela_wire_2698)
    );

    bfr new_Jinkela_buffer_4588 (
        .din(new_Jinkela_wire_6284),
        .dout(new_Jinkela_wire_6285)
    );

    spl4L new_Jinkela_splitter_171 (
        .a(new_Jinkela_wire_877),
        .d(new_Jinkela_wire_878),
        .e(new_Jinkela_wire_879),
        .b(new_Jinkela_wire_880),
        .c(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_1668 (
        .din(new_Jinkela_wire_2679),
        .dout(new_Jinkela_wire_2680)
    );

    bfr new_Jinkela_buffer_4570 (
        .din(new_Jinkela_wire_6262),
        .dout(new_Jinkela_wire_6263)
    );

    spl2 new_Jinkela_splitter_153 (
        .a(new_Jinkela_wire_810),
        .b(new_Jinkela_wire_811),
        .c(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_2748 (
        .din(new_Jinkela_wire_4056),
        .dout(new_Jinkela_wire_4057)
    );

    bfr new_Jinkela_buffer_2693 (
        .din(new_Jinkela_wire_3976),
        .dout(new_Jinkela_wire_3977)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    bfr new_Jinkela_buffer_2712 (
        .din(new_Jinkela_wire_4001),
        .dout(new_Jinkela_wire_4002)
    );

    bfr new_Jinkela_buffer_2694 (
        .din(new_Jinkela_wire_3977),
        .dout(new_Jinkela_wire_3978)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    bfr new_Jinkela_buffer_2737 (
        .din(new_Jinkela_wire_4039),
        .dout(new_Jinkela_wire_4040)
    );

    spl2 new_Jinkela_splitter_486 (
        .a(new_Jinkela_wire_3978),
        .b(new_Jinkela_wire_3979),
        .c(new_Jinkela_wire_3980)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_2695 (
        .din(new_Jinkela_wire_3980),
        .dout(new_Jinkela_wire_3981)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_2713 (
        .din(new_Jinkela_wire_4002),
        .dout(new_Jinkela_wire_4003)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    spl2 new_Jinkela_splitter_495 (
        .a(_0174_),
        .b(new_Jinkela_wire_4077),
        .c(new_Jinkela_wire_4078)
    );

    spl2 new_Jinkela_splitter_487 (
        .a(new_Jinkela_wire_3981),
        .b(new_Jinkela_wire_3982),
        .c(new_Jinkela_wire_3983)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    spl2 new_Jinkela_splitter_488 (
        .a(new_Jinkela_wire_3983),
        .b(new_Jinkela_wire_3984),
        .c(new_Jinkela_wire_3985)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    spl2 new_Jinkela_splitter_496 (
        .a(new_net_15),
        .b(new_Jinkela_wire_4079),
        .c(new_Jinkela_wire_4080)
    );

    bfr new_Jinkela_buffer_330 (
        .din(G4),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    bfr new_Jinkela_buffer_2714 (
        .din(new_Jinkela_wire_4003),
        .dout(new_Jinkela_wire_4004)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    bfr new_Jinkela_buffer_2715 (
        .din(new_Jinkela_wire_4004),
        .dout(new_Jinkela_wire_4005)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_2738 (
        .din(new_Jinkela_wire_4040),
        .dout(new_Jinkela_wire_4041)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_2767 (
        .din(new_Jinkela_wire_4075),
        .dout(new_Jinkela_wire_4076)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    bfr new_Jinkela_buffer_2716 (
        .din(new_Jinkela_wire_4005),
        .dout(new_Jinkela_wire_4006)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_2739 (
        .din(new_Jinkela_wire_4041),
        .dout(new_Jinkela_wire_4042)
    );

    bfr new_Jinkela_buffer_2717 (
        .din(new_Jinkela_wire_4006),
        .dout(new_Jinkela_wire_4007)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    bfr new_Jinkela_buffer_2749 (
        .din(new_Jinkela_wire_4057),
        .dout(new_Jinkela_wire_4058)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(new_Jinkela_wire_709),
        .b(new_Jinkela_wire_710),
        .c(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_2718 (
        .din(new_Jinkela_wire_4007),
        .dout(new_Jinkela_wire_4008)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    bfr new_Jinkela_buffer_2740 (
        .din(new_Jinkela_wire_4042),
        .dout(new_Jinkela_wire_4043)
    );

    bfr new_Jinkela_buffer_2719 (
        .din(new_Jinkela_wire_4008),
        .dout(new_Jinkela_wire_4009)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_2720 (
        .din(new_Jinkela_wire_4009),
        .dout(new_Jinkela_wire_4010)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    bfr new_Jinkela_buffer_2741 (
        .din(new_Jinkela_wire_4043),
        .dout(new_Jinkela_wire_4044)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    bfr new_Jinkela_buffer_2721 (
        .din(new_Jinkela_wire_4010),
        .dout(new_Jinkela_wire_4011)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_2750 (
        .din(new_Jinkela_wire_4058),
        .dout(new_Jinkela_wire_4059)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_2722 (
        .din(new_Jinkela_wire_4011),
        .dout(new_Jinkela_wire_4012)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_2742 (
        .din(new_Jinkela_wire_4044),
        .dout(new_Jinkela_wire_4045)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    bfr new_Jinkela_buffer_2723 (
        .din(new_Jinkela_wire_4012),
        .dout(new_Jinkela_wire_4013)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_617),
        .dout(new_Jinkela_wire_618)
    );

    bfr new_Jinkela_buffer_2796 (
        .din(_1161_),
        .dout(new_Jinkela_wire_4109)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_2724 (
        .din(new_Jinkela_wire_4013),
        .dout(new_Jinkela_wire_4014)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_618),
        .dout(new_Jinkela_wire_619)
    );

    bfr new_Jinkela_buffer_2743 (
        .din(new_Jinkela_wire_4045),
        .dout(new_Jinkela_wire_4046)
    );

    bfr new_Jinkela_buffer_2725 (
        .din(new_Jinkela_wire_4014),
        .dout(new_Jinkela_wire_4015)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_619),
        .dout(new_Jinkela_wire_620)
    );

    bfr new_Jinkela_buffer_2751 (
        .din(new_Jinkela_wire_4059),
        .dout(new_Jinkela_wire_4060)
    );

    bfr new_Jinkela_buffer_2726 (
        .din(new_Jinkela_wire_4015),
        .dout(new_Jinkela_wire_4016)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_620),
        .dout(new_Jinkela_wire_621)
    );

    bfr new_Jinkela_buffer_2744 (
        .din(new_Jinkela_wire_4046),
        .dout(new_Jinkela_wire_4047)
    );

    spl2 new_Jinkela_splitter_136 (
        .a(new_Jinkela_wire_716),
        .b(new_Jinkela_wire_717),
        .c(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_2727 (
        .din(new_Jinkela_wire_4016),
        .dout(new_Jinkela_wire_4017)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    bfr new_Jinkela_buffer_327 (
        .din(G14),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_2768 (
        .din(new_Jinkela_wire_4080),
        .dout(new_Jinkela_wire_4081)
    );

    bfr new_Jinkela_buffer_2799 (
        .din(_0270_),
        .dout(new_Jinkela_wire_4114)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_2728 (
        .din(new_Jinkela_wire_4017),
        .dout(new_Jinkela_wire_4018)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(G150),
        .b(new_Jinkela_wire_729),
        .c(new_Jinkela_wire_730)
    );

    bfr new_Jinkela_buffer_2745 (
        .din(new_Jinkela_wire_4047),
        .dout(new_Jinkela_wire_4048)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_2729 (
        .din(new_Jinkela_wire_4018),
        .dout(new_Jinkela_wire_4019)
    );

    bfr new_Jinkela_buffer_5460 (
        .din(new_Jinkela_wire_7392),
        .dout(new_Jinkela_wire_7393)
    );

    bfr new_Jinkela_buffer_5394 (
        .din(new_Jinkela_wire_7326),
        .dout(new_Jinkela_wire_7327)
    );

    bfr new_Jinkela_buffer_5425 (
        .din(new_Jinkela_wire_7357),
        .dout(new_Jinkela_wire_7358)
    );

    bfr new_Jinkela_buffer_5395 (
        .din(new_Jinkela_wire_7327),
        .dout(new_Jinkela_wire_7328)
    );

    bfr new_Jinkela_buffer_5441 (
        .din(new_Jinkela_wire_7373),
        .dout(new_Jinkela_wire_7374)
    );

    bfr new_Jinkela_buffer_5396 (
        .din(new_Jinkela_wire_7328),
        .dout(new_Jinkela_wire_7329)
    );

    bfr new_Jinkela_buffer_5426 (
        .din(new_Jinkela_wire_7358),
        .dout(new_Jinkela_wire_7359)
    );

    bfr new_Jinkela_buffer_5397 (
        .din(new_Jinkela_wire_7329),
        .dout(new_Jinkela_wire_7330)
    );

    spl2 new_Jinkela_splitter_745 (
        .a(new_net_12),
        .b(new_Jinkela_wire_7433),
        .c(new_Jinkela_wire_7435)
    );

    bfr new_Jinkela_buffer_5523 (
        .din(_0264_),
        .dout(new_Jinkela_wire_7462)
    );

    bfr new_Jinkela_buffer_5398 (
        .din(new_Jinkela_wire_7330),
        .dout(new_Jinkela_wire_7331)
    );

    bfr new_Jinkela_buffer_5427 (
        .din(new_Jinkela_wire_7359),
        .dout(new_Jinkela_wire_7360)
    );

    bfr new_Jinkela_buffer_5399 (
        .din(new_Jinkela_wire_7331),
        .dout(new_Jinkela_wire_7332)
    );

    bfr new_Jinkela_buffer_5442 (
        .din(new_Jinkela_wire_7374),
        .dout(new_Jinkela_wire_7375)
    );

    bfr new_Jinkela_buffer_5400 (
        .din(new_Jinkela_wire_7332),
        .dout(new_Jinkela_wire_7333)
    );

    bfr new_Jinkela_buffer_5428 (
        .din(new_Jinkela_wire_7360),
        .dout(new_Jinkela_wire_7361)
    );

    bfr new_Jinkela_buffer_5401 (
        .din(new_Jinkela_wire_7333),
        .dout(new_Jinkela_wire_7334)
    );

    bfr new_Jinkela_buffer_5461 (
        .din(new_Jinkela_wire_7393),
        .dout(new_Jinkela_wire_7394)
    );

    bfr new_Jinkela_buffer_5402 (
        .din(new_Jinkela_wire_7334),
        .dout(new_Jinkela_wire_7335)
    );

    bfr new_Jinkela_buffer_5429 (
        .din(new_Jinkela_wire_7361),
        .dout(new_Jinkela_wire_7362)
    );

    bfr new_Jinkela_buffer_5403 (
        .din(new_Jinkela_wire_7335),
        .dout(new_Jinkela_wire_7336)
    );

    bfr new_Jinkela_buffer_5443 (
        .din(new_Jinkela_wire_7375),
        .dout(new_Jinkela_wire_7376)
    );

    bfr new_Jinkela_buffer_5404 (
        .din(new_Jinkela_wire_7336),
        .dout(new_Jinkela_wire_7337)
    );

    bfr new_Jinkela_buffer_5430 (
        .din(new_Jinkela_wire_7362),
        .dout(new_Jinkela_wire_7363)
    );

    bfr new_Jinkela_buffer_5405 (
        .din(new_Jinkela_wire_7337),
        .dout(new_Jinkela_wire_7338)
    );

    bfr new_Jinkela_buffer_5406 (
        .din(new_Jinkela_wire_7338),
        .dout(new_Jinkela_wire_7339)
    );

    bfr new_Jinkela_buffer_5431 (
        .din(new_Jinkela_wire_7363),
        .dout(new_Jinkela_wire_7364)
    );

    bfr new_Jinkela_buffer_5407 (
        .din(new_Jinkela_wire_7339),
        .dout(new_Jinkela_wire_7340)
    );

    bfr new_Jinkela_buffer_5444 (
        .din(new_Jinkela_wire_7376),
        .dout(new_Jinkela_wire_7377)
    );

    bfr new_Jinkela_buffer_5408 (
        .din(new_Jinkela_wire_7340),
        .dout(new_Jinkela_wire_7341)
    );

    bfr new_Jinkela_buffer_5432 (
        .din(new_Jinkela_wire_7364),
        .dout(new_Jinkela_wire_7365)
    );

    bfr new_Jinkela_buffer_5409 (
        .din(new_Jinkela_wire_7341),
        .dout(new_Jinkela_wire_7342)
    );

    bfr new_Jinkela_buffer_5462 (
        .din(new_Jinkela_wire_7394),
        .dout(new_Jinkela_wire_7395)
    );

    bfr new_Jinkela_buffer_5410 (
        .din(new_Jinkela_wire_7342),
        .dout(new_Jinkela_wire_7343)
    );

    bfr new_Jinkela_buffer_5433 (
        .din(new_Jinkela_wire_7365),
        .dout(new_Jinkela_wire_7366)
    );

    bfr new_Jinkela_buffer_5411 (
        .din(new_Jinkela_wire_7343),
        .dout(new_Jinkela_wire_7344)
    );

    bfr new_Jinkela_buffer_5445 (
        .din(new_Jinkela_wire_7377),
        .dout(new_Jinkela_wire_7378)
    );

    bfr new_Jinkela_buffer_5412 (
        .din(new_Jinkela_wire_7344),
        .dout(new_Jinkela_wire_7345)
    );

    bfr new_Jinkela_buffer_5434 (
        .din(new_Jinkela_wire_7366),
        .dout(new_Jinkela_wire_7367)
    );

    bfr new_Jinkela_buffer_5413 (
        .din(new_Jinkela_wire_7345),
        .dout(new_Jinkela_wire_7346)
    );

    spl4L new_Jinkela_splitter_746 (
        .a(new_Jinkela_wire_7435),
        .d(new_Jinkela_wire_7436),
        .e(new_Jinkela_wire_7437),
        .b(new_Jinkela_wire_7438),
        .c(new_Jinkela_wire_7439)
    );

    bfr new_Jinkela_buffer_5414 (
        .din(new_Jinkela_wire_7346),
        .dout(new_Jinkela_wire_7347)
    );

    and_ii _1949_ (
        .a(_1237_),
        .b(_1236_),
        .c(_1238_)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_2602),
        .dout(new_Jinkela_wire_2603)
    );

    bfr new_Jinkela_buffer_4489 (
        .din(new_Jinkela_wire_6158),
        .dout(new_Jinkela_wire_6159)
    );

    or_bi _1950_ (
        .a(new_Jinkela_wire_3747),
        .b(new_Jinkela_wire_3103),
        .c(_1239_)
    );

    bfr new_Jinkela_buffer_1622 (
        .din(new_Jinkela_wire_2633),
        .dout(new_Jinkela_wire_2634)
    );

    bfr new_Jinkela_buffer_4536 (
        .din(_0870_),
        .dout(new_Jinkela_wire_6212)
    );

    bfr new_Jinkela_buffer_4518 (
        .din(new_Jinkela_wire_6193),
        .dout(new_Jinkela_wire_6194)
    );

    and_bi _1951_ (
        .a(new_Jinkela_wire_3748),
        .b(new_Jinkela_wire_3104),
        .c(_1240_)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_2603),
        .dout(new_Jinkela_wire_2604)
    );

    bfr new_Jinkela_buffer_4490 (
        .din(new_Jinkela_wire_6159),
        .dout(new_Jinkela_wire_6160)
    );

    and_bi _1952_ (
        .a(_1239_),
        .b(_1240_),
        .c(_1241_)
    );

    bfr new_Jinkela_buffer_1632 (
        .din(new_Jinkela_wire_2643),
        .dout(new_Jinkela_wire_2644)
    );

    bfr new_Jinkela_buffer_4505 (
        .din(new_Jinkela_wire_6174),
        .dout(new_Jinkela_wire_6175)
    );

    or_bb _1953_ (
        .a(new_Jinkela_wire_7196),
        .b(new_Jinkela_wire_3310),
        .c(_1242_)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_2604),
        .dout(new_Jinkela_wire_2605)
    );

    bfr new_Jinkela_buffer_4491 (
        .din(new_Jinkela_wire_6160),
        .dout(new_Jinkela_wire_6161)
    );

    and_bi _1954_ (
        .a(new_Jinkela_wire_5635),
        .b(new_Jinkela_wire_6765),
        .c(_1243_)
    );

    bfr new_Jinkela_buffer_1623 (
        .din(new_Jinkela_wire_2634),
        .dout(new_Jinkela_wire_2635)
    );

    or_bb _1955_ (
        .a(_1243_),
        .b(new_Jinkela_wire_5299),
        .c(_1244_)
    );

    bfr new_Jinkela_buffer_1596 (
        .din(new_Jinkela_wire_2605),
        .dout(new_Jinkela_wire_2606)
    );

    bfr new_Jinkela_buffer_4492 (
        .din(new_Jinkela_wire_6161),
        .dout(new_Jinkela_wire_6162)
    );

    and_bi _1956_ (
        .a(new_Jinkela_wire_7110),
        .b(new_Jinkela_wire_2778),
        .c(_1245_)
    );

    bfr new_Jinkela_buffer_1674 (
        .din(new_Jinkela_wire_2685),
        .dout(new_Jinkela_wire_2686)
    );

    bfr new_Jinkela_buffer_4506 (
        .din(new_Jinkela_wire_6175),
        .dout(new_Jinkela_wire_6176)
    );

    and_bi _1957_ (
        .a(new_Jinkela_wire_2777),
        .b(new_Jinkela_wire_7108),
        .c(_1246_)
    );

    bfr new_Jinkela_buffer_1597 (
        .din(new_Jinkela_wire_2606),
        .dout(new_Jinkela_wire_2607)
    );

    bfr new_Jinkela_buffer_4493 (
        .din(new_Jinkela_wire_6162),
        .dout(new_Jinkela_wire_6163)
    );

    and_ii _1958_ (
        .a(_1246_),
        .b(_1245_),
        .c(_1247_)
    );

    bfr new_Jinkela_buffer_1624 (
        .din(new_Jinkela_wire_2635),
        .dout(new_Jinkela_wire_2636)
    );

    bfr new_Jinkela_buffer_4519 (
        .din(new_Jinkela_wire_6194),
        .dout(new_Jinkela_wire_6195)
    );

    or_bb _1959_ (
        .a(new_Jinkela_wire_7593),
        .b(new_Jinkela_wire_2263),
        .c(_0000_)
    );

    bfr new_Jinkela_buffer_1598 (
        .din(new_Jinkela_wire_2607),
        .dout(new_Jinkela_wire_2608)
    );

    bfr new_Jinkela_buffer_4494 (
        .din(new_Jinkela_wire_6163),
        .dout(new_Jinkela_wire_6164)
    );

    and_bb _1960_ (
        .a(new_Jinkela_wire_7594),
        .b(new_Jinkela_wire_2264),
        .c(_0001_)
    );

    bfr new_Jinkela_buffer_1633 (
        .din(new_Jinkela_wire_2644),
        .dout(new_Jinkela_wire_2645)
    );

    bfr new_Jinkela_buffer_4507 (
        .din(new_Jinkela_wire_6176),
        .dout(new_Jinkela_wire_6177)
    );

    and_bi _1961_ (
        .a(_0000_),
        .b(_0001_),
        .c(_0002_)
    );

    bfr new_Jinkela_buffer_1599 (
        .din(new_Jinkela_wire_2608),
        .dout(new_Jinkela_wire_2609)
    );

    bfr new_Jinkela_buffer_4495 (
        .din(new_Jinkela_wire_6164),
        .dout(new_Jinkela_wire_6165)
    );

    and_bi _1962_ (
        .a(new_Jinkela_wire_3309),
        .b(new_Jinkela_wire_2939),
        .c(_0003_)
    );

    bfr new_Jinkela_buffer_1625 (
        .din(new_Jinkela_wire_2636),
        .dout(new_Jinkela_wire_2637)
    );

    bfr new_Jinkela_buffer_4521 (
        .din(new_Jinkela_wire_6196),
        .dout(new_Jinkela_wire_6197)
    );

    and_bi _1963_ (
        .a(_1242_),
        .b(_0003_),
        .c(_0004_)
    );

    bfr new_Jinkela_buffer_1600 (
        .din(new_Jinkela_wire_2609),
        .dout(new_Jinkela_wire_2610)
    );

    bfr new_Jinkela_buffer_4496 (
        .din(new_Jinkela_wire_6165),
        .dout(new_Jinkela_wire_6166)
    );

    and_bi _1964_ (
        .a(new_Jinkela_wire_7239),
        .b(new_Jinkela_wire_5824),
        .c(_0005_)
    );

    bfr new_Jinkela_buffer_1644 (
        .din(new_Jinkela_wire_2655),
        .dout(new_Jinkela_wire_2656)
    );

    bfr new_Jinkela_buffer_4508 (
        .din(new_Jinkela_wire_6177),
        .dout(new_Jinkela_wire_6178)
    );

    and_bi _1965_ (
        .a(new_Jinkela_wire_3832),
        .b(new_Jinkela_wire_7236),
        .c(_0006_)
    );

    bfr new_Jinkela_buffer_1601 (
        .din(new_Jinkela_wire_2610),
        .dout(new_Jinkela_wire_2611)
    );

    bfr new_Jinkela_buffer_4497 (
        .din(new_Jinkela_wire_6166),
        .dout(new_Jinkela_wire_6167)
    );

    and_ii _1966_ (
        .a(_0006_),
        .b(_0005_),
        .c(_0007_)
    );

    bfr new_Jinkela_buffer_1626 (
        .din(new_Jinkela_wire_2637),
        .dout(new_Jinkela_wire_2638)
    );

    spl2 new_Jinkela_splitter_642 (
        .a(_0599_),
        .b(new_Jinkela_wire_6225),
        .c(new_Jinkela_wire_6226)
    );

    bfr new_Jinkela_buffer_4551 (
        .din(_0147_),
        .dout(new_Jinkela_wire_6229)
    );

    or_bi _1967_ (
        .a(new_Jinkela_wire_6020),
        .b(new_Jinkela_wire_1123),
        .c(_0008_)
    );

    bfr new_Jinkela_buffer_1602 (
        .din(new_Jinkela_wire_2611),
        .dout(new_Jinkela_wire_2612)
    );

    bfr new_Jinkela_buffer_4509 (
        .din(new_Jinkela_wire_6178),
        .dout(new_Jinkela_wire_6179)
    );

    and_bi _1968_ (
        .a(new_Jinkela_wire_4531),
        .b(new_Jinkela_wire_6283),
        .c(_0009_)
    );

    bfr new_Jinkela_buffer_1634 (
        .din(new_Jinkela_wire_2645),
        .dout(new_Jinkela_wire_2646)
    );

    bfr new_Jinkela_buffer_4522 (
        .din(new_Jinkela_wire_6197),
        .dout(new_Jinkela_wire_6198)
    );

    and_ii _1969_ (
        .a(new_Jinkela_wire_4529),
        .b(new_Jinkela_wire_1126),
        .c(_0010_)
    );

    bfr new_Jinkela_buffer_1603 (
        .din(new_Jinkela_wire_2612),
        .dout(new_Jinkela_wire_2613)
    );

    bfr new_Jinkela_buffer_4510 (
        .din(new_Jinkela_wire_6179),
        .dout(new_Jinkela_wire_6180)
    );

    or_bb _1970_ (
        .a(new_Jinkela_wire_7935),
        .b(new_Jinkela_wire_5903),
        .c(_0011_)
    );

    spl4L new_Jinkela_splitter_379 (
        .a(_0580_),
        .d(new_Jinkela_wire_2765),
        .e(new_Jinkela_wire_2766),
        .b(new_Jinkela_wire_2767),
        .c(new_Jinkela_wire_2771)
    );

    bfr new_Jinkela_buffer_4537 (
        .din(new_Jinkela_wire_6212),
        .dout(new_Jinkela_wire_6213)
    );

    bfr new_Jinkela_buffer_1754 (
        .din(_0642_),
        .dout(new_Jinkela_wire_2779)
    );

    or_bb _1971_ (
        .a(_0011_),
        .b(new_Jinkela_wire_7784),
        .c(_0012_)
    );

    bfr new_Jinkela_buffer_1604 (
        .din(new_Jinkela_wire_2613),
        .dout(new_Jinkela_wire_2614)
    );

    bfr new_Jinkela_buffer_4511 (
        .din(new_Jinkela_wire_6180),
        .dout(new_Jinkela_wire_6181)
    );

    or_bb _1972_ (
        .a(new_Jinkela_wire_4346),
        .b(new_Jinkela_wire_2808),
        .c(_0013_)
    );

    bfr new_Jinkela_buffer_1635 (
        .din(new_Jinkela_wire_2646),
        .dout(new_Jinkela_wire_2647)
    );

    bfr new_Jinkela_buffer_4523 (
        .din(new_Jinkela_wire_6198),
        .dout(new_Jinkela_wire_6199)
    );

    and_bb _1973_ (
        .a(new_Jinkela_wire_4348),
        .b(new_Jinkela_wire_2807),
        .c(_0014_)
    );

    bfr new_Jinkela_buffer_1605 (
        .din(new_Jinkela_wire_2614),
        .dout(new_Jinkela_wire_2615)
    );

    bfr new_Jinkela_buffer_4512 (
        .din(new_Jinkela_wire_6181),
        .dout(new_Jinkela_wire_6182)
    );

    and_bi _1974_ (
        .a(_0013_),
        .b(_0014_),
        .c(_0015_)
    );

    bfr new_Jinkela_buffer_1645 (
        .din(new_Jinkela_wire_2656),
        .dout(new_Jinkela_wire_2657)
    );

    bfr new_Jinkela_buffer_4549 (
        .din(new_Jinkela_wire_6226),
        .dout(new_Jinkela_wire_6227)
    );

    or_bb _1975_ (
        .a(new_Jinkela_wire_5731),
        .b(new_Jinkela_wire_6752),
        .c(_0016_)
    );

    bfr new_Jinkela_buffer_1606 (
        .din(new_Jinkela_wire_2615),
        .dout(new_Jinkela_wire_2616)
    );

    bfr new_Jinkela_buffer_4513 (
        .din(new_Jinkela_wire_6182),
        .dout(new_Jinkela_wire_6183)
    );

    and_bb _1976_ (
        .a(new_Jinkela_wire_5732),
        .b(new_Jinkela_wire_6753),
        .c(_0017_)
    );

    bfr new_Jinkela_buffer_1636 (
        .din(new_Jinkela_wire_2647),
        .dout(new_Jinkela_wire_2648)
    );

    bfr new_Jinkela_buffer_4524 (
        .din(new_Jinkela_wire_6199),
        .dout(new_Jinkela_wire_6200)
    );

    or_bi _1977_ (
        .a(_0017_),
        .b(_0016_),
        .c(_0018_)
    );

    bfr new_Jinkela_buffer_1607 (
        .din(new_Jinkela_wire_2616),
        .dout(new_Jinkela_wire_2617)
    );

    bfr new_Jinkela_buffer_4514 (
        .din(new_Jinkela_wire_6183),
        .dout(new_Jinkela_wire_6184)
    );

    or_bb _1978_ (
        .a(new_Jinkela_wire_2209),
        .b(new_Jinkela_wire_5283),
        .c(_0019_)
    );

    bfr new_Jinkela_buffer_1675 (
        .din(new_Jinkela_wire_2686),
        .dout(new_Jinkela_wire_2687)
    );

    bfr new_Jinkela_buffer_4538 (
        .din(new_Jinkela_wire_6213),
        .dout(new_Jinkela_wire_6214)
    );

    and_bi _1979_ (
        .a(new_Jinkela_wire_2210),
        .b(new_Jinkela_wire_5695),
        .c(_0020_)
    );

    bfr new_Jinkela_buffer_1608 (
        .din(new_Jinkela_wire_2617),
        .dout(new_Jinkela_wire_2618)
    );

    bfr new_Jinkela_buffer_4525 (
        .din(new_Jinkela_wire_6200),
        .dout(new_Jinkela_wire_6201)
    );

    and_bi _1980_ (
        .a(_0019_),
        .b(_0020_),
        .c(_0021_)
    );

    bfr new_Jinkela_buffer_1637 (
        .din(new_Jinkela_wire_2648),
        .dout(new_Jinkela_wire_2649)
    );

    and_bi _1981_ (
        .a(new_Jinkela_wire_6072),
        .b(new_Jinkela_wire_5435),
        .c(_0022_)
    );

    bfr new_Jinkela_buffer_1609 (
        .din(new_Jinkela_wire_2618),
        .dout(new_Jinkela_wire_2619)
    );

    bfr new_Jinkela_buffer_4526 (
        .din(new_Jinkela_wire_6201),
        .dout(new_Jinkela_wire_6202)
    );

    and_bi _1982_ (
        .a(new_Jinkela_wire_5436),
        .b(new_Jinkela_wire_6073),
        .c(_0023_)
    );

    bfr new_Jinkela_buffer_1646 (
        .din(new_Jinkela_wire_2657),
        .dout(new_Jinkela_wire_2658)
    );

    bfr new_Jinkela_buffer_4539 (
        .din(new_Jinkela_wire_6214),
        .dout(new_Jinkela_wire_6215)
    );

    or_bb _1983_ (
        .a(_0023_),
        .b(_0022_),
        .c(_0024_)
    );

    bfr new_Jinkela_buffer_1610 (
        .din(new_Jinkela_wire_2619),
        .dout(new_Jinkela_wire_2620)
    );

    bfr new_Jinkela_buffer_4527 (
        .din(new_Jinkela_wire_6202),
        .dout(new_Jinkela_wire_6203)
    );

    and_ii _1984_ (
        .a(new_Jinkela_wire_5196),
        .b(new_Jinkela_wire_2197),
        .c(_0025_)
    );

    bfr new_Jinkela_buffer_1638 (
        .din(new_Jinkela_wire_2649),
        .dout(new_Jinkela_wire_2650)
    );

    bfr new_Jinkela_buffer_4552 (
        .din(_0228_),
        .dout(new_Jinkela_wire_6232)
    );

    and_bb _1985_ (
        .a(new_Jinkela_wire_5197),
        .b(new_Jinkela_wire_2198),
        .c(_0026_)
    );

    bfr new_Jinkela_buffer_1611 (
        .din(new_Jinkela_wire_2620),
        .dout(new_Jinkela_wire_2621)
    );

    bfr new_Jinkela_buffer_4528 (
        .din(new_Jinkela_wire_6203),
        .dout(new_Jinkela_wire_6204)
    );

    or_bb _1986_ (
        .a(_0026_),
        .b(new_Jinkela_wire_1090),
        .c(_0027_)
    );

    bfr new_Jinkela_buffer_1714 (
        .din(new_Jinkela_wire_2725),
        .dout(new_Jinkela_wire_2726)
    );

    bfr new_Jinkela_buffer_4540 (
        .din(new_Jinkela_wire_6215),
        .dout(new_Jinkela_wire_6216)
    );

    or_bb _1987_ (
        .a(_0027_),
        .b(new_Jinkela_wire_5433),
        .c(_0028_)
    );

    bfr new_Jinkela_buffer_1639 (
        .din(new_Jinkela_wire_2650),
        .dout(new_Jinkela_wire_2651)
    );

    bfr new_Jinkela_buffer_4529 (
        .din(new_Jinkela_wire_6204),
        .dout(new_Jinkela_wire_6205)
    );

    and_bi _1988_ (
        .a(new_Jinkela_wire_1529),
        .b(new_Jinkela_wire_1105),
        .c(_0029_)
    );

    bfr new_Jinkela_buffer_1647 (
        .din(new_Jinkela_wire_2658),
        .dout(new_Jinkela_wire_2659)
    );

    spl2 new_Jinkela_splitter_644 (
        .a(_0941_),
        .b(new_Jinkela_wire_6234),
        .c(new_Jinkela_wire_6235)
    );

    bfr new_Jinkela_buffer_4550 (
        .din(new_Jinkela_wire_6227),
        .dout(new_Jinkela_wire_6228)
    );

    and_bi _1989_ (
        .a(new_Jinkela_wire_1102),
        .b(new_Jinkela_wire_49),
        .c(_0030_)
    );

    bfr new_Jinkela_buffer_1640 (
        .din(new_Jinkela_wire_2651),
        .dout(new_Jinkela_wire_2652)
    );

    bfr new_Jinkela_buffer_4530 (
        .din(new_Jinkela_wire_6205),
        .dout(new_Jinkela_wire_6206)
    );

    and_ii _1990_ (
        .a(_0030_),
        .b(_0029_),
        .c(_0031_)
    );

    bfr new_Jinkela_buffer_1676 (
        .din(new_Jinkela_wire_2687),
        .dout(new_Jinkela_wire_2688)
    );

    bfr new_Jinkela_buffer_4541 (
        .din(new_Jinkela_wire_6216),
        .dout(new_Jinkela_wire_6217)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_5435 (
        .din(new_Jinkela_wire_7367),
        .dout(new_Jinkela_wire_7368)
    );

    bfr new_Jinkela_buffer_5415 (
        .din(new_Jinkela_wire_7347),
        .dout(new_Jinkela_wire_7348)
    );

    spl4L new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_872),
        .d(new_Jinkela_wire_873),
        .e(new_Jinkela_wire_874),
        .b(new_Jinkela_wire_875),
        .c(new_Jinkela_wire_876)
    );

    spl2 new_Jinkela_splitter_174 (
        .a(new_Jinkela_wire_891),
        .b(new_Jinkela_wire_892),
        .c(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_5446 (
        .din(new_Jinkela_wire_7378),
        .dout(new_Jinkela_wire_7379)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_5416 (
        .din(new_Jinkela_wire_7348),
        .dout(new_Jinkela_wire_7349)
    );

    spl4L new_Jinkela_splitter_172 (
        .a(new_Jinkela_wire_882),
        .d(new_Jinkela_wire_883),
        .e(new_Jinkela_wire_884),
        .b(new_Jinkela_wire_885),
        .c(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_5436 (
        .din(new_Jinkela_wire_7368),
        .dout(new_Jinkela_wire_7369)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_5417 (
        .din(new_Jinkela_wire_7349),
        .dout(new_Jinkela_wire_7350)
    );

    spl4L new_Jinkela_splitter_173 (
        .a(new_Jinkela_wire_887),
        .d(new_Jinkela_wire_888),
        .e(new_Jinkela_wire_889),
        .b(new_Jinkela_wire_890),
        .c(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_5463 (
        .din(new_Jinkela_wire_7395),
        .dout(new_Jinkela_wire_7396)
    );

    spl2 new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_815),
        .b(new_Jinkela_wire_816),
        .c(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_5418 (
        .din(new_Jinkela_wire_7350),
        .dout(new_Jinkela_wire_7351)
    );

    spl2 new_Jinkela_splitter_155 (
        .a(new_Jinkela_wire_817),
        .b(new_Jinkela_wire_818),
        .c(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_5437 (
        .din(new_Jinkela_wire_7369),
        .dout(new_Jinkela_wire_7370)
    );

    bfr new_Jinkela_buffer_442 (
        .din(G146),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_5447 (
        .din(new_Jinkela_wire_7379),
        .dout(new_Jinkela_wire_7380)
    );

    spl2 new_Jinkela_splitter_156 (
        .a(new_Jinkela_wire_819),
        .b(new_Jinkela_wire_820),
        .c(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_5500 (
        .din(new_Jinkela_wire_7433),
        .dout(new_Jinkela_wire_7434)
    );

    bfr new_Jinkela_buffer_446 (
        .din(G32),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_5448 (
        .din(new_Jinkela_wire_7380),
        .dout(new_Jinkela_wire_7381)
    );

    spl3L new_Jinkela_splitter_157 (
        .a(new_Jinkela_wire_821),
        .d(new_Jinkela_wire_822),
        .b(new_Jinkela_wire_823),
        .c(new_Jinkela_wire_824)
    );

    bfr new_Jinkela_buffer_5464 (
        .din(new_Jinkela_wire_7396),
        .dout(new_Jinkela_wire_7397)
    );

    bfr new_Jinkela_buffer_450 (
        .din(G85),
        .dout(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_5449 (
        .din(new_Jinkela_wire_7381),
        .dout(new_Jinkela_wire_7382)
    );

    bfr new_Jinkela_buffer_453 (
        .din(G47),
        .dout(new_Jinkela_wire_963)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_5526 (
        .din(new_net_2405),
        .dout(new_Jinkela_wire_7465)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_5450 (
        .din(new_Jinkela_wire_7382),
        .dout(new_Jinkela_wire_7383)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_5465 (
        .din(new_Jinkela_wire_7397),
        .dout(new_Jinkela_wire_7398)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_5451 (
        .din(new_Jinkela_wire_7383),
        .dout(new_Jinkela_wire_7384)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_5501 (
        .din(new_Jinkela_wire_7439),
        .dout(new_Jinkela_wire_7440)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_5452 (
        .din(new_Jinkela_wire_7384),
        .dout(new_Jinkela_wire_7385)
    );

    or_bb _2464_ (
        .a(_0457_),
        .b(new_Jinkela_wire_3521),
        .c(_0458_)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_5466 (
        .din(new_Jinkela_wire_7398),
        .dout(new_Jinkela_wire_7399)
    );

    and_bi _2463_ (
        .a(new_Jinkela_wire_6794),
        .b(new_Jinkela_wire_1479),
        .c(_0457_)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_5453 (
        .din(new_Jinkela_wire_7385),
        .dout(new_Jinkela_wire_7386)
    );

    bfr new_Jinkela_buffer_5524 (
        .din(new_Jinkela_wire_7462),
        .dout(new_Jinkela_wire_7463)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_5454 (
        .din(new_Jinkela_wire_7386),
        .dout(new_Jinkela_wire_7387)
    );

    or_ii _2462_ (
        .a(new_Jinkela_wire_5778),
        .b(new_Jinkela_wire_1477),
        .c(_0456_)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_5467 (
        .din(new_Jinkela_wire_7399),
        .dout(new_Jinkela_wire_7400)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_5455 (
        .din(new_Jinkela_wire_7387),
        .dout(new_Jinkela_wire_7388)
    );

    spl3L new_Jinkela_splitter_747 (
        .a(_0952_),
        .d(new_Jinkela_wire_7469),
        .b(new_Jinkela_wire_7470),
        .c(new_Jinkela_wire_7471)
    );

    bfr new_Jinkela_buffer_5530 (
        .din(_0476_),
        .dout(new_Jinkela_wire_7472)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_5456 (
        .din(new_Jinkela_wire_7388),
        .dout(new_Jinkela_wire_7389)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_5468 (
        .din(new_Jinkela_wire_7400),
        .dout(new_Jinkela_wire_7401)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_5457 (
        .din(new_Jinkela_wire_7389),
        .dout(new_Jinkela_wire_7390)
    );

    bfr new_Jinkela_buffer_5502 (
        .din(new_Jinkela_wire_7440),
        .dout(new_Jinkela_wire_7441)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_5458 (
        .din(new_Jinkela_wire_7390),
        .dout(new_Jinkela_wire_7391)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_5469 (
        .din(new_Jinkela_wire_7401),
        .dout(new_Jinkela_wire_7402)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_5525 (
        .din(new_Jinkela_wire_7463),
        .dout(new_Jinkela_wire_7464)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_955),
        .dout(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_5470 (
        .din(new_Jinkela_wire_7402),
        .dout(new_Jinkela_wire_7403)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_5503 (
        .din(new_Jinkela_wire_7441),
        .dout(new_Jinkela_wire_7442)
    );

    spl3L new_Jinkela_splitter_177 (
        .a(new_Jinkela_wire_948),
        .d(new_Jinkela_wire_949),
        .b(new_Jinkela_wire_950),
        .c(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_5471 (
        .din(new_Jinkela_wire_7403),
        .dout(new_Jinkela_wire_7404)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_5527 (
        .din(new_Jinkela_wire_7465),
        .dout(new_Jinkela_wire_7466)
    );

    bfr new_Jinkela_buffer_458 (
        .din(G95),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_5472 (
        .din(new_Jinkela_wire_7404),
        .dout(new_Jinkela_wire_7405)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_5504 (
        .din(new_Jinkela_wire_7442),
        .dout(new_Jinkela_wire_7443)
    );

    spl2 new_Jinkela_splitter_178 (
        .a(new_Jinkela_wire_951),
        .b(new_Jinkela_wire_952),
        .c(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_5473 (
        .din(new_Jinkela_wire_7405),
        .dout(new_Jinkela_wire_7406)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_3409 (
        .din(new_Jinkela_wire_4802),
        .dout(new_Jinkela_wire_4803)
    );

    bfr new_Jinkela_buffer_4459 (
        .din(new_Jinkela_wire_6109),
        .dout(new_Jinkela_wire_6110)
    );

    bfr new_Jinkela_buffer_3359 (
        .din(new_Jinkela_wire_4750),
        .dout(new_Jinkela_wire_4751)
    );

    bfr new_Jinkela_buffer_3386 (
        .din(new_Jinkela_wire_4779),
        .dout(new_Jinkela_wire_4780)
    );

    bfr new_Jinkela_buffer_4470 (
        .din(new_Jinkela_wire_6120),
        .dout(new_Jinkela_wire_6121)
    );

    bfr new_Jinkela_buffer_4460 (
        .din(new_Jinkela_wire_6110),
        .dout(new_Jinkela_wire_6111)
    );

    bfr new_Jinkela_buffer_3360 (
        .din(new_Jinkela_wire_4751),
        .dout(new_Jinkela_wire_4752)
    );

    bfr new_Jinkela_buffer_4461 (
        .din(new_Jinkela_wire_6111),
        .dout(new_Jinkela_wire_6112)
    );

    bfr new_Jinkela_buffer_3435 (
        .din(new_Jinkela_wire_4857),
        .dout(new_Jinkela_wire_4858)
    );

    bfr new_Jinkela_buffer_3361 (
        .din(new_Jinkela_wire_4752),
        .dout(new_Jinkela_wire_4753)
    );

    bfr new_Jinkela_buffer_3387 (
        .din(new_Jinkela_wire_4780),
        .dout(new_Jinkela_wire_4781)
    );

    bfr new_Jinkela_buffer_4473 (
        .din(new_Jinkela_wire_6138),
        .dout(new_Jinkela_wire_6139)
    );

    bfr new_Jinkela_buffer_4462 (
        .din(new_Jinkela_wire_6112),
        .dout(new_Jinkela_wire_6113)
    );

    bfr new_Jinkela_buffer_3362 (
        .din(new_Jinkela_wire_4753),
        .dout(new_Jinkela_wire_4754)
    );

    spl2 new_Jinkela_splitter_636 (
        .a(new_Jinkela_wire_6125),
        .b(new_Jinkela_wire_6126),
        .c(new_Jinkela_wire_6127)
    );

    bfr new_Jinkela_buffer_3410 (
        .din(new_Jinkela_wire_4803),
        .dout(new_Jinkela_wire_4804)
    );

    bfr new_Jinkela_buffer_4463 (
        .din(new_Jinkela_wire_6113),
        .dout(new_Jinkela_wire_6114)
    );

    bfr new_Jinkela_buffer_3388 (
        .din(new_Jinkela_wire_4781),
        .dout(new_Jinkela_wire_4782)
    );

    bfr new_Jinkela_buffer_4476 (
        .din(new_net_2373),
        .dout(new_Jinkela_wire_6146)
    );

    spl4L new_Jinkela_splitter_637 (
        .a(new_Jinkela_wire_6128),
        .d(new_Jinkela_wire_6129),
        .e(new_Jinkela_wire_6130),
        .b(new_Jinkela_wire_6131),
        .c(new_Jinkela_wire_6132)
    );

    bfr new_Jinkela_buffer_4464 (
        .din(new_Jinkela_wire_6114),
        .dout(new_Jinkela_wire_6115)
    );

    bfr new_Jinkela_buffer_3389 (
        .din(new_Jinkela_wire_4782),
        .dout(new_Jinkela_wire_4783)
    );

    bfr new_Jinkela_buffer_3411 (
        .din(new_Jinkela_wire_4804),
        .dout(new_Jinkela_wire_4805)
    );

    spl4L new_Jinkela_splitter_638 (
        .a(new_Jinkela_wire_6133),
        .d(new_Jinkela_wire_6134),
        .e(new_Jinkela_wire_6135),
        .b(new_Jinkela_wire_6136),
        .c(new_Jinkela_wire_6137)
    );

    bfr new_Jinkela_buffer_4465 (
        .din(new_Jinkela_wire_6115),
        .dout(new_Jinkela_wire_6116)
    );

    bfr new_Jinkela_buffer_3390 (
        .din(new_Jinkela_wire_4783),
        .dout(new_Jinkela_wire_4784)
    );

    bfr new_Jinkela_buffer_3436 (
        .din(new_Jinkela_wire_4858),
        .dout(new_Jinkela_wire_4859)
    );

    bfr new_Jinkela_buffer_4477 (
        .din(new_Jinkela_wire_6146),
        .dout(new_Jinkela_wire_6147)
    );

    bfr new_Jinkela_buffer_3437 (
        .din(new_Jinkela_wire_4859),
        .dout(new_Jinkela_wire_4860)
    );

    bfr new_Jinkela_buffer_3391 (
        .din(new_Jinkela_wire_4784),
        .dout(new_Jinkela_wire_4785)
    );

    spl4L new_Jinkela_splitter_639 (
        .a(new_Jinkela_wire_6139),
        .d(new_Jinkela_wire_6140),
        .e(new_Jinkela_wire_6141),
        .b(new_Jinkela_wire_6142),
        .c(new_Jinkela_wire_6143)
    );

    bfr new_Jinkela_buffer_3412 (
        .din(new_Jinkela_wire_4805),
        .dout(new_Jinkela_wire_4806)
    );

    bfr new_Jinkela_buffer_4498 (
        .din(_0451_),
        .dout(new_Jinkela_wire_6168)
    );

    bfr new_Jinkela_buffer_4474 (
        .din(new_Jinkela_wire_6143),
        .dout(new_Jinkela_wire_6144)
    );

    bfr new_Jinkela_buffer_3392 (
        .din(new_Jinkela_wire_4785),
        .dout(new_Jinkela_wire_4786)
    );

    bfr new_Jinkela_buffer_3445 (
        .din(new_net_2397),
        .dout(new_Jinkela_wire_4868)
    );

    bfr new_Jinkela_buffer_4515 (
        .din(_0645_),
        .dout(new_Jinkela_wire_6185)
    );

    spl2 new_Jinkela_splitter_641 (
        .a(_0934_),
        .b(new_Jinkela_wire_6191),
        .c(new_Jinkela_wire_6192)
    );

    bfr new_Jinkela_buffer_3422 (
        .din(new_Jinkela_wire_4817),
        .dout(new_Jinkela_wire_4818)
    );

    bfr new_Jinkela_buffer_3393 (
        .din(new_Jinkela_wire_4786),
        .dout(new_Jinkela_wire_4787)
    );

    bfr new_Jinkela_buffer_4478 (
        .din(new_Jinkela_wire_6147),
        .dout(new_Jinkela_wire_6148)
    );

    bfr new_Jinkela_buffer_4475 (
        .din(new_Jinkela_wire_6144),
        .dout(new_Jinkela_wire_6145)
    );

    bfr new_Jinkela_buffer_3413 (
        .din(new_Jinkela_wire_4806),
        .dout(new_Jinkela_wire_4807)
    );

    bfr new_Jinkela_buffer_3394 (
        .din(new_Jinkela_wire_4787),
        .dout(new_Jinkela_wire_4788)
    );

    bfr new_Jinkela_buffer_4499 (
        .din(new_Jinkela_wire_6168),
        .dout(new_Jinkela_wire_6169)
    );

    bfr new_Jinkela_buffer_4479 (
        .din(new_Jinkela_wire_6148),
        .dout(new_Jinkela_wire_6149)
    );

    spl4L new_Jinkela_splitter_532 (
        .a(new_Jinkela_wire_4819),
        .d(new_Jinkela_wire_4820),
        .e(new_Jinkela_wire_4821),
        .b(new_Jinkela_wire_4822),
        .c(new_Jinkela_wire_4823)
    );

    bfr new_Jinkela_buffer_3395 (
        .din(new_Jinkela_wire_4788),
        .dout(new_Jinkela_wire_4789)
    );

    bfr new_Jinkela_buffer_4516 (
        .din(new_Jinkela_wire_6185),
        .dout(new_Jinkela_wire_6186)
    );

    bfr new_Jinkela_buffer_3414 (
        .din(new_Jinkela_wire_4807),
        .dout(new_Jinkela_wire_4808)
    );

    bfr new_Jinkela_buffer_4480 (
        .din(new_Jinkela_wire_6149),
        .dout(new_Jinkela_wire_6150)
    );

    bfr new_Jinkela_buffer_3396 (
        .din(new_Jinkela_wire_4789),
        .dout(new_Jinkela_wire_4790)
    );

    bfr new_Jinkela_buffer_4500 (
        .din(new_Jinkela_wire_6169),
        .dout(new_Jinkela_wire_6170)
    );

    bfr new_Jinkela_buffer_4481 (
        .din(new_Jinkela_wire_6150),
        .dout(new_Jinkela_wire_6151)
    );

    bfr new_Jinkela_buffer_3397 (
        .din(new_Jinkela_wire_4790),
        .dout(new_Jinkela_wire_4791)
    );

    bfr new_Jinkela_buffer_4517 (
        .din(_0101_),
        .dout(new_Jinkela_wire_6193)
    );

    bfr new_Jinkela_buffer_3415 (
        .din(new_Jinkela_wire_4808),
        .dout(new_Jinkela_wire_4809)
    );

    bfr new_Jinkela_buffer_4482 (
        .din(new_Jinkela_wire_6151),
        .dout(new_Jinkela_wire_6152)
    );

    bfr new_Jinkela_buffer_3398 (
        .din(new_Jinkela_wire_4791),
        .dout(new_Jinkela_wire_4792)
    );

    bfr new_Jinkela_buffer_4501 (
        .din(new_Jinkela_wire_6170),
        .dout(new_Jinkela_wire_6171)
    );

    bfr new_Jinkela_buffer_4483 (
        .din(new_Jinkela_wire_6152),
        .dout(new_Jinkela_wire_6153)
    );

    bfr new_Jinkela_buffer_3399 (
        .din(new_Jinkela_wire_4792),
        .dout(new_Jinkela_wire_4793)
    );

    spl4L new_Jinkela_splitter_640 (
        .a(new_Jinkela_wire_6186),
        .d(new_Jinkela_wire_6187),
        .e(new_Jinkela_wire_6188),
        .b(new_Jinkela_wire_6189),
        .c(new_Jinkela_wire_6190)
    );

    bfr new_Jinkela_buffer_3416 (
        .din(new_Jinkela_wire_4809),
        .dout(new_Jinkela_wire_4810)
    );

    bfr new_Jinkela_buffer_4484 (
        .din(new_Jinkela_wire_6153),
        .dout(new_Jinkela_wire_6154)
    );

    bfr new_Jinkela_buffer_3400 (
        .din(new_Jinkela_wire_4793),
        .dout(new_Jinkela_wire_4794)
    );

    bfr new_Jinkela_buffer_4502 (
        .din(new_Jinkela_wire_6171),
        .dout(new_Jinkela_wire_6172)
    );

    spl3L new_Jinkela_splitter_533 (
        .a(new_Jinkela_wire_4823),
        .d(new_Jinkela_wire_4824),
        .b(new_Jinkela_wire_4825),
        .c(new_Jinkela_wire_4828)
    );

    bfr new_Jinkela_buffer_4485 (
        .din(new_Jinkela_wire_6154),
        .dout(new_Jinkela_wire_6155)
    );

    bfr new_Jinkela_buffer_3401 (
        .din(new_Jinkela_wire_4794),
        .dout(new_Jinkela_wire_4795)
    );

    bfr new_Jinkela_buffer_3417 (
        .din(new_Jinkela_wire_4810),
        .dout(new_Jinkela_wire_4811)
    );

    bfr new_Jinkela_buffer_4486 (
        .din(new_Jinkela_wire_6155),
        .dout(new_Jinkela_wire_6156)
    );

    bfr new_Jinkela_buffer_3423 (
        .din(new_Jinkela_wire_4818),
        .dout(new_Jinkela_wire_4819)
    );

    bfr new_Jinkela_buffer_4503 (
        .din(new_Jinkela_wire_6172),
        .dout(new_Jinkela_wire_6173)
    );

    bfr new_Jinkela_buffer_3418 (
        .din(new_Jinkela_wire_4811),
        .dout(new_Jinkela_wire_4812)
    );

    bfr new_Jinkela_buffer_4487 (
        .din(new_Jinkela_wire_6156),
        .dout(new_Jinkela_wire_6157)
    );

    bfr new_Jinkela_buffer_3443 (
        .din(new_Jinkela_wire_4865),
        .dout(new_Jinkela_wire_4866)
    );

    bfr new_Jinkela_buffer_4520 (
        .din(new_net_2365),
        .dout(new_Jinkela_wire_6196)
    );

    bfr new_Jinkela_buffer_3419 (
        .din(new_Jinkela_wire_4812),
        .dout(new_Jinkela_wire_4813)
    );

    bfr new_Jinkela_buffer_4488 (
        .din(new_Jinkela_wire_6157),
        .dout(new_Jinkela_wire_6158)
    );

    bfr new_Jinkela_buffer_3464 (
        .din(_0700_),
        .dout(new_Jinkela_wire_4887)
    );

    bfr new_Jinkela_buffer_4504 (
        .din(new_Jinkela_wire_6173),
        .dout(new_Jinkela_wire_6174)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(new_Jinkela_wire_2580),
        .dout(new_Jinkela_wire_2581)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_2559),
        .dout(new_Jinkela_wire_2560)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_2560),
        .dout(new_Jinkela_wire_2561)
    );

    bfr new_Jinkela_buffer_1614 (
        .din(new_Jinkela_wire_2625),
        .dout(new_Jinkela_wire_2626)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_2561),
        .dout(new_Jinkela_wire_2562)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(new_Jinkela_wire_2587),
        .dout(new_Jinkela_wire_2588)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_2562),
        .dout(new_Jinkela_wire_2563)
    );

    bfr new_Jinkela_buffer_1628 (
        .din(new_Jinkela_wire_2639),
        .dout(new_Jinkela_wire_2640)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_2563),
        .dout(new_Jinkela_wire_2564)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_2588),
        .dout(new_Jinkela_wire_2589)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_2564),
        .dout(new_Jinkela_wire_2565)
    );

    bfr new_Jinkela_buffer_1615 (
        .din(new_Jinkela_wire_2626),
        .dout(new_Jinkela_wire_2627)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_2565),
        .dout(new_Jinkela_wire_2566)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(new_Jinkela_wire_2589),
        .dout(new_Jinkela_wire_2590)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_2566),
        .dout(new_Jinkela_wire_2567)
    );

    bfr new_Jinkela_buffer_1673 (
        .din(new_net_2465),
        .dout(new_Jinkela_wire_2685)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_2567),
        .dout(new_Jinkela_wire_2568)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_2590),
        .dout(new_Jinkela_wire_2591)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(new_Jinkela_wire_2568),
        .dout(new_Jinkela_wire_2569)
    );

    bfr new_Jinkela_buffer_1616 (
        .din(new_Jinkela_wire_2627),
        .dout(new_Jinkela_wire_2628)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_2591),
        .dout(new_Jinkela_wire_2592)
    );

    bfr new_Jinkela_buffer_1629 (
        .din(new_Jinkela_wire_2640),
        .dout(new_Jinkela_wire_2641)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(new_Jinkela_wire_2592),
        .dout(new_Jinkela_wire_2593)
    );

    bfr new_Jinkela_buffer_1617 (
        .din(new_Jinkela_wire_2628),
        .dout(new_Jinkela_wire_2629)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_Jinkela_wire_2593),
        .dout(new_Jinkela_wire_2594)
    );

    bfr new_Jinkela_buffer_1642 (
        .din(new_Jinkela_wire_2653),
        .dout(new_Jinkela_wire_2654)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_Jinkela_wire_2594),
        .dout(new_Jinkela_wire_2595)
    );

    bfr new_Jinkela_buffer_1618 (
        .din(new_Jinkela_wire_2629),
        .dout(new_Jinkela_wire_2630)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_2595),
        .dout(new_Jinkela_wire_2596)
    );

    bfr new_Jinkela_buffer_1630 (
        .din(new_Jinkela_wire_2641),
        .dout(new_Jinkela_wire_2642)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_2596),
        .dout(new_Jinkela_wire_2597)
    );

    bfr new_Jinkela_buffer_1619 (
        .din(new_Jinkela_wire_2630),
        .dout(new_Jinkela_wire_2631)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_2597),
        .dout(new_Jinkela_wire_2598)
    );

    bfr new_Jinkela_buffer_1713 (
        .din(new_net_2463),
        .dout(new_Jinkela_wire_2725)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(new_Jinkela_wire_2598),
        .dout(new_Jinkela_wire_2599)
    );

    bfr new_Jinkela_buffer_1620 (
        .din(new_Jinkela_wire_2631),
        .dout(new_Jinkela_wire_2632)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(new_Jinkela_wire_2599),
        .dout(new_Jinkela_wire_2600)
    );

    bfr new_Jinkela_buffer_1631 (
        .din(new_Jinkela_wire_2642),
        .dout(new_Jinkela_wire_2643)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(new_Jinkela_wire_2600),
        .dout(new_Jinkela_wire_2601)
    );

    bfr new_Jinkela_buffer_1621 (
        .din(new_Jinkela_wire_2632),
        .dout(new_Jinkela_wire_2633)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_2601),
        .dout(new_Jinkela_wire_2602)
    );

    bfr new_Jinkela_buffer_1643 (
        .din(new_Jinkela_wire_2654),
        .dout(new_Jinkela_wire_2655)
    );

    bfr new_Jinkela_buffer_4696 (
        .din(new_Jinkela_wire_6428),
        .dout(new_Jinkela_wire_6429)
    );

    bfr new_Jinkela_buffer_4679 (
        .din(new_Jinkela_wire_6396),
        .dout(new_Jinkela_wire_6397)
    );

    bfr new_Jinkela_buffer_4703 (
        .din(new_Jinkela_wire_6435),
        .dout(new_Jinkela_wire_6436)
    );

    bfr new_Jinkela_buffer_4680 (
        .din(new_Jinkela_wire_6397),
        .dout(new_Jinkela_wire_6398)
    );

    bfr new_Jinkela_buffer_4697 (
        .din(new_Jinkela_wire_6429),
        .dout(new_Jinkela_wire_6430)
    );

    bfr new_Jinkela_buffer_4681 (
        .din(new_Jinkela_wire_6398),
        .dout(new_Jinkela_wire_6399)
    );

    bfr new_Jinkela_buffer_4682 (
        .din(new_Jinkela_wire_6399),
        .dout(new_Jinkela_wire_6400)
    );

    bfr new_Jinkela_buffer_4698 (
        .din(new_Jinkela_wire_6430),
        .dout(new_Jinkela_wire_6431)
    );

    bfr new_Jinkela_buffer_4683 (
        .din(new_Jinkela_wire_6400),
        .dout(new_Jinkela_wire_6401)
    );

    bfr new_Jinkela_buffer_4704 (
        .din(new_Jinkela_wire_6436),
        .dout(new_Jinkela_wire_6437)
    );

    bfr new_Jinkela_buffer_4684 (
        .din(new_Jinkela_wire_6401),
        .dout(new_Jinkela_wire_6402)
    );

    bfr new_Jinkela_buffer_4699 (
        .din(new_Jinkela_wire_6431),
        .dout(new_Jinkela_wire_6432)
    );

    bfr new_Jinkela_buffer_4685 (
        .din(new_Jinkela_wire_6402),
        .dout(new_Jinkela_wire_6403)
    );

    bfr new_Jinkela_buffer_4738 (
        .din(new_Jinkela_wire_6472),
        .dout(new_Jinkela_wire_6473)
    );

    bfr new_Jinkela_buffer_4686 (
        .din(new_Jinkela_wire_6403),
        .dout(new_Jinkela_wire_6404)
    );

    bfr new_Jinkela_buffer_4700 (
        .din(new_Jinkela_wire_6432),
        .dout(new_Jinkela_wire_6433)
    );

    bfr new_Jinkela_buffer_4687 (
        .din(new_Jinkela_wire_6404),
        .dout(new_Jinkela_wire_6405)
    );

    bfr new_Jinkela_buffer_4705 (
        .din(new_Jinkela_wire_6437),
        .dout(new_Jinkela_wire_6438)
    );

    bfr new_Jinkela_buffer_4688 (
        .din(new_Jinkela_wire_6405),
        .dout(new_Jinkela_wire_6406)
    );

    bfr new_Jinkela_buffer_4701 (
        .din(new_Jinkela_wire_6433),
        .dout(new_Jinkela_wire_6434)
    );

    bfr new_Jinkela_buffer_4761 (
        .din(new_net_2381),
        .dout(new_Jinkela_wire_6496)
    );

    bfr new_Jinkela_buffer_4706 (
        .din(new_Jinkela_wire_6438),
        .dout(new_Jinkela_wire_6439)
    );

    spl2 new_Jinkela_splitter_665 (
        .a(_0931_),
        .b(new_Jinkela_wire_6498),
        .c(new_Jinkela_wire_6499)
    );

    spl2 new_Jinkela_splitter_666 (
        .a(new_net_0),
        .b(new_Jinkela_wire_6500),
        .c(new_Jinkela_wire_6504)
    );

    bfr new_Jinkela_buffer_4707 (
        .din(new_Jinkela_wire_6439),
        .dout(new_Jinkela_wire_6440)
    );

    bfr new_Jinkela_buffer_4739 (
        .din(new_Jinkela_wire_6473),
        .dout(new_Jinkela_wire_6474)
    );

    bfr new_Jinkela_buffer_4708 (
        .din(new_Jinkela_wire_6440),
        .dout(new_Jinkela_wire_6441)
    );

    bfr new_Jinkela_buffer_4762 (
        .din(new_Jinkela_wire_6496),
        .dout(new_Jinkela_wire_6497)
    );

    bfr new_Jinkela_buffer_4709 (
        .din(new_Jinkela_wire_6441),
        .dout(new_Jinkela_wire_6442)
    );

    bfr new_Jinkela_buffer_4740 (
        .din(new_Jinkela_wire_6474),
        .dout(new_Jinkela_wire_6475)
    );

    bfr new_Jinkela_buffer_4710 (
        .din(new_Jinkela_wire_6442),
        .dout(new_Jinkela_wire_6443)
    );

    spl2 new_Jinkela_splitter_670 (
        .a(_1143_),
        .b(new_Jinkela_wire_6549),
        .c(new_Jinkela_wire_6550)
    );

    bfr new_Jinkela_buffer_4711 (
        .din(new_Jinkela_wire_6443),
        .dout(new_Jinkela_wire_6444)
    );

    bfr new_Jinkela_buffer_4741 (
        .din(new_Jinkela_wire_6475),
        .dout(new_Jinkela_wire_6476)
    );

    bfr new_Jinkela_buffer_4712 (
        .din(new_Jinkela_wire_6444),
        .dout(new_Jinkela_wire_6445)
    );

    bfr new_Jinkela_buffer_4713 (
        .din(new_Jinkela_wire_6445),
        .dout(new_Jinkela_wire_6446)
    );

    bfr new_Jinkela_buffer_4742 (
        .din(new_Jinkela_wire_6476),
        .dout(new_Jinkela_wire_6477)
    );

    bfr new_Jinkela_buffer_4714 (
        .din(new_Jinkela_wire_6446),
        .dout(new_Jinkela_wire_6447)
    );

    bfr new_Jinkela_buffer_4800 (
        .din(new_net_2493),
        .dout(new_Jinkela_wire_6551)
    );

    bfr new_Jinkela_buffer_4715 (
        .din(new_Jinkela_wire_6447),
        .dout(new_Jinkela_wire_6448)
    );

    bfr new_Jinkela_buffer_4743 (
        .din(new_Jinkela_wire_6477),
        .dout(new_Jinkela_wire_6478)
    );

    bfr new_Jinkela_buffer_5567 (
        .din(_0198_),
        .dout(new_Jinkela_wire_7511)
    );

    bfr new_Jinkela_buffer_5474 (
        .din(new_Jinkela_wire_7406),
        .dout(new_Jinkela_wire_7407)
    );

    bfr new_Jinkela_buffer_5505 (
        .din(new_Jinkela_wire_7443),
        .dout(new_Jinkela_wire_7444)
    );

    bfr new_Jinkela_buffer_5475 (
        .din(new_Jinkela_wire_7407),
        .dout(new_Jinkela_wire_7408)
    );

    bfr new_Jinkela_buffer_5528 (
        .din(new_Jinkela_wire_7466),
        .dout(new_Jinkela_wire_7467)
    );

    bfr new_Jinkela_buffer_5476 (
        .din(new_Jinkela_wire_7408),
        .dout(new_Jinkela_wire_7409)
    );

    bfr new_Jinkela_buffer_5506 (
        .din(new_Jinkela_wire_7444),
        .dout(new_Jinkela_wire_7445)
    );

    bfr new_Jinkela_buffer_5477 (
        .din(new_Jinkela_wire_7409),
        .dout(new_Jinkela_wire_7410)
    );

    spl2 new_Jinkela_splitter_748 (
        .a(_0932_),
        .b(new_Jinkela_wire_7501),
        .c(new_Jinkela_wire_7502)
    );

    bfr new_Jinkela_buffer_5478 (
        .din(new_Jinkela_wire_7410),
        .dout(new_Jinkela_wire_7411)
    );

    bfr new_Jinkela_buffer_5507 (
        .din(new_Jinkela_wire_7445),
        .dout(new_Jinkela_wire_7446)
    );

    bfr new_Jinkela_buffer_5479 (
        .din(new_Jinkela_wire_7411),
        .dout(new_Jinkela_wire_7412)
    );

    bfr new_Jinkela_buffer_5529 (
        .din(new_Jinkela_wire_7467),
        .dout(new_Jinkela_wire_7468)
    );

    bfr new_Jinkela_buffer_5480 (
        .din(new_Jinkela_wire_7412),
        .dout(new_Jinkela_wire_7413)
    );

    bfr new_Jinkela_buffer_5508 (
        .din(new_Jinkela_wire_7446),
        .dout(new_Jinkela_wire_7447)
    );

    bfr new_Jinkela_buffer_5481 (
        .din(new_Jinkela_wire_7413),
        .dout(new_Jinkela_wire_7414)
    );

    bfr new_Jinkela_buffer_5531 (
        .din(new_Jinkela_wire_7472),
        .dout(new_Jinkela_wire_7473)
    );

    bfr new_Jinkela_buffer_5482 (
        .din(new_Jinkela_wire_7414),
        .dout(new_Jinkela_wire_7415)
    );

    bfr new_Jinkela_buffer_5509 (
        .din(new_Jinkela_wire_7447),
        .dout(new_Jinkela_wire_7448)
    );

    bfr new_Jinkela_buffer_5483 (
        .din(new_Jinkela_wire_7415),
        .dout(new_Jinkela_wire_7416)
    );

    bfr new_Jinkela_buffer_5559 (
        .din(new_Jinkela_wire_7502),
        .dout(new_Jinkela_wire_7503)
    );

    bfr new_Jinkela_buffer_5484 (
        .din(new_Jinkela_wire_7416),
        .dout(new_Jinkela_wire_7417)
    );

    bfr new_Jinkela_buffer_5510 (
        .din(new_Jinkela_wire_7448),
        .dout(new_Jinkela_wire_7449)
    );

    bfr new_Jinkela_buffer_5485 (
        .din(new_Jinkela_wire_7417),
        .dout(new_Jinkela_wire_7418)
    );

    bfr new_Jinkela_buffer_5532 (
        .din(new_Jinkela_wire_7473),
        .dout(new_Jinkela_wire_7474)
    );

    bfr new_Jinkela_buffer_5486 (
        .din(new_Jinkela_wire_7418),
        .dout(new_Jinkela_wire_7419)
    );

    bfr new_Jinkela_buffer_5511 (
        .din(new_Jinkela_wire_7449),
        .dout(new_Jinkela_wire_7450)
    );

    bfr new_Jinkela_buffer_5487 (
        .din(new_Jinkela_wire_7419),
        .dout(new_Jinkela_wire_7420)
    );

    spl2 new_Jinkela_splitter_750 (
        .a(_0071_),
        .b(new_Jinkela_wire_7517),
        .c(new_Jinkela_wire_7518)
    );

    bfr new_Jinkela_buffer_5488 (
        .din(new_Jinkela_wire_7420),
        .dout(new_Jinkela_wire_7421)
    );

    bfr new_Jinkela_buffer_5512 (
        .din(new_Jinkela_wire_7450),
        .dout(new_Jinkela_wire_7451)
    );

    bfr new_Jinkela_buffer_5489 (
        .din(new_Jinkela_wire_7421),
        .dout(new_Jinkela_wire_7422)
    );

    bfr new_Jinkela_buffer_5533 (
        .din(new_Jinkela_wire_7474),
        .dout(new_Jinkela_wire_7475)
    );

    bfr new_Jinkela_buffer_5490 (
        .din(new_Jinkela_wire_7422),
        .dout(new_Jinkela_wire_7423)
    );

    bfr new_Jinkela_buffer_5513 (
        .din(new_Jinkela_wire_7451),
        .dout(new_Jinkela_wire_7452)
    );

    bfr new_Jinkela_buffer_5491 (
        .din(new_Jinkela_wire_7423),
        .dout(new_Jinkela_wire_7424)
    );

    bfr new_Jinkela_buffer_5492 (
        .din(new_Jinkela_wire_7424),
        .dout(new_Jinkela_wire_7425)
    );

    bfr new_Jinkela_buffer_5514 (
        .din(new_Jinkela_wire_7452),
        .dout(new_Jinkela_wire_7453)
    );

    bfr new_Jinkela_buffer_5493 (
        .din(new_Jinkela_wire_7425),
        .dout(new_Jinkela_wire_7426)
    );

    bfr new_Jinkela_buffer_5534 (
        .din(new_Jinkela_wire_7475),
        .dout(new_Jinkela_wire_7476)
    );

    bfr new_Jinkela_buffer_5494 (
        .din(new_Jinkela_wire_7426),
        .dout(new_Jinkela_wire_7427)
    );

    bfr new_Jinkela_buffer_5515 (
        .din(new_Jinkela_wire_7453),
        .dout(new_Jinkela_wire_7454)
    );

    bfr new_Jinkela_buffer_4430 (
        .din(new_Jinkela_wire_6070),
        .dout(new_Jinkela_wire_6071)
    );

    bfr new_Jinkela_buffer_4419 (
        .din(new_Jinkela_wire_6055),
        .dout(new_Jinkela_wire_6056)
    );

    spl2 new_Jinkela_splitter_632 (
        .a(_0761_),
        .b(new_Jinkela_wire_6096),
        .c(new_Jinkela_wire_6097)
    );

    bfr new_Jinkela_buffer_4434 (
        .din(new_Jinkela_wire_6076),
        .dout(new_Jinkela_wire_6077)
    );

    bfr new_Jinkela_buffer_4420 (
        .din(new_Jinkela_wire_6056),
        .dout(new_Jinkela_wire_6057)
    );

    bfr new_Jinkela_buffer_4450 (
        .din(new_Jinkela_wire_6092),
        .dout(new_Jinkela_wire_6093)
    );

    bfr new_Jinkela_buffer_4421 (
        .din(new_Jinkela_wire_6057),
        .dout(new_Jinkela_wire_6058)
    );

    bfr new_Jinkela_buffer_4435 (
        .din(new_Jinkela_wire_6077),
        .dout(new_Jinkela_wire_6078)
    );

    bfr new_Jinkela_buffer_4422 (
        .din(new_Jinkela_wire_6058),
        .dout(new_Jinkela_wire_6059)
    );

    bfr new_Jinkela_buffer_4423 (
        .din(new_Jinkela_wire_6059),
        .dout(new_Jinkela_wire_6060)
    );

    bfr new_Jinkela_buffer_4436 (
        .din(new_Jinkela_wire_6078),
        .dout(new_Jinkela_wire_6079)
    );

    bfr new_Jinkela_buffer_4424 (
        .din(new_Jinkela_wire_6060),
        .dout(new_Jinkela_wire_6061)
    );

    bfr new_Jinkela_buffer_4425 (
        .din(new_Jinkela_wire_6061),
        .dout(new_Jinkela_wire_6062)
    );

    bfr new_Jinkela_buffer_4437 (
        .din(new_Jinkela_wire_6079),
        .dout(new_Jinkela_wire_6080)
    );

    spl2 new_Jinkela_splitter_628 (
        .a(new_Jinkela_wire_6062),
        .b(new_Jinkela_wire_6063),
        .c(new_Jinkela_wire_6064)
    );

    bfr new_Jinkela_buffer_4451 (
        .din(new_Jinkela_wire_6097),
        .dout(new_Jinkela_wire_6098)
    );

    bfr new_Jinkela_buffer_4438 (
        .din(new_Jinkela_wire_6080),
        .dout(new_Jinkela_wire_6081)
    );

    spl4L new_Jinkela_splitter_633 (
        .a(_0955_),
        .d(new_Jinkela_wire_6100),
        .e(new_Jinkela_wire_6101),
        .b(new_Jinkela_wire_6102),
        .c(new_Jinkela_wire_6103)
    );

    bfr new_Jinkela_buffer_4466 (
        .din(_1048_),
        .dout(new_Jinkela_wire_6117)
    );

    bfr new_Jinkela_buffer_4439 (
        .din(new_Jinkela_wire_6081),
        .dout(new_Jinkela_wire_6082)
    );

    spl2 new_Jinkela_splitter_634 (
        .a(_0180_),
        .b(new_Jinkela_wire_6122),
        .c(new_Jinkela_wire_6123)
    );

    bfr new_Jinkela_buffer_4452 (
        .din(new_Jinkela_wire_6098),
        .dout(new_Jinkela_wire_6099)
    );

    bfr new_Jinkela_buffer_4440 (
        .din(new_Jinkela_wire_6082),
        .dout(new_Jinkela_wire_6083)
    );

    bfr new_Jinkela_buffer_4454 (
        .din(new_Jinkela_wire_6104),
        .dout(new_Jinkela_wire_6105)
    );

    bfr new_Jinkela_buffer_4441 (
        .din(new_Jinkela_wire_6083),
        .dout(new_Jinkela_wire_6084)
    );

    bfr new_Jinkela_buffer_4453 (
        .din(new_Jinkela_wire_6103),
        .dout(new_Jinkela_wire_6104)
    );

    bfr new_Jinkela_buffer_4442 (
        .din(new_Jinkela_wire_6084),
        .dout(new_Jinkela_wire_6085)
    );

    bfr new_Jinkela_buffer_4471 (
        .din(_0591_),
        .dout(new_Jinkela_wire_6124)
    );

    bfr new_Jinkela_buffer_4467 (
        .din(new_Jinkela_wire_6117),
        .dout(new_Jinkela_wire_6118)
    );

    bfr new_Jinkela_buffer_4443 (
        .din(new_Jinkela_wire_6085),
        .dout(new_Jinkela_wire_6086)
    );

    bfr new_Jinkela_buffer_4444 (
        .din(new_Jinkela_wire_6086),
        .dout(new_Jinkela_wire_6087)
    );

    spl3L new_Jinkela_splitter_635 (
        .a(_0093_),
        .d(new_Jinkela_wire_6125),
        .b(new_Jinkela_wire_6128),
        .c(new_Jinkela_wire_6133)
    );

    bfr new_Jinkela_buffer_4455 (
        .din(new_Jinkela_wire_6105),
        .dout(new_Jinkela_wire_6106)
    );

    bfr new_Jinkela_buffer_4445 (
        .din(new_Jinkela_wire_6087),
        .dout(new_Jinkela_wire_6088)
    );

    bfr new_Jinkela_buffer_4472 (
        .din(_0614_),
        .dout(new_Jinkela_wire_6138)
    );

    bfr new_Jinkela_buffer_4446 (
        .din(new_Jinkela_wire_6088),
        .dout(new_Jinkela_wire_6089)
    );

    bfr new_Jinkela_buffer_4468 (
        .din(new_Jinkela_wire_6118),
        .dout(new_Jinkela_wire_6119)
    );

    bfr new_Jinkela_buffer_4456 (
        .din(new_Jinkela_wire_6106),
        .dout(new_Jinkela_wire_6107)
    );

    bfr new_Jinkela_buffer_4447 (
        .din(new_Jinkela_wire_6089),
        .dout(new_Jinkela_wire_6090)
    );

    bfr new_Jinkela_buffer_4448 (
        .din(new_Jinkela_wire_6090),
        .dout(new_Jinkela_wire_6091)
    );

    bfr new_Jinkela_buffer_4457 (
        .din(new_Jinkela_wire_6107),
        .dout(new_Jinkela_wire_6108)
    );

    bfr new_Jinkela_buffer_4469 (
        .din(new_Jinkela_wire_6119),
        .dout(new_Jinkela_wire_6120)
    );

    bfr new_Jinkela_buffer_4458 (
        .din(new_Jinkela_wire_6108),
        .dout(new_Jinkela_wire_6109)
    );

    inv _1274_ (
        .din(new_Jinkela_wire_1147),
        .dout(new_net_25)
    );

    and_ii _1991_ (
        .a(new_Jinkela_wire_2536),
        .b(new_Jinkela_wire_4978),
        .c(_0032_)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(new_Jinkela_wire_477),
        .b(new_Jinkela_wire_478),
        .c(new_Jinkela_wire_479)
    );

    inv _1275_ (
        .din(new_Jinkela_wire_970),
        .dout(new_net_26)
    );

    and_bb _1992_ (
        .a(new_Jinkela_wire_2537),
        .b(new_Jinkela_wire_4976),
        .c(_0033_)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    or_ii _1276_ (
        .a(new_Jinkela_wire_1549),
        .b(new_Jinkela_wire_1564),
        .c(_0586_)
    );

    or_bb _1993_ (
        .a(_0033_),
        .b(_0032_),
        .c(_0034_)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    and_bi _1277_ (
        .a(new_Jinkela_wire_1551),
        .b(new_Jinkela_wire_1555),
        .c(_0587_)
    );

    or_bb _1994_ (
        .a(new_Jinkela_wire_96),
        .b(new_Jinkela_wire_63),
        .c(_0035_)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(new_Jinkela_wire_534),
        .b(new_Jinkela_wire_535),
        .c(new_Jinkela_wire_536)
    );

    and_bi _1278_ (
        .a(_0586_),
        .b(_0587_),
        .c(_0588_)
    );

    and_bi _1995_ (
        .a(new_Jinkela_wire_102),
        .b(new_Jinkela_wire_412),
        .c(_0036_)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    or_bb _1279_ (
        .a(new_Jinkela_wire_5705),
        .b(new_Jinkela_wire_6510),
        .c(new_net_2507)
    );

    and_bi _1996_ (
        .a(_0035_),
        .b(_0036_),
        .c(_0037_)
    );

    or_ii _1280_ (
        .a(new_Jinkela_wire_704),
        .b(new_Jinkela_wire_1565),
        .c(_0589_)
    );

    and_bi _1997_ (
        .a(new_Jinkela_wire_1230),
        .b(_0037_),
        .c(_0038_)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    and_bi _1281_ (
        .a(new_Jinkela_wire_1384),
        .b(new_Jinkela_wire_1556),
        .c(_0590_)
    );

    or_ii _1998_ (
        .a(new_Jinkela_wire_97),
        .b(new_Jinkela_wire_1206),
        .c(_0039_)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(G92),
        .b(new_Jinkela_wire_552),
        .c(new_Jinkela_wire_554)
    );

    and_bi _1282_ (
        .a(_0589_),
        .b(_0590_),
        .c(_0591_)
    );

    and_bi _1999_ (
        .a(new_Jinkela_wire_1534),
        .b(new_Jinkela_wire_98),
        .c(_0040_)
    );

    spl3L new_Jinkela_splitter_99 (
        .a(new_Jinkela_wire_482),
        .d(new_Jinkela_wire_483),
        .b(new_Jinkela_wire_484),
        .c(new_Jinkela_wire_485)
    );

    or_bb _1283_ (
        .a(new_Jinkela_wire_6124),
        .b(new_Jinkela_wire_6509),
        .c(new_net_27)
    );

    and_bi _2000_ (
        .a(_0039_),
        .b(_0040_),
        .c(_0041_)
    );

    spl3L new_Jinkela_splitter_120 (
        .a(G66),
        .d(new_Jinkela_wire_573),
        .b(new_Jinkela_wire_574),
        .c(new_Jinkela_wire_575)
    );

    or_bi _1284_ (
        .a(new_Jinkela_wire_6506),
        .b(new_Jinkela_wire_957),
        .c(new_net_2495)
    );

    and_bi _2001_ (
        .a(new_Jinkela_wire_7186),
        .b(_0041_),
        .c(_0042_)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    spl2 new_Jinkela_splitter_100 (
        .a(new_Jinkela_wire_485),
        .b(new_Jinkela_wire_486),
        .c(new_Jinkela_wire_487)
    );

    or_bi _1285_ (
        .a(new_Jinkela_wire_1401),
        .b(new_Jinkela_wire_1030),
        .c(_0592_)
    );

    and_ii _2002_ (
        .a(_0042_),
        .b(_0038_),
        .c(_0043_)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    and_bi _1286_ (
        .a(new_Jinkela_wire_1488),
        .b(new_Jinkela_wire_6683),
        .c(_0593_)
    );

    or_bi _2003_ (
        .a(new_Jinkela_wire_5217),
        .b(new_Jinkela_wire_4601),
        .c(_0044_)
    );

    and_bb _1287_ (
        .a(new_Jinkela_wire_1367),
        .b(new_Jinkela_wire_874),
        .c(_0594_)
    );

    and_bi _2004_ (
        .a(new_Jinkela_wire_5218),
        .b(new_Jinkela_wire_4602),
        .c(_0045_)
    );

    and_bi _1288_ (
        .a(new_Jinkela_wire_776),
        .b(new_Jinkela_wire_890),
        .c(_0595_)
    );

    and_bi _2005_ (
        .a(_0044_),
        .b(_0045_),
        .c(_0046_)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_488),
        .dout(new_Jinkela_wire_489)
    );

    and_ii _1289_ (
        .a(_0595_),
        .b(_0594_),
        .c(_0596_)
    );

    or_bb _2006_ (
        .a(new_Jinkela_wire_289),
        .b(new_Jinkela_wire_58),
        .c(_0047_)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    or_bb _1290_ (
        .a(new_Jinkela_wire_6018),
        .b(new_Jinkela_wire_1500),
        .c(_0597_)
    );

    and_bi _2007_ (
        .a(new_Jinkela_wire_292),
        .b(new_Jinkela_wire_417),
        .c(_0048_)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_489),
        .dout(new_Jinkela_wire_490)
    );

    and_bb _1291_ (
        .a(new_Jinkela_wire_6019),
        .b(new_Jinkela_wire_1501),
        .c(_0598_)
    );

    and_bi _2008_ (
        .a(_0047_),
        .b(_0048_),
        .c(_0049_)
    );

    and_bi _1292_ (
        .a(_0597_),
        .b(_0598_),
        .c(_0599_)
    );

    and_bi _2009_ (
        .a(new_Jinkela_wire_734),
        .b(_0049_),
        .c(_0050_)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    spl2 new_Jinkela_splitter_101 (
        .a(new_Jinkela_wire_490),
        .b(new_Jinkela_wire_491),
        .c(new_Jinkela_wire_492)
    );

    or_bb _1293_ (
        .a(new_Jinkela_wire_6225),
        .b(new_Jinkela_wire_1062),
        .c(_0600_)
    );

    or_ii _2010_ (
        .a(new_Jinkela_wire_285),
        .b(new_Jinkela_wire_1201),
        .c(_0051_)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(new_Jinkela_wire_492),
        .b(new_Jinkela_wire_493),
        .c(new_Jinkela_wire_494)
    );

    and_ii _1297_ (
        .a(_0603_),
        .b(_0602_),
        .c(_0604_)
    );

    and_bi _2011_ (
        .a(new_Jinkela_wire_1537),
        .b(new_Jinkela_wire_294),
        .c(_0052_)
    );

    and_bi _1298_ (
        .a(new_Jinkela_wire_1038),
        .b(new_Jinkela_wire_4977),
        .c(_0605_)
    );

    and_bi _2012_ (
        .a(_0051_),
        .b(_0052_),
        .c(_0053_)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(new_Jinkela_wire_494),
        .b(new_Jinkela_wire_495),
        .c(new_Jinkela_wire_496)
    );

    or_bb _1299_ (
        .a(_0605_),
        .b(new_Jinkela_wire_4822),
        .c(_0606_)
    );

    and_bi _2013_ (
        .a(new_Jinkela_wire_6142),
        .b(_0053_),
        .c(_0054_)
    );

    and_bi _1300_ (
        .a(_0600_),
        .b(new_Jinkela_wire_6255),
        .c(_0607_)
    );

    or_bb _2014_ (
        .a(_0054_),
        .b(_0050_),
        .c(_0055_)
    );

    spl3L new_Jinkela_splitter_104 (
        .a(new_Jinkela_wire_496),
        .d(new_Jinkela_wire_497),
        .b(new_Jinkela_wire_498),
        .c(new_Jinkela_wire_499)
    );

    and_ii _1301_ (
        .a(_0607_),
        .b(new_Jinkela_wire_2460),
        .c(new_net_4)
    );

    or_bb _2015_ (
        .a(new_Jinkela_wire_428),
        .b(new_Jinkela_wire_45),
        .c(_0056_)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_568),
        .dout(new_Jinkela_wire_569)
    );

    and_bi _1302_ (
        .a(new_Jinkela_wire_1601),
        .b(new_Jinkela_wire_6698),
        .c(_0608_)
    );

    and_bi _2016_ (
        .a(new_Jinkela_wire_434),
        .b(new_Jinkela_wire_402),
        .c(_0057_)
    );

    spl2 new_Jinkela_splitter_115 (
        .a(new_Jinkela_wire_545),
        .b(new_Jinkela_wire_546),
        .c(new_Jinkela_wire_547)
    );

    inv _1303_ (
        .din(new_Jinkela_wire_6016),
        .dout(_0609_)
    );

    and_bi _2017_ (
        .a(_0056_),
        .b(_0057_),
        .c(_0058_)
    );

    spl4L new_Jinkela_splitter_117 (
        .a(new_Jinkela_wire_554),
        .d(new_Jinkela_wire_555),
        .e(new_Jinkela_wire_556),
        .b(new_Jinkela_wire_558),
        .c(new_Jinkela_wire_563)
    );

    or_ii _1304_ (
        .a(new_Jinkela_wire_296),
        .b(new_Jinkela_wire_893),
        .c(_0610_)
    );

    and_bi _2018_ (
        .a(new_Jinkela_wire_1132),
        .b(_0058_),
        .c(_0059_)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    and_bi _1305_ (
        .a(new_Jinkela_wire_1238),
        .b(new_Jinkela_wire_886),
        .c(_0611_)
    );

    or_ii _2019_ (
        .a(new_Jinkela_wire_425),
        .b(new_Jinkela_wire_1199),
        .c(_0060_)
    );

    bfr new_Jinkela_buffer_222 (
        .din(G56),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_267 (
        .din(G9),
        .dout(new_Jinkela_wire_622)
    );

    and_bi _1306_ (
        .a(_0610_),
        .b(new_Jinkela_wire_3411),
        .c(_0612_)
    );

    and_bi _2020_ (
        .a(new_Jinkela_wire_1532),
        .b(new_Jinkela_wire_432),
        .c(_0061_)
    );

    and_bi _1307_ (
        .a(new_Jinkela_wire_737),
        .b(new_Jinkela_wire_4918),
        .c(_0613_)
    );

    and_bi _2021_ (
        .a(_0060_),
        .b(_0061_),
        .c(_0062_)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    spl4L new_Jinkela_splitter_118 (
        .a(new_Jinkela_wire_558),
        .d(new_Jinkela_wire_559),
        .e(new_Jinkela_wire_560),
        .b(new_Jinkela_wire_561),
        .c(new_Jinkela_wire_562)
    );

    inv _1308_ (
        .din(new_Jinkela_wire_729),
        .dout(_0614_)
    );

    and_bi _2022_ (
        .a(new_Jinkela_wire_3585),
        .b(_0062_),
        .c(_0063_)
    );

    or_ii _1309_ (
        .a(new_Jinkela_wire_4917),
        .b(new_Jinkela_wire_6145),
        .c(_0615_)
    );

    or_bb _2023_ (
        .a(_0063_),
        .b(_0059_),
        .c(_0064_)
    );

    spl4L new_Jinkela_splitter_119 (
        .a(new_Jinkela_wire_563),
        .d(new_Jinkela_wire_564),
        .e(new_Jinkela_wire_565),
        .b(new_Jinkela_wire_566),
        .c(new_Jinkela_wire_567)
    );

    and_bi _1310_ (
        .a(new_Jinkela_wire_4530),
        .b(new_Jinkela_wire_6356),
        .c(_0616_)
    );

    and_ii _2024_ (
        .a(new_Jinkela_wire_4756),
        .b(new_Jinkela_wire_6890),
        .c(_0065_)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    and_bi _1311_ (
        .a(new_Jinkela_wire_2901),
        .b(_0616_),
        .c(_0617_)
    );

    and_bb _2025_ (
        .a(new_Jinkela_wire_4757),
        .b(new_Jinkela_wire_6891),
        .c(_0066_)
    );

    bfr new_Jinkela_buffer_269 (
        .din(G112),
        .dout(new_Jinkela_wire_624)
    );

    and_bi _1312_ (
        .a(new_Jinkela_wire_6023),
        .b(new_Jinkela_wire_6355),
        .c(_0618_)
    );

    and_ii _2026_ (
        .a(_0066_),
        .b(_0065_),
        .c(_0067_)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    and_bb _1313_ (
        .a(new_Jinkela_wire_5902),
        .b(new_Jinkela_wire_4534),
        .c(_0619_)
    );

    or_bb _2027_ (
        .a(new_Jinkela_wire_1969),
        .b(new_Jinkela_wire_5706),
        .c(_0068_)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    or_bb _1314_ (
        .a(new_Jinkela_wire_2407),
        .b(new_Jinkela_wire_5901),
        .c(_0620_)
    );

    and_bb _2028_ (
        .a(new_Jinkela_wire_1970),
        .b(new_Jinkela_wire_5707),
        .c(_0069_)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_622),
        .dout(new_Jinkela_wire_623)
    );

    or_bb _1315_ (
        .a(new_Jinkela_wire_4343),
        .b(new_Jinkela_wire_1069),
        .c(_0621_)
    );

    and_bi _2029_ (
        .a(_0068_),
        .b(_0069_),
        .c(_0070_)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    or_bb _1316_ (
        .a(new_Jinkela_wire_293),
        .b(new_Jinkela_wire_318),
        .c(_0622_)
    );

    and_ii _2030_ (
        .a(new_Jinkela_wire_4706),
        .b(new_Jinkela_wire_7145),
        .c(_0071_)
    );

    bfr new_Jinkela_buffer_271 (
        .din(G171),
        .dout(new_Jinkela_wire_626)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    and_bi _1317_ (
        .a(new_Jinkela_wire_288),
        .b(new_Jinkela_wire_217),
        .c(_0623_)
    );

    and_bb _2031_ (
        .a(new_Jinkela_wire_4708),
        .b(new_Jinkela_wire_7146),
        .c(_0072_)
    );

    and_bi _1318_ (
        .a(_0622_),
        .b(_0623_),
        .c(_0624_)
    );

    and_ii _2032_ (
        .a(new_Jinkela_wire_5489),
        .b(new_Jinkela_wire_7517),
        .c(_0073_)
    );

    bfr new_Jinkela_buffer_4716 (
        .din(new_Jinkela_wire_6448),
        .dout(new_Jinkela_wire_6449)
    );

    spl4L new_Jinkela_splitter_668 (
        .a(new_Jinkela_wire_6504),
        .d(new_Jinkela_wire_6505),
        .e(new_Jinkela_wire_6506),
        .b(new_Jinkela_wire_6507),
        .c(new_Jinkela_wire_6508)
    );

    bfr new_Jinkela_buffer_4803 (
        .din(_0220_),
        .dout(new_Jinkela_wire_6556)
    );

    bfr new_Jinkela_buffer_4717 (
        .din(new_Jinkela_wire_6449),
        .dout(new_Jinkela_wire_6450)
    );

    bfr new_Jinkela_buffer_4744 (
        .din(new_Jinkela_wire_6478),
        .dout(new_Jinkela_wire_6479)
    );

    bfr new_Jinkela_buffer_4718 (
        .din(new_Jinkela_wire_6450),
        .dout(new_Jinkela_wire_6451)
    );

    spl3L new_Jinkela_splitter_667 (
        .a(new_Jinkela_wire_6500),
        .d(new_Jinkela_wire_6501),
        .b(new_Jinkela_wire_6502),
        .c(new_Jinkela_wire_6503)
    );

    bfr new_Jinkela_buffer_4719 (
        .din(new_Jinkela_wire_6451),
        .dout(new_Jinkela_wire_6452)
    );

    bfr new_Jinkela_buffer_4745 (
        .din(new_Jinkela_wire_6479),
        .dout(new_Jinkela_wire_6480)
    );

    bfr new_Jinkela_buffer_4720 (
        .din(new_Jinkela_wire_6452),
        .dout(new_Jinkela_wire_6453)
    );

    spl3L new_Jinkela_splitter_669 (
        .a(new_Jinkela_wire_6508),
        .d(new_Jinkela_wire_6509),
        .b(new_Jinkela_wire_6510),
        .c(new_Jinkela_wire_6511)
    );

    bfr new_Jinkela_buffer_4721 (
        .din(new_Jinkela_wire_6453),
        .dout(new_Jinkela_wire_6454)
    );

    bfr new_Jinkela_buffer_4746 (
        .din(new_Jinkela_wire_6480),
        .dout(new_Jinkela_wire_6481)
    );

    bfr new_Jinkela_buffer_4722 (
        .din(new_Jinkela_wire_6454),
        .dout(new_Jinkela_wire_6455)
    );

    spl2 new_Jinkela_splitter_671 (
        .a(_0654_),
        .b(new_Jinkela_wire_6554),
        .c(new_Jinkela_wire_6555)
    );

    bfr new_Jinkela_buffer_4723 (
        .din(new_Jinkela_wire_6455),
        .dout(new_Jinkela_wire_6456)
    );

    bfr new_Jinkela_buffer_4747 (
        .din(new_Jinkela_wire_6481),
        .dout(new_Jinkela_wire_6482)
    );

    bfr new_Jinkela_buffer_4724 (
        .din(new_Jinkela_wire_6456),
        .dout(new_Jinkela_wire_6457)
    );

    spl3L new_Jinkela_splitter_672 (
        .a(_0747_),
        .d(new_Jinkela_wire_6558),
        .b(new_Jinkela_wire_6559),
        .c(new_Jinkela_wire_6560)
    );

    bfr new_Jinkela_buffer_4725 (
        .din(new_Jinkela_wire_6457),
        .dout(new_Jinkela_wire_6458)
    );

    bfr new_Jinkela_buffer_4748 (
        .din(new_Jinkela_wire_6482),
        .dout(new_Jinkela_wire_6483)
    );

    bfr new_Jinkela_buffer_4726 (
        .din(new_Jinkela_wire_6458),
        .dout(new_Jinkela_wire_6459)
    );

    bfr new_Jinkela_buffer_4801 (
        .din(new_Jinkela_wire_6551),
        .dout(new_Jinkela_wire_6552)
    );

    bfr new_Jinkela_buffer_4806 (
        .din(_1027_),
        .dout(new_Jinkela_wire_6564)
    );

    bfr new_Jinkela_buffer_4727 (
        .din(new_Jinkela_wire_6459),
        .dout(new_Jinkela_wire_6460)
    );

    bfr new_Jinkela_buffer_4749 (
        .din(new_Jinkela_wire_6483),
        .dout(new_Jinkela_wire_6484)
    );

    bfr new_Jinkela_buffer_4728 (
        .din(new_Jinkela_wire_6460),
        .dout(new_Jinkela_wire_6461)
    );

    bfr new_Jinkela_buffer_4763 (
        .din(new_Jinkela_wire_6511),
        .dout(new_Jinkela_wire_6512)
    );

    bfr new_Jinkela_buffer_4729 (
        .din(new_Jinkela_wire_6461),
        .dout(new_Jinkela_wire_6462)
    );

    bfr new_Jinkela_buffer_4750 (
        .din(new_Jinkela_wire_6484),
        .dout(new_Jinkela_wire_6485)
    );

    bfr new_Jinkela_buffer_4730 (
        .din(new_Jinkela_wire_6462),
        .dout(new_Jinkela_wire_6463)
    );

    bfr new_Jinkela_buffer_4802 (
        .din(new_Jinkela_wire_6552),
        .dout(new_Jinkela_wire_6553)
    );

    bfr new_Jinkela_buffer_4731 (
        .din(new_Jinkela_wire_6463),
        .dout(new_Jinkela_wire_6464)
    );

    bfr new_Jinkela_buffer_4751 (
        .din(new_Jinkela_wire_6485),
        .dout(new_Jinkela_wire_6486)
    );

    bfr new_Jinkela_buffer_4732 (
        .din(new_Jinkela_wire_6464),
        .dout(new_Jinkela_wire_6465)
    );

    bfr new_Jinkela_buffer_4764 (
        .din(new_Jinkela_wire_6512),
        .dout(new_Jinkela_wire_6513)
    );

    bfr new_Jinkela_buffer_4733 (
        .din(new_Jinkela_wire_6465),
        .dout(new_Jinkela_wire_6466)
    );

    bfr new_Jinkela_buffer_4752 (
        .din(new_Jinkela_wire_6486),
        .dout(new_Jinkela_wire_6487)
    );

    bfr new_Jinkela_buffer_4734 (
        .din(new_Jinkela_wire_6466),
        .dout(new_Jinkela_wire_6467)
    );

    bfr new_Jinkela_buffer_4735 (
        .din(new_Jinkela_wire_6467),
        .dout(new_Jinkela_wire_6468)
    );

    bfr new_Jinkela_buffer_4753 (
        .din(new_Jinkela_wire_6487),
        .dout(new_Jinkela_wire_6488)
    );

    bfr new_Jinkela_buffer_4736 (
        .din(new_Jinkela_wire_6468),
        .dout(new_Jinkela_wire_6469)
    );

    bfr new_Jinkela_buffer_4765 (
        .din(new_Jinkela_wire_6513),
        .dout(new_Jinkela_wire_6514)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_1447),
        .dout(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_5495 (
        .din(new_Jinkela_wire_7427),
        .dout(new_Jinkela_wire_7428)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    spl2 new_Jinkela_splitter_751 (
        .a(_0074_),
        .b(new_Jinkela_wire_7520),
        .c(new_Jinkela_wire_7521)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(new_Jinkela_wire_1066),
        .b(new_Jinkela_wire_1067),
        .c(new_Jinkela_wire_1068)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_1494),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_5560 (
        .din(new_Jinkela_wire_7503),
        .dout(new_Jinkela_wire_7504)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_1448),
        .dout(new_Jinkela_wire_1449)
    );

    bfr new_Jinkela_buffer_5496 (
        .din(new_Jinkela_wire_7428),
        .dout(new_Jinkela_wire_7429)
    );

    spl2 new_Jinkela_splitter_194 (
        .a(new_Jinkela_wire_1068),
        .b(new_Jinkela_wire_1069),
        .c(new_Jinkela_wire_1070)
    );

    bfr new_Jinkela_buffer_5516 (
        .din(new_Jinkela_wire_7454),
        .dout(new_Jinkela_wire_7455)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_1130),
        .dout(new_Jinkela_wire_1131)
    );

    spl2 new_Jinkela_splitter_270 (
        .a(new_Jinkela_wire_1491),
        .b(new_Jinkela_wire_1492),
        .c(new_Jinkela_wire_1493)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_1449),
        .dout(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_5497 (
        .din(new_Jinkela_wire_7429),
        .dout(new_Jinkela_wire_7430)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_1070),
        .dout(new_Jinkela_wire_1071)
    );

    bfr new_Jinkela_buffer_5535 (
        .din(new_Jinkela_wire_7476),
        .dout(new_Jinkela_wire_7477)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(new_Jinkela_wire_1122),
        .b(new_Jinkela_wire_1123),
        .c(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_1495),
        .dout(new_Jinkela_wire_1496)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_1450),
        .dout(new_Jinkela_wire_1451)
    );

    bfr new_Jinkela_buffer_5498 (
        .din(new_Jinkela_wire_7430),
        .dout(new_Jinkela_wire_7431)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    bfr new_Jinkela_buffer_5517 (
        .din(new_Jinkela_wire_7455),
        .dout(new_Jinkela_wire_7456)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_1451),
        .dout(new_Jinkela_wire_1452)
    );

    bfr new_Jinkela_buffer_591 (
        .din(G26),
        .dout(new_Jinkela_wire_1190)
    );

    bfr new_Jinkela_buffer_5568 (
        .din(new_Jinkela_wire_7511),
        .dout(new_Jinkela_wire_7512)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_1139),
        .dout(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_5518 (
        .din(new_Jinkela_wire_7456),
        .dout(new_Jinkela_wire_7457)
    );

    spl3L new_Jinkela_splitter_195 (
        .a(new_Jinkela_wire_1072),
        .d(new_Jinkela_wire_1073),
        .b(new_Jinkela_wire_1074),
        .c(new_Jinkela_wire_1075)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_1502),
        .dout(new_Jinkela_wire_1503)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_1452),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_5536 (
        .din(new_Jinkela_wire_7477),
        .dout(new_Jinkela_wire_7478)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_1131),
        .dout(new_Jinkela_wire_1132)
    );

    bfr new_Jinkela_buffer_5519 (
        .din(new_Jinkela_wire_7457),
        .dout(new_Jinkela_wire_7458)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_1075),
        .dout(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_1496),
        .dout(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_1453),
        .dout(new_Jinkela_wire_1454)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    bfr new_Jinkela_buffer_5561 (
        .din(new_Jinkela_wire_7504),
        .dout(new_Jinkela_wire_7505)
    );

    bfr new_Jinkela_buffer_5520 (
        .din(new_Jinkela_wire_7458),
        .dout(new_Jinkela_wire_7459)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(new_Jinkela_wire_1076),
        .b(new_Jinkela_wire_1077),
        .c(new_Jinkela_wire_1078)
    );

    bfr new_Jinkela_buffer_763 (
        .din(G34),
        .dout(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_5537 (
        .din(new_Jinkela_wire_7478),
        .dout(new_Jinkela_wire_7479)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    bfr new_Jinkela_buffer_5521 (
        .din(new_Jinkela_wire_7459),
        .dout(new_Jinkela_wire_7460)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_1497),
        .dout(new_Jinkela_wire_1498)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_1138),
        .dout(new_Jinkela_wire_1139)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_1148),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_5522 (
        .din(new_Jinkela_wire_7460),
        .dout(new_Jinkela_wire_7461)
    );

    spl4L new_Jinkela_splitter_197 (
        .a(new_Jinkela_wire_1079),
        .d(new_Jinkela_wire_1080),
        .e(new_Jinkela_wire_1081),
        .b(new_Jinkela_wire_1082),
        .c(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_1503),
        .dout(new_Jinkela_wire_1504)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_5538 (
        .din(new_Jinkela_wire_7479),
        .dout(new_Jinkela_wire_7480)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(new_Jinkela_wire_1083),
        .b(new_Jinkela_wire_1084),
        .c(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_1498),
        .dout(new_Jinkela_wire_1499)
    );

    bfr new_Jinkela_buffer_5562 (
        .din(new_Jinkela_wire_7505),
        .dout(new_Jinkela_wire_7506)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_5539 (
        .din(new_Jinkela_wire_7480),
        .dout(new_Jinkela_wire_7481)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_1085),
        .dout(new_Jinkela_wire_1086)
    );

    spl3L new_Jinkela_splitter_212 (
        .a(G1),
        .d(new_Jinkela_wire_1146),
        .b(new_Jinkela_wire_1147),
        .c(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_5569 (
        .din(new_Jinkela_wire_7512),
        .dout(new_Jinkela_wire_7513)
    );

    bfr new_Jinkela_buffer_597 (
        .din(G17),
        .dout(new_Jinkela_wire_1220)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    bfr new_Jinkela_buffer_5540 (
        .din(new_Jinkela_wire_7481),
        .dout(new_Jinkela_wire_7482)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_1140),
        .dout(new_Jinkela_wire_1141)
    );

    spl2 new_Jinkela_splitter_277 (
        .a(G98),
        .b(new_Jinkela_wire_1527),
        .c(new_Jinkela_wire_1531)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_1086),
        .dout(new_Jinkela_wire_1087)
    );

    spl2 new_Jinkela_splitter_271 (
        .a(new_Jinkela_wire_1499),
        .b(new_Jinkela_wire_1500),
        .c(new_Jinkela_wire_1501)
    );

    bfr new_Jinkela_buffer_5563 (
        .din(new_Jinkela_wire_7506),
        .dout(new_Jinkela_wire_7507)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_5541 (
        .din(new_Jinkela_wire_7482),
        .dout(new_Jinkela_wire_7483)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    spl2 new_Jinkela_splitter_199 (
        .a(new_Jinkela_wire_1087),
        .b(new_Jinkela_wire_1088),
        .c(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_1523),
        .dout(new_Jinkela_wire_1524)
    );

    bfr new_Jinkela_buffer_5571 (
        .din(new_Jinkela_wire_7518),
        .dout(new_Jinkela_wire_7519)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_5542 (
        .din(new_Jinkela_wire_7483),
        .dout(new_Jinkela_wire_7484)
    );

    spl3L new_Jinkela_splitter_200 (
        .a(new_Jinkela_wire_1089),
        .d(new_Jinkela_wire_1090),
        .b(new_Jinkela_wire_1091),
        .c(new_Jinkela_wire_1092)
    );

    spl2 new_Jinkela_splitter_752 (
        .a(_1134_),
        .b(new_Jinkela_wire_7522),
        .c(new_Jinkela_wire_7523)
    );

    spl2 new_Jinkela_splitter_272 (
        .a(new_Jinkela_wire_1504),
        .b(new_Jinkela_wire_1505),
        .c(new_Jinkela_wire_1506)
    );

    bfr new_Jinkela_buffer_5564 (
        .din(new_Jinkela_wire_7507),
        .dout(new_Jinkela_wire_7508)
    );

    bfr new_Jinkela_buffer_594 (
        .din(G70),
        .dout(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_5543 (
        .din(new_Jinkela_wire_7484),
        .dout(new_Jinkela_wire_7485)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(G102),
        .b(new_Jinkela_wire_1195),
        .c(new_Jinkela_wire_1198)
    );

    spl3L new_Jinkela_splitter_211 (
        .a(new_Jinkela_wire_1141),
        .d(new_Jinkela_wire_1142),
        .b(new_Jinkela_wire_1143),
        .c(new_Jinkela_wire_1144)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    bfr new_Jinkela_buffer_5570 (
        .din(new_Jinkela_wire_7513),
        .dout(new_Jinkela_wire_7514)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    bfr new_Jinkela_buffer_5544 (
        .din(new_Jinkela_wire_7485),
        .dout(new_Jinkela_wire_7486)
    );

    spl3L new_Jinkela_splitter_201 (
        .a(new_Jinkela_wire_1093),
        .d(new_Jinkela_wire_1094),
        .b(new_Jinkela_wire_1095),
        .c(new_Jinkela_wire_1096)
    );

    bfr new_Jinkela_buffer_5565 (
        .din(new_Jinkela_wire_7508),
        .dout(new_Jinkela_wire_7509)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_5545 (
        .din(new_Jinkela_wire_7486),
        .dout(new_Jinkela_wire_7487)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_1190),
        .dout(new_Jinkela_wire_1191)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_1144),
        .dout(new_Jinkela_wire_1145)
    );

    spl3L new_Jinkela_splitter_202 (
        .a(new_Jinkela_wire_1096),
        .d(new_Jinkela_wire_1097),
        .b(new_Jinkela_wire_1098),
        .c(new_Jinkela_wire_1099)
    );

    bfr new_Jinkela_buffer_765 (
        .din(G33),
        .dout(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_5546 (
        .din(new_Jinkela_wire_7487),
        .dout(new_Jinkela_wire_7488)
    );

    bfr new_Jinkela_buffer_760 (
        .din(G71),
        .dout(new_Jinkela_wire_1522)
    );

    spl2 new_Jinkela_splitter_753 (
        .a(_0162_),
        .b(new_Jinkela_wire_7524),
        .c(new_Jinkela_wire_7525)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_1099),
        .dout(new_Jinkela_wire_1100)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_5566 (
        .din(new_Jinkela_wire_7509),
        .dout(new_Jinkela_wire_7510)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_1465),
        .dout(new_Jinkela_wire_1466)
    );

    bfr new_Jinkela_buffer_5547 (
        .din(new_Jinkela_wire_7488),
        .dout(new_Jinkela_wire_7489)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    spl2 new_Jinkela_splitter_749 (
        .a(new_Jinkela_wire_7514),
        .b(new_Jinkela_wire_7515),
        .c(new_Jinkela_wire_7516)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_1466),
        .dout(new_Jinkela_wire_1467)
    );

    bfr new_Jinkela_buffer_5548 (
        .din(new_Jinkela_wire_7489),
        .dout(new_Jinkela_wire_7490)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_1151),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_1522),
        .dout(new_Jinkela_wire_1523)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_1191),
        .dout(new_Jinkela_wire_1192)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_1511),
        .dout(new_Jinkela_wire_1512)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_1467),
        .dout(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_5549 (
        .din(new_Jinkela_wire_7490),
        .dout(new_Jinkela_wire_7491)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_1152),
        .dout(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_5572 (
        .din(new_net_24),
        .dout(new_Jinkela_wire_7526)
    );

    bfr new_Jinkela_buffer_3655 (
        .din(_0566_),
        .dout(new_Jinkela_wire_5116)
    );

    bfr new_Jinkela_buffer_4372 (
        .din(new_Jinkela_wire_5995),
        .dout(new_Jinkela_wire_5996)
    );

    bfr new_Jinkela_buffer_4449 (
        .din(_0399_),
        .dout(new_Jinkela_wire_6092)
    );

    bfr new_Jinkela_buffer_4401 (
        .din(new_Jinkela_wire_6032),
        .dout(new_Jinkela_wire_6033)
    );

    bfr new_Jinkela_buffer_4373 (
        .din(new_Jinkela_wire_5996),
        .dout(new_Jinkela_wire_5997)
    );

    bfr new_Jinkela_buffer_4427 (
        .din(new_Jinkela_wire_6067),
        .dout(new_Jinkela_wire_6068)
    );

    bfr new_Jinkela_buffer_4374 (
        .din(new_Jinkela_wire_5997),
        .dout(new_Jinkela_wire_5998)
    );

    bfr new_Jinkela_buffer_4402 (
        .din(new_Jinkela_wire_6033),
        .dout(new_Jinkela_wire_6034)
    );

    bfr new_Jinkela_buffer_4375 (
        .din(new_Jinkela_wire_5998),
        .dout(new_Jinkela_wire_5999)
    );

    bfr new_Jinkela_buffer_4413 (
        .din(new_Jinkela_wire_6049),
        .dout(new_Jinkela_wire_6050)
    );

    bfr new_Jinkela_buffer_4376 (
        .din(new_Jinkela_wire_5999),
        .dout(new_Jinkela_wire_6000)
    );

    bfr new_Jinkela_buffer_4403 (
        .din(new_Jinkela_wire_6034),
        .dout(new_Jinkela_wire_6035)
    );

    bfr new_Jinkela_buffer_4377 (
        .din(new_Jinkela_wire_6000),
        .dout(new_Jinkela_wire_6001)
    );

    bfr new_Jinkela_buffer_4378 (
        .din(new_Jinkela_wire_6001),
        .dout(new_Jinkela_wire_6002)
    );

    bfr new_Jinkela_buffer_4432 (
        .din(_0444_),
        .dout(new_Jinkela_wire_6075)
    );

    bfr new_Jinkela_buffer_4404 (
        .din(new_Jinkela_wire_6035),
        .dout(new_Jinkela_wire_6036)
    );

    bfr new_Jinkela_buffer_4379 (
        .din(new_Jinkela_wire_6002),
        .dout(new_Jinkela_wire_6003)
    );

    bfr new_Jinkela_buffer_4414 (
        .din(new_Jinkela_wire_6050),
        .dout(new_Jinkela_wire_6051)
    );

    bfr new_Jinkela_buffer_4380 (
        .din(new_Jinkela_wire_6003),
        .dout(new_Jinkela_wire_6004)
    );

    bfr new_Jinkela_buffer_4405 (
        .din(new_Jinkela_wire_6036),
        .dout(new_Jinkela_wire_6037)
    );

    bfr new_Jinkela_buffer_4381 (
        .din(new_Jinkela_wire_6004),
        .dout(new_Jinkela_wire_6005)
    );

    bfr new_Jinkela_buffer_4428 (
        .din(new_Jinkela_wire_6068),
        .dout(new_Jinkela_wire_6069)
    );

    bfr new_Jinkela_buffer_4382 (
        .din(new_Jinkela_wire_6005),
        .dout(new_Jinkela_wire_6006)
    );

    bfr new_Jinkela_buffer_4406 (
        .din(new_Jinkela_wire_6037),
        .dout(new_Jinkela_wire_6038)
    );

    bfr new_Jinkela_buffer_4383 (
        .din(new_Jinkela_wire_6006),
        .dout(new_Jinkela_wire_6007)
    );

    bfr new_Jinkela_buffer_4415 (
        .din(new_Jinkela_wire_6051),
        .dout(new_Jinkela_wire_6052)
    );

    bfr new_Jinkela_buffer_4384 (
        .din(new_Jinkela_wire_6007),
        .dout(new_Jinkela_wire_6008)
    );

    bfr new_Jinkela_buffer_4407 (
        .din(new_Jinkela_wire_6038),
        .dout(new_Jinkela_wire_6039)
    );

    bfr new_Jinkela_buffer_4385 (
        .din(new_Jinkela_wire_6008),
        .dout(new_Jinkela_wire_6009)
    );

    bfr new_Jinkela_buffer_4386 (
        .din(new_Jinkela_wire_6009),
        .dout(new_Jinkela_wire_6010)
    );

    bfr new_Jinkela_buffer_4433 (
        .din(new_Jinkela_wire_6075),
        .dout(new_Jinkela_wire_6076)
    );

    bfr new_Jinkela_buffer_4408 (
        .din(new_Jinkela_wire_6039),
        .dout(new_Jinkela_wire_6040)
    );

    bfr new_Jinkela_buffer_4387 (
        .din(new_Jinkela_wire_6010),
        .dout(new_Jinkela_wire_6011)
    );

    bfr new_Jinkela_buffer_4416 (
        .din(new_Jinkela_wire_6052),
        .dout(new_Jinkela_wire_6053)
    );

    bfr new_Jinkela_buffer_4388 (
        .din(new_Jinkela_wire_6011),
        .dout(new_Jinkela_wire_6012)
    );

    bfr new_Jinkela_buffer_4409 (
        .din(new_Jinkela_wire_6040),
        .dout(new_Jinkela_wire_6041)
    );

    bfr new_Jinkela_buffer_4389 (
        .din(new_Jinkela_wire_6012),
        .dout(new_Jinkela_wire_6013)
    );

    bfr new_Jinkela_buffer_4429 (
        .din(new_Jinkela_wire_6069),
        .dout(new_Jinkela_wire_6070)
    );

    bfr new_Jinkela_buffer_4390 (
        .din(new_Jinkela_wire_6013),
        .dout(new_Jinkela_wire_6014)
    );

    bfr new_Jinkela_buffer_4410 (
        .din(new_Jinkela_wire_6041),
        .dout(new_Jinkela_wire_6042)
    );

    bfr new_Jinkela_buffer_4417 (
        .din(new_Jinkela_wire_6053),
        .dout(new_Jinkela_wire_6054)
    );

    spl2 new_Jinkela_splitter_631 (
        .a(_0715_),
        .b(new_Jinkela_wire_6094),
        .c(new_Jinkela_wire_6095)
    );

    bfr new_Jinkela_buffer_4418 (
        .din(new_Jinkela_wire_6054),
        .dout(new_Jinkela_wire_6055)
    );

    bfr new_Jinkela_buffer_4754 (
        .din(new_Jinkela_wire_6488),
        .dout(new_Jinkela_wire_6489)
    );

    bfr new_Jinkela_buffer_5550 (
        .din(new_Jinkela_wire_7491),
        .dout(new_Jinkela_wire_7492)
    );

    bfr new_Jinkela_buffer_4804 (
        .din(new_Jinkela_wire_6556),
        .dout(new_Jinkela_wire_6557)
    );

    bfr new_Jinkela_buffer_5612 (
        .din(new_net_2425),
        .dout(new_Jinkela_wire_7569)
    );

    bfr new_Jinkela_buffer_4755 (
        .din(new_Jinkela_wire_6489),
        .dout(new_Jinkela_wire_6490)
    );

    bfr new_Jinkela_buffer_5551 (
        .din(new_Jinkela_wire_7492),
        .dout(new_Jinkela_wire_7493)
    );

    bfr new_Jinkela_buffer_4766 (
        .din(new_Jinkela_wire_6514),
        .dout(new_Jinkela_wire_6515)
    );

    bfr new_Jinkela_buffer_5573 (
        .din(new_Jinkela_wire_7526),
        .dout(new_Jinkela_wire_7527)
    );

    bfr new_Jinkela_buffer_4756 (
        .din(new_Jinkela_wire_6490),
        .dout(new_Jinkela_wire_6491)
    );

    bfr new_Jinkela_buffer_5552 (
        .din(new_Jinkela_wire_7493),
        .dout(new_Jinkela_wire_7494)
    );

    spl2 new_Jinkela_splitter_756 (
        .a(_0942_),
        .b(new_Jinkela_wire_7595),
        .c(new_Jinkela_wire_7596)
    );

    bfr new_Jinkela_buffer_4757 (
        .din(new_Jinkela_wire_6491),
        .dout(new_Jinkela_wire_6492)
    );

    bfr new_Jinkela_buffer_5553 (
        .din(new_Jinkela_wire_7494),
        .dout(new_Jinkela_wire_7495)
    );

    bfr new_Jinkela_buffer_4767 (
        .din(new_Jinkela_wire_6515),
        .dout(new_Jinkela_wire_6516)
    );

    bfr new_Jinkela_buffer_5613 (
        .din(new_Jinkela_wire_7569),
        .dout(new_Jinkela_wire_7570)
    );

    bfr new_Jinkela_buffer_5574 (
        .din(new_Jinkela_wire_7527),
        .dout(new_Jinkela_wire_7528)
    );

    bfr new_Jinkela_buffer_4758 (
        .din(new_Jinkela_wire_6492),
        .dout(new_Jinkela_wire_6493)
    );

    bfr new_Jinkela_buffer_5554 (
        .din(new_Jinkela_wire_7495),
        .dout(new_Jinkela_wire_7496)
    );

    bfr new_Jinkela_buffer_4759 (
        .din(new_Jinkela_wire_6493),
        .dout(new_Jinkela_wire_6494)
    );

    bfr new_Jinkela_buffer_5555 (
        .din(new_Jinkela_wire_7496),
        .dout(new_Jinkela_wire_7497)
    );

    bfr new_Jinkela_buffer_4768 (
        .din(new_Jinkela_wire_6516),
        .dout(new_Jinkela_wire_6517)
    );

    bfr new_Jinkela_buffer_5575 (
        .din(new_Jinkela_wire_7528),
        .dout(new_Jinkela_wire_7529)
    );

    bfr new_Jinkela_buffer_4760 (
        .din(new_Jinkela_wire_6494),
        .dout(new_Jinkela_wire_6495)
    );

    bfr new_Jinkela_buffer_5556 (
        .din(new_Jinkela_wire_7497),
        .dout(new_Jinkela_wire_7498)
    );

    bfr new_Jinkela_buffer_4833 (
        .din(new_Jinkela_wire_6590),
        .dout(new_Jinkela_wire_6591)
    );

    bfr new_Jinkela_buffer_4807 (
        .din(new_Jinkela_wire_6564),
        .dout(new_Jinkela_wire_6565)
    );

    bfr new_Jinkela_buffer_5637 (
        .din(new_Jinkela_wire_7597),
        .dout(new_Jinkela_wire_7598)
    );

    bfr new_Jinkela_buffer_4769 (
        .din(new_Jinkela_wire_6517),
        .dout(new_Jinkela_wire_6518)
    );

    bfr new_Jinkela_buffer_5557 (
        .din(new_Jinkela_wire_7498),
        .dout(new_Jinkela_wire_7499)
    );

    bfr new_Jinkela_buffer_5614 (
        .din(new_Jinkela_wire_7570),
        .dout(new_Jinkela_wire_7571)
    );

    bfr new_Jinkela_buffer_4805 (
        .din(new_Jinkela_wire_6560),
        .dout(new_Jinkela_wire_6561)
    );

    bfr new_Jinkela_buffer_5576 (
        .din(new_Jinkela_wire_7529),
        .dout(new_Jinkela_wire_7530)
    );

    bfr new_Jinkela_buffer_4770 (
        .din(new_Jinkela_wire_6518),
        .dout(new_Jinkela_wire_6519)
    );

    bfr new_Jinkela_buffer_5558 (
        .din(new_Jinkela_wire_7499),
        .dout(new_Jinkela_wire_7500)
    );

    spl2 new_Jinkela_splitter_673 (
        .a(new_Jinkela_wire_6561),
        .b(new_Jinkela_wire_6562),
        .c(new_Jinkela_wire_6563)
    );

    bfr new_Jinkela_buffer_4771 (
        .din(new_Jinkela_wire_6519),
        .dout(new_Jinkela_wire_6520)
    );

    bfr new_Jinkela_buffer_5577 (
        .din(new_Jinkela_wire_7530),
        .dout(new_Jinkela_wire_7531)
    );

    bfr new_Jinkela_buffer_4808 (
        .din(new_Jinkela_wire_6565),
        .dout(new_Jinkela_wire_6566)
    );

    bfr new_Jinkela_buffer_4772 (
        .din(new_Jinkela_wire_6520),
        .dout(new_Jinkela_wire_6521)
    );

    bfr new_Jinkela_buffer_5615 (
        .din(new_Jinkela_wire_7571),
        .dout(new_Jinkela_wire_7572)
    );

    bfr new_Jinkela_buffer_5578 (
        .din(new_Jinkela_wire_7531),
        .dout(new_Jinkela_wire_7532)
    );

    spl2 new_Jinkela_splitter_675 (
        .a(new_Jinkela_wire_6624),
        .b(new_Jinkela_wire_6625),
        .c(new_Jinkela_wire_6626)
    );

    bfr new_Jinkela_buffer_4773 (
        .din(new_Jinkela_wire_6521),
        .dout(new_Jinkela_wire_6522)
    );

    spl2 new_Jinkela_splitter_758 (
        .a(_1224_),
        .b(new_Jinkela_wire_7605),
        .c(new_Jinkela_wire_7606)
    );

    bfr new_Jinkela_buffer_5579 (
        .din(new_Jinkela_wire_7532),
        .dout(new_Jinkela_wire_7533)
    );

    bfr new_Jinkela_buffer_4834 (
        .din(new_Jinkela_wire_6591),
        .dout(new_Jinkela_wire_6592)
    );

    bfr new_Jinkela_buffer_5636 (
        .din(new_Jinkela_wire_7596),
        .dout(new_Jinkela_wire_7597)
    );

    bfr new_Jinkela_buffer_4774 (
        .din(new_Jinkela_wire_6522),
        .dout(new_Jinkela_wire_6523)
    );

    bfr new_Jinkela_buffer_5616 (
        .din(new_Jinkela_wire_7572),
        .dout(new_Jinkela_wire_7573)
    );

    bfr new_Jinkela_buffer_5580 (
        .din(new_Jinkela_wire_7533),
        .dout(new_Jinkela_wire_7534)
    );

    bfr new_Jinkela_buffer_4809 (
        .din(new_Jinkela_wire_6566),
        .dout(new_Jinkela_wire_6567)
    );

    bfr new_Jinkela_buffer_4775 (
        .din(new_Jinkela_wire_6523),
        .dout(new_Jinkela_wire_6524)
    );

    bfr new_Jinkela_buffer_5642 (
        .din(_1046_),
        .dout(new_Jinkela_wire_7607)
    );

    bfr new_Jinkela_buffer_5581 (
        .din(new_Jinkela_wire_7534),
        .dout(new_Jinkela_wire_7535)
    );

    bfr new_Jinkela_buffer_4776 (
        .din(new_Jinkela_wire_6524),
        .dout(new_Jinkela_wire_6525)
    );

    bfr new_Jinkela_buffer_5617 (
        .din(new_Jinkela_wire_7573),
        .dout(new_Jinkela_wire_7574)
    );

    bfr new_Jinkela_buffer_5582 (
        .din(new_Jinkela_wire_7535),
        .dout(new_Jinkela_wire_7536)
    );

    bfr new_Jinkela_buffer_4810 (
        .din(new_Jinkela_wire_6567),
        .dout(new_Jinkela_wire_6568)
    );

    spl2 new_Jinkela_splitter_755 (
        .a(_1247_),
        .b(new_Jinkela_wire_7593),
        .c(new_Jinkela_wire_7594)
    );

    bfr new_Jinkela_buffer_5583 (
        .din(new_Jinkela_wire_7536),
        .dout(new_Jinkela_wire_7537)
    );

    bfr new_Jinkela_buffer_4777 (
        .din(new_Jinkela_wire_6525),
        .dout(new_Jinkela_wire_6526)
    );

    bfr new_Jinkela_buffer_4888 (
        .din(new_Jinkela_wire_6649),
        .dout(new_Jinkela_wire_6650)
    );

    bfr new_Jinkela_buffer_4835 (
        .din(new_Jinkela_wire_6592),
        .dout(new_Jinkela_wire_6593)
    );

    spl2 new_Jinkela_splitter_760 (
        .a(_0660_),
        .b(new_Jinkela_wire_7646),
        .c(new_Jinkela_wire_7647)
    );

    bfr new_Jinkela_buffer_4778 (
        .din(new_Jinkela_wire_6526),
        .dout(new_Jinkela_wire_6527)
    );

    bfr new_Jinkela_buffer_5618 (
        .din(new_Jinkela_wire_7574),
        .dout(new_Jinkela_wire_7575)
    );

    bfr new_Jinkela_buffer_5584 (
        .din(new_Jinkela_wire_7537),
        .dout(new_Jinkela_wire_7538)
    );

    bfr new_Jinkela_buffer_4811 (
        .din(new_Jinkela_wire_6568),
        .dout(new_Jinkela_wire_6569)
    );

    bfr new_Jinkela_buffer_4779 (
        .din(new_Jinkela_wire_6527),
        .dout(new_Jinkela_wire_6528)
    );

    bfr new_Jinkela_buffer_5585 (
        .din(new_Jinkela_wire_7538),
        .dout(new_Jinkela_wire_7539)
    );

    spl3L new_Jinkela_splitter_677 (
        .a(_0771_),
        .d(new_Jinkela_wire_6676),
        .b(new_Jinkela_wire_6677),
        .c(new_Jinkela_wire_6678)
    );

    bfr new_Jinkela_buffer_5679 (
        .din(_0246_),
        .dout(new_Jinkela_wire_7648)
    );

    bfr new_Jinkela_buffer_4780 (
        .din(new_Jinkela_wire_6528),
        .dout(new_Jinkela_wire_6529)
    );

    bfr new_Jinkela_buffer_5619 (
        .din(new_Jinkela_wire_7575),
        .dout(new_Jinkela_wire_7576)
    );

    bfr new_Jinkela_buffer_5586 (
        .din(new_Jinkela_wire_7539),
        .dout(new_Jinkela_wire_7540)
    );

    bfr new_Jinkela_buffer_4812 (
        .din(new_Jinkela_wire_6569),
        .dout(new_Jinkela_wire_6570)
    );

    bfr new_Jinkela_buffer_4781 (
        .din(new_Jinkela_wire_6529),
        .dout(new_Jinkela_wire_6530)
    );

    bfr new_Jinkela_buffer_5587 (
        .din(new_Jinkela_wire_7540),
        .dout(new_Jinkela_wire_7541)
    );

    bfr new_Jinkela_buffer_4867 (
        .din(new_Jinkela_wire_6628),
        .dout(new_Jinkela_wire_6629)
    );

    bfr new_Jinkela_buffer_4836 (
        .din(new_Jinkela_wire_6593),
        .dout(new_Jinkela_wire_6594)
    );

    bfr new_Jinkela_buffer_5643 (
        .din(new_Jinkela_wire_7607),
        .dout(new_Jinkela_wire_7608)
    );

    bfr new_Jinkela_buffer_4782 (
        .din(new_Jinkela_wire_6530),
        .dout(new_Jinkela_wire_6531)
    );

    bfr new_Jinkela_buffer_5620 (
        .din(new_Jinkela_wire_7576),
        .dout(new_Jinkela_wire_7577)
    );

    bfr new_Jinkela_buffer_5588 (
        .din(new_Jinkela_wire_7541),
        .dout(new_Jinkela_wire_7542)
    );

    bfr new_Jinkela_buffer_4813 (
        .din(new_Jinkela_wire_6570),
        .dout(new_Jinkela_wire_6571)
    );

    bfr new_Jinkela_buffer_1814 (
        .din(new_Jinkela_wire_2852),
        .dout(new_Jinkela_wire_2853)
    );

    bfr new_Jinkela_buffer_1800 (
        .din(new_Jinkela_wire_2833),
        .dout(new_Jinkela_wire_2834)
    );

    bfr new_Jinkela_buffer_1801 (
        .din(new_Jinkela_wire_2834),
        .dout(new_Jinkela_wire_2835)
    );

    bfr new_Jinkela_buffer_1822 (
        .din(new_Jinkela_wire_2877),
        .dout(new_Jinkela_wire_2878)
    );

    bfr new_Jinkela_buffer_1844 (
        .din(new_net_2453),
        .dout(new_Jinkela_wire_2903)
    );

    bfr new_Jinkela_buffer_1802 (
        .din(new_Jinkela_wire_2835),
        .dout(new_Jinkela_wire_2836)
    );

    bfr new_Jinkela_buffer_1820 (
        .din(_0321_),
        .dout(new_Jinkela_wire_2876)
    );

    bfr new_Jinkela_buffer_1803 (
        .din(new_Jinkela_wire_2836),
        .dout(new_Jinkela_wire_2837)
    );

    bfr new_Jinkela_buffer_1843 (
        .din(_0609_),
        .dout(new_Jinkela_wire_2899)
    );

    bfr new_Jinkela_buffer_1804 (
        .din(new_Jinkela_wire_2837),
        .dout(new_Jinkela_wire_2838)
    );

    spl2 new_Jinkela_splitter_391 (
        .a(new_Jinkela_wire_2863),
        .b(new_Jinkela_wire_2864),
        .c(new_Jinkela_wire_2865)
    );

    bfr new_Jinkela_buffer_1805 (
        .din(new_Jinkela_wire_2838),
        .dout(new_Jinkela_wire_2839)
    );

    spl4L new_Jinkela_splitter_392 (
        .a(new_Jinkela_wire_2866),
        .d(new_Jinkela_wire_2867),
        .e(new_Jinkela_wire_2868),
        .b(new_Jinkela_wire_2869),
        .c(new_Jinkela_wire_2870)
    );

    bfr new_Jinkela_buffer_1806 (
        .din(new_Jinkela_wire_2839),
        .dout(new_Jinkela_wire_2840)
    );

    spl4L new_Jinkela_splitter_393 (
        .a(new_Jinkela_wire_2871),
        .d(new_Jinkela_wire_2872),
        .e(new_Jinkela_wire_2873),
        .b(new_Jinkela_wire_2874),
        .c(new_Jinkela_wire_2875)
    );

    bfr new_Jinkela_buffer_1821 (
        .din(new_Jinkela_wire_2876),
        .dout(new_Jinkela_wire_2877)
    );

    spl3L new_Jinkela_splitter_395 (
        .a(_0953_),
        .d(new_Jinkela_wire_2904),
        .b(new_Jinkela_wire_2905),
        .c(new_Jinkela_wire_2906)
    );

    bfr new_Jinkela_buffer_1823 (
        .din(new_Jinkela_wire_2878),
        .dout(new_Jinkela_wire_2879)
    );

    spl3L new_Jinkela_splitter_398 (
        .a(_0637_),
        .d(new_Jinkela_wire_2926),
        .b(new_Jinkela_wire_2927),
        .c(new_Jinkela_wire_2928)
    );

    spl2 new_Jinkela_splitter_397 (
        .a(_0836_),
        .b(new_Jinkela_wire_2924),
        .c(new_Jinkela_wire_2925)
    );

    bfr new_Jinkela_buffer_1824 (
        .din(new_Jinkela_wire_2879),
        .dout(new_Jinkela_wire_2880)
    );

    spl3L new_Jinkela_splitter_394 (
        .a(new_Jinkela_wire_2899),
        .d(new_Jinkela_wire_2900),
        .b(new_Jinkela_wire_2901),
        .c(new_Jinkela_wire_2902)
    );

    bfr new_Jinkela_buffer_1825 (
        .din(new_Jinkela_wire_2880),
        .dout(new_Jinkela_wire_2881)
    );

    spl2 new_Jinkela_splitter_399 (
        .a(new_Jinkela_wire_2928),
        .b(new_Jinkela_wire_2929),
        .c(new_Jinkela_wire_2930)
    );

    bfr new_Jinkela_buffer_1826 (
        .din(new_Jinkela_wire_2881),
        .dout(new_Jinkela_wire_2882)
    );

    bfr new_Jinkela_buffer_1845 (
        .din(new_Jinkela_wire_2906),
        .dout(new_Jinkela_wire_2907)
    );

    bfr new_Jinkela_buffer_1827 (
        .din(new_Jinkela_wire_2882),
        .dout(new_Jinkela_wire_2883)
    );

    bfr new_Jinkela_buffer_1860 (
        .din(_0002_),
        .dout(new_Jinkela_wire_2931)
    );

    bfr new_Jinkela_buffer_1828 (
        .din(new_Jinkela_wire_2883),
        .dout(new_Jinkela_wire_2884)
    );

    bfr new_Jinkela_buffer_1846 (
        .din(new_Jinkela_wire_2907),
        .dout(new_Jinkela_wire_2908)
    );

    bfr new_Jinkela_buffer_1829 (
        .din(new_Jinkela_wire_2884),
        .dout(new_Jinkela_wire_2885)
    );

    bfr new_Jinkela_buffer_1861 (
        .din(new_Jinkela_wire_2931),
        .dout(new_Jinkela_wire_2932)
    );

    bfr new_Jinkela_buffer_1830 (
        .din(new_Jinkela_wire_2885),
        .dout(new_Jinkela_wire_2886)
    );

    bfr new_Jinkela_buffer_1847 (
        .din(new_Jinkela_wire_2908),
        .dout(new_Jinkela_wire_2909)
    );

    bfr new_Jinkela_buffer_1831 (
        .din(new_Jinkela_wire_2886),
        .dout(new_Jinkela_wire_2887)
    );

    bfr new_Jinkela_buffer_1832 (
        .din(new_Jinkela_wire_2887),
        .dout(new_Jinkela_wire_2888)
    );

    bfr new_Jinkela_buffer_1848 (
        .din(new_Jinkela_wire_2909),
        .dout(new_Jinkela_wire_2910)
    );

    bfr new_Jinkela_buffer_1833 (
        .din(new_Jinkela_wire_2888),
        .dout(new_Jinkela_wire_2889)
    );

    bfr new_Jinkela_buffer_1871 (
        .din(new_net_2349),
        .dout(new_Jinkela_wire_2944)
    );

    bfr new_Jinkela_buffer_1869 (
        .din(_1098_),
        .dout(new_Jinkela_wire_2940)
    );

    bfr new_Jinkela_buffer_1834 (
        .din(new_Jinkela_wire_2889),
        .dout(new_Jinkela_wire_2890)
    );

    bfr new_Jinkela_buffer_1849 (
        .din(new_Jinkela_wire_2910),
        .dout(new_Jinkela_wire_2911)
    );

    spl2 new_Jinkela_splitter_289 (
        .a(new_Jinkela_wire_1577),
        .b(new_Jinkela_wire_1578),
        .c(new_Jinkela_wire_1579)
    );

    or_bi _2033_ (
        .a(new_Jinkela_wire_4339),
        .b(new_Jinkela_wire_2419),
        .c(_0074_)
    );

    bfr new_Jinkela_buffer_4338 (
        .din(new_Jinkela_wire_5961),
        .dout(new_Jinkela_wire_5962)
    );

    spl4L new_Jinkela_splitter_292 (
        .a(new_Jinkela_wire_1587),
        .d(new_Jinkela_wire_1588),
        .e(new_Jinkela_wire_1589),
        .b(new_Jinkela_wire_1590),
        .c(new_Jinkela_wire_1591)
    );

    and_bi _2034_ (
        .a(new_Jinkela_wire_4338),
        .b(new_Jinkela_wire_2417),
        .c(_0075_)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    spl2 new_Jinkela_splitter_625 (
        .a(new_Jinkela_wire_6024),
        .b(new_Jinkela_wire_6025),
        .c(new_Jinkela_wire_6026)
    );

    or_bi _2035_ (
        .a(new_Jinkela_wire_5730),
        .b(new_Jinkela_wire_7520),
        .c(_0076_)
    );

    bfr new_Jinkela_buffer_4339 (
        .din(new_Jinkela_wire_5962),
        .dout(new_Jinkela_wire_5963)
    );

    spl3L new_Jinkela_splitter_291 (
        .a(new_Jinkela_wire_1583),
        .d(new_Jinkela_wire_1584),
        .b(new_Jinkela_wire_1585),
        .c(new_Jinkela_wire_1586)
    );

    and_ii _2036_ (
        .a(new_Jinkela_wire_6258),
        .b(new_Jinkela_wire_5300),
        .c(_0077_)
    );

    bfr new_Jinkela_buffer_4358 (
        .din(new_Jinkela_wire_5981),
        .dout(new_Jinkela_wire_5982)
    );

    bfr new_Jinkela_buffer_782 (
        .din(G79),
        .dout(new_Jinkela_wire_1602)
    );

    and_bb _2037_ (
        .a(new_Jinkela_wire_6259),
        .b(new_Jinkela_wire_5301),
        .c(_0078_)
    );

    bfr new_Jinkela_buffer_785 (
        .din(G25),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_4340 (
        .din(new_Jinkela_wire_5963),
        .dout(new_Jinkela_wire_5964)
    );

    and_ii _2038_ (
        .a(_0078_),
        .b(_0077_),
        .c(_0079_)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_4395 (
        .din(new_Jinkela_wire_6026),
        .dout(new_Jinkela_wire_6027)
    );

    or_bb _2039_ (
        .a(new_Jinkela_wire_6768),
        .b(new_Jinkela_wire_2316),
        .c(_0080_)
    );

    bfr new_Jinkela_buffer_4341 (
        .din(new_Jinkela_wire_5964),
        .dout(new_Jinkela_wire_5965)
    );

    spl2 new_Jinkela_splitter_296 (
        .a(_0910_),
        .b(new_Jinkela_wire_1612),
        .c(new_Jinkela_wire_1614)
    );

    and_bb _2040_ (
        .a(new_Jinkela_wire_6769),
        .b(new_Jinkela_wire_2317),
        .c(_0081_)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_4359 (
        .din(new_Jinkela_wire_5982),
        .dout(new_Jinkela_wire_5983)
    );

    or_bb _2041_ (
        .a(_0081_),
        .b(new_Jinkela_wire_7696),
        .c(_0082_)
    );

    bfr new_Jinkela_buffer_4342 (
        .din(new_Jinkela_wire_5965),
        .dout(new_Jinkela_wire_5966)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    and_bi _2042_ (
        .a(new_Jinkela_wire_7432),
        .b(_0082_),
        .c(_0083_)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_4393 (
        .din(new_Jinkela_wire_6022),
        .dout(new_Jinkela_wire_6023)
    );

    or_bb _2043_ (
        .a(_0083_),
        .b(new_Jinkela_wire_4853),
        .c(_0084_)
    );

    bfr new_Jinkela_buffer_789 (
        .din(_0632_),
        .dout(new_Jinkela_wire_1619)
    );

    bfr new_Jinkela_buffer_4343 (
        .din(new_Jinkela_wire_5966),
        .dout(new_Jinkela_wire_5967)
    );

    and_bi _2044_ (
        .a(_0028_),
        .b(new_Jinkela_wire_4546),
        .c(_0085_)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_4360 (
        .din(new_Jinkela_wire_5983),
        .dout(new_Jinkela_wire_5984)
    );

    and_bi _2045_ (
        .a(new_Jinkela_wire_115),
        .b(new_Jinkela_wire_1403),
        .c(_0086_)
    );

    bfr new_Jinkela_buffer_4344 (
        .din(new_Jinkela_wire_5967),
        .dout(new_Jinkela_wire_5968)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    or_bb _2046_ (
        .a(new_Jinkela_wire_1943),
        .b(new_Jinkela_wire_1681),
        .c(_0087_)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1607),
        .dout(new_Jinkela_wire_1608)
    );

    and_bi _2047_ (
        .a(new_Jinkela_wire_493),
        .b(new_Jinkela_wire_3751),
        .c(_0088_)
    );

    bfr new_Jinkela_buffer_4345 (
        .din(new_Jinkela_wire_5968),
        .dout(new_Jinkela_wire_5969)
    );

    spl2 new_Jinkela_splitter_294 (
        .a(new_Jinkela_wire_1604),
        .b(new_Jinkela_wire_1605),
        .c(new_Jinkela_wire_1606)
    );

    or_bb _2048_ (
        .a(_0088_),
        .b(new_Jinkela_wire_1747),
        .c(_0089_)
    );

    bfr new_Jinkela_buffer_4361 (
        .din(new_Jinkela_wire_5984),
        .dout(new_Jinkela_wire_5985)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1608),
        .dout(new_Jinkela_wire_1609)
    );

    or_bb _2049_ (
        .a(new_Jinkela_wire_1977),
        .b(_1227_),
        .c(_0090_)
    );

    bfr new_Jinkela_buffer_4346 (
        .din(new_Jinkela_wire_5969),
        .dout(new_Jinkela_wire_5970)
    );

    or_bb _2050_ (
        .a(new_Jinkela_wire_453),
        .b(new_Jinkela_wire_835),
        .c(_0091_)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    bfr new_Jinkela_buffer_4411 (
        .din(new_Jinkela_wire_6045),
        .dout(new_Jinkela_wire_6046)
    );

    spl4L new_Jinkela_splitter_297 (
        .a(new_Jinkela_wire_1614),
        .d(new_Jinkela_wire_1615),
        .e(new_Jinkela_wire_1616),
        .b(new_Jinkela_wire_1617),
        .c(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_4431 (
        .din(new_net_2357),
        .dout(new_Jinkela_wire_6074)
    );

    and_bi _2051_ (
        .a(new_Jinkela_wire_1605),
        .b(new_Jinkela_wire_7921),
        .c(_0092_)
    );

    spl2 new_Jinkela_splitter_298 (
        .a(_0963_),
        .b(new_Jinkela_wire_1625),
        .c(new_Jinkela_wire_1628)
    );

    bfr new_Jinkela_buffer_4347 (
        .din(new_Jinkela_wire_5970),
        .dout(new_Jinkela_wire_5971)
    );

    spl2 new_Jinkela_splitter_295 (
        .a(new_Jinkela_wire_1609),
        .b(new_Jinkela_wire_1610),
        .c(new_Jinkela_wire_1611)
    );

    or_bi _2052_ (
        .a(new_Jinkela_wire_837),
        .b(new_Jinkela_wire_454),
        .c(_0093_)
    );

    bfr new_Jinkela_buffer_4362 (
        .din(new_Jinkela_wire_5985),
        .dout(new_Jinkela_wire_5986)
    );

    and_bi _2053_ (
        .a(new_Jinkela_wire_246),
        .b(new_Jinkela_wire_6135),
        .c(_0094_)
    );

    bfr new_Jinkela_buffer_4348 (
        .din(new_Jinkela_wire_5971),
        .dout(new_Jinkela_wire_5972)
    );

    or_bb _2054_ (
        .a(_0094_),
        .b(_0092_),
        .c(_0095_)
    );

    spl2 new_Jinkela_splitter_630 (
        .a(_0021_),
        .b(new_Jinkela_wire_6072),
        .c(new_Jinkela_wire_6073)
    );

    bfr new_Jinkela_buffer_795 (
        .din(_1047_),
        .dout(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_4396 (
        .din(new_Jinkela_wire_6027),
        .dout(new_Jinkela_wire_6028)
    );

    and_bi _2055_ (
        .a(_0090_),
        .b(new_Jinkela_wire_3249),
        .c(_0096_)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1619),
        .dout(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_4349 (
        .din(new_Jinkela_wire_5972),
        .dout(new_Jinkela_wire_5973)
    );

    or_bb _2056_ (
        .a(_0096_),
        .b(new_Jinkela_wire_7644),
        .c(new_net_2453)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1620),
        .dout(new_Jinkela_wire_1621)
    );

    bfr new_Jinkela_buffer_4363 (
        .din(new_Jinkela_wire_5986),
        .dout(new_Jinkela_wire_5987)
    );

    inv _2057_ (
        .din(new_Jinkela_wire_777),
        .dout(_0097_)
    );

    bfr new_Jinkela_buffer_825 (
        .din(_0335_),
        .dout(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_4350 (
        .din(new_Jinkela_wire_5973),
        .dout(new_Jinkela_wire_5974)
    );

    and_bi _2058_ (
        .a(new_Jinkela_wire_6846),
        .b(new_Jinkela_wire_3414),
        .c(_0098_)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1621),
        .dout(new_Jinkela_wire_1622)
    );

    bfr new_Jinkela_buffer_4426 (
        .din(new_Jinkela_wire_6066),
        .dout(new_Jinkela_wire_6067)
    );

    inv _2059_ (
        .din(new_Jinkela_wire_501),
        .dout(_0099_)
    );

    bfr new_Jinkela_buffer_4364 (
        .din(new_Jinkela_wire_5987),
        .dout(new_Jinkela_wire_5988)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1677),
        .dout(new_Jinkela_wire_1678)
    );

    and_bi _2060_ (
        .a(new_Jinkela_wire_818),
        .b(new_Jinkela_wire_3752),
        .c(_0100_)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1622),
        .dout(new_Jinkela_wire_1623)
    );

    bfr new_Jinkela_buffer_4397 (
        .din(new_Jinkela_wire_6028),
        .dout(new_Jinkela_wire_6029)
    );

    or_bb _2061_ (
        .a(_0100_),
        .b(new_Jinkela_wire_5592),
        .c(_0101_)
    );

    spl2 new_Jinkela_splitter_299 (
        .a(new_Jinkela_wire_1625),
        .b(new_Jinkela_wire_1626),
        .c(new_Jinkela_wire_1627)
    );

    bfr new_Jinkela_buffer_4365 (
        .din(new_Jinkela_wire_5988),
        .dout(new_Jinkela_wire_5989)
    );

    or_bb _2062_ (
        .a(new_Jinkela_wire_6195),
        .b(_0098_),
        .c(_0102_)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1623),
        .dout(new_Jinkela_wire_1624)
    );

    or_bb _2063_ (
        .a(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_779),
        .c(_0103_)
    );

    spl4L new_Jinkela_splitter_300 (
        .a(new_Jinkela_wire_1628),
        .d(new_Jinkela_wire_1629),
        .e(new_Jinkela_wire_1630),
        .b(new_Jinkela_wire_1631),
        .c(new_Jinkela_wire_1632)
    );

    bfr new_Jinkela_buffer_4366 (
        .din(new_Jinkela_wire_5989),
        .dout(new_Jinkela_wire_5990)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_1676),
        .dout(new_Jinkela_wire_1677)
    );

    and_bi _2064_ (
        .a(new_Jinkela_wire_1606),
        .b(new_Jinkela_wire_3383),
        .c(_0104_)
    );

    spl2 new_Jinkela_splitter_627 (
        .a(new_Jinkela_wire_6046),
        .b(new_Jinkela_wire_6047),
        .c(new_Jinkela_wire_6048)
    );

    bfr new_Jinkela_buffer_4398 (
        .din(new_Jinkela_wire_6029),
        .dout(new_Jinkela_wire_6030)
    );

    or_bi _2065_ (
        .a(new_Jinkela_wire_500),
        .b(new_Jinkela_wire_778),
        .c(_0105_)
    );

    bfr new_Jinkela_buffer_4367 (
        .din(new_Jinkela_wire_5990),
        .dout(new_Jinkela_wire_5991)
    );

    and_bi _2066_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_4026),
        .c(_0106_)
    );

    spl2 new_Jinkela_splitter_310 (
        .a(_0085_),
        .b(new_Jinkela_wire_1681),
        .c(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_822 (
        .din(_1182_),
        .dout(new_Jinkela_wire_1676)
    );

    or_bb _2067_ (
        .a(_0106_),
        .b(_0104_),
        .c(_0107_)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_4368 (
        .din(new_Jinkela_wire_5991),
        .dout(new_Jinkela_wire_5992)
    );

    and_bi _2068_ (
        .a(_0102_),
        .b(new_Jinkela_wire_5113),
        .c(_0108_)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    bfr new_Jinkela_buffer_4399 (
        .din(new_Jinkela_wire_6030),
        .dout(new_Jinkela_wire_6031)
    );

    or_bb _2069_ (
        .a(_0108_),
        .b(new_Jinkela_wire_7645),
        .c(new_net_2357)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    bfr new_Jinkela_buffer_4369 (
        .din(new_Jinkela_wire_5992),
        .dout(new_Jinkela_wire_5993)
    );

    and_bb _2070_ (
        .a(new_Jinkela_wire_90),
        .b(new_Jinkela_wire_1146),
        .c(new_net_2435)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1636),
        .dout(new_Jinkela_wire_1637)
    );

    spl2 new_Jinkela_splitter_309 (
        .a(new_Jinkela_wire_1678),
        .b(new_Jinkela_wire_1679),
        .c(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_4412 (
        .din(new_Jinkela_wire_6048),
        .dout(new_Jinkela_wire_6049)
    );

    and_ii _2071_ (
        .a(new_Jinkela_wire_524),
        .b(new_Jinkela_wire_1395),
        .c(_0109_)
    );

    bfr new_Jinkela_buffer_874 (
        .din(_0930_),
        .dout(new_Jinkela_wire_1752)
    );

    bfr new_Jinkela_buffer_4370 (
        .din(new_Jinkela_wire_5993),
        .dout(new_Jinkela_wire_5994)
    );

    and_bb _2072_ (
        .a(new_Jinkela_wire_523),
        .b(new_Jinkela_wire_1393),
        .c(_0110_)
    );

    bfr new_Jinkela_buffer_849 (
        .din(_1228_),
        .dout(new_Jinkela_wire_1709)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_1635),
        .dout(new_Jinkela_wire_1636)
    );

    bfr new_Jinkela_buffer_4400 (
        .din(new_Jinkela_wire_6031),
        .dout(new_Jinkela_wire_6032)
    );

    and_ii _2073_ (
        .a(_0110_),
        .b(_0109_),
        .c(_0111_)
    );

    bfr new_Jinkela_buffer_4371 (
        .din(new_Jinkela_wire_5994),
        .dout(new_Jinkela_wire_5995)
    );

    spl2 new_Jinkela_splitter_311 (
        .a(_1108_),
        .b(new_Jinkela_wire_1683),
        .c(new_Jinkela_wire_1684)
    );

    and_bi _2074_ (
        .a(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_826),
        .c(_0112_)
    );

    or_bb _1319_ (
        .a(_0624_),
        .b(new_Jinkela_wire_6140),
        .c(_0625_)
    );

    bfr new_Jinkela_buffer_4783 (
        .din(new_Jinkela_wire_6531),
        .dout(new_Jinkela_wire_6532)
    );

    or_ii _1320_ (
        .a(new_Jinkela_wire_1586),
        .b(new_Jinkela_wire_290),
        .c(_0626_)
    );

    bfr new_Jinkela_buffer_4862 (
        .din(_0153_),
        .dout(new_Jinkela_wire_6622)
    );

    and_bi _1321_ (
        .a(new_Jinkela_wire_1283),
        .b(new_Jinkela_wire_287),
        .c(_0627_)
    );

    bfr new_Jinkela_buffer_4784 (
        .din(new_Jinkela_wire_6532),
        .dout(new_Jinkela_wire_6533)
    );

    and_bi _1322_ (
        .a(_0626_),
        .b(_0627_),
        .c(_0628_)
    );

    bfr new_Jinkela_buffer_4814 (
        .din(new_Jinkela_wire_6571),
        .dout(new_Jinkela_wire_6572)
    );

    and_bi _1323_ (
        .a(new_Jinkela_wire_6141),
        .b(_0628_),
        .c(_0629_)
    );

    bfr new_Jinkela_buffer_4785 (
        .din(new_Jinkela_wire_6533),
        .dout(new_Jinkela_wire_6534)
    );

    and_bi _1324_ (
        .a(_0625_),
        .b(_0629_),
        .c(_0630_)
    );

    bfr new_Jinkela_buffer_4865 (
        .din(new_net_2371),
        .dout(new_Jinkela_wire_6627)
    );

    and_bi _1325_ (
        .a(new_Jinkela_wire_1057),
        .b(new_Jinkela_wire_6376),
        .c(_0631_)
    );

    bfr new_Jinkela_buffer_4786 (
        .din(new_Jinkela_wire_6534),
        .dout(new_Jinkela_wire_6535)
    );

    or_bb _1326_ (
        .a(_0631_),
        .b(new_Jinkela_wire_4832),
        .c(_0632_)
    );

    bfr new_Jinkela_buffer_4815 (
        .din(new_Jinkela_wire_6572),
        .dout(new_Jinkela_wire_6573)
    );

    and_bi _1327_ (
        .a(_0621_),
        .b(new_Jinkela_wire_1624),
        .c(_0633_)
    );

    bfr new_Jinkela_buffer_4787 (
        .din(new_Jinkela_wire_6535),
        .dout(new_Jinkela_wire_6536)
    );

    and_ii _1328_ (
        .a(_0633_),
        .b(new_Jinkela_wire_5295),
        .c(new_net_12)
    );

    bfr new_Jinkela_buffer_4828 (
        .din(new_Jinkela_wire_6585),
        .dout(new_Jinkela_wire_6586)
    );

    and_bi _1329_ (
        .a(new_Jinkela_wire_35),
        .b(new_Jinkela_wire_6688),
        .c(_0634_)
    );

    bfr new_Jinkela_buffer_4788 (
        .din(new_Jinkela_wire_6536),
        .dout(new_Jinkela_wire_6537)
    );

    or_ii _1330_ (
        .a(new_Jinkela_wire_20),
        .b(new_Jinkela_wire_752),
        .c(_0635_)
    );

    bfr new_Jinkela_buffer_4816 (
        .din(new_Jinkela_wire_6573),
        .dout(new_Jinkela_wire_6574)
    );

    and_bi _1331_ (
        .a(new_Jinkela_wire_65),
        .b(new_Jinkela_wire_6),
        .c(_0636_)
    );

    bfr new_Jinkela_buffer_4789 (
        .din(new_Jinkela_wire_6537),
        .dout(new_Jinkela_wire_6538)
    );

    and_bi _1332_ (
        .a(_0635_),
        .b(new_Jinkela_wire_2092),
        .c(_0637_)
    );

    bfr new_Jinkela_buffer_4887 (
        .din(new_net_2421),
        .dout(new_Jinkela_wire_6649)
    );

    and_bi _1333_ (
        .a(new_Jinkela_wire_546),
        .b(new_Jinkela_wire_2926),
        .c(_0638_)
    );

    bfr new_Jinkela_buffer_4790 (
        .din(new_Jinkela_wire_6538),
        .dout(new_Jinkela_wire_6539)
    );

    and_bi _1334_ (
        .a(new_Jinkela_wire_2927),
        .b(new_Jinkela_wire_547),
        .c(_0639_)
    );

    bfr new_Jinkela_buffer_4817 (
        .din(new_Jinkela_wire_6574),
        .dout(new_Jinkela_wire_6575)
    );

    or_bb _1335_ (
        .a(new_Jinkela_wire_2204),
        .b(new_Jinkela_wire_7036),
        .c(_0640_)
    );

    bfr new_Jinkela_buffer_4791 (
        .din(new_Jinkela_wire_6539),
        .dout(new_Jinkela_wire_6540)
    );

    and_bi _1336_ (
        .a(new_Jinkela_wire_1413),
        .b(new_Jinkela_wire_7206),
        .c(_0641_)
    );

    bfr new_Jinkela_buffer_4829 (
        .din(new_Jinkela_wire_6586),
        .dout(new_Jinkela_wire_6587)
    );

    and_bi _1337_ (
        .a(new_Jinkela_wire_7207),
        .b(new_Jinkela_wire_1414),
        .c(_0642_)
    );

    bfr new_Jinkela_buffer_4792 (
        .din(new_Jinkela_wire_6540),
        .dout(new_Jinkela_wire_6541)
    );

    and_ii _1338_ (
        .a(new_Jinkela_wire_2779),
        .b(new_Jinkela_wire_5864),
        .c(_0643_)
    );

    bfr new_Jinkela_buffer_4818 (
        .din(new_Jinkela_wire_6575),
        .dout(new_Jinkela_wire_6576)
    );

    or_bb _1339_ (
        .a(new_Jinkela_wire_4606),
        .b(new_Jinkela_wire_1067),
        .c(_0644_)
    );

    bfr new_Jinkela_buffer_4793 (
        .din(new_Jinkela_wire_6541),
        .dout(new_Jinkela_wire_6542)
    );

    inv _1340_ (
        .din(new_Jinkela_wire_540),
        .dout(_0645_)
    );

    bfr new_Jinkela_buffer_4863 (
        .din(new_Jinkela_wire_6622),
        .dout(new_Jinkela_wire_6623)
    );

    or_bb _1341_ (
        .a(new_Jinkela_wire_754),
        .b(new_Jinkela_wire_316),
        .c(_0646_)
    );

    bfr new_Jinkela_buffer_4794 (
        .din(new_Jinkela_wire_6542),
        .dout(new_Jinkela_wire_6543)
    );

    and_bi _1342_ (
        .a(new_Jinkela_wire_748),
        .b(new_Jinkela_wire_214),
        .c(_0647_)
    );

    bfr new_Jinkela_buffer_4819 (
        .din(new_Jinkela_wire_6576),
        .dout(new_Jinkela_wire_6577)
    );

    and_bi _1343_ (
        .a(_0646_),
        .b(_0647_),
        .c(_0648_)
    );

    bfr new_Jinkela_buffer_4795 (
        .din(new_Jinkela_wire_6543),
        .dout(new_Jinkela_wire_6544)
    );

    or_bb _1344_ (
        .a(_0648_),
        .b(new_Jinkela_wire_6188),
        .c(_0649_)
    );

    bfr new_Jinkela_buffer_4830 (
        .din(new_Jinkela_wire_6587),
        .dout(new_Jinkela_wire_6588)
    );

    or_ii _1345_ (
        .a(new_Jinkela_wire_1585),
        .b(new_Jinkela_wire_750),
        .c(_0650_)
    );

    bfr new_Jinkela_buffer_4796 (
        .din(new_Jinkela_wire_6544),
        .dout(new_Jinkela_wire_6545)
    );

    and_bi _1346_ (
        .a(new_Jinkela_wire_1290),
        .b(new_Jinkela_wire_753),
        .c(_0651_)
    );

    bfr new_Jinkela_buffer_4820 (
        .din(new_Jinkela_wire_6577),
        .dout(new_Jinkela_wire_6578)
    );

    and_bi _1347_ (
        .a(_0650_),
        .b(_0651_),
        .c(_0652_)
    );

    bfr new_Jinkela_buffer_4797 (
        .din(new_Jinkela_wire_6545),
        .dout(new_Jinkela_wire_6546)
    );

    and_bi _1348_ (
        .a(new_Jinkela_wire_6190),
        .b(_0652_),
        .c(_0653_)
    );

    bfr new_Jinkela_buffer_4866 (
        .din(new_Jinkela_wire_6627),
        .dout(new_Jinkela_wire_6628)
    );

    and_bi _1349_ (
        .a(_0649_),
        .b(_0653_),
        .c(_0654_)
    );

    bfr new_Jinkela_buffer_4798 (
        .din(new_Jinkela_wire_6546),
        .dout(new_Jinkela_wire_6547)
    );

    and_bi _1350_ (
        .a(new_Jinkela_wire_1049),
        .b(new_Jinkela_wire_6554),
        .c(_0655_)
    );

    bfr new_Jinkela_buffer_4821 (
        .din(new_Jinkela_wire_6578),
        .dout(new_Jinkela_wire_6579)
    );

    or_bb _1351_ (
        .a(_0655_),
        .b(new_Jinkela_wire_4833),
        .c(_0656_)
    );

    bfr new_Jinkela_buffer_4799 (
        .din(new_Jinkela_wire_6547),
        .dout(new_Jinkela_wire_6548)
    );

    and_bi _1352_ (
        .a(_0644_),
        .b(new_Jinkela_wire_4762),
        .c(_0657_)
    );

    bfr new_Jinkela_buffer_4831 (
        .din(new_Jinkela_wire_6588),
        .dout(new_Jinkela_wire_6589)
    );

    and_ii _1353_ (
        .a(_0657_),
        .b(new_Jinkela_wire_4463),
        .c(new_net_3)
    );

    bfr new_Jinkela_buffer_4822 (
        .din(new_Jinkela_wire_6579),
        .dout(new_Jinkela_wire_6580)
    );

    and_bi _1354_ (
        .a(new_Jinkela_wire_842),
        .b(new_Jinkela_wire_6681),
        .c(_0658_)
    );

    bfr new_Jinkela_buffer_4864 (
        .din(new_Jinkela_wire_6623),
        .dout(new_Jinkela_wire_6624)
    );

    and_ii _1355_ (
        .a(new_Jinkela_wire_1348),
        .b(new_Jinkela_wire_880),
        .c(_0659_)
    );

    bfr new_Jinkela_buffer_4823 (
        .din(new_Jinkela_wire_6580),
        .dout(new_Jinkela_wire_6581)
    );

    and_bi _1356_ (
        .a(new_Jinkela_wire_1110),
        .b(new_Jinkela_wire_4167),
        .c(_0660_)
    );

    bfr new_Jinkela_buffer_4832 (
        .din(new_Jinkela_wire_6589),
        .dout(new_Jinkela_wire_6590)
    );

    and_bi _1357_ (
        .a(new_Jinkela_wire_4168),
        .b(new_Jinkela_wire_1111),
        .c(_0661_)
    );

    bfr new_Jinkela_buffer_4824 (
        .din(new_Jinkela_wire_6581),
        .dout(new_Jinkela_wire_6582)
    );

    and_ii _1358_ (
        .a(new_Jinkela_wire_3820),
        .b(new_Jinkela_wire_7646),
        .c(_0662_)
    );

    bfr new_Jinkela_buffer_4909 (
        .din(_0127_),
        .dout(new_Jinkela_wire_6671)
    );

    inv _1359_ (
        .din(new_Jinkela_wire_1128),
        .dout(_0663_)
    );

    bfr new_Jinkela_buffer_4825 (
        .din(new_Jinkela_wire_6582),
        .dout(new_Jinkela_wire_6583)
    );

    and_bb _1360_ (
        .a(new_Jinkela_wire_436),
        .b(new_Jinkela_wire_878),
        .c(_0664_)
    );

    bfr new_Jinkela_buffer_4827 (
        .din(new_net_27),
        .dout(new_Jinkela_wire_6585)
    );

    bfr new_Jinkela_buffer_5638 (
        .din(new_Jinkela_wire_7598),
        .dout(new_Jinkela_wire_7599)
    );

    bfr new_Jinkela_buffer_5589 (
        .din(new_Jinkela_wire_7542),
        .dout(new_Jinkela_wire_7543)
    );

    bfr new_Jinkela_buffer_5621 (
        .din(new_Jinkela_wire_7577),
        .dout(new_Jinkela_wire_7578)
    );

    bfr new_Jinkela_buffer_5590 (
        .din(new_Jinkela_wire_7543),
        .dout(new_Jinkela_wire_7544)
    );

    bfr new_Jinkela_buffer_5591 (
        .din(new_Jinkela_wire_7544),
        .dout(new_Jinkela_wire_7545)
    );

    spl2 new_Jinkela_splitter_763 (
        .a(_0135_),
        .b(new_Jinkela_wire_7654),
        .c(new_Jinkela_wire_7655)
    );

    bfr new_Jinkela_buffer_5622 (
        .din(new_Jinkela_wire_7578),
        .dout(new_Jinkela_wire_7579)
    );

    bfr new_Jinkela_buffer_5592 (
        .din(new_Jinkela_wire_7545),
        .dout(new_Jinkela_wire_7546)
    );

    spl2 new_Jinkela_splitter_757 (
        .a(new_Jinkela_wire_7599),
        .b(new_Jinkela_wire_7600),
        .c(new_Jinkela_wire_7601)
    );

    bfr new_Jinkela_buffer_5593 (
        .din(new_Jinkela_wire_7546),
        .dout(new_Jinkela_wire_7547)
    );

    bfr new_Jinkela_buffer_5623 (
        .din(new_Jinkela_wire_7579),
        .dout(new_Jinkela_wire_7580)
    );

    bfr new_Jinkela_buffer_5594 (
        .din(new_Jinkela_wire_7547),
        .dout(new_Jinkela_wire_7548)
    );

    bfr new_Jinkela_buffer_5639 (
        .din(new_Jinkela_wire_7601),
        .dout(new_Jinkela_wire_7602)
    );

    bfr new_Jinkela_buffer_5595 (
        .din(new_Jinkela_wire_7548),
        .dout(new_Jinkela_wire_7549)
    );

    bfr new_Jinkela_buffer_5624 (
        .din(new_Jinkela_wire_7580),
        .dout(new_Jinkela_wire_7581)
    );

    bfr new_Jinkela_buffer_5596 (
        .din(new_Jinkela_wire_7549),
        .dout(new_Jinkela_wire_7550)
    );

    bfr new_Jinkela_buffer_5597 (
        .din(new_Jinkela_wire_7550),
        .dout(new_Jinkela_wire_7551)
    );

    bfr new_Jinkela_buffer_5644 (
        .din(new_Jinkela_wire_7608),
        .dout(new_Jinkela_wire_7609)
    );

    bfr new_Jinkela_buffer_5625 (
        .din(new_Jinkela_wire_7581),
        .dout(new_Jinkela_wire_7582)
    );

    bfr new_Jinkela_buffer_5598 (
        .din(new_Jinkela_wire_7551),
        .dout(new_Jinkela_wire_7552)
    );

    bfr new_Jinkela_buffer_5599 (
        .din(new_Jinkela_wire_7552),
        .dout(new_Jinkela_wire_7553)
    );

    spl2 new_Jinkela_splitter_762 (
        .a(_0124_),
        .b(new_Jinkela_wire_7652),
        .c(new_Jinkela_wire_7653)
    );

    bfr new_Jinkela_buffer_5626 (
        .din(new_Jinkela_wire_7582),
        .dout(new_Jinkela_wire_7583)
    );

    bfr new_Jinkela_buffer_5600 (
        .din(new_Jinkela_wire_7553),
        .dout(new_Jinkela_wire_7554)
    );

    bfr new_Jinkela_buffer_5640 (
        .din(new_Jinkela_wire_7602),
        .dout(new_Jinkela_wire_7603)
    );

    bfr new_Jinkela_buffer_5601 (
        .din(new_Jinkela_wire_7554),
        .dout(new_Jinkela_wire_7555)
    );

    bfr new_Jinkela_buffer_5627 (
        .din(new_Jinkela_wire_7583),
        .dout(new_Jinkela_wire_7584)
    );

    bfr new_Jinkela_buffer_5602 (
        .din(new_Jinkela_wire_7555),
        .dout(new_Jinkela_wire_7556)
    );

    bfr new_Jinkela_buffer_5680 (
        .din(new_Jinkela_wire_7648),
        .dout(new_Jinkela_wire_7649)
    );

    bfr new_Jinkela_buffer_5603 (
        .din(new_Jinkela_wire_7556),
        .dout(new_Jinkela_wire_7557)
    );

    bfr new_Jinkela_buffer_5645 (
        .din(new_Jinkela_wire_7609),
        .dout(new_Jinkela_wire_7610)
    );

    bfr new_Jinkela_buffer_5628 (
        .din(new_Jinkela_wire_7584),
        .dout(new_Jinkela_wire_7585)
    );

    bfr new_Jinkela_buffer_5604 (
        .din(new_Jinkela_wire_7557),
        .dout(new_Jinkela_wire_7558)
    );

    bfr new_Jinkela_buffer_5641 (
        .din(new_Jinkela_wire_7603),
        .dout(new_Jinkela_wire_7604)
    );

    bfr new_Jinkela_buffer_5605 (
        .din(new_Jinkela_wire_7558),
        .dout(new_Jinkela_wire_7559)
    );

    bfr new_Jinkela_buffer_5629 (
        .din(new_Jinkela_wire_7585),
        .dout(new_Jinkela_wire_7586)
    );

    bfr new_Jinkela_buffer_5606 (
        .din(new_Jinkela_wire_7559),
        .dout(new_Jinkela_wire_7560)
    );

    bfr new_Jinkela_buffer_5607 (
        .din(new_Jinkela_wire_7560),
        .dout(new_Jinkela_wire_7561)
    );

    bfr new_Jinkela_buffer_5630 (
        .din(new_Jinkela_wire_7586),
        .dout(new_Jinkela_wire_7587)
    );

    bfr new_Jinkela_buffer_5608 (
        .din(new_Jinkela_wire_7561),
        .dout(new_Jinkela_wire_7562)
    );

    bfr new_Jinkela_buffer_5609 (
        .din(new_Jinkela_wire_7562),
        .dout(new_Jinkela_wire_7563)
    );

    bfr new_Jinkela_buffer_510 (
        .din(G111),
        .dout(new_Jinkela_wire_1026)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(new_Jinkela_wire_1016),
        .b(new_Jinkela_wire_1017),
        .c(new_Jinkela_wire_1018)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    spl2 new_Jinkela_splitter_176 (
        .a(new_Jinkela_wire_937),
        .b(new_Jinkela_wire_938),
        .c(new_Jinkela_wire_939)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    spl3L new_Jinkela_splitter_184 (
        .a(G176),
        .d(new_Jinkela_wire_1030),
        .b(new_Jinkela_wire_1031),
        .c(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_980),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

    spl2 new_Jinkela_splitter_203 (
        .a(G148),
        .b(new_Jinkela_wire_1101),
        .c(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_1022),
        .dout(new_Jinkela_wire_1023)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    spl3L new_Jinkela_splitter_183 (
        .a(new_Jinkela_wire_1026),
        .d(new_Jinkela_wire_1027),
        .b(new_Jinkela_wire_1028),
        .c(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    spl4L new_Jinkela_splitter_204 (
        .a(new_Jinkela_wire_1103),
        .d(new_Jinkela_wire_1104),
        .e(new_Jinkela_wire_1105),
        .b(new_Jinkela_wire_1106),
        .c(new_Jinkela_wire_1107)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_542 (
        .din(G63),
        .dout(new_Jinkela_wire_1127)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_534 (
        .din(G162),
        .dout(new_Jinkela_wire_1117)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(new_Jinkela_wire_1109),
        .b(new_Jinkela_wire_1110),
        .c(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_991),
        .dout(new_Jinkela_wire_992)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_529 (
        .din(G51),
        .dout(new_Jinkela_wire_1112)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_994),
        .dout(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_1101),
        .dout(new_Jinkela_wire_1102)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_1835 (
        .din(new_Jinkela_wire_2890),
        .dout(new_Jinkela_wire_2891)
    );

    spl2 new_Jinkela_splitter_623 (
        .a(_0596_),
        .b(new_Jinkela_wire_6015),
        .c(new_Jinkela_wire_6017)
    );

    bfr new_Jinkela_buffer_4394 (
        .din(_1013_),
        .dout(new_Jinkela_wire_6024)
    );

    bfr new_Jinkela_buffer_4299 (
        .din(new_Jinkela_wire_5922),
        .dout(new_Jinkela_wire_5923)
    );

    bfr new_Jinkela_buffer_1836 (
        .din(new_Jinkela_wire_2891),
        .dout(new_Jinkela_wire_2892)
    );

    bfr new_Jinkela_buffer_4312 (
        .din(new_Jinkela_wire_5935),
        .dout(new_Jinkela_wire_5936)
    );

    spl2 new_Jinkela_splitter_396 (
        .a(new_Jinkela_wire_2911),
        .b(new_Jinkela_wire_2912),
        .c(new_Jinkela_wire_2913)
    );

    bfr new_Jinkela_buffer_4300 (
        .din(new_Jinkela_wire_5923),
        .dout(new_Jinkela_wire_5924)
    );

    bfr new_Jinkela_buffer_1837 (
        .din(new_Jinkela_wire_2892),
        .dout(new_Jinkela_wire_2893)
    );

    bfr new_Jinkela_buffer_4327 (
        .din(new_Jinkela_wire_5950),
        .dout(new_Jinkela_wire_5951)
    );

    bfr new_Jinkela_buffer_1850 (
        .din(new_Jinkela_wire_2913),
        .dout(new_Jinkela_wire_2914)
    );

    bfr new_Jinkela_buffer_4301 (
        .din(new_Jinkela_wire_5924),
        .dout(new_Jinkela_wire_5925)
    );

    bfr new_Jinkela_buffer_1838 (
        .din(new_Jinkela_wire_2893),
        .dout(new_Jinkela_wire_2894)
    );

    bfr new_Jinkela_buffer_4313 (
        .din(new_Jinkela_wire_5936),
        .dout(new_Jinkela_wire_5937)
    );

    bfr new_Jinkela_buffer_1862 (
        .din(new_Jinkela_wire_2932),
        .dout(new_Jinkela_wire_2933)
    );

    bfr new_Jinkela_buffer_4302 (
        .din(new_Jinkela_wire_5925),
        .dout(new_Jinkela_wire_5926)
    );

    bfr new_Jinkela_buffer_1839 (
        .din(new_Jinkela_wire_2894),
        .dout(new_Jinkela_wire_2895)
    );

    bfr new_Jinkela_buffer_4352 (
        .din(new_Jinkela_wire_5975),
        .dout(new_Jinkela_wire_5976)
    );

    bfr new_Jinkela_buffer_1873 (
        .din(new_net_2379),
        .dout(new_Jinkela_wire_2946)
    );

    bfr new_Jinkela_buffer_4303 (
        .din(new_Jinkela_wire_5926),
        .dout(new_Jinkela_wire_5927)
    );

    bfr new_Jinkela_buffer_1870 (
        .din(new_Jinkela_wire_2940),
        .dout(new_Jinkela_wire_2941)
    );

    bfr new_Jinkela_buffer_1840 (
        .din(new_Jinkela_wire_2895),
        .dout(new_Jinkela_wire_2896)
    );

    bfr new_Jinkela_buffer_4314 (
        .din(new_Jinkela_wire_5937),
        .dout(new_Jinkela_wire_5938)
    );

    bfr new_Jinkela_buffer_1851 (
        .din(new_Jinkela_wire_2914),
        .dout(new_Jinkela_wire_2915)
    );

    bfr new_Jinkela_buffer_4304 (
        .din(new_Jinkela_wire_5927),
        .dout(new_Jinkela_wire_5928)
    );

    bfr new_Jinkela_buffer_1841 (
        .din(new_Jinkela_wire_2896),
        .dout(new_Jinkela_wire_2897)
    );

    bfr new_Jinkela_buffer_4328 (
        .din(new_Jinkela_wire_5951),
        .dout(new_Jinkela_wire_5952)
    );

    bfr new_Jinkela_buffer_1863 (
        .din(new_Jinkela_wire_2933),
        .dout(new_Jinkela_wire_2934)
    );

    bfr new_Jinkela_buffer_4315 (
        .din(new_Jinkela_wire_5938),
        .dout(new_Jinkela_wire_5939)
    );

    bfr new_Jinkela_buffer_1842 (
        .din(new_Jinkela_wire_2897),
        .dout(new_Jinkela_wire_2898)
    );

    spl3L new_Jinkela_splitter_626 (
        .a(_0964_),
        .d(new_Jinkela_wire_6043),
        .b(new_Jinkela_wire_6044),
        .c(new_Jinkela_wire_6045)
    );

    bfr new_Jinkela_buffer_4392 (
        .din(new_Jinkela_wire_6021),
        .dout(new_Jinkela_wire_6022)
    );

    bfr new_Jinkela_buffer_1852 (
        .din(new_Jinkela_wire_2915),
        .dout(new_Jinkela_wire_2916)
    );

    bfr new_Jinkela_buffer_4316 (
        .din(new_Jinkela_wire_5939),
        .dout(new_Jinkela_wire_5940)
    );

    bfr new_Jinkela_buffer_4329 (
        .din(new_Jinkela_wire_5952),
        .dout(new_Jinkela_wire_5953)
    );

    bfr new_Jinkela_buffer_1853 (
        .din(new_Jinkela_wire_2916),
        .dout(new_Jinkela_wire_2917)
    );

    bfr new_Jinkela_buffer_4317 (
        .din(new_Jinkela_wire_5940),
        .dout(new_Jinkela_wire_5941)
    );

    bfr new_Jinkela_buffer_1864 (
        .din(new_Jinkela_wire_2934),
        .dout(new_Jinkela_wire_2935)
    );

    bfr new_Jinkela_buffer_4353 (
        .din(new_Jinkela_wire_5976),
        .dout(new_Jinkela_wire_5977)
    );

    bfr new_Jinkela_buffer_1854 (
        .din(new_Jinkela_wire_2917),
        .dout(new_Jinkela_wire_2918)
    );

    bfr new_Jinkela_buffer_4318 (
        .din(new_Jinkela_wire_5941),
        .dout(new_Jinkela_wire_5942)
    );

    bfr new_Jinkela_buffer_1872 (
        .din(new_Jinkela_wire_2944),
        .dout(new_Jinkela_wire_2945)
    );

    bfr new_Jinkela_buffer_4330 (
        .din(new_Jinkela_wire_5953),
        .dout(new_Jinkela_wire_5954)
    );

    spl2 new_Jinkela_splitter_400 (
        .a(new_Jinkela_wire_2941),
        .b(new_Jinkela_wire_2942),
        .c(new_Jinkela_wire_2943)
    );

    bfr new_Jinkela_buffer_1855 (
        .din(new_Jinkela_wire_2918),
        .dout(new_Jinkela_wire_2919)
    );

    bfr new_Jinkela_buffer_4319 (
        .din(new_Jinkela_wire_5942),
        .dout(new_Jinkela_wire_5943)
    );

    bfr new_Jinkela_buffer_1865 (
        .din(new_Jinkela_wire_2935),
        .dout(new_Jinkela_wire_2936)
    );

    bfr new_Jinkela_buffer_4391 (
        .din(new_Jinkela_wire_6015),
        .dout(new_Jinkela_wire_6016)
    );

    spl4L new_Jinkela_splitter_624 (
        .a(new_Jinkela_wire_6017),
        .d(new_Jinkela_wire_6018),
        .e(new_Jinkela_wire_6019),
        .b(new_Jinkela_wire_6020),
        .c(new_Jinkela_wire_6021)
    );

    bfr new_Jinkela_buffer_1856 (
        .din(new_Jinkela_wire_2919),
        .dout(new_Jinkela_wire_2920)
    );

    bfr new_Jinkela_buffer_4320 (
        .din(new_Jinkela_wire_5943),
        .dout(new_Jinkela_wire_5944)
    );

    bfr new_Jinkela_buffer_4331 (
        .din(new_Jinkela_wire_5954),
        .dout(new_Jinkela_wire_5955)
    );

    bfr new_Jinkela_buffer_1913 (
        .din(new_net_2487),
        .dout(new_Jinkela_wire_2989)
    );

    bfr new_Jinkela_buffer_1857 (
        .din(new_Jinkela_wire_2920),
        .dout(new_Jinkela_wire_2921)
    );

    bfr new_Jinkela_buffer_4321 (
        .din(new_Jinkela_wire_5944),
        .dout(new_Jinkela_wire_5945)
    );

    bfr new_Jinkela_buffer_1866 (
        .din(new_Jinkela_wire_2936),
        .dout(new_Jinkela_wire_2937)
    );

    bfr new_Jinkela_buffer_4354 (
        .din(new_Jinkela_wire_5977),
        .dout(new_Jinkela_wire_5978)
    );

    bfr new_Jinkela_buffer_1858 (
        .din(new_Jinkela_wire_2921),
        .dout(new_Jinkela_wire_2922)
    );

    bfr new_Jinkela_buffer_4322 (
        .din(new_Jinkela_wire_5945),
        .dout(new_Jinkela_wire_5946)
    );

    bfr new_Jinkela_buffer_1874 (
        .din(new_Jinkela_wire_2946),
        .dout(new_Jinkela_wire_2947)
    );

    bfr new_Jinkela_buffer_4332 (
        .din(new_Jinkela_wire_5955),
        .dout(new_Jinkela_wire_5956)
    );

    bfr new_Jinkela_buffer_1859 (
        .din(new_Jinkela_wire_2922),
        .dout(new_Jinkela_wire_2923)
    );

    bfr new_Jinkela_buffer_4323 (
        .din(new_Jinkela_wire_5946),
        .dout(new_Jinkela_wire_5947)
    );

    bfr new_Jinkela_buffer_1867 (
        .din(new_Jinkela_wire_2937),
        .dout(new_Jinkela_wire_2938)
    );

    spl2 new_Jinkela_splitter_629 (
        .a(_0954_),
        .b(new_Jinkela_wire_6065),
        .c(new_Jinkela_wire_6066)
    );

    spl3L new_Jinkela_splitter_401 (
        .a(_0745_),
        .d(new_Jinkela_wire_2986),
        .b(new_Jinkela_wire_2987),
        .c(new_Jinkela_wire_2988)
    );

    bfr new_Jinkela_buffer_4324 (
        .din(new_Jinkela_wire_5947),
        .dout(new_Jinkela_wire_5948)
    );

    bfr new_Jinkela_buffer_1868 (
        .din(new_Jinkela_wire_2938),
        .dout(new_Jinkela_wire_2939)
    );

    bfr new_Jinkela_buffer_4333 (
        .din(new_Jinkela_wire_5956),
        .dout(new_Jinkela_wire_5957)
    );

    bfr new_Jinkela_buffer_4355 (
        .din(new_Jinkela_wire_5978),
        .dout(new_Jinkela_wire_5979)
    );

    spl4L new_Jinkela_splitter_402 (
        .a(_0757_),
        .d(new_Jinkela_wire_3028),
        .e(new_Jinkela_wire_3029),
        .b(new_Jinkela_wire_3030),
        .c(new_Jinkela_wire_3031)
    );

    bfr new_Jinkela_buffer_1875 (
        .din(new_Jinkela_wire_2947),
        .dout(new_Jinkela_wire_2948)
    );

    bfr new_Jinkela_buffer_4334 (
        .din(new_Jinkela_wire_5957),
        .dout(new_Jinkela_wire_5958)
    );

    bfr new_Jinkela_buffer_1952 (
        .din(_0563_),
        .dout(new_Jinkela_wire_3032)
    );

    bfr new_Jinkela_buffer_1876 (
        .din(new_Jinkela_wire_2948),
        .dout(new_Jinkela_wire_2949)
    );

    bfr new_Jinkela_buffer_4335 (
        .din(new_Jinkela_wire_5958),
        .dout(new_Jinkela_wire_5959)
    );

    bfr new_Jinkela_buffer_1914 (
        .din(new_Jinkela_wire_2989),
        .dout(new_Jinkela_wire_2990)
    );

    bfr new_Jinkela_buffer_4356 (
        .din(new_Jinkela_wire_5979),
        .dout(new_Jinkela_wire_5980)
    );

    bfr new_Jinkela_buffer_1877 (
        .din(new_Jinkela_wire_2949),
        .dout(new_Jinkela_wire_2950)
    );

    bfr new_Jinkela_buffer_4336 (
        .din(new_Jinkela_wire_5959),
        .dout(new_Jinkela_wire_5960)
    );

    bfr new_Jinkela_buffer_1878 (
        .din(new_Jinkela_wire_2950),
        .dout(new_Jinkela_wire_2951)
    );

    bfr new_Jinkela_buffer_4337 (
        .din(new_Jinkela_wire_5960),
        .dout(new_Jinkela_wire_5961)
    );

    bfr new_Jinkela_buffer_1915 (
        .din(new_Jinkela_wire_2990),
        .dout(new_Jinkela_wire_2991)
    );

    bfr new_Jinkela_buffer_4357 (
        .din(new_Jinkela_wire_5980),
        .dout(new_Jinkela_wire_5981)
    );

    bfr new_Jinkela_buffer_5646 (
        .din(new_Jinkela_wire_7610),
        .dout(new_Jinkela_wire_7611)
    );

    bfr new_Jinkela_buffer_4826 (
        .din(new_Jinkela_wire_6583),
        .dout(new_Jinkela_wire_6584)
    );

    bfr new_Jinkela_buffer_5631 (
        .din(new_Jinkela_wire_7587),
        .dout(new_Jinkela_wire_7588)
    );

    bfr new_Jinkela_buffer_5610 (
        .din(new_Jinkela_wire_7563),
        .dout(new_Jinkela_wire_7564)
    );

    bfr new_Jinkela_buffer_4868 (
        .din(new_Jinkela_wire_6629),
        .dout(new_Jinkela_wire_6630)
    );

    bfr new_Jinkela_buffer_4837 (
        .din(new_Jinkela_wire_6594),
        .dout(new_Jinkela_wire_6595)
    );

    bfr new_Jinkela_buffer_5611 (
        .din(new_Jinkela_wire_7564),
        .dout(new_Jinkela_wire_7565)
    );

    bfr new_Jinkela_buffer_4838 (
        .din(new_Jinkela_wire_6595),
        .dout(new_Jinkela_wire_6596)
    );

    bfr new_Jinkela_buffer_5682 (
        .din(new_Jinkela_wire_7656),
        .dout(new_Jinkela_wire_7657)
    );

    bfr new_Jinkela_buffer_5632 (
        .din(new_Jinkela_wire_7588),
        .dout(new_Jinkela_wire_7589)
    );

    spl3L new_Jinkela_splitter_754 (
        .a(new_Jinkela_wire_7565),
        .d(new_Jinkela_wire_7566),
        .b(new_Jinkela_wire_7567),
        .c(new_Jinkela_wire_7568)
    );

    bfr new_Jinkela_buffer_4869 (
        .din(new_Jinkela_wire_6630),
        .dout(new_Jinkela_wire_6631)
    );

    bfr new_Jinkela_buffer_4839 (
        .din(new_Jinkela_wire_6596),
        .dout(new_Jinkela_wire_6597)
    );

    bfr new_Jinkela_buffer_5647 (
        .din(new_Jinkela_wire_7611),
        .dout(new_Jinkela_wire_7612)
    );

    bfr new_Jinkela_buffer_4889 (
        .din(new_Jinkela_wire_6650),
        .dout(new_Jinkela_wire_6651)
    );

    bfr new_Jinkela_buffer_5633 (
        .din(new_Jinkela_wire_7589),
        .dout(new_Jinkela_wire_7590)
    );

    bfr new_Jinkela_buffer_4840 (
        .din(new_Jinkela_wire_6597),
        .dout(new_Jinkela_wire_6598)
    );

    spl2 new_Jinkela_splitter_761 (
        .a(new_Jinkela_wire_7649),
        .b(new_Jinkela_wire_7650),
        .c(new_Jinkela_wire_7651)
    );

    bfr new_Jinkela_buffer_4870 (
        .din(new_Jinkela_wire_6631),
        .dout(new_Jinkela_wire_6632)
    );

    bfr new_Jinkela_buffer_5634 (
        .din(new_Jinkela_wire_7590),
        .dout(new_Jinkela_wire_7591)
    );

    bfr new_Jinkela_buffer_4841 (
        .din(new_Jinkela_wire_6598),
        .dout(new_Jinkela_wire_6599)
    );

    bfr new_Jinkela_buffer_5648 (
        .din(new_Jinkela_wire_7612),
        .dout(new_Jinkela_wire_7613)
    );

    spl2 new_Jinkela_splitter_678 (
        .a(_0592_),
        .b(new_Jinkela_wire_6679),
        .c(new_Jinkela_wire_6685)
    );

    bfr new_Jinkela_buffer_5635 (
        .din(new_Jinkela_wire_7591),
        .dout(new_Jinkela_wire_7592)
    );

    bfr new_Jinkela_buffer_4842 (
        .din(new_Jinkela_wire_6599),
        .dout(new_Jinkela_wire_6600)
    );

    bfr new_Jinkela_buffer_4910 (
        .din(new_Jinkela_wire_6671),
        .dout(new_Jinkela_wire_6672)
    );

    bfr new_Jinkela_buffer_5798 (
        .din(_0009_),
        .dout(new_Jinkela_wire_7783)
    );

    bfr new_Jinkela_buffer_4871 (
        .din(new_Jinkela_wire_6632),
        .dout(new_Jinkela_wire_6633)
    );

    bfr new_Jinkela_buffer_5707 (
        .din(_0851_),
        .dout(new_Jinkela_wire_7682)
    );

    bfr new_Jinkela_buffer_4843 (
        .din(new_Jinkela_wire_6600),
        .dout(new_Jinkela_wire_6601)
    );

    bfr new_Jinkela_buffer_5649 (
        .din(new_Jinkela_wire_7613),
        .dout(new_Jinkela_wire_7614)
    );

    bfr new_Jinkela_buffer_4890 (
        .din(new_Jinkela_wire_6651),
        .dout(new_Jinkela_wire_6652)
    );

    bfr new_Jinkela_buffer_5681 (
        .din(_0928_),
        .dout(new_Jinkela_wire_7656)
    );

    bfr new_Jinkela_buffer_4844 (
        .din(new_Jinkela_wire_6601),
        .dout(new_Jinkela_wire_6602)
    );

    bfr new_Jinkela_buffer_5650 (
        .din(new_Jinkela_wire_7614),
        .dout(new_Jinkela_wire_7615)
    );

    bfr new_Jinkela_buffer_4872 (
        .din(new_Jinkela_wire_6633),
        .dout(new_Jinkela_wire_6634)
    );

    bfr new_Jinkela_buffer_4845 (
        .din(new_Jinkela_wire_6602),
        .dout(new_Jinkela_wire_6603)
    );

    bfr new_Jinkela_buffer_5651 (
        .din(new_Jinkela_wire_7615),
        .dout(new_Jinkela_wire_7616)
    );

    bfr new_Jinkela_buffer_5733 (
        .din(new_Jinkela_wire_7715),
        .dout(new_Jinkela_wire_7716)
    );

    bfr new_Jinkela_buffer_5683 (
        .din(new_Jinkela_wire_7657),
        .dout(new_Jinkela_wire_7658)
    );

    bfr new_Jinkela_buffer_4846 (
        .din(new_Jinkela_wire_6603),
        .dout(new_Jinkela_wire_6604)
    );

    bfr new_Jinkela_buffer_5652 (
        .din(new_Jinkela_wire_7616),
        .dout(new_Jinkela_wire_7617)
    );

    bfr new_Jinkela_buffer_4873 (
        .din(new_Jinkela_wire_6634),
        .dout(new_Jinkela_wire_6635)
    );

    bfr new_Jinkela_buffer_4847 (
        .din(new_Jinkela_wire_6604),
        .dout(new_Jinkela_wire_6605)
    );

    bfr new_Jinkela_buffer_5653 (
        .din(new_Jinkela_wire_7617),
        .dout(new_Jinkela_wire_7618)
    );

    bfr new_Jinkela_buffer_5708 (
        .din(new_Jinkela_wire_7682),
        .dout(new_Jinkela_wire_7683)
    );

    bfr new_Jinkela_buffer_4891 (
        .din(new_Jinkela_wire_6652),
        .dout(new_Jinkela_wire_6653)
    );

    bfr new_Jinkela_buffer_5684 (
        .din(new_Jinkela_wire_7658),
        .dout(new_Jinkela_wire_7659)
    );

    bfr new_Jinkela_buffer_4848 (
        .din(new_Jinkela_wire_6605),
        .dout(new_Jinkela_wire_6606)
    );

    bfr new_Jinkela_buffer_5654 (
        .din(new_Jinkela_wire_7618),
        .dout(new_Jinkela_wire_7619)
    );

    bfr new_Jinkela_buffer_4874 (
        .din(new_Jinkela_wire_6635),
        .dout(new_Jinkela_wire_6636)
    );

    bfr new_Jinkela_buffer_4849 (
        .din(new_Jinkela_wire_6606),
        .dout(new_Jinkela_wire_6607)
    );

    bfr new_Jinkela_buffer_5655 (
        .din(new_Jinkela_wire_7619),
        .dout(new_Jinkela_wire_7620)
    );

    bfr new_Jinkela_buffer_4913 (
        .din(_0742_),
        .dout(new_Jinkela_wire_6706)
    );

    bfr new_Jinkela_buffer_5685 (
        .din(new_Jinkela_wire_7659),
        .dout(new_Jinkela_wire_7660)
    );

    bfr new_Jinkela_buffer_4850 (
        .din(new_Jinkela_wire_6607),
        .dout(new_Jinkela_wire_6608)
    );

    bfr new_Jinkela_buffer_5656 (
        .din(new_Jinkela_wire_7620),
        .dout(new_Jinkela_wire_7621)
    );

    bfr new_Jinkela_buffer_4911 (
        .din(new_Jinkela_wire_6672),
        .dout(new_Jinkela_wire_6673)
    );

    bfr new_Jinkela_buffer_4875 (
        .din(new_Jinkela_wire_6636),
        .dout(new_Jinkela_wire_6637)
    );

    spl2 new_Jinkela_splitter_768 (
        .a(new_net_13),
        .b(new_Jinkela_wire_7741),
        .c(new_Jinkela_wire_7742)
    );

    bfr new_Jinkela_buffer_4851 (
        .din(new_Jinkela_wire_6608),
        .dout(new_Jinkela_wire_6609)
    );

    bfr new_Jinkela_buffer_5657 (
        .din(new_Jinkela_wire_7621),
        .dout(new_Jinkela_wire_7622)
    );

    bfr new_Jinkela_buffer_5709 (
        .din(new_Jinkela_wire_7683),
        .dout(new_Jinkela_wire_7684)
    );

    bfr new_Jinkela_buffer_4892 (
        .din(new_Jinkela_wire_6653),
        .dout(new_Jinkela_wire_6654)
    );

    bfr new_Jinkela_buffer_5686 (
        .din(new_Jinkela_wire_7660),
        .dout(new_Jinkela_wire_7661)
    );

    bfr new_Jinkela_buffer_4852 (
        .din(new_Jinkela_wire_6609),
        .dout(new_Jinkela_wire_6610)
    );

    bfr new_Jinkela_buffer_5658 (
        .din(new_Jinkela_wire_7622),
        .dout(new_Jinkela_wire_7623)
    );

    bfr new_Jinkela_buffer_4876 (
        .din(new_Jinkela_wire_6637),
        .dout(new_Jinkela_wire_6638)
    );

    bfr new_Jinkela_buffer_4853 (
        .din(new_Jinkela_wire_6610),
        .dout(new_Jinkela_wire_6611)
    );

    bfr new_Jinkela_buffer_5659 (
        .din(new_Jinkela_wire_7623),
        .dout(new_Jinkela_wire_7624)
    );

    bfr new_Jinkela_buffer_5687 (
        .din(new_Jinkela_wire_7661),
        .dout(new_Jinkela_wire_7662)
    );

    bfr new_Jinkela_buffer_4854 (
        .din(new_Jinkela_wire_6611),
        .dout(new_Jinkela_wire_6612)
    );

    bfr new_Jinkela_buffer_5660 (
        .din(new_Jinkela_wire_7624),
        .dout(new_Jinkela_wire_7625)
    );

    bfr new_Jinkela_buffer_4914 (
        .din(_0245_),
        .dout(new_Jinkela_wire_6709)
    );

    bfr new_Jinkela_buffer_4877 (
        .din(new_Jinkela_wire_6638),
        .dout(new_Jinkela_wire_6639)
    );

    spl2 new_Jinkela_splitter_767 (
        .a(_0914_),
        .b(new_Jinkela_wire_7713),
        .c(new_Jinkela_wire_7714)
    );

    bfr new_Jinkela_buffer_4855 (
        .din(new_Jinkela_wire_6612),
        .dout(new_Jinkela_wire_6613)
    );

    bfr new_Jinkela_buffer_5661 (
        .din(new_Jinkela_wire_7625),
        .dout(new_Jinkela_wire_7626)
    );

    bfr new_Jinkela_buffer_4893 (
        .din(new_Jinkela_wire_6654),
        .dout(new_Jinkela_wire_6655)
    );

    bfr new_Jinkela_buffer_5688 (
        .din(new_Jinkela_wire_7662),
        .dout(new_Jinkela_wire_7663)
    );

    bfr new_Jinkela_buffer_4856 (
        .din(new_Jinkela_wire_6613),
        .dout(new_Jinkela_wire_6614)
    );

    bfr new_Jinkela_buffer_5662 (
        .din(new_Jinkela_wire_7626),
        .dout(new_Jinkela_wire_7627)
    );

    bfr new_Jinkela_buffer_4878 (
        .din(new_Jinkela_wire_6639),
        .dout(new_Jinkela_wire_6640)
    );

    bfr new_Jinkela_buffer_5732 (
        .din(new_net_2485),
        .dout(new_Jinkela_wire_7715)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    spl3L new_Jinkela_splitter_186 (
        .a(new_Jinkela_wire_1039),
        .d(new_Jinkela_wire_1040),
        .b(new_Jinkela_wire_1041),
        .c(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(G156),
        .b(new_Jinkela_wire_1133),
        .c(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(G149),
        .b(new_Jinkela_wire_1128),
        .c(new_Jinkela_wire_1129)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    spl4L new_Jinkela_splitter_188 (
        .a(new_Jinkela_wire_1044),
        .d(new_Jinkela_wire_1045),
        .e(new_Jinkela_wire_1046),
        .b(new_Jinkela_wire_1051),
        .c(new_Jinkela_wire_1056)
    );

    spl4L new_Jinkela_splitter_185 (
        .a(new_Jinkela_wire_1035),
        .d(new_Jinkela_wire_1036),
        .e(new_Jinkela_wire_1037),
        .b(new_Jinkela_wire_1038),
        .c(new_Jinkela_wire_1039)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_1129),
        .dout(new_Jinkela_wire_1130)
    );

    spl4L new_Jinkela_splitter_189 (
        .a(new_Jinkela_wire_1046),
        .d(new_Jinkela_wire_1047),
        .e(new_Jinkela_wire_1048),
        .b(new_Jinkela_wire_1049),
        .c(new_Jinkela_wire_1050)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_1060),
        .dout(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    spl4L new_Jinkela_splitter_191 (
        .a(new_Jinkela_wire_1056),
        .d(new_Jinkela_wire_1057),
        .e(new_Jinkela_wire_1058),
        .b(new_Jinkela_wire_1059),
        .c(new_Jinkela_wire_1060)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    spl2 new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_1041),
        .b(new_Jinkela_wire_1042),
        .c(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_1011),
        .dout(new_Jinkela_wire_1012)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    spl4L new_Jinkela_splitter_190 (
        .a(new_Jinkela_wire_1051),
        .d(new_Jinkela_wire_1052),
        .e(new_Jinkela_wire_1053),
        .b(new_Jinkela_wire_1054),
        .c(new_Jinkela_wire_1055)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(G155),
        .b(new_Jinkela_wire_1135),
        .c(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(new_Jinkela_wire_1061),
        .b(new_Jinkela_wire_1062),
        .c(new_Jinkela_wire_1063)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(G144),
        .b(new_Jinkela_wire_1137),
        .c(new_Jinkela_wire_1138)
    );

    and_bi _2075_ (
        .a(new_Jinkela_wire_827),
        .b(new_Jinkela_wire_168),
        .c(_0113_)
    );

    and_ii _2076_ (
        .a(_0113_),
        .b(_0112_),
        .c(_0114_)
    );

    and_ii _2077_ (
        .a(new_Jinkela_wire_2532),
        .b(new_Jinkela_wire_7189),
        .c(_0115_)
    );

    and_bb _2078_ (
        .a(new_Jinkela_wire_2533),
        .b(new_Jinkela_wire_7190),
        .c(_0116_)
    );

    and_ii _2079_ (
        .a(_0116_),
        .b(_0115_),
        .c(_0117_)
    );

    inv _2080_ (
        .din(_0117_),
        .dout(_0118_)
    );

    and_bi _2081_ (
        .a(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_77),
        .c(_0119_)
    );

    and_bi _2082_ (
        .a(new_Jinkela_wire_76),
        .b(new_Jinkela_wire_1361),
        .c(_0120_)
    );

    or_bb _2083_ (
        .a(_0120_),
        .b(_0119_),
        .c(_0121_)
    );

    and_bi _2084_ (
        .a(new_Jinkela_wire_107),
        .b(new_Jinkela_wire_5392),
        .c(_0122_)
    );

    and_bi _2085_ (
        .a(new_Jinkela_wire_5393),
        .b(new_Jinkela_wire_106),
        .c(_0123_)
    );

    and_ii _2086_ (
        .a(_0123_),
        .b(_0122_),
        .c(_0124_)
    );

    and_bi _2087_ (
        .a(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_281),
        .c(_0125_)
    );

    and_bi _2088_ (
        .a(new_Jinkela_wire_283),
        .b(new_Jinkela_wire_424),
        .c(_0126_)
    );

    and_ii _2089_ (
        .a(_0126_),
        .b(_0125_),
        .c(_0127_)
    );

    and_bi _2090_ (
        .a(new_Jinkela_wire_6674),
        .b(new_Jinkela_wire_7652),
        .c(_0128_)
    );

    and_bi _2091_ (
        .a(new_Jinkela_wire_7653),
        .b(new_Jinkela_wire_6675),
        .c(_0129_)
    );

    and_ii _2092_ (
        .a(_0129_),
        .b(_0128_),
        .c(_0130_)
    );

    and_bi _2093_ (
        .a(new_Jinkela_wire_7824),
        .b(new_Jinkela_wire_5552),
        .c(_0131_)
    );

    and_bi _2094_ (
        .a(new_Jinkela_wire_5553),
        .b(new_Jinkela_wire_7825),
        .c(_0132_)
    );

    or_bb _2095_ (
        .a(_0132_),
        .b(_0131_),
        .c(new_net_15)
    );

    and_ii _2096_ (
        .a(new_Jinkela_wire_256),
        .b(new_Jinkela_wire_1337),
        .c(_0133_)
    );

    and_bb _2097_ (
        .a(new_Jinkela_wire_262),
        .b(new_Jinkela_wire_1331),
        .c(_0134_)
    );

    and_ii _2098_ (
        .a(_0134_),
        .b(_0133_),
        .c(_0135_)
    );

    and_bi _2099_ (
        .a(new_Jinkela_wire_555),
        .b(new_Jinkela_wire_847),
        .c(_0136_)
    );

    and_bi _2100_ (
        .a(new_Jinkela_wire_858),
        .b(new_Jinkela_wire_553),
        .c(_0137_)
    );

    and_ii _2101_ (
        .a(_0137_),
        .b(_0136_),
        .c(_0138_)
    );

    and_ii _2102_ (
        .a(new_Jinkela_wire_1972),
        .b(new_Jinkela_wire_7654),
        .c(_0139_)
    );

    and_bb _2103_ (
        .a(new_Jinkela_wire_1973),
        .b(new_Jinkela_wire_7655),
        .c(_0140_)
    );

    and_ii _2104_ (
        .a(_0140_),
        .b(_0139_),
        .c(_0141_)
    );

    and_ii _2105_ (
        .a(new_Jinkela_wire_445),
        .b(new_Jinkela_wire_205),
        .c(_0142_)
    );

    and_bb _2106_ (
        .a(new_Jinkela_wire_446),
        .b(new_Jinkela_wire_195),
        .c(_0143_)
    );

    and_ii _2107_ (
        .a(_0143_),
        .b(_0142_),
        .c(_0144_)
    );

    and_bi _2108_ (
        .a(new_Jinkela_wire_741),
        .b(new_Jinkela_wire_1028),
        .c(_0145_)
    );

    and_bi _2109_ (
        .a(new_Jinkela_wire_1027),
        .b(new_Jinkela_wire_743),
        .c(_0146_)
    );

    and_ii _2110_ (
        .a(_0146_),
        .b(_0145_),
        .c(_0147_)
    );

    and_bi _2111_ (
        .a(new_Jinkela_wire_6230),
        .b(new_Jinkela_wire_2313),
        .c(_0148_)
    );

    and_bi _2112_ (
        .a(new_Jinkela_wire_2314),
        .b(new_Jinkela_wire_6231),
        .c(_0149_)
    );

    or_bb _2113_ (
        .a(_0149_),
        .b(_0148_),
        .c(_0150_)
    );

    and_bi _2114_ (
        .a(new_Jinkela_wire_155),
        .b(new_Jinkela_wire_1321),
        .c(_0151_)
    );

    and_bi _2115_ (
        .a(new_Jinkela_wire_1320),
        .b(new_Jinkela_wire_160),
        .c(_0152_)
    );

    or_bb _2116_ (
        .a(_0152_),
        .b(_0151_),
        .c(_0153_)
    );

    and_bi _1361_ (
        .a(new_Jinkela_wire_1432),
        .b(new_Jinkela_wire_881),
        .c(_0665_)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1774),
        .dout(new_Jinkela_wire_1775)
    );

    bfr new_Jinkela_buffer_4249 (
        .din(new_Jinkela_wire_5852),
        .dout(new_Jinkela_wire_5853)
    );

    or_bb _1362_ (
        .a(_0665_),
        .b(_0664_),
        .c(_0666_)
    );

    bfr new_Jinkela_buffer_971 (
        .din(_0225_),
        .dout(new_Jinkela_wire_1860)
    );

    bfr new_Jinkela_buffer_4274 (
        .din(new_Jinkela_wire_5885),
        .dout(new_Jinkela_wire_5886)
    );

    and_bi _1363_ (
        .a(new_Jinkela_wire_7890),
        .b(new_Jinkela_wire_3589),
        .c(_0667_)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1775),
        .dout(new_Jinkela_wire_1776)
    );

    bfr new_Jinkela_buffer_4250 (
        .din(new_Jinkela_wire_5853),
        .dout(new_Jinkela_wire_5854)
    );

    and_bi _1364_ (
        .a(new_Jinkela_wire_3590),
        .b(new_Jinkela_wire_7889),
        .c(_0668_)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1797),
        .dout(new_Jinkela_wire_1798)
    );

    bfr new_Jinkela_buffer_4271 (
        .din(new_Jinkela_wire_5876),
        .dout(new_Jinkela_wire_5877)
    );

    and_ii _1365_ (
        .a(new_Jinkela_wire_4712),
        .b(new_Jinkela_wire_3416),
        .c(_0669_)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1776),
        .dout(new_Jinkela_wire_1777)
    );

    bfr new_Jinkela_buffer_4251 (
        .din(new_Jinkela_wire_5854),
        .dout(new_Jinkela_wire_5855)
    );

    inv _1366_ (
        .din(new_Jinkela_wire_5273),
        .dout(_0670_)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    spl2 new_Jinkela_splitter_620 (
        .a(_1084_),
        .b(new_Jinkela_wire_5906),
        .c(new_Jinkela_wire_5907)
    );

    or_bi _1367_ (
        .a(new_Jinkela_wire_5690),
        .b(new_Jinkela_wire_2408),
        .c(_0671_)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_1777),
        .dout(new_Jinkela_wire_1778)
    );

    bfr new_Jinkela_buffer_4252 (
        .din(new_Jinkela_wire_5855),
        .dout(new_Jinkela_wire_5856)
    );

    and_bi _1368_ (
        .a(new_Jinkela_wire_2813),
        .b(new_Jinkela_wire_6470),
        .c(_0672_)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_1798),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_4275 (
        .din(new_Jinkela_wire_5886),
        .dout(new_Jinkela_wire_5887)
    );

    inv _1369_ (
        .din(new_Jinkela_wire_7647),
        .dout(_0673_)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1778),
        .dout(new_Jinkela_wire_1779)
    );

    bfr new_Jinkela_buffer_4253 (
        .din(new_Jinkela_wire_5856),
        .dout(new_Jinkela_wire_5857)
    );

    and_bi _1370_ (
        .a(new_Jinkela_wire_6357),
        .b(new_Jinkela_wire_4714),
        .c(_0674_)
    );

    spl3L new_Jinkela_splitter_330 (
        .a(_0969_),
        .d(new_Jinkela_wire_1889),
        .b(new_Jinkela_wire_1890),
        .c(new_Jinkela_wire_1891)
    );

    spl3L new_Jinkela_splitter_324 (
        .a(new_Jinkela_wire_1854),
        .d(new_Jinkela_wire_1855),
        .b(new_Jinkela_wire_1856),
        .c(new_Jinkela_wire_1857)
    );

    or_bb _1371_ (
        .a(_0674_),
        .b(new_Jinkela_wire_3419),
        .c(_0675_)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1779),
        .dout(new_Jinkela_wire_1780)
    );

    bfr new_Jinkela_buffer_4276 (
        .din(new_Jinkela_wire_5887),
        .dout(new_Jinkela_wire_5888)
    );

    or_bi _1372_ (
        .a(new_Jinkela_wire_6951),
        .b(new_Jinkela_wire_5818),
        .c(_0676_)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    spl2 new_Jinkela_splitter_621 (
        .a(new_net_5),
        .b(new_Jinkela_wire_5908),
        .c(new_Jinkela_wire_5910)
    );

    bfr new_Jinkela_buffer_4291 (
        .din(new_Jinkela_wire_5914),
        .dout(new_Jinkela_wire_5915)
    );

    and_bi _1373_ (
        .a(_0676_),
        .b(new_Jinkela_wire_3827),
        .c(_0677_)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1780),
        .dout(new_Jinkela_wire_1781)
    );

    bfr new_Jinkela_buffer_4277 (
        .din(new_Jinkela_wire_5888),
        .dout(new_Jinkela_wire_5889)
    );

    or_bb _1374_ (
        .a(new_Jinkela_wire_1966),
        .b(new_Jinkela_wire_4569),
        .c(_0678_)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1826),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_4305 (
        .din(_0765_),
        .dout(new_Jinkela_wire_5929)
    );

    or_bb _1375_ (
        .a(new_Jinkela_wire_1324),
        .b(new_Jinkela_wire_888),
        .c(_0679_)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1781),
        .dout(new_Jinkela_wire_1782)
    );

    bfr new_Jinkela_buffer_4278 (
        .din(new_Jinkela_wire_5889),
        .dout(new_Jinkela_wire_5890)
    );

    and_bi _1376_ (
        .a(new_Jinkela_wire_892),
        .b(new_Jinkela_wire_104),
        .c(_0680_)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    or_bi _1377_ (
        .a(_0680_),
        .b(new_Jinkela_wire_1849),
        .c(_0681_)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1782),
        .dout(new_Jinkela_wire_1783)
    );

    bfr new_Jinkela_buffer_4279 (
        .din(new_Jinkela_wire_5890),
        .dout(new_Jinkela_wire_5891)
    );

    and_bi _1378_ (
        .a(new_Jinkela_wire_1233),
        .b(new_Jinkela_wire_7084),
        .c(_0682_)
    );

    spl4L new_Jinkela_splitter_622 (
        .a(new_Jinkela_wire_5910),
        .d(new_Jinkela_wire_5911),
        .e(new_Jinkela_wire_5912),
        .b(new_Jinkela_wire_5913),
        .c(new_Jinkela_wire_5914)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1853),
        .dout(new_Jinkela_wire_1854)
    );

    and_bi _1379_ (
        .a(new_Jinkela_wire_7083),
        .b(new_Jinkela_wire_1234),
        .c(_0683_)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    bfr new_Jinkela_buffer_4280 (
        .din(new_Jinkela_wire_5891),
        .dout(new_Jinkela_wire_5892)
    );

    or_bb _1380_ (
        .a(new_Jinkela_wire_5404),
        .b(new_Jinkela_wire_6921),
        .c(_0684_)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    bfr new_Jinkela_buffer_4308 (
        .din(_0524_),
        .dout(new_Jinkela_wire_5932)
    );

    bfr new_Jinkela_buffer_4290 (
        .din(new_Jinkela_wire_5908),
        .dout(new_Jinkela_wire_5909)
    );

    and_bi _1381_ (
        .a(new_Jinkela_wire_4357),
        .b(new_Jinkela_wire_1953),
        .c(_0685_)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    bfr new_Jinkela_buffer_4281 (
        .din(new_Jinkela_wire_5892),
        .dout(new_Jinkela_wire_5893)
    );

    and_bi _1382_ (
        .a(new_Jinkela_wire_1952),
        .b(new_Jinkela_wire_4358),
        .c(_0686_)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    bfr new_Jinkela_buffer_4306 (
        .din(new_Jinkela_wire_5929),
        .dout(new_Jinkela_wire_5930)
    );

    or_bb _1383_ (
        .a(_0686_),
        .b(_0685_),
        .c(_0687_)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1785),
        .dout(new_Jinkela_wire_1786)
    );

    bfr new_Jinkela_buffer_4282 (
        .din(new_Jinkela_wire_5893),
        .dout(new_Jinkela_wire_5894)
    );

    or_bb _1384_ (
        .a(new_Jinkela_wire_6755),
        .b(new_Jinkela_wire_1082),
        .c(_0688_)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_1802),
        .dout(new_Jinkela_wire_1803)
    );

    bfr new_Jinkela_buffer_4325 (
        .din(new_net_2411),
        .dout(new_Jinkela_wire_5949)
    );

    inv _1385_ (
        .din(new_Jinkela_wire_1225),
        .dout(_0689_)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1786),
        .dout(new_Jinkela_wire_1787)
    );

    bfr new_Jinkela_buffer_4283 (
        .din(new_Jinkela_wire_5894),
        .dout(new_Jinkela_wire_5895)
    );

    or_bb _1386_ (
        .a(new_Jinkela_wire_100),
        .b(new_Jinkela_wire_325),
        .c(_0690_)
    );

    bfr new_Jinkela_buffer_4292 (
        .din(new_Jinkela_wire_5915),
        .dout(new_Jinkela_wire_5916)
    );

    bfr new_Jinkela_buffer_986 (
        .din(_0897_),
        .dout(new_Jinkela_wire_1879)
    );

    and_bi _1387_ (
        .a(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_222),
        .c(_0691_)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1803),
        .dout(new_Jinkela_wire_1804)
    );

    bfr new_Jinkela_buffer_4284 (
        .din(new_Jinkela_wire_5895),
        .dout(new_Jinkela_wire_5896)
    );

    and_bi _1388_ (
        .a(_0690_),
        .b(_0691_),
        .c(_0692_)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    bfr new_Jinkela_buffer_4307 (
        .din(new_Jinkela_wire_5930),
        .dout(new_Jinkela_wire_5931)
    );

    or_bb _1389_ (
        .a(_0692_),
        .b(new_Jinkela_wire_7187),
        .c(_0693_)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_1804),
        .dout(new_Jinkela_wire_1805)
    );

    bfr new_Jinkela_buffer_4285 (
        .din(new_Jinkela_wire_5896),
        .dout(new_Jinkela_wire_5897)
    );

    or_ii _1390_ (
        .a(new_Jinkela_wire_93),
        .b(new_Jinkela_wire_1588),
        .c(_0694_)
    );

    spl2 new_Jinkela_splitter_326 (
        .a(_0871_),
        .b(new_Jinkela_wire_1861),
        .c(new_Jinkela_wire_1862)
    );

    bfr new_Jinkela_buffer_4293 (
        .din(new_Jinkela_wire_5916),
        .dout(new_Jinkela_wire_5917)
    );

    and_bi _1391_ (
        .a(new_Jinkela_wire_1288),
        .b(new_Jinkela_wire_95),
        .c(_0695_)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1805),
        .dout(new_Jinkela_wire_1806)
    );

    bfr new_Jinkela_buffer_4286 (
        .din(new_Jinkela_wire_5897),
        .dout(new_Jinkela_wire_5898)
    );

    and_bi _1392_ (
        .a(_0694_),
        .b(_0695_),
        .c(_0696_)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    bfr new_Jinkela_buffer_4309 (
        .din(new_Jinkela_wire_5932),
        .dout(new_Jinkela_wire_5933)
    );

    and_bi _1393_ (
        .a(new_Jinkela_wire_7188),
        .b(_0696_),
        .c(_0697_)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1806),
        .dout(new_Jinkela_wire_1807)
    );

    bfr new_Jinkela_buffer_4287 (
        .din(new_Jinkela_wire_5898),
        .dout(new_Jinkela_wire_5899)
    );

    and_bi _1394_ (
        .a(_0693_),
        .b(_0697_),
        .c(_0698_)
    );

    bfr new_Jinkela_buffer_4294 (
        .din(new_Jinkela_wire_5917),
        .dout(new_Jinkela_wire_5918)
    );

    spl2 new_Jinkela_splitter_331 (
        .a(_0962_),
        .b(new_Jinkela_wire_1904),
        .c(new_Jinkela_wire_1905)
    );

    and_bi _1395_ (
        .a(new_Jinkela_wire_1053),
        .b(new_Jinkela_wire_4464),
        .c(_0699_)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    bfr new_Jinkela_buffer_4351 (
        .din(new_net_2429),
        .dout(new_Jinkela_wire_5975)
    );

    or_bb _1396_ (
        .a(_0699_),
        .b(new_Jinkela_wire_4831),
        .c(_0700_)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1830),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_4295 (
        .din(new_Jinkela_wire_5918),
        .dout(new_Jinkela_wire_5919)
    );

    and_bi _1397_ (
        .a(_0688_),
        .b(new_Jinkela_wire_4899),
        .c(_0701_)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    bfr new_Jinkela_buffer_4310 (
        .din(new_Jinkela_wire_5933),
        .dout(new_Jinkela_wire_5934)
    );

    and_ii _1398_ (
        .a(_0701_),
        .b(new_Jinkela_wire_4376),
        .c(new_net_6)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1862),
        .dout(new_Jinkela_wire_1863)
    );

    bfr new_Jinkela_buffer_4296 (
        .din(new_Jinkela_wire_5919),
        .dout(new_Jinkela_wire_5920)
    );

    and_bi _1399_ (
        .a(new_Jinkela_wire_1571),
        .b(new_Jinkela_wire_6700),
        .c(_0702_)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    bfr new_Jinkela_buffer_4326 (
        .din(new_Jinkela_wire_5949),
        .dout(new_Jinkela_wire_5950)
    );

    and_bi _1400_ (
        .a(new_Jinkela_wire_6471),
        .b(new_Jinkela_wire_6955),
        .c(_0703_)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    bfr new_Jinkela_buffer_4297 (
        .din(new_Jinkela_wire_5920),
        .dout(new_Jinkela_wire_5921)
    );

    or_bb _1401_ (
        .a(new_Jinkela_wire_7237),
        .b(new_Jinkela_wire_2817),
        .c(_0704_)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1810),
        .dout(new_Jinkela_wire_1811)
    );

    bfr new_Jinkela_buffer_4311 (
        .din(new_Jinkela_wire_5934),
        .dout(new_Jinkela_wire_5935)
    );

    and_bb _1402_ (
        .a(new_Jinkela_wire_7238),
        .b(new_Jinkela_wire_2816),
        .c(_0705_)
    );

    bfr new_Jinkela_buffer_4298 (
        .din(new_Jinkela_wire_5921),
        .dout(new_Jinkela_wire_5922)
    );

    bfr new_Jinkela_buffer_4857 (
        .din(new_Jinkela_wire_6614),
        .dout(new_Jinkela_wire_6615)
    );

    bfr new_Jinkela_buffer_5663 (
        .din(new_Jinkela_wire_7627),
        .dout(new_Jinkela_wire_7628)
    );

    spl2 new_Jinkela_splitter_685 (
        .a(new_Jinkela_wire_6706),
        .b(new_Jinkela_wire_6707),
        .c(new_Jinkela_wire_6708)
    );

    bfr new_Jinkela_buffer_5689 (
        .din(new_Jinkela_wire_7663),
        .dout(new_Jinkela_wire_7664)
    );

    bfr new_Jinkela_buffer_4858 (
        .din(new_Jinkela_wire_6615),
        .dout(new_Jinkela_wire_6616)
    );

    bfr new_Jinkela_buffer_5664 (
        .din(new_Jinkela_wire_7628),
        .dout(new_Jinkela_wire_7629)
    );

    spl2 new_Jinkela_splitter_676 (
        .a(new_Jinkela_wire_6673),
        .b(new_Jinkela_wire_6674),
        .c(new_Jinkela_wire_6675)
    );

    bfr new_Jinkela_buffer_4879 (
        .din(new_Jinkela_wire_6640),
        .dout(new_Jinkela_wire_6641)
    );

    bfr new_Jinkela_buffer_5710 (
        .din(new_Jinkela_wire_7684),
        .dout(new_Jinkela_wire_7685)
    );

    bfr new_Jinkela_buffer_4859 (
        .din(new_Jinkela_wire_6616),
        .dout(new_Jinkela_wire_6617)
    );

    bfr new_Jinkela_buffer_5665 (
        .din(new_Jinkela_wire_7629),
        .dout(new_Jinkela_wire_7630)
    );

    bfr new_Jinkela_buffer_5758 (
        .din(new_Jinkela_wire_7742),
        .dout(new_Jinkela_wire_7743)
    );

    bfr new_Jinkela_buffer_4894 (
        .din(new_Jinkela_wire_6655),
        .dout(new_Jinkela_wire_6656)
    );

    bfr new_Jinkela_buffer_5690 (
        .din(new_Jinkela_wire_7664),
        .dout(new_Jinkela_wire_7665)
    );

    bfr new_Jinkela_buffer_4860 (
        .din(new_Jinkela_wire_6617),
        .dout(new_Jinkela_wire_6618)
    );

    bfr new_Jinkela_buffer_5666 (
        .din(new_Jinkela_wire_7630),
        .dout(new_Jinkela_wire_7631)
    );

    bfr new_Jinkela_buffer_4880 (
        .din(new_Jinkela_wire_6641),
        .dout(new_Jinkela_wire_6642)
    );

    bfr new_Jinkela_buffer_5711 (
        .din(new_Jinkela_wire_7685),
        .dout(new_Jinkela_wire_7686)
    );

    bfr new_Jinkela_buffer_4861 (
        .din(new_Jinkela_wire_6618),
        .dout(new_Jinkela_wire_6619)
    );

    bfr new_Jinkela_buffer_5667 (
        .din(new_Jinkela_wire_7631),
        .dout(new_Jinkela_wire_7632)
    );

    bfr new_Jinkela_buffer_5691 (
        .din(new_Jinkela_wire_7665),
        .dout(new_Jinkela_wire_7666)
    );

    spl2 new_Jinkela_splitter_674 (
        .a(new_Jinkela_wire_6619),
        .b(new_Jinkela_wire_6620),
        .c(new_Jinkela_wire_6621)
    );

    bfr new_Jinkela_buffer_5668 (
        .din(new_Jinkela_wire_7632),
        .dout(new_Jinkela_wire_7633)
    );

    bfr new_Jinkela_buffer_4895 (
        .din(new_Jinkela_wire_6656),
        .dout(new_Jinkela_wire_6657)
    );

    bfr new_Jinkela_buffer_4912 (
        .din(new_Jinkela_wire_6679),
        .dout(new_Jinkela_wire_6680)
    );

    bfr new_Jinkela_buffer_5669 (
        .din(new_Jinkela_wire_7633),
        .dout(new_Jinkela_wire_7634)
    );

    bfr new_Jinkela_buffer_4881 (
        .din(new_Jinkela_wire_6642),
        .dout(new_Jinkela_wire_6643)
    );

    bfr new_Jinkela_buffer_5734 (
        .din(new_Jinkela_wire_7716),
        .dout(new_Jinkela_wire_7717)
    );

    bfr new_Jinkela_buffer_4882 (
        .din(new_Jinkela_wire_6643),
        .dout(new_Jinkela_wire_6644)
    );

    bfr new_Jinkela_buffer_5692 (
        .din(new_Jinkela_wire_7666),
        .dout(new_Jinkela_wire_7667)
    );

    bfr new_Jinkela_buffer_5670 (
        .din(new_Jinkela_wire_7634),
        .dout(new_Jinkela_wire_7635)
    );

    bfr new_Jinkela_buffer_4883 (
        .din(new_Jinkela_wire_6644),
        .dout(new_Jinkela_wire_6645)
    );

    bfr new_Jinkela_buffer_5712 (
        .din(new_Jinkela_wire_7686),
        .dout(new_Jinkela_wire_7687)
    );

    bfr new_Jinkela_buffer_5671 (
        .din(new_Jinkela_wire_7635),
        .dout(new_Jinkela_wire_7636)
    );

    bfr new_Jinkela_buffer_4896 (
        .din(new_Jinkela_wire_6657),
        .dout(new_Jinkela_wire_6658)
    );

    bfr new_Jinkela_buffer_4884 (
        .din(new_Jinkela_wire_6645),
        .dout(new_Jinkela_wire_6646)
    );

    bfr new_Jinkela_buffer_5693 (
        .din(new_Jinkela_wire_7667),
        .dout(new_Jinkela_wire_7668)
    );

    bfr new_Jinkela_buffer_5672 (
        .din(new_Jinkela_wire_7636),
        .dout(new_Jinkela_wire_7637)
    );

    bfr new_Jinkela_buffer_4885 (
        .din(new_Jinkela_wire_6646),
        .dout(new_Jinkela_wire_6647)
    );

    bfr new_Jinkela_buffer_5673 (
        .din(new_Jinkela_wire_7637),
        .dout(new_Jinkela_wire_7638)
    );

    bfr new_Jinkela_buffer_4897 (
        .din(new_Jinkela_wire_6658),
        .dout(new_Jinkela_wire_6659)
    );

    bfr new_Jinkela_buffer_4886 (
        .din(new_Jinkela_wire_6647),
        .dout(new_Jinkela_wire_6648)
    );

    bfr new_Jinkela_buffer_5694 (
        .din(new_Jinkela_wire_7668),
        .dout(new_Jinkela_wire_7669)
    );

    bfr new_Jinkela_buffer_5674 (
        .din(new_Jinkela_wire_7638),
        .dout(new_Jinkela_wire_7639)
    );

    bfr new_Jinkela_buffer_4915 (
        .din(_0278_),
        .dout(new_Jinkela_wire_6710)
    );

    bfr new_Jinkela_buffer_4898 (
        .din(new_Jinkela_wire_6659),
        .dout(new_Jinkela_wire_6660)
    );

    bfr new_Jinkela_buffer_5735 (
        .din(new_Jinkela_wire_7717),
        .dout(new_Jinkela_wire_7718)
    );

    bfr new_Jinkela_buffer_5675 (
        .din(new_Jinkela_wire_7639),
        .dout(new_Jinkela_wire_7640)
    );

    spl4L new_Jinkela_splitter_680 (
        .a(new_Jinkela_wire_6685),
        .d(new_Jinkela_wire_6686),
        .e(new_Jinkela_wire_6691),
        .b(new_Jinkela_wire_6696),
        .c(new_Jinkela_wire_6701)
    );

    bfr new_Jinkela_buffer_5713 (
        .din(new_Jinkela_wire_7687),
        .dout(new_Jinkela_wire_7688)
    );

    bfr new_Jinkela_buffer_4899 (
        .din(new_Jinkela_wire_6660),
        .dout(new_Jinkela_wire_6661)
    );

    bfr new_Jinkela_buffer_5695 (
        .din(new_Jinkela_wire_7669),
        .dout(new_Jinkela_wire_7670)
    );

    bfr new_Jinkela_buffer_5676 (
        .din(new_Jinkela_wire_7640),
        .dout(new_Jinkela_wire_7641)
    );

    bfr new_Jinkela_buffer_4916 (
        .din(new_Jinkela_wire_6710),
        .dout(new_Jinkela_wire_6711)
    );

    spl4L new_Jinkela_splitter_679 (
        .a(new_Jinkela_wire_6680),
        .d(new_Jinkela_wire_6681),
        .e(new_Jinkela_wire_6682),
        .b(new_Jinkela_wire_6683),
        .c(new_Jinkela_wire_6684)
    );

    bfr new_Jinkela_buffer_4900 (
        .din(new_Jinkela_wire_6661),
        .dout(new_Jinkela_wire_6662)
    );

    bfr new_Jinkela_buffer_5677 (
        .din(new_Jinkela_wire_7641),
        .dout(new_Jinkela_wire_7642)
    );

    spl4L new_Jinkela_splitter_681 (
        .a(new_Jinkela_wire_6686),
        .d(new_Jinkela_wire_6687),
        .e(new_Jinkela_wire_6688),
        .b(new_Jinkela_wire_6689),
        .c(new_Jinkela_wire_6690)
    );

    bfr new_Jinkela_buffer_4901 (
        .din(new_Jinkela_wire_6662),
        .dout(new_Jinkela_wire_6663)
    );

    bfr new_Jinkela_buffer_5696 (
        .din(new_Jinkela_wire_7670),
        .dout(new_Jinkela_wire_7671)
    );

    bfr new_Jinkela_buffer_5678 (
        .din(new_Jinkela_wire_7642),
        .dout(new_Jinkela_wire_7643)
    );

    spl4L new_Jinkela_splitter_682 (
        .a(new_Jinkela_wire_6691),
        .d(new_Jinkela_wire_6692),
        .e(new_Jinkela_wire_6693),
        .b(new_Jinkela_wire_6694),
        .c(new_Jinkela_wire_6695)
    );

    bfr new_Jinkela_buffer_4902 (
        .din(new_Jinkela_wire_6663),
        .dout(new_Jinkela_wire_6664)
    );

    spl2 new_Jinkela_splitter_769 (
        .a(new_net_1),
        .b(new_Jinkela_wire_7785),
        .c(new_Jinkela_wire_7788)
    );

    spl2 new_Jinkela_splitter_759 (
        .a(new_Jinkela_wire_7643),
        .b(new_Jinkela_wire_7644),
        .c(new_Jinkela_wire_7645)
    );

    bfr new_Jinkela_buffer_4926 (
        .din(_0504_),
        .dout(new_Jinkela_wire_6721)
    );

    bfr new_Jinkela_buffer_4903 (
        .din(new_Jinkela_wire_6664),
        .dout(new_Jinkela_wire_6665)
    );

    bfr new_Jinkela_buffer_5714 (
        .din(new_Jinkela_wire_7688),
        .dout(new_Jinkela_wire_7689)
    );

    bfr new_Jinkela_buffer_5697 (
        .din(new_Jinkela_wire_7671),
        .dout(new_Jinkela_wire_7672)
    );

    spl4L new_Jinkela_splitter_683 (
        .a(new_Jinkela_wire_6696),
        .d(new_Jinkela_wire_6697),
        .e(new_Jinkela_wire_6698),
        .b(new_Jinkela_wire_6699),
        .c(new_Jinkela_wire_6700)
    );

    bfr new_Jinkela_buffer_5830 (
        .din(_1109_),
        .dout(new_Jinkela_wire_7823)
    );

    bfr new_Jinkela_buffer_4904 (
        .din(new_Jinkela_wire_6665),
        .dout(new_Jinkela_wire_6666)
    );

    bfr new_Jinkela_buffer_5698 (
        .din(new_Jinkela_wire_7672),
        .dout(new_Jinkela_wire_7673)
    );

    bfr new_Jinkela_buffer_5736 (
        .din(new_Jinkela_wire_7718),
        .dout(new_Jinkela_wire_7719)
    );

    spl4L new_Jinkela_splitter_684 (
        .a(new_Jinkela_wire_6701),
        .d(new_Jinkela_wire_6702),
        .e(new_Jinkela_wire_6703),
        .b(new_Jinkela_wire_6704),
        .c(new_Jinkela_wire_6705)
    );

    bfr new_Jinkela_buffer_5715 (
        .din(new_Jinkela_wire_7689),
        .dout(new_Jinkela_wire_7690)
    );

    bfr new_Jinkela_buffer_4905 (
        .din(new_Jinkela_wire_6666),
        .dout(new_Jinkela_wire_6667)
    );

    bfr new_Jinkela_buffer_5699 (
        .din(new_Jinkela_wire_7673),
        .dout(new_Jinkela_wire_7674)
    );

    bfr new_Jinkela_buffer_4906 (
        .din(new_Jinkela_wire_6667),
        .dout(new_Jinkela_wire_6668)
    );

    bfr new_Jinkela_buffer_5700 (
        .din(new_Jinkela_wire_7674),
        .dout(new_Jinkela_wire_7675)
    );

    bfr new_Jinkela_buffer_4917 (
        .din(_0848_),
        .dout(new_Jinkela_wire_6712)
    );

    bfr new_Jinkela_buffer_5799 (
        .din(new_Jinkela_wire_7783),
        .dout(new_Jinkela_wire_7784)
    );

    spl2 new_Jinkela_splitter_764 (
        .a(new_Jinkela_wire_7690),
        .b(new_Jinkela_wire_7691),
        .c(new_Jinkela_wire_7692)
    );

    bfr new_Jinkela_buffer_4907 (
        .din(new_Jinkela_wire_6668),
        .dout(new_Jinkela_wire_6669)
    );

    bfr new_Jinkela_buffer_5701 (
        .din(new_Jinkela_wire_7675),
        .dout(new_Jinkela_wire_7676)
    );

    bfr new_Jinkela_buffer_1879 (
        .din(new_Jinkela_wire_2951),
        .dout(new_Jinkela_wire_2952)
    );

    bfr new_Jinkela_buffer_4228 (
        .din(new_Jinkela_wire_5831),
        .dout(new_Jinkela_wire_5832)
    );

    bfr new_Jinkela_buffer_1953 (
        .din(new_Jinkela_wire_3032),
        .dout(new_Jinkela_wire_3033)
    );

    bfr new_Jinkela_buffer_4261 (
        .din(new_Jinkela_wire_5866),
        .dout(new_Jinkela_wire_5867)
    );

    bfr new_Jinkela_buffer_4262 (
        .din(_0730_),
        .dout(new_Jinkela_wire_5868)
    );

    spl2 new_Jinkela_splitter_409 (
        .a(_1116_),
        .b(new_Jinkela_wire_3094),
        .c(new_Jinkela_wire_3095)
    );

    bfr new_Jinkela_buffer_1880 (
        .din(new_Jinkela_wire_2952),
        .dout(new_Jinkela_wire_2953)
    );

    bfr new_Jinkela_buffer_4229 (
        .din(new_Jinkela_wire_5832),
        .dout(new_Jinkela_wire_5833)
    );

    bfr new_Jinkela_buffer_1916 (
        .din(new_Jinkela_wire_2991),
        .dout(new_Jinkela_wire_2992)
    );

    bfr new_Jinkela_buffer_4257 (
        .din(new_Jinkela_wire_5860),
        .dout(new_Jinkela_wire_5861)
    );

    bfr new_Jinkela_buffer_1881 (
        .din(new_Jinkela_wire_2953),
        .dout(new_Jinkela_wire_2954)
    );

    bfr new_Jinkela_buffer_4230 (
        .din(new_Jinkela_wire_5833),
        .dout(new_Jinkela_wire_5834)
    );

    spl3L new_Jinkela_splitter_404 (
        .a(_0936_),
        .d(new_Jinkela_wire_3063),
        .b(new_Jinkela_wire_3064),
        .c(new_Jinkela_wire_3065)
    );

    bfr new_Jinkela_buffer_1882 (
        .din(new_Jinkela_wire_2954),
        .dout(new_Jinkela_wire_2955)
    );

    bfr new_Jinkela_buffer_4231 (
        .din(new_Jinkela_wire_5834),
        .dout(new_Jinkela_wire_5835)
    );

    bfr new_Jinkela_buffer_1917 (
        .din(new_Jinkela_wire_2992),
        .dout(new_Jinkela_wire_2993)
    );

    bfr new_Jinkela_buffer_4258 (
        .din(new_Jinkela_wire_5861),
        .dout(new_Jinkela_wire_5862)
    );

    bfr new_Jinkela_buffer_1883 (
        .din(new_Jinkela_wire_2955),
        .dout(new_Jinkela_wire_2956)
    );

    bfr new_Jinkela_buffer_4232 (
        .din(new_Jinkela_wire_5835),
        .dout(new_Jinkela_wire_5836)
    );

    spl2 new_Jinkela_splitter_403 (
        .a(_1011_),
        .b(new_Jinkela_wire_3061),
        .c(new_Jinkela_wire_3062)
    );

    spl2 new_Jinkela_splitter_616 (
        .a(new_net_7),
        .b(new_Jinkela_wire_5878),
        .c(new_Jinkela_wire_5880)
    );

    bfr new_Jinkela_buffer_4288 (
        .din(_0617_),
        .dout(new_Jinkela_wire_5900)
    );

    bfr new_Jinkela_buffer_1884 (
        .din(new_Jinkela_wire_2956),
        .dout(new_Jinkela_wire_2957)
    );

    bfr new_Jinkela_buffer_4233 (
        .din(new_Jinkela_wire_5836),
        .dout(new_Jinkela_wire_5837)
    );

    bfr new_Jinkela_buffer_1918 (
        .din(new_Jinkela_wire_2993),
        .dout(new_Jinkela_wire_2994)
    );

    bfr new_Jinkela_buffer_4259 (
        .din(new_Jinkela_wire_5862),
        .dout(new_Jinkela_wire_5863)
    );

    bfr new_Jinkela_buffer_1885 (
        .din(new_Jinkela_wire_2957),
        .dout(new_Jinkela_wire_2958)
    );

    bfr new_Jinkela_buffer_4234 (
        .din(new_Jinkela_wire_5837),
        .dout(new_Jinkela_wire_5838)
    );

    bfr new_Jinkela_buffer_1954 (
        .din(new_Jinkela_wire_3033),
        .dout(new_Jinkela_wire_3034)
    );

    bfr new_Jinkela_buffer_4263 (
        .din(new_Jinkela_wire_5868),
        .dout(new_Jinkela_wire_5869)
    );

    bfr new_Jinkela_buffer_1886 (
        .din(new_Jinkela_wire_2958),
        .dout(new_Jinkela_wire_2959)
    );

    bfr new_Jinkela_buffer_4235 (
        .din(new_Jinkela_wire_5838),
        .dout(new_Jinkela_wire_5839)
    );

    bfr new_Jinkela_buffer_1919 (
        .din(new_Jinkela_wire_2994),
        .dout(new_Jinkela_wire_2995)
    );

    spl2 new_Jinkela_splitter_619 (
        .a(_0171_),
        .b(new_Jinkela_wire_5904),
        .c(new_Jinkela_wire_5905)
    );

    bfr new_Jinkela_buffer_4273 (
        .din(new_Jinkela_wire_5884),
        .dout(new_Jinkela_wire_5885)
    );

    bfr new_Jinkela_buffer_1887 (
        .din(new_Jinkela_wire_2959),
        .dout(new_Jinkela_wire_2960)
    );

    bfr new_Jinkela_buffer_4236 (
        .din(new_Jinkela_wire_5839),
        .dout(new_Jinkela_wire_5840)
    );

    bfr new_Jinkela_buffer_4264 (
        .din(new_Jinkela_wire_5869),
        .dout(new_Jinkela_wire_5870)
    );

    bfr new_Jinkela_buffer_1995 (
        .din(_1083_),
        .dout(new_Jinkela_wire_3084)
    );

    bfr new_Jinkela_buffer_1888 (
        .din(new_Jinkela_wire_2960),
        .dout(new_Jinkela_wire_2961)
    );

    bfr new_Jinkela_buffer_4237 (
        .din(new_Jinkela_wire_5840),
        .dout(new_Jinkela_wire_5841)
    );

    bfr new_Jinkela_buffer_1920 (
        .din(new_Jinkela_wire_2995),
        .dout(new_Jinkela_wire_2996)
    );

    bfr new_Jinkela_buffer_4272 (
        .din(new_Jinkela_wire_5878),
        .dout(new_Jinkela_wire_5879)
    );

    spl4L new_Jinkela_splitter_617 (
        .a(new_Jinkela_wire_5880),
        .d(new_Jinkela_wire_5881),
        .e(new_Jinkela_wire_5882),
        .b(new_Jinkela_wire_5883),
        .c(new_Jinkela_wire_5884)
    );

    bfr new_Jinkela_buffer_1889 (
        .din(new_Jinkela_wire_2961),
        .dout(new_Jinkela_wire_2962)
    );

    bfr new_Jinkela_buffer_4238 (
        .din(new_Jinkela_wire_5841),
        .dout(new_Jinkela_wire_5842)
    );

    bfr new_Jinkela_buffer_1955 (
        .din(new_Jinkela_wire_3034),
        .dout(new_Jinkela_wire_3035)
    );

    bfr new_Jinkela_buffer_4265 (
        .din(new_Jinkela_wire_5870),
        .dout(new_Jinkela_wire_5871)
    );

    bfr new_Jinkela_buffer_1890 (
        .din(new_Jinkela_wire_2962),
        .dout(new_Jinkela_wire_2963)
    );

    bfr new_Jinkela_buffer_4239 (
        .din(new_Jinkela_wire_5842),
        .dout(new_Jinkela_wire_5843)
    );

    bfr new_Jinkela_buffer_1921 (
        .din(new_Jinkela_wire_2996),
        .dout(new_Jinkela_wire_2997)
    );

    spl2 new_Jinkela_splitter_618 (
        .a(_0618_),
        .b(new_Jinkela_wire_5902),
        .c(new_Jinkela_wire_5903)
    );

    bfr new_Jinkela_buffer_1891 (
        .din(new_Jinkela_wire_2963),
        .dout(new_Jinkela_wire_2964)
    );

    bfr new_Jinkela_buffer_4240 (
        .din(new_Jinkela_wire_5843),
        .dout(new_Jinkela_wire_5844)
    );

    bfr new_Jinkela_buffer_4266 (
        .din(new_Jinkela_wire_5871),
        .dout(new_Jinkela_wire_5872)
    );

    spl3L new_Jinkela_splitter_408 (
        .a(_0947_),
        .d(new_Jinkela_wire_3089),
        .b(new_Jinkela_wire_3090),
        .c(new_Jinkela_wire_3091)
    );

    bfr new_Jinkela_buffer_1892 (
        .din(new_Jinkela_wire_2964),
        .dout(new_Jinkela_wire_2965)
    );

    bfr new_Jinkela_buffer_4241 (
        .din(new_Jinkela_wire_5844),
        .dout(new_Jinkela_wire_5845)
    );

    bfr new_Jinkela_buffer_1922 (
        .din(new_Jinkela_wire_2997),
        .dout(new_Jinkela_wire_2998)
    );

    bfr new_Jinkela_buffer_1893 (
        .din(new_Jinkela_wire_2965),
        .dout(new_Jinkela_wire_2966)
    );

    bfr new_Jinkela_buffer_4242 (
        .din(new_Jinkela_wire_5845),
        .dout(new_Jinkela_wire_5846)
    );

    bfr new_Jinkela_buffer_1956 (
        .din(new_Jinkela_wire_3035),
        .dout(new_Jinkela_wire_3036)
    );

    bfr new_Jinkela_buffer_4267 (
        .din(new_Jinkela_wire_5872),
        .dout(new_Jinkela_wire_5873)
    );

    bfr new_Jinkela_buffer_1894 (
        .din(new_Jinkela_wire_2966),
        .dout(new_Jinkela_wire_2967)
    );

    bfr new_Jinkela_buffer_4243 (
        .din(new_Jinkela_wire_5846),
        .dout(new_Jinkela_wire_5847)
    );

    bfr new_Jinkela_buffer_1923 (
        .din(new_Jinkela_wire_2998),
        .dout(new_Jinkela_wire_2999)
    );

    bfr new_Jinkela_buffer_1895 (
        .din(new_Jinkela_wire_2967),
        .dout(new_Jinkela_wire_2968)
    );

    bfr new_Jinkela_buffer_4244 (
        .din(new_Jinkela_wire_5847),
        .dout(new_Jinkela_wire_5848)
    );

    bfr new_Jinkela_buffer_1981 (
        .din(new_Jinkela_wire_3065),
        .dout(new_Jinkela_wire_3066)
    );

    bfr new_Jinkela_buffer_4268 (
        .din(new_Jinkela_wire_5873),
        .dout(new_Jinkela_wire_5874)
    );

    bfr new_Jinkela_buffer_1896 (
        .din(new_Jinkela_wire_2968),
        .dout(new_Jinkela_wire_2969)
    );

    bfr new_Jinkela_buffer_4245 (
        .din(new_Jinkela_wire_5848),
        .dout(new_Jinkela_wire_5849)
    );

    bfr new_Jinkela_buffer_1924 (
        .din(new_Jinkela_wire_2999),
        .dout(new_Jinkela_wire_3000)
    );

    bfr new_Jinkela_buffer_4289 (
        .din(new_Jinkela_wire_5900),
        .dout(new_Jinkela_wire_5901)
    );

    bfr new_Jinkela_buffer_1897 (
        .din(new_Jinkela_wire_2969),
        .dout(new_Jinkela_wire_2970)
    );

    bfr new_Jinkela_buffer_4246 (
        .din(new_Jinkela_wire_5849),
        .dout(new_Jinkela_wire_5850)
    );

    bfr new_Jinkela_buffer_1957 (
        .din(new_Jinkela_wire_3036),
        .dout(new_Jinkela_wire_3037)
    );

    bfr new_Jinkela_buffer_4269 (
        .din(new_Jinkela_wire_5874),
        .dout(new_Jinkela_wire_5875)
    );

    bfr new_Jinkela_buffer_1898 (
        .din(new_Jinkela_wire_2970),
        .dout(new_Jinkela_wire_2971)
    );

    bfr new_Jinkela_buffer_4247 (
        .din(new_Jinkela_wire_5850),
        .dout(new_Jinkela_wire_5851)
    );

    bfr new_Jinkela_buffer_1925 (
        .din(new_Jinkela_wire_3000),
        .dout(new_Jinkela_wire_3001)
    );

    bfr new_Jinkela_buffer_1899 (
        .din(new_Jinkela_wire_2971),
        .dout(new_Jinkela_wire_2972)
    );

    bfr new_Jinkela_buffer_4248 (
        .din(new_Jinkela_wire_5851),
        .dout(new_Jinkela_wire_5852)
    );

    bfr new_Jinkela_buffer_4270 (
        .din(new_Jinkela_wire_5875),
        .dout(new_Jinkela_wire_5876)
    );

    spl3L new_Jinkela_splitter_328 (
        .a(new_Jinkela_wire_1879),
        .d(new_Jinkela_wire_1880),
        .b(new_Jinkela_wire_1881),
        .c(new_Jinkela_wire_1882)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1811),
        .dout(new_Jinkela_wire_1812)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1832),
        .dout(new_Jinkela_wire_1833)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1863),
        .dout(new_Jinkela_wire_1864)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1833),
        .dout(new_Jinkela_wire_1834)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1814),
        .dout(new_Jinkela_wire_1815)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1891),
        .dout(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1815),
        .dout(new_Jinkela_wire_1816)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1834),
        .dout(new_Jinkela_wire_1835)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1864),
        .dout(new_Jinkela_wire_1865)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1817),
        .dout(new_Jinkela_wire_1818)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1818),
        .dout(new_Jinkela_wire_1819)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1882),
        .dout(new_Jinkela_wire_1883)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1819),
        .dout(new_Jinkela_wire_1820)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1865),
        .dout(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    spl2 new_Jinkela_splitter_334 (
        .a(_1179_),
        .b(new_Jinkela_wire_1944),
        .c(new_Jinkela_wire_1945)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1838),
        .dout(new_Jinkela_wire_1839)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1866),
        .dout(new_Jinkela_wire_1867)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1839),
        .dout(new_Jinkela_wire_1840)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1892),
        .dout(new_Jinkela_wire_1893)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1840),
        .dout(new_Jinkela_wire_1841)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1867),
        .dout(new_Jinkela_wire_1868)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1841),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_988 (
        .din(new_Jinkela_wire_1883),
        .dout(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1842),
        .dout(new_Jinkela_wire_1843)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1868),
        .dout(new_Jinkela_wire_1869)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1843),
        .dout(new_Jinkela_wire_1844)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(_0086_),
        .dout(new_Jinkela_wire_1915)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1844),
        .dout(new_Jinkela_wire_1845)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1869),
        .dout(new_Jinkela_wire_1870)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1845),
        .dout(new_Jinkela_wire_1846)
    );

    spl2 new_Jinkela_splitter_329 (
        .a(new_Jinkela_wire_1884),
        .b(new_Jinkela_wire_1885),
        .c(new_Jinkela_wire_1886)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1846),
        .dout(new_Jinkela_wire_1847)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1870),
        .dout(new_Jinkela_wire_1871)
    );

    and_bi _2465_ (
        .a(new_Jinkela_wire_5653),
        .b(_0458_),
        .c(_0459_)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1847),
        .dout(new_Jinkela_wire_1848)
    );

    inv _1294_ (
        .din(new_Jinkela_wire_1402),
        .dout(_0601_)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1886),
        .dout(new_Jinkela_wire_1887)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1871),
        .dout(new_Jinkela_wire_1872)
    );

    bfr new_Jinkela_buffer_1900 (
        .din(new_Jinkela_wire_2972),
        .dout(new_Jinkela_wire_2973)
    );

    bfr new_Jinkela_buffer_4918 (
        .din(new_Jinkela_wire_6712),
        .dout(new_Jinkela_wire_6713)
    );

    bfr new_Jinkela_buffer_5716 (
        .din(new_Jinkela_wire_7692),
        .dout(new_Jinkela_wire_7693)
    );

    bfr new_Jinkela_buffer_1926 (
        .din(new_Jinkela_wire_3001),
        .dout(new_Jinkela_wire_3002)
    );

    bfr new_Jinkela_buffer_4908 (
        .din(new_Jinkela_wire_6669),
        .dout(new_Jinkela_wire_6670)
    );

    bfr new_Jinkela_buffer_5702 (
        .din(new_Jinkela_wire_7676),
        .dout(new_Jinkela_wire_7677)
    );

    bfr new_Jinkela_buffer_1901 (
        .din(new_Jinkela_wire_2973),
        .dout(new_Jinkela_wire_2974)
    );

    spl2 new_Jinkela_splitter_686 (
        .a(_1170_),
        .b(new_Jinkela_wire_6750),
        .c(new_Jinkela_wire_6751)
    );

    spl2 new_Jinkela_splitter_687 (
        .a(_0012_),
        .b(new_Jinkela_wire_6752),
        .c(new_Jinkela_wire_6753)
    );

    bfr new_Jinkela_buffer_5759 (
        .din(new_Jinkela_wire_7743),
        .dout(new_Jinkela_wire_7744)
    );

    bfr new_Jinkela_buffer_1958 (
        .din(new_Jinkela_wire_3037),
        .dout(new_Jinkela_wire_3038)
    );

    bfr new_Jinkela_buffer_4919 (
        .din(new_Jinkela_wire_6713),
        .dout(new_Jinkela_wire_6714)
    );

    bfr new_Jinkela_buffer_5703 (
        .din(new_Jinkela_wire_7677),
        .dout(new_Jinkela_wire_7678)
    );

    bfr new_Jinkela_buffer_1902 (
        .din(new_Jinkela_wire_2974),
        .dout(new_Jinkela_wire_2975)
    );

    bfr new_Jinkela_buffer_4927 (
        .din(new_Jinkela_wire_6721),
        .dout(new_Jinkela_wire_6722)
    );

    bfr new_Jinkela_buffer_5737 (
        .din(new_Jinkela_wire_7719),
        .dout(new_Jinkela_wire_7720)
    );

    bfr new_Jinkela_buffer_1927 (
        .din(new_Jinkela_wire_3002),
        .dout(new_Jinkela_wire_3003)
    );

    bfr new_Jinkela_buffer_4920 (
        .din(new_Jinkela_wire_6714),
        .dout(new_Jinkela_wire_6715)
    );

    bfr new_Jinkela_buffer_5704 (
        .din(new_Jinkela_wire_7678),
        .dout(new_Jinkela_wire_7679)
    );

    bfr new_Jinkela_buffer_1903 (
        .din(new_Jinkela_wire_2975),
        .dout(new_Jinkela_wire_2976)
    );

    spl3L new_Jinkela_splitter_690 (
        .a(_0863_),
        .d(new_Jinkela_wire_6764),
        .b(new_Jinkela_wire_6765),
        .c(new_Jinkela_wire_6766)
    );

    bfr new_Jinkela_buffer_5717 (
        .din(new_Jinkela_wire_7693),
        .dout(new_Jinkela_wire_7694)
    );

    bfr new_Jinkela_buffer_1982 (
        .din(new_Jinkela_wire_3066),
        .dout(new_Jinkela_wire_3067)
    );

    bfr new_Jinkela_buffer_4921 (
        .din(new_Jinkela_wire_6715),
        .dout(new_Jinkela_wire_6716)
    );

    bfr new_Jinkela_buffer_5705 (
        .din(new_Jinkela_wire_7679),
        .dout(new_Jinkela_wire_7680)
    );

    bfr new_Jinkela_buffer_1904 (
        .din(new_Jinkela_wire_2976),
        .dout(new_Jinkela_wire_2977)
    );

    bfr new_Jinkela_buffer_4928 (
        .din(new_Jinkela_wire_6722),
        .dout(new_Jinkela_wire_6723)
    );

    bfr new_Jinkela_buffer_1928 (
        .din(new_Jinkela_wire_3003),
        .dout(new_Jinkela_wire_3004)
    );

    bfr new_Jinkela_buffer_4922 (
        .din(new_Jinkela_wire_6716),
        .dout(new_Jinkela_wire_6717)
    );

    bfr new_Jinkela_buffer_5706 (
        .din(new_Jinkela_wire_7680),
        .dout(new_Jinkela_wire_7681)
    );

    bfr new_Jinkela_buffer_1905 (
        .din(new_Jinkela_wire_2977),
        .dout(new_Jinkela_wire_2978)
    );

    bfr new_Jinkela_buffer_5738 (
        .din(new_Jinkela_wire_7720),
        .dout(new_Jinkela_wire_7721)
    );

    bfr new_Jinkela_buffer_5718 (
        .din(new_Jinkela_wire_7694),
        .dout(new_Jinkela_wire_7695)
    );

    bfr new_Jinkela_buffer_1959 (
        .din(new_Jinkela_wire_3038),
        .dout(new_Jinkela_wire_3039)
    );

    bfr new_Jinkela_buffer_4923 (
        .din(new_Jinkela_wire_6717),
        .dout(new_Jinkela_wire_6718)
    );

    spl2 new_Jinkela_splitter_82 (
        .a(G101),
        .b(new_Jinkela_wire_400),
        .c(new_Jinkela_wire_405)
    );

    bfr new_Jinkela_buffer_1906 (
        .din(new_Jinkela_wire_2978),
        .dout(new_Jinkela_wire_2979)
    );

    bfr new_Jinkela_buffer_4929 (
        .din(new_Jinkela_wire_6723),
        .dout(new_Jinkela_wire_6724)
    );

    spl2 new_Jinkela_splitter_765 (
        .a(new_Jinkela_wire_7695),
        .b(new_Jinkela_wire_7696),
        .c(new_Jinkela_wire_7697)
    );

    spl2 new_Jinkela_splitter_772 (
        .a(_0130_),
        .b(new_Jinkela_wire_7824),
        .c(new_Jinkela_wire_7825)
    );

    bfr new_Jinkela_buffer_1929 (
        .din(new_Jinkela_wire_3004),
        .dout(new_Jinkela_wire_3005)
    );

    bfr new_Jinkela_buffer_4924 (
        .din(new_Jinkela_wire_6718),
        .dout(new_Jinkela_wire_6719)
    );

    bfr new_Jinkela_buffer_5719 (
        .din(new_Jinkela_wire_7697),
        .dout(new_Jinkela_wire_7698)
    );

    bfr new_Jinkela_buffer_1907 (
        .din(new_Jinkela_wire_2979),
        .dout(new_Jinkela_wire_2980)
    );

    bfr new_Jinkela_buffer_4955 (
        .din(_0734_),
        .dout(new_Jinkela_wire_6754)
    );

    bfr new_Jinkela_buffer_4956 (
        .din(_0338_),
        .dout(new_Jinkela_wire_6757)
    );

    bfr new_Jinkela_buffer_5760 (
        .din(new_Jinkela_wire_7744),
        .dout(new_Jinkela_wire_7745)
    );

    bfr new_Jinkela_buffer_1996 (
        .din(new_Jinkela_wire_3084),
        .dout(new_Jinkela_wire_3085)
    );

    bfr new_Jinkela_buffer_4925 (
        .din(new_Jinkela_wire_6719),
        .dout(new_Jinkela_wire_6720)
    );

    bfr new_Jinkela_buffer_5739 (
        .din(new_Jinkela_wire_7721),
        .dout(new_Jinkela_wire_7722)
    );

    bfr new_Jinkela_buffer_1908 (
        .din(new_Jinkela_wire_2980),
        .dout(new_Jinkela_wire_2981)
    );

    bfr new_Jinkela_buffer_4930 (
        .din(new_Jinkela_wire_6724),
        .dout(new_Jinkela_wire_6725)
    );

    or_bi _1273_ (
        .a(new_Jinkela_wire_6503),
        .b(new_Jinkela_wire_551),
        .c(new_net_2351)
    );

    spl2 new_Jinkela_splitter_766 (
        .a(new_Jinkela_wire_7698),
        .b(new_Jinkela_wire_7699),
        .c(new_Jinkela_wire_7700)
    );

    bfr new_Jinkela_buffer_1930 (
        .din(new_Jinkela_wire_3005),
        .dout(new_Jinkela_wire_3006)
    );

    spl2 new_Jinkela_splitter_688 (
        .a(_0687_),
        .b(new_Jinkela_wire_6755),
        .c(new_Jinkela_wire_6756)
    );

    and_bb _1251_ (
        .a(new_Jinkela_wire_1399),
        .b(new_Jinkela_wire_870),
        .c(_0581_)
    );

    bfr new_Jinkela_buffer_4958 (
        .din(new_Jinkela_wire_6758),
        .dout(new_Jinkela_wire_6759)
    );

    bfr new_Jinkela_buffer_5720 (
        .din(new_Jinkela_wire_7700),
        .dout(new_Jinkela_wire_7701)
    );

    and_bi _1249_ (
        .a(new_Jinkela_wire_973),
        .b(new_Jinkela_wire_884),
        .c(_0579_)
    );

    bfr new_Jinkela_buffer_1909 (
        .din(new_Jinkela_wire_2981),
        .dout(new_Jinkela_wire_2982)
    );

    bfr new_Jinkela_buffer_4931 (
        .din(new_Jinkela_wire_6725),
        .dout(new_Jinkela_wire_6726)
    );

    and_ii _1250_ (
        .a(_0579_),
        .b(_0578_),
        .c(_0580_)
    );

    bfr new_Jinkela_buffer_1960 (
        .din(new_Jinkela_wire_3039),
        .dout(new_Jinkela_wire_3040)
    );

    bfr new_Jinkela_buffer_5740 (
        .din(new_Jinkela_wire_7722),
        .dout(new_Jinkela_wire_7723)
    );

    and_bb _1248_ (
        .a(new_Jinkela_wire_526),
        .b(new_Jinkela_wire_875),
        .c(_0578_)
    );

    bfr new_Jinkela_buffer_1910 (
        .din(new_Jinkela_wire_2982),
        .dout(new_Jinkela_wire_2983)
    );

    bfr new_Jinkela_buffer_4932 (
        .din(new_Jinkela_wire_6726),
        .dout(new_Jinkela_wire_6727)
    );

    and_bi _1252_ (
        .a(new_Jinkela_wire_1379),
        .b(new_Jinkela_wire_873),
        .c(_0582_)
    );

    bfr new_Jinkela_buffer_5721 (
        .din(new_Jinkela_wire_7701),
        .dout(new_Jinkela_wire_7702)
    );

    bfr new_Jinkela_buffer_1931 (
        .din(new_Jinkela_wire_3006),
        .dout(new_Jinkela_wire_3007)
    );

    bfr new_Jinkela_buffer_4957 (
        .din(_0933_),
        .dout(new_Jinkela_wire_6758)
    );

    and_bi _1256_ (
        .a(new_Jinkela_wire_2841),
        .b(new_Jinkela_wire_5284),
        .c(new_net_1)
    );

    bfr new_Jinkela_buffer_5761 (
        .din(new_Jinkela_wire_7745),
        .dout(new_Jinkela_wire_7746)
    );

    bfr new_Jinkela_buffer_1911 (
        .din(new_Jinkela_wire_2983),
        .dout(new_Jinkela_wire_2984)
    );

    bfr new_Jinkela_buffer_4933 (
        .din(new_Jinkela_wire_6727),
        .dout(new_Jinkela_wire_6728)
    );

    bfr new_Jinkela_buffer_5741 (
        .din(new_Jinkela_wire_7723),
        .dout(new_Jinkela_wire_7724)
    );

    and_ii _1255_ (
        .a(new_Jinkela_wire_4577),
        .b(new_Jinkela_wire_2773),
        .c(_0585_)
    );

    bfr new_Jinkela_buffer_5722 (
        .din(new_Jinkela_wire_7702),
        .dout(new_Jinkela_wire_7703)
    );

    spl2 new_Jinkela_splitter_691 (
        .a(_0079_),
        .b(new_Jinkela_wire_6768),
        .c(new_Jinkela_wire_6769)
    );

    and_ii _1253_ (
        .a(_0582_),
        .b(_0581_),
        .c(_0583_)
    );

    spl2 new_Jinkela_splitter_405 (
        .a(new_Jinkela_wire_3067),
        .b(new_Jinkela_wire_3068),
        .c(new_Jinkela_wire_3069)
    );

    bfr new_Jinkela_buffer_1912 (
        .din(new_Jinkela_wire_2984),
        .dout(new_Jinkela_wire_2985)
    );

    bfr new_Jinkela_buffer_4934 (
        .din(new_Jinkela_wire_6728),
        .dout(new_Jinkela_wire_6729)
    );

    bfr new_Jinkela_buffer_5723 (
        .din(new_Jinkela_wire_7703),
        .dout(new_Jinkela_wire_7704)
    );

    inv _1265_ (
        .din(new_Jinkela_wire_1235),
        .dout(new_net_2465)
    );

    bfr new_Jinkela_buffer_1932 (
        .din(new_Jinkela_wire_3007),
        .dout(new_Jinkela_wire_3008)
    );

    or_ii _1254_ (
        .a(new_Jinkela_wire_4578),
        .b(new_Jinkela_wire_2772),
        .c(_0584_)
    );

    bfr new_Jinkela_buffer_4990 (
        .din(_0097_),
        .dout(new_Jinkela_wire_6804)
    );

    inv _1257_ (
        .din(new_Jinkela_wire_573),
        .dout(new_net_2379)
    );

    bfr new_Jinkela_buffer_1961 (
        .din(new_Jinkela_wire_3040),
        .dout(new_Jinkela_wire_3041)
    );

    bfr new_Jinkela_buffer_4935 (
        .din(new_Jinkela_wire_6729),
        .dout(new_Jinkela_wire_6730)
    );

    bfr new_Jinkela_buffer_5724 (
        .din(new_Jinkela_wire_7704),
        .dout(new_Jinkela_wire_7705)
    );

    bfr new_Jinkela_buffer_5742 (
        .din(new_Jinkela_wire_7724),
        .dout(new_Jinkela_wire_7725)
    );

    inv _1258_ (
        .din(new_Jinkela_wire_522),
        .dout(new_net_2487)
    );

    bfr new_Jinkela_buffer_1933 (
        .din(new_Jinkela_wire_3008),
        .dout(new_Jinkela_wire_3009)
    );

    bfr new_Jinkela_buffer_4961 (
        .din(new_Jinkela_wire_6766),
        .dout(new_Jinkela_wire_6767)
    );

    spl2 new_Jinkela_splitter_689 (
        .a(new_Jinkela_wire_6759),
        .b(new_Jinkela_wire_6760),
        .c(new_Jinkela_wire_6761)
    );

    inv _1259_ (
        .din(new_Jinkela_wire_116),
        .dout(new_net_2415)
    );

    bfr new_Jinkela_buffer_4936 (
        .din(new_Jinkela_wire_6730),
        .dout(new_Jinkela_wire_6731)
    );

    bfr new_Jinkela_buffer_1983 (
        .din(new_Jinkela_wire_3069),
        .dout(new_Jinkela_wire_3070)
    );

    bfr new_Jinkela_buffer_5725 (
        .din(new_Jinkela_wire_7705),
        .dout(new_Jinkela_wire_7706)
    );

    inv _1260_ (
        .din(G151),
        .dout(new_net_24)
    );

    bfr new_Jinkela_buffer_1934 (
        .din(new_Jinkela_wire_3009),
        .dout(new_Jinkela_wire_3010)
    );

    bfr new_Jinkela_buffer_4959 (
        .din(new_Jinkela_wire_6761),
        .dout(new_Jinkela_wire_6762)
    );

    bfr new_Jinkela_buffer_5762 (
        .din(new_Jinkela_wire_7746),
        .dout(new_Jinkela_wire_7747)
    );

    inv _1261_ (
        .din(new_Jinkela_wire_1429),
        .dout(new_net_2359)
    );

    bfr new_Jinkela_buffer_1962 (
        .din(new_Jinkela_wire_3041),
        .dout(new_Jinkela_wire_3042)
    );

    bfr new_Jinkela_buffer_4937 (
        .din(new_Jinkela_wire_6731),
        .dout(new_Jinkela_wire_6732)
    );

    bfr new_Jinkela_buffer_5726 (
        .din(new_Jinkela_wire_7706),
        .dout(new_Jinkela_wire_7707)
    );

    bfr new_Jinkela_buffer_5743 (
        .din(new_Jinkela_wire_7725),
        .dout(new_Jinkela_wire_7726)
    );

    inv _1262_ (
        .din(new_Jinkela_wire_773),
        .dout(new_net_2463)
    );

    bfr new_Jinkela_buffer_1935 (
        .din(new_Jinkela_wire_3010),
        .dout(new_Jinkela_wire_3011)
    );

    inv _1263_ (
        .din(new_Jinkela_wire_896),
        .dout(new_net_2429)
    );

    bfr new_Jinkela_buffer_4938 (
        .din(new_Jinkela_wire_6732),
        .dout(new_Jinkela_wire_6733)
    );

    bfr new_Jinkela_buffer_1997 (
        .din(new_Jinkela_wire_3085),
        .dout(new_Jinkela_wire_3086)
    );

    bfr new_Jinkela_buffer_5727 (
        .din(new_Jinkela_wire_7707),
        .dout(new_Jinkela_wire_7708)
    );

    inv _1264_ (
        .din(new_Jinkela_wire_1345),
        .dout(new_net_2)
    );

    bfr new_Jinkela_buffer_1936 (
        .din(new_Jinkela_wire_3011),
        .dout(new_Jinkela_wire_3012)
    );

    bfr new_Jinkela_buffer_4963 (
        .din(new_Jinkela_wire_6770),
        .dout(new_Jinkela_wire_6771)
    );

    spl4L new_Jinkela_splitter_771 (
        .a(new_Jinkela_wire_7788),
        .d(new_Jinkela_wire_7789),
        .e(new_Jinkela_wire_7790),
        .b(new_Jinkela_wire_7791),
        .c(new_Jinkela_wire_7792)
    );

    bfr new_Jinkela_buffer_1963 (
        .din(new_Jinkela_wire_3042),
        .dout(new_Jinkela_wire_3043)
    );

    bfr new_Jinkela_buffer_4939 (
        .din(new_Jinkela_wire_6733),
        .dout(new_Jinkela_wire_6734)
    );

    bfr new_Jinkela_buffer_5744 (
        .din(new_Jinkela_wire_7726),
        .dout(new_Jinkela_wire_7727)
    );

    inv _1266_ (
        .din(new_Jinkela_wire_88),
        .dout(new_net_2441)
    );

    bfr new_Jinkela_buffer_5728 (
        .din(new_Jinkela_wire_7708),
        .dout(new_Jinkela_wire_7709)
    );

    bfr new_Jinkela_buffer_1937 (
        .din(new_Jinkela_wire_3012),
        .dout(new_Jinkela_wire_3013)
    );

    bfr new_Jinkela_buffer_4962 (
        .din(new_net_2509),
        .dout(new_Jinkela_wire_6770)
    );

    inv _1267_ (
        .din(new_Jinkela_wire_297),
        .dout(new_net_2403)
    );

    bfr new_Jinkela_buffer_4960 (
        .din(new_Jinkela_wire_6762),
        .dout(new_Jinkela_wire_6763)
    );

    bfr new_Jinkela_buffer_4940 (
        .din(new_Jinkela_wire_6734),
        .dout(new_Jinkela_wire_6735)
    );

    spl2 new_Jinkela_splitter_770 (
        .a(new_Jinkela_wire_7785),
        .b(new_Jinkela_wire_7786),
        .c(new_Jinkela_wire_7787)
    );

    inv _1268_ (
        .din(new_Jinkela_wire_1133),
        .dout(new_net_2419)
    );

    spl3L new_Jinkela_splitter_410 (
        .a(_1238_),
        .d(new_Jinkela_wire_3096),
        .b(new_Jinkela_wire_3097),
        .c(new_Jinkela_wire_3098)
    );

    bfr new_Jinkela_buffer_5729 (
        .din(new_Jinkela_wire_7709),
        .dout(new_Jinkela_wire_7710)
    );

    bfr new_Jinkela_buffer_1938 (
        .din(new_Jinkela_wire_3013),
        .dout(new_Jinkela_wire_3014)
    );

    inv _1269_ (
        .din(new_Jinkela_wire_1135),
        .dout(new_net_2375)
    );

    bfr new_Jinkela_buffer_5763 (
        .din(new_Jinkela_wire_7747),
        .dout(new_Jinkela_wire_7748)
    );

    bfr new_Jinkela_buffer_1964 (
        .din(new_Jinkela_wire_3043),
        .dout(new_Jinkela_wire_3044)
    );

    bfr new_Jinkela_buffer_4941 (
        .din(new_Jinkela_wire_6735),
        .dout(new_Jinkela_wire_6736)
    );

    bfr new_Jinkela_buffer_5745 (
        .din(new_Jinkela_wire_7727),
        .dout(new_Jinkela_wire_7728)
    );

    or_bi _1270_ (
        .a(new_Jinkela_wire_1368),
        .b(new_Jinkela_wire_843),
        .c(new_net_2389)
    );

    bfr new_Jinkela_buffer_5730 (
        .din(new_Jinkela_wire_7710),
        .dout(new_Jinkela_wire_7711)
    );

    bfr new_Jinkela_buffer_1939 (
        .din(new_Jinkela_wire_3014),
        .dout(new_Jinkela_wire_3015)
    );

    spl2 new_Jinkela_splitter_692 (
        .a(new_net_20),
        .b(new_Jinkela_wire_6790),
        .c(new_Jinkela_wire_6792)
    );

    or_ii _1271_ (
        .a(G154),
        .b(G136),
        .c(new_net_13)
    );

    bfr new_Jinkela_buffer_1998 (
        .din(new_Jinkela_wire_3091),
        .dout(new_Jinkela_wire_3092)
    );

    bfr new_Jinkela_buffer_4942 (
        .din(new_Jinkela_wire_6736),
        .dout(new_Jinkela_wire_6737)
    );

    or_ii _1272_ (
        .a(new_Jinkela_wire_844),
        .b(new_Jinkela_wire_248),
        .c(new_net_0)
    );

    bfr new_Jinkela_buffer_1984 (
        .din(new_Jinkela_wire_3070),
        .dout(new_Jinkela_wire_3071)
    );

    bfr new_Jinkela_buffer_5731 (
        .din(new_Jinkela_wire_7711),
        .dout(new_Jinkela_wire_7712)
    );

    bfr new_Jinkela_buffer_1940 (
        .din(new_Jinkela_wire_3015),
        .dout(new_Jinkela_wire_3016)
    );

    and_bi _1403_ (
        .a(_0704_),
        .b(_0705_),
        .c(_0706_)
    );

    and_ii _2117_ (
        .a(new_Jinkela_wire_6625),
        .b(new_Jinkela_wire_4254),
        .c(_0154_)
    );

    or_bb _1404_ (
        .a(new_Jinkela_wire_5052),
        .b(new_Jinkela_wire_1077),
        .c(_0707_)
    );

    and_bb _2118_ (
        .a(new_Jinkela_wire_6626),
        .b(new_Jinkela_wire_4255),
        .c(_0155_)
    );

    or_bi _1405_ (
        .a(new_Jinkela_wire_1104),
        .b(new_Jinkela_wire_1281),
        .c(_0708_)
    );

    and_ii _2119_ (
        .a(_0155_),
        .b(_0154_),
        .c(_0156_)
    );

    and_bi _1406_ (
        .a(new_Jinkela_wire_1106),
        .b(new_Jinkela_wire_311),
        .c(_0709_)
    );

    and_ii _2120_ (
        .a(new_Jinkela_wire_4974),
        .b(new_Jinkela_wire_2402),
        .c(_0157_)
    );

    and_bi _1407_ (
        .a(_0708_),
        .b(_0709_),
        .c(_0710_)
    );

    and_bb _2121_ (
        .a(new_Jinkela_wire_4975),
        .b(new_Jinkela_wire_2403),
        .c(_0158_)
    );

    and_bi _1408_ (
        .a(new_Jinkela_wire_1037),
        .b(new_Jinkela_wire_1851),
        .c(_0711_)
    );

    and_ii _2122_ (
        .a(_0158_),
        .b(_0157_),
        .c(_0159_)
    );

    or_bb _1409_ (
        .a(_0711_),
        .b(new_Jinkela_wire_4821),
        .c(_0712_)
    );

    inv _2123_ (
        .din(new_Jinkela_wire_5129),
        .dout(new_net_2411)
    );

    and_bi _1410_ (
        .a(_0707_),
        .b(new_Jinkela_wire_5232),
        .c(_0713_)
    );

    and_ii _2124_ (
        .a(new_Jinkela_wire_3174),
        .b(new_Jinkela_wire_4572),
        .c(_0160_)
    );

    and_ii _1411_ (
        .a(_0713_),
        .b(new_Jinkela_wire_4049),
        .c(new_net_8)
    );

    and_bb _2125_ (
        .a(new_Jinkela_wire_3173),
        .b(new_Jinkela_wire_4574),
        .c(_0161_)
    );

    and_bi _1412_ (
        .a(new_Jinkela_wire_341),
        .b(new_Jinkela_wire_6687),
        .c(_0714_)
    );

    or_bb _2126_ (
        .a(_0161_),
        .b(_0160_),
        .c(_0162_)
    );

    and_ii _1413_ (
        .a(new_Jinkela_wire_2406),
        .b(new_Jinkela_wire_6362),
        .c(_0715_)
    );

    or_bb _2127_ (
        .a(new_Jinkela_wire_7524),
        .b(new_Jinkela_wire_3097),
        .c(_0163_)
    );

    and_bi _1414_ (
        .a(new_Jinkela_wire_6094),
        .b(new_Jinkela_wire_5279),
        .c(_0716_)
    );

    and_bb _2128_ (
        .a(new_Jinkela_wire_7525),
        .b(new_Jinkela_wire_3096),
        .c(_0164_)
    );

    and_bi _1415_ (
        .a(new_Jinkela_wire_5280),
        .b(new_Jinkela_wire_6095),
        .c(_0717_)
    );

    and_bi _2129_ (
        .a(_0163_),
        .b(_0164_),
        .c(_0165_)
    );

    or_bb _1416_ (
        .a(_0717_),
        .b(_0716_),
        .c(_0718_)
    );

    and_bb _2130_ (
        .a(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_889),
        .c(_0166_)
    );

    or_bb _1417_ (
        .a(new_Jinkela_wire_1858),
        .b(new_Jinkela_wire_1074),
        .c(_0719_)
    );

    and_bi _2131_ (
        .a(new_Jinkela_wire_1382),
        .b(new_Jinkela_wire_876),
        .c(_0167_)
    );

    or_bb _1418_ (
        .a(new_Jinkela_wire_429),
        .b(new_Jinkela_wire_314),
        .c(_0720_)
    );

    and_ii _2132_ (
        .a(_0167_),
        .b(_0166_),
        .c(_0168_)
    );

    and_bi _1419_ (
        .a(new_Jinkela_wire_427),
        .b(new_Jinkela_wire_208),
        .c(_0721_)
    );

    and_bi _2133_ (
        .a(new_Jinkela_wire_4920),
        .b(new_Jinkela_wire_7892),
        .c(_0169_)
    );

    and_bi _1420_ (
        .a(_0720_),
        .b(_0721_),
        .c(_0722_)
    );

    and_bi _2134_ (
        .a(new_Jinkela_wire_7893),
        .b(new_Jinkela_wire_4919),
        .c(_0170_)
    );

    or_bb _1421_ (
        .a(_0722_),
        .b(new_Jinkela_wire_3586),
        .c(_0723_)
    );

    and_ii _2135_ (
        .a(_0170_),
        .b(_0169_),
        .c(_0171_)
    );

    or_ii _1422_ (
        .a(new_Jinkela_wire_1579),
        .b(new_Jinkela_wire_433),
        .c(_0724_)
    );

    and_bi _2136_ (
        .a(new_Jinkela_wire_6411),
        .b(new_Jinkela_wire_5904),
        .c(_0172_)
    );

    and_bi _1423_ (
        .a(new_Jinkela_wire_1278),
        .b(new_Jinkela_wire_423),
        .c(_0725_)
    );

    and_bi _2137_ (
        .a(new_Jinkela_wire_5905),
        .b(new_Jinkela_wire_6412),
        .c(_0173_)
    );

    and_bi _1424_ (
        .a(_0724_),
        .b(_0725_),
        .c(_0726_)
    );

    or_bb _2138_ (
        .a(_0173_),
        .b(_0172_),
        .c(_0174_)
    );

    and_bi _1425_ (
        .a(new_Jinkela_wire_3584),
        .b(_0726_),
        .c(_0727_)
    );

    and_ii _2139_ (
        .a(new_Jinkela_wire_7085),
        .b(new_Jinkela_wire_4171),
        .c(_0175_)
    );

    and_bi _1426_ (
        .a(_0723_),
        .b(_0727_),
        .c(_0728_)
    );

    and_bi _2140_ (
        .a(new_Jinkela_wire_6849),
        .b(new_Jinkela_wire_1850),
        .c(_0176_)
    );

    and_bi _1427_ (
        .a(new_Jinkela_wire_1045),
        .b(new_Jinkela_wire_4814),
        .c(_0729_)
    );

    and_ii _2141_ (
        .a(new_Jinkela_wire_6364),
        .b(_0175_),
        .c(_0177_)
    );

    or_bb _1428_ (
        .a(_0729_),
        .b(new_Jinkela_wire_4829),
        .c(_0730_)
    );

    and_bi _2142_ (
        .a(new_Jinkela_wire_2404),
        .b(new_Jinkela_wire_2900),
        .c(_0178_)
    );

    and_bi _1429_ (
        .a(_0719_),
        .b(new_Jinkela_wire_5877),
        .c(_0731_)
    );

    and_bi _2143_ (
        .a(new_Jinkela_wire_2902),
        .b(new_Jinkela_wire_2405),
        .c(_0179_)
    );

    and_ii _1430_ (
        .a(_0731_),
        .b(new_Jinkela_wire_5331),
        .c(new_net_10)
    );

    or_bb _2144_ (
        .a(_0179_),
        .b(_0178_),
        .c(_0180_)
    );

    and_bi _1431_ (
        .a(new_Jinkela_wire_70),
        .b(new_Jinkela_wire_6702),
        .c(_0732_)
    );

    and_ii _2145_ (
        .a(new_Jinkela_wire_6122),
        .b(new_Jinkela_wire_4077),
        .c(_0181_)
    );

    or_ii _1432_ (
        .a(new_Jinkela_wire_22),
        .b(new_Jinkela_wire_201),
        .c(_0733_)
    );

    and_bb _2146_ (
        .a(new_Jinkela_wire_6123),
        .b(new_Jinkela_wire_4078),
        .c(_0182_)
    );

    and_bi _1433_ (
        .a(new_Jinkela_wire_539),
        .b(new_Jinkela_wire_11),
        .c(_0734_)
    );

    and_ii _2147_ (
        .a(_0182_),
        .b(_0181_),
        .c(_0183_)
    );

    and_bi _1434_ (
        .a(_0733_),
        .b(new_Jinkela_wire_6754),
        .c(_0735_)
    );

    and_bi _2148_ (
        .a(new_Jinkela_wire_4202),
        .b(new_Jinkela_wire_2090),
        .c(_0184_)
    );

    and_bi _1435_ (
        .a(new_Jinkela_wire_1257),
        .b(new_Jinkela_wire_7079),
        .c(_0736_)
    );

    and_bi _2149_ (
        .a(new_Jinkela_wire_2091),
        .b(new_Jinkela_wire_4203),
        .c(_0185_)
    );

    and_bi _1436_ (
        .a(new_Jinkela_wire_7078),
        .b(new_Jinkela_wire_1258),
        .c(_0737_)
    );

    or_bb _2150_ (
        .a(_0185_),
        .b(_0184_),
        .c(_0186_)
    );

    or_bb _1437_ (
        .a(new_Jinkela_wire_4308),
        .b(new_Jinkela_wire_3610),
        .c(_0738_)
    );

    inv _2151_ (
        .din(new_Jinkela_wire_5421),
        .dout(new_net_2505)
    );

    inv _1438_ (
        .din(new_Jinkela_wire_2845),
        .dout(_0739_)
    );

    or_bb _2152_ (
        .a(new_Jinkela_wire_3030),
        .b(new_Jinkela_wire_2453),
        .c(_0187_)
    );

    inv _1439_ (
        .din(new_Jinkela_wire_765),
        .dout(_0740_)
    );

    and_bb _2153_ (
        .a(new_Jinkela_wire_3031),
        .b(new_Jinkela_wire_2454),
        .c(_0188_)
    );

    or_ii _1440_ (
        .a(new_Jinkela_wire_25),
        .b(new_Jinkela_wire_1318),
        .c(_0741_)
    );

    and_bi _2154_ (
        .a(_0187_),
        .b(_0188_),
        .c(_0189_)
    );

    and_bi _1441_ (
        .a(new_Jinkela_wire_530),
        .b(new_Jinkela_wire_1),
        .c(_0742_)
    );

    and_bi _2155_ (
        .a(new_Jinkela_wire_2930),
        .b(new_Jinkela_wire_2988),
        .c(_0190_)
    );

    or_bi _1442_ (
        .a(new_Jinkela_wire_6707),
        .b(new_Jinkela_wire_4603),
        .c(_0743_)
    );

    and_bi _2156_ (
        .a(new_Jinkela_wire_2986),
        .b(new_Jinkela_wire_2929),
        .c(_0191_)
    );

    and_bi _1443_ (
        .a(new_Jinkela_wire_5704),
        .b(_0743_),
        .c(_0744_)
    );

    and_ii _2157_ (
        .a(_0191_),
        .b(_0190_),
        .c(_0192_)
    );

    and_bi _1444_ (
        .a(new_Jinkela_wire_4604),
        .b(new_Jinkela_wire_6708),
        .c(_0745_)
    );

    or_bi _2158_ (
        .a(new_Jinkela_wire_3678),
        .b(new_Jinkela_wire_2154),
        .c(_0193_)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1905),
        .dout(new_Jinkela_wire_1906)
    );

    bfr new_Jinkela_buffer_4211 (
        .din(new_Jinkela_wire_5795),
        .dout(new_Jinkela_wire_5796)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1872),
        .dout(new_Jinkela_wire_1873)
    );

    bfr new_Jinkela_buffer_4181 (
        .din(new_Jinkela_wire_5754),
        .dout(new_Jinkela_wire_5755)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(_0244_),
        .dout(new_Jinkela_wire_1946)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1893),
        .dout(new_Jinkela_wire_1894)
    );

    bfr new_Jinkela_buffer_4217 (
        .din(new_Jinkela_wire_5816),
        .dout(new_Jinkela_wire_5817)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1873),
        .dout(new_Jinkela_wire_1874)
    );

    bfr new_Jinkela_buffer_4182 (
        .din(new_Jinkela_wire_5755),
        .dout(new_Jinkela_wire_5756)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1887),
        .dout(new_Jinkela_wire_1888)
    );

    bfr new_Jinkela_buffer_4224 (
        .din(new_Jinkela_wire_5827),
        .dout(new_Jinkela_wire_5828)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1874),
        .dout(new_Jinkela_wire_1875)
    );

    bfr new_Jinkela_buffer_4183 (
        .din(new_Jinkela_wire_5756),
        .dout(new_Jinkela_wire_5757)
    );

    bfr new_Jinkela_buffer_4216 (
        .din(new_Jinkela_wire_5815),
        .dout(new_Jinkela_wire_5816)
    );

    bfr new_Jinkela_buffer_4212 (
        .din(new_Jinkela_wire_5796),
        .dout(new_Jinkela_wire_5797)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1875),
        .dout(new_Jinkela_wire_1876)
    );

    bfr new_Jinkela_buffer_4184 (
        .din(new_Jinkela_wire_5757),
        .dout(new_Jinkela_wire_5758)
    );

    spl3L new_Jinkela_splitter_332 (
        .a(new_Jinkela_wire_1906),
        .d(new_Jinkela_wire_1907),
        .b(new_Jinkela_wire_1908),
        .c(new_Jinkela_wire_1909)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1894),
        .dout(new_Jinkela_wire_1895)
    );

    spl2 new_Jinkela_splitter_327 (
        .a(new_Jinkela_wire_1876),
        .b(new_Jinkela_wire_1877),
        .c(new_Jinkela_wire_1878)
    );

    bfr new_Jinkela_buffer_4185 (
        .din(new_Jinkela_wire_5758),
        .dout(new_Jinkela_wire_5759)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1915),
        .dout(new_Jinkela_wire_1916)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1895),
        .dout(new_Jinkela_wire_1896)
    );

    bfr new_Jinkela_buffer_4213 (
        .din(new_Jinkela_wire_5797),
        .dout(new_Jinkela_wire_5798)
    );

    bfr new_Jinkela_buffer_4186 (
        .din(new_Jinkela_wire_5759),
        .dout(new_Jinkela_wire_5760)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(new_Jinkela_wire_1948),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_4187 (
        .din(new_Jinkela_wire_5760),
        .dout(new_Jinkela_wire_5761)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1896),
        .dout(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_4214 (
        .din(new_Jinkela_wire_5798),
        .dout(new_Jinkela_wire_5799)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(new_Jinkela_wire_1916),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_4188 (
        .din(new_Jinkela_wire_5761),
        .dout(new_Jinkela_wire_5762)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1897),
        .dout(new_Jinkela_wire_1898)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1909),
        .dout(new_Jinkela_wire_1910)
    );

    bfr new_Jinkela_buffer_4189 (
        .din(new_Jinkela_wire_5762),
        .dout(new_Jinkela_wire_5763)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1898),
        .dout(new_Jinkela_wire_1899)
    );

    bfr new_Jinkela_buffer_4254 (
        .din(new_net_2409),
        .dout(new_Jinkela_wire_5858)
    );

    spl2 new_Jinkela_splitter_608 (
        .a(new_Jinkela_wire_5799),
        .b(new_Jinkela_wire_5800),
        .c(new_Jinkela_wire_5801)
    );

    bfr new_Jinkela_buffer_4190 (
        .din(new_Jinkela_wire_5763),
        .dout(new_Jinkela_wire_5764)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1899),
        .dout(new_Jinkela_wire_1900)
    );

    spl2 new_Jinkela_splitter_333 (
        .a(new_Jinkela_wire_1910),
        .b(new_Jinkela_wire_1911),
        .c(new_Jinkela_wire_1912)
    );

    bfr new_Jinkela_buffer_4218 (
        .din(new_Jinkela_wire_5819),
        .dout(new_Jinkela_wire_5820)
    );

    bfr new_Jinkela_buffer_4191 (
        .din(new_Jinkela_wire_5764),
        .dout(new_Jinkela_wire_5765)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(new_Jinkela_wire_1912),
        .dout(new_Jinkela_wire_1913)
    );

    spl2 new_Jinkela_splitter_613 (
        .a(new_Jinkela_wire_5817),
        .b(new_Jinkela_wire_5818),
        .c(new_Jinkela_wire_5819)
    );

    bfr new_Jinkela_buffer_4192 (
        .din(new_Jinkela_wire_5765),
        .dout(new_Jinkela_wire_5766)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    spl3L new_Jinkela_splitter_337 (
        .a(_0678_),
        .d(new_Jinkela_wire_1952),
        .b(new_Jinkela_wire_1953),
        .c(new_Jinkela_wire_1954)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1917),
        .dout(new_Jinkela_wire_1918)
    );

    bfr new_Jinkela_buffer_4193 (
        .din(new_Jinkela_wire_5766),
        .dout(new_Jinkela_wire_5767)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    spl2 new_Jinkela_splitter_615 (
        .a(_0641_),
        .b(new_Jinkela_wire_5864),
        .c(new_Jinkela_wire_5865)
    );

    bfr new_Jinkela_buffer_4260 (
        .din(_0546_),
        .dout(new_Jinkela_wire_5866)
    );

    bfr new_Jinkela_buffer_4194 (
        .din(new_Jinkela_wire_5767),
        .dout(new_Jinkela_wire_5768)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1913),
        .dout(new_Jinkela_wire_1914)
    );

    bfr new_Jinkela_buffer_4225 (
        .din(new_Jinkela_wire_5828),
        .dout(new_Jinkela_wire_5829)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(_0739_),
        .dout(new_Jinkela_wire_1955)
    );

    bfr new_Jinkela_buffer_4219 (
        .din(new_Jinkela_wire_5820),
        .dout(new_Jinkela_wire_5821)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1918),
        .dout(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_4195 (
        .din(new_Jinkela_wire_5768),
        .dout(new_Jinkela_wire_5769)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(_0677_),
        .dout(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1919),
        .dout(new_Jinkela_wire_1920)
    );

    bfr new_Jinkela_buffer_4196 (
        .din(new_Jinkela_wire_5769),
        .dout(new_Jinkela_wire_5770)
    );

    bfr new_Jinkela_buffer_4255 (
        .din(new_Jinkela_wire_5858),
        .dout(new_Jinkela_wire_5859)
    );

    spl2 new_Jinkela_splitter_335 (
        .a(new_Jinkela_wire_1946),
        .b(new_Jinkela_wire_1947),
        .c(new_Jinkela_wire_1948)
    );

    bfr new_Jinkela_buffer_4220 (
        .din(new_Jinkela_wire_5821),
        .dout(new_Jinkela_wire_5822)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1920),
        .dout(new_Jinkela_wire_1921)
    );

    bfr new_Jinkela_buffer_4197 (
        .din(new_Jinkela_wire_5770),
        .dout(new_Jinkela_wire_5771)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1955),
        .dout(new_Jinkela_wire_1956)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1921),
        .dout(new_Jinkela_wire_1922)
    );

    bfr new_Jinkela_buffer_4198 (
        .din(new_Jinkela_wire_5771),
        .dout(new_Jinkela_wire_5772)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(_0367_),
        .dout(new_Jinkela_wire_1967)
    );

    bfr new_Jinkela_buffer_4226 (
        .din(new_Jinkela_wire_5829),
        .dout(new_Jinkela_wire_5830)
    );

    bfr new_Jinkela_buffer_4221 (
        .din(new_Jinkela_wire_5822),
        .dout(new_Jinkela_wire_5823)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1922),
        .dout(new_Jinkela_wire_1923)
    );

    spl2 new_Jinkela_splitter_336 (
        .a(new_Jinkela_wire_1949),
        .b(new_Jinkela_wire_1950),
        .c(new_Jinkela_wire_1951)
    );

    bfr new_Jinkela_buffer_4222 (
        .din(new_Jinkela_wire_5823),
        .dout(new_Jinkela_wire_5824)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1923),
        .dout(new_Jinkela_wire_1924)
    );

    bfr new_Jinkela_buffer_4227 (
        .din(new_Jinkela_wire_5830),
        .dout(new_Jinkela_wire_5831)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1924),
        .dout(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_4256 (
        .din(new_Jinkela_wire_5859),
        .dout(new_Jinkela_wire_5860)
    );

    bfr new_Jinkela_buffer_5831 (
        .din(_0834_),
        .dout(new_Jinkela_wire_7826)
    );

    bfr new_Jinkela_buffer_5746 (
        .din(new_Jinkela_wire_7728),
        .dout(new_Jinkela_wire_7729)
    );

    and_ii _1295_ (
        .a(new_Jinkela_wire_1364),
        .b(new_Jinkela_wire_47),
        .c(_0602_)
    );

    bfr new_Jinkela_buffer_5764 (
        .din(new_Jinkela_wire_7748),
        .dout(new_Jinkela_wire_7749)
    );

    bfr new_Jinkela_buffer_5747 (
        .din(new_Jinkela_wire_7729),
        .dout(new_Jinkela_wire_7730)
    );

    bfr new_Jinkela_buffer_5800 (
        .din(new_Jinkela_wire_7792),
        .dout(new_Jinkela_wire_7793)
    );

    bfr new_Jinkela_buffer_5748 (
        .din(new_Jinkela_wire_7730),
        .dout(new_Jinkela_wire_7731)
    );

    spl2 new_Jinkela_splitter_774 (
        .a(_1004_),
        .b(new_Jinkela_wire_7848),
        .c(new_Jinkela_wire_7849)
    );

    bfr new_Jinkela_buffer_5765 (
        .din(new_Jinkela_wire_7749),
        .dout(new_Jinkela_wire_7750)
    );

    bfr new_Jinkela_buffer_5749 (
        .din(new_Jinkela_wire_7731),
        .dout(new_Jinkela_wire_7732)
    );

    bfr new_Jinkela_buffer_5832 (
        .din(new_Jinkela_wire_7826),
        .dout(new_Jinkela_wire_7827)
    );

    spl4L new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_400),
        .d(new_Jinkela_wire_401),
        .e(new_Jinkela_wire_402),
        .b(new_Jinkela_wire_403),
        .c(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_5750 (
        .din(new_Jinkela_wire_7732),
        .dout(new_Jinkela_wire_7733)
    );

    bfr new_Jinkela_buffer_5766 (
        .din(new_Jinkela_wire_7750),
        .dout(new_Jinkela_wire_7751)
    );

    bfr new_Jinkela_buffer_5751 (
        .din(new_Jinkela_wire_7733),
        .dout(new_Jinkela_wire_7734)
    );

    bfr new_Jinkela_buffer_5752 (
        .din(new_Jinkela_wire_7734),
        .dout(new_Jinkela_wire_7735)
    );

    spl2 new_Jinkela_splitter_773 (
        .a(_0758_),
        .b(new_Jinkela_wire_7840),
        .c(new_Jinkela_wire_7841)
    );

    bfr new_Jinkela_buffer_5767 (
        .din(new_Jinkela_wire_7751),
        .dout(new_Jinkela_wire_7752)
    );

    bfr new_Jinkela_buffer_5753 (
        .din(new_Jinkela_wire_7735),
        .dout(new_Jinkela_wire_7736)
    );

    bfr new_Jinkela_buffer_5801 (
        .din(new_Jinkela_wire_7793),
        .dout(new_Jinkela_wire_7794)
    );

    bfr new_Jinkela_buffer_5754 (
        .din(new_Jinkela_wire_7736),
        .dout(new_Jinkela_wire_7737)
    );

    bfr new_Jinkela_buffer_5768 (
        .din(new_Jinkela_wire_7752),
        .dout(new_Jinkela_wire_7753)
    );

    bfr new_Jinkela_buffer_5755 (
        .din(new_Jinkela_wire_7737),
        .dout(new_Jinkela_wire_7738)
    );

    bfr new_Jinkela_buffer_5756 (
        .din(new_Jinkela_wire_7738),
        .dout(new_Jinkela_wire_7739)
    );

    bfr new_Jinkela_buffer_5845 (
        .din(new_Jinkela_wire_7841),
        .dout(new_Jinkela_wire_7842)
    );

    bfr new_Jinkela_buffer_5769 (
        .din(new_Jinkela_wire_7753),
        .dout(new_Jinkela_wire_7754)
    );

    bfr new_Jinkela_buffer_5757 (
        .din(new_Jinkela_wire_7739),
        .dout(new_Jinkela_wire_7740)
    );

    bfr new_Jinkela_buffer_5802 (
        .din(new_Jinkela_wire_7794),
        .dout(new_Jinkela_wire_7795)
    );

    bfr new_Jinkela_buffer_5770 (
        .din(new_Jinkela_wire_7754),
        .dout(new_Jinkela_wire_7755)
    );

    bfr new_Jinkela_buffer_5833 (
        .din(new_Jinkela_wire_7827),
        .dout(new_Jinkela_wire_7828)
    );

    bfr new_Jinkela_buffer_5771 (
        .din(new_Jinkela_wire_7755),
        .dout(new_Jinkela_wire_7756)
    );

    bfr new_Jinkela_buffer_5803 (
        .din(new_Jinkela_wire_7795),
        .dout(new_Jinkela_wire_7796)
    );

    bfr new_Jinkela_buffer_5772 (
        .din(new_Jinkela_wire_7756),
        .dout(new_Jinkela_wire_7757)
    );

    bfr new_Jinkela_buffer_5773 (
        .din(new_Jinkela_wire_7757),
        .dout(new_Jinkela_wire_7758)
    );

    bfr new_Jinkela_buffer_5804 (
        .din(new_Jinkela_wire_7796),
        .dout(new_Jinkela_wire_7797)
    );

    bfr new_Jinkela_buffer_5774 (
        .din(new_Jinkela_wire_7758),
        .dout(new_Jinkela_wire_7759)
    );

    bfr new_Jinkela_buffer_5851 (
        .din(_0415_),
        .dout(new_Jinkela_wire_7850)
    );

    bfr new_Jinkela_buffer_5834 (
        .din(new_Jinkela_wire_7828),
        .dout(new_Jinkela_wire_7829)
    );

    bfr new_Jinkela_buffer_5775 (
        .din(new_Jinkela_wire_7759),
        .dout(new_Jinkela_wire_7760)
    );

    bfr new_Jinkela_buffer_5805 (
        .din(new_Jinkela_wire_7797),
        .dout(new_Jinkela_wire_7798)
    );

    bfr new_Jinkela_buffer_5776 (
        .din(new_Jinkela_wire_7760),
        .dout(new_Jinkela_wire_7761)
    );

    bfr new_Jinkela_buffer_5777 (
        .din(new_Jinkela_wire_7761),
        .dout(new_Jinkela_wire_7762)
    );

    bfr new_Jinkela_buffer_5806 (
        .din(new_Jinkela_wire_7798),
        .dout(new_Jinkela_wire_7799)
    );

    bfr new_Jinkela_buffer_5778 (
        .din(new_Jinkela_wire_7762),
        .dout(new_Jinkela_wire_7763)
    );

    bfr new_Jinkela_buffer_1965 (
        .din(new_Jinkela_wire_3044),
        .dout(new_Jinkela_wire_3045)
    );

    bfr new_Jinkela_buffer_4164 (
        .din(new_Jinkela_wire_5737),
        .dout(new_Jinkela_wire_5738)
    );

    bfr new_Jinkela_buffer_1941 (
        .din(new_Jinkela_wire_3016),
        .dout(new_Jinkela_wire_3017)
    );

    bfr new_Jinkela_buffer_4149 (
        .din(new_Jinkela_wire_5720),
        .dout(new_Jinkela_wire_5721)
    );

    bfr new_Jinkela_buffer_4200 (
        .din(new_Jinkela_wire_5779),
        .dout(new_Jinkela_wire_5780)
    );

    spl2 new_Jinkela_splitter_407 (
        .a(new_Jinkela_wire_3086),
        .b(new_Jinkela_wire_3087),
        .c(new_Jinkela_wire_3088)
    );

    bfr new_Jinkela_buffer_1942 (
        .din(new_Jinkela_wire_3017),
        .dout(new_Jinkela_wire_3018)
    );

    bfr new_Jinkela_buffer_4150 (
        .din(new_Jinkela_wire_5721),
        .dout(new_Jinkela_wire_5722)
    );

    bfr new_Jinkela_buffer_1966 (
        .din(new_Jinkela_wire_3045),
        .dout(new_Jinkela_wire_3046)
    );

    bfr new_Jinkela_buffer_4165 (
        .din(new_Jinkela_wire_5738),
        .dout(new_Jinkela_wire_5739)
    );

    bfr new_Jinkela_buffer_1943 (
        .din(new_Jinkela_wire_3018),
        .dout(new_Jinkela_wire_3019)
    );

    bfr new_Jinkela_buffer_4151 (
        .din(new_Jinkela_wire_5722),
        .dout(new_Jinkela_wire_5723)
    );

    spl2 new_Jinkela_splitter_614 (
        .a(_0929_),
        .b(new_Jinkela_wire_5825),
        .c(new_Jinkela_wire_5826)
    );

    bfr new_Jinkela_buffer_1985 (
        .din(new_Jinkela_wire_3071),
        .dout(new_Jinkela_wire_3072)
    );

    bfr new_Jinkela_buffer_4208 (
        .din(new_Jinkela_wire_5790),
        .dout(new_Jinkela_wire_5791)
    );

    bfr new_Jinkela_buffer_1944 (
        .din(new_Jinkela_wire_3019),
        .dout(new_Jinkela_wire_3020)
    );

    bfr new_Jinkela_buffer_4152 (
        .din(new_Jinkela_wire_5723),
        .dout(new_Jinkela_wire_5724)
    );

    bfr new_Jinkela_buffer_1967 (
        .din(new_Jinkela_wire_3046),
        .dout(new_Jinkela_wire_3047)
    );

    bfr new_Jinkela_buffer_4166 (
        .din(new_Jinkela_wire_5739),
        .dout(new_Jinkela_wire_5740)
    );

    bfr new_Jinkela_buffer_1945 (
        .din(new_Jinkela_wire_3020),
        .dout(new_Jinkela_wire_3021)
    );

    bfr new_Jinkela_buffer_4153 (
        .din(new_Jinkela_wire_5724),
        .dout(new_Jinkela_wire_5725)
    );

    bfr new_Jinkela_buffer_1999 (
        .din(new_Jinkela_wire_3092),
        .dout(new_Jinkela_wire_3093)
    );

    bfr new_Jinkela_buffer_1946 (
        .din(new_Jinkela_wire_3021),
        .dout(new_Jinkela_wire_3022)
    );

    bfr new_Jinkela_buffer_4154 (
        .din(new_Jinkela_wire_5725),
        .dout(new_Jinkela_wire_5726)
    );

    bfr new_Jinkela_buffer_1968 (
        .din(new_Jinkela_wire_3047),
        .dout(new_Jinkela_wire_3048)
    );

    bfr new_Jinkela_buffer_4167 (
        .din(new_Jinkela_wire_5740),
        .dout(new_Jinkela_wire_5741)
    );

    bfr new_Jinkela_buffer_1947 (
        .din(new_Jinkela_wire_3022),
        .dout(new_Jinkela_wire_3023)
    );

    bfr new_Jinkela_buffer_4155 (
        .din(new_Jinkela_wire_5726),
        .dout(new_Jinkela_wire_5727)
    );

    bfr new_Jinkela_buffer_4201 (
        .din(new_Jinkela_wire_5780),
        .dout(new_Jinkela_wire_5781)
    );

    bfr new_Jinkela_buffer_1986 (
        .din(new_Jinkela_wire_3072),
        .dout(new_Jinkela_wire_3073)
    );

    bfr new_Jinkela_buffer_1948 (
        .din(new_Jinkela_wire_3023),
        .dout(new_Jinkela_wire_3024)
    );

    bfr new_Jinkela_buffer_4156 (
        .din(new_Jinkela_wire_5727),
        .dout(new_Jinkela_wire_5728)
    );

    bfr new_Jinkela_buffer_1969 (
        .din(new_Jinkela_wire_3048),
        .dout(new_Jinkela_wire_3049)
    );

    bfr new_Jinkela_buffer_4168 (
        .din(new_Jinkela_wire_5741),
        .dout(new_Jinkela_wire_5742)
    );

    bfr new_Jinkela_buffer_1949 (
        .din(new_Jinkela_wire_3024),
        .dout(new_Jinkela_wire_3025)
    );

    bfr new_Jinkela_buffer_4157 (
        .din(new_Jinkela_wire_5728),
        .dout(new_Jinkela_wire_5729)
    );

    spl4L new_Jinkela_splitter_611 (
        .a(new_Jinkela_wire_5805),
        .d(new_Jinkela_wire_5806),
        .e(new_Jinkela_wire_5807),
        .b(new_Jinkela_wire_5808),
        .c(new_Jinkela_wire_5809)
    );

    bfr new_Jinkela_buffer_1950 (
        .din(new_Jinkela_wire_3025),
        .dout(new_Jinkela_wire_3026)
    );

    bfr new_Jinkela_buffer_4169 (
        .din(new_Jinkela_wire_5742),
        .dout(new_Jinkela_wire_5743)
    );

    bfr new_Jinkela_buffer_1970 (
        .din(new_Jinkela_wire_3049),
        .dout(new_Jinkela_wire_3050)
    );

    bfr new_Jinkela_buffer_4202 (
        .din(new_Jinkela_wire_5781),
        .dout(new_Jinkela_wire_5782)
    );

    bfr new_Jinkela_buffer_1951 (
        .din(new_Jinkela_wire_3026),
        .dout(new_Jinkela_wire_3027)
    );

    bfr new_Jinkela_buffer_4170 (
        .din(new_Jinkela_wire_5743),
        .dout(new_Jinkela_wire_5744)
    );

    bfr new_Jinkela_buffer_2000 (
        .din(new_Jinkela_wire_3098),
        .dout(new_Jinkela_wire_3099)
    );

    bfr new_Jinkela_buffer_4223 (
        .din(_0490_),
        .dout(new_Jinkela_wire_5827)
    );

    bfr new_Jinkela_buffer_1987 (
        .din(new_Jinkela_wire_3073),
        .dout(new_Jinkela_wire_3074)
    );

    bfr new_Jinkela_buffer_4209 (
        .din(new_Jinkela_wire_5791),
        .dout(new_Jinkela_wire_5792)
    );

    bfr new_Jinkela_buffer_1971 (
        .din(new_Jinkela_wire_3050),
        .dout(new_Jinkela_wire_3051)
    );

    bfr new_Jinkela_buffer_4171 (
        .din(new_Jinkela_wire_5744),
        .dout(new_Jinkela_wire_5745)
    );

    bfr new_Jinkela_buffer_4203 (
        .din(new_Jinkela_wire_5782),
        .dout(new_Jinkela_wire_5783)
    );

    bfr new_Jinkela_buffer_1972 (
        .din(new_Jinkela_wire_3051),
        .dout(new_Jinkela_wire_3052)
    );

    bfr new_Jinkela_buffer_4172 (
        .din(new_Jinkela_wire_5745),
        .dout(new_Jinkela_wire_5746)
    );

    bfr new_Jinkela_buffer_2004 (
        .din(_0455_),
        .dout(new_Jinkela_wire_3105)
    );

    bfr new_Jinkela_buffer_1988 (
        .din(new_Jinkela_wire_3074),
        .dout(new_Jinkela_wire_3075)
    );

    bfr new_Jinkela_buffer_1973 (
        .din(new_Jinkela_wire_3052),
        .dout(new_Jinkela_wire_3053)
    );

    bfr new_Jinkela_buffer_4173 (
        .din(new_Jinkela_wire_5746),
        .dout(new_Jinkela_wire_5747)
    );

    bfr new_Jinkela_buffer_4204 (
        .din(new_Jinkela_wire_5783),
        .dout(new_Jinkela_wire_5784)
    );

    bfr new_Jinkela_buffer_2005 (
        .din(new_Jinkela_wire_3105),
        .dout(new_Jinkela_wire_3106)
    );

    bfr new_Jinkela_buffer_1974 (
        .din(new_Jinkela_wire_3053),
        .dout(new_Jinkela_wire_3054)
    );

    bfr new_Jinkela_buffer_4174 (
        .din(new_Jinkela_wire_5747),
        .dout(new_Jinkela_wire_5748)
    );

    spl2 new_Jinkela_splitter_610 (
        .a(new_Jinkela_wire_5802),
        .b(new_Jinkela_wire_5803),
        .c(new_Jinkela_wire_5804)
    );

    bfr new_Jinkela_buffer_1989 (
        .din(new_Jinkela_wire_3075),
        .dout(new_Jinkela_wire_3076)
    );

    bfr new_Jinkela_buffer_4210 (
        .din(new_Jinkela_wire_5792),
        .dout(new_Jinkela_wire_5793)
    );

    bfr new_Jinkela_buffer_1975 (
        .din(new_Jinkela_wire_3054),
        .dout(new_Jinkela_wire_3055)
    );

    bfr new_Jinkela_buffer_4175 (
        .din(new_Jinkela_wire_5748),
        .dout(new_Jinkela_wire_5749)
    );

    bfr new_Jinkela_buffer_4205 (
        .din(new_Jinkela_wire_5784),
        .dout(new_Jinkela_wire_5785)
    );

    bfr new_Jinkela_buffer_1976 (
        .din(new_Jinkela_wire_3055),
        .dout(new_Jinkela_wire_3056)
    );

    bfr new_Jinkela_buffer_4176 (
        .din(new_Jinkela_wire_5749),
        .dout(new_Jinkela_wire_5750)
    );

    bfr new_Jinkela_buffer_2035 (
        .din(_0363_),
        .dout(new_Jinkela_wire_3136)
    );

    bfr new_Jinkela_buffer_1990 (
        .din(new_Jinkela_wire_3076),
        .dout(new_Jinkela_wire_3077)
    );

    spl4L new_Jinkela_splitter_612 (
        .a(new_Jinkela_wire_5810),
        .d(new_Jinkela_wire_5811),
        .e(new_Jinkela_wire_5812),
        .b(new_Jinkela_wire_5813),
        .c(new_Jinkela_wire_5814)
    );

    bfr new_Jinkela_buffer_1977 (
        .din(new_Jinkela_wire_3056),
        .dout(new_Jinkela_wire_3057)
    );

    bfr new_Jinkela_buffer_4177 (
        .din(new_Jinkela_wire_5750),
        .dout(new_Jinkela_wire_5751)
    );

    bfr new_Jinkela_buffer_4206 (
        .din(new_Jinkela_wire_5785),
        .dout(new_Jinkela_wire_5786)
    );

    bfr new_Jinkela_buffer_1978 (
        .din(new_Jinkela_wire_3057),
        .dout(new_Jinkela_wire_3058)
    );

    bfr new_Jinkela_buffer_4178 (
        .din(new_Jinkela_wire_5751),
        .dout(new_Jinkela_wire_5752)
    );

    bfr new_Jinkela_buffer_2001 (
        .din(new_Jinkela_wire_3099),
        .dout(new_Jinkela_wire_3100)
    );

    bfr new_Jinkela_buffer_1991 (
        .din(new_Jinkela_wire_3077),
        .dout(new_Jinkela_wire_3078)
    );

    spl2 new_Jinkela_splitter_607 (
        .a(new_Jinkela_wire_5793),
        .b(new_Jinkela_wire_5794),
        .c(new_Jinkela_wire_5795)
    );

    bfr new_Jinkela_buffer_1979 (
        .din(new_Jinkela_wire_3058),
        .dout(new_Jinkela_wire_3059)
    );

    bfr new_Jinkela_buffer_4179 (
        .din(new_Jinkela_wire_5752),
        .dout(new_Jinkela_wire_5753)
    );

    bfr new_Jinkela_buffer_4207 (
        .din(new_Jinkela_wire_5786),
        .dout(new_Jinkela_wire_5787)
    );

    bfr new_Jinkela_buffer_1980 (
        .din(new_Jinkela_wire_3059),
        .dout(new_Jinkela_wire_3060)
    );

    bfr new_Jinkela_buffer_4180 (
        .din(new_Jinkela_wire_5753),
        .dout(new_Jinkela_wire_5754)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_Jinkela_wire_1925),
        .dout(new_Jinkela_wire_1926)
    );

    spl2 new_Jinkela_splitter_340 (
        .a(_0067_),
        .b(new_Jinkela_wire_1969),
        .c(new_Jinkela_wire_1970)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1956),
        .dout(new_Jinkela_wire_1957)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1926),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1964),
        .dout(new_Jinkela_wire_1965)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(_0138_),
        .dout(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1928),
        .dout(new_Jinkela_wire_1929)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1929),
        .dout(new_Jinkela_wire_1930)
    );

    spl3L new_Jinkela_splitter_338 (
        .a(new_Jinkela_wire_1958),
        .d(new_Jinkela_wire_1959),
        .b(new_Jinkela_wire_1960),
        .c(new_Jinkela_wire_1961)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1930),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1967),
        .dout(new_Jinkela_wire_1968)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1931),
        .dout(new_Jinkela_wire_1932)
    );

    spl2 new_Jinkela_splitter_339 (
        .a(new_Jinkela_wire_1961),
        .b(new_Jinkela_wire_1962),
        .c(new_Jinkela_wire_1963)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1932),
        .dout(new_Jinkela_wire_1933)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(_1122_),
        .dout(new_Jinkela_wire_1974)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1933),
        .dout(new_Jinkela_wire_1934)
    );

    spl2 new_Jinkela_splitter_341 (
        .a(new_Jinkela_wire_1971),
        .b(new_Jinkela_wire_1972),
        .c(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1934),
        .dout(new_Jinkela_wire_1935)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(_0089_),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1935),
        .dout(new_Jinkela_wire_1936)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1936),
        .dout(new_Jinkela_wire_1937)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(new_Jinkela_wire_1975),
        .dout(new_Jinkela_wire_1976)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1937),
        .dout(new_Jinkela_wire_1938)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(_0514_),
        .dout(new_Jinkela_wire_1978)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1938),
        .dout(new_Jinkela_wire_1939)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(_0375_),
        .dout(new_Jinkela_wire_1980)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1939),
        .dout(new_Jinkela_wire_1940)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1976),
        .dout(new_Jinkela_wire_1977)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1940),
        .dout(new_Jinkela_wire_1941)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1978),
        .dout(new_Jinkela_wire_1979)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(new_Jinkela_wire_1941),
        .dout(new_Jinkela_wire_1942)
    );

    spl2 new_Jinkela_splitter_342 (
        .a(_1070_),
        .b(new_Jinkela_wire_1983),
        .c(new_Jinkela_wire_1984)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(_0217_),
        .dout(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1942),
        .dout(new_Jinkela_wire_1943)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1980),
        .dout(new_Jinkela_wire_1981)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_net_2445),
        .dout(new_Jinkela_wire_1989)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1981),
        .dout(new_Jinkela_wire_1982)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(_0573_),
        .dout(new_Jinkela_wire_1986)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1986),
        .dout(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_700 (
        .din(G27),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_5835 (
        .din(new_Jinkela_wire_7829),
        .dout(new_Jinkela_wire_7830)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_1404),
        .dout(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_5779 (
        .din(new_Jinkela_wire_7763),
        .dout(new_Jinkela_wire_7764)
    );

    bfr new_Jinkela_buffer_5807 (
        .din(new_Jinkela_wire_7799),
        .dout(new_Jinkela_wire_7800)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_1405),
        .dout(new_Jinkela_wire_1406)
    );

    bfr new_Jinkela_buffer_5780 (
        .din(new_Jinkela_wire_7764),
        .dout(new_Jinkela_wire_7765)
    );

    spl3L new_Jinkela_splitter_775 (
        .a(_0268_),
        .d(new_Jinkela_wire_7867),
        .b(new_Jinkela_wire_7870),
        .c(new_Jinkela_wire_7875)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_1406),
        .dout(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_5781 (
        .din(new_Jinkela_wire_7765),
        .dout(new_Jinkela_wire_7766)
    );

    bfr new_Jinkela_buffer_5808 (
        .din(new_Jinkela_wire_7800),
        .dout(new_Jinkela_wire_7801)
    );

    spl4L new_Jinkela_splitter_264 (
        .a(G173),
        .d(new_Jinkela_wire_1438),
        .e(new_Jinkela_wire_1439),
        .b(new_Jinkela_wire_1440),
        .c(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_1407),
        .dout(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_5782 (
        .din(new_Jinkela_wire_7766),
        .dout(new_Jinkela_wire_7767)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_1484),
        .dout(new_Jinkela_wire_1485)
    );

    bfr new_Jinkela_buffer_5846 (
        .din(new_Jinkela_wire_7842),
        .dout(new_Jinkela_wire_7843)
    );

    bfr new_Jinkela_buffer_734 (
        .din(G60),
        .dout(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_5836 (
        .din(new_Jinkela_wire_7830),
        .dout(new_Jinkela_wire_7831)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_5783 (
        .din(new_Jinkela_wire_7767),
        .dout(new_Jinkela_wire_7768)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_5809 (
        .din(new_Jinkela_wire_7801),
        .dout(new_Jinkela_wire_7802)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_5784 (
        .din(new_Jinkela_wire_7768),
        .dout(new_Jinkela_wire_7769)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_1410),
        .dout(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_5785 (
        .din(new_Jinkela_wire_7769),
        .dout(new_Jinkela_wire_7770)
    );

    bfr new_Jinkela_buffer_5810 (
        .din(new_Jinkela_wire_7802),
        .dout(new_Jinkela_wire_7803)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_1411),
        .dout(new_Jinkela_wire_1412)
    );

    bfr new_Jinkela_buffer_5786 (
        .din(new_Jinkela_wire_7770),
        .dout(new_Jinkela_wire_7771)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_5837 (
        .din(new_Jinkela_wire_7831),
        .dout(new_Jinkela_wire_7832)
    );

    spl3L new_Jinkela_splitter_259 (
        .a(new_Jinkela_wire_1412),
        .d(new_Jinkela_wire_1413),
        .b(new_Jinkela_wire_1414),
        .c(new_Jinkela_wire_1415)
    );

    bfr new_Jinkela_buffer_5787 (
        .din(new_Jinkela_wire_7771),
        .dout(new_Jinkela_wire_7772)
    );

    bfr new_Jinkela_buffer_5811 (
        .din(new_Jinkela_wire_7803),
        .dout(new_Jinkela_wire_7804)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_5788 (
        .din(new_Jinkela_wire_7772),
        .dout(new_Jinkela_wire_7773)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(new_Jinkela_wire_1435),
        .b(new_Jinkela_wire_1436),
        .c(new_Jinkela_wire_1437)
    );

    bfr new_Jinkela_buffer_5852 (
        .din(new_net_2369),
        .dout(new_Jinkela_wire_7851)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    bfr new_Jinkela_buffer_5789 (
        .din(new_Jinkela_wire_7773),
        .dout(new_Jinkela_wire_7774)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_5812 (
        .din(new_Jinkela_wire_7804),
        .dout(new_Jinkela_wire_7805)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    bfr new_Jinkela_buffer_5790 (
        .din(new_Jinkela_wire_7774),
        .dout(new_Jinkela_wire_7775)
    );

    bfr new_Jinkela_buffer_742 (
        .din(G21),
        .dout(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_5847 (
        .din(new_Jinkela_wire_7843),
        .dout(new_Jinkela_wire_7844)
    );

    spl2 new_Jinkela_splitter_273 (
        .a(G170),
        .b(new_Jinkela_wire_1507),
        .c(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_5838 (
        .din(new_Jinkela_wire_7832),
        .dout(new_Jinkela_wire_7833)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(new_Jinkela_wire_1418),
        .b(new_Jinkela_wire_1419),
        .c(new_Jinkela_wire_1420)
    );

    bfr new_Jinkela_buffer_5791 (
        .din(new_Jinkela_wire_7775),
        .dout(new_Jinkela_wire_7776)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_5813 (
        .din(new_Jinkela_wire_7805),
        .dout(new_Jinkela_wire_7806)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_1485),
        .dout(new_Jinkela_wire_1486)
    );

    bfr new_Jinkela_buffer_5792 (
        .din(new_Jinkela_wire_7776),
        .dout(new_Jinkela_wire_7777)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_1442),
        .dout(new_Jinkela_wire_1443)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(new_Jinkela_wire_1421),
        .b(new_Jinkela_wire_1422),
        .c(new_Jinkela_wire_1423)
    );

    bfr new_Jinkela_buffer_5793 (
        .din(new_Jinkela_wire_7777),
        .dout(new_Jinkela_wire_7778)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    bfr new_Jinkela_buffer_5814 (
        .din(new_Jinkela_wire_7806),
        .dout(new_Jinkela_wire_7807)
    );

    bfr new_Jinkela_buffer_748 (
        .din(G23),
        .dout(new_Jinkela_wire_1502)
    );

    bfr new_Jinkela_buffer_5794 (
        .din(new_Jinkela_wire_7778),
        .dout(new_Jinkela_wire_7779)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_1443),
        .dout(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_5868 (
        .din(_1111_),
        .dout(new_Jinkela_wire_7880)
    );

    bfr new_Jinkela_buffer_5839 (
        .din(new_Jinkela_wire_7833),
        .dout(new_Jinkela_wire_7834)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_5795 (
        .din(new_Jinkela_wire_7779),
        .dout(new_Jinkela_wire_7780)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_5815 (
        .din(new_Jinkela_wire_7807),
        .dout(new_Jinkela_wire_7808)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_5796 (
        .din(new_Jinkela_wire_7780),
        .dout(new_Jinkela_wire_7781)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_1444),
        .dout(new_Jinkela_wire_1445)
    );

    bfr new_Jinkela_buffer_5853 (
        .din(new_Jinkela_wire_7851),
        .dout(new_Jinkela_wire_7852)
    );

    bfr new_Jinkela_buffer_5797 (
        .din(new_Jinkela_wire_7781),
        .dout(new_Jinkela_wire_7782)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_1445),
        .dout(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_5816 (
        .din(new_Jinkela_wire_7808),
        .dout(new_Jinkela_wire_7809)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_1487),
        .dout(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_5848 (
        .din(new_Jinkela_wire_7844),
        .dout(new_Jinkela_wire_7845)
    );

    bfr new_Jinkela_buffer_5840 (
        .din(new_Jinkela_wire_7834),
        .dout(new_Jinkela_wire_7835)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_1446),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_5817 (
        .din(new_Jinkela_wire_7809),
        .dout(new_Jinkela_wire_7810)
    );

    bfr new_Jinkela_buffer_739 (
        .din(G22),
        .dout(new_Jinkela_wire_1489)
    );

    and_bi _1445_ (
        .a(new_Jinkela_wire_772),
        .b(new_Jinkela_wire_2987),
        .c(_0746_)
    );

    and_bi _2159_ (
        .a(new_Jinkela_wire_3679),
        .b(new_Jinkela_wire_2155),
        .c(_0194_)
    );

    bfr new_Jinkela_buffer_3502 (
        .din(new_Jinkela_wire_4928),
        .dout(new_Jinkela_wire_4929)
    );

    and_ii _1446_ (
        .a(new_Jinkela_wire_4985),
        .b(new_Jinkela_wire_2203),
        .c(_0747_)
    );

    and_bi _2160_ (
        .a(_0193_),
        .b(_0194_),
        .c(_0195_)
    );

    spl2 new_Jinkela_splitter_548 (
        .a(new_net_18),
        .b(new_Jinkela_wire_4999),
        .c(new_Jinkela_wire_5001)
    );

    or_bi _1447_ (
        .a(new_Jinkela_wire_7211),
        .b(new_Jinkela_wire_6558),
        .c(_0748_)
    );

    and_ii _2161_ (
        .a(new_Jinkela_wire_5127),
        .b(new_Jinkela_wire_5051),
        .c(_0196_)
    );

    bfr new_Jinkela_buffer_3503 (
        .din(new_Jinkela_wire_4929),
        .dout(new_Jinkela_wire_4930)
    );

    or_ii _1448_ (
        .a(new_Jinkela_wire_23),
        .b(new_Jinkela_wire_163),
        .c(_0749_)
    );

    and_bb _2162_ (
        .a(new_Jinkela_wire_5125),
        .b(new_Jinkela_wire_5050),
        .c(_0197_)
    );

    bfr new_Jinkela_buffer_3511 (
        .din(new_Jinkela_wire_4937),
        .dout(new_Jinkela_wire_4938)
    );

    and_bi _1449_ (
        .a(new_Jinkela_wire_739),
        .b(new_Jinkela_wire_7),
        .c(_0750_)
    );

    and_ii _2163_ (
        .a(_0197_),
        .b(_0196_),
        .c(_0198_)
    );

    bfr new_Jinkela_buffer_3504 (
        .din(new_Jinkela_wire_4930),
        .dout(new_Jinkela_wire_4931)
    );

    and_bi _1450_ (
        .a(_0749_),
        .b(new_Jinkela_wire_2538),
        .c(_0751_)
    );

    and_bb _2164_ (
        .a(new_Jinkela_wire_10),
        .b(new_Jinkela_wire_1029),
        .c(_0199_)
    );

    spl2 new_Jinkela_splitter_545 (
        .a(_0746_),
        .b(new_Jinkela_wire_4984),
        .c(new_Jinkela_wire_4986)
    );

    bfr new_Jinkela_buffer_3554 (
        .din(new_Jinkela_wire_4999),
        .dout(new_Jinkela_wire_5000)
    );

    and_bi _1451_ (
        .a(new_Jinkela_wire_514),
        .b(new_Jinkela_wire_2452),
        .c(_0752_)
    );

    and_bi _2165_ (
        .a(new_Jinkela_wire_625),
        .b(new_Jinkela_wire_5),
        .c(_0200_)
    );

    bfr new_Jinkela_buffer_3505 (
        .din(new_Jinkela_wire_4931),
        .dout(new_Jinkela_wire_4932)
    );

    and_bi _1452_ (
        .a(new_Jinkela_wire_2451),
        .b(new_Jinkela_wire_515),
        .c(_0753_)
    );

    and_ii _2166_ (
        .a(_0200_),
        .b(_0199_),
        .c(_0201_)
    );

    bfr new_Jinkela_buffer_3512 (
        .din(new_Jinkela_wire_4938),
        .dout(new_Jinkela_wire_4939)
    );

    or_bb _1453_ (
        .a(new_Jinkela_wire_7964),
        .b(new_Jinkela_wire_4424),
        .c(_0754_)
    );

    and_bi _2167_ (
        .a(new_Jinkela_wire_3768),
        .b(new_Jinkela_wire_7469),
        .c(_0202_)
    );

    bfr new_Jinkela_buffer_3506 (
        .din(new_Jinkela_wire_4932),
        .dout(new_Jinkela_wire_4933)
    );

    or_ii _1454_ (
        .a(new_Jinkela_wire_17),
        .b(new_Jinkela_wire_439),
        .c(_0755_)
    );

    and_bi _2168_ (
        .a(new_Jinkela_wire_7471),
        .b(new_Jinkela_wire_3769),
        .c(_0203_)
    );

    and_bi _1455_ (
        .a(new_Jinkela_wire_1428),
        .b(new_Jinkela_wire_9),
        .c(_0756_)
    );

    or_bb _2169_ (
        .a(_0203_),
        .b(_0202_),
        .c(_0204_)
    );

    bfr new_Jinkela_buffer_3513 (
        .din(new_Jinkela_wire_4939),
        .dout(new_Jinkela_wire_4940)
    );

    and_bi _1456_ (
        .a(_0755_),
        .b(new_Jinkela_wire_4605),
        .c(_0757_)
    );

    or_ii _2170_ (
        .a(new_Jinkela_wire_6192),
        .b(new_Jinkela_wire_7082),
        .c(_0205_)
    );

    bfr new_Jinkela_buffer_3547 (
        .din(new_Jinkela_wire_4984),
        .dout(new_Jinkela_wire_4985)
    );

    and_bi _1457_ (
        .a(new_Jinkela_wire_3029),
        .b(new_Jinkela_wire_278),
        .c(_0758_)
    );

    and_bi _2171_ (
        .a(new_Jinkela_wire_6499),
        .b(new_Jinkela_wire_7081),
        .c(_0206_)
    );

    bfr new_Jinkela_buffer_3514 (
        .din(new_Jinkela_wire_4940),
        .dout(new_Jinkela_wire_4941)
    );

    and_bi _1458_ (
        .a(new_Jinkela_wire_279),
        .b(new_Jinkela_wire_3028),
        .c(_0759_)
    );

    and_bi _2172_ (
        .a(_0205_),
        .b(_0206_),
        .c(_0207_)
    );

    bfr new_Jinkela_buffer_3555 (
        .din(new_Jinkela_wire_5005),
        .dout(new_Jinkela_wire_5006)
    );

    or_bb _1459_ (
        .a(new_Jinkela_wire_3194),
        .b(new_Jinkela_wire_7840),
        .c(_0760_)
    );

    and_ii _2173_ (
        .a(new_Jinkela_wire_3465),
        .b(new_Jinkela_wire_7928),
        .c(_0208_)
    );

    bfr new_Jinkela_buffer_3515 (
        .din(new_Jinkela_wire_4941),
        .dout(new_Jinkela_wire_4942)
    );

    or_bb _1460_ (
        .a(new_Jinkela_wire_3250),
        .b(new_Jinkela_wire_5788),
        .c(_0761_)
    );

    and_bb _2174_ (
        .a(new_Jinkela_wire_3466),
        .b(new_Jinkela_wire_7929),
        .c(_0209_)
    );

    spl4L new_Jinkela_splitter_546 (
        .a(new_Jinkela_wire_4986),
        .d(new_Jinkela_wire_4987),
        .e(new_Jinkela_wire_4988),
        .b(new_Jinkela_wire_4989),
        .c(new_Jinkela_wire_4990)
    );

    spl2 new_Jinkela_splitter_551 (
        .a(_0706_),
        .b(new_Jinkela_wire_5052),
        .c(new_Jinkela_wire_5053)
    );

    or_bb _1461_ (
        .a(new_Jinkela_wire_6099),
        .b(new_Jinkela_wire_4613),
        .c(_0762_)
    );

    and_ii _2175_ (
        .a(_0209_),
        .b(_0208_),
        .c(_0210_)
    );

    bfr new_Jinkela_buffer_3516 (
        .din(new_Jinkela_wire_4942),
        .dout(new_Jinkela_wire_4943)
    );

    or_bi _1462_ (
        .a(new_Jinkela_wire_7884),
        .b(new_Jinkela_wire_1959),
        .c(_0763_)
    );

    and_ii _2176_ (
        .a(new_Jinkela_wire_5123),
        .b(new_Jinkela_wire_7515),
        .c(_0211_)
    );

    bfr new_Jinkela_buffer_3580 (
        .din(_0556_),
        .dout(new_Jinkela_wire_5031)
    );

    spl2 new_Jinkela_splitter_547 (
        .a(new_Jinkela_wire_4990),
        .b(new_Jinkela_wire_4991),
        .c(new_Jinkela_wire_4992)
    );

    and_bi _1463_ (
        .a(new_Jinkela_wire_1426),
        .b(new_Jinkela_wire_3163),
        .c(_0764_)
    );

    and_bb _2177_ (
        .a(new_Jinkela_wire_5124),
        .b(new_Jinkela_wire_7516),
        .c(_0212_)
    );

    bfr new_Jinkela_buffer_3517 (
        .din(new_Jinkela_wire_4943),
        .dout(new_Jinkela_wire_4944)
    );

    or_bi _1464_ (
        .a(new_Jinkela_wire_7883),
        .b(new_Jinkela_wire_1422),
        .c(_0765_)
    );

    and_ii _2178_ (
        .a(_0212_),
        .b(_0211_),
        .c(_0213_)
    );

    spl4L new_Jinkela_splitter_549 (
        .a(new_Jinkela_wire_5001),
        .d(new_Jinkela_wire_5002),
        .e(new_Jinkela_wire_5003),
        .b(new_Jinkela_wire_5004),
        .c(new_Jinkela_wire_5005)
    );

    and_bi _1465_ (
        .a(new_Jinkela_wire_7037),
        .b(new_Jinkela_wire_2200),
        .c(_0766_)
    );

    or_bb _2179_ (
        .a(new_Jinkela_wire_5687),
        .b(new_Jinkela_wire_4313),
        .c(_0214_)
    );

    bfr new_Jinkela_buffer_3518 (
        .din(new_Jinkela_wire_4944),
        .dout(new_Jinkela_wire_4945)
    );

    and_ii _1466_ (
        .a(new_Jinkela_wire_4427),
        .b(new_Jinkela_wire_4989),
        .c(_0767_)
    );

    and_bb _2180_ (
        .a(new_Jinkela_wire_5688),
        .b(new_Jinkela_wire_4314),
        .c(_0215_)
    );

    spl4L new_Jinkela_splitter_550 (
        .a(_0940_),
        .d(new_Jinkela_wire_5048),
        .e(new_Jinkela_wire_5049),
        .b(new_Jinkela_wire_5050),
        .c(new_Jinkela_wire_5051)
    );

    bfr new_Jinkela_buffer_3548 (
        .din(new_Jinkela_wire_4992),
        .dout(new_Jinkela_wire_4993)
    );

    and_bi _1467_ (
        .a(_0767_),
        .b(new_Jinkela_wire_3215),
        .c(_0768_)
    );

    and_bi _2181_ (
        .a(_0214_),
        .b(_0215_),
        .c(new_net_16)
    );

    bfr new_Jinkela_buffer_3519 (
        .din(new_Jinkela_wire_4945),
        .dout(new_Jinkela_wire_4946)
    );

    or_bb _1468_ (
        .a(_0768_),
        .b(new_Jinkela_wire_7969),
        .c(_0769_)
    );

    and_bb _2182_ (
        .a(new_Jinkela_wire_1134),
        .b(new_Jinkela_wire_298),
        .c(new_net_14)
    );

    and_ii _1469_ (
        .a(new_Jinkela_wire_3524),
        .b(new_Jinkela_wire_7847),
        .c(_0770_)
    );

    and_bb _2183_ (
        .a(new_Jinkela_wire_421),
        .b(new_Jinkela_wire_574),
        .c(new_net_2367)
    );

    bfr new_Jinkela_buffer_3520 (
        .din(new_Jinkela_wire_4946),
        .dout(new_Jinkela_wire_4947)
    );

    or_bb _1470_ (
        .a(_0770_),
        .b(new_Jinkela_wire_3202),
        .c(_0771_)
    );

    and_bi _2184_ (
        .a(new_Jinkela_wire_1127),
        .b(new_Jinkela_wire_117),
        .c(new_net_2393)
    );

    and_bi _1471_ (
        .a(new_Jinkela_wire_6677),
        .b(new_Jinkela_wire_1962),
        .c(_0772_)
    );

    or_bi _2185_ (
        .a(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_623),
        .c(_0216_)
    );

    bfr new_Jinkela_buffer_3521 (
        .din(new_Jinkela_wire_4947),
        .dout(new_Jinkela_wire_4948)
    );

    and_bi _1472_ (
        .a(new_Jinkela_wire_1963),
        .b(new_Jinkela_wire_6678),
        .c(_0773_)
    );

    and_bb _2186_ (
        .a(new_Jinkela_wire_270),
        .b(new_Jinkela_wire_1559),
        .c(_0217_)
    );

    bfr new_Jinkela_buffer_3549 (
        .din(new_Jinkela_wire_4993),
        .dout(new_Jinkela_wire_4994)
    );

    or_bb _1473_ (
        .a(_0773_),
        .b(_0772_),
        .c(_0774_)
    );

    or_bb _2187_ (
        .a(new_Jinkela_wire_1985),
        .b(new_Jinkela_wire_6505),
        .c(_0218_)
    );

    bfr new_Jinkela_buffer_3522 (
        .din(new_Jinkela_wire_4948),
        .dout(new_Jinkela_wire_4949)
    );

    and_bi _1474_ (
        .a(new_Jinkela_wire_5931),
        .b(new_Jinkela_wire_3372),
        .c(_0775_)
    );

    and_bi _2188_ (
        .a(new_Jinkela_wire_2422),
        .b(_0218_),
        .c(_0219_)
    );

    or_bb _1475_ (
        .a(_0775_),
        .b(new_Jinkela_wire_5114),
        .c(_0776_)
    );

    and_bi _2189_ (
        .a(new_Jinkela_wire_583),
        .b(_0219_),
        .c(new_net_2399)
    );

    bfr new_Jinkela_buffer_3523 (
        .din(new_Jinkela_wire_4949),
        .dout(new_Jinkela_wire_4950)
    );

    or_bb _1476_ (
        .a(new_Jinkela_wire_5233),
        .b(new_Jinkela_wire_1084),
        .c(_0777_)
    );

    or_bi _2190_ (
        .a(new_Jinkela_wire_1560),
        .b(new_Jinkela_wire_1025),
        .c(_0220_)
    );

    bfr new_Jinkela_buffer_3581 (
        .din(new_Jinkela_wire_5031),
        .dout(new_Jinkela_wire_5032)
    );

    bfr new_Jinkela_buffer_3550 (
        .din(new_Jinkela_wire_4994),
        .dout(new_Jinkela_wire_4995)
    );

    inv _1477_ (
        .din(new_Jinkela_wire_1251),
        .dout(_0778_)
    );

    and_bb _2191_ (
        .a(new_Jinkela_wire_1371),
        .b(new_Jinkela_wire_1563),
        .c(_0221_)
    );

    bfr new_Jinkela_buffer_3524 (
        .din(new_Jinkela_wire_4950),
        .dout(new_Jinkela_wire_4951)
    );

    or_bb _1478_ (
        .a(new_Jinkela_wire_200),
        .b(new_Jinkela_wire_319),
        .c(_0779_)
    );

    or_bb _2192_ (
        .a(new_Jinkela_wire_4600),
        .b(new_Jinkela_wire_6502),
        .c(_0222_)
    );

    and_bi _1479_ (
        .a(new_Jinkela_wire_204),
        .b(new_Jinkela_wire_221),
        .c(_0780_)
    );

    and_bi _2193_ (
        .a(new_Jinkela_wire_6557),
        .b(_0222_),
        .c(_0223_)
    );

    bfr new_Jinkela_buffer_3525 (
        .din(new_Jinkela_wire_4951),
        .dout(new_Jinkela_wire_4952)
    );

    and_bi _1480_ (
        .a(_0779_),
        .b(_0780_),
        .c(_0781_)
    );

    and_bi _2194_ (
        .a(new_Jinkela_wire_582),
        .b(_0223_),
        .c(new_net_2503)
    );

    bfr new_Jinkela_buffer_3551 (
        .din(new_Jinkela_wire_4995),
        .dout(new_Jinkela_wire_4996)
    );

    or_bb _1481_ (
        .a(_0781_),
        .b(new_Jinkela_wire_6352),
        .c(_0782_)
    );

    or_bi _2195_ (
        .a(new_Jinkela_wire_1566),
        .b(new_Jinkela_wire_1391),
        .c(_0224_)
    );

    bfr new_Jinkela_buffer_3526 (
        .din(new_Jinkela_wire_4952),
        .dout(new_Jinkela_wire_4953)
    );

    or_ii _1482_ (
        .a(new_Jinkela_wire_1581),
        .b(new_Jinkela_wire_193),
        .c(_0783_)
    );

    and_bb _2196_ (
        .a(new_Jinkela_wire_1596),
        .b(new_Jinkela_wire_1561),
        .c(_0225_)
    );

    and_bi _1483_ (
        .a(new_Jinkela_wire_1292),
        .b(new_Jinkela_wire_203),
        .c(_0784_)
    );

    or_bb _2197_ (
        .a(new_Jinkela_wire_1860),
        .b(new_Jinkela_wire_6507),
        .c(_0226_)
    );

    bfr new_Jinkela_buffer_3527 (
        .din(new_Jinkela_wire_4953),
        .dout(new_Jinkela_wire_4954)
    );

    and_bi _1484_ (
        .a(new_Jinkela_wire_6892),
        .b(_0784_),
        .c(_0785_)
    );

    and_bi _2198_ (
        .a(new_Jinkela_wire_3468),
        .b(_0226_),
        .c(_0227_)
    );

    bfr new_Jinkela_buffer_3556 (
        .din(new_Jinkela_wire_5006),
        .dout(new_Jinkela_wire_5007)
    );

    bfr new_Jinkela_buffer_3552 (
        .din(new_Jinkela_wire_4996),
        .dout(new_Jinkela_wire_4997)
    );

    and_bi _1485_ (
        .a(new_Jinkela_wire_6351),
        .b(_0785_),
        .c(_0786_)
    );

    and_bi _2199_ (
        .a(new_Jinkela_wire_584),
        .b(_0227_),
        .c(new_net_2459)
    );

    bfr new_Jinkela_buffer_3528 (
        .din(new_Jinkela_wire_4954),
        .dout(new_Jinkela_wire_4955)
    );

    and_bi _1486_ (
        .a(_0782_),
        .b(_0786_),
        .c(_0787_)
    );

    or_bi _2200_ (
        .a(new_Jinkela_wire_1558),
        .b(new_Jinkela_wire_1355),
        .c(_0228_)
    );

    bfr new_Jinkela_buffer_4130 (
        .din(new_Jinkela_wire_5693),
        .dout(new_Jinkela_wire_5694)
    );

    bfr new_Jinkela_buffer_4114 (
        .din(new_Jinkela_wire_5673),
        .dout(new_Jinkela_wire_5674)
    );

    bfr new_Jinkela_buffer_4133 (
        .din(new_Jinkela_wire_5697),
        .dout(new_Jinkela_wire_5698)
    );

    bfr new_Jinkela_buffer_4115 (
        .din(new_Jinkela_wire_5674),
        .dout(new_Jinkela_wire_5675)
    );

    bfr new_Jinkela_buffer_4131 (
        .din(new_Jinkela_wire_5694),
        .dout(new_Jinkela_wire_5695)
    );

    bfr new_Jinkela_buffer_4116 (
        .din(new_Jinkela_wire_5675),
        .dout(new_Jinkela_wire_5676)
    );

    bfr new_Jinkela_buffer_4117 (
        .din(new_Jinkela_wire_5676),
        .dout(new_Jinkela_wire_5677)
    );

    bfr new_Jinkela_buffer_4118 (
        .din(new_Jinkela_wire_5677),
        .dout(new_Jinkela_wire_5678)
    );

    bfr new_Jinkela_buffer_4134 (
        .din(new_Jinkela_wire_5703),
        .dout(new_Jinkela_wire_5704)
    );

    bfr new_Jinkela_buffer_4119 (
        .din(new_Jinkela_wire_5678),
        .dout(new_Jinkela_wire_5679)
    );

    bfr new_Jinkela_buffer_4137 (
        .din(new_Jinkela_wire_5708),
        .dout(new_Jinkela_wire_5709)
    );

    bfr new_Jinkela_buffer_4120 (
        .din(new_Jinkela_wire_5679),
        .dout(new_Jinkela_wire_5680)
    );

    bfr new_Jinkela_buffer_4158 (
        .din(_0075_),
        .dout(new_Jinkela_wire_5730)
    );

    bfr new_Jinkela_buffer_4121 (
        .din(new_Jinkela_wire_5680),
        .dout(new_Jinkela_wire_5681)
    );

    spl2 new_Jinkela_splitter_603 (
        .a(_0015_),
        .b(new_Jinkela_wire_5731),
        .c(new_Jinkela_wire_5732)
    );

    bfr new_Jinkela_buffer_4159 (
        .din(new_net_2415),
        .dout(new_Jinkela_wire_5733)
    );

    bfr new_Jinkela_buffer_4122 (
        .din(new_Jinkela_wire_5681),
        .dout(new_Jinkela_wire_5682)
    );

    bfr new_Jinkela_buffer_4138 (
        .din(new_Jinkela_wire_5709),
        .dout(new_Jinkela_wire_5710)
    );

    bfr new_Jinkela_buffer_4123 (
        .din(new_Jinkela_wire_5682),
        .dout(new_Jinkela_wire_5683)
    );

    spl3L new_Jinkela_splitter_606 (
        .a(_0754_),
        .d(new_Jinkela_wire_5788),
        .b(new_Jinkela_wire_5789),
        .c(new_Jinkela_wire_5790)
    );

    bfr new_Jinkela_buffer_4160 (
        .din(new_Jinkela_wire_5733),
        .dout(new_Jinkela_wire_5734)
    );

    bfr new_Jinkela_buffer_4124 (
        .din(new_Jinkela_wire_5683),
        .dout(new_Jinkela_wire_5684)
    );

    bfr new_Jinkela_buffer_4139 (
        .din(new_Jinkela_wire_5710),
        .dout(new_Jinkela_wire_5711)
    );

    bfr new_Jinkela_buffer_4125 (
        .din(new_Jinkela_wire_5684),
        .dout(new_Jinkela_wire_5685)
    );

    bfr new_Jinkela_buffer_4126 (
        .din(new_Jinkela_wire_5685),
        .dout(new_Jinkela_wire_5686)
    );

    bfr new_Jinkela_buffer_4140 (
        .din(new_Jinkela_wire_5711),
        .dout(new_Jinkela_wire_5712)
    );

    spl2 new_Jinkela_splitter_604 (
        .a(new_net_19),
        .b(new_Jinkela_wire_5773),
        .c(new_Jinkela_wire_5775)
    );

    bfr new_Jinkela_buffer_4141 (
        .din(new_Jinkela_wire_5712),
        .dout(new_Jinkela_wire_5713)
    );

    bfr new_Jinkela_buffer_4215 (
        .din(_0673_),
        .dout(new_Jinkela_wire_5815)
    );

    bfr new_Jinkela_buffer_4142 (
        .din(new_Jinkela_wire_5713),
        .dout(new_Jinkela_wire_5714)
    );

    bfr new_Jinkela_buffer_4161 (
        .din(new_Jinkela_wire_5734),
        .dout(new_Jinkela_wire_5735)
    );

    bfr new_Jinkela_buffer_4143 (
        .din(new_Jinkela_wire_5714),
        .dout(new_Jinkela_wire_5715)
    );

    spl4L new_Jinkela_splitter_605 (
        .a(new_Jinkela_wire_5775),
        .d(new_Jinkela_wire_5776),
        .e(new_Jinkela_wire_5777),
        .b(new_Jinkela_wire_5778),
        .c(new_Jinkela_wire_5779)
    );

    bfr new_Jinkela_buffer_4144 (
        .din(new_Jinkela_wire_5715),
        .dout(new_Jinkela_wire_5716)
    );

    bfr new_Jinkela_buffer_4162 (
        .din(new_Jinkela_wire_5735),
        .dout(new_Jinkela_wire_5736)
    );

    bfr new_Jinkela_buffer_4145 (
        .din(new_Jinkela_wire_5716),
        .dout(new_Jinkela_wire_5717)
    );

    bfr new_Jinkela_buffer_4146 (
        .din(new_Jinkela_wire_5717),
        .dout(new_Jinkela_wire_5718)
    );

    bfr new_Jinkela_buffer_4163 (
        .din(new_Jinkela_wire_5736),
        .dout(new_Jinkela_wire_5737)
    );

    bfr new_Jinkela_buffer_4147 (
        .din(new_Jinkela_wire_5718),
        .dout(new_Jinkela_wire_5719)
    );

    spl3L new_Jinkela_splitter_609 (
        .a(_0266_),
        .d(new_Jinkela_wire_5802),
        .b(new_Jinkela_wire_5805),
        .c(new_Jinkela_wire_5810)
    );

    bfr new_Jinkela_buffer_4199 (
        .din(new_Jinkela_wire_5773),
        .dout(new_Jinkela_wire_5774)
    );

    bfr new_Jinkela_buffer_4148 (
        .din(new_Jinkela_wire_5719),
        .dout(new_Jinkela_wire_5720)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_net_2399),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1987),
        .dout(new_Jinkela_wire_1988)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1989),
        .dout(new_Jinkela_wire_1990)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_net_2447),
        .dout(new_Jinkela_wire_2034)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1990),
        .dout(new_Jinkela_wire_1991)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1991),
        .dout(new_Jinkela_wire_1992)
    );

    spl2 new_Jinkela_splitter_343 (
        .a(new_net_6),
        .b(new_Jinkela_wire_2064),
        .c(new_Jinkela_wire_2066)
    );

    spl2 new_Jinkela_splitter_345 (
        .a(_1086_),
        .b(new_Jinkela_wire_2086),
        .c(new_Jinkela_wire_2087)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_2000),
        .dout(new_Jinkela_wire_2001)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1993),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_2034),
        .dout(new_Jinkela_wire_2035)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_2001),
        .dout(new_Jinkela_wire_2002)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    and_bi _1296_ (
        .a(new_Jinkela_wire_1365),
        .b(new_Jinkela_wire_401),
        .c(_0603_)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_2070),
        .dout(new_Jinkela_wire_2071)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1996),
        .dout(new_Jinkela_wire_1997)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_2002),
        .dout(new_Jinkela_wire_2003)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1997),
        .dout(new_Jinkela_wire_1998)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_2035),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(new_Jinkela_wire_2003),
        .dout(new_Jinkela_wire_2004)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_2064),
        .dout(new_Jinkela_wire_2065)
    );

    spl4L new_Jinkela_splitter_344 (
        .a(new_Jinkela_wire_2066),
        .d(new_Jinkela_wire_2067),
        .e(new_Jinkela_wire_2068),
        .b(new_Jinkela_wire_2069),
        .c(new_Jinkela_wire_2070)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_Jinkela_wire_2004),
        .dout(new_Jinkela_wire_2005)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_2036),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_2005),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_2087),
        .dout(new_Jinkela_wire_2088)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_2006),
        .dout(new_Jinkela_wire_2007)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_2007),
        .dout(new_Jinkela_wire_2008)
    );

    spl2 new_Jinkela_splitter_346 (
        .a(_0183_),
        .b(new_Jinkela_wire_2090),
        .c(new_Jinkela_wire_2091)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_2008),
        .dout(new_Jinkela_wire_2009)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_2009),
        .dout(new_Jinkela_wire_2010)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_2010),
        .dout(new_Jinkela_wire_2011)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_2011),
        .dout(new_Jinkela_wire_2012)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_2012),
        .dout(new_Jinkela_wire_2013)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(new_Jinkela_wire_2013),
        .dout(new_Jinkela_wire_2014)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(_0636_),
        .dout(new_Jinkela_wire_2092)
    );

    bfr new_Jinkela_buffer_654 (
        .din(G74),
        .dout(new_Jinkela_wire_1356)
    );

    spl2 new_Jinkela_splitter_412 (
        .a(_0763_),
        .b(new_Jinkela_wire_3160),
        .c(new_Jinkela_wire_3162)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_1347),
        .dout(new_Jinkela_wire_1348)
    );

    bfr new_Jinkela_buffer_1992 (
        .din(new_Jinkela_wire_3078),
        .dout(new_Jinkela_wire_3079)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_1349),
        .dout(new_Jinkela_wire_1350)
    );

    spl3L new_Jinkela_splitter_414 (
        .a(_0867_),
        .d(new_Jinkela_wire_3170),
        .b(new_Jinkela_wire_3171),
        .c(new_Jinkela_wire_3172)
    );

    bfr new_Jinkela_buffer_2002 (
        .din(new_Jinkela_wire_3100),
        .dout(new_Jinkela_wire_3101)
    );

    spl3L new_Jinkela_splitter_252 (
        .a(G130),
        .d(new_Jinkela_wire_1361),
        .b(new_Jinkela_wire_1362),
        .c(new_Jinkela_wire_1363)
    );

    bfr new_Jinkela_buffer_1993 (
        .din(new_Jinkela_wire_3079),
        .dout(new_Jinkela_wire_3080)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_1354),
        .dout(new_Jinkela_wire_1355)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_1350),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_2006 (
        .din(new_Jinkela_wire_3106),
        .dout(new_Jinkela_wire_3107)
    );

    bfr new_Jinkela_buffer_1994 (
        .din(new_Jinkela_wire_3080),
        .dout(new_Jinkela_wire_3081)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(new_Jinkela_wire_1351),
        .b(new_Jinkela_wire_1352),
        .c(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_2003 (
        .din(new_Jinkela_wire_3101),
        .dout(new_Jinkela_wire_3102)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_1356),
        .dout(new_Jinkela_wire_1357)
    );

    spl2 new_Jinkela_splitter_406 (
        .a(new_Jinkela_wire_3081),
        .b(new_Jinkela_wire_3082),
        .c(new_Jinkela_wire_3083)
    );

    spl3L new_Jinkela_splitter_253 (
        .a(new_Jinkela_wire_1363),
        .d(new_Jinkela_wire_1364),
        .b(new_Jinkela_wire_1365),
        .c(new_Jinkela_wire_1366)
    );

    bfr new_Jinkela_buffer_658 (
        .din(G164),
        .dout(new_Jinkela_wire_1368)
    );

    spl2 new_Jinkela_splitter_411 (
        .a(new_Jinkela_wire_3102),
        .b(new_Jinkela_wire_3103),
        .c(new_Jinkela_wire_3104)
    );

    bfr new_Jinkela_buffer_2036 (
        .din(new_Jinkela_wire_3136),
        .dout(new_Jinkela_wire_3137)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_1357),
        .dout(new_Jinkela_wire_1358)
    );

    bfr new_Jinkela_buffer_2063 (
        .din(_0791_),
        .dout(new_Jinkela_wire_3175)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_1366),
        .dout(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_2060 (
        .din(new_Jinkela_wire_3166),
        .dout(new_Jinkela_wire_3167)
    );

    bfr new_Jinkela_buffer_659 (
        .din(G38),
        .dout(new_Jinkela_wire_1369)
    );

    bfr new_Jinkela_buffer_2007 (
        .din(new_Jinkela_wire_3107),
        .dout(new_Jinkela_wire_3108)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(new_Jinkela_wire_1358),
        .b(new_Jinkela_wire_1359),
        .c(new_Jinkela_wire_1360)
    );

    bfr new_Jinkela_buffer_2008 (
        .din(new_Jinkela_wire_3108),
        .dout(new_Jinkela_wire_3109)
    );

    bfr new_Jinkela_buffer_662 (
        .din(G76),
        .dout(new_Jinkela_wire_1372)
    );

    bfr new_Jinkela_buffer_2037 (
        .din(new_Jinkela_wire_3137),
        .dout(new_Jinkela_wire_3138)
    );

    bfr new_Jinkela_buffer_2009 (
        .din(new_Jinkela_wire_3109),
        .dout(new_Jinkela_wire_3110)
    );

    bfr new_Jinkela_buffer_660 (
        .din(G10),
        .dout(new_Jinkela_wire_1370)
    );

    bfr new_Jinkela_buffer_2059 (
        .din(new_Jinkela_wire_3160),
        .dout(new_Jinkela_wire_3161)
    );

    bfr new_Jinkela_buffer_665 (
        .din(G116),
        .dout(new_Jinkela_wire_1377)
    );

    spl4L new_Jinkela_splitter_413 (
        .a(new_Jinkela_wire_3162),
        .d(new_Jinkela_wire_3163),
        .e(new_Jinkela_wire_3164),
        .b(new_Jinkela_wire_3165),
        .c(new_Jinkela_wire_3166)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_1370),
        .dout(new_Jinkela_wire_1371)
    );

    bfr new_Jinkela_buffer_2010 (
        .din(new_Jinkela_wire_3110),
        .dout(new_Jinkela_wire_3111)
    );

    bfr new_Jinkela_buffer_2038 (
        .din(new_Jinkela_wire_3138),
        .dout(new_Jinkela_wire_3139)
    );

    bfr new_Jinkela_buffer_668 (
        .din(G133),
        .dout(new_Jinkela_wire_1380)
    );

    bfr new_Jinkela_buffer_2011 (
        .din(new_Jinkela_wire_3111),
        .dout(new_Jinkela_wire_3112)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_1372),
        .dout(new_Jinkela_wire_1373)
    );

    spl3L new_Jinkela_splitter_416 (
        .a(_0759_),
        .d(new_Jinkela_wire_3193),
        .b(new_Jinkela_wire_3194),
        .c(new_Jinkela_wire_3195)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    bfr new_Jinkela_buffer_2012 (
        .din(new_Jinkela_wire_3112),
        .dout(new_Jinkela_wire_3113)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_1373),
        .dout(new_Jinkela_wire_1374)
    );

    bfr new_Jinkela_buffer_2039 (
        .din(new_Jinkela_wire_3139),
        .dout(new_Jinkela_wire_3140)
    );

    bfr new_Jinkela_buffer_671 (
        .din(G35),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_2013 (
        .din(new_Jinkela_wire_3113),
        .dout(new_Jinkela_wire_3114)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(new_Jinkela_wire_1374),
        .b(new_Jinkela_wire_1375),
        .c(new_Jinkela_wire_1376)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    bfr new_Jinkela_buffer_2014 (
        .din(new_Jinkela_wire_3114),
        .dout(new_Jinkela_wire_3115)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_1378),
        .dout(new_Jinkela_wire_1379)
    );

    bfr new_Jinkela_buffer_2040 (
        .din(new_Jinkela_wire_3140),
        .dout(new_Jinkela_wire_3141)
    );

    bfr new_Jinkela_buffer_673 (
        .din(G40),
        .dout(new_Jinkela_wire_1385)
    );

    bfr new_Jinkela_buffer_2015 (
        .din(new_Jinkela_wire_3115),
        .dout(new_Jinkela_wire_3116)
    );

    bfr new_Jinkela_buffer_676 (
        .din(G7),
        .dout(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_1383),
        .dout(new_Jinkela_wire_1384)
    );

    bfr new_Jinkela_buffer_2016 (
        .din(new_Jinkela_wire_3116),
        .dout(new_Jinkela_wire_3117)
    );

    bfr new_Jinkela_buffer_2041 (
        .din(new_Jinkela_wire_3141),
        .dout(new_Jinkela_wire_3142)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(G115),
        .b(new_Jinkela_wire_1392),
        .c(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_2017 (
        .din(new_Jinkela_wire_3117),
        .dout(new_Jinkela_wire_3118)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_1385),
        .dout(new_Jinkela_wire_1386)
    );

    spl4L new_Jinkela_splitter_258 (
        .a(G177),
        .d(new_Jinkela_wire_1400),
        .e(new_Jinkela_wire_1401),
        .b(new_Jinkela_wire_1402),
        .c(new_Jinkela_wire_1403)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_1390),
        .dout(new_Jinkela_wire_1391)
    );

    bfr new_Jinkela_buffer_2018 (
        .din(new_Jinkela_wire_3118),
        .dout(new_Jinkela_wire_3119)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_1386),
        .dout(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_2042 (
        .din(new_Jinkela_wire_3142),
        .dout(new_Jinkela_wire_3143)
    );

    bfr new_Jinkela_buffer_680 (
        .din(G2),
        .dout(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_2019 (
        .din(new_Jinkela_wire_3119),
        .dout(new_Jinkela_wire_3120)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(new_Jinkela_wire_1387),
        .b(new_Jinkela_wire_1388),
        .c(new_Jinkela_wire_1389)
    );

    bfr new_Jinkela_buffer_2088 (
        .din(new_net_2431),
        .dout(new_Jinkela_wire_3203)
    );

    spl4L new_Jinkela_splitter_257 (
        .a(new_Jinkela_wire_1394),
        .d(new_Jinkela_wire_1395),
        .e(new_Jinkela_wire_1396),
        .b(new_Jinkela_wire_1397),
        .c(new_Jinkela_wire_1398)
    );

    spl2 new_Jinkela_splitter_415 (
        .a(new_Jinkela_wire_3172),
        .b(new_Jinkela_wire_3173),
        .c(new_Jinkela_wire_3174)
    );

    bfr new_Jinkela_buffer_2020 (
        .din(new_Jinkela_wire_3120),
        .dout(new_Jinkela_wire_3121)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_1398),
        .dout(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_1392),
        .dout(new_Jinkela_wire_1393)
    );

    bfr new_Jinkela_buffer_2043 (
        .din(new_Jinkela_wire_3143),
        .dout(new_Jinkela_wire_3144)
    );

    bfr new_Jinkela_buffer_2021 (
        .din(new_Jinkela_wire_3121),
        .dout(new_Jinkela_wire_3122)
    );

    bfr new_Jinkela_buffer_2061 (
        .din(new_Jinkela_wire_3167),
        .dout(new_Jinkela_wire_3168)
    );

    bfr new_Jinkela_buffer_2022 (
        .din(new_Jinkela_wire_3122),
        .dout(new_Jinkela_wire_3123)
    );

    bfr new_Jinkela_buffer_696 (
        .din(G104),
        .dout(new_Jinkela_wire_1427)
    );

    spl2 new_Jinkela_splitter_262 (
        .a(G127),
        .b(new_Jinkela_wire_1429),
        .c(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_2044 (
        .din(new_Jinkela_wire_3144),
        .dout(new_Jinkela_wire_3145)
    );

    bfr new_Jinkela_buffer_5818 (
        .din(new_Jinkela_wire_7810),
        .dout(new_Jinkela_wire_7811)
    );

    bfr new_Jinkela_buffer_3507 (
        .din(new_net_2389),
        .dout(new_Jinkela_wire_4934)
    );

    bfr new_Jinkela_buffer_3496 (
        .din(new_Jinkela_wire_4922),
        .dout(new_Jinkela_wire_4923)
    );

    bfr new_Jinkela_buffer_3457 (
        .din(new_Jinkela_wire_4879),
        .dout(new_Jinkela_wire_4880)
    );

    bfr new_Jinkela_buffer_5841 (
        .din(new_Jinkela_wire_7835),
        .dout(new_Jinkela_wire_7836)
    );

    bfr new_Jinkela_buffer_5819 (
        .din(new_Jinkela_wire_7811),
        .dout(new_Jinkela_wire_7812)
    );

    bfr new_Jinkela_buffer_3470 (
        .din(new_Jinkela_wire_4892),
        .dout(new_Jinkela_wire_4893)
    );

    bfr new_Jinkela_buffer_3458 (
        .din(new_Jinkela_wire_4880),
        .dout(new_Jinkela_wire_4881)
    );

    spl3L new_Jinkela_splitter_779 (
        .a(_0762_),
        .d(new_Jinkela_wire_7883),
        .b(new_Jinkela_wire_7884),
        .c(new_Jinkela_wire_7885)
    );

    bfr new_Jinkela_buffer_5820 (
        .din(new_Jinkela_wire_7812),
        .dout(new_Jinkela_wire_7813)
    );

    bfr new_Jinkela_buffer_3480 (
        .din(new_Jinkela_wire_4902),
        .dout(new_Jinkela_wire_4903)
    );

    bfr new_Jinkela_buffer_5849 (
        .din(new_Jinkela_wire_7845),
        .dout(new_Jinkela_wire_7846)
    );

    bfr new_Jinkela_buffer_3459 (
        .din(new_Jinkela_wire_4881),
        .dout(new_Jinkela_wire_4882)
    );

    bfr new_Jinkela_buffer_5842 (
        .din(new_Jinkela_wire_7836),
        .dout(new_Jinkela_wire_7837)
    );

    bfr new_Jinkela_buffer_5821 (
        .din(new_Jinkela_wire_7813),
        .dout(new_Jinkela_wire_7814)
    );

    bfr new_Jinkela_buffer_3471 (
        .din(new_Jinkela_wire_4893),
        .dout(new_Jinkela_wire_4894)
    );

    bfr new_Jinkela_buffer_3460 (
        .din(new_Jinkela_wire_4882),
        .dout(new_Jinkela_wire_4883)
    );

    bfr new_Jinkela_buffer_5822 (
        .din(new_Jinkela_wire_7814),
        .dout(new_Jinkela_wire_7815)
    );

    bfr new_Jinkela_buffer_3461 (
        .din(new_Jinkela_wire_4883),
        .dout(new_Jinkela_wire_4884)
    );

    bfr new_Jinkela_buffer_5843 (
        .din(new_Jinkela_wire_7837),
        .dout(new_Jinkela_wire_7838)
    );

    bfr new_Jinkela_buffer_5823 (
        .din(new_Jinkela_wire_7815),
        .dout(new_Jinkela_wire_7816)
    );

    bfr new_Jinkela_buffer_3472 (
        .din(new_Jinkela_wire_4894),
        .dout(new_Jinkela_wire_4895)
    );

    bfr new_Jinkela_buffer_3462 (
        .din(new_Jinkela_wire_4884),
        .dout(new_Jinkela_wire_4885)
    );

    bfr new_Jinkela_buffer_5854 (
        .din(new_Jinkela_wire_7852),
        .dout(new_Jinkela_wire_7853)
    );

    bfr new_Jinkela_buffer_5824 (
        .din(new_Jinkela_wire_7816),
        .dout(new_Jinkela_wire_7817)
    );

    bfr new_Jinkela_buffer_3481 (
        .din(new_Jinkela_wire_4903),
        .dout(new_Jinkela_wire_4904)
    );

    bfr new_Jinkela_buffer_5850 (
        .din(new_Jinkela_wire_7846),
        .dout(new_Jinkela_wire_7847)
    );

    bfr new_Jinkela_buffer_3463 (
        .din(new_Jinkela_wire_4885),
        .dout(new_Jinkela_wire_4886)
    );

    bfr new_Jinkela_buffer_5844 (
        .din(new_Jinkela_wire_7838),
        .dout(new_Jinkela_wire_7839)
    );

    bfr new_Jinkela_buffer_5825 (
        .din(new_Jinkela_wire_7817),
        .dout(new_Jinkela_wire_7818)
    );

    bfr new_Jinkela_buffer_3473 (
        .din(new_Jinkela_wire_4895),
        .dout(new_Jinkela_wire_4896)
    );

    bfr new_Jinkela_buffer_3495 (
        .din(new_net_2467),
        .dout(new_Jinkela_wire_4922)
    );

    bfr new_Jinkela_buffer_5826 (
        .din(new_Jinkela_wire_7818),
        .dout(new_Jinkela_wire_7819)
    );

    bfr new_Jinkela_buffer_3474 (
        .din(new_Jinkela_wire_4896),
        .dout(new_Jinkela_wire_4897)
    );

    bfr new_Jinkela_buffer_3482 (
        .din(new_Jinkela_wire_4904),
        .dout(new_Jinkela_wire_4905)
    );

    bfr new_Jinkela_buffer_5870 (
        .din(new_Jinkela_wire_7881),
        .dout(new_Jinkela_wire_7882)
    );

    bfr new_Jinkela_buffer_5827 (
        .din(new_Jinkela_wire_7819),
        .dout(new_Jinkela_wire_7820)
    );

    bfr new_Jinkela_buffer_3475 (
        .din(new_Jinkela_wire_4897),
        .dout(new_Jinkela_wire_4898)
    );

    spl2 new_Jinkela_splitter_541 (
        .a(_0156_),
        .b(new_Jinkela_wire_4974),
        .c(new_Jinkela_wire_4975)
    );

    bfr new_Jinkela_buffer_5855 (
        .din(new_Jinkela_wire_7853),
        .dout(new_Jinkela_wire_7854)
    );

    bfr new_Jinkela_buffer_5828 (
        .din(new_Jinkela_wire_7820),
        .dout(new_Jinkela_wire_7821)
    );

    spl4L new_Jinkela_splitter_542 (
        .a(_0604_),
        .d(new_Jinkela_wire_4976),
        .e(new_Jinkela_wire_4977),
        .b(new_Jinkela_wire_4978),
        .c(new_Jinkela_wire_4979)
    );

    bfr new_Jinkela_buffer_3476 (
        .din(new_Jinkela_wire_4898),
        .dout(new_Jinkela_wire_4899)
    );

    bfr new_Jinkela_buffer_3483 (
        .din(new_Jinkela_wire_4905),
        .dout(new_Jinkela_wire_4906)
    );

    bfr new_Jinkela_buffer_5872 (
        .din(_0283_),
        .dout(new_Jinkela_wire_7887)
    );

    bfr new_Jinkela_buffer_5829 (
        .din(new_Jinkela_wire_7821),
        .dout(new_Jinkela_wire_7822)
    );

    bfr new_Jinkela_buffer_3497 (
        .din(new_Jinkela_wire_4923),
        .dout(new_Jinkela_wire_4924)
    );

    spl2 new_Jinkela_splitter_776 (
        .a(new_Jinkela_wire_7867),
        .b(new_Jinkela_wire_7868),
        .c(new_Jinkela_wire_7869)
    );

    bfr new_Jinkela_buffer_3484 (
        .din(new_Jinkela_wire_4906),
        .dout(new_Jinkela_wire_4907)
    );

    bfr new_Jinkela_buffer_5856 (
        .din(new_Jinkela_wire_7854),
        .dout(new_Jinkela_wire_7855)
    );

    bfr new_Jinkela_buffer_3508 (
        .din(new_Jinkela_wire_4934),
        .dout(new_Jinkela_wire_4935)
    );

    bfr new_Jinkela_buffer_3485 (
        .din(new_Jinkela_wire_4907),
        .dout(new_Jinkela_wire_4908)
    );

    bfr new_Jinkela_buffer_5857 (
        .din(new_Jinkela_wire_7855),
        .dout(new_Jinkela_wire_7856)
    );

    bfr new_Jinkela_buffer_3498 (
        .din(new_Jinkela_wire_4924),
        .dout(new_Jinkela_wire_4925)
    );

    spl4L new_Jinkela_splitter_777 (
        .a(new_Jinkela_wire_7870),
        .d(new_Jinkela_wire_7871),
        .e(new_Jinkela_wire_7872),
        .b(new_Jinkela_wire_7873),
        .c(new_Jinkela_wire_7874)
    );

    bfr new_Jinkela_buffer_3486 (
        .din(new_Jinkela_wire_4908),
        .dout(new_Jinkela_wire_4909)
    );

    bfr new_Jinkela_buffer_5858 (
        .din(new_Jinkela_wire_7856),
        .dout(new_Jinkela_wire_7857)
    );

    spl2 new_Jinkela_splitter_543 (
        .a(_1146_),
        .b(new_Jinkela_wire_4980),
        .c(new_Jinkela_wire_4981)
    );

    spl4L new_Jinkela_splitter_778 (
        .a(new_Jinkela_wire_7875),
        .d(new_Jinkela_wire_7876),
        .e(new_Jinkela_wire_7877),
        .b(new_Jinkela_wire_7878),
        .c(new_Jinkela_wire_7879)
    );

    spl2 new_Jinkela_splitter_544 (
        .a(_1209_),
        .b(new_Jinkela_wire_4982),
        .c(new_Jinkela_wire_4983)
    );

    bfr new_Jinkela_buffer_3487 (
        .din(new_Jinkela_wire_4909),
        .dout(new_Jinkela_wire_4910)
    );

    bfr new_Jinkela_buffer_5859 (
        .din(new_Jinkela_wire_7857),
        .dout(new_Jinkela_wire_7858)
    );

    bfr new_Jinkela_buffer_3499 (
        .din(new_Jinkela_wire_4925),
        .dout(new_Jinkela_wire_4926)
    );

    bfr new_Jinkela_buffer_5869 (
        .din(new_Jinkela_wire_7880),
        .dout(new_Jinkela_wire_7881)
    );

    bfr new_Jinkela_buffer_3488 (
        .din(new_Jinkela_wire_4910),
        .dout(new_Jinkela_wire_4911)
    );

    bfr new_Jinkela_buffer_5860 (
        .din(new_Jinkela_wire_7858),
        .dout(new_Jinkela_wire_7859)
    );

    bfr new_Jinkela_buffer_3509 (
        .din(new_Jinkela_wire_4935),
        .dout(new_Jinkela_wire_4936)
    );

    spl3L new_Jinkela_splitter_780 (
        .a(_0666_),
        .d(new_Jinkela_wire_7889),
        .b(new_Jinkela_wire_7890),
        .c(new_Jinkela_wire_7891)
    );

    bfr new_Jinkela_buffer_3489 (
        .din(new_Jinkela_wire_4911),
        .dout(new_Jinkela_wire_4912)
    );

    bfr new_Jinkela_buffer_5861 (
        .din(new_Jinkela_wire_7859),
        .dout(new_Jinkela_wire_7860)
    );

    bfr new_Jinkela_buffer_3500 (
        .din(new_Jinkela_wire_4926),
        .dout(new_Jinkela_wire_4927)
    );

    bfr new_Jinkela_buffer_5871 (
        .din(new_Jinkela_wire_7885),
        .dout(new_Jinkela_wire_7886)
    );

    bfr new_Jinkela_buffer_5874 (
        .din(_0813_),
        .dout(new_Jinkela_wire_7894)
    );

    bfr new_Jinkela_buffer_3490 (
        .din(new_Jinkela_wire_4912),
        .dout(new_Jinkela_wire_4913)
    );

    bfr new_Jinkela_buffer_5862 (
        .din(new_Jinkela_wire_7860),
        .dout(new_Jinkela_wire_7861)
    );

    bfr new_Jinkela_buffer_3491 (
        .din(new_Jinkela_wire_4913),
        .dout(new_Jinkela_wire_4914)
    );

    bfr new_Jinkela_buffer_5863 (
        .din(new_Jinkela_wire_7861),
        .dout(new_Jinkela_wire_7862)
    );

    bfr new_Jinkela_buffer_3501 (
        .din(new_Jinkela_wire_4927),
        .dout(new_Jinkela_wire_4928)
    );

    bfr new_Jinkela_buffer_5873 (
        .din(new_Jinkela_wire_7887),
        .dout(new_Jinkela_wire_7888)
    );

    bfr new_Jinkela_buffer_3492 (
        .din(new_Jinkela_wire_4914),
        .dout(new_Jinkela_wire_4915)
    );

    bfr new_Jinkela_buffer_5864 (
        .din(new_Jinkela_wire_7862),
        .dout(new_Jinkela_wire_7863)
    );

    bfr new_Jinkela_buffer_3510 (
        .din(new_Jinkela_wire_4936),
        .dout(new_Jinkela_wire_4937)
    );

    bfr new_Jinkela_buffer_3493 (
        .din(new_Jinkela_wire_4915),
        .dout(new_Jinkela_wire_4916)
    );

    bfr new_Jinkela_buffer_5865 (
        .din(new_Jinkela_wire_7863),
        .dout(new_Jinkela_wire_7864)
    );

    bfr new_Jinkela_buffer_4096 (
        .din(new_Jinkela_wire_5655),
        .dout(new_Jinkela_wire_5656)
    );

    bfr new_Jinkela_buffer_4074 (
        .din(new_Jinkela_wire_5625),
        .dout(new_Jinkela_wire_5626)
    );

    bfr new_Jinkela_buffer_4081 (
        .din(new_Jinkela_wire_5638),
        .dout(new_Jinkela_wire_5639)
    );

    bfr new_Jinkela_buffer_4082 (
        .din(new_Jinkela_wire_5639),
        .dout(new_Jinkela_wire_5640)
    );

    bfr new_Jinkela_buffer_4104 (
        .din(_0887_),
        .dout(new_Jinkela_wire_5664)
    );

    bfr new_Jinkela_buffer_4083 (
        .din(new_Jinkela_wire_5640),
        .dout(new_Jinkela_wire_5641)
    );

    spl2 new_Jinkela_splitter_598 (
        .a(_0213_),
        .b(new_Jinkela_wire_5687),
        .c(new_Jinkela_wire_5688)
    );

    bfr new_Jinkela_buffer_4097 (
        .din(new_Jinkela_wire_5656),
        .dout(new_Jinkela_wire_5657)
    );

    bfr new_Jinkela_buffer_4084 (
        .din(new_Jinkela_wire_5641),
        .dout(new_Jinkela_wire_5642)
    );

    bfr new_Jinkela_buffer_4127 (
        .din(_0670_),
        .dout(new_Jinkela_wire_5689)
    );

    bfr new_Jinkela_buffer_4085 (
        .din(new_Jinkela_wire_5642),
        .dout(new_Jinkela_wire_5643)
    );

    bfr new_Jinkela_buffer_4105 (
        .din(new_Jinkela_wire_5664),
        .dout(new_Jinkela_wire_5665)
    );

    bfr new_Jinkela_buffer_4098 (
        .din(new_Jinkela_wire_5657),
        .dout(new_Jinkela_wire_5658)
    );

    bfr new_Jinkela_buffer_4086 (
        .din(new_Jinkela_wire_5643),
        .dout(new_Jinkela_wire_5644)
    );

    bfr new_Jinkela_buffer_4087 (
        .din(new_Jinkela_wire_5644),
        .dout(new_Jinkela_wire_5645)
    );

    spl2 new_Jinkela_splitter_599 (
        .a(new_Jinkela_wire_5689),
        .b(new_Jinkela_wire_5690),
        .c(new_Jinkela_wire_5691)
    );

    bfr new_Jinkela_buffer_4099 (
        .din(new_Jinkela_wire_5658),
        .dout(new_Jinkela_wire_5659)
    );

    bfr new_Jinkela_buffer_4088 (
        .din(new_Jinkela_wire_5645),
        .dout(new_Jinkela_wire_5646)
    );

    bfr new_Jinkela_buffer_4089 (
        .din(new_Jinkela_wire_5646),
        .dout(new_Jinkela_wire_5647)
    );

    bfr new_Jinkela_buffer_4106 (
        .din(new_Jinkela_wire_5665),
        .dout(new_Jinkela_wire_5666)
    );

    bfr new_Jinkela_buffer_4100 (
        .din(new_Jinkela_wire_5659),
        .dout(new_Jinkela_wire_5660)
    );

    bfr new_Jinkela_buffer_4090 (
        .din(new_Jinkela_wire_5647),
        .dout(new_Jinkela_wire_5648)
    );

    bfr new_Jinkela_buffer_4091 (
        .din(new_Jinkela_wire_5648),
        .dout(new_Jinkela_wire_5649)
    );

    bfr new_Jinkela_buffer_4101 (
        .din(new_Jinkela_wire_5660),
        .dout(new_Jinkela_wire_5661)
    );

    bfr new_Jinkela_buffer_4092 (
        .din(new_Jinkela_wire_5649),
        .dout(new_Jinkela_wire_5650)
    );

    bfr new_Jinkela_buffer_4093 (
        .din(new_Jinkela_wire_5650),
        .dout(new_Jinkela_wire_5651)
    );

    spl2 new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_1),
        .c(new_Jinkela_wire_2)
    );

    bfr new_Jinkela_buffer_4107 (
        .din(new_Jinkela_wire_5666),
        .dout(new_Jinkela_wire_5667)
    );

    spl4L new_Jinkela_splitter_0 (
        .a(G124),
        .d(new_Jinkela_wire_0),
        .e(new_Jinkela_wire_3),
        .b(new_Jinkela_wire_8),
        .c(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_4102 (
        .din(new_Jinkela_wire_5661),
        .dout(new_Jinkela_wire_5662)
    );

    bfr new_Jinkela_buffer_0 (
        .din(G52),
        .dout(new_Jinkela_wire_26)
    );

    spl4L new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_3),
        .d(new_Jinkela_wire_4),
        .e(new_Jinkela_wire_5),
        .b(new_Jinkela_wire_6),
        .c(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_4132 (
        .din(_0740_),
        .dout(new_Jinkela_wire_5696)
    );

    bfr new_Jinkela_buffer_4108 (
        .din(new_Jinkela_wire_5667),
        .dout(new_Jinkela_wire_5668)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    bfr new_Jinkela_buffer_4135 (
        .din(_0588_),
        .dout(new_Jinkela_wire_5705)
    );

    bfr new_Jinkela_buffer_5 (
        .din(G48),
        .dout(new_Jinkela_wire_31)
    );

    bfr new_Jinkela_buffer_4128 (
        .din(new_Jinkela_wire_5691),
        .dout(new_Jinkela_wire_5692)
    );

    bfr new_Jinkela_buffer_4109 (
        .din(new_Jinkela_wire_5668),
        .dout(new_Jinkela_wire_5669)
    );

    bfr new_Jinkela_buffer_10 (
        .din(G72),
        .dout(new_Jinkela_wire_36)
    );

    spl4L new_Jinkela_splitter_6 (
        .a(new_Jinkela_wire_21),
        .d(new_Jinkela_wire_22),
        .e(new_Jinkela_wire_23),
        .b(new_Jinkela_wire_24),
        .c(new_Jinkela_wire_25)
    );

    spl2 new_Jinkela_splitter_602 (
        .a(_0046_),
        .b(new_Jinkela_wire_5706),
        .c(new_Jinkela_wire_5707)
    );

    bfr new_Jinkela_buffer_4110 (
        .din(new_Jinkela_wire_5669),
        .dout(new_Jinkela_wire_5670)
    );

    spl4L new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_8),
        .d(new_Jinkela_wire_9),
        .e(new_Jinkela_wire_10),
        .b(new_Jinkela_wire_11),
        .c(new_Jinkela_wire_12)
    );

    spl4L new_Jinkela_splitter_601 (
        .a(new_Jinkela_wire_5699),
        .d(new_Jinkela_wire_5700),
        .e(new_Jinkela_wire_5701),
        .b(new_Jinkela_wire_5702),
        .c(new_Jinkela_wire_5703)
    );

    spl4L new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_13),
        .d(new_Jinkela_wire_14),
        .e(new_Jinkela_wire_15),
        .b(new_Jinkela_wire_16),
        .c(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_4136 (
        .din(new_net_2505),
        .dout(new_Jinkela_wire_5708)
    );

    bfr new_Jinkela_buffer_4111 (
        .din(new_Jinkela_wire_5670),
        .dout(new_Jinkela_wire_5671)
    );

    spl3L new_Jinkela_splitter_8 (
        .a(G100),
        .d(new_Jinkela_wire_41),
        .b(new_Jinkela_wire_43),
        .c(new_Jinkela_wire_48)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    spl4L new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_16),
        .d(new_Jinkela_wire_17),
        .e(new_Jinkela_wire_18),
        .b(new_Jinkela_wire_19),
        .c(new_Jinkela_wire_20)
    );

    bfr new_Jinkela_buffer_4129 (
        .din(new_Jinkela_wire_5692),
        .dout(new_Jinkela_wire_5693)
    );

    bfr new_Jinkela_buffer_4112 (
        .din(new_Jinkela_wire_5671),
        .dout(new_Jinkela_wire_5672)
    );

    spl2 new_Jinkela_splitter_600 (
        .a(new_Jinkela_wire_5696),
        .b(new_Jinkela_wire_5697),
        .c(new_Jinkela_wire_5699)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_31),
        .dout(new_Jinkela_wire_32)
    );

    bfr new_Jinkela_buffer_4113 (
        .din(new_Jinkela_wire_5672),
        .dout(new_Jinkela_wire_5673)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(G64),
        .b(new_Jinkela_wire_641),
        .c(new_Jinkela_wire_642)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_1268),
        .dout(new_Jinkela_wire_1269)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_624),
        .dout(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_1272),
        .dout(new_Jinkela_wire_1273)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(new_Jinkela_wire_1269),
        .b(new_Jinkela_wire_1270),
        .c(new_Jinkela_wire_1271)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(new_Jinkela_wire_578),
        .b(new_Jinkela_wire_579),
        .c(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_1273),
        .dout(new_Jinkela_wire_1274)
    );

    spl4L new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_581),
        .d(new_Jinkela_wire_582),
        .e(new_Jinkela_wire_583),
        .b(new_Jinkela_wire_584),
        .c(new_Jinkela_wire_585)
    );

    spl2 new_Jinkela_splitter_238 (
        .a(G143),
        .b(new_Jinkela_wire_1299),
        .c(new_Jinkela_wire_1300)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_630 (
        .din(G20),
        .dout(new_Jinkela_wire_1294)
    );

    spl2 new_Jinkela_splitter_134 (
        .a(G142),
        .b(new_Jinkela_wire_705),
        .c(new_Jinkela_wire_706)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(new_Jinkela_wire_1274),
        .b(new_Jinkela_wire_1275),
        .c(new_Jinkela_wire_1276)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(new_Jinkela_wire_1277),
        .b(new_Jinkela_wire_1278),
        .c(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_626),
        .dout(new_Jinkela_wire_627)
    );

    bfr new_Jinkela_buffer_639 (
        .din(G107),
        .dout(new_Jinkela_wire_1307)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_1294),
        .dout(new_Jinkela_wire_1295)
    );

    spl4L new_Jinkela_splitter_235 (
        .a(new_Jinkela_wire_1280),
        .d(new_Jinkela_wire_1281),
        .e(new_Jinkela_wire_1282),
        .b(new_Jinkela_wire_1284),
        .c(new_Jinkela_wire_1289)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_586),
        .dout(new_Jinkela_wire_587)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_1282),
        .dout(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_627),
        .dout(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    spl4L new_Jinkela_splitter_236 (
        .a(new_Jinkela_wire_1284),
        .d(new_Jinkela_wire_1285),
        .e(new_Jinkela_wire_1286),
        .b(new_Jinkela_wire_1287),
        .c(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    spl4L new_Jinkela_splitter_237 (
        .a(new_Jinkela_wire_1289),
        .d(new_Jinkela_wire_1290),
        .e(new_Jinkela_wire_1291),
        .b(new_Jinkela_wire_1292),
        .c(new_Jinkela_wire_1293)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_588),
        .dout(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_1296),
        .dout(new_Jinkela_wire_1297)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_628),
        .dout(new_Jinkela_wire_629)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_1295),
        .dout(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_589),
        .dout(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_1300),
        .dout(new_Jinkela_wire_1301)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_590),
        .dout(new_Jinkela_wire_591)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_1297),
        .dout(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_629),
        .dout(new_Jinkela_wire_630)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_1301),
        .dout(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    bfr new_Jinkela_buffer_324 (
        .din(G69),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_317 (
        .din(G13),
        .dout(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_640 (
        .din(G122),
        .dout(new_Jinkela_wire_1322)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_592),
        .dout(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_1302),
        .dout(new_Jinkela_wire_1303)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_630),
        .dout(new_Jinkela_wire_631)
    );

    spl4L new_Jinkela_splitter_242 (
        .a(new_Jinkela_wire_1312),
        .d(new_Jinkela_wire_1313),
        .e(new_Jinkela_wire_1314),
        .b(new_Jinkela_wire_1315),
        .c(new_Jinkela_wire_1316)
    );

    spl4L new_Jinkela_splitter_243 (
        .a(new_Jinkela_wire_1317),
        .d(new_Jinkela_wire_1318),
        .e(new_Jinkela_wire_1319),
        .b(new_Jinkela_wire_1320),
        .c(new_Jinkela_wire_1321)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_593),
        .dout(new_Jinkela_wire_594)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(new_Jinkela_wire_1303),
        .b(new_Jinkela_wire_1304),
        .c(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_1305),
        .dout(new_Jinkela_wire_1306)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_594),
        .dout(new_Jinkela_wire_595)
    );

    bfr new_Jinkela_buffer_643 (
        .din(G90),
        .dout(new_Jinkela_wire_1325)
    );

    spl3L new_Jinkela_splitter_241 (
        .a(new_Jinkela_wire_1308),
        .d(new_Jinkela_wire_1309),
        .b(new_Jinkela_wire_1310),
        .c(new_Jinkela_wire_1311)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_631),
        .dout(new_Jinkela_wire_632)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_595),
        .dout(new_Jinkela_wire_596)
    );

    spl3L new_Jinkela_splitter_240 (
        .a(new_Jinkela_wire_1307),
        .d(new_Jinkela_wire_1308),
        .b(new_Jinkela_wire_1312),
        .c(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_644 (
        .din(G77),
        .dout(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_596),
        .dout(new_Jinkela_wire_597)
    );

    spl2 new_Jinkela_splitter_123 (
        .a(new_Jinkela_wire_632),
        .b(new_Jinkela_wire_633),
        .c(new_Jinkela_wire_634)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_1323),
        .dout(new_Jinkela_wire_1324)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_597),
        .dout(new_Jinkela_wire_598)
    );

    spl3L new_Jinkela_splitter_244 (
        .a(new_Jinkela_wire_1325),
        .d(new_Jinkela_wire_1326),
        .b(new_Jinkela_wire_1330),
        .c(new_Jinkela_wire_1335)
    );

    spl3L new_Jinkela_splitter_245 (
        .a(new_Jinkela_wire_1326),
        .d(new_Jinkela_wire_1327),
        .b(new_Jinkela_wire_1328),
        .c(new_Jinkela_wire_1329)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_634),
        .dout(new_Jinkela_wire_635)
    );

    spl4L new_Jinkela_splitter_246 (
        .a(new_Jinkela_wire_1330),
        .d(new_Jinkela_wire_1331),
        .e(new_Jinkela_wire_1332),
        .b(new_Jinkela_wire_1333),
        .c(new_Jinkela_wire_1334)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_598),
        .dout(new_Jinkela_wire_599)
    );

    spl2 new_Jinkela_splitter_249 (
        .a(G125),
        .b(new_Jinkela_wire_1345),
        .c(new_Jinkela_wire_1346)
    );

    bfr new_Jinkela_buffer_649 (
        .din(G82),
        .dout(new_Jinkela_wire_1349)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_1340),
        .dout(new_Jinkela_wire_1341)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_599),
        .dout(new_Jinkela_wire_600)
    );

    spl4L new_Jinkela_splitter_247 (
        .a(new_Jinkela_wire_1335),
        .d(new_Jinkela_wire_1336),
        .e(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_1338),
        .c(new_Jinkela_wire_1339)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_1346),
        .dout(new_Jinkela_wire_1347)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_600),
        .dout(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_1341),
        .dout(new_Jinkela_wire_1342)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_652 (
        .din(G29),
        .dout(new_Jinkela_wire_1354)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(new_Jinkela_wire_1342),
        .b(new_Jinkela_wire_1343),
        .c(new_Jinkela_wire_1344)
    );

    and_bb _2201_ (
        .a(new_Jinkela_wire_1250),
        .b(new_Jinkela_wire_1553),
        .c(_0229_)
    );

    or_bb _2202_ (
        .a(new_Jinkela_wire_4342),
        .b(new_Jinkela_wire_6501),
        .c(_0230_)
    );

    and_bi _2203_ (
        .a(new_Jinkela_wire_6233),
        .b(_0230_),
        .c(_0231_)
    );

    and_bi _2204_ (
        .a(new_Jinkela_wire_580),
        .b(_0231_),
        .c(new_net_2477)
    );

    or_bb _2205_ (
        .a(new_Jinkela_wire_1852),
        .b(new_Jinkela_wire_4979),
        .c(_0232_)
    );

    or_bb _2206_ (
        .a(new_Jinkela_wire_2398),
        .b(new_Jinkela_wire_7521),
        .c(_0233_)
    );

    or_bb _2207_ (
        .a(_0233_),
        .b(new_Jinkela_wire_6378),
        .c(_0234_)
    );

    or_bb _2208_ (
        .a(new_Jinkela_wire_4816),
        .b(new_Jinkela_wire_4465),
        .c(_0235_)
    );

    or_bb _2209_ (
        .a(new_Jinkela_wire_6426),
        .b(_0234_),
        .c(_0236_)
    );

    and_bi _2210_ (
        .a(new_Jinkela_wire_7519),
        .b(_0236_),
        .c(new_net_2447)
    );

    and_ii _2211_ (
        .a(new_Jinkela_wire_3391),
        .b(new_Jinkela_wire_7849),
        .c(_0237_)
    );

    and_bi _2212_ (
        .a(_0237_),
        .b(new_Jinkela_wire_2416),
        .c(_0238_)
    );

    or_bb _2213_ (
        .a(new_Jinkela_wire_4178),
        .b(new_Jinkela_wire_6555),
        .c(_0239_)
    );

    or_bb _2214_ (
        .a(new_Jinkela_wire_3836),
        .b(new_Jinkela_wire_2308),
        .c(_0240_)
    );

    or_bb _2215_ (
        .a(new_Jinkela_wire_5244),
        .b(new_Jinkela_wire_5055),
        .c(_0241_)
    );

    or_bb _2216_ (
        .a(_0241_),
        .b(_0240_),
        .c(_0242_)
    );

    or_bb _2217_ (
        .a(_0242_),
        .b(new_Jinkela_wire_5663),
        .c(_0243_)
    );

    and_bi _2218_ (
        .a(new_Jinkela_wire_5434),
        .b(_0243_),
        .c(new_net_2499)
    );

    or_bi _2219_ (
        .a(new_Jinkela_wire_6937),
        .b(new_Jinkela_wire_3068),
        .c(_0244_)
    );

    and_ii _2220_ (
        .a(new_Jinkela_wire_1950),
        .b(new_Jinkela_wire_3164),
        .c(new_net_2371)
    );

    and_ii _2221_ (
        .a(new_Jinkela_wire_4347),
        .b(new_Jinkela_wire_2844),
        .c(_0245_)
    );

    or_ii _2222_ (
        .a(new_Jinkela_wire_6709),
        .b(new_Jinkela_wire_2570),
        .c(_0246_)
    );

    and_bi _2223_ (
        .a(new_Jinkela_wire_4568),
        .b(new_Jinkela_wire_7650),
        .c(new_net_2425)
    );

    and_bi _2224_ (
        .a(new_Jinkela_wire_1904),
        .b(new_Jinkela_wire_1947),
        .c(_0247_)
    );

    and_ii _2225_ (
        .a(new_Jinkela_wire_3877),
        .b(new_Jinkela_wire_5662),
        .c(_0248_)
    );

    or_bb _2226_ (
        .a(_0248_),
        .b(new_Jinkela_wire_7510),
        .c(_0249_)
    );

    or_bb _2227_ (
        .a(new_Jinkela_wire_7128),
        .b(new_Jinkela_wire_6888),
        .c(new_net_2373)
    );

    or_bi _2228_ (
        .a(new_Jinkela_wire_4576),
        .b(new_Jinkela_wire_2768),
        .c(new_net_2443)
    );

    inv _2229_ (
        .din(new_Jinkela_wire_1438),
        .dout(_0250_)
    );

    or_ii _2230_ (
        .a(new_Jinkela_wire_3277),
        .b(new_Jinkela_wire_3438),
        .c(_0251_)
    );

    inv _2231_ (
        .din(new_Jinkela_wire_1260),
        .dout(_0252_)
    );

    and_bi _2232_ (
        .a(new_Jinkela_wire_4382),
        .b(new_Jinkela_wire_3432),
        .c(_0253_)
    );

    or_bb _2233_ (
        .a(_0253_),
        .b(new_Jinkela_wire_3493),
        .c(_0254_)
    );

    and_bi _2234_ (
        .a(_0251_),
        .b(new_Jinkela_wire_5200),
        .c(_0255_)
    );

    or_bi _2235_ (
        .a(new_Jinkela_wire_1259),
        .b(new_Jinkela_wire_1440),
        .c(_0256_)
    );

    and_bi _2236_ (
        .a(new_Jinkela_wire_231),
        .b(new_Jinkela_wire_2867),
        .c(_0257_)
    );

    or_bb _2237_ (
        .a(new_Jinkela_wire_1261),
        .b(new_Jinkela_wire_1439),
        .c(_0258_)
    );

    and_bi _2238_ (
        .a(new_Jinkela_wire_1492),
        .b(new_Jinkela_wire_6418),
        .c(_0259_)
    );

    or_bb _2239_ (
        .a(_0259_),
        .b(_0257_),
        .c(_0260_)
    );

    or_bb _2240_ (
        .a(new_Jinkela_wire_4193),
        .b(_0255_),
        .c(new_net_2509)
    );

    or_bi _2241_ (
        .a(new_Jinkela_wire_364),
        .b(new_Jinkela_wire_3279),
        .c(_0261_)
    );

    inv _2242_ (
        .din(new_Jinkela_wire_1593),
        .dout(_0262_)
    );

    and_bi _1487_ (
        .a(new_Jinkela_wire_1054),
        .b(new_Jinkela_wire_4177),
        .c(_0788_)
    );

    or_bb _1488_ (
        .a(_0788_),
        .b(new_Jinkela_wire_4838),
        .c(_0789_)
    );

    and_bi _1489_ (
        .a(_0777_),
        .b(new_Jinkela_wire_2652),
        .c(_0790_)
    );

    and_ii _1490_ (
        .a(_0790_),
        .b(new_Jinkela_wire_5390),
        .c(new_net_5)
    );

    and_bi _1491_ (
        .a(new_Jinkela_wire_268),
        .b(new_Jinkela_wire_6684),
        .c(_0791_)
    );

    or_bb _1492_ (
        .a(new_Jinkela_wire_5794),
        .b(new_Jinkela_wire_4612),
        .c(_0792_)
    );

    and_bb _1493_ (
        .a(new_Jinkela_wire_3527),
        .b(_0792_),
        .c(_0793_)
    );

    or_bi _1494_ (
        .a(new_Jinkela_wire_1419),
        .b(new_Jinkela_wire_3523),
        .c(_0794_)
    );

    and_bi _1495_ (
        .a(new_Jinkela_wire_7913),
        .b(new_Jinkela_wire_6245),
        .c(_0795_)
    );

    or_ii _1496_ (
        .a(new_Jinkela_wire_7012),
        .b(new_Jinkela_wire_3262),
        .c(_0796_)
    );

    and_ii _1497_ (
        .a(new_Jinkela_wire_7013),
        .b(new_Jinkela_wire_3263),
        .c(_0797_)
    );

    and_bi _1498_ (
        .a(_0796_),
        .b(_0797_),
        .c(_0798_)
    );

    or_bb _1499_ (
        .a(new_Jinkela_wire_5271),
        .b(new_Jinkela_wire_1080),
        .c(_0799_)
    );

    inv _1500_ (
        .din(new_Jinkela_wire_271),
        .dout(_0800_)
    );

    or_bb _1501_ (
        .a(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_321),
        .c(_0801_)
    );

    and_bi _1502_ (
        .a(new_Jinkela_wire_441),
        .b(new_Jinkela_wire_219),
        .c(_0802_)
    );

    and_bi _1503_ (
        .a(_0801_),
        .b(_0802_),
        .c(_0803_)
    );

    or_bb _1504_ (
        .a(_0803_),
        .b(new_Jinkela_wire_1856),
        .c(_0804_)
    );

    or_ii _1505_ (
        .a(new_Jinkela_wire_1584),
        .b(new_Jinkela_wire_444),
        .c(_0805_)
    );

    and_bi _1506_ (
        .a(new_Jinkela_wire_1285),
        .b(new_Jinkela_wire_451),
        .c(_0806_)
    );

    and_bi _1507_ (
        .a(_0805_),
        .b(_0806_),
        .c(_0807_)
    );

    and_bi _1508_ (
        .a(new_Jinkela_wire_1855),
        .b(_0807_),
        .c(_0808_)
    );

    and_bi _1509_ (
        .a(_0804_),
        .b(_0808_),
        .c(_0809_)
    );

    and_bi _1510_ (
        .a(new_Jinkela_wire_1055),
        .b(new_Jinkela_wire_5054),
        .c(_0810_)
    );

    or_bb _1511_ (
        .a(_0810_),
        .b(new_Jinkela_wire_4841),
        .c(_0811_)
    );

    and_bi _1512_ (
        .a(_0799_),
        .b(new_Jinkela_wire_5626),
        .c(_0812_)
    );

    and_ii _1513_ (
        .a(_0812_),
        .b(new_Jinkela_wire_3192),
        .c(new_net_7)
    );

    and_bi _1514_ (
        .a(new_Jinkela_wire_572),
        .b(new_Jinkela_wire_6705),
        .c(_0813_)
    );

    and_ii _1515_ (
        .a(new_Jinkela_wire_5865),
        .b(new_Jinkela_wire_7043),
        .c(_0814_)
    );

    and_bi _1516_ (
        .a(new_Jinkela_wire_6563),
        .b(new_Jinkela_wire_3942),
        .c(_0815_)
    );

    and_ii _1517_ (
        .a(new_Jinkela_wire_7963),
        .b(new_Jinkela_wire_4998),
        .c(_0816_)
    );

    or_ii _1518_ (
        .a(new_Jinkela_wire_6901),
        .b(new_Jinkela_wire_5801),
        .c(_0817_)
    );

    or_bb _1519_ (
        .a(new_Jinkela_wire_6902),
        .b(new_Jinkela_wire_5800),
        .c(_0818_)
    );

    or_ii _1520_ (
        .a(_0818_),
        .b(_0817_),
        .c(_0819_)
    );

    or_bb _1521_ (
        .a(new_Jinkela_wire_6934),
        .b(new_Jinkela_wire_1081),
        .c(_0820_)
    );

    inv _1522_ (
        .din(new_Jinkela_wire_508),
        .dout(_0821_)
    );

    or_bb _1523_ (
        .a(new_Jinkela_wire_156),
        .b(new_Jinkela_wire_326),
        .c(_0822_)
    );

    and_bi _1524_ (
        .a(new_Jinkela_wire_165),
        .b(new_Jinkela_wire_220),
        .c(_0823_)
    );

    and_bi _1525_ (
        .a(_0822_),
        .b(_0823_),
        .c(_0824_)
    );

    or_bb _1526_ (
        .a(_0824_),
        .b(new_Jinkela_wire_7009),
        .c(_0825_)
    );

    or_ii _1527_ (
        .a(new_Jinkela_wire_1578),
        .b(new_Jinkela_wire_153),
        .c(_0826_)
    );

    and_bi _1528_ (
        .a(new_Jinkela_wire_1291),
        .b(new_Jinkela_wire_161),
        .c(_0827_)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_2431),
        .dout(new_Jinkela_wire_2432)
    );

    bfr new_Jinkela_buffer_2023 (
        .din(new_Jinkela_wire_3123),
        .dout(new_Jinkela_wire_3124)
    );

    bfr new_Jinkela_buffer_3529 (
        .din(new_Jinkela_wire_4955),
        .dout(new_Jinkela_wire_4956)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_2374),
        .dout(new_Jinkela_wire_2375)
    );

    bfr new_Jinkela_buffer_2081 (
        .din(new_Jinkela_wire_3195),
        .dout(new_Jinkela_wire_3196)
    );

    bfr new_Jinkela_buffer_3582 (
        .din(new_Jinkela_wire_5032),
        .dout(new_Jinkela_wire_5033)
    );

    bfr new_Jinkela_buffer_3553 (
        .din(new_Jinkela_wire_4997),
        .dout(new_Jinkela_wire_4998)
    );

    bfr new_Jinkela_buffer_2024 (
        .din(new_Jinkela_wire_3124),
        .dout(new_Jinkela_wire_3125)
    );

    bfr new_Jinkela_buffer_3530 (
        .din(new_Jinkela_wire_4956),
        .dout(new_Jinkela_wire_4957)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(new_Jinkela_wire_2375),
        .dout(new_Jinkela_wire_2376)
    );

    bfr new_Jinkela_buffer_2045 (
        .din(new_Jinkela_wire_3145),
        .dout(new_Jinkela_wire_3146)
    );

    spl4L new_Jinkela_splitter_373 (
        .a(_0751_),
        .d(new_Jinkela_wire_2451),
        .e(new_Jinkela_wire_2452),
        .b(new_Jinkela_wire_2453),
        .c(new_Jinkela_wire_2454)
    );

    bfr new_Jinkela_buffer_2025 (
        .din(new_Jinkela_wire_3125),
        .dout(new_Jinkela_wire_3126)
    );

    bfr new_Jinkela_buffer_3531 (
        .din(new_Jinkela_wire_4957),
        .dout(new_Jinkela_wire_4958)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(new_Jinkela_wire_2376),
        .dout(new_Jinkela_wire_2377)
    );

    bfr new_Jinkela_buffer_2062 (
        .din(new_Jinkela_wire_3168),
        .dout(new_Jinkela_wire_3169)
    );

    bfr new_Jinkela_buffer_3557 (
        .din(new_Jinkela_wire_5007),
        .dout(new_Jinkela_wire_5008)
    );

    bfr new_Jinkela_buffer_2026 (
        .din(new_Jinkela_wire_3126),
        .dout(new_Jinkela_wire_3127)
    );

    bfr new_Jinkela_buffer_3532 (
        .din(new_Jinkela_wire_4958),
        .dout(new_Jinkela_wire_4959)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_2377),
        .dout(new_Jinkela_wire_2378)
    );

    bfr new_Jinkela_buffer_2046 (
        .din(new_Jinkela_wire_3146),
        .dout(new_Jinkela_wire_3147)
    );

    bfr new_Jinkela_buffer_3597 (
        .din(_0562_),
        .dout(new_Jinkela_wire_5056)
    );

    spl4L new_Jinkela_splitter_372 (
        .a(new_Jinkela_wire_2427),
        .d(new_Jinkela_wire_2428),
        .e(new_Jinkela_wire_2429),
        .b(new_Jinkela_wire_2430),
        .c(new_Jinkela_wire_2431)
    );

    bfr new_Jinkela_buffer_2027 (
        .din(new_Jinkela_wire_3127),
        .dout(new_Jinkela_wire_3128)
    );

    bfr new_Jinkela_buffer_3533 (
        .din(new_Jinkela_wire_4959),
        .dout(new_Jinkela_wire_4960)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_Jinkela_wire_2378),
        .dout(new_Jinkela_wire_2379)
    );

    bfr new_Jinkela_buffer_2064 (
        .din(new_Jinkela_wire_3175),
        .dout(new_Jinkela_wire_3176)
    );

    bfr new_Jinkela_buffer_3558 (
        .din(new_Jinkela_wire_5008),
        .dout(new_Jinkela_wire_5009)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(_0593_),
        .dout(new_Jinkela_wire_2455)
    );

    bfr new_Jinkela_buffer_2028 (
        .din(new_Jinkela_wire_3128),
        .dout(new_Jinkela_wire_3129)
    );

    bfr new_Jinkela_buffer_3534 (
        .din(new_Jinkela_wire_4960),
        .dout(new_Jinkela_wire_4961)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_2379),
        .dout(new_Jinkela_wire_2380)
    );

    bfr new_Jinkela_buffer_2047 (
        .din(new_Jinkela_wire_3147),
        .dout(new_Jinkela_wire_3148)
    );

    bfr new_Jinkela_buffer_3583 (
        .din(new_Jinkela_wire_5033),
        .dout(new_Jinkela_wire_5034)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_2425),
        .dout(new_Jinkela_wire_2426)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(_0448_),
        .dout(new_Jinkela_wire_2501)
    );

    bfr new_Jinkela_buffer_2029 (
        .din(new_Jinkela_wire_3129),
        .dout(new_Jinkela_wire_3130)
    );

    bfr new_Jinkela_buffer_3535 (
        .din(new_Jinkela_wire_4961),
        .dout(new_Jinkela_wire_4962)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_2380),
        .dout(new_Jinkela_wire_2381)
    );

    bfr new_Jinkela_buffer_2065 (
        .din(new_Jinkela_wire_3176),
        .dout(new_Jinkela_wire_3177)
    );

    bfr new_Jinkela_buffer_3559 (
        .din(new_Jinkela_wire_5009),
        .dout(new_Jinkela_wire_5010)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(new_Jinkela_wire_2455),
        .dout(new_Jinkela_wire_2456)
    );

    bfr new_Jinkela_buffer_2030 (
        .din(new_Jinkela_wire_3130),
        .dout(new_Jinkela_wire_3131)
    );

    bfr new_Jinkela_buffer_3536 (
        .din(new_Jinkela_wire_4962),
        .dout(new_Jinkela_wire_4963)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_2381),
        .dout(new_Jinkela_wire_2382)
    );

    bfr new_Jinkela_buffer_2048 (
        .din(new_Jinkela_wire_3148),
        .dout(new_Jinkela_wire_3149)
    );

    bfr new_Jinkela_buffer_3598 (
        .din(new_Jinkela_wire_5056),
        .dout(new_Jinkela_wire_5057)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_net_2441),
        .dout(new_Jinkela_wire_2461)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_2432),
        .dout(new_Jinkela_wire_2433)
    );

    bfr new_Jinkela_buffer_2031 (
        .din(new_Jinkela_wire_3131),
        .dout(new_Jinkela_wire_3132)
    );

    bfr new_Jinkela_buffer_3537 (
        .din(new_Jinkela_wire_4963),
        .dout(new_Jinkela_wire_4964)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_2382),
        .dout(new_Jinkela_wire_2383)
    );

    bfr new_Jinkela_buffer_2099 (
        .din(_0766_),
        .dout(new_Jinkela_wire_3214)
    );

    bfr new_Jinkela_buffer_3560 (
        .din(new_Jinkela_wire_5010),
        .dout(new_Jinkela_wire_5011)
    );

    bfr new_Jinkela_buffer_2100 (
        .din(_0095_),
        .dout(new_Jinkela_wire_3217)
    );

    bfr new_Jinkela_buffer_2032 (
        .din(new_Jinkela_wire_3132),
        .dout(new_Jinkela_wire_3133)
    );

    bfr new_Jinkela_buffer_3538 (
        .din(new_Jinkela_wire_4964),
        .dout(new_Jinkela_wire_4965)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_2383),
        .dout(new_Jinkela_wire_2384)
    );

    bfr new_Jinkela_buffer_2049 (
        .din(new_Jinkela_wire_3149),
        .dout(new_Jinkela_wire_3150)
    );

    bfr new_Jinkela_buffer_3584 (
        .din(new_Jinkela_wire_5034),
        .dout(new_Jinkela_wire_5035)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_2433),
        .dout(new_Jinkela_wire_2434)
    );

    bfr new_Jinkela_buffer_2033 (
        .din(new_Jinkela_wire_3133),
        .dout(new_Jinkela_wire_3134)
    );

    bfr new_Jinkela_buffer_3539 (
        .din(new_Jinkela_wire_4965),
        .dout(new_Jinkela_wire_4966)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(new_Jinkela_wire_2384),
        .dout(new_Jinkela_wire_2385)
    );

    bfr new_Jinkela_buffer_2066 (
        .din(new_Jinkela_wire_3177),
        .dout(new_Jinkela_wire_3178)
    );

    bfr new_Jinkela_buffer_3561 (
        .din(new_Jinkela_wire_5011),
        .dout(new_Jinkela_wire_5012)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(new_Jinkela_wire_2456),
        .dout(new_Jinkela_wire_2457)
    );

    bfr new_Jinkela_buffer_2034 (
        .din(new_Jinkela_wire_3134),
        .dout(new_Jinkela_wire_3135)
    );

    bfr new_Jinkela_buffer_3540 (
        .din(new_Jinkela_wire_4966),
        .dout(new_Jinkela_wire_4967)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_Jinkela_wire_2385),
        .dout(new_Jinkela_wire_2386)
    );

    bfr new_Jinkela_buffer_2050 (
        .din(new_Jinkela_wire_3150),
        .dout(new_Jinkela_wire_3151)
    );

    spl2 new_Jinkela_splitter_552 (
        .a(_0809_),
        .b(new_Jinkela_wire_5054),
        .c(new_Jinkela_wire_5055)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_2434),
        .dout(new_Jinkela_wire_2435)
    );

    bfr new_Jinkela_buffer_3541 (
        .din(new_Jinkela_wire_4967),
        .dout(new_Jinkela_wire_4968)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_2386),
        .dout(new_Jinkela_wire_2387)
    );

    bfr new_Jinkela_buffer_2051 (
        .din(new_Jinkela_wire_3151),
        .dout(new_Jinkela_wire_3152)
    );

    bfr new_Jinkela_buffer_3562 (
        .din(new_Jinkela_wire_5012),
        .dout(new_Jinkela_wire_5013)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(new_Jinkela_wire_2461),
        .dout(new_Jinkela_wire_2462)
    );

    bfr new_Jinkela_buffer_2067 (
        .din(new_Jinkela_wire_3178),
        .dout(new_Jinkela_wire_3179)
    );

    bfr new_Jinkela_buffer_3542 (
        .din(new_Jinkela_wire_4968),
        .dout(new_Jinkela_wire_4969)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_2387),
        .dout(new_Jinkela_wire_2388)
    );

    bfr new_Jinkela_buffer_2052 (
        .din(new_Jinkela_wire_3152),
        .dout(new_Jinkela_wire_3153)
    );

    bfr new_Jinkela_buffer_3585 (
        .din(new_Jinkela_wire_5035),
        .dout(new_Jinkela_wire_5036)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(new_Jinkela_wire_2435),
        .dout(new_Jinkela_wire_2436)
    );

    bfr new_Jinkela_buffer_2089 (
        .din(new_Jinkela_wire_3203),
        .dout(new_Jinkela_wire_3204)
    );

    bfr new_Jinkela_buffer_3543 (
        .din(new_Jinkela_wire_4969),
        .dout(new_Jinkela_wire_4970)
    );

    bfr new_Jinkela_buffer_2082 (
        .din(new_Jinkela_wire_3196),
        .dout(new_Jinkela_wire_3197)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_2388),
        .dout(new_Jinkela_wire_2389)
    );

    bfr new_Jinkela_buffer_2053 (
        .din(new_Jinkela_wire_3153),
        .dout(new_Jinkela_wire_3154)
    );

    bfr new_Jinkela_buffer_3563 (
        .din(new_Jinkela_wire_5013),
        .dout(new_Jinkela_wire_5014)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_2457),
        .dout(new_Jinkela_wire_2458)
    );

    bfr new_Jinkela_buffer_2068 (
        .din(new_Jinkela_wire_3179),
        .dout(new_Jinkela_wire_3180)
    );

    bfr new_Jinkela_buffer_3544 (
        .din(new_Jinkela_wire_4970),
        .dout(new_Jinkela_wire_4971)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_2389),
        .dout(new_Jinkela_wire_2390)
    );

    bfr new_Jinkela_buffer_2054 (
        .din(new_Jinkela_wire_3154),
        .dout(new_Jinkela_wire_3155)
    );

    bfr new_Jinkela_buffer_3622 (
        .din(_0107_),
        .dout(new_Jinkela_wire_5081)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_2436),
        .dout(new_Jinkela_wire_2437)
    );

    bfr new_Jinkela_buffer_3545 (
        .din(new_Jinkela_wire_4971),
        .dout(new_Jinkela_wire_4972)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_2390),
        .dout(new_Jinkela_wire_2391)
    );

    bfr new_Jinkela_buffer_2055 (
        .din(new_Jinkela_wire_3155),
        .dout(new_Jinkela_wire_3156)
    );

    bfr new_Jinkela_buffer_3564 (
        .din(new_Jinkela_wire_5014),
        .dout(new_Jinkela_wire_5015)
    );

    spl2 new_Jinkela_splitter_374 (
        .a(_0114_),
        .b(new_Jinkela_wire_2532),
        .c(new_Jinkela_wire_2533)
    );

    bfr new_Jinkela_buffer_2069 (
        .din(new_Jinkela_wire_3180),
        .dout(new_Jinkela_wire_3181)
    );

    bfr new_Jinkela_buffer_3546 (
        .din(new_Jinkela_wire_4972),
        .dout(new_Jinkela_wire_4973)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(new_Jinkela_wire_2391),
        .dout(new_Jinkela_wire_2392)
    );

    bfr new_Jinkela_buffer_2056 (
        .din(new_Jinkela_wire_3156),
        .dout(new_Jinkela_wire_3157)
    );

    bfr new_Jinkela_buffer_3586 (
        .din(new_Jinkela_wire_5036),
        .dout(new_Jinkela_wire_5037)
    );

    spl2 new_Jinkela_splitter_375 (
        .a(_1032_),
        .b(new_Jinkela_wire_2534),
        .c(new_Jinkela_wire_2535)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_2437),
        .dout(new_Jinkela_wire_2438)
    );

    bfr new_Jinkela_buffer_3565 (
        .din(new_Jinkela_wire_5015),
        .dout(new_Jinkela_wire_5016)
    );

    bfr new_Jinkela_buffer_2083 (
        .din(new_Jinkela_wire_3197),
        .dout(new_Jinkela_wire_3198)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(new_Jinkela_wire_2392),
        .dout(new_Jinkela_wire_2393)
    );

    bfr new_Jinkela_buffer_2057 (
        .din(new_Jinkela_wire_3157),
        .dout(new_Jinkela_wire_3158)
    );

    spl2 new_Jinkela_splitter_553 (
        .a(_0764_),
        .b(new_Jinkela_wire_5114),
        .c(new_Jinkela_wire_5115)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_2458),
        .dout(new_Jinkela_wire_2459)
    );

    bfr new_Jinkela_buffer_2070 (
        .din(new_Jinkela_wire_3181),
        .dout(new_Jinkela_wire_3182)
    );

    bfr new_Jinkela_buffer_3566 (
        .din(new_Jinkela_wire_5016),
        .dout(new_Jinkela_wire_5017)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_2393),
        .dout(new_Jinkela_wire_2394)
    );

    bfr new_Jinkela_buffer_2058 (
        .din(new_Jinkela_wire_3158),
        .dout(new_Jinkela_wire_3159)
    );

    bfr new_Jinkela_buffer_3587 (
        .din(new_Jinkela_wire_5037),
        .dout(new_Jinkela_wire_5038)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(new_Jinkela_wire_2438),
        .dout(new_Jinkela_wire_2439)
    );

    bfr new_Jinkela_buffer_3567 (
        .din(new_Jinkela_wire_5017),
        .dout(new_Jinkela_wire_5018)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_2394),
        .dout(new_Jinkela_wire_2395)
    );

    bfr new_Jinkela_buffer_2071 (
        .din(new_Jinkela_wire_3182),
        .dout(new_Jinkela_wire_3183)
    );

    bfr new_Jinkela_buffer_3599 (
        .din(new_Jinkela_wire_5057),
        .dout(new_Jinkela_wire_5058)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_1237),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_2553 (
        .din(new_Jinkela_wire_3812),
        .dout(new_Jinkela_wire_3813)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_1174),
        .dout(new_Jinkela_wire_1175)
    );

    bfr new_Jinkela_buffer_2565 (
        .din(new_Jinkela_wire_3828),
        .dout(new_Jinkela_wire_3829)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(new_Jinkela_wire_1229),
        .b(new_Jinkela_wire_1230),
        .c(new_Jinkela_wire_1231)
    );

    bfr new_Jinkela_buffer_2554 (
        .din(new_Jinkela_wire_3813),
        .dout(new_Jinkela_wire_3814)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_1175),
        .dout(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_2572 (
        .din(new_Jinkela_wire_3839),
        .dout(new_Jinkela_wire_3840)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_1231),
        .dout(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_2555 (
        .din(new_Jinkela_wire_3814),
        .dout(new_Jinkela_wire_3815)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_1176),
        .dout(new_Jinkela_wire_1177)
    );

    bfr new_Jinkela_buffer_2620 (
        .din(new_net_2481),
        .dout(new_Jinkela_wire_3890)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_1239),
        .dout(new_Jinkela_wire_1240)
    );

    bfr new_Jinkela_buffer_2556 (
        .din(new_Jinkela_wire_3815),
        .dout(new_Jinkela_wire_3816)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_1177),
        .dout(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_2566 (
        .din(new_Jinkela_wire_3829),
        .dout(new_Jinkela_wire_3830)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(G141),
        .b(new_Jinkela_wire_1251),
        .c(new_Jinkela_wire_1252)
    );

    bfr new_Jinkela_buffer_2557 (
        .din(new_Jinkela_wire_3816),
        .dout(new_Jinkela_wire_3817)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_1178),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_2573 (
        .din(new_Jinkela_wire_3840),
        .dout(new_Jinkela_wire_3841)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(new_Jinkela_wire_1232),
        .b(new_Jinkela_wire_1233),
        .c(new_Jinkela_wire_1234)
    );

    bfr new_Jinkela_buffer_2558 (
        .din(new_Jinkela_wire_3817),
        .dout(new_Jinkela_wire_3818)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_1179),
        .dout(new_Jinkela_wire_1180)
    );

    bfr new_Jinkela_buffer_2567 (
        .din(new_Jinkela_wire_3830),
        .dout(new_Jinkela_wire_3831)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    bfr new_Jinkela_buffer_2559 (
        .din(new_Jinkela_wire_3818),
        .dout(new_Jinkela_wire_3819)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_2619 (
        .din(new_Jinkela_wire_3888),
        .dout(new_Jinkela_wire_3889)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_1240),
        .dout(new_Jinkela_wire_1241)
    );

    bfr new_Jinkela_buffer_2610 (
        .din(new_Jinkela_wire_3879),
        .dout(new_Jinkela_wire_3880)
    );

    bfr new_Jinkela_buffer_2568 (
        .din(new_Jinkela_wire_3831),
        .dout(new_Jinkela_wire_3832)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_1181),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_2574 (
        .din(new_Jinkela_wire_3841),
        .dout(new_Jinkela_wire_3842)
    );

    spl2 new_Jinkela_splitter_226 (
        .a(new_Jinkela_wire_1241),
        .b(new_Jinkela_wire_1242),
        .c(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_1182),
        .dout(new_Jinkela_wire_1183)
    );

    bfr new_Jinkela_buffer_2575 (
        .din(new_Jinkela_wire_3842),
        .dout(new_Jinkela_wire_3843)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_2632 (
        .din(new_net_2375),
        .dout(new_Jinkela_wire_3902)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_1183),
        .dout(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_2611 (
        .din(new_Jinkela_wire_3880),
        .dout(new_Jinkela_wire_3881)
    );

    bfr new_Jinkela_buffer_2576 (
        .din(new_Jinkela_wire_3843),
        .dout(new_Jinkela_wire_3844)
    );

    spl3L new_Jinkela_splitter_230 (
        .a(G172),
        .d(new_Jinkela_wire_1259),
        .b(new_Jinkela_wire_1260),
        .c(new_Jinkela_wire_1261)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_1184),
        .dout(new_Jinkela_wire_1185)
    );

    bfr new_Jinkela_buffer_2577 (
        .din(new_Jinkela_wire_3844),
        .dout(new_Jinkela_wire_3845)
    );

    bfr new_Jinkela_buffer_2621 (
        .din(new_Jinkela_wire_3890),
        .dout(new_Jinkela_wire_3891)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_1185),
        .dout(new_Jinkela_wire_1186)
    );

    bfr new_Jinkela_buffer_2612 (
        .din(new_Jinkela_wire_3881),
        .dout(new_Jinkela_wire_3882)
    );

    bfr new_Jinkela_buffer_2578 (
        .din(new_Jinkela_wire_3845),
        .dout(new_Jinkela_wire_3846)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(new_Jinkela_wire_1246),
        .b(new_Jinkela_wire_1247),
        .c(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_1186),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_2579 (
        .din(new_Jinkela_wire_3846),
        .dout(new_Jinkela_wire_3847)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_1252),
        .dout(new_Jinkela_wire_1253)
    );

    spl2 new_Jinkela_splitter_479 (
        .a(_0814_),
        .b(new_Jinkela_wire_3942),
        .c(new_Jinkela_wire_3943)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_1187),
        .dout(new_Jinkela_wire_1188)
    );

    bfr new_Jinkela_buffer_2613 (
        .din(new_Jinkela_wire_3882),
        .dout(new_Jinkela_wire_3883)
    );

    bfr new_Jinkela_buffer_2580 (
        .din(new_Jinkela_wire_3847),
        .dout(new_Jinkela_wire_3848)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_1253),
        .dout(new_Jinkela_wire_1254)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_1188),
        .dout(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_2672 (
        .din(_0262_),
        .dout(new_Jinkela_wire_3944)
    );

    bfr new_Jinkela_buffer_2581 (
        .din(new_Jinkela_wire_3848),
        .dout(new_Jinkela_wire_3849)
    );

    bfr new_Jinkela_buffer_618 (
        .din(G49),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_626 (
        .din(G84),
        .dout(new_Jinkela_wire_1272)
    );

    bfr new_Jinkela_buffer_2622 (
        .din(new_Jinkela_wire_3891),
        .dout(new_Jinkela_wire_3892)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_2614 (
        .din(new_Jinkela_wire_3883),
        .dout(new_Jinkela_wire_3884)
    );

    bfr new_Jinkela_buffer_2582 (
        .din(new_Jinkela_wire_3849),
        .dout(new_Jinkela_wire_3850)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_1254),
        .dout(new_Jinkela_wire_1255)
    );

    bfr new_Jinkela_buffer_2583 (
        .din(new_Jinkela_wire_3850),
        .dout(new_Jinkela_wire_3851)
    );

    bfr new_Jinkela_buffer_2633 (
        .din(new_Jinkela_wire_3902),
        .dout(new_Jinkela_wire_3903)
    );

    bfr new_Jinkela_buffer_623 (
        .din(G41),
        .dout(new_Jinkela_wire_1267)
    );

    bfr new_Jinkela_buffer_2615 (
        .din(new_Jinkela_wire_3884),
        .dout(new_Jinkela_wire_3885)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_1255),
        .dout(new_Jinkela_wire_1256)
    );

    bfr new_Jinkela_buffer_2584 (
        .din(new_Jinkela_wire_3851),
        .dout(new_Jinkela_wire_3852)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    spl2 new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_1256),
        .b(new_Jinkela_wire_1257),
        .c(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_2585 (
        .din(new_Jinkela_wire_3852),
        .dout(new_Jinkela_wire_3853)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_1264),
        .dout(new_Jinkela_wire_1265)
    );

    bfr new_Jinkela_buffer_2623 (
        .din(new_Jinkela_wire_3892),
        .dout(new_Jinkela_wire_3893)
    );

    bfr new_Jinkela_buffer_2616 (
        .din(new_Jinkela_wire_3885),
        .dout(new_Jinkela_wire_3886)
    );

    spl2 new_Jinkela_splitter_233 (
        .a(G166),
        .b(new_Jinkela_wire_1277),
        .c(new_Jinkela_wire_1280)
    );

    bfr new_Jinkela_buffer_2586 (
        .din(new_Jinkela_wire_3853),
        .dout(new_Jinkela_wire_3854)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_1267),
        .dout(new_Jinkela_wire_1268)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_1265),
        .dout(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_2587 (
        .din(new_Jinkela_wire_3854),
        .dout(new_Jinkela_wire_3855)
    );

    or_bb _2325_ (
        .a(new_Jinkela_wire_1708),
        .b(_0332_),
        .c(new_net_2473)
    );

    or_bi _2326_ (
        .a(new_Jinkela_wire_379),
        .b(new_Jinkela_wire_5879),
        .c(_0336_)
    );

    spl2 new_Jinkela_splitter_534 (
        .a(new_Jinkela_wire_4825),
        .b(new_Jinkela_wire_4826),
        .c(new_Jinkela_wire_4827)
    );

    spl4L new_Jinkela_splitter_535 (
        .a(new_Jinkela_wire_4828),
        .d(new_Jinkela_wire_4829),
        .e(new_Jinkela_wire_4830),
        .b(new_Jinkela_wire_4835),
        .c(new_Jinkela_wire_4840)
    );

    spl4L new_Jinkela_splitter_536 (
        .a(new_Jinkela_wire_4830),
        .d(new_Jinkela_wire_4831),
        .e(new_Jinkela_wire_4832),
        .b(new_Jinkela_wire_4833),
        .c(new_Jinkela_wire_4834)
    );

    bfr new_Jinkela_buffer_3438 (
        .din(new_Jinkela_wire_4860),
        .dout(new_Jinkela_wire_4861)
    );

    spl4L new_Jinkela_splitter_537 (
        .a(new_Jinkela_wire_4835),
        .d(new_Jinkela_wire_4836),
        .e(new_Jinkela_wire_4837),
        .b(new_Jinkela_wire_4838),
        .c(new_Jinkela_wire_4839)
    );

    bfr new_Jinkela_buffer_3424 (
        .din(new_Jinkela_wire_4844),
        .dout(new_Jinkela_wire_4845)
    );

    spl4L new_Jinkela_splitter_538 (
        .a(new_Jinkela_wire_4840),
        .d(new_Jinkela_wire_4841),
        .e(new_Jinkela_wire_4842),
        .b(new_Jinkela_wire_4843),
        .c(new_Jinkela_wire_4844)
    );

    bfr new_Jinkela_buffer_3444 (
        .din(new_Jinkela_wire_4866),
        .dout(new_Jinkela_wire_4867)
    );

    bfr new_Jinkela_buffer_3439 (
        .din(new_Jinkela_wire_4861),
        .dout(new_Jinkela_wire_4862)
    );

    bfr new_Jinkela_buffer_3446 (
        .din(new_Jinkela_wire_4868),
        .dout(new_Jinkela_wire_4869)
    );

    bfr new_Jinkela_buffer_3425 (
        .din(new_Jinkela_wire_4845),
        .dout(new_Jinkela_wire_4846)
    );

    bfr new_Jinkela_buffer_3440 (
        .din(new_Jinkela_wire_4862),
        .dout(new_Jinkela_wire_4863)
    );

    bfr new_Jinkela_buffer_3426 (
        .din(new_Jinkela_wire_4846),
        .dout(new_Jinkela_wire_4847)
    );

    bfr new_Jinkela_buffer_3477 (
        .din(_0926_),
        .dout(new_Jinkela_wire_4900)
    );

    bfr new_Jinkela_buffer_3427 (
        .din(new_Jinkela_wire_4847),
        .dout(new_Jinkela_wire_4848)
    );

    bfr new_Jinkela_buffer_3441 (
        .din(new_Jinkela_wire_4863),
        .dout(new_Jinkela_wire_4864)
    );

    bfr new_Jinkela_buffer_3428 (
        .din(new_Jinkela_wire_4848),
        .dout(new_Jinkela_wire_4849)
    );

    bfr new_Jinkela_buffer_3447 (
        .din(new_Jinkela_wire_4869),
        .dout(new_Jinkela_wire_4870)
    );

    bfr new_Jinkela_buffer_3429 (
        .din(new_Jinkela_wire_4849),
        .dout(new_Jinkela_wire_4850)
    );

    bfr new_Jinkela_buffer_3465 (
        .din(new_Jinkela_wire_4887),
        .dout(new_Jinkela_wire_4888)
    );

    bfr new_Jinkela_buffer_3430 (
        .din(new_Jinkela_wire_4850),
        .dout(new_Jinkela_wire_4851)
    );

    bfr new_Jinkela_buffer_3448 (
        .din(new_Jinkela_wire_4870),
        .dout(new_Jinkela_wire_4871)
    );

    bfr new_Jinkela_buffer_3431 (
        .din(new_Jinkela_wire_4851),
        .dout(new_Jinkela_wire_4852)
    );

    spl4L new_Jinkela_splitter_540 (
        .a(_0612_),
        .d(new_Jinkela_wire_4917),
        .e(new_Jinkela_wire_4918),
        .b(new_Jinkela_wire_4919),
        .c(new_Jinkela_wire_4920)
    );

    bfr new_Jinkela_buffer_3494 (
        .din(_0280_),
        .dout(new_Jinkela_wire_4921)
    );

    spl2 new_Jinkela_splitter_539 (
        .a(new_Jinkela_wire_4852),
        .b(new_Jinkela_wire_4853),
        .c(new_Jinkela_wire_4854)
    );

    bfr new_Jinkela_buffer_3432 (
        .din(new_Jinkela_wire_4854),
        .dout(new_Jinkela_wire_4855)
    );

    bfr new_Jinkela_buffer_3449 (
        .din(new_Jinkela_wire_4871),
        .dout(new_Jinkela_wire_4872)
    );

    bfr new_Jinkela_buffer_3466 (
        .din(new_Jinkela_wire_4888),
        .dout(new_Jinkela_wire_4889)
    );

    bfr new_Jinkela_buffer_3433 (
        .din(new_Jinkela_wire_4855),
        .dout(new_Jinkela_wire_4856)
    );

    bfr new_Jinkela_buffer_3450 (
        .din(new_Jinkela_wire_4872),
        .dout(new_Jinkela_wire_4873)
    );

    bfr new_Jinkela_buffer_3478 (
        .din(new_Jinkela_wire_4900),
        .dout(new_Jinkela_wire_4901)
    );

    bfr new_Jinkela_buffer_3451 (
        .din(new_Jinkela_wire_4873),
        .dout(new_Jinkela_wire_4874)
    );

    bfr new_Jinkela_buffer_3467 (
        .din(new_Jinkela_wire_4889),
        .dout(new_Jinkela_wire_4890)
    );

    bfr new_Jinkela_buffer_3452 (
        .din(new_Jinkela_wire_4874),
        .dout(new_Jinkela_wire_4875)
    );

    bfr new_Jinkela_buffer_3453 (
        .din(new_Jinkela_wire_4875),
        .dout(new_Jinkela_wire_4876)
    );

    bfr new_Jinkela_buffer_3468 (
        .din(new_Jinkela_wire_4890),
        .dout(new_Jinkela_wire_4891)
    );

    bfr new_Jinkela_buffer_3454 (
        .din(new_Jinkela_wire_4876),
        .dout(new_Jinkela_wire_4877)
    );

    bfr new_Jinkela_buffer_3479 (
        .din(new_Jinkela_wire_4901),
        .dout(new_Jinkela_wire_4902)
    );

    bfr new_Jinkela_buffer_3455 (
        .din(new_Jinkela_wire_4877),
        .dout(new_Jinkela_wire_4878)
    );

    bfr new_Jinkela_buffer_3469 (
        .din(new_Jinkela_wire_4891),
        .dout(new_Jinkela_wire_4892)
    );

    bfr new_Jinkela_buffer_3456 (
        .din(new_Jinkela_wire_4878),
        .dout(new_Jinkela_wire_4879)
    );

    spl4L new_Jinkela_splitter_216 (
        .a(new_Jinkela_wire_1198),
        .d(new_Jinkela_wire_1199),
        .e(new_Jinkela_wire_1200),
        .b(new_Jinkela_wire_1205),
        .c(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_1215),
        .dout(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_2462),
        .dout(new_Jinkela_wire_2463)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_1153),
        .dout(new_Jinkela_wire_1154)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_2395),
        .dout(new_Jinkela_wire_2396)
    );

    spl2 new_Jinkela_splitter_213 (
        .a(new_Jinkela_wire_1192),
        .b(new_Jinkela_wire_1193),
        .c(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(new_Jinkela_wire_2439),
        .dout(new_Jinkela_wire_2440)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_1154),
        .dout(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(new_Jinkela_wire_2459),
        .dout(new_Jinkela_wire_2460)
    );

    spl4L new_Jinkela_splitter_217 (
        .a(new_Jinkela_wire_1200),
        .d(new_Jinkela_wire_1201),
        .e(new_Jinkela_wire_1202),
        .b(new_Jinkela_wire_1203),
        .c(new_Jinkela_wire_1204)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(new_Jinkela_wire_2440),
        .dout(new_Jinkela_wire_2441)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_1155),
        .dout(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(new_Jinkela_wire_2501),
        .dout(new_Jinkela_wire_2502)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(new_Jinkela_wire_2441),
        .dout(new_Jinkela_wire_2442)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_1156),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(new_Jinkela_wire_2463),
        .dout(new_Jinkela_wire_2464)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_2442),
        .dout(new_Jinkela_wire_2443)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    spl2 new_Jinkela_splitter_222 (
        .a(G147),
        .b(new_Jinkela_wire_1225),
        .c(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(new_Jinkela_wire_2443),
        .dout(new_Jinkela_wire_2444)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(new_Jinkela_wire_2464),
        .dout(new_Jinkela_wire_2465)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(new_Jinkela_wire_1195),
        .b(new_Jinkela_wire_1196),
        .c(new_Jinkela_wire_1197)
    );

    spl4L new_Jinkela_splitter_218 (
        .a(new_Jinkela_wire_1205),
        .d(new_Jinkela_wire_1206),
        .e(new_Jinkela_wire_1207),
        .b(new_Jinkela_wire_1208),
        .c(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_2444),
        .dout(new_Jinkela_wire_2445)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_1159),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_Jinkela_wire_2502),
        .dout(new_Jinkela_wire_2503)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(new_Jinkela_wire_1217),
        .b(new_Jinkela_wire_1218),
        .c(new_Jinkela_wire_1219)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_Jinkela_wire_2445),
        .dout(new_Jinkela_wire_2446)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(new_Jinkela_wire_2465),
        .dout(new_Jinkela_wire_2466)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_1236),
        .dout(new_Jinkela_wire_1237)
    );

    spl4L new_Jinkela_splitter_219 (
        .a(new_Jinkela_wire_1210),
        .d(new_Jinkela_wire_1211),
        .e(new_Jinkela_wire_1212),
        .b(new_Jinkela_wire_1213),
        .c(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_2446),
        .dout(new_Jinkela_wire_2447)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    spl2 new_Jinkela_splitter_376 (
        .a(_0031_),
        .b(new_Jinkela_wire_2536),
        .c(new_Jinkela_wire_2537)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(new_Jinkela_wire_2447),
        .dout(new_Jinkela_wire_2448)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_Jinkela_wire_2466),
        .dout(new_Jinkela_wire_2467)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(new_Jinkela_wire_2448),
        .dout(new_Jinkela_wire_2449)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_1163),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_2503),
        .dout(new_Jinkela_wire_2504)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(new_Jinkela_wire_2449),
        .dout(new_Jinkela_wire_2450)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_1164),
        .dout(new_Jinkela_wire_1165)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(new_Jinkela_wire_2467),
        .dout(new_Jinkela_wire_2468)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    spl2 new_Jinkela_splitter_377 (
        .a(_0874_),
        .b(new_Jinkela_wire_2570),
        .c(new_Jinkela_wire_2571)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_1165),
        .dout(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(_0750_),
        .dout(new_Jinkela_wire_2538)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(new_Jinkela_wire_2468),
        .dout(new_Jinkela_wire_2469)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_2504),
        .dout(new_Jinkela_wire_2505)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_1166),
        .dout(new_Jinkela_wire_1167)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_2469),
        .dout(new_Jinkela_wire_2470)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_1226),
        .dout(new_Jinkela_wire_1227)
    );

    bfr new_Jinkela_buffer_606 (
        .din(G15),
        .dout(new_Jinkela_wire_1239)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_1167),
        .dout(new_Jinkela_wire_1168)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(new_Jinkela_wire_2470),
        .dout(new_Jinkela_wire_2471)
    );

    spl2 new_Jinkela_splitter_221 (
        .a(new_Jinkela_wire_1222),
        .b(new_Jinkela_wire_1223),
        .c(new_Jinkela_wire_1224)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_2505),
        .dout(new_Jinkela_wire_2506)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_1168),
        .dout(new_Jinkela_wire_1169)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(new_Jinkela_wire_2471),
        .dout(new_Jinkela_wire_2472)
    );

    bfr new_Jinkela_buffer_609 (
        .din(G24),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_612 (
        .din(G31),
        .dout(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(_0528_),
        .dout(new_Jinkela_wire_2539)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_1169),
        .dout(new_Jinkela_wire_1170)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_net_2419),
        .dout(new_Jinkela_wire_2582)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_2472),
        .dout(new_Jinkela_wire_2473)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(new_Jinkela_wire_2506),
        .dout(new_Jinkela_wire_2507)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_1170),
        .dout(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(new_Jinkela_wire_2473),
        .dout(new_Jinkela_wire_2474)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_1227),
        .dout(new_Jinkela_wire_1228)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(new_Jinkela_wire_2539),
        .dout(new_Jinkela_wire_2540)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_1171),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(new_Jinkela_wire_2474),
        .dout(new_Jinkela_wire_2475)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(G129),
        .b(new_Jinkela_wire_1235),
        .c(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_1228),
        .dout(new_Jinkela_wire_1229)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(new_Jinkela_wire_2507),
        .dout(new_Jinkela_wire_2508)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_1172),
        .dout(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(new_Jinkela_wire_2475),
        .dout(new_Jinkela_wire_2476)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(new_Jinkela_wire_2571),
        .dout(new_Jinkela_wire_2572)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_1173),
        .dout(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_2476),
        .dout(new_Jinkela_wire_2477)
    );

    and_bi _1529_ (
        .a(new_Jinkela_wire_7995),
        .b(_0827_),
        .c(_0828_)
    );

    and_bb _2243_ (
        .a(new_Jinkela_wire_4378),
        .b(new_Jinkela_wire_358),
        .c(_0263_)
    );

    bfr new_Jinkela_buffer_2521 (
        .din(new_Jinkela_wire_3780),
        .dout(new_Jinkela_wire_3781)
    );

    and_bi _1530_ (
        .a(new_Jinkela_wire_7010),
        .b(_0828_),
        .c(_0829_)
    );

    or_bb _2244_ (
        .a(_0263_),
        .b(new_Jinkela_wire_3957),
        .c(_0264_)
    );

    bfr new_Jinkela_buffer_2541 (
        .din(new_Jinkela_wire_3800),
        .dout(new_Jinkela_wire_3801)
    );

    and_bi _1531_ (
        .a(_0825_),
        .b(_0829_),
        .c(_0830_)
    );

    and_bi _2245_ (
        .a(_0261_),
        .b(new_Jinkela_wire_7464),
        .c(_0265_)
    );

    bfr new_Jinkela_buffer_2522 (
        .din(new_Jinkela_wire_3781),
        .dout(new_Jinkela_wire_3782)
    );

    and_bi _1532_ (
        .a(new_Jinkela_wire_1058),
        .b(new_Jinkela_wire_5243),
        .c(_0831_)
    );

    or_bi _2246_ (
        .a(new_Jinkela_wire_1592),
        .b(new_Jinkela_wire_342),
        .c(_0266_)
    );

    bfr new_Jinkela_buffer_2560 (
        .din(new_Jinkela_wire_3821),
        .dout(new_Jinkela_wire_3822)
    );

    or_bb _1533_ (
        .a(_0831_),
        .b(new_Jinkela_wire_4839),
        .c(_0832_)
    );

    and_bi _2247_ (
        .a(new_Jinkela_wire_232),
        .b(new_Jinkela_wire_5812),
        .c(_0267_)
    );

    bfr new_Jinkela_buffer_2523 (
        .din(new_Jinkela_wire_3782),
        .dout(new_Jinkela_wire_3783)
    );

    and_bi _1534_ (
        .a(_0820_),
        .b(new_Jinkela_wire_3766),
        .c(_0833_)
    );

    or_bb _2248_ (
        .a(new_Jinkela_wire_1594),
        .b(new_Jinkela_wire_343),
        .c(_0268_)
    );

    bfr new_Jinkela_buffer_2542 (
        .din(new_Jinkela_wire_3801),
        .dout(new_Jinkela_wire_3802)
    );

    and_ii _1535_ (
        .a(_0833_),
        .b(new_Jinkela_wire_7911),
        .c(new_net_9)
    );

    and_bi _2249_ (
        .a(new_Jinkela_wire_1493),
        .b(new_Jinkela_wire_7869),
        .c(_0269_)
    );

    bfr new_Jinkela_buffer_2524 (
        .din(new_Jinkela_wire_3783),
        .dout(new_Jinkela_wire_3784)
    );

    and_bi _1536_ (
        .a(new_Jinkela_wire_87),
        .b(new_Jinkela_wire_6704),
        .c(_0834_)
    );

    or_bb _2250_ (
        .a(_0269_),
        .b(_0267_),
        .c(_0270_)
    );

    bfr new_Jinkela_buffer_2618 (
        .din(_0279_),
        .dout(new_Jinkela_wire_3888)
    );

    and_bi _1537_ (
        .a(new_Jinkela_wire_3943),
        .b(new_Jinkela_wire_6562),
        .c(_0835_)
    );

    or_bb _2251_ (
        .a(new_Jinkela_wire_4128),
        .b(_0265_),
        .c(new_net_2451)
    );

    bfr new_Jinkela_buffer_2525 (
        .din(new_Jinkela_wire_3784),
        .dout(new_Jinkela_wire_3785)
    );

    or_bb _1538_ (
        .a(new_Jinkela_wire_2265),
        .b(new_Jinkela_wire_7961),
        .c(_0836_)
    );

    or_bb _2252_ (
        .a(new_Jinkela_wire_2925),
        .b(new_Jinkela_wire_4611),
        .c(_0271_)
    );

    bfr new_Jinkela_buffer_2543 (
        .din(new_Jinkela_wire_3802),
        .dout(new_Jinkela_wire_3803)
    );

    or_bb _1539_ (
        .a(new_Jinkela_wire_2924),
        .b(new_Jinkela_wire_1073),
        .c(_0837_)
    );

    or_bb _2253_ (
        .a(new_Jinkela_wire_5215),
        .b(new_Jinkela_wire_5272),
        .c(_0272_)
    );

    bfr new_Jinkela_buffer_2526 (
        .din(new_Jinkela_wire_3785),
        .dout(new_Jinkela_wire_3786)
    );

    or_bb _1540_ (
        .a(new_Jinkela_wire_1311),
        .b(new_Jinkela_wire_320),
        .c(_0838_)
    );

    or_bb _2254_ (
        .a(_0272_),
        .b(new_Jinkela_wire_6936),
        .c(_0273_)
    );

    and_bi _1541_ (
        .a(new_Jinkela_wire_1319),
        .b(new_Jinkela_wire_215),
        .c(_0839_)
    );

    or_bb _2255_ (
        .a(_0273_),
        .b(new_Jinkela_wire_5235),
        .c(_0274_)
    );

    bfr new_Jinkela_buffer_2527 (
        .din(new_Jinkela_wire_3786),
        .dout(new_Jinkela_wire_3787)
    );

    and_bi _1542_ (
        .a(_0838_),
        .b(_0839_),
        .c(_0840_)
    );

    or_bb _2256_ (
        .a(new_Jinkela_wire_5333),
        .b(new_Jinkela_wire_2535),
        .c(_0275_)
    );

    bfr new_Jinkela_buffer_2544 (
        .din(new_Jinkela_wire_3803),
        .dout(new_Jinkela_wire_3804)
    );

    or_bb _1543_ (
        .a(_0840_),
        .b(new_Jinkela_wire_5698),
        .c(_0841_)
    );

    and_bi _2257_ (
        .a(new_Jinkela_wire_7106),
        .b(new_Jinkela_wire_5120),
        .c(_0276_)
    );

    bfr new_Jinkela_buffer_2528 (
        .din(new_Jinkela_wire_3787),
        .dout(new_Jinkela_wire_3788)
    );

    or_ii _1544_ (
        .a(new_Jinkela_wire_1590),
        .b(new_Jinkela_wire_1316),
        .c(_0842_)
    );

    or_bb _2258_ (
        .a(new_Jinkela_wire_6251),
        .b(new_Jinkela_wire_4412),
        .c(_0277_)
    );

    bfr new_Jinkela_buffer_2561 (
        .din(new_Jinkela_wire_3822),
        .dout(new_Jinkela_wire_3823)
    );

    and_bi _1545_ (
        .a(new_Jinkela_wire_1293),
        .b(new_Jinkela_wire_1309),
        .c(_0843_)
    );

    and_bi _2259_ (
        .a(_0276_),
        .b(_0277_),
        .c(new_net_2417)
    );

    bfr new_Jinkela_buffer_2529 (
        .din(new_Jinkela_wire_3788),
        .dout(new_Jinkela_wire_3789)
    );

    and_bi _1546_ (
        .a(_0842_),
        .b(_0843_),
        .c(_0844_)
    );

    or_bi _2260_ (
        .a(new_Jinkela_wire_6228),
        .b(new_Jinkela_wire_7786),
        .c(_0278_)
    );

    bfr new_Jinkela_buffer_2545 (
        .din(new_Jinkela_wire_3804),
        .dout(new_Jinkela_wire_3805)
    );

    and_bi _1547_ (
        .a(new_Jinkela_wire_5701),
        .b(_0844_),
        .c(_0845_)
    );

    or_bb _2261_ (
        .a(new_Jinkela_wire_6711),
        .b(new_Jinkela_wire_4344),
        .c(_0279_)
    );

    bfr new_Jinkela_buffer_2530 (
        .din(new_Jinkela_wire_3789),
        .dout(new_Jinkela_wire_3790)
    );

    and_bi _1548_ (
        .a(_0841_),
        .b(_0845_),
        .c(_0846_)
    );

    or_bb _2262_ (
        .a(new_Jinkela_wire_3889),
        .b(new_Jinkela_wire_1859),
        .c(_0280_)
    );

    bfr new_Jinkela_buffer_2609 (
        .din(new_Jinkela_wire_3878),
        .dout(new_Jinkela_wire_3879)
    );

    spl2 new_Jinkela_splitter_478 (
        .a(_0957_),
        .b(new_Jinkela_wire_3877),
        .c(new_Jinkela_wire_3878)
    );

    or_bb _2263_ (
        .a(new_Jinkela_wire_4921),
        .b(new_Jinkela_wire_5053),
        .c(_0281_)
    );

    and_bi _1549_ (
        .a(new_Jinkela_wire_1059),
        .b(new_Jinkela_wire_2307),
        .c(_0847_)
    );

    bfr new_Jinkela_buffer_2531 (
        .din(new_Jinkela_wire_3790),
        .dout(new_Jinkela_wire_3791)
    );

    or_bb _1550_ (
        .a(_0847_),
        .b(new_Jinkela_wire_4842),
        .c(_0848_)
    );

    or_bb _2264_ (
        .a(new_Jinkela_wire_6375),
        .b(new_Jinkela_wire_6756),
        .c(_0282_)
    );

    bfr new_Jinkela_buffer_2546 (
        .din(new_Jinkela_wire_3805),
        .dout(new_Jinkela_wire_3806)
    );

    and_bi _1551_ (
        .a(_0837_),
        .b(new_Jinkela_wire_6720),
        .c(_0849_)
    );

    or_bb _2265_ (
        .a(new_Jinkela_wire_5439),
        .b(new_Jinkela_wire_7714),
        .c(_0283_)
    );

    bfr new_Jinkela_buffer_2532 (
        .din(new_Jinkela_wire_3791),
        .dout(new_Jinkela_wire_3792)
    );

    and_ii _1552_ (
        .a(_0849_),
        .b(new_Jinkela_wire_7839),
        .c(new_net_11)
    );

    and_ii _2266_ (
        .a(new_Jinkela_wire_7888),
        .b(new_Jinkela_wire_5237),
        .c(_0284_)
    );

    bfr new_Jinkela_buffer_2562 (
        .din(new_Jinkela_wire_3823),
        .dout(new_Jinkela_wire_3824)
    );

    and_bi _1553_ (
        .a(new_Jinkela_wire_304),
        .b(new_Jinkela_wire_6697),
        .c(_0850_)
    );

    and_bi _2267_ (
        .a(_0284_),
        .b(new_Jinkela_wire_5397),
        .c(new_net_2469)
    );

    bfr new_Jinkela_buffer_2533 (
        .din(new_Jinkela_wire_3792),
        .dout(new_Jinkela_wire_3793)
    );

    and_bi _2268_ (
        .a(new_Jinkela_wire_3280),
        .b(new_Jinkela_wire_473),
        .c(_0285_)
    );

    inv _1554_ (
        .din(new_Jinkela_wire_1031),
        .dout(_0851_)
    );

    bfr new_Jinkela_buffer_2547 (
        .din(new_Jinkela_wire_3806),
        .dout(new_Jinkela_wire_3807)
    );

    or_ii _1555_ (
        .a(new_Jinkela_wire_7791),
        .b(new_Jinkela_wire_7691),
        .c(_0852_)
    );

    and_bi _2269_ (
        .a(new_Jinkela_wire_4381),
        .b(new_Jinkela_wire_1645),
        .c(_0286_)
    );

    bfr new_Jinkela_buffer_2534 (
        .din(new_Jinkela_wire_3793),
        .dout(new_Jinkela_wire_3794)
    );

    or_bb _1556_ (
        .a(new_Jinkela_wire_527),
        .b(new_Jinkela_wire_1539),
        .c(_0853_)
    );

    or_bb _2270_ (
        .a(_0286_),
        .b(new_Jinkela_wire_1722),
        .c(_0287_)
    );

    bfr new_Jinkela_buffer_2570 (
        .din(new_Jinkela_wire_3837),
        .dout(new_Jinkela_wire_3838)
    );

    and_bi _1557_ (
        .a(new_Jinkela_wire_528),
        .b(new_Jinkela_wire_1214),
        .c(_0854_)
    );

    or_bb _2271_ (
        .a(new_Jinkela_wire_3579),
        .b(_0285_),
        .c(_0288_)
    );

    bfr new_Jinkela_buffer_2535 (
        .din(new_Jinkela_wire_3794),
        .dout(new_Jinkela_wire_3795)
    );

    and_bi _1558_ (
        .a(_0853_),
        .b(_0854_),
        .c(_0855_)
    );

    and_bi _2272_ (
        .a(new_Jinkela_wire_1017),
        .b(new_Jinkela_wire_7920),
        .c(_0289_)
    );

    bfr new_Jinkela_buffer_2548 (
        .din(new_Jinkela_wire_3807),
        .dout(new_Jinkela_wire_3808)
    );

    and_bi _1559_ (
        .a(new_Jinkela_wire_1040),
        .b(new_Jinkela_wire_2418),
        .c(_0856_)
    );

    and_bi _2273_ (
        .a(new_Jinkela_wire_74),
        .b(new_Jinkela_wire_6130),
        .c(_0290_)
    );

    bfr new_Jinkela_buffer_2536 (
        .din(new_Jinkela_wire_3795),
        .dout(new_Jinkela_wire_3796)
    );

    or_bb _1560_ (
        .a(_0856_),
        .b(new_Jinkela_wire_4824),
        .c(_0857_)
    );

    or_bb _2274_ (
        .a(_0290_),
        .b(_0289_),
        .c(_0291_)
    );

    bfr new_Jinkela_buffer_2563 (
        .din(new_Jinkela_wire_3824),
        .dout(new_Jinkela_wire_3825)
    );

    and_bi _1561_ (
        .a(_0852_),
        .b(new_Jinkela_wire_5420),
        .c(_0858_)
    );

    and_bi _2275_ (
        .a(_0288_),
        .b(new_Jinkela_wire_5613),
        .c(_0292_)
    );

    bfr new_Jinkela_buffer_2537 (
        .din(new_Jinkela_wire_3796),
        .dout(new_Jinkela_wire_3797)
    );

    and_ii _1562_ (
        .a(_0858_),
        .b(new_Jinkela_wire_6434),
        .c(new_net_18)
    );

    and_bi _2276_ (
        .a(new_Jinkela_wire_663),
        .b(_0292_),
        .c(new_net_2427)
    );

    bfr new_Jinkela_buffer_2549 (
        .din(new_Jinkela_wire_3808),
        .dout(new_Jinkela_wire_3809)
    );

    and_bi _2277_ (
        .a(new_Jinkela_wire_3281),
        .b(new_Jinkela_wire_798),
        .c(_0293_)
    );

    and_bi _1563_ (
        .a(new_Jinkela_wire_30),
        .b(new_Jinkela_wire_6695),
        .c(_0859_)
    );

    bfr new_Jinkela_buffer_2538 (
        .din(new_Jinkela_wire_3797),
        .dout(new_Jinkela_wire_3798)
    );

    and_bb _1564_ (
        .a(new_Jinkela_wire_176),
        .b(new_Jinkela_wire_885),
        .c(_0860_)
    );

    and_bi _2278_ (
        .a(new_Jinkela_wire_4380),
        .b(new_Jinkela_wire_6816),
        .c(_0294_)
    );

    bfr new_Jinkela_buffer_2571 (
        .din(new_Jinkela_wire_3838),
        .dout(new_Jinkela_wire_3839)
    );

    and_bi _1565_ (
        .a(new_Jinkela_wire_307),
        .b(new_Jinkela_wire_883),
        .c(_0861_)
    );

    or_bb _2279_ (
        .a(_0294_),
        .b(new_Jinkela_wire_5567),
        .c(_0295_)
    );

    bfr new_Jinkela_buffer_2550 (
        .din(new_Jinkela_wire_3809),
        .dout(new_Jinkela_wire_3810)
    );

    and_ii _1566_ (
        .a(_0861_),
        .b(_0860_),
        .c(_0862_)
    );

    or_bb _2280_ (
        .a(new_Jinkela_wire_4867),
        .b(_0293_),
        .c(_0296_)
    );

    bfr new_Jinkela_buffer_2564 (
        .din(new_Jinkela_wire_3825),
        .dout(new_Jinkela_wire_3826)
    );

    and_bi _1567_ (
        .a(new_Jinkela_wire_763),
        .b(new_Jinkela_wire_6319),
        .c(_0863_)
    );

    and_bi _2281_ (
        .a(new_Jinkela_wire_1018),
        .b(new_Jinkela_wire_3381),
        .c(_0297_)
    );

    bfr new_Jinkela_buffer_2551 (
        .din(new_Jinkela_wire_3810),
        .dout(new_Jinkela_wire_3811)
    );

    and_bi _1568_ (
        .a(new_Jinkela_wire_6322),
        .b(new_Jinkela_wire_764),
        .c(_0864_)
    );

    and_bi _2282_ (
        .a(new_Jinkela_wire_75),
        .b(new_Jinkela_wire_4025),
        .c(_0298_)
    );

    or_bb _2283_ (
        .a(_0298_),
        .b(_0297_),
        .c(_0299_)
    );

    and_bb _1569_ (
        .a(new_Jinkela_wire_832),
        .b(new_Jinkela_wire_869),
        .c(_0865_)
    );

    bfr new_Jinkela_buffer_2552 (
        .din(new_Jinkela_wire_3811),
        .dout(new_Jinkela_wire_3812)
    );

    and_bi _2284_ (
        .a(_0296_),
        .b(new_Jinkela_wire_4813),
        .c(_0300_)
    );

    and_bi _1570_ (
        .a(new_Jinkela_wire_861),
        .b(new_Jinkela_wire_879),
        .c(_0866_)
    );

    spl2 new_Jinkela_splitter_476 (
        .a(new_Jinkela_wire_3826),
        .b(new_Jinkela_wire_3827),
        .c(new_Jinkela_wire_3828)
    );

    bfr new_Jinkela_buffer_2090 (
        .din(new_Jinkela_wire_3204),
        .dout(new_Jinkela_wire_3205)
    );

    bfr new_Jinkela_buffer_2084 (
        .din(new_Jinkela_wire_3198),
        .dout(new_Jinkela_wire_3199)
    );

    bfr new_Jinkela_buffer_2072 (
        .din(new_Jinkela_wire_3183),
        .dout(new_Jinkela_wire_3184)
    );

    bfr new_Jinkela_buffer_2073 (
        .din(new_Jinkela_wire_3184),
        .dout(new_Jinkela_wire_3185)
    );

    spl4L new_Jinkela_splitter_418 (
        .a(_0760_),
        .d(new_Jinkela_wire_3250),
        .e(new_Jinkela_wire_3251),
        .b(new_Jinkela_wire_3252),
        .c(new_Jinkela_wire_3253)
    );

    bfr new_Jinkela_buffer_2085 (
        .din(new_Jinkela_wire_3199),
        .dout(new_Jinkela_wire_3200)
    );

    bfr new_Jinkela_buffer_2074 (
        .din(new_Jinkela_wire_3185),
        .dout(new_Jinkela_wire_3186)
    );

    spl2 new_Jinkela_splitter_417 (
        .a(new_Jinkela_wire_3214),
        .b(new_Jinkela_wire_3215),
        .c(new_Jinkela_wire_3216)
    );

    bfr new_Jinkela_buffer_2075 (
        .din(new_Jinkela_wire_3186),
        .dout(new_Jinkela_wire_3187)
    );

    bfr new_Jinkela_buffer_2091 (
        .din(new_Jinkela_wire_3205),
        .dout(new_Jinkela_wire_3206)
    );

    bfr new_Jinkela_buffer_2086 (
        .din(new_Jinkela_wire_3200),
        .dout(new_Jinkela_wire_3201)
    );

    bfr new_Jinkela_buffer_2076 (
        .din(new_Jinkela_wire_3187),
        .dout(new_Jinkela_wire_3188)
    );

    bfr new_Jinkela_buffer_2077 (
        .din(new_Jinkela_wire_3188),
        .dout(new_Jinkela_wire_3189)
    );

    bfr new_Jinkela_buffer_2087 (
        .din(new_Jinkela_wire_3201),
        .dout(new_Jinkela_wire_3202)
    );

    bfr new_Jinkela_buffer_2078 (
        .din(new_Jinkela_wire_3189),
        .dout(new_Jinkela_wire_3190)
    );

    bfr new_Jinkela_buffer_2079 (
        .din(new_Jinkela_wire_3190),
        .dout(new_Jinkela_wire_3191)
    );

    bfr new_Jinkela_buffer_2092 (
        .din(new_Jinkela_wire_3206),
        .dout(new_Jinkela_wire_3207)
    );

    bfr new_Jinkela_buffer_2080 (
        .din(new_Jinkela_wire_3191),
        .dout(new_Jinkela_wire_3192)
    );

    bfr new_Jinkela_buffer_2133 (
        .din(new_Jinkela_wire_3253),
        .dout(new_Jinkela_wire_3254)
    );

    bfr new_Jinkela_buffer_2141 (
        .din(new_net_2353),
        .dout(new_Jinkela_wire_3264)
    );

    bfr new_Jinkela_buffer_2093 (
        .din(new_Jinkela_wire_3207),
        .dout(new_Jinkela_wire_3208)
    );

    bfr new_Jinkela_buffer_2101 (
        .din(new_Jinkela_wire_3217),
        .dout(new_Jinkela_wire_3218)
    );

    bfr new_Jinkela_buffer_2094 (
        .din(new_Jinkela_wire_3208),
        .dout(new_Jinkela_wire_3209)
    );

    bfr new_Jinkela_buffer_2102 (
        .din(new_Jinkela_wire_3218),
        .dout(new_Jinkela_wire_3219)
    );

    bfr new_Jinkela_buffer_2095 (
        .din(new_Jinkela_wire_3209),
        .dout(new_Jinkela_wire_3210)
    );

    bfr new_Jinkela_buffer_2096 (
        .din(new_Jinkela_wire_3210),
        .dout(new_Jinkela_wire_3211)
    );

    bfr new_Jinkela_buffer_2103 (
        .din(new_Jinkela_wire_3219),
        .dout(new_Jinkela_wire_3220)
    );

    bfr new_Jinkela_buffer_2097 (
        .din(new_Jinkela_wire_3211),
        .dout(new_Jinkela_wire_3212)
    );

    spl2 new_Jinkela_splitter_420 (
        .a(_1200_),
        .b(new_Jinkela_wire_3274),
        .c(new_Jinkela_wire_3275)
    );

    bfr new_Jinkela_buffer_2098 (
        .din(new_Jinkela_wire_3212),
        .dout(new_Jinkela_wire_3213)
    );

    bfr new_Jinkela_buffer_2104 (
        .din(new_Jinkela_wire_3220),
        .dout(new_Jinkela_wire_3221)
    );

    spl2 new_Jinkela_splitter_421 (
        .a(new_net_3),
        .b(new_Jinkela_wire_3276),
        .c(new_Jinkela_wire_3278)
    );

    bfr new_Jinkela_buffer_2105 (
        .din(new_Jinkela_wire_3221),
        .dout(new_Jinkela_wire_3222)
    );

    bfr new_Jinkela_buffer_2134 (
        .din(new_Jinkela_wire_3254),
        .dout(new_Jinkela_wire_3255)
    );

    bfr new_Jinkela_buffer_2106 (
        .din(new_Jinkela_wire_3222),
        .dout(new_Jinkela_wire_3223)
    );

    bfr new_Jinkela_buffer_2107 (
        .din(new_Jinkela_wire_3223),
        .dout(new_Jinkela_wire_3224)
    );

    bfr new_Jinkela_buffer_2135 (
        .din(new_Jinkela_wire_3255),
        .dout(new_Jinkela_wire_3256)
    );

    bfr new_Jinkela_buffer_2143 (
        .din(new_Jinkela_wire_3265),
        .dout(new_Jinkela_wire_3266)
    );

    bfr new_Jinkela_buffer_2108 (
        .din(new_Jinkela_wire_3224),
        .dout(new_Jinkela_wire_3225)
    );

    bfr new_Jinkela_buffer_2142 (
        .din(new_Jinkela_wire_3264),
        .dout(new_Jinkela_wire_3265)
    );

    bfr new_Jinkela_buffer_2109 (
        .din(new_Jinkela_wire_3225),
        .dout(new_Jinkela_wire_3226)
    );

    bfr new_Jinkela_buffer_2136 (
        .din(new_Jinkela_wire_3256),
        .dout(new_Jinkela_wire_3257)
    );

    bfr new_Jinkela_buffer_3568 (
        .din(new_Jinkela_wire_5018),
        .dout(new_Jinkela_wire_5019)
    );

    bfr new_Jinkela_buffer_3588 (
        .din(new_Jinkela_wire_5038),
        .dout(new_Jinkela_wire_5039)
    );

    bfr new_Jinkela_buffer_3569 (
        .din(new_Jinkela_wire_5019),
        .dout(new_Jinkela_wire_5020)
    );

    bfr new_Jinkela_buffer_3623 (
        .din(new_Jinkela_wire_5081),
        .dout(new_Jinkela_wire_5082)
    );

    bfr new_Jinkela_buffer_3570 (
        .din(new_Jinkela_wire_5020),
        .dout(new_Jinkela_wire_5021)
    );

    bfr new_Jinkela_buffer_3589 (
        .din(new_Jinkela_wire_5039),
        .dout(new_Jinkela_wire_5040)
    );

    bfr new_Jinkela_buffer_3571 (
        .din(new_Jinkela_wire_5021),
        .dout(new_Jinkela_wire_5022)
    );

    bfr new_Jinkela_buffer_3600 (
        .din(new_Jinkela_wire_5058),
        .dout(new_Jinkela_wire_5059)
    );

    bfr new_Jinkela_buffer_3572 (
        .din(new_Jinkela_wire_5022),
        .dout(new_Jinkela_wire_5023)
    );

    bfr new_Jinkela_buffer_3590 (
        .din(new_Jinkela_wire_5040),
        .dout(new_Jinkela_wire_5041)
    );

    bfr new_Jinkela_buffer_3573 (
        .din(new_Jinkela_wire_5023),
        .dout(new_Jinkela_wire_5024)
    );

    bfr new_Jinkela_buffer_3574 (
        .din(new_Jinkela_wire_5024),
        .dout(new_Jinkela_wire_5025)
    );

    bfr new_Jinkela_buffer_3591 (
        .din(new_Jinkela_wire_5041),
        .dout(new_Jinkela_wire_5042)
    );

    bfr new_Jinkela_buffer_3575 (
        .din(new_Jinkela_wire_5025),
        .dout(new_Jinkela_wire_5026)
    );

    bfr new_Jinkela_buffer_3601 (
        .din(new_Jinkela_wire_5059),
        .dout(new_Jinkela_wire_5060)
    );

    bfr new_Jinkela_buffer_3576 (
        .din(new_Jinkela_wire_5026),
        .dout(new_Jinkela_wire_5027)
    );

    bfr new_Jinkela_buffer_3592 (
        .din(new_Jinkela_wire_5042),
        .dout(new_Jinkela_wire_5043)
    );

    bfr new_Jinkela_buffer_3577 (
        .din(new_Jinkela_wire_5027),
        .dout(new_Jinkela_wire_5028)
    );

    bfr new_Jinkela_buffer_3624 (
        .din(new_Jinkela_wire_5082),
        .dout(new_Jinkela_wire_5083)
    );

    bfr new_Jinkela_buffer_3578 (
        .din(new_Jinkela_wire_5028),
        .dout(new_Jinkela_wire_5029)
    );

    bfr new_Jinkela_buffer_3593 (
        .din(new_Jinkela_wire_5043),
        .dout(new_Jinkela_wire_5044)
    );

    bfr new_Jinkela_buffer_3579 (
        .din(new_Jinkela_wire_5029),
        .dout(new_Jinkela_wire_5030)
    );

    bfr new_Jinkela_buffer_3602 (
        .din(new_Jinkela_wire_5060),
        .dout(new_Jinkela_wire_5061)
    );

    bfr new_Jinkela_buffer_3594 (
        .din(new_Jinkela_wire_5044),
        .dout(new_Jinkela_wire_5045)
    );

    bfr new_Jinkela_buffer_3656 (
        .din(new_Jinkela_wire_5116),
        .dout(new_Jinkela_wire_5117)
    );

    bfr new_Jinkela_buffer_3595 (
        .din(new_Jinkela_wire_5045),
        .dout(new_Jinkela_wire_5046)
    );

    bfr new_Jinkela_buffer_3603 (
        .din(new_Jinkela_wire_5061),
        .dout(new_Jinkela_wire_5062)
    );

    bfr new_Jinkela_buffer_3596 (
        .din(new_Jinkela_wire_5046),
        .dout(new_Jinkela_wire_5047)
    );

    bfr new_Jinkela_buffer_3625 (
        .din(new_Jinkela_wire_5083),
        .dout(new_Jinkela_wire_5084)
    );

    bfr new_Jinkela_buffer_3604 (
        .din(new_Jinkela_wire_5062),
        .dout(new_Jinkela_wire_5063)
    );

    bfr new_Jinkela_buffer_3658 (
        .din(_0275_),
        .dout(new_Jinkela_wire_5119)
    );

    bfr new_Jinkela_buffer_3605 (
        .din(new_Jinkela_wire_5063),
        .dout(new_Jinkela_wire_5064)
    );

    bfr new_Jinkela_buffer_3626 (
        .din(new_Jinkela_wire_5084),
        .dout(new_Jinkela_wire_5085)
    );

    bfr new_Jinkela_buffer_3606 (
        .din(new_Jinkela_wire_5064),
        .dout(new_Jinkela_wire_5065)
    );

    spl2 new_Jinkela_splitter_554 (
        .a(_1121_),
        .b(new_Jinkela_wire_5121),
        .c(new_Jinkela_wire_5122)
    );

    spl2 new_Jinkela_splitter_555 (
        .a(_0210_),
        .b(new_Jinkela_wire_5123),
        .c(new_Jinkela_wire_5124)
    );

    bfr new_Jinkela_buffer_3607 (
        .din(new_Jinkela_wire_5065),
        .dout(new_Jinkela_wire_5066)
    );

    bfr new_Jinkela_buffer_3627 (
        .din(new_Jinkela_wire_5085),
        .dout(new_Jinkela_wire_5086)
    );

    bfr new_Jinkela_buffer_3608 (
        .din(new_Jinkela_wire_5066),
        .dout(new_Jinkela_wire_5067)
    );

    bfr new_Jinkela_buffer_3657 (
        .din(new_Jinkela_wire_5117),
        .dout(new_Jinkela_wire_5118)
    );

    bfr new_Jinkela_buffer_3609 (
        .din(new_Jinkela_wire_5067),
        .dout(new_Jinkela_wire_5068)
    );

    bfr new_Jinkela_buffer_3628 (
        .din(new_Jinkela_wire_5086),
        .dout(new_Jinkela_wire_5087)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_2508),
        .dout(new_Jinkela_wire_2509)
    );

    bfr new_Jinkela_buffer_2461 (
        .din(new_Jinkela_wire_3706),
        .dout(new_Jinkela_wire_3707)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_2477),
        .dout(new_Jinkela_wire_2478)
    );

    bfr new_Jinkela_buffer_2481 (
        .din(new_Jinkela_wire_3728),
        .dout(new_Jinkela_wire_3729)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_2540),
        .dout(new_Jinkela_wire_2541)
    );

    bfr new_Jinkela_buffer_2462 (
        .din(new_Jinkela_wire_3707),
        .dout(new_Jinkela_wire_3708)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_2478),
        .dout(new_Jinkela_wire_2479)
    );

    bfr new_Jinkela_buffer_2505 (
        .din(new_Jinkela_wire_3758),
        .dout(new_Jinkela_wire_3759)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_2509),
        .dout(new_Jinkela_wire_2510)
    );

    bfr new_Jinkela_buffer_2463 (
        .din(new_Jinkela_wire_3708),
        .dout(new_Jinkela_wire_3709)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(new_Jinkela_wire_2479),
        .dout(new_Jinkela_wire_2480)
    );

    bfr new_Jinkela_buffer_2482 (
        .din(new_Jinkela_wire_3729),
        .dout(new_Jinkela_wire_3730)
    );

    bfr new_Jinkela_buffer_2464 (
        .din(new_Jinkela_wire_3709),
        .dout(new_Jinkela_wire_3710)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(new_Jinkela_wire_2480),
        .dout(new_Jinkela_wire_2481)
    );

    spl4L new_Jinkela_splitter_474 (
        .a(new_Jinkela_wire_3770),
        .d(new_Jinkela_wire_3771),
        .e(new_Jinkela_wire_3772),
        .b(new_Jinkela_wire_3773),
        .c(new_Jinkela_wire_3774)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_2510),
        .dout(new_Jinkela_wire_2511)
    );

    bfr new_Jinkela_buffer_2465 (
        .din(new_Jinkela_wire_3710),
        .dout(new_Jinkela_wire_3711)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_2481),
        .dout(new_Jinkela_wire_2482)
    );

    bfr new_Jinkela_buffer_2483 (
        .din(new_Jinkela_wire_3730),
        .dout(new_Jinkela_wire_3731)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_2541),
        .dout(new_Jinkela_wire_2542)
    );

    bfr new_Jinkela_buffer_2466 (
        .din(new_Jinkela_wire_3711),
        .dout(new_Jinkela_wire_3712)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(new_Jinkela_wire_2482),
        .dout(new_Jinkela_wire_2483)
    );

    bfr new_Jinkela_buffer_2506 (
        .din(new_Jinkela_wire_3759),
        .dout(new_Jinkela_wire_3760)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_2511),
        .dout(new_Jinkela_wire_2512)
    );

    bfr new_Jinkela_buffer_2467 (
        .din(new_Jinkela_wire_3712),
        .dout(new_Jinkela_wire_3713)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(new_Jinkela_wire_2483),
        .dout(new_Jinkela_wire_2484)
    );

    bfr new_Jinkela_buffer_2484 (
        .din(new_Jinkela_wire_3731),
        .dout(new_Jinkela_wire_3732)
    );

    spl2 new_Jinkela_splitter_378 (
        .a(_0972_),
        .b(new_Jinkela_wire_2622),
        .c(new_Jinkela_wire_2623)
    );

    bfr new_Jinkela_buffer_2515 (
        .din(new_Jinkela_wire_3774),
        .dout(new_Jinkela_wire_3775)
    );

    bfr new_Jinkela_buffer_1612 (
        .din(new_net_2407),
        .dout(new_Jinkela_wire_2624)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(new_Jinkela_wire_2484),
        .dout(new_Jinkela_wire_2485)
    );

    bfr new_Jinkela_buffer_2485 (
        .din(new_Jinkela_wire_3732),
        .dout(new_Jinkela_wire_3733)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_2512),
        .dout(new_Jinkela_wire_2513)
    );

    bfr new_Jinkela_buffer_2507 (
        .din(new_Jinkela_wire_3760),
        .dout(new_Jinkela_wire_3761)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_2485),
        .dout(new_Jinkela_wire_2486)
    );

    bfr new_Jinkela_buffer_2486 (
        .din(new_Jinkela_wire_3733),
        .dout(new_Jinkela_wire_3734)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_2542),
        .dout(new_Jinkela_wire_2543)
    );

    bfr new_Jinkela_buffer_2518 (
        .din(new_Jinkela_wire_3777),
        .dout(new_Jinkela_wire_3778)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(new_Jinkela_wire_2486),
        .dout(new_Jinkela_wire_2487)
    );

    bfr new_Jinkela_buffer_2487 (
        .din(new_Jinkela_wire_3734),
        .dout(new_Jinkela_wire_3735)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_2513),
        .dout(new_Jinkela_wire_2514)
    );

    bfr new_Jinkela_buffer_2508 (
        .din(new_Jinkela_wire_3761),
        .dout(new_Jinkela_wire_3762)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(new_Jinkela_wire_2487),
        .dout(new_Jinkela_wire_2488)
    );

    bfr new_Jinkela_buffer_2488 (
        .din(new_Jinkela_wire_3735),
        .dout(new_Jinkela_wire_3736)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(new_Jinkela_wire_2582),
        .dout(new_Jinkela_wire_2583)
    );

    spl2 new_Jinkela_splitter_475 (
        .a(_0661_),
        .b(new_Jinkela_wire_3820),
        .c(new_Jinkela_wire_3821)
    );

    bfr new_Jinkela_buffer_2516 (
        .din(new_Jinkela_wire_3775),
        .dout(new_Jinkela_wire_3776)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_2572),
        .dout(new_Jinkela_wire_2573)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(new_Jinkela_wire_2488),
        .dout(new_Jinkela_wire_2489)
    );

    bfr new_Jinkela_buffer_2489 (
        .din(new_Jinkela_wire_3736),
        .dout(new_Jinkela_wire_3737)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_2514),
        .dout(new_Jinkela_wire_2515)
    );

    bfr new_Jinkela_buffer_2509 (
        .din(new_Jinkela_wire_3762),
        .dout(new_Jinkela_wire_3763)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(new_Jinkela_wire_2489),
        .dout(new_Jinkela_wire_2490)
    );

    bfr new_Jinkela_buffer_2490 (
        .din(new_Jinkela_wire_3737),
        .dout(new_Jinkela_wire_3738)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(new_Jinkela_wire_2543),
        .dout(new_Jinkela_wire_2544)
    );

    spl4L new_Jinkela_splitter_477 (
        .a(_0985_),
        .d(new_Jinkela_wire_3833),
        .e(new_Jinkela_wire_3834),
        .b(new_Jinkela_wire_3835),
        .c(new_Jinkela_wire_3836)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_2490),
        .dout(new_Jinkela_wire_2491)
    );

    bfr new_Jinkela_buffer_2491 (
        .din(new_Jinkela_wire_3738),
        .dout(new_Jinkela_wire_3739)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_2515),
        .dout(new_Jinkela_wire_2516)
    );

    bfr new_Jinkela_buffer_2510 (
        .din(new_Jinkela_wire_3763),
        .dout(new_Jinkela_wire_3764)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(new_Jinkela_wire_2491),
        .dout(new_Jinkela_wire_2492)
    );

    bfr new_Jinkela_buffer_2492 (
        .din(new_Jinkela_wire_3739),
        .dout(new_Jinkela_wire_3740)
    );

    bfr new_Jinkela_buffer_2519 (
        .din(new_Jinkela_wire_3778),
        .dout(new_Jinkela_wire_3779)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_2492),
        .dout(new_Jinkela_wire_2493)
    );

    bfr new_Jinkela_buffer_2493 (
        .din(new_Jinkela_wire_3740),
        .dout(new_Jinkela_wire_3741)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_2516),
        .dout(new_Jinkela_wire_2517)
    );

    bfr new_Jinkela_buffer_2511 (
        .din(new_Jinkela_wire_3764),
        .dout(new_Jinkela_wire_3765)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_2493),
        .dout(new_Jinkela_wire_2494)
    );

    bfr new_Jinkela_buffer_2494 (
        .din(new_Jinkela_wire_3741),
        .dout(new_Jinkela_wire_3742)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_2544),
        .dout(new_Jinkela_wire_2545)
    );

    bfr new_Jinkela_buffer_2540 (
        .din(new_Jinkela_wire_3799),
        .dout(new_Jinkela_wire_3800)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(new_Jinkela_wire_2494),
        .dout(new_Jinkela_wire_2495)
    );

    bfr new_Jinkela_buffer_2495 (
        .din(new_Jinkela_wire_3742),
        .dout(new_Jinkela_wire_3743)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_2517),
        .dout(new_Jinkela_wire_2518)
    );

    bfr new_Jinkela_buffer_2512 (
        .din(new_Jinkela_wire_3765),
        .dout(new_Jinkela_wire_3766)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(new_Jinkela_wire_2495),
        .dout(new_Jinkela_wire_2496)
    );

    bfr new_Jinkela_buffer_2496 (
        .din(new_Jinkela_wire_3743),
        .dout(new_Jinkela_wire_3744)
    );

    bfr new_Jinkela_buffer_2520 (
        .din(new_Jinkela_wire_3779),
        .dout(new_Jinkela_wire_3780)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_2573),
        .dout(new_Jinkela_wire_2574)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(new_Jinkela_wire_2496),
        .dout(new_Jinkela_wire_2497)
    );

    bfr new_Jinkela_buffer_2497 (
        .din(new_Jinkela_wire_3744),
        .dout(new_Jinkela_wire_3745)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_2518),
        .dout(new_Jinkela_wire_2519)
    );

    bfr new_Jinkela_buffer_2569 (
        .din(new_net_2403),
        .dout(new_Jinkela_wire_3837)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_2497),
        .dout(new_Jinkela_wire_2498)
    );

    bfr new_Jinkela_buffer_2498 (
        .din(new_Jinkela_wire_3745),
        .dout(new_Jinkela_wire_3746)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1664),
        .dout(new_Jinkela_wire_1665)
    );

    bfr new_Jinkela_buffer_3610 (
        .din(new_Jinkela_wire_5068),
        .dout(new_Jinkela_wire_5069)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1696),
        .dout(new_Jinkela_wire_1697)
    );

    bfr new_Jinkela_buffer_3659 (
        .din(new_Jinkela_wire_5119),
        .dout(new_Jinkela_wire_5120)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_1665),
        .dout(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_3611 (
        .din(new_Jinkela_wire_5069),
        .dout(new_Jinkela_wire_5070)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1788),
        .dout(new_Jinkela_wire_1789)
    );

    bfr new_Jinkela_buffer_3629 (
        .din(new_Jinkela_wire_5087),
        .dout(new_Jinkela_wire_5088)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1713),
        .dout(new_Jinkela_wire_1714)
    );

    spl2 new_Jinkela_splitter_307 (
        .a(new_Jinkela_wire_1666),
        .b(new_Jinkela_wire_1667),
        .c(new_Jinkela_wire_1668)
    );

    bfr new_Jinkela_buffer_3612 (
        .din(new_Jinkela_wire_5070),
        .dout(new_Jinkela_wire_5071)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1668),
        .dout(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_3685 (
        .din(new_net_2497),
        .dout(new_Jinkela_wire_5158)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1697),
        .dout(new_Jinkela_wire_1698)
    );

    bfr new_Jinkela_buffer_3613 (
        .din(new_Jinkela_wire_5071),
        .dout(new_Jinkela_wire_5072)
    );

    bfr new_Jinkela_buffer_3630 (
        .din(new_Jinkela_wire_5088),
        .dout(new_Jinkela_wire_5089)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_3614 (
        .din(new_Jinkela_wire_5072),
        .dout(new_Jinkela_wire_5073)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_1698),
        .dout(new_Jinkela_wire_1699)
    );

    spl4L new_Jinkela_splitter_556 (
        .a(_0946_),
        .d(new_Jinkela_wire_5125),
        .e(new_Jinkela_wire_5126),
        .b(new_Jinkela_wire_5127),
        .c(new_Jinkela_wire_5128)
    );

    spl2 new_Jinkela_splitter_308 (
        .a(new_Jinkela_wire_1670),
        .b(new_Jinkela_wire_1671),
        .c(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_3615 (
        .din(new_Jinkela_wire_5073),
        .dout(new_Jinkela_wire_5074)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1672),
        .dout(new_Jinkela_wire_1673)
    );

    bfr new_Jinkela_buffer_3631 (
        .din(new_Jinkela_wire_5089),
        .dout(new_Jinkela_wire_5090)
    );

    bfr new_Jinkela_buffer_3616 (
        .din(new_Jinkela_wire_5074),
        .dout(new_Jinkela_wire_5075)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1758),
        .dout(new_Jinkela_wire_1759)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1699),
        .dout(new_Jinkela_wire_1700)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1673),
        .dout(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_3617 (
        .din(new_Jinkela_wire_5075),
        .dout(new_Jinkela_wire_5076)
    );

    spl2 new_Jinkela_splitter_323 (
        .a(_0710_),
        .b(new_Jinkela_wire_1851),
        .c(new_Jinkela_wire_1852)
    );

    bfr new_Jinkela_buffer_3632 (
        .din(new_Jinkela_wire_5090),
        .dout(new_Jinkela_wire_5091)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1712),
        .dout(new_Jinkela_wire_1713)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_1674),
        .dout(new_Jinkela_wire_1675)
    );

    bfr new_Jinkela_buffer_3618 (
        .din(new_Jinkela_wire_5076),
        .dout(new_Jinkela_wire_5077)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_1700),
        .dout(new_Jinkela_wire_1701)
    );

    spl2 new_Jinkela_splitter_557 (
        .a(_0159_),
        .b(new_Jinkela_wire_5129),
        .c(new_Jinkela_wire_5130)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1714),
        .dout(new_Jinkela_wire_1715)
    );

    bfr new_Jinkela_buffer_3619 (
        .din(new_Jinkela_wire_5077),
        .dout(new_Jinkela_wire_5078)
    );

    spl2 new_Jinkela_splitter_322 (
        .a(_0679_),
        .b(new_Jinkela_wire_1849),
        .c(new_Jinkela_wire_1850)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_1701),
        .dout(new_Jinkela_wire_1702)
    );

    bfr new_Jinkela_buffer_3633 (
        .din(new_Jinkela_wire_5091),
        .dout(new_Jinkela_wire_5092)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1715),
        .dout(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_3620 (
        .din(new_Jinkela_wire_5078),
        .dout(new_Jinkela_wire_5079)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1702),
        .dout(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_3660 (
        .din(_0889_),
        .dout(new_Jinkela_wire_5131)
    );

    bfr new_Jinkela_buffer_3661 (
        .din(new_Jinkela_wire_5131),
        .dout(new_Jinkela_wire_5132)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1759),
        .dout(new_Jinkela_wire_1760)
    );

    bfr new_Jinkela_buffer_3621 (
        .din(new_Jinkela_wire_5079),
        .dout(new_Jinkela_wire_5080)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1703),
        .dout(new_Jinkela_wire_1704)
    );

    bfr new_Jinkela_buffer_3634 (
        .din(new_Jinkela_wire_5092),
        .dout(new_Jinkela_wire_5093)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    spl2 new_Jinkela_splitter_558 (
        .a(_0991_),
        .b(new_Jinkela_wire_5156),
        .c(new_Jinkela_wire_5157)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1704),
        .dout(new_Jinkela_wire_1705)
    );

    bfr new_Jinkela_buffer_3635 (
        .din(new_Jinkela_wire_5093),
        .dout(new_Jinkela_wire_5094)
    );

    bfr new_Jinkela_buffer_3686 (
        .din(new_Jinkela_wire_5158),
        .dout(new_Jinkela_wire_5159)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1705),
        .dout(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_3636 (
        .din(new_Jinkela_wire_5094),
        .dout(new_Jinkela_wire_5095)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_1760),
        .dout(new_Jinkela_wire_1761)
    );

    bfr new_Jinkela_buffer_3662 (
        .din(new_Jinkela_wire_5132),
        .dout(new_Jinkela_wire_5133)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1717),
        .dout(new_Jinkela_wire_1718)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1706),
        .dout(new_Jinkela_wire_1707)
    );

    bfr new_Jinkela_buffer_3637 (
        .din(new_Jinkela_wire_5095),
        .dout(new_Jinkela_wire_5096)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1707),
        .dout(new_Jinkela_wire_1708)
    );

    bfr new_Jinkela_buffer_3638 (
        .din(new_Jinkela_wire_5096),
        .dout(new_Jinkela_wire_5097)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1716),
        .dout(new_Jinkela_wire_1717)
    );

    bfr new_Jinkela_buffer_3663 (
        .din(new_Jinkela_wire_5133),
        .dout(new_Jinkela_wire_5134)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1718),
        .dout(new_Jinkela_wire_1719)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_1761),
        .dout(new_Jinkela_wire_1762)
    );

    bfr new_Jinkela_buffer_3639 (
        .din(new_Jinkela_wire_5097),
        .dout(new_Jinkela_wire_5098)
    );

    bfr new_Jinkela_buffer_3719 (
        .din(_1075_),
        .dout(new_Jinkela_wire_5192)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1789),
        .dout(new_Jinkela_wire_1790)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1719),
        .dout(new_Jinkela_wire_1720)
    );

    bfr new_Jinkela_buffer_3640 (
        .din(new_Jinkela_wire_5098),
        .dout(new_Jinkela_wire_5099)
    );

    bfr new_Jinkela_buffer_3664 (
        .din(new_Jinkela_wire_5134),
        .dout(new_Jinkela_wire_5135)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1790),
        .dout(new_Jinkela_wire_1791)
    );

    bfr new_Jinkela_buffer_3641 (
        .din(new_Jinkela_wire_5099),
        .dout(new_Jinkela_wire_5100)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1720),
        .dout(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_3720 (
        .din(_0024_),
        .dout(new_Jinkela_wire_5193)
    );

    bfr new_Jinkela_buffer_3723 (
        .din(_0254_),
        .dout(new_Jinkela_wire_5198)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1762),
        .dout(new_Jinkela_wire_1763)
    );

    bfr new_Jinkela_buffer_3642 (
        .din(new_Jinkela_wire_5100),
        .dout(new_Jinkela_wire_5101)
    );

    spl2 new_Jinkela_splitter_312 (
        .a(new_Jinkela_wire_1721),
        .b(new_Jinkela_wire_1722),
        .c(new_Jinkela_wire_1723)
    );

    bfr new_Jinkela_buffer_3665 (
        .din(new_Jinkela_wire_5135),
        .dout(new_Jinkela_wire_5136)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1723),
        .dout(new_Jinkela_wire_1724)
    );

    bfr new_Jinkela_buffer_3643 (
        .din(new_Jinkela_wire_5101),
        .dout(new_Jinkela_wire_5102)
    );

    spl3L new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_437),
        .d(new_Jinkela_wire_438),
        .b(new_Jinkela_wire_442),
        .c(new_Jinkela_wire_447)
    );

    bfr new_Jinkela_buffer_2110 (
        .din(new_Jinkela_wire_3226),
        .dout(new_Jinkela_wire_3227)
    );

    bfr new_Jinkela_buffer_3226 (
        .din(new_Jinkela_wire_4607),
        .dout(new_Jinkela_wire_4608)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_3191 (
        .din(new_Jinkela_wire_4552),
        .dout(new_Jinkela_wire_4553)
    );

    bfr new_Jinkela_buffer_2175 (
        .din(new_net_2489),
        .dout(new_Jinkela_wire_3306)
    );

    bfr new_Jinkela_buffer_2111 (
        .din(new_Jinkela_wire_3227),
        .dout(new_Jinkela_wire_3228)
    );

    spl4L new_Jinkela_splitter_91 (
        .a(new_Jinkela_wire_431),
        .d(new_Jinkela_wire_432),
        .e(new_Jinkela_wire_433),
        .b(new_Jinkela_wire_434),
        .c(new_Jinkela_wire_435)
    );

    spl3L new_Jinkela_splitter_520 (
        .a(new_Jinkela_wire_4571),
        .d(new_Jinkela_wire_4572),
        .b(new_Jinkela_wire_4573),
        .c(new_Jinkela_wire_4574)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_350),
        .dout(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_2137 (
        .din(new_Jinkela_wire_3257),
        .dout(new_Jinkela_wire_3258)
    );

    bfr new_Jinkela_buffer_3192 (
        .din(new_Jinkela_wire_4553),
        .dout(new_Jinkela_wire_4554)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_2112 (
        .din(new_Jinkela_wire_3228),
        .dout(new_Jinkela_wire_3229)
    );

    bfr new_Jinkela_buffer_3206 (
        .din(new_Jinkela_wire_4579),
        .dout(new_Jinkela_wire_4580)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_2144 (
        .din(new_Jinkela_wire_3266),
        .dout(new_Jinkela_wire_3267)
    );

    bfr new_Jinkela_buffer_3193 (
        .din(new_Jinkela_wire_4554),
        .dout(new_Jinkela_wire_4555)
    );

    bfr new_Jinkela_buffer_2113 (
        .din(new_Jinkela_wire_3229),
        .dout(new_Jinkela_wire_3230)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_2138 (
        .din(new_Jinkela_wire_3258),
        .dout(new_Jinkela_wire_3259)
    );

    bfr new_Jinkela_buffer_3194 (
        .din(new_Jinkela_wire_4555),
        .dout(new_Jinkela_wire_4556)
    );

    bfr new_Jinkela_buffer_2114 (
        .din(new_Jinkela_wire_3230),
        .dout(new_Jinkela_wire_3231)
    );

    bfr new_Jinkela_buffer_3225 (
        .din(_0756_),
        .dout(new_Jinkela_wire_4605)
    );

    spl3L new_Jinkela_splitter_526 (
        .a(_0748_),
        .d(new_Jinkela_wire_4612),
        .b(new_Jinkela_wire_4613),
        .c(new_Jinkela_wire_4614)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    bfr new_Jinkela_buffer_2152 (
        .din(new_Jinkela_wire_3282),
        .dout(new_Jinkela_wire_3283)
    );

    bfr new_Jinkela_buffer_3195 (
        .din(new_Jinkela_wire_4556),
        .dout(new_Jinkela_wire_4557)
    );

    spl3L new_Jinkela_splitter_93 (
        .a(new_Jinkela_wire_438),
        .d(new_Jinkela_wire_439),
        .b(new_Jinkela_wire_440),
        .c(new_Jinkela_wire_441)
    );

    bfr new_Jinkela_buffer_2115 (
        .din(new_Jinkela_wire_3231),
        .dout(new_Jinkela_wire_3232)
    );

    bfr new_Jinkela_buffer_3207 (
        .din(new_Jinkela_wire_4580),
        .dout(new_Jinkela_wire_4581)
    );

    bfr new_Jinkela_buffer_201 (
        .din(G68),
        .dout(new_Jinkela_wire_516)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_354),
        .dout(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_2139 (
        .din(new_Jinkela_wire_3259),
        .dout(new_Jinkela_wire_3260)
    );

    bfr new_Jinkela_buffer_3196 (
        .din(new_Jinkela_wire_4557),
        .dout(new_Jinkela_wire_4558)
    );

    bfr new_Jinkela_buffer_2116 (
        .din(new_Jinkela_wire_3232),
        .dout(new_Jinkela_wire_3233)
    );

    spl2 new_Jinkela_splitter_525 (
        .a(_0643_),
        .b(new_Jinkela_wire_4606),
        .c(new_Jinkela_wire_4607)
    );

    spl4L new_Jinkela_splitter_95 (
        .a(new_Jinkela_wire_447),
        .d(new_Jinkela_wire_448),
        .e(new_Jinkela_wire_449),
        .b(new_Jinkela_wire_450),
        .c(new_Jinkela_wire_451)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_2145 (
        .din(new_Jinkela_wire_3267),
        .dout(new_Jinkela_wire_3268)
    );

    bfr new_Jinkela_buffer_3197 (
        .din(new_Jinkela_wire_4558),
        .dout(new_Jinkela_wire_4559)
    );

    bfr new_Jinkela_buffer_2117 (
        .din(new_Jinkela_wire_3233),
        .dout(new_Jinkela_wire_3234)
    );

    bfr new_Jinkela_buffer_3208 (
        .din(new_Jinkela_wire_4581),
        .dout(new_Jinkela_wire_4582)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_2140 (
        .din(new_Jinkela_wire_3260),
        .dout(new_Jinkela_wire_3261)
    );

    bfr new_Jinkela_buffer_3198 (
        .din(new_Jinkela_wire_4559),
        .dout(new_Jinkela_wire_4560)
    );

    spl4L new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_442),
        .d(new_Jinkela_wire_443),
        .e(new_Jinkela_wire_444),
        .b(new_Jinkela_wire_445),
        .c(new_Jinkela_wire_446)
    );

    bfr new_Jinkela_buffer_2118 (
        .din(new_Jinkela_wire_3234),
        .dout(new_Jinkela_wire_3235)
    );

    bfr new_Jinkela_buffer_3230 (
        .din(new_net_26),
        .dout(new_Jinkela_wire_4615)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(new_Jinkela_wire_357),
        .b(new_Jinkela_wire_358),
        .c(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_3199 (
        .din(new_Jinkela_wire_4560),
        .dout(new_Jinkela_wire_4561)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_359),
        .dout(new_Jinkela_wire_360)
    );

    bfr new_Jinkela_buffer_2119 (
        .din(new_Jinkela_wire_3235),
        .dout(new_Jinkela_wire_3236)
    );

    bfr new_Jinkela_buffer_3209 (
        .din(new_Jinkela_wire_4582),
        .dout(new_Jinkela_wire_4583)
    );

    spl2 new_Jinkela_splitter_419 (
        .a(new_Jinkela_wire_3261),
        .b(new_Jinkela_wire_3262),
        .c(new_Jinkela_wire_3263)
    );

    bfr new_Jinkela_buffer_3200 (
        .din(new_Jinkela_wire_4561),
        .dout(new_Jinkela_wire_4562)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_503),
        .dout(new_Jinkela_wire_504)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(G138),
        .b(new_Jinkela_wire_508),
        .c(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_2120 (
        .din(new_Jinkela_wire_3236),
        .dout(new_Jinkela_wire_3237)
    );

    bfr new_Jinkela_buffer_3269 (
        .din(new_net_2461),
        .dout(new_Jinkela_wire_4656)
    );

    spl2 new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_360),
        .b(new_Jinkela_wire_361),
        .c(new_Jinkela_wire_362)
    );

    spl4L new_Jinkela_splitter_422 (
        .a(new_Jinkela_wire_3278),
        .d(new_Jinkela_wire_3279),
        .e(new_Jinkela_wire_3280),
        .b(new_Jinkela_wire_3281),
        .c(new_Jinkela_wire_3282)
    );

    bfr new_Jinkela_buffer_3201 (
        .din(new_Jinkela_wire_4562),
        .dout(new_Jinkela_wire_4563)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    bfr new_Jinkela_buffer_2121 (
        .din(new_Jinkela_wire_3237),
        .dout(new_Jinkela_wire_3238)
    );

    bfr new_Jinkela_buffer_3210 (
        .din(new_Jinkela_wire_4583),
        .dout(new_Jinkela_wire_4584)
    );

    bfr new_Jinkela_buffer_194 (
        .din(G86),
        .dout(new_Jinkela_wire_503)
    );

    bfr new_Jinkela_buffer_2146 (
        .din(new_Jinkela_wire_3268),
        .dout(new_Jinkela_wire_3269)
    );

    bfr new_Jinkela_buffer_3202 (
        .din(new_Jinkela_wire_4563),
        .dout(new_Jinkela_wire_4564)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_2122 (
        .din(new_Jinkela_wire_3238),
        .dout(new_Jinkela_wire_3239)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    bfr new_Jinkela_buffer_3227 (
        .din(new_Jinkela_wire_4608),
        .dout(new_Jinkela_wire_4609)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_363),
        .b(new_Jinkela_wire_364),
        .c(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_2147 (
        .din(new_Jinkela_wire_3269),
        .dout(new_Jinkela_wire_3270)
    );

    bfr new_Jinkela_buffer_3203 (
        .din(new_Jinkela_wire_4564),
        .dout(new_Jinkela_wire_4565)
    );

    spl2 new_Jinkela_splitter_72 (
        .a(new_Jinkela_wire_365),
        .b(new_Jinkela_wire_366),
        .c(new_Jinkela_wire_367)
    );

    bfr new_Jinkela_buffer_2123 (
        .din(new_Jinkela_wire_3239),
        .dout(new_Jinkela_wire_3240)
    );

    bfr new_Jinkela_buffer_3211 (
        .din(new_Jinkela_wire_4584),
        .dout(new_Jinkela_wire_4585)
    );

    spl2 new_Jinkela_splitter_423 (
        .a(_0876_),
        .b(new_Jinkela_wire_3308),
        .c(new_Jinkela_wire_3312)
    );

    bfr new_Jinkela_buffer_3204 (
        .din(new_Jinkela_wire_4565),
        .dout(new_Jinkela_wire_4566)
    );

    bfr new_Jinkela_buffer_204 (
        .din(G113),
        .dout(new_Jinkela_wire_521)
    );

    bfr new_Jinkela_buffer_2151 (
        .din(new_Jinkela_wire_3276),
        .dout(new_Jinkela_wire_3277)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    bfr new_Jinkela_buffer_2124 (
        .din(new_Jinkela_wire_3240),
        .dout(new_Jinkela_wire_3241)
    );

    bfr new_Jinkela_buffer_3231 (
        .din(new_Jinkela_wire_4615),
        .dout(new_Jinkela_wire_4616)
    );

    bfr new_Jinkela_buffer_2148 (
        .din(new_Jinkela_wire_3270),
        .dout(new_Jinkela_wire_3271)
    );

    bfr new_Jinkela_buffer_3205 (
        .din(new_Jinkela_wire_4566),
        .dout(new_Jinkela_wire_4567)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    bfr new_Jinkela_buffer_2125 (
        .din(new_Jinkela_wire_3241),
        .dout(new_Jinkela_wire_3242)
    );

    bfr new_Jinkela_buffer_3212 (
        .din(new_Jinkela_wire_4585),
        .dout(new_Jinkela_wire_4586)
    );

    spl2 new_Jinkela_splitter_106 (
        .a(new_Jinkela_wire_505),
        .b(new_Jinkela_wire_506),
        .c(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_2176 (
        .din(new_Jinkela_wire_3306),
        .dout(new_Jinkela_wire_3307)
    );

    bfr new_Jinkela_buffer_3279 (
        .din(new_net_2359),
        .dout(new_Jinkela_wire_4666)
    );

    bfr new_Jinkela_buffer_3228 (
        .din(new_Jinkela_wire_4609),
        .dout(new_Jinkela_wire_4610)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    bfr new_Jinkela_buffer_2126 (
        .din(new_Jinkela_wire_3242),
        .dout(new_Jinkela_wire_3243)
    );

    bfr new_Jinkela_buffer_3213 (
        .din(new_Jinkela_wire_4586),
        .dout(new_Jinkela_wire_4587)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    spl3L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_369),
        .d(new_Jinkela_wire_370),
        .b(new_Jinkela_wire_371),
        .c(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_2149 (
        .din(new_Jinkela_wire_3271),
        .dout(new_Jinkela_wire_3272)
    );

    bfr new_Jinkela_buffer_2127 (
        .din(new_Jinkela_wire_3243),
        .dout(new_Jinkela_wire_3244)
    );

    bfr new_Jinkela_buffer_3214 (
        .din(new_Jinkela_wire_4587),
        .dout(new_Jinkela_wire_4588)
    );

    bfr new_Jinkela_buffer_205 (
        .din(G108),
        .dout(new_Jinkela_wire_529)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_2177 (
        .din(_0345_),
        .dout(new_Jinkela_wire_3317)
    );

    bfr new_Jinkela_buffer_3229 (
        .din(new_Jinkela_wire_4610),
        .dout(new_Jinkela_wire_4611)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_2128 (
        .din(new_Jinkela_wire_3244),
        .dout(new_Jinkela_wire_3245)
    );

    bfr new_Jinkela_buffer_3215 (
        .din(new_Jinkela_wire_4588),
        .dout(new_Jinkela_wire_4589)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_373),
        .b(new_Jinkela_wire_374),
        .c(new_Jinkela_wire_375)
    );

    bfr new_Jinkela_buffer_2150 (
        .din(new_Jinkela_wire_3272),
        .dout(new_Jinkela_wire_3273)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_2129 (
        .din(new_Jinkela_wire_3245),
        .dout(new_Jinkela_wire_3246)
    );

    bfr new_Jinkela_buffer_3216 (
        .din(new_Jinkela_wire_4589),
        .dout(new_Jinkela_wire_4590)
    );

    bfr new_Jinkela_buffer_2153 (
        .din(new_Jinkela_wire_3283),
        .dout(new_Jinkela_wire_3284)
    );

    bfr new_Jinkela_buffer_3270 (
        .din(new_Jinkela_wire_4656),
        .dout(new_Jinkela_wire_4657)
    );

    bfr new_Jinkela_buffer_3232 (
        .din(new_Jinkela_wire_4616),
        .dout(new_Jinkela_wire_4617)
    );

    bfr new_Jinkela_buffer_2130 (
        .din(new_Jinkela_wire_3246),
        .dout(new_Jinkela_wire_3247)
    );

    bfr new_Jinkela_buffer_3217 (
        .din(new_Jinkela_wire_4590),
        .dout(new_Jinkela_wire_4591)
    );

    spl4L new_Jinkela_splitter_75 (
        .a(new_Jinkela_wire_376),
        .d(new_Jinkela_wire_377),
        .e(new_Jinkela_wire_378),
        .b(new_Jinkela_wire_379),
        .c(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_2180 (
        .din(new_net_2507),
        .dout(new_Jinkela_wire_3320)
    );

    and_ii _1571_ (
        .a(_0866_),
        .b(_0865_),
        .c(_0867_)
    );

    and_bi _2285_ (
        .a(new_Jinkela_wire_664),
        .b(_0300_),
        .c(new_net_2397)
    );

    and_bi _1572_ (
        .a(new_Jinkela_wire_952),
        .b(new_Jinkela_wire_3171),
        .c(_0868_)
    );

    or_ii _2286_ (
        .a(new_Jinkela_wire_5913),
        .b(new_Jinkela_wire_3455),
        .c(_0301_)
    );

    or_bi _1573_ (
        .a(new_Jinkela_wire_5297),
        .b(new_Jinkela_wire_5634),
        .c(_0869_)
    );

    and_bi _2287_ (
        .a(new_Jinkela_wire_2068),
        .b(new_Jinkela_wire_3451),
        .c(_0302_)
    );

    and_bi _1574_ (
        .a(_0869_),
        .b(new_Jinkela_wire_6767),
        .c(_0870_)
    );

    or_bb _2288_ (
        .a(_0302_),
        .b(new_Jinkela_wire_3510),
        .c(_0303_)
    );

    and_ii _1575_ (
        .a(new_Jinkela_wire_5296),
        .b(new_Jinkela_wire_6764),
        .c(_0871_)
    );

    and_bi _2289_ (
        .a(_0301_),
        .b(_0303_),
        .c(_0304_)
    );

    and_bi _1576_ (
        .a(new_Jinkela_wire_3170),
        .b(new_Jinkela_wire_953),
        .c(_0872_)
    );

    and_bi _2290_ (
        .a(new_Jinkela_wire_180),
        .b(new_Jinkela_wire_2874),
        .c(_0305_)
    );

    and_ii _1577_ (
        .a(new_Jinkela_wire_7111),
        .b(new_Jinkela_wire_5632),
        .c(_0873_)
    );

    and_bi _2291_ (
        .a(new_Jinkela_wire_722),
        .b(new_Jinkela_wire_6423),
        .c(_0306_)
    );

    and_bb _1578_ (
        .a(new_Jinkela_wire_3356),
        .b(new_Jinkela_wire_1861),
        .c(_0874_)
    );

    or_bb _2292_ (
        .a(_0306_),
        .b(_0305_),
        .c(_0307_)
    );

    and_bi _1579_ (
        .a(new_Jinkela_wire_1954),
        .b(new_Jinkela_wire_5415),
        .c(_0875_)
    );

    or_bb _2293_ (
        .a(new_Jinkela_wire_5357),
        .b(_0304_),
        .c(new_net_2437)
    );

    and_ii _1580_ (
        .a(_0875_),
        .b(new_Jinkela_wire_6933),
        .c(_0876_)
    );

    or_ii _2294_ (
        .a(new_Jinkela_wire_5883),
        .b(new_Jinkela_wire_3453),
        .c(_0308_)
    );

    and_bi _1581_ (
        .a(new_Jinkela_wire_2581),
        .b(new_Jinkela_wire_3314),
        .c(_0877_)
    );

    and_bi _2295_ (
        .a(new_Jinkela_wire_4054),
        .b(new_Jinkela_wire_3448),
        .c(_0309_)
    );

    and_bi _1582_ (
        .a(new_Jinkela_wire_6224),
        .b(_0877_),
        .c(_0878_)
    );

    or_bb _2296_ (
        .a(_0309_),
        .b(new_Jinkela_wire_3507),
        .c(_0310_)
    );

    or_ii _1583_ (
        .a(new_Jinkela_wire_4340),
        .b(new_Jinkela_wire_4598),
        .c(_0879_)
    );

    and_bi _2297_ (
        .a(_0308_),
        .b(new_Jinkela_wire_3664),
        .c(_0311_)
    );

    and_ii _1584_ (
        .a(new_Jinkela_wire_4341),
        .b(new_Jinkela_wire_4599),
        .c(_0880_)
    );

    and_bi _2298_ (
        .a(new_Jinkela_wire_241),
        .b(new_Jinkela_wire_6415),
        .c(_0312_)
    );

    and_bi _1585_ (
        .a(_0879_),
        .b(_0880_),
        .c(_0881_)
    );

    and_bi _2299_ (
        .a(new_Jinkela_wire_1436),
        .b(new_Jinkela_wire_2869),
        .c(_0313_)
    );

    or_bb _1586_ (
        .a(new_Jinkela_wire_5236),
        .b(new_Jinkela_wire_1094),
        .c(_0882_)
    );

    or_bb _2300_ (
        .a(_0313_),
        .b(_0312_),
        .c(_0314_)
    );

    or_bb _2301_ (
        .a(new_Jinkela_wire_7992),
        .b(_0311_),
        .c(new_net_2501)
    );

    or_bb _1587_ (
        .a(new_Jinkela_wire_1396),
        .b(new_Jinkela_wire_42),
        .c(_0883_)
    );

    or_ii _2302_ (
        .a(new_Jinkela_wire_7941),
        .b(new_Jinkela_wire_3452),
        .c(_0315_)
    );

    and_bi _1588_ (
        .a(new_Jinkela_wire_1397),
        .b(new_Jinkela_wire_403),
        .c(_0884_)
    );

    and_bi _2303_ (
        .a(new_Jinkela_wire_7293),
        .b(new_Jinkela_wire_3444),
        .c(_0316_)
    );

    and_bi _1589_ (
        .a(_0883_),
        .b(_0884_),
        .c(_0885_)
    );

    or_bb _2304_ (
        .a(_0316_),
        .b(new_Jinkela_wire_3504),
        .c(_0317_)
    );

    and_bi _1590_ (
        .a(new_Jinkela_wire_1036),
        .b(new_Jinkela_wire_4336),
        .c(_0886_)
    );

    and_bi _2305_ (
        .a(_0315_),
        .b(new_Jinkela_wire_6249),
        .c(_0318_)
    );

    or_bb _1591_ (
        .a(_0886_),
        .b(new_Jinkela_wire_4820),
        .c(_0887_)
    );

    and_bi _2306_ (
        .a(new_Jinkela_wire_1193),
        .b(new_Jinkela_wire_2872),
        .c(_0319_)
    );

    and_bi _1592_ (
        .a(_0882_),
        .b(new_Jinkela_wire_5686),
        .c(_0888_)
    );

    and_bi _2307_ (
        .a(new_Jinkela_wire_150),
        .b(new_Jinkela_wire_6422),
        .c(_0320_)
    );

    and_ii _1593_ (
        .a(_0888_),
        .b(new_Jinkela_wire_6406),
        .c(new_net_19)
    );

    or_bb _2308_ (
        .a(_0320_),
        .b(_0319_),
        .c(_0321_)
    );

    and_bi _1594_ (
        .a(new_Jinkela_wire_967),
        .b(new_Jinkela_wire_6690),
        .c(_0889_)
    );

    and_ii _1595_ (
        .a(new_Jinkela_wire_3316),
        .b(new_Jinkela_wire_7127),
        .c(_0890_)
    );

    or_bb _2309_ (
        .a(new_Jinkela_wire_2898),
        .b(_0318_),
        .c(new_net_2383)
    );

    or_ii _2310_ (
        .a(new_Jinkela_wire_2428),
        .b(new_Jinkela_wire_3445),
        .c(_0322_)
    );

    and_bi _1596_ (
        .a(new_Jinkela_wire_3313),
        .b(new_Jinkela_wire_5651),
        .c(_0891_)
    );

    and_bi _2311_ (
        .a(new_Jinkela_wire_7438),
        .b(new_Jinkela_wire_3440),
        .c(_0323_)
    );

    or_bb _1597_ (
        .a(_0891_),
        .b(_0890_),
        .c(_0892_)
    );

    or_bb _2312_ (
        .a(_0323_),
        .b(new_Jinkela_wire_3500),
        .c(_0324_)
    );

    or_bi _1598_ (
        .a(new_Jinkela_wire_5245),
        .b(new_Jinkela_wire_1877),
        .c(_0893_)
    );

    and_bi _2313_ (
        .a(_0322_),
        .b(new_Jinkela_wire_5488),
        .c(_0325_)
    );

    and_bi _1599_ (
        .a(new_Jinkela_wire_5246),
        .b(new_Jinkela_wire_1878),
        .c(_0894_)
    );

    and_bi _2314_ (
        .a(new_Jinkela_wire_1247),
        .b(new_Jinkela_wire_2875),
        .c(_0326_)
    );

    and_bi _1600_ (
        .a(_0893_),
        .b(_0894_),
        .c(_0895_)
    );

    and_bi _2315_ (
        .a(new_Jinkela_wire_1610),
        .b(new_Jinkela_wire_6425),
        .c(_0327_)
    );

    or_bb _1601_ (
        .a(new_Jinkela_wire_5395),
        .b(new_Jinkela_wire_1095),
        .c(_0896_)
    );

    or_bb _2316_ (
        .a(_0327_),
        .b(_0326_),
        .c(_0328_)
    );

    inv _1602_ (
        .din(new_Jinkela_wire_756),
        .dout(_0897_)
    );

    or_bb _2317_ (
        .a(new_Jinkela_wire_3609),
        .b(_0325_),
        .c(new_net_2369)
    );

    or_bb _1603_ (
        .a(new_Jinkela_wire_170),
        .b(new_Jinkela_wire_44),
        .c(_0898_)
    );

    or_bi _2318_ (
        .a(new_Jinkela_wire_381),
        .b(new_Jinkela_wire_5911),
        .c(_0329_)
    );

    and_bi _1604_ (
        .a(new_Jinkela_wire_174),
        .b(new_Jinkela_wire_404),
        .c(_0899_)
    );

    and_bb _2319_ (
        .a(new_Jinkela_wire_2065),
        .b(new_Jinkela_wire_378),
        .c(_0330_)
    );

    and_bi _1605_ (
        .a(_0898_),
        .b(_0899_),
        .c(_0900_)
    );

    or_bb _2320_ (
        .a(_0330_),
        .b(new_Jinkela_wire_3974),
        .c(_0331_)
    );

    or_bb _1606_ (
        .a(_0900_),
        .b(new_Jinkela_wire_1881),
        .c(_0901_)
    );

    and_bi _2321_ (
        .a(_0329_),
        .b(_0331_),
        .c(_0332_)
    );

    or_ii _1607_ (
        .a(new_Jinkela_wire_169),
        .b(new_Jinkela_wire_1196),
        .c(_0902_)
    );

    and_bi _2322_ (
        .a(new_Jinkela_wire_723),
        .b(new_Jinkela_wire_7871),
        .c(_0333_)
    );

    and_bi _1608_ (
        .a(new_Jinkela_wire_1528),
        .b(new_Jinkela_wire_173),
        .c(_0903_)
    );

    and_bi _2323_ (
        .a(new_Jinkela_wire_181),
        .b(new_Jinkela_wire_5809),
        .c(_0334_)
    );

    and_bi _1609_ (
        .a(_0902_),
        .b(_0903_),
        .c(_0904_)
    );

    and_bi _1610_ (
        .a(new_Jinkela_wire_1880),
        .b(_0904_),
        .c(_0905_)
    );

    or_bb _2324_ (
        .a(_0334_),
        .b(_0333_),
        .c(_0335_)
    );

    and_bi _1611_ (
        .a(_0901_),
        .b(_0905_),
        .c(_0906_)
    );

    and_bi _1612_ (
        .a(new_Jinkela_wire_1043),
        .b(new_Jinkela_wire_7143),
        .c(_0907_)
    );

endmodule
