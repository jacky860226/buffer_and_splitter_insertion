module c432(N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432);
	wire new_net_346;
	wire new_net_762;
	wire new_net_721;
	wire new_net_802;
	wire new_net_810;
	wire new_net_556;
	wire new_net_603;
	wire new_net_729;
	wire _011_;
	wire _095_;
	wire new_net_2;
	wire new_net_17;
	wire new_net_50;
	wire new_net_65;
	wire new_net_131;
	wire new_net_146;
	wire new_net_390;
	wire new_net_424;
	wire new_net_518;
	wire new_net_814;
	wire new_net_801;
	wire new_net_365;
	wire new_net_737;
	wire new_net_525;
	wire new_net_696;
	wire new_net_822;
	wire new_net_655;
	wire _032_;
	wire _074_;
	wire _116_;
	wire new_net_41;
	wire new_net_122;
	wire new_net_104;
	wire new_net_188;
	wire new_net_396;
	wire new_net_418;
	wire new_net_430;
	wire new_net_497;
	wire new_net_866;
	wire _053_;
	wire new_net_96;
	wire new_net_380;
	wire new_net_402;
	wire new_net_413;
	wire new_net_436;
	wire new_net_459;
	wire new_net_493;
	wire new_net_526;
	wire new_net_537;
	wire new_net_663;
	wire new_net_750;
	wire new_net_917;
	wire new_net_582;
	wire new_net_958;
	wire new_net_191;
	wire new_net_796;
	wire new_net_342;
	wire new_net_460;
	wire new_net_385;
	wire new_net_407;
	wire new_net_442;
	wire new_net_476;
	wire new_net_510;
	wire new_net_521;
	wire new_net_542;
	wire new_net_565;
	wire new_net_599;
	wire new_net_634;
	wire new_net_676;
	wire _012_;
	wire _096_;
	wire new_net_183;
	wire new_net_250;
	wire new_net_261;
	wire new_net_272;
	wire new_net_283;
	wire new_net_513;
	wire new_net_596;
	wire new_net_640;
	wire new_net_359;
	wire new_net_649;
	wire new_net_73;
	wire new_net_139;
	wire _033_;
	wire _075_;
	wire new_net_10;
	wire new_net_25;
	wire new_net_58;
	wire new_net_154;
	wire new_net_206;
	wire new_net_245;
	wire new_net_439;
	wire new_net_562;
	wire new_net_688;
	wire new_net_861;
	wire new_net_859;
	wire _054_;
	wire new_net_921;
	wire new_net_775;
	wire new_net_933;
	wire new_net_657;
	wire new_net_905;
	wire new_net_945;
	wire new_net_864;
	wire new_net_576;
	wire new_net_743;
	wire new_net_952;
	wire new_net_702;
	wire new_net_372;
	wire new_net_828;
	wire new_net_574;
	wire new_net_168;
	wire new_net_200;
	wire new_net_927;
	wire new_net_939;
	wire new_net_972;
	wire new_net_793;
	wire new_net_990;
	wire new_net_709;
	wire _013_;
	wire _097_;
	wire new_net_18;
	wire new_net_33;
	wire new_net_66;
	wire new_net_81;
	wire new_net_147;
	wire new_net_515;
	wire new_net_835;
	wire new_net_590;
	wire new_net_885;
	wire new_net_966;
	wire new_net_42;
	wire new_net_123;
	wire _034_;
	wire _076_;
	wire new_net_105;
	wire new_net_178;
	wire new_net_374;
	wire new_net_682;
	wire new_net_767;
	wire new_net_889;
	wire _055_;
	wire new_net_210;
	wire new_net_226;
	wire new_net_237;
	wire new_net_293;
	wire new_net_321;
	wire new_net_332;
	wire new_net_353;
	wire new_net_364;
	wire new_net_561;
	wire new_net_855;
	wire new_net_734;
	wire new_net_902;
	wire new_net_445;
	wire new_net_286;
	wire new_net_221;
	wire new_net_266;
	wire new_net_305;
	wire new_net_316;
	wire new_net_337;
	wire new_net_348;
	wire new_net_369;
	wire new_net_781;
	wire new_net_616;
	wire new_net_787;
	wire new_net_530;
	wire _056_;
	wire _014_;
	wire _098_;
	wire new_net_241;
	wire new_net_300;
	wire new_net_453;
	wire new_net_624;
	wire new_net_704;
	wire new_net_716;
	wire new_net_715;
	wire new_net_871;
	wire new_net_911;
	wire new_net_841;
	wire new_net_960;
	wire new_net_89;
	wire new_net_155;
	wire _035_;
	wire _077_;
	wire new_net_26;
	wire new_net_74;
	wire new_net_162;
	wire new_net_165;
	wire new_net_201;
	wire new_net_202;
	wire new_net_345;
	wire new_net_504;
	wire new_net_587;
	wire new_net_761;
	wire new_net_549;
	wire new_net_720;
	wire new_net_3;
	wire new_net_51;
	wire new_net_132;
	wire new_net_391;
	wire new_net_425;
	wire new_net_448;
	wire new_net_471;
	wire new_net_482;
	wire new_net_505;
	wire new_net_560;
	wire new_net_809;
	wire new_net_749;
	wire new_net_969;
	wire new_net_606;
	wire new_net_602;
	wire new_net_728;
	wire new_net_896;
	wire new_net_517;
	wire new_net_813;
	wire new_net_397;
	wire new_net_419;
	wire new_net_431;
	wire new_net_454;
	wire new_net_465;
	wire new_net_488;
	wire new_net_499;
	wire new_net_554;
	wire new_net_577;
	wire new_net_589;
	wire new_net_695;
	wire new_net_821;
	wire new_net_97;
	wire new_net_115;
	wire new_net_170;
	wire new_net_82;
	wire _015_;
	wire _099_;
	wire new_net_34;
	wire new_net_215;
	wire new_net_288;
	wire new_net_310;
	wire new_net_654;
	wire new_net_865;
	wire new_net_492;
	wire new_net_536;
	wire new_net_662;
	wire new_net_189;
	wire _078_;
	wire new_net_43;
	wire new_net_106;
	wire new_net_124;
	wire new_net_231;
	wire new_net_326;
	wire new_net_358;
	wire new_net_375;
	wire new_net_386;
	wire new_net_498;
	wire new_net_581;
	wire new_net_622;
	wire new_net_747;
	wire new_net_957;
	wire new_net_543;
	wire _057_;
	wire new_net_211;
	wire new_net_251;
	wire new_net_262;
	wire new_net_273;
	wire new_net_294;
	wire new_net_618;
	wire new_net_628;
	wire new_net_641;
	wire new_net_664;
	wire new_net_675;
	wire new_net_595;
	wire _036_;
	wire new_net_11;
	wire new_net_59;
	wire new_net_140;
	wire new_net_207;
	wire new_net_246;
	wire new_net_257;
	wire new_net_267;
	wire new_net_278;
	wire new_net_289;
	wire _016_;
	wire _100_;
	wire new_net_184;
	wire new_net_196;
	wire new_net_314;
	wire new_net_648;
	wire new_net_774;
	wire new_net_922;
	wire new_net_687;
	wire new_net_934;
	wire new_net_795;
	wire new_net_858;
	wire new_net_944;
	wire _037_;
	wire _079_;
	wire new_net_90;
	wire new_net_167;
	wire new_net_928;
	wire new_net_940;
	wire new_net_973;
	wire new_net_951;
	wire new_net_701;
	wire _058_;
	wire new_net_4;
	wire new_net_19;
	wire new_net_52;
	wire new_net_67;
	wire new_net_133;
	wire new_net_148;
	wire new_net_172;
	wire new_net_827;
	wire new_net_897;
	wire new_net_792;
	wire new_net_670;
	wire new_net_989;
	wire new_net_834;
	wire new_net_877;
	wire new_net_668;
	wire new_net_671;
	wire new_net_916;
	wire new_net_532;
	wire new_net_983;
	wire new_net_995;
	wire new_net_884;
	wire new_net_846;
	wire _017_;
	wire _101_;
	wire new_net_98;
	wire new_net_216;
	wire new_net_227;
	wire new_net_238;
	wire new_net_311;
	wire new_net_322;
	wire new_net_333;
	wire new_net_229;
	wire new_net_681;
	wire new_net_847;
	wire new_net_930;
	wire new_net_766;
	wire new_net_738;
	wire new_net_853;
	wire _038_;
	wire _080_;
	wire new_net_44;
	wire new_net_107;
	wire new_net_179;
	wire new_net_125;
	wire new_net_232;
	wire new_net_306;
	wire new_net_317;
	wire new_net_327;
	wire new_net_733;
	wire new_net_901;
	wire _059_;
	wire new_net_978;
	wire new_net_780;
	wire new_net_368;
	wire new_net_615;
	wire new_net_786;
	wire new_net_405;
	wire new_net_529;
	wire new_net_700;
	wire new_net_256;
	wire new_net_299;
	wire new_net_703;
	wire new_net_910;
	wire new_net_870;
	wire new_net_12;
	wire new_net_27;
	wire new_net_60;
	wire new_net_75;
	wire new_net_141;
	wire new_net_156;
	wire new_net_642;
	wire new_net_171;
	wire _018_;
	wire _102_;
	wire new_net_174;
	wire new_net_392;
	wire new_net_426;
	wire new_net_449;
	wire new_net_472;
	wire new_net_483;
	wire new_net_503;
	wire new_net_588;
	wire new_net_959;
	wire new_net_586;
	wire new_net_344;
	wire new_net_388;
	wire new_net_760;
	wire new_net_548;
	wire new_net_719;
	wire new_net_800;
	wire new_net_633;
	wire new_net_758;
	wire new_net_636;
	wire new_net_808;
	wire _039_;
	wire _081_;
	wire new_net_398;
	wire new_net_420;
	wire new_net_432;
	wire new_net_466;
	wire new_net_470;
	wire new_net_489;
	wire new_net_500;
	wire new_net_555;
	wire new_net_601;
	wire new_net_727;
	wire new_net_754;
	wire new_net_895;
	wire new_net_516;
	wire new_net_812;
	wire _060_;
	wire new_net_20;
	wire new_net_35;
	wire new_net_68;
	wire new_net_83;
	wire new_net_116;
	wire new_net_149;
	wire new_net_404;
	wire new_net_438;
	wire new_net_495;
	wire new_net_970;
	wire new_net_783;
	wire new_net_357;
	wire new_net_694;
	wire new_net_820;
	wire new_net_653;
	wire new_net_376;
	wire new_net_387;
	wire new_net_409;
	wire new_net_455;
	wire new_net_478;
	wire new_net_512;
	wire new_net_523;
	wire new_net_533;
	wire new_net_544;
	wire new_net_567;
	wire new_net_661;
	wire new_net_909;
	wire _019_;
	wire _103_;
	wire new_net_212;
	wire new_net_252;
	wire new_net_263;
	wire new_net_274;
	wire new_net_295;
	wire new_net_619;
	wire new_net_623;
	wire new_net_665;
	wire new_net_748;
	wire new_net_580;
	wire new_net_621;
	wire new_net_746;
	wire new_net_956;
	wire new_net_794;
	wire new_net_627;
	wire new_net_108;
	wire new_net_190;
	wire _040_;
	wire _082_;
	wire new_net_45;
	wire new_net_126;
	wire new_net_208;
	wire new_net_247;
	wire new_net_268;
	wire new_net_279;
	wire new_net_464;
	wire new_net_674;
	wire new_net_713;
	wire new_net_881;
	wire new_net_511;
	wire _061_;
	wire new_net_635;
	wire new_net_923;
	wire new_net_594;
	wire new_net_935;
	wire new_net_313;
	wire new_net_647;
	wire new_net_773;
	wire new_net_437;
	wire new_net_686;
	wire new_net_28;
	wire new_net_76;
	wire new_net_91;
	wire new_net_157;
	wire new_net_929;
	wire new_net_941;
	wire new_net_974;
	wire new_net_857;
	wire new_net_185;
	wire new_net_134;
	wire _020_;
	wire _104_;
	wire new_net_5;
	wire new_net_53;
	wire new_net_240;
	wire new_net_325;
	wire new_net_381;
	wire new_net_943;
	wire new_net_741;
	wire new_net_950;
	wire new_net_826;
	wire new_net_370;
	wire new_net_572;
	wire new_net_414;
	wire _041_;
	wire _083_;
	wire new_net_984;
	wire new_net_791;
	wire new_net_996;
	wire new_net_669;
	wire new_net_988;
	wire new_net_833;
	wire new_net_876;
	wire new_net_297;
	wire _062_;
	wire new_net_36;
	wire new_net_84;
	wire new_net_99;
	wire new_net_117;
	wire new_net_203;
	wire new_net_217;
	wire new_net_228;
	wire new_net_239;
	wire new_net_284;
	wire new_net_883;
	wire new_net_845;
	wire new_net_964;
	wire new_net_680;
	wire new_net_233;
	wire new_net_307;
	wire new_net_328;
	wire new_net_339;
	wire new_net_360;
	wire new_net_371;
	wire new_net_765;
	wire new_net_724;
	wire new_net_852;
	wire _021_;
	wire _105_;
	wire new_net_559;
	wire new_net_979;
	wire new_net_732;
	wire new_net_900;
	wire new_net_965;
	wire new_net_779;
	wire _000_;
	wire _042_;
	wire _084_;
	wire new_net_13;
	wire new_net_46;
	wire new_net_61;
	wire new_net_109;
	wire new_net_127;
	wire new_net_142;
	wire new_net_180;
	wire new_net_367;
	wire new_net_528;
	wire new_net_614;
	wire new_net_699;
	wire new_net_977;
	wire _063_;
	wire new_net_393;
	wire new_net_415;
	wire new_net_427;
	wire new_net_450;
	wire new_net_484;
	wire new_net_507;
	wire new_net_573;
	wire new_net_585;
	wire new_net_607;
	wire new_net_829;
	wire new_net_869;
	wire new_net_872;
	wire new_net_496;
	wire new_net_540;
	wire new_net_915;
	wire new_net_714;
	wire new_net_839;
	wire new_net_502;
	wire new_net_92;
	wire new_net_399;
	wire new_net_421;
	wire new_net_433;
	wire new_net_343;
	wire new_net_444;
	wire new_net_467;
	wire new_net_490;
	wire new_net_501;
	wire new_net_547;
	wire new_net_718;
	wire new_net_759;
	wire new_net_799;
	wire new_net_632;
	wire new_net_757;
	wire _022_;
	wire _106_;
	wire new_net_6;
	wire new_net_21;
	wire new_net_54;
	wire new_net_175;
	wire new_net_135;
	wire new_net_150;
	wire new_net_69;
	wire new_net_382;
	wire new_net_469;
	wire new_net_553;
	wire new_net_551;
	wire new_net_600;
	wire new_net_726;
	wire new_net_894;
	wire _043_;
	wire _001_;
	wire _085_;
	wire new_net_163;
	wire new_net_166;
	wire new_net_222;
	wire new_net_377;
	wire new_net_410;
	wire new_net_456;
	wire new_net_356;
	wire new_net_693;
	wire new_net_819;
	wire new_net_652;
	wire _064_;
	wire new_net_100;
	wire new_net_204;
	wire new_net_213;
	wire new_net_253;
	wire new_net_264;
	wire new_net_285;
	wire new_net_296;
	wire new_net_620;
	wire new_net_666;
	wire new_net_534;
	wire new_net_660;
	wire new_net_908;
	wire new_net_209;
	wire new_net_248;
	wire new_net_269;
	wire new_net_280;
	wire new_net_291;
	wire new_net_338;
	wire new_net_461;
	wire new_net_579;
	wire new_net_637;
	wire new_net_706;
	wire new_net_752;
	wire new_net_955;
	wire new_net_626;
	wire _065_;
	wire _023_;
	wire _107_;
	wire new_net_198;
	wire new_net_924;
	wire new_net_936;
	wire new_net_712;
	wire new_net_593;
	wire new_net_926;
	wire _002_;
	wire _044_;
	wire _086_;
	wire new_net_14;
	wire new_net_29;
	wire new_net_62;
	wire new_net_77;
	wire new_net_110;
	wire new_net_143;
	wire new_net_158;
	wire new_net_805;
	wire new_net_849;
	wire new_net_312;
	wire new_net_477;
	wire new_net_479;
	wire new_net_646;
	wire new_net_772;
	wire new_net_685;
	wire new_net_991;
	wire new_net_770;
	wire new_net_892;
	wire new_net_856;
	wire new_net_481;
	wire new_net_942;
	wire new_net_324;
	wire new_net_985;
	wire new_net_997;
	wire new_net_740;
	wire new_net_949;
	wire new_net_825;
	wire new_net_571;
	wire new_net_85;
	wire new_net_151;
	wire new_net_70;
	wire _024_;
	wire _066_;
	wire _108_;
	wire new_net_22;
	wire new_net_37;
	wire new_net_118;
	wire new_net_186;
	wire new_net_785;
	wire new_net_790;
	wire new_net_707;
	wire new_net_832;
	wire new_net_875;
	wire new_net_914;
	wire new_net_708;
	wire new_net_550;
	wire _003_;
	wire _045_;
	wire _087_;
	wire new_net_223;
	wire new_net_234;
	wire new_net_258;
	wire new_net_308;
	wire new_net_329;
	wire new_net_340;
	wire new_net_361;
	wire new_net_629;
	wire new_net_844;
	wire new_net_882;
	wire new_net_963;
	wire new_net_101;
	wire new_net_753;
	wire new_net_811;
	wire new_net_980;
	wire new_net_967;
	wire new_net_764;
	wire new_net_723;
	wire new_net_851;
	wire new_net_558;
	wire new_net_0;
	wire new_net_47;
	wire new_net_128;
	wire new_net_605;
	wire new_net_679;
	wire new_net_731;
	wire new_net_782;
	wire new_net_899;
	wire new_net_644;
	wire new_net_816;
	wire new_net_778;
	wire _067_;
	wire _025_;
	wire _109_;
	wire new_net_394;
	wire new_net_416;
	wire new_net_428;
	wire new_net_451;
	wire new_net_462;
	wire new_net_485;
	wire new_net_508;
	wire new_net_609;
	wire new_net_613;
	wire new_net_784;
	wire new_net_975;
	wire new_net_403;
	wire new_net_527;
	wire new_net_698;
	wire new_net_868;
	wire new_net_181;
	wire _004_;
	wire _046_;
	wire _088_;
	wire new_net_30;
	wire new_net_78;
	wire new_net_93;
	wire new_net_111;
	wire new_net_159;
	wire new_net_422;
	wire new_net_539;
	wire new_net_7;
	wire new_net_55;
	wire new_net_136;
	wire new_net_302;
	wire new_net_334;
	wire new_net_366;
	wire new_net_383;
	wire new_net_440;
	wire new_net_474;
	wire new_net_519;
	wire new_net_584;
	wire new_net_336;
	wire new_net_717;
	wire new_net_798;
	wire new_net_631;
	wire new_net_667;
	wire new_net_756;
	wire new_net_806;
	wire new_net_468;
	wire new_net_678;
	wire new_net_318;
	wire new_net_350;
	wire new_net_378;
	wire new_net_400;
	wire new_net_411;
	wire new_net_457;
	wire new_net_491;
	wire new_net_514;
	wire new_net_535;
	wire new_net_546;
	wire new_net_725;
	wire new_net_893;
	wire new_net_176;
	wire new_net_119;
	wire _068_;
	wire _026_;
	wire _110_;
	wire new_net_38;
	wire new_net_86;
	wire new_net_243;
	wire new_net_254;
	wire new_net_265;
	wire new_net_355;
	wire new_net_522;
	wire new_net_568;
	wire new_net_692;
	wire new_net_818;
	wire new_net_651;
	wire new_net_690;
	wire new_net_878;
	wire _047_;
	wire _005_;
	wire _089_;
	wire new_net_173;
	wire new_net_259;
	wire new_net_270;
	wire new_net_281;
	wire new_net_292;
	wire new_net_611;
	wire new_net_638;
	wire new_net_659;
	wire new_net_907;
	wire new_net_925;
	wire new_net_937;
	wire new_net_578;
	wire new_net_954;
	wire new_net_625;
	wire new_net_15;
	wire new_net_48;
	wire new_net_63;
	wire new_net_129;
	wire new_net_144;
	wire new_net_672;
	wire new_net_711;
	wire new_net_837;
	wire new_net_919;
	wire new_net_931;
	wire new_net_592;
	wire new_net_838;
	wire _069_;
	wire _027_;
	wire _111_;
	wire new_net_164;
	wire new_net_161;
	wire new_net_597;
	wire new_net_992;
	wire new_net_887;
	wire new_net_804;
	wire new_net_848;
	wire new_net_645;
	wire new_net_771;
	wire new_net_684;
	wire new_net_769;
	wire new_net_891;
	wire _006_;
	wire _090_;
	wire new_net_94;
	wire new_net_524;
	wire new_net_986;
	wire new_net_998;
	wire new_net_480;
	wire new_net_323;
	wire new_net_566;
	wire new_net_8;
	wire new_net_23;
	wire new_net_56;
	wire new_net_71;
	wire new_net_137;
	wire new_net_152;
	wire new_net_219;
	wire new_net_230;
	wire new_net_275;
	wire new_net_303;
	wire new_net_736;
	wire new_net_739;
	wire new_net_807;
	wire new_net_904;
	wire new_net_948;
	wire new_net_824;
	wire new_net_447;
	wire new_net_570;
	wire new_net_789;
	wire _048_;
	wire new_net_224;
	wire new_net_235;
	wire new_net_309;
	wire new_net_319;
	wire new_net_330;
	wire new_net_341;
	wire new_net_351;
	wire new_net_362;
	wire new_net_373;
	wire new_net_831;
	wire new_net_874;
	wire new_net_913;
	wire _028_;
	wire _070_;
	wire _112_;
	wire new_net_39;
	wire new_net_102;
	wire new_net_120;
	wire new_net_187;
	wire new_net_888;
	wire new_net_981;
	wire new_net_994;
	wire new_net_843;
	wire new_net_962;
	wire new_net_506;
	wire new_net_347;
	wire new_net_763;
	wire _007_;
	wire _049_;
	wire _091_;
	wire new_net_722;
	wire new_net_803;
	wire new_net_850;
	wire new_net_434;
	wire new_net_557;
	wire new_net_854;
	wire _072_;
	wire new_net_169;
	wire new_net_395;
	wire new_net_417;
	wire new_net_429;
	wire new_net_452;
	wire new_net_463;
	wire new_net_486;
	wire new_net_552;
	wire new_net_575;
	wire new_net_604;
	wire new_net_730;
	wire new_net_898;
	wire new_net_643;
	wire new_net_815;
	wire new_net_947;
	wire new_net_777;
	wire new_net_608;
	wire new_net_612;
	wire new_net_16;
	wire new_net_31;
	wire new_net_64;
	wire new_net_79;
	wire new_net_112;
	wire new_net_145;
	wire new_net_242;
	wire new_net_389;
	wire new_net_423;
	wire new_net_435;
	wire new_net_656;
	wire new_net_290;
	wire new_net_697;
	wire new_net_867;
	wire _029_;
	wire _113_;
	wire new_net_384;
	wire new_net_441;
	wire new_net_475;
	wire new_net_509;
	wire new_net_520;
	wire new_net_531;
	wire new_net_564;
	wire new_net_598;
	wire new_net_946;
	wire new_net_494;
	wire new_net_538;
	wire new_net_751;
	wire new_net_583;
	wire _008_;
	wire _050_;
	wire _092_;
	wire new_net_182;
	wire new_net_192;
	wire new_net_335;
	wire new_net_379;
	wire new_net_401;
	wire new_net_412;
	wire new_net_458;
	wire new_net_545;
	wire new_net_630;
	wire new_net_755;
	wire new_net_797;
	wire new_net_840;
	wire _071_;
	wire new_net_24;
	wire new_net_72;
	wire new_net_87;
	wire new_net_153;
	wire new_net_244;
	wire new_net_255;
	wire new_net_276;
	wire new_net_287;
	wire new_net_298;
	wire new_net_677;
	wire new_net_277;
	wire new_net_260;
	wire new_net_271;
	wire new_net_282;
	wire new_net_639;
	wire new_net_354;
	wire new_net_673;
	wire new_net_691;
	wire new_net_742;
	wire new_net_776;
	wire new_net_650;
	wire new_net_817;
	wire new_net_938;
	wire new_net_563;
	wire new_net_689;
	wire new_net_121;
	wire new_net_160;
	wire _030_;
	wire _114_;
	wire new_net_40;
	wire new_net_103;
	wire new_net_177;
	wire new_net_610;
	wire new_net_862;
	wire new_net_860;
	wire new_net_863;
	wire new_net_408;
	wire new_net_658;
	wire new_net_906;
	wire new_net_744;
	wire new_net_49;
	wire new_net_130;
	wire _051_;
	wire _009_;
	wire _093_;
	wire new_net_1;
	wire new_net_194;
	wire new_net_920;
	wire new_net_932;
	wire new_net_745;
	wire new_net_953;
	wire new_net_406;
	wire new_net_541;
	wire new_net_993;
	wire new_net_710;
	wire new_net_836;
	wire new_net_879;
	wire new_net_880;
	wire new_net_591;
	wire new_net_32;
	wire new_net_80;
	wire new_net_95;
	wire new_net_113;
	wire new_net_886;
	wire new_net_349;
	wire new_net_987;
	wire new_net_999;
	wire new_net_683;
	wire new_net_138;
	wire _031_;
	wire _115_;
	wire new_net_9;
	wire new_net_57;
	wire new_net_205;
	wire new_net_214;
	wire new_net_220;
	wire new_net_304;
	wire new_net_315;
	wire new_net_473;
	wire new_net_768;
	wire new_net_890;
	wire new_net_971;
	wire new_net_735;
	wire new_net_903;
	wire _010_;
	wire _094_;
	wire new_net_225;
	wire new_net_236;
	wire new_net_249;
	wire new_net_320;
	wire new_net_331;
	wire new_net_352;
	wire new_net_363;
	wire new_net_443;
	wire new_net_446;
	wire new_net_487;
	wire new_net_569;
	wire new_net_823;
	wire _073_;
	wire new_net_88;
	wire new_net_982;
	wire new_net_617;
	wire new_net_788;
	wire new_net_968;
	wire new_net_301;
	wire new_net_705;
	wire new_net_830;
	wire new_net_873;
	wire new_net_912;
	wire new_net_918;
	wire new_net_218;
	wire _052_;
	wire new_net_976;
	wire new_net_842;
	wire new_net_961;
	input N1;
	input N102;
	input N105;
	input N108;
	input N11;
	input N112;
	input N115;
	input N14;
	input N17;
	input N21;
	input N24;
	input N27;
	input N30;
	input N34;
	input N37;
	input N4;
	input N40;
	input N43;
	input N47;
	input N50;
	input N53;
	input N56;
	input N60;
	input N63;
	input N66;
	input N69;
	input N73;
	input N76;
	input N79;
	input N8;
	input N82;
	input N86;
	input N89;
	input N92;
	input N95;
	input N99;
	output N223;
	output N329;
	output N370;
	output N421;
	output N430;
	output N431;
	output N432;

	or_bi _117_ (
		.a(new_net_169),
		.b(new_net_134),
		.c(_061_)
	);

	and_bi _118_ (
		.a(new_net_148),
		.b(new_net_73),
		.c(_062_)
	);

	and_bi _119_ (
		.a(new_net_116),
		.b(new_net_170),
		.c(_063_)
	);

	and_bi _120_ (
		.a(new_net_146),
		.b(new_net_53),
		.c(_064_)
	);

	and_bi _121_ (
		.a(new_net_27),
		.b(new_net_132),
		.c(_065_)
	);

	and_bi _122_ (
		.a(new_net_57),
		.b(new_net_138),
		.c(_066_)
	);

	or_bb _123_ (
		.a(_066_),
		.b(_065_),
		.c(_067_)
	);

	or_bb _124_ (
		.a(_067_),
		.b(new_net_171),
		.c(_068_)
	);

	and_bi _125_ (
		.a(new_net_35),
		.b(new_net_172),
		.c(_069_)
	);

	and_bi _126_ (
		.a(new_net_63),
		.b(new_net_75),
		.c(_070_)
	);

	or_bb _127_ (
		.a(new_net_173),
		.b(new_net_9),
		.c(_071_)
	);

	and_bi _128_ (
		.a(new_net_112),
		.b(new_net_49),
		.c(_072_)
	);

	and_bi _129_ (
		.a(new_net_142),
		.b(new_net_17),
		.c(_073_)
	);

	or_bb _130_ (
		.a(_073_),
		.b(_072_),
		.c(_074_)
	);

	or_bb _131_ (
		.a(new_net_174),
		.b(_071_),
		.c(_075_)
	);

	or_bb _132_ (
		.a(_075_),
		.b(new_net_175),
		.c(_076_)
	);

	and_bi _133_ (
		.a(new_net_176),
		.b(_076_),
		.c(_077_)
	);

	or_ii _134_ (
		.a(new_net_122),
		.b(new_net_135),
		.c(_078_)
	);

	and_bb _135_ (
		.a(_078_),
		.b(new_net_117),
		.c(_079_)
	);

	or_bi _136_ (
		.a(new_net_124),
		.b(new_net_74),
		.c(_080_)
	);

	or_ii _137_ (
		.a(_080_),
		.b(new_net_149),
		.c(_081_)
	);

	or_bb _138_ (
		.a(new_net_65),
		.b(new_net_47),
		.c(_082_)
	);

	or_bi _139_ (
		.a(new_net_118),
		.b(new_net_139),
		.c(_083_)
	);

	or_ii _140_ (
		.a(_083_),
		.b(new_net_58),
		.c(_084_)
	);

	and_ii _141_ (
		.a(new_net_3),
		.b(new_net_81),
		.c(_085_)
	);

	and_bi _142_ (
		.a(_082_),
		.b(_085_),
		.c(_086_)
	);

	and_ii _143_ (
		.a(new_net_19),
		.b(new_net_25),
		.c(_087_)
	);

	or_bi _144_ (
		.a(new_net_123),
		.b(new_net_18),
		.c(_088_)
	);

	or_ii _145_ (
		.a(_088_),
		.b(new_net_143),
		.c(_089_)
	);

	and_ii _146_ (
		.a(new_net_154),
		.b(new_net_7),
		.c(_090_)
	);

	or_bb _147_ (
		.a(_090_),
		.b(_087_),
		.c(_091_)
	);

	and_bi _148_ (
		.a(_086_),
		.b(_091_),
		.c(_092_)
	);

	or_bi _149_ (
		.a(new_net_119),
		.b(new_net_54),
		.c(_093_)
	);

	or_ii _150_ (
		.a(_093_),
		.b(new_net_147),
		.c(_094_)
	);

	and_ii _151_ (
		.a(new_net_150),
		.b(new_net_31),
		.c(_095_)
	);

	or_bi _152_ (
		.a(new_net_125),
		.b(new_net_133),
		.c(_096_)
	);

	or_ii _153_ (
		.a(_096_),
		.b(new_net_28),
		.c(_097_)
	);

	and_ii _154_ (
		.a(new_net_67),
		.b(new_net_55),
		.c(_098_)
	);

	or_bb _155_ (
		.a(_098_),
		.b(_095_),
		.c(_099_)
	);

	or_bi _156_ (
		.a(new_net_126),
		.b(new_net_50),
		.c(_100_)
	);

	or_ii _157_ (
		.a(_100_),
		.b(new_net_113),
		.c(_101_)
	);

	and_ii _158_ (
		.a(new_net_33),
		.b(new_net_144),
		.c(_102_)
	);

	or_ii _159_ (
		.a(new_net_120),
		.b(new_net_36),
		.c(_103_)
	);

	and_bi _160_ (
		.a(_103_),
		.b(new_net_10),
		.c(_104_)
	);

	and_ii _161_ (
		.a(new_net_136),
		.b(new_net_91),
		.c(_105_)
	);

	or_bi _162_ (
		.a(new_net_127),
		.b(new_net_76),
		.c(_106_)
	);

	or_ii _163_ (
		.a(_106_),
		.b(new_net_64),
		.c(_107_)
	);

	and_ii _164_ (
		.a(new_net_51),
		.b(new_net_21),
		.c(_108_)
	);

	or_bb _165_ (
		.a(_108_),
		.b(_105_),
		.c(_109_)
	);

	or_bb _166_ (
		.a(_109_),
		.b(new_net_177),
		.c(_110_)
	);

	or_bb _167_ (
		.a(_110_),
		.b(new_net_178),
		.c(_111_)
	);

	and_bi _168_ (
		.a(new_net_179),
		.b(_111_),
		.c(_112_)
	);

	and_bi _169_ (
		.a(new_net_26),
		.b(new_net_37),
		.c(_113_)
	);

	or_bb _170_ (
		.a(_113_),
		.b(new_net_20),
		.c(_114_)
	);

	or_bb _171_ (
		.a(new_net_97),
		.b(new_net_15),
		.c(_115_)
	);

	and_bi _172_ (
		.a(new_net_56),
		.b(new_net_43),
		.c(_116_)
	);

	or_bb _173_ (
		.a(_116_),
		.b(new_net_68),
		.c(_000_)
	);

	and_ii _174_ (
		.a(new_net_1),
		.b(new_net_93),
		.c(_001_)
	);

	and_bi _175_ (
		.a(new_net_8),
		.b(new_net_39),
		.c(_002_)
	);

	or_bb _176_ (
		.a(_002_),
		.b(new_net_155),
		.c(_003_)
	);

	and_ii _177_ (
		.a(new_net_85),
		.b(new_net_89),
		.c(_004_)
	);

	or_bb _178_ (
		.a(_004_),
		.b(_001_),
		.c(_005_)
	);

	and_bi _179_ (
		.a(new_net_180),
		.b(_005_),
		.c(_006_)
	);

	and_bi _180_ (
		.a(new_net_32),
		.b(new_net_42),
		.c(_007_)
	);

	or_bb _181_ (
		.a(_007_),
		.b(new_net_151),
		.c(_008_)
	);

	and_ii _182_ (
		.a(new_net_77),
		.b(new_net_95),
		.c(_009_)
	);

	and_bi _183_ (
		.a(new_net_82),
		.b(new_net_38),
		.c(_010_)
	);

	or_bb _184_ (
		.a(_010_),
		.b(new_net_4),
		.c(_011_)
	);

	and_ii _185_ (
		.a(new_net_11),
		.b(new_net_152),
		.c(_012_)
	);

	or_bb _186_ (
		.a(_012_),
		.b(_009_),
		.c(_013_)
	);

	and_bi _187_ (
		.a(new_net_92),
		.b(new_net_40),
		.c(_014_)
	);

	or_bb _188_ (
		.a(_014_),
		.b(new_net_137),
		.c(_015_)
	);

	and_ii _189_ (
		.a(new_net_140),
		.b(new_net_158),
		.c(_016_)
	);

	and_bi _190_ (
		.a(new_net_145),
		.b(new_net_44),
		.c(_017_)
	);

	or_bb _191_ (
		.a(_017_),
		.b(new_net_34),
		.c(_018_)
	);

	and_ii _192_ (
		.a(new_net_59),
		.b(new_net_181),
		.c(_019_)
	);

	or_bb _193_ (
		.a(new_net_83),
		.b(new_net_182),
		.c(_020_)
	);

	and_bi _194_ (
		.a(new_net_22),
		.b(new_net_45),
		.c(_021_)
	);

	or_bb _195_ (
		.a(_021_),
		.b(new_net_52),
		.c(_022_)
	);

	and_ii _196_ (
		.a(new_net_29),
		.b(new_net_71),
		.c(_023_)
	);

	and_bi _197_ (
		.a(new_net_48),
		.b(new_net_41),
		.c(_024_)
	);

	or_bb _198_ (
		.a(_024_),
		.b(new_net_66),
		.c(_025_)
	);

	and_ii _199_ (
		.a(new_net_130),
		.b(new_net_69),
		.c(_026_)
	);

	or_bb _200_ (
		.a(_026_),
		.b(_023_),
		.c(_027_)
	);

	or_bb _201_ (
		.a(new_net_183),
		.b(_020_),
		.c(_028_)
	);

	or_bb _202_ (
		.a(_028_),
		.b(new_net_184),
		.c(_029_)
	);

	and_bi _203_ (
		.a(new_net_185),
		.b(_029_),
		.c(_030_)
	);

	inv _204_ (
		.din(new_net_107),
		.dout(new_net_198)
	);

	inv _205_ (
		.din(new_net_121),
		.dout(new_net_192)
	);

	and_bi _206_ (
		.a(new_net_16),
		.b(new_net_108),
		.c(_031_)
	);

	or_bb _207_ (
		.a(_031_),
		.b(new_net_98),
		.c(_032_)
	);

	or_bi _208_ (
		.a(new_net_109),
		.b(new_net_90),
		.c(_033_)
	);

	and_bi _209_ (
		.a(_033_),
		.b(new_net_86),
		.c(_034_)
	);

	or_bi _210_ (
		.a(new_net_79),
		.b(new_net_23),
		.c(_035_)
	);

	and_bi _211_ (
		.a(new_net_72),
		.b(new_net_102),
		.c(_036_)
	);

	and_ii _212_ (
		.a(_036_),
		.b(new_net_30),
		.c(_037_)
	);

	and_bi _213_ (
		.a(new_net_103),
		.b(new_net_60),
		.c(_038_)
	);

	or_bb _214_ (
		.a(_038_),
		.b(new_net_84),
		.c(_039_)
	);

	or_bb _215_ (
		.a(new_net_186),
		.b(new_net_13),
		.c(_040_)
	);

	or_bb _216_ (
		.a(new_net_99),
		.b(new_net_128),
		.c(new_net_0)
	);

	and_bi _217_ (
		.a(new_net_153),
		.b(new_net_104),
		.c(_041_)
	);

	or_bb _218_ (
		.a(_041_),
		.b(new_net_12),
		.c(_042_)
	);

	and_bi _219_ (
		.a(new_net_159),
		.b(new_net_105),
		.c(_043_)
	);

	and_ii _220_ (
		.a(_043_),
		.b(new_net_141),
		.c(_044_)
	);

	or_bi _221_ (
		.a(new_net_61),
		.b(new_net_5),
		.c(_045_)
	);

	and_bi _222_ (
		.a(new_net_94),
		.b(new_net_110),
		.c(_046_)
	);

	or_bb _223_ (
		.a(_046_),
		.b(new_net_2),
		.c(_047_)
	);

	and_bi _224_ (
		.a(new_net_70),
		.b(new_net_111),
		.c(_048_)
	);

	or_bb _225_ (
		.a(_048_),
		.b(new_net_131),
		.c(_049_)
	);

	or_ii _226_ (
		.a(new_net_187),
		.b(new_net_156),
		.c(_050_)
	);

	or_bb _227_ (
		.a(new_net_188),
		.b(new_net_87),
		.c(_051_)
	);

	or_bb _228_ (
		.a(new_net_189),
		.b(new_net_115),
		.c(_052_)
	);

	or_bi _229_ (
		.a(new_net_106),
		.b(new_net_96),
		.c(_053_)
	);

	and_bi _230_ (
		.a(_053_),
		.b(new_net_78),
		.c(_054_)
	);

	and_bi _231_ (
		.a(_052_),
		.b(new_net_190),
		.c(N421)
	);

	and_bi _232_ (
		.a(new_net_88),
		.b(new_net_101),
		.c(_055_)
	);

	or_bb _233_ (
		.a(_055_),
		.b(new_net_129),
		.c(new_net_196)
	);

	or_bi _234_ (
		.a(new_net_100),
		.b(new_net_62),
		.c(_056_)
	);

	and_bi _235_ (
		.a(new_net_6),
		.b(new_net_157),
		.c(_057_)
	);

	or_bb _236_ (
		.a(_057_),
		.b(new_net_14),
		.c(_058_)
	);

	and_bi _237_ (
		.a(_056_),
		.b(new_net_191),
		.c(_059_)
	);

	and_bi _238_ (
		.a(new_net_24),
		.b(_059_),
		.c(_060_)
	);

	or_bb _239_ (
		.a(_060_),
		.b(new_net_80),
		.c(N432)
	);

	inv _240_ (
		.din(new_net_46),
		.dout(new_net_194)
	);

	bfr new_net_200_bfr_before (
		.din(new_net_200),
		.dout(N430)
	);

	bfr new_net_201_bfr_before (
		.din(new_net_201),
		.dout(new_net_200)
	);

	spl2 new_net_0_v_fanout (
		.a(new_net_0),
		.b(new_net_201),
		.c(new_net_115)
	);

	bfr new_net_202_bfr_before (
		.din(new_net_202),
		.dout(new_net_129)
	);

	spl2 _035__v_fanout (
		.a(_035_),
		.b(new_net_128),
		.c(new_net_202)
	);

	spl2 _045__v_fanout (
		.a(_045_),
		.b(new_net_87),
		.c(new_net_88)
	);

	spl3L _040__v_fanout (
		.a(_040_),
		.b(new_net_101),
		.c(new_net_100),
		.d(new_net_99)
	);

	spl2 _047__v_fanout (
		.a(_047_),
		.b(new_net_156),
		.c(new_net_157)
	);

	bfr new_net_203_bfr_before (
		.din(new_net_203),
		.dout(new_net_62)
	);

	bfr new_net_204_bfr_before (
		.din(new_net_204),
		.dout(new_net_203)
	);

	spl2 _044__v_fanout (
		.a(_044_),
		.b(new_net_61),
		.c(new_net_204)
	);

	bfr new_net_205_bfr_before (
		.din(new_net_205),
		.dout(new_net_80)
	);

	bfr new_net_206_bfr_before (
		.din(new_net_206),
		.dout(new_net_205)
	);

	bfr new_net_207_bfr_before (
		.din(new_net_207),
		.dout(new_net_206)
	);

	bfr new_net_208_bfr_before (
		.din(new_net_208),
		.dout(new_net_207)
	);

	bfr new_net_209_bfr_before (
		.din(new_net_209),
		.dout(new_net_208)
	);

	spl2 _034__v_fanout (
		.a(_034_),
		.b(new_net_79),
		.c(new_net_209)
	);

	spl2 _042__v_fanout (
		.a(_042_),
		.b(new_net_5),
		.c(new_net_6)
	);

	bfr new_net_210_bfr_before (
		.din(new_net_210),
		.dout(new_net_24)
	);

	bfr new_net_211_bfr_before (
		.din(new_net_211),
		.dout(new_net_210)
	);

	bfr new_net_212_bfr_before (
		.din(new_net_212),
		.dout(new_net_211)
	);

	bfr new_net_213_bfr_before (
		.din(new_net_213),
		.dout(new_net_212)
	);

	spl2 _032__v_fanout (
		.a(_032_),
		.b(new_net_23),
		.c(new_net_213)
	);

	bfr new_net_214_bfr_before (
		.din(new_net_214),
		.dout(new_net_14)
	);

	spl2 _037__v_fanout (
		.a(_037_),
		.b(new_net_13),
		.c(new_net_214)
	);

	spl4L new_net_168_v_fanout (
		.a(new_net_168),
		.b(new_net_110),
		.c(new_net_111),
		.d(new_net_108),
		.e(new_net_109)
	);

	spl2 new_net_166_v_fanout (
		.a(new_net_166),
		.b(new_net_102),
		.c(new_net_106)
	);

	spl4L new_net_167_v_fanout (
		.a(new_net_167),
		.b(new_net_104),
		.c(new_net_103),
		.d(new_net_105),
		.e(new_net_107)
	);

	spl3L _030__v_fanout (
		.a(_030_),
		.b(new_net_167),
		.c(new_net_168),
		.d(new_net_166)
	);

	bfr new_net_215_bfr_before (
		.din(new_net_215),
		.dout(new_net_84)
	);

	bfr new_net_216_bfr_before (
		.din(new_net_216),
		.dout(new_net_215)
	);

	bfr new_net_217_bfr_before (
		.din(new_net_217),
		.dout(new_net_216)
	);

	bfr new_net_218_bfr_before (
		.din(new_net_218),
		.dout(new_net_217)
	);

	bfr new_net_219_bfr_before (
		.din(new_net_219),
		.dout(new_net_218)
	);

	bfr new_net_220_bfr_before (
		.din(new_net_220),
		.dout(new_net_219)
	);

	bfr new_net_221_bfr_before (
		.din(new_net_221),
		.dout(new_net_220)
	);

	spl2 _019__v_fanout (
		.a(_019_),
		.b(new_net_83),
		.c(new_net_221)
	);

	bfr new_net_222_bfr_before (
		.din(new_net_222),
		.dout(new_net_98)
	);

	bfr new_net_223_bfr_before (
		.din(new_net_223),
		.dout(new_net_222)
	);

	bfr new_net_224_bfr_before (
		.din(new_net_224),
		.dout(new_net_223)
	);

	bfr new_net_225_bfr_before (
		.din(new_net_225),
		.dout(new_net_224)
	);

	bfr new_net_226_bfr_before (
		.din(new_net_226),
		.dout(new_net_225)
	);

	bfr new_net_227_bfr_before (
		.din(new_net_227),
		.dout(new_net_226)
	);

	bfr new_net_228_bfr_before (
		.din(new_net_228),
		.dout(new_net_227)
	);

	bfr new_net_229_bfr_before (
		.din(new_net_229),
		.dout(new_net_228)
	);

	bfr new_net_230_bfr_before (
		.din(new_net_230),
		.dout(new_net_229)
	);

	spl2 _114__v_fanout (
		.a(_114_),
		.b(new_net_97),
		.c(new_net_230)
	);

	bfr new_net_231_bfr_before (
		.din(new_net_231),
		.dout(new_net_86)
	);

	bfr new_net_232_bfr_before (
		.din(new_net_232),
		.dout(new_net_231)
	);

	bfr new_net_233_bfr_before (
		.din(new_net_233),
		.dout(new_net_232)
	);

	bfr new_net_234_bfr_before (
		.din(new_net_234),
		.dout(new_net_233)
	);

	bfr new_net_235_bfr_before (
		.din(new_net_235),
		.dout(new_net_234)
	);

	bfr new_net_236_bfr_before (
		.din(new_net_236),
		.dout(new_net_235)
	);

	bfr new_net_237_bfr_before (
		.din(new_net_237),
		.dout(new_net_236)
	);

	bfr new_net_238_bfr_before (
		.din(new_net_238),
		.dout(new_net_237)
	);

	bfr new_net_239_bfr_before (
		.din(new_net_239),
		.dout(new_net_238)
	);

	spl2 _003__v_fanout (
		.a(_003_),
		.b(new_net_85),
		.c(new_net_239)
	);

	bfr new_net_240_bfr_before (
		.din(new_net_240),
		.dout(new_net_141)
	);

	bfr new_net_241_bfr_before (
		.din(new_net_241),
		.dout(new_net_240)
	);

	bfr new_net_242_bfr_before (
		.din(new_net_242),
		.dout(new_net_241)
	);

	bfr new_net_243_bfr_before (
		.din(new_net_243),
		.dout(new_net_242)
	);

	bfr new_net_244_bfr_before (
		.din(new_net_244),
		.dout(new_net_243)
	);

	bfr new_net_245_bfr_before (
		.din(new_net_245),
		.dout(new_net_244)
	);

	bfr new_net_246_bfr_before (
		.din(new_net_246),
		.dout(new_net_245)
	);

	bfr new_net_247_bfr_before (
		.din(new_net_247),
		.dout(new_net_246)
	);

	bfr new_net_248_bfr_before (
		.din(new_net_248),
		.dout(new_net_247)
	);

	spl2 _015__v_fanout (
		.a(_015_),
		.b(new_net_140),
		.c(new_net_248)
	);

	bfr new_net_249_bfr_before (
		.din(new_net_249),
		.dout(new_net_2)
	);

	bfr new_net_250_bfr_before (
		.din(new_net_250),
		.dout(new_net_249)
	);

	bfr new_net_251_bfr_before (
		.din(new_net_251),
		.dout(new_net_250)
	);

	bfr new_net_252_bfr_before (
		.din(new_net_252),
		.dout(new_net_251)
	);

	bfr new_net_253_bfr_before (
		.din(new_net_253),
		.dout(new_net_252)
	);

	bfr new_net_254_bfr_before (
		.din(new_net_254),
		.dout(new_net_253)
	);

	bfr new_net_255_bfr_before (
		.din(new_net_255),
		.dout(new_net_254)
	);

	bfr new_net_256_bfr_before (
		.din(new_net_256),
		.dout(new_net_255)
	);

	bfr new_net_257_bfr_before (
		.din(new_net_257),
		.dout(new_net_256)
	);

	spl2 _000__v_fanout (
		.a(_000_),
		.b(new_net_1),
		.c(new_net_257)
	);

	bfr new_net_258_bfr_before (
		.din(new_net_258),
		.dout(new_net_60)
	);

	bfr new_net_259_bfr_before (
		.din(new_net_259),
		.dout(new_net_258)
	);

	bfr new_net_260_bfr_before (
		.din(new_net_260),
		.dout(new_net_259)
	);

	bfr new_net_261_bfr_before (
		.din(new_net_261),
		.dout(new_net_260)
	);

	bfr new_net_262_bfr_before (
		.din(new_net_262),
		.dout(new_net_261)
	);

	bfr new_net_263_bfr_before (
		.din(new_net_263),
		.dout(new_net_262)
	);

	bfr new_net_264_bfr_before (
		.din(new_net_264),
		.dout(new_net_263)
	);

	bfr new_net_265_bfr_before (
		.din(new_net_265),
		.dout(new_net_264)
	);

	spl2 _018__v_fanout (
		.a(_018_),
		.b(new_net_59),
		.c(new_net_265)
	);

	bfr new_net_266_bfr_before (
		.din(new_net_266),
		.dout(new_net_131)
	);

	bfr new_net_267_bfr_before (
		.din(new_net_267),
		.dout(new_net_266)
	);

	bfr new_net_268_bfr_before (
		.din(new_net_268),
		.dout(new_net_267)
	);

	bfr new_net_269_bfr_before (
		.din(new_net_269),
		.dout(new_net_268)
	);

	bfr new_net_270_bfr_before (
		.din(new_net_270),
		.dout(new_net_269)
	);

	bfr new_net_271_bfr_before (
		.din(new_net_271),
		.dout(new_net_270)
	);

	bfr new_net_272_bfr_before (
		.din(new_net_272),
		.dout(new_net_271)
	);

	bfr new_net_273_bfr_before (
		.din(new_net_273),
		.dout(new_net_272)
	);

	bfr new_net_274_bfr_before (
		.din(new_net_274),
		.dout(new_net_273)
	);

	spl2 _025__v_fanout (
		.a(_025_),
		.b(new_net_130),
		.c(new_net_274)
	);

	bfr new_net_275_bfr_before (
		.din(new_net_275),
		.dout(new_net_78)
	);

	bfr new_net_276_bfr_before (
		.din(new_net_276),
		.dout(new_net_275)
	);

	bfr new_net_277_bfr_before (
		.din(new_net_277),
		.dout(new_net_276)
	);

	bfr new_net_278_bfr_before (
		.din(new_net_278),
		.dout(new_net_277)
	);

	bfr new_net_279_bfr_before (
		.din(new_net_279),
		.dout(new_net_278)
	);

	bfr new_net_280_bfr_before (
		.din(new_net_280),
		.dout(new_net_279)
	);

	bfr new_net_281_bfr_before (
		.din(new_net_281),
		.dout(new_net_280)
	);

	bfr new_net_282_bfr_before (
		.din(new_net_282),
		.dout(new_net_281)
	);

	bfr new_net_283_bfr_before (
		.din(new_net_283),
		.dout(new_net_282)
	);

	spl2 _008__v_fanout (
		.a(_008_),
		.b(new_net_77),
		.c(new_net_283)
	);

	bfr new_net_284_bfr_before (
		.din(new_net_284),
		.dout(new_net_12)
	);

	bfr new_net_285_bfr_before (
		.din(new_net_285),
		.dout(new_net_284)
	);

	bfr new_net_286_bfr_before (
		.din(new_net_286),
		.dout(new_net_285)
	);

	bfr new_net_287_bfr_before (
		.din(new_net_287),
		.dout(new_net_286)
	);

	bfr new_net_288_bfr_before (
		.din(new_net_288),
		.dout(new_net_287)
	);

	bfr new_net_289_bfr_before (
		.din(new_net_289),
		.dout(new_net_288)
	);

	bfr new_net_290_bfr_before (
		.din(new_net_290),
		.dout(new_net_289)
	);

	bfr new_net_291_bfr_before (
		.din(new_net_291),
		.dout(new_net_290)
	);

	bfr new_net_292_bfr_before (
		.din(new_net_292),
		.dout(new_net_291)
	);

	spl2 _011__v_fanout (
		.a(_011_),
		.b(new_net_11),
		.c(new_net_292)
	);

	bfr new_net_293_bfr_before (
		.din(new_net_293),
		.dout(new_net_30)
	);

	bfr new_net_294_bfr_before (
		.din(new_net_294),
		.dout(new_net_293)
	);

	bfr new_net_295_bfr_before (
		.din(new_net_295),
		.dout(new_net_294)
	);

	bfr new_net_296_bfr_before (
		.din(new_net_296),
		.dout(new_net_295)
	);

	bfr new_net_297_bfr_before (
		.din(new_net_297),
		.dout(new_net_296)
	);

	bfr new_net_298_bfr_before (
		.din(new_net_298),
		.dout(new_net_297)
	);

	bfr new_net_299_bfr_before (
		.din(new_net_299),
		.dout(new_net_298)
	);

	bfr new_net_300_bfr_before (
		.din(new_net_300),
		.dout(new_net_299)
	);

	bfr new_net_301_bfr_before (
		.din(new_net_301),
		.dout(new_net_300)
	);

	spl2 _022__v_fanout (
		.a(_022_),
		.b(new_net_29),
		.c(new_net_301)
	);

	spl4L new_net_164_v_fanout (
		.a(new_net_164),
		.b(new_net_41),
		.c(new_net_40),
		.d(new_net_39),
		.e(new_net_42)
	);

	spl4L new_net_165_v_fanout (
		.a(new_net_165),
		.b(new_net_44),
		.c(new_net_46),
		.d(new_net_43),
		.e(new_net_45)
	);

	spl2 new_net_163_v_fanout (
		.a(new_net_163),
		.b(new_net_37),
		.c(new_net_38)
	);

	spl3L _112__v_fanout (
		.a(_112_),
		.b(new_net_164),
		.c(new_net_165),
		.d(new_net_163)
	);

	bfr new_net_302_bfr_before (
		.din(new_net_302),
		.dout(new_net_66)
	);

	bfr new_net_303_bfr_before (
		.din(new_net_303),
		.dout(new_net_302)
	);

	bfr new_net_304_bfr_before (
		.din(new_net_304),
		.dout(new_net_303)
	);

	bfr new_net_305_bfr_before (
		.din(new_net_305),
		.dout(new_net_304)
	);

	bfr new_net_306_bfr_before (
		.din(new_net_306),
		.dout(new_net_305)
	);

	bfr new_net_307_bfr_before (
		.din(new_net_307),
		.dout(new_net_306)
	);

	bfr new_net_308_bfr_before (
		.din(new_net_308),
		.dout(new_net_307)
	);

	bfr new_net_309_bfr_before (
		.din(new_net_309),
		.dout(new_net_308)
	);

	spl2 _081__v_fanout (
		.a(_081_),
		.b(new_net_65),
		.c(new_net_309)
	);

	bfr new_net_310_bfr_before (
		.din(new_net_310),
		.dout(new_net_155)
	);

	bfr new_net_311_bfr_before (
		.din(new_net_311),
		.dout(new_net_310)
	);

	bfr new_net_312_bfr_before (
		.din(new_net_312),
		.dout(new_net_311)
	);

	bfr new_net_313_bfr_before (
		.din(new_net_313),
		.dout(new_net_312)
	);

	bfr new_net_314_bfr_before (
		.din(new_net_314),
		.dout(new_net_313)
	);

	bfr new_net_315_bfr_before (
		.din(new_net_315),
		.dout(new_net_314)
	);

	bfr new_net_316_bfr_before (
		.din(new_net_316),
		.dout(new_net_315)
	);

	bfr new_net_317_bfr_before (
		.din(new_net_317),
		.dout(new_net_316)
	);

	spl2 _089__v_fanout (
		.a(_089_),
		.b(new_net_154),
		.c(new_net_317)
	);

	bfr new_net_318_bfr_before (
		.din(new_net_318),
		.dout(new_net_137)
	);

	bfr new_net_319_bfr_before (
		.din(new_net_319),
		.dout(new_net_318)
	);

	bfr new_net_320_bfr_before (
		.din(new_net_320),
		.dout(new_net_319)
	);

	bfr new_net_321_bfr_before (
		.din(new_net_321),
		.dout(new_net_320)
	);

	bfr new_net_322_bfr_before (
		.din(new_net_322),
		.dout(new_net_321)
	);

	bfr new_net_323_bfr_before (
		.din(new_net_323),
		.dout(new_net_322)
	);

	bfr new_net_324_bfr_before (
		.din(new_net_324),
		.dout(new_net_323)
	);

	bfr new_net_325_bfr_before (
		.din(new_net_325),
		.dout(new_net_324)
	);

	spl2 _104__v_fanout (
		.a(_104_),
		.b(new_net_136),
		.c(new_net_325)
	);

	bfr new_net_326_bfr_before (
		.din(new_net_326),
		.dout(new_net_34)
	);

	bfr new_net_327_bfr_before (
		.din(new_net_327),
		.dout(new_net_326)
	);

	bfr new_net_328_bfr_before (
		.din(new_net_328),
		.dout(new_net_327)
	);

	bfr new_net_329_bfr_before (
		.din(new_net_329),
		.dout(new_net_328)
	);

	bfr new_net_330_bfr_before (
		.din(new_net_330),
		.dout(new_net_329)
	);

	bfr new_net_331_bfr_before (
		.din(new_net_331),
		.dout(new_net_330)
	);

	bfr new_net_332_bfr_before (
		.din(new_net_332),
		.dout(new_net_331)
	);

	bfr new_net_333_bfr_before (
		.din(new_net_333),
		.dout(new_net_332)
	);

	spl2 _101__v_fanout (
		.a(_101_),
		.b(new_net_33),
		.c(new_net_333)
	);

	bfr new_net_334_bfr_before (
		.din(new_net_334),
		.dout(new_net_20)
	);

	bfr new_net_335_bfr_before (
		.din(new_net_335),
		.dout(new_net_334)
	);

	bfr new_net_336_bfr_before (
		.din(new_net_336),
		.dout(new_net_335)
	);

	bfr new_net_337_bfr_before (
		.din(new_net_337),
		.dout(new_net_336)
	);

	bfr new_net_338_bfr_before (
		.din(new_net_338),
		.dout(new_net_337)
	);

	bfr new_net_339_bfr_before (
		.din(new_net_339),
		.dout(new_net_338)
	);

	bfr new_net_340_bfr_before (
		.din(new_net_340),
		.dout(new_net_339)
	);

	bfr new_net_341_bfr_before (
		.din(new_net_341),
		.dout(new_net_340)
	);

	spl2 _079__v_fanout (
		.a(_079_),
		.b(new_net_19),
		.c(new_net_341)
	);

	bfr new_net_342_bfr_before (
		.din(new_net_342),
		.dout(new_net_4)
	);

	bfr new_net_343_bfr_before (
		.din(new_net_343),
		.dout(new_net_342)
	);

	bfr new_net_344_bfr_before (
		.din(new_net_344),
		.dout(new_net_343)
	);

	bfr new_net_345_bfr_before (
		.din(new_net_345),
		.dout(new_net_344)
	);

	bfr new_net_346_bfr_before (
		.din(new_net_346),
		.dout(new_net_345)
	);

	bfr new_net_347_bfr_before (
		.din(new_net_347),
		.dout(new_net_346)
	);

	bfr new_net_348_bfr_before (
		.din(new_net_348),
		.dout(new_net_347)
	);

	bfr new_net_349_bfr_before (
		.din(new_net_349),
		.dout(new_net_348)
	);

	spl2 _084__v_fanout (
		.a(_084_),
		.b(new_net_3),
		.c(new_net_349)
	);

	bfr new_net_350_bfr_before (
		.din(new_net_350),
		.dout(new_net_68)
	);

	bfr new_net_351_bfr_before (
		.din(new_net_351),
		.dout(new_net_350)
	);

	bfr new_net_352_bfr_before (
		.din(new_net_352),
		.dout(new_net_351)
	);

	bfr new_net_353_bfr_before (
		.din(new_net_353),
		.dout(new_net_352)
	);

	bfr new_net_354_bfr_before (
		.din(new_net_354),
		.dout(new_net_353)
	);

	bfr new_net_355_bfr_before (
		.din(new_net_355),
		.dout(new_net_354)
	);

	bfr new_net_356_bfr_before (
		.din(new_net_356),
		.dout(new_net_355)
	);

	bfr new_net_357_bfr_before (
		.din(new_net_357),
		.dout(new_net_356)
	);

	spl2 _097__v_fanout (
		.a(_097_),
		.b(new_net_67),
		.c(new_net_357)
	);

	bfr new_net_358_bfr_before (
		.din(new_net_358),
		.dout(new_net_151)
	);

	bfr new_net_359_bfr_before (
		.din(new_net_359),
		.dout(new_net_358)
	);

	bfr new_net_360_bfr_before (
		.din(new_net_360),
		.dout(new_net_359)
	);

	bfr new_net_361_bfr_before (
		.din(new_net_361),
		.dout(new_net_360)
	);

	bfr new_net_362_bfr_before (
		.din(new_net_362),
		.dout(new_net_361)
	);

	bfr new_net_363_bfr_before (
		.din(new_net_363),
		.dout(new_net_362)
	);

	bfr new_net_364_bfr_before (
		.din(new_net_364),
		.dout(new_net_363)
	);

	bfr new_net_365_bfr_before (
		.din(new_net_365),
		.dout(new_net_364)
	);

	spl2 _094__v_fanout (
		.a(_094_),
		.b(new_net_150),
		.c(new_net_365)
	);

	bfr new_net_366_bfr_before (
		.din(new_net_366),
		.dout(new_net_52)
	);

	bfr new_net_367_bfr_before (
		.din(new_net_367),
		.dout(new_net_366)
	);

	bfr new_net_368_bfr_before (
		.din(new_net_368),
		.dout(new_net_367)
	);

	bfr new_net_369_bfr_before (
		.din(new_net_369),
		.dout(new_net_368)
	);

	bfr new_net_370_bfr_before (
		.din(new_net_370),
		.dout(new_net_369)
	);

	bfr new_net_371_bfr_before (
		.din(new_net_371),
		.dout(new_net_370)
	);

	bfr new_net_372_bfr_before (
		.din(new_net_372),
		.dout(new_net_371)
	);

	bfr new_net_373_bfr_before (
		.din(new_net_373),
		.dout(new_net_372)
	);

	spl2 _107__v_fanout (
		.a(_107_),
		.b(new_net_51),
		.c(new_net_373)
	);

	spl4L new_net_161_v_fanout (
		.a(new_net_161),
		.b(new_net_123),
		.c(new_net_121),
		.d(new_net_120),
		.e(new_net_122)
	);

	spl4L new_net_162_v_fanout (
		.a(new_net_162),
		.b(new_net_125),
		.c(new_net_127),
		.d(new_net_124),
		.e(new_net_126)
	);

	spl2 new_net_160_v_fanout (
		.a(new_net_160),
		.b(new_net_118),
		.c(new_net_119)
	);

	spl3L _077__v_fanout (
		.a(_077_),
		.b(new_net_161),
		.c(new_net_162),
		.d(new_net_160)
	);

	bfr new_net_374_bfr_before (
		.din(new_net_374),
		.dout(new_net_117)
	);

	bfr new_net_375_bfr_before (
		.din(new_net_375),
		.dout(new_net_374)
	);

	bfr new_net_376_bfr_before (
		.din(new_net_376),
		.dout(new_net_375)
	);

	bfr new_net_377_bfr_before (
		.din(new_net_377),
		.dout(new_net_376)
	);

	bfr new_net_378_bfr_before (
		.din(new_net_378),
		.dout(new_net_377)
	);

	bfr new_net_379_bfr_before (
		.din(new_net_379),
		.dout(new_net_378)
	);

	bfr new_net_380_bfr_before (
		.din(new_net_380),
		.dout(new_net_379)
	);

	spl2 _061__v_fanout (
		.a(_061_),
		.b(new_net_116),
		.c(new_net_380)
	);

	bfr new_net_381_bfr_before (
		.din(new_net_381),
		.dout(new_net_10)
	);

	bfr new_net_382_bfr_before (
		.din(new_net_382),
		.dout(new_net_381)
	);

	bfr new_net_383_bfr_before (
		.din(new_net_383),
		.dout(new_net_382)
	);

	bfr new_net_384_bfr_before (
		.din(new_net_384),
		.dout(new_net_383)
	);

	bfr new_net_385_bfr_before (
		.din(new_net_385),
		.dout(new_net_384)
	);

	bfr new_net_386_bfr_before (
		.din(new_net_386),
		.dout(new_net_385)
	);

	bfr new_net_387_bfr_before (
		.din(new_net_387),
		.dout(new_net_386)
	);

	spl2 _069__v_fanout (
		.a(_069_),
		.b(new_net_9),
		.c(new_net_387)
	);

	bfr new_net_388_bfr_after (
		.din(N112),
		.dout(new_net_388)
	);

	bfr new_net_389_bfr_after (
		.din(new_net_388),
		.dout(new_net_389)
	);

	bfr new_net_390_bfr_after (
		.din(new_net_389),
		.dout(new_net_390)
	);

	bfr new_net_391_bfr_after (
		.din(new_net_390),
		.dout(new_net_391)
	);

	bfr new_net_392_bfr_after (
		.din(new_net_391),
		.dout(new_net_392)
	);

	bfr new_net_393_bfr_after (
		.din(new_net_392),
		.dout(new_net_393)
	);

	bfr new_net_394_bfr_after (
		.din(new_net_393),
		.dout(new_net_394)
	);

	bfr new_net_395_bfr_after (
		.din(new_net_394),
		.dout(new_net_395)
	);

	bfr new_net_396_bfr_after (
		.din(new_net_395),
		.dout(new_net_396)
	);

	bfr new_net_397_bfr_after (
		.din(new_net_396),
		.dout(new_net_397)
	);

	bfr new_net_398_bfr_after (
		.din(new_net_397),
		.dout(new_net_398)
	);

	bfr new_net_399_bfr_before (
		.din(new_net_399),
		.dout(new_net_48)
	);

	bfr new_net_400_bfr_before (
		.din(new_net_400),
		.dout(new_net_399)
	);

	bfr new_net_401_bfr_before (
		.din(new_net_401),
		.dout(new_net_400)
	);

	bfr new_net_402_bfr_before (
		.din(new_net_402),
		.dout(new_net_401)
	);

	bfr new_net_403_bfr_before (
		.din(new_net_403),
		.dout(new_net_402)
	);

	bfr new_net_404_bfr_before (
		.din(new_net_404),
		.dout(new_net_403)
	);

	bfr new_net_405_bfr_before (
		.din(new_net_405),
		.dout(new_net_404)
	);

	spl2 N112_v_fanout (
		.a(new_net_398),
		.b(new_net_47),
		.c(new_net_405)
	);

	bfr new_net_406_bfr_before (
		.din(new_net_406),
		.dout(new_net_50)
	);

	bfr new_net_407_bfr_before (
		.din(new_net_407),
		.dout(new_net_406)
	);

	bfr new_net_408_bfr_before (
		.din(new_net_408),
		.dout(new_net_407)
	);

	bfr new_net_409_bfr_before (
		.din(new_net_409),
		.dout(new_net_408)
	);

	bfr new_net_410_bfr_before (
		.din(new_net_410),
		.dout(new_net_409)
	);

	bfr new_net_411_bfr_before (
		.din(new_net_411),
		.dout(new_net_410)
	);

	bfr new_net_412_bfr_before (
		.din(new_net_412),
		.dout(new_net_411)
	);

	bfr new_net_413_bfr_before (
		.din(new_net_413),
		.dout(new_net_412)
	);

	spl2 N50_v_fanout (
		.a(N50),
		.b(new_net_49),
		.c(new_net_413)
	);

	bfr new_net_414_bfr_after (
		.din(N105),
		.dout(new_net_414)
	);

	bfr new_net_415_bfr_after (
		.din(new_net_414),
		.dout(new_net_415)
	);

	bfr new_net_416_bfr_after (
		.din(new_net_415),
		.dout(new_net_416)
	);

	bfr new_net_417_bfr_after (
		.din(new_net_416),
		.dout(new_net_417)
	);

	bfr new_net_418_bfr_after (
		.din(new_net_417),
		.dout(new_net_418)
	);

	bfr new_net_419_bfr_after (
		.din(new_net_418),
		.dout(new_net_419)
	);

	bfr new_net_420_bfr_after (
		.din(new_net_419),
		.dout(new_net_420)
	);

	bfr new_net_421_bfr_after (
		.din(new_net_420),
		.dout(new_net_421)
	);

	bfr new_net_422_bfr_after (
		.din(new_net_421),
		.dout(new_net_422)
	);

	bfr new_net_423_bfr_after (
		.din(new_net_422),
		.dout(new_net_423)
	);

	bfr new_net_424_bfr_after (
		.din(new_net_423),
		.dout(new_net_424)
	);

	bfr new_net_425_bfr_after (
		.din(new_net_424),
		.dout(new_net_425)
	);

	bfr new_net_426_bfr_after (
		.din(new_net_425),
		.dout(new_net_426)
	);

	bfr new_net_427_bfr_after (
		.din(new_net_426),
		.dout(new_net_427)
	);

	bfr new_net_428_bfr_after (
		.din(new_net_427),
		.dout(new_net_428)
	);

	bfr new_net_429_bfr_after (
		.din(new_net_428),
		.dout(new_net_429)
	);

	bfr new_net_430_bfr_after (
		.din(new_net_429),
		.dout(new_net_430)
	);

	bfr new_net_431_bfr_after (
		.din(new_net_430),
		.dout(new_net_431)
	);

	bfr new_net_432_bfr_after (
		.din(new_net_431),
		.dout(new_net_432)
	);

	bfr new_net_433_bfr_after (
		.din(new_net_432),
		.dout(new_net_433)
	);

	bfr new_net_434_bfr_after (
		.din(new_net_433),
		.dout(new_net_434)
	);

	bfr new_net_435_bfr_before (
		.din(new_net_435),
		.dout(new_net_94)
	);

	bfr new_net_436_bfr_before (
		.din(new_net_436),
		.dout(new_net_435)
	);

	bfr new_net_437_bfr_before (
		.din(new_net_437),
		.dout(new_net_436)
	);

	bfr new_net_438_bfr_before (
		.din(new_net_438),
		.dout(new_net_437)
	);

	bfr new_net_439_bfr_before (
		.din(new_net_439),
		.dout(new_net_438)
	);

	bfr new_net_440_bfr_before (
		.din(new_net_440),
		.dout(new_net_439)
	);

	bfr new_net_441_bfr_before (
		.din(new_net_441),
		.dout(new_net_440)
	);

	bfr new_net_442_bfr_before (
		.din(new_net_442),
		.dout(new_net_441)
	);

	spl2 N105_v_fanout (
		.a(new_net_434),
		.b(new_net_93),
		.c(new_net_442)
	);

	bfr new_net_443_bfr_after (
		.din(N86),
		.dout(new_net_443)
	);

	bfr new_net_444_bfr_after (
		.din(new_net_443),
		.dout(new_net_444)
	);

	bfr new_net_445_bfr_after (
		.din(new_net_444),
		.dout(new_net_445)
	);

	bfr new_net_446_bfr_after (
		.din(new_net_445),
		.dout(new_net_446)
	);

	bfr new_net_447_bfr_after (
		.din(new_net_446),
		.dout(new_net_447)
	);

	bfr new_net_448_bfr_after (
		.din(new_net_447),
		.dout(new_net_448)
	);

	bfr new_net_449_bfr_after (
		.din(new_net_448),
		.dout(new_net_449)
	);

	bfr new_net_450_bfr_after (
		.din(new_net_449),
		.dout(new_net_450)
	);

	bfr new_net_451_bfr_after (
		.din(new_net_450),
		.dout(new_net_451)
	);

	bfr new_net_452_bfr_after (
		.din(new_net_451),
		.dout(new_net_452)
	);

	bfr new_net_453_bfr_after (
		.din(new_net_452),
		.dout(new_net_453)
	);

	bfr new_net_454_bfr_before (
		.din(new_net_454),
		.dout(new_net_82)
	);

	bfr new_net_455_bfr_before (
		.din(new_net_455),
		.dout(new_net_454)
	);

	bfr new_net_456_bfr_before (
		.din(new_net_456),
		.dout(new_net_455)
	);

	bfr new_net_457_bfr_before (
		.din(new_net_457),
		.dout(new_net_456)
	);

	bfr new_net_458_bfr_before (
		.din(new_net_458),
		.dout(new_net_457)
	);

	bfr new_net_459_bfr_before (
		.din(new_net_459),
		.dout(new_net_458)
	);

	bfr new_net_460_bfr_before (
		.din(new_net_460),
		.dout(new_net_459)
	);

	spl2 N86_v_fanout (
		.a(new_net_453),
		.b(new_net_81),
		.c(new_net_460)
	);

	bfr new_net_461_bfr_after (
		.din(N21),
		.dout(new_net_461)
	);

	bfr new_net_462_bfr_after (
		.din(new_net_461),
		.dout(new_net_462)
	);

	bfr new_net_463_bfr_after (
		.din(new_net_462),
		.dout(new_net_463)
	);

	bfr new_net_464_bfr_after (
		.din(new_net_463),
		.dout(new_net_464)
	);

	bfr new_net_465_bfr_after (
		.din(new_net_464),
		.dout(new_net_465)
	);

	bfr new_net_466_bfr_after (
		.din(new_net_465),
		.dout(new_net_466)
	);

	bfr new_net_467_bfr_after (
		.din(new_net_466),
		.dout(new_net_467)
	);

	bfr new_net_468_bfr_after (
		.din(new_net_467),
		.dout(new_net_468)
	);

	bfr new_net_469_bfr_after (
		.din(new_net_468),
		.dout(new_net_469)
	);

	bfr new_net_470_bfr_after (
		.din(new_net_469),
		.dout(new_net_470)
	);

	bfr new_net_471_bfr_after (
		.din(new_net_470),
		.dout(new_net_471)
	);

	bfr new_net_472_bfr_before (
		.din(new_net_472),
		.dout(new_net_8)
	);

	bfr new_net_473_bfr_before (
		.din(new_net_473),
		.dout(new_net_472)
	);

	bfr new_net_474_bfr_before (
		.din(new_net_474),
		.dout(new_net_473)
	);

	bfr new_net_475_bfr_before (
		.din(new_net_475),
		.dout(new_net_474)
	);

	bfr new_net_476_bfr_before (
		.din(new_net_476),
		.dout(new_net_475)
	);

	bfr new_net_477_bfr_before (
		.din(new_net_477),
		.dout(new_net_476)
	);

	bfr new_net_478_bfr_before (
		.din(new_net_478),
		.dout(new_net_477)
	);

	spl2 N21_v_fanout (
		.a(new_net_471),
		.b(new_net_7),
		.c(new_net_478)
	);

	bfr new_net_479_bfr_after (
		.din(N47),
		.dout(new_net_479)
	);

	bfr new_net_480_bfr_after (
		.din(new_net_479),
		.dout(new_net_480)
	);

	bfr new_net_481_bfr_after (
		.din(new_net_480),
		.dout(new_net_481)
	);

	bfr new_net_482_bfr_after (
		.din(new_net_481),
		.dout(new_net_482)
	);

	bfr new_net_483_bfr_after (
		.din(new_net_482),
		.dout(new_net_483)
	);

	bfr new_net_484_bfr_after (
		.din(new_net_483),
		.dout(new_net_484)
	);

	bfr new_net_485_bfr_after (
		.din(new_net_484),
		.dout(new_net_485)
	);

	bfr new_net_486_bfr_after (
		.din(new_net_485),
		.dout(new_net_486)
	);

	bfr new_net_487_bfr_after (
		.din(new_net_486),
		.dout(new_net_487)
	);

	bfr new_net_488_bfr_after (
		.din(new_net_487),
		.dout(new_net_488)
	);

	bfr new_net_489_bfr_after (
		.din(new_net_488),
		.dout(new_net_489)
	);

	bfr new_net_490_bfr_before (
		.din(new_net_490),
		.dout(new_net_22)
	);

	bfr new_net_491_bfr_before (
		.din(new_net_491),
		.dout(new_net_490)
	);

	bfr new_net_492_bfr_before (
		.din(new_net_492),
		.dout(new_net_491)
	);

	bfr new_net_493_bfr_before (
		.din(new_net_493),
		.dout(new_net_492)
	);

	bfr new_net_494_bfr_before (
		.din(new_net_494),
		.dout(new_net_493)
	);

	bfr new_net_495_bfr_before (
		.din(new_net_495),
		.dout(new_net_494)
	);

	bfr new_net_496_bfr_before (
		.din(new_net_496),
		.dout(new_net_495)
	);

	spl2 N47_v_fanout (
		.a(new_net_489),
		.b(new_net_21),
		.c(new_net_496)
	);

	bfr new_net_497_bfr_after (
		.din(N60),
		.dout(new_net_497)
	);

	bfr new_net_498_bfr_after (
		.din(new_net_497),
		.dout(new_net_498)
	);

	bfr new_net_499_bfr_after (
		.din(new_net_498),
		.dout(new_net_499)
	);

	bfr new_net_500_bfr_after (
		.din(new_net_499),
		.dout(new_net_500)
	);

	bfr new_net_501_bfr_after (
		.din(new_net_500),
		.dout(new_net_501)
	);

	bfr new_net_502_bfr_after (
		.din(new_net_501),
		.dout(new_net_502)
	);

	bfr new_net_503_bfr_after (
		.din(new_net_502),
		.dout(new_net_503)
	);

	bfr new_net_504_bfr_after (
		.din(new_net_503),
		.dout(new_net_504)
	);

	bfr new_net_505_bfr_after (
		.din(new_net_504),
		.dout(new_net_505)
	);

	bfr new_net_506_bfr_after (
		.din(new_net_505),
		.dout(new_net_506)
	);

	bfr new_net_507_bfr_after (
		.din(new_net_506),
		.dout(new_net_507)
	);

	bfr new_net_508_bfr_before (
		.din(new_net_508),
		.dout(new_net_145)
	);

	bfr new_net_509_bfr_before (
		.din(new_net_509),
		.dout(new_net_508)
	);

	bfr new_net_510_bfr_before (
		.din(new_net_510),
		.dout(new_net_509)
	);

	bfr new_net_511_bfr_before (
		.din(new_net_511),
		.dout(new_net_510)
	);

	bfr new_net_512_bfr_before (
		.din(new_net_512),
		.dout(new_net_511)
	);

	bfr new_net_513_bfr_before (
		.din(new_net_513),
		.dout(new_net_512)
	);

	bfr new_net_514_bfr_before (
		.din(new_net_514),
		.dout(new_net_513)
	);

	spl2 N60_v_fanout (
		.a(new_net_507),
		.b(new_net_144),
		.c(new_net_514)
	);

	bfr new_net_515_bfr_before (
		.din(new_net_515),
		.dout(new_net_147)
	);

	bfr new_net_516_bfr_before (
		.din(new_net_516),
		.dout(new_net_515)
	);

	bfr new_net_517_bfr_before (
		.din(new_net_517),
		.dout(new_net_516)
	);

	bfr new_net_518_bfr_before (
		.din(new_net_518),
		.dout(new_net_517)
	);

	bfr new_net_519_bfr_before (
		.din(new_net_519),
		.dout(new_net_518)
	);

	bfr new_net_520_bfr_before (
		.din(new_net_520),
		.dout(new_net_519)
	);

	bfr new_net_521_bfr_before (
		.din(new_net_521),
		.dout(new_net_520)
	);

	bfr new_net_522_bfr_before (
		.din(new_net_522),
		.dout(new_net_521)
	);

	bfr new_net_523_bfr_before (
		.din(new_net_523),
		.dout(new_net_522)
	);

	spl2 N4_v_fanout (
		.a(N4),
		.b(new_net_146),
		.c(new_net_523)
	);

	bfr new_net_524_bfr_before (
		.din(new_net_524),
		.dout(new_net_18)
	);

	bfr new_net_525_bfr_before (
		.din(new_net_525),
		.dout(new_net_524)
	);

	bfr new_net_526_bfr_before (
		.din(new_net_526),
		.dout(new_net_525)
	);

	bfr new_net_527_bfr_before (
		.din(new_net_527),
		.dout(new_net_526)
	);

	bfr new_net_528_bfr_before (
		.din(new_net_528),
		.dout(new_net_527)
	);

	bfr new_net_529_bfr_before (
		.din(new_net_529),
		.dout(new_net_528)
	);

	bfr new_net_530_bfr_before (
		.din(new_net_530),
		.dout(new_net_529)
	);

	bfr new_net_531_bfr_before (
		.din(new_net_531),
		.dout(new_net_530)
	);

	spl2 N11_v_fanout (
		.a(N11),
		.b(new_net_17),
		.c(new_net_531)
	);

	bfr new_net_532_bfr_before (
		.din(new_net_532),
		.dout(new_net_28)
	);

	bfr new_net_533_bfr_before (
		.din(new_net_533),
		.dout(new_net_532)
	);

	bfr new_net_534_bfr_before (
		.din(new_net_534),
		.dout(new_net_533)
	);

	bfr new_net_535_bfr_before (
		.din(new_net_535),
		.dout(new_net_534)
	);

	bfr new_net_536_bfr_before (
		.din(new_net_536),
		.dout(new_net_535)
	);

	bfr new_net_537_bfr_before (
		.din(new_net_537),
		.dout(new_net_536)
	);

	bfr new_net_538_bfr_before (
		.din(new_net_538),
		.dout(new_net_537)
	);

	bfr new_net_539_bfr_before (
		.din(new_net_539),
		.dout(new_net_538)
	);

	bfr new_net_540_bfr_before (
		.din(new_net_540),
		.dout(new_net_539)
	);

	spl2 N95_v_fanout (
		.a(N95),
		.b(new_net_27),
		.c(new_net_540)
	);

	bfr new_net_541_bfr_before (
		.din(new_net_541),
		.dout(new_net_149)
	);

	bfr new_net_542_bfr_before (
		.din(new_net_542),
		.dout(new_net_541)
	);

	bfr new_net_543_bfr_before (
		.din(new_net_543),
		.dout(new_net_542)
	);

	bfr new_net_544_bfr_before (
		.din(new_net_544),
		.dout(new_net_543)
	);

	bfr new_net_545_bfr_before (
		.din(new_net_545),
		.dout(new_net_544)
	);

	bfr new_net_546_bfr_before (
		.din(new_net_546),
		.dout(new_net_545)
	);

	bfr new_net_547_bfr_before (
		.din(new_net_547),
		.dout(new_net_546)
	);

	bfr new_net_548_bfr_before (
		.din(new_net_548),
		.dout(new_net_547)
	);

	bfr new_net_549_bfr_before (
		.din(new_net_549),
		.dout(new_net_548)
	);

	spl2 N108_v_fanout (
		.a(N108),
		.b(new_net_148),
		.c(new_net_549)
	);

	bfr new_net_550_bfr_after (
		.din(N99),
		.dout(new_net_550)
	);

	bfr new_net_551_bfr_after (
		.din(new_net_550),
		.dout(new_net_551)
	);

	bfr new_net_552_bfr_after (
		.din(new_net_551),
		.dout(new_net_552)
	);

	bfr new_net_553_bfr_after (
		.din(new_net_552),
		.dout(new_net_553)
	);

	bfr new_net_554_bfr_after (
		.din(new_net_553),
		.dout(new_net_554)
	);

	bfr new_net_555_bfr_after (
		.din(new_net_554),
		.dout(new_net_555)
	);

	bfr new_net_556_bfr_after (
		.din(new_net_555),
		.dout(new_net_556)
	);

	bfr new_net_557_bfr_after (
		.din(new_net_556),
		.dout(new_net_557)
	);

	bfr new_net_558_bfr_after (
		.din(new_net_557),
		.dout(new_net_558)
	);

	bfr new_net_559_bfr_after (
		.din(new_net_558),
		.dout(new_net_559)
	);

	bfr new_net_560_bfr_after (
		.din(new_net_559),
		.dout(new_net_560)
	);

	bfr new_net_561_bfr_before (
		.din(new_net_561),
		.dout(new_net_56)
	);

	bfr new_net_562_bfr_before (
		.din(new_net_562),
		.dout(new_net_561)
	);

	bfr new_net_563_bfr_before (
		.din(new_net_563),
		.dout(new_net_562)
	);

	bfr new_net_564_bfr_before (
		.din(new_net_564),
		.dout(new_net_563)
	);

	bfr new_net_565_bfr_before (
		.din(new_net_565),
		.dout(new_net_564)
	);

	bfr new_net_566_bfr_before (
		.din(new_net_566),
		.dout(new_net_565)
	);

	bfr new_net_567_bfr_before (
		.din(new_net_567),
		.dout(new_net_566)
	);

	spl2 N99_v_fanout (
		.a(new_net_560),
		.b(new_net_55),
		.c(new_net_567)
	);

	bfr new_net_568_bfr_after (
		.din(N92),
		.dout(new_net_568)
	);

	bfr new_net_569_bfr_after (
		.din(new_net_568),
		.dout(new_net_569)
	);

	bfr new_net_570_bfr_after (
		.din(new_net_569),
		.dout(new_net_570)
	);

	bfr new_net_571_bfr_after (
		.din(new_net_570),
		.dout(new_net_571)
	);

	bfr new_net_572_bfr_after (
		.din(new_net_571),
		.dout(new_net_572)
	);

	bfr new_net_573_bfr_after (
		.din(new_net_572),
		.dout(new_net_573)
	);

	bfr new_net_574_bfr_after (
		.din(new_net_573),
		.dout(new_net_574)
	);

	bfr new_net_575_bfr_after (
		.din(new_net_574),
		.dout(new_net_575)
	);

	bfr new_net_576_bfr_after (
		.din(new_net_575),
		.dout(new_net_576)
	);

	bfr new_net_577_bfr_after (
		.din(new_net_576),
		.dout(new_net_577)
	);

	bfr new_net_578_bfr_after (
		.din(new_net_577),
		.dout(new_net_578)
	);

	bfr new_net_579_bfr_after (
		.din(new_net_578),
		.dout(new_net_579)
	);

	bfr new_net_580_bfr_after (
		.din(new_net_579),
		.dout(new_net_580)
	);

	bfr new_net_581_bfr_after (
		.din(new_net_580),
		.dout(new_net_581)
	);

	bfr new_net_582_bfr_after (
		.din(new_net_581),
		.dout(new_net_582)
	);

	bfr new_net_583_bfr_after (
		.din(new_net_582),
		.dout(new_net_583)
	);

	bfr new_net_584_bfr_after (
		.din(new_net_583),
		.dout(new_net_584)
	);

	bfr new_net_585_bfr_after (
		.din(new_net_584),
		.dout(new_net_585)
	);

	bfr new_net_586_bfr_after (
		.din(new_net_585),
		.dout(new_net_586)
	);

	bfr new_net_587_bfr_after (
		.din(new_net_586),
		.dout(new_net_587)
	);

	bfr new_net_588_bfr_after (
		.din(new_net_587),
		.dout(new_net_588)
	);

	bfr new_net_589_bfr_before (
		.din(new_net_589),
		.dout(new_net_153)
	);

	bfr new_net_590_bfr_before (
		.din(new_net_590),
		.dout(new_net_589)
	);

	bfr new_net_591_bfr_before (
		.din(new_net_591),
		.dout(new_net_590)
	);

	bfr new_net_592_bfr_before (
		.din(new_net_592),
		.dout(new_net_591)
	);

	bfr new_net_593_bfr_before (
		.din(new_net_593),
		.dout(new_net_592)
	);

	bfr new_net_594_bfr_before (
		.din(new_net_594),
		.dout(new_net_593)
	);

	bfr new_net_595_bfr_before (
		.din(new_net_595),
		.dout(new_net_594)
	);

	bfr new_net_596_bfr_before (
		.din(new_net_596),
		.dout(new_net_595)
	);

	spl2 N92_v_fanout (
		.a(new_net_588),
		.b(new_net_152),
		.c(new_net_596)
	);

	bfr new_net_597_bfr_before (
		.din(new_net_597),
		.dout(new_net_58)
	);

	bfr new_net_598_bfr_before (
		.din(new_net_598),
		.dout(new_net_597)
	);

	bfr new_net_599_bfr_before (
		.din(new_net_599),
		.dout(new_net_598)
	);

	bfr new_net_600_bfr_before (
		.din(new_net_600),
		.dout(new_net_599)
	);

	bfr new_net_601_bfr_before (
		.din(new_net_601),
		.dout(new_net_600)
	);

	bfr new_net_602_bfr_before (
		.din(new_net_602),
		.dout(new_net_601)
	);

	bfr new_net_603_bfr_before (
		.din(new_net_603),
		.dout(new_net_602)
	);

	bfr new_net_604_bfr_before (
		.din(new_net_604),
		.dout(new_net_603)
	);

	bfr new_net_605_bfr_before (
		.din(new_net_605),
		.dout(new_net_604)
	);

	spl2 N82_v_fanout (
		.a(N82),
		.b(new_net_57),
		.c(new_net_605)
	);

	bfr new_net_606_bfr_after (
		.din(N8),
		.dout(new_net_606)
	);

	bfr new_net_607_bfr_after (
		.din(new_net_606),
		.dout(new_net_607)
	);

	bfr new_net_608_bfr_after (
		.din(new_net_607),
		.dout(new_net_608)
	);

	bfr new_net_609_bfr_after (
		.din(new_net_608),
		.dout(new_net_609)
	);

	bfr new_net_610_bfr_after (
		.din(new_net_609),
		.dout(new_net_610)
	);

	bfr new_net_611_bfr_after (
		.din(new_net_610),
		.dout(new_net_611)
	);

	bfr new_net_612_bfr_after (
		.din(new_net_611),
		.dout(new_net_612)
	);

	bfr new_net_613_bfr_after (
		.din(new_net_612),
		.dout(new_net_613)
	);

	bfr new_net_614_bfr_after (
		.din(new_net_613),
		.dout(new_net_614)
	);

	bfr new_net_615_bfr_after (
		.din(new_net_614),
		.dout(new_net_615)
	);

	bfr new_net_616_bfr_after (
		.din(new_net_615),
		.dout(new_net_616)
	);

	bfr new_net_617_bfr_before (
		.din(new_net_617),
		.dout(new_net_32)
	);

	bfr new_net_618_bfr_before (
		.din(new_net_618),
		.dout(new_net_617)
	);

	bfr new_net_619_bfr_before (
		.din(new_net_619),
		.dout(new_net_618)
	);

	bfr new_net_620_bfr_before (
		.din(new_net_620),
		.dout(new_net_619)
	);

	bfr new_net_621_bfr_before (
		.din(new_net_621),
		.dout(new_net_620)
	);

	bfr new_net_622_bfr_before (
		.din(new_net_622),
		.dout(new_net_621)
	);

	bfr new_net_623_bfr_before (
		.din(new_net_623),
		.dout(new_net_622)
	);

	spl2 N8_v_fanout (
		.a(new_net_616),
		.b(new_net_31),
		.c(new_net_623)
	);

	bfr new_net_624_bfr_after (
		.din(N34),
		.dout(new_net_624)
	);

	bfr new_net_625_bfr_after (
		.din(new_net_624),
		.dout(new_net_625)
	);

	bfr new_net_626_bfr_after (
		.din(new_net_625),
		.dout(new_net_626)
	);

	bfr new_net_627_bfr_after (
		.din(new_net_626),
		.dout(new_net_627)
	);

	bfr new_net_628_bfr_after (
		.din(new_net_627),
		.dout(new_net_628)
	);

	bfr new_net_629_bfr_after (
		.din(new_net_628),
		.dout(new_net_629)
	);

	bfr new_net_630_bfr_after (
		.din(new_net_629),
		.dout(new_net_630)
	);

	bfr new_net_631_bfr_after (
		.din(new_net_630),
		.dout(new_net_631)
	);

	bfr new_net_632_bfr_after (
		.din(new_net_631),
		.dout(new_net_632)
	);

	bfr new_net_633_bfr_after (
		.din(new_net_632),
		.dout(new_net_633)
	);

	bfr new_net_634_bfr_after (
		.din(new_net_633),
		.dout(new_net_634)
	);

	bfr new_net_635_bfr_before (
		.din(new_net_635),
		.dout(new_net_26)
	);

	bfr new_net_636_bfr_before (
		.din(new_net_636),
		.dout(new_net_635)
	);

	bfr new_net_637_bfr_before (
		.din(new_net_637),
		.dout(new_net_636)
	);

	bfr new_net_638_bfr_before (
		.din(new_net_638),
		.dout(new_net_637)
	);

	bfr new_net_639_bfr_before (
		.din(new_net_639),
		.dout(new_net_638)
	);

	bfr new_net_640_bfr_before (
		.din(new_net_640),
		.dout(new_net_639)
	);

	bfr new_net_641_bfr_before (
		.din(new_net_641),
		.dout(new_net_640)
	);

	spl2 N34_v_fanout (
		.a(new_net_634),
		.b(new_net_25),
		.c(new_net_641)
	);

	bfr new_net_642_bfr_after (
		.din(N115),
		.dout(new_net_642)
	);

	bfr new_net_643_bfr_after (
		.din(new_net_642),
		.dout(new_net_643)
	);

	bfr new_net_644_bfr_after (
		.din(new_net_643),
		.dout(new_net_644)
	);

	bfr new_net_645_bfr_after (
		.din(new_net_644),
		.dout(new_net_645)
	);

	bfr new_net_646_bfr_after (
		.din(new_net_645),
		.dout(new_net_646)
	);

	bfr new_net_647_bfr_after (
		.din(new_net_646),
		.dout(new_net_647)
	);

	bfr new_net_648_bfr_after (
		.din(new_net_647),
		.dout(new_net_648)
	);

	bfr new_net_649_bfr_after (
		.din(new_net_648),
		.dout(new_net_649)
	);

	bfr new_net_650_bfr_after (
		.din(new_net_649),
		.dout(new_net_650)
	);

	bfr new_net_651_bfr_after (
		.din(new_net_650),
		.dout(new_net_651)
	);

	bfr new_net_652_bfr_after (
		.din(new_net_651),
		.dout(new_net_652)
	);

	bfr new_net_653_bfr_after (
		.din(new_net_652),
		.dout(new_net_653)
	);

	bfr new_net_654_bfr_after (
		.din(new_net_653),
		.dout(new_net_654)
	);

	bfr new_net_655_bfr_after (
		.din(new_net_654),
		.dout(new_net_655)
	);

	bfr new_net_656_bfr_after (
		.din(new_net_655),
		.dout(new_net_656)
	);

	bfr new_net_657_bfr_after (
		.din(new_net_656),
		.dout(new_net_657)
	);

	bfr new_net_658_bfr_after (
		.din(new_net_657),
		.dout(new_net_658)
	);

	bfr new_net_659_bfr_after (
		.din(new_net_658),
		.dout(new_net_659)
	);

	bfr new_net_660_bfr_after (
		.din(new_net_659),
		.dout(new_net_660)
	);

	bfr new_net_661_bfr_after (
		.din(new_net_660),
		.dout(new_net_661)
	);

	bfr new_net_662_bfr_after (
		.din(new_net_661),
		.dout(new_net_662)
	);

	bfr new_net_663_bfr_before (
		.din(new_net_663),
		.dout(new_net_70)
	);

	bfr new_net_664_bfr_before (
		.din(new_net_664),
		.dout(new_net_663)
	);

	bfr new_net_665_bfr_before (
		.din(new_net_665),
		.dout(new_net_664)
	);

	bfr new_net_666_bfr_before (
		.din(new_net_666),
		.dout(new_net_665)
	);

	bfr new_net_667_bfr_before (
		.din(new_net_667),
		.dout(new_net_666)
	);

	bfr new_net_668_bfr_before (
		.din(new_net_668),
		.dout(new_net_667)
	);

	bfr new_net_669_bfr_before (
		.din(new_net_669),
		.dout(new_net_668)
	);

	bfr new_net_670_bfr_before (
		.din(new_net_670),
		.dout(new_net_669)
	);

	spl2 N115_v_fanout (
		.a(new_net_662),
		.b(new_net_69),
		.c(new_net_670)
	);

	bfr new_net_671_bfr_before (
		.din(new_net_671),
		.dout(new_net_139)
	);

	bfr new_net_672_bfr_before (
		.din(new_net_672),
		.dout(new_net_671)
	);

	bfr new_net_673_bfr_before (
		.din(new_net_673),
		.dout(new_net_672)
	);

	bfr new_net_674_bfr_before (
		.din(new_net_674),
		.dout(new_net_673)
	);

	bfr new_net_675_bfr_before (
		.din(new_net_675),
		.dout(new_net_674)
	);

	bfr new_net_676_bfr_before (
		.din(new_net_676),
		.dout(new_net_675)
	);

	bfr new_net_677_bfr_before (
		.din(new_net_677),
		.dout(new_net_676)
	);

	bfr new_net_678_bfr_before (
		.din(new_net_678),
		.dout(new_net_677)
	);

	spl2 N76_v_fanout (
		.a(N76),
		.b(new_net_138),
		.c(new_net_678)
	);

	bfr new_net_679_bfr_after (
		.din(N40),
		.dout(new_net_679)
	);

	bfr new_net_680_bfr_after (
		.din(new_net_679),
		.dout(new_net_680)
	);

	bfr new_net_681_bfr_after (
		.din(new_net_680),
		.dout(new_net_681)
	);

	bfr new_net_682_bfr_after (
		.din(new_net_681),
		.dout(new_net_682)
	);

	bfr new_net_683_bfr_after (
		.din(new_net_682),
		.dout(new_net_683)
	);

	bfr new_net_684_bfr_after (
		.din(new_net_683),
		.dout(new_net_684)
	);

	bfr new_net_685_bfr_after (
		.din(new_net_684),
		.dout(new_net_685)
	);

	bfr new_net_686_bfr_after (
		.din(new_net_685),
		.dout(new_net_686)
	);

	bfr new_net_687_bfr_after (
		.din(new_net_686),
		.dout(new_net_687)
	);

	bfr new_net_688_bfr_after (
		.din(new_net_687),
		.dout(new_net_688)
	);

	bfr new_net_689_bfr_after (
		.din(new_net_688),
		.dout(new_net_689)
	);

	bfr new_net_690_bfr_after (
		.din(new_net_689),
		.dout(new_net_690)
	);

	bfr new_net_691_bfr_after (
		.din(new_net_690),
		.dout(new_net_691)
	);

	bfr new_net_692_bfr_after (
		.din(new_net_691),
		.dout(new_net_692)
	);

	bfr new_net_693_bfr_after (
		.din(new_net_692),
		.dout(new_net_693)
	);

	bfr new_net_694_bfr_after (
		.din(new_net_693),
		.dout(new_net_694)
	);

	bfr new_net_695_bfr_after (
		.din(new_net_694),
		.dout(new_net_695)
	);

	bfr new_net_696_bfr_after (
		.din(new_net_695),
		.dout(new_net_696)
	);

	bfr new_net_697_bfr_after (
		.din(new_net_696),
		.dout(new_net_697)
	);

	bfr new_net_698_bfr_after (
		.din(new_net_697),
		.dout(new_net_698)
	);

	bfr new_net_699_bfr_after (
		.din(new_net_698),
		.dout(new_net_699)
	);

	bfr new_net_700_bfr_before (
		.din(new_net_700),
		.dout(new_net_16)
	);

	bfr new_net_701_bfr_before (
		.din(new_net_701),
		.dout(new_net_700)
	);

	bfr new_net_702_bfr_before (
		.din(new_net_702),
		.dout(new_net_701)
	);

	bfr new_net_703_bfr_before (
		.din(new_net_703),
		.dout(new_net_702)
	);

	bfr new_net_704_bfr_before (
		.din(new_net_704),
		.dout(new_net_703)
	);

	bfr new_net_705_bfr_before (
		.din(new_net_705),
		.dout(new_net_704)
	);

	bfr new_net_706_bfr_before (
		.din(new_net_706),
		.dout(new_net_705)
	);

	bfr new_net_707_bfr_before (
		.din(new_net_707),
		.dout(new_net_706)
	);

	spl2 N40_v_fanout (
		.a(new_net_699),
		.b(new_net_15),
		.c(new_net_707)
	);

	bfr new_net_708_bfr_before (
		.din(new_net_708),
		.dout(new_net_54)
	);

	bfr new_net_709_bfr_before (
		.din(new_net_709),
		.dout(new_net_708)
	);

	bfr new_net_710_bfr_before (
		.din(new_net_710),
		.dout(new_net_709)
	);

	bfr new_net_711_bfr_before (
		.din(new_net_711),
		.dout(new_net_710)
	);

	bfr new_net_712_bfr_before (
		.din(new_net_712),
		.dout(new_net_711)
	);

	bfr new_net_713_bfr_before (
		.din(new_net_713),
		.dout(new_net_712)
	);

	bfr new_net_714_bfr_before (
		.din(new_net_714),
		.dout(new_net_713)
	);

	bfr new_net_715_bfr_before (
		.din(new_net_715),
		.dout(new_net_714)
	);

	spl2 N1_v_fanout (
		.a(N1),
		.b(new_net_53),
		.c(new_net_715)
	);

	bfr new_net_716_bfr_after (
		.din(N14),
		.dout(new_net_716)
	);

	bfr new_net_717_bfr_after (
		.din(new_net_716),
		.dout(new_net_717)
	);

	bfr new_net_718_bfr_after (
		.din(new_net_717),
		.dout(new_net_718)
	);

	bfr new_net_719_bfr_after (
		.din(new_net_718),
		.dout(new_net_719)
	);

	bfr new_net_720_bfr_after (
		.din(new_net_719),
		.dout(new_net_720)
	);

	bfr new_net_721_bfr_after (
		.din(new_net_720),
		.dout(new_net_721)
	);

	bfr new_net_722_bfr_after (
		.din(new_net_721),
		.dout(new_net_722)
	);

	bfr new_net_723_bfr_after (
		.din(new_net_722),
		.dout(new_net_723)
	);

	bfr new_net_724_bfr_after (
		.din(new_net_723),
		.dout(new_net_724)
	);

	bfr new_net_725_bfr_after (
		.din(new_net_724),
		.dout(new_net_725)
	);

	bfr new_net_726_bfr_after (
		.din(new_net_725),
		.dout(new_net_726)
	);

	bfr new_net_727_bfr_after (
		.din(new_net_726),
		.dout(new_net_727)
	);

	bfr new_net_728_bfr_after (
		.din(new_net_727),
		.dout(new_net_728)
	);

	bfr new_net_729_bfr_after (
		.din(new_net_728),
		.dout(new_net_729)
	);

	bfr new_net_730_bfr_after (
		.din(new_net_729),
		.dout(new_net_730)
	);

	bfr new_net_731_bfr_after (
		.din(new_net_730),
		.dout(new_net_731)
	);

	bfr new_net_732_bfr_after (
		.din(new_net_731),
		.dout(new_net_732)
	);

	bfr new_net_733_bfr_after (
		.din(new_net_732),
		.dout(new_net_733)
	);

	bfr new_net_734_bfr_after (
		.din(new_net_733),
		.dout(new_net_734)
	);

	bfr new_net_735_bfr_after (
		.din(new_net_734),
		.dout(new_net_735)
	);

	bfr new_net_736_bfr_after (
		.din(new_net_735),
		.dout(new_net_736)
	);

	bfr new_net_737_bfr_before (
		.din(new_net_737),
		.dout(new_net_96)
	);

	bfr new_net_738_bfr_before (
		.din(new_net_738),
		.dout(new_net_737)
	);

	bfr new_net_739_bfr_before (
		.din(new_net_739),
		.dout(new_net_738)
	);

	bfr new_net_740_bfr_before (
		.din(new_net_740),
		.dout(new_net_739)
	);

	bfr new_net_741_bfr_before (
		.din(new_net_741),
		.dout(new_net_740)
	);

	bfr new_net_742_bfr_before (
		.din(new_net_742),
		.dout(new_net_741)
	);

	bfr new_net_743_bfr_before (
		.din(new_net_743),
		.dout(new_net_742)
	);

	bfr new_net_744_bfr_before (
		.din(new_net_744),
		.dout(new_net_743)
	);

	spl2 N14_v_fanout (
		.a(new_net_736),
		.b(new_net_95),
		.c(new_net_744)
	);

	bfr new_net_745_bfr_before (
		.din(new_net_745),
		.dout(new_net_133)
	);

	bfr new_net_746_bfr_before (
		.din(new_net_746),
		.dout(new_net_745)
	);

	bfr new_net_747_bfr_before (
		.din(new_net_747),
		.dout(new_net_746)
	);

	bfr new_net_748_bfr_before (
		.din(new_net_748),
		.dout(new_net_747)
	);

	bfr new_net_749_bfr_before (
		.din(new_net_749),
		.dout(new_net_748)
	);

	bfr new_net_750_bfr_before (
		.din(new_net_750),
		.dout(new_net_749)
	);

	bfr new_net_751_bfr_before (
		.din(new_net_751),
		.dout(new_net_750)
	);

	bfr new_net_752_bfr_before (
		.din(new_net_752),
		.dout(new_net_751)
	);

	spl2 N89_v_fanout (
		.a(N89),
		.b(new_net_132),
		.c(new_net_752)
	);

	bfr new_net_753_bfr_after (
		.din(N79),
		.dout(new_net_753)
	);

	bfr new_net_754_bfr_after (
		.din(new_net_753),
		.dout(new_net_754)
	);

	bfr new_net_755_bfr_after (
		.din(new_net_754),
		.dout(new_net_755)
	);

	bfr new_net_756_bfr_after (
		.din(new_net_755),
		.dout(new_net_756)
	);

	bfr new_net_757_bfr_after (
		.din(new_net_756),
		.dout(new_net_757)
	);

	bfr new_net_758_bfr_after (
		.din(new_net_757),
		.dout(new_net_758)
	);

	bfr new_net_759_bfr_after (
		.din(new_net_758),
		.dout(new_net_759)
	);

	bfr new_net_760_bfr_after (
		.din(new_net_759),
		.dout(new_net_760)
	);

	bfr new_net_761_bfr_after (
		.din(new_net_760),
		.dout(new_net_761)
	);

	bfr new_net_762_bfr_after (
		.din(new_net_761),
		.dout(new_net_762)
	);

	bfr new_net_763_bfr_after (
		.din(new_net_762),
		.dout(new_net_763)
	);

	bfr new_net_764_bfr_after (
		.din(new_net_763),
		.dout(new_net_764)
	);

	bfr new_net_765_bfr_after (
		.din(new_net_764),
		.dout(new_net_765)
	);

	bfr new_net_766_bfr_after (
		.din(new_net_765),
		.dout(new_net_766)
	);

	bfr new_net_767_bfr_after (
		.din(new_net_766),
		.dout(new_net_767)
	);

	bfr new_net_768_bfr_after (
		.din(new_net_767),
		.dout(new_net_768)
	);

	bfr new_net_769_bfr_after (
		.din(new_net_768),
		.dout(new_net_769)
	);

	bfr new_net_770_bfr_after (
		.din(new_net_769),
		.dout(new_net_770)
	);

	bfr new_net_771_bfr_after (
		.din(new_net_770),
		.dout(new_net_771)
	);

	bfr new_net_772_bfr_after (
		.din(new_net_771),
		.dout(new_net_772)
	);

	bfr new_net_773_bfr_after (
		.din(new_net_772),
		.dout(new_net_773)
	);

	bfr new_net_774_bfr_before (
		.din(new_net_774),
		.dout(new_net_159)
	);

	bfr new_net_775_bfr_before (
		.din(new_net_775),
		.dout(new_net_774)
	);

	bfr new_net_776_bfr_before (
		.din(new_net_776),
		.dout(new_net_775)
	);

	bfr new_net_777_bfr_before (
		.din(new_net_777),
		.dout(new_net_776)
	);

	bfr new_net_778_bfr_before (
		.din(new_net_778),
		.dout(new_net_777)
	);

	bfr new_net_779_bfr_before (
		.din(new_net_779),
		.dout(new_net_778)
	);

	bfr new_net_780_bfr_before (
		.din(new_net_780),
		.dout(new_net_779)
	);

	bfr new_net_781_bfr_before (
		.din(new_net_781),
		.dout(new_net_780)
	);

	spl2 N79_v_fanout (
		.a(new_net_773),
		.b(new_net_158),
		.c(new_net_781)
	);

	bfr new_net_782_bfr_after (
		.din(N53),
		.dout(new_net_782)
	);

	bfr new_net_783_bfr_after (
		.din(new_net_782),
		.dout(new_net_783)
	);

	bfr new_net_784_bfr_after (
		.din(new_net_783),
		.dout(new_net_784)
	);

	bfr new_net_785_bfr_after (
		.din(new_net_784),
		.dout(new_net_785)
	);

	bfr new_net_786_bfr_after (
		.din(new_net_785),
		.dout(new_net_786)
	);

	bfr new_net_787_bfr_after (
		.din(new_net_786),
		.dout(new_net_787)
	);

	bfr new_net_788_bfr_after (
		.din(new_net_787),
		.dout(new_net_788)
	);

	bfr new_net_789_bfr_after (
		.din(new_net_788),
		.dout(new_net_789)
	);

	bfr new_net_790_bfr_after (
		.din(new_net_789),
		.dout(new_net_790)
	);

	bfr new_net_791_bfr_after (
		.din(new_net_790),
		.dout(new_net_791)
	);

	bfr new_net_792_bfr_after (
		.din(new_net_791),
		.dout(new_net_792)
	);

	bfr new_net_793_bfr_after (
		.din(new_net_792),
		.dout(new_net_793)
	);

	bfr new_net_794_bfr_after (
		.din(new_net_793),
		.dout(new_net_794)
	);

	bfr new_net_795_bfr_after (
		.din(new_net_794),
		.dout(new_net_795)
	);

	bfr new_net_796_bfr_after (
		.din(new_net_795),
		.dout(new_net_796)
	);

	bfr new_net_797_bfr_after (
		.din(new_net_796),
		.dout(new_net_797)
	);

	bfr new_net_798_bfr_after (
		.din(new_net_797),
		.dout(new_net_798)
	);

	bfr new_net_799_bfr_after (
		.din(new_net_798),
		.dout(new_net_799)
	);

	bfr new_net_800_bfr_after (
		.din(new_net_799),
		.dout(new_net_800)
	);

	bfr new_net_801_bfr_after (
		.din(new_net_800),
		.dout(new_net_801)
	);

	bfr new_net_802_bfr_after (
		.din(new_net_801),
		.dout(new_net_802)
	);

	bfr new_net_803_bfr_before (
		.din(new_net_803),
		.dout(new_net_72)
	);

	bfr new_net_804_bfr_before (
		.din(new_net_804),
		.dout(new_net_803)
	);

	bfr new_net_805_bfr_before (
		.din(new_net_805),
		.dout(new_net_804)
	);

	bfr new_net_806_bfr_before (
		.din(new_net_806),
		.dout(new_net_805)
	);

	bfr new_net_807_bfr_before (
		.din(new_net_807),
		.dout(new_net_806)
	);

	bfr new_net_808_bfr_before (
		.din(new_net_808),
		.dout(new_net_807)
	);

	bfr new_net_809_bfr_before (
		.din(new_net_809),
		.dout(new_net_808)
	);

	bfr new_net_810_bfr_before (
		.din(new_net_810),
		.dout(new_net_809)
	);

	spl2 N53_v_fanout (
		.a(new_net_802),
		.b(new_net_71),
		.c(new_net_810)
	);

	bfr new_net_811_bfr_after (
		.din(N73),
		.dout(new_net_811)
	);

	bfr new_net_812_bfr_after (
		.din(new_net_811),
		.dout(new_net_812)
	);

	bfr new_net_813_bfr_after (
		.din(new_net_812),
		.dout(new_net_813)
	);

	bfr new_net_814_bfr_after (
		.din(new_net_813),
		.dout(new_net_814)
	);

	bfr new_net_815_bfr_after (
		.din(new_net_814),
		.dout(new_net_815)
	);

	bfr new_net_816_bfr_after (
		.din(new_net_815),
		.dout(new_net_816)
	);

	bfr new_net_817_bfr_after (
		.din(new_net_816),
		.dout(new_net_817)
	);

	bfr new_net_818_bfr_after (
		.din(new_net_817),
		.dout(new_net_818)
	);

	bfr new_net_819_bfr_after (
		.din(new_net_818),
		.dout(new_net_819)
	);

	bfr new_net_820_bfr_after (
		.din(new_net_819),
		.dout(new_net_820)
	);

	bfr new_net_821_bfr_after (
		.din(new_net_820),
		.dout(new_net_821)
	);

	bfr new_net_822_bfr_before (
		.din(new_net_822),
		.dout(new_net_92)
	);

	bfr new_net_823_bfr_before (
		.din(new_net_823),
		.dout(new_net_822)
	);

	bfr new_net_824_bfr_before (
		.din(new_net_824),
		.dout(new_net_823)
	);

	bfr new_net_825_bfr_before (
		.din(new_net_825),
		.dout(new_net_824)
	);

	bfr new_net_826_bfr_before (
		.din(new_net_826),
		.dout(new_net_825)
	);

	bfr new_net_827_bfr_before (
		.din(new_net_827),
		.dout(new_net_826)
	);

	bfr new_net_828_bfr_before (
		.din(new_net_828),
		.dout(new_net_827)
	);

	spl2 N73_v_fanout (
		.a(new_net_821),
		.b(new_net_91),
		.c(new_net_828)
	);

	bfr new_net_829_bfr_before (
		.din(new_net_829),
		.dout(new_net_113)
	);

	bfr new_net_830_bfr_before (
		.din(new_net_830),
		.dout(new_net_829)
	);

	bfr new_net_831_bfr_before (
		.din(new_net_831),
		.dout(new_net_830)
	);

	bfr new_net_832_bfr_before (
		.din(new_net_832),
		.dout(new_net_831)
	);

	bfr new_net_833_bfr_before (
		.din(new_net_833),
		.dout(new_net_832)
	);

	bfr new_net_834_bfr_before (
		.din(new_net_834),
		.dout(new_net_833)
	);

	bfr new_net_835_bfr_before (
		.din(new_net_835),
		.dout(new_net_834)
	);

	bfr new_net_836_bfr_before (
		.din(new_net_836),
		.dout(new_net_835)
	);

	bfr new_net_837_bfr_before (
		.din(new_net_837),
		.dout(new_net_836)
	);

	spl2 N56_v_fanout (
		.a(N56),
		.b(new_net_112),
		.c(new_net_837)
	);

	bfr new_net_838_bfr_before (
		.din(new_net_838),
		.dout(new_net_143)
	);

	bfr new_net_839_bfr_before (
		.din(new_net_839),
		.dout(new_net_838)
	);

	bfr new_net_840_bfr_before (
		.din(new_net_840),
		.dout(new_net_839)
	);

	bfr new_net_841_bfr_before (
		.din(new_net_841),
		.dout(new_net_840)
	);

	bfr new_net_842_bfr_before (
		.din(new_net_842),
		.dout(new_net_841)
	);

	bfr new_net_843_bfr_before (
		.din(new_net_843),
		.dout(new_net_842)
	);

	bfr new_net_844_bfr_before (
		.din(new_net_844),
		.dout(new_net_843)
	);

	bfr new_net_845_bfr_before (
		.din(new_net_845),
		.dout(new_net_844)
	);

	bfr new_net_846_bfr_before (
		.din(new_net_846),
		.dout(new_net_845)
	);

	spl2 N17_v_fanout (
		.a(N17),
		.b(new_net_142),
		.c(new_net_846)
	);

	bfr new_net_847_bfr_before (
		.din(new_net_847),
		.dout(new_net_74)
	);

	bfr new_net_848_bfr_before (
		.din(new_net_848),
		.dout(new_net_847)
	);

	bfr new_net_849_bfr_before (
		.din(new_net_849),
		.dout(new_net_848)
	);

	bfr new_net_850_bfr_before (
		.din(new_net_850),
		.dout(new_net_849)
	);

	bfr new_net_851_bfr_before (
		.din(new_net_851),
		.dout(new_net_850)
	);

	bfr new_net_852_bfr_before (
		.din(new_net_852),
		.dout(new_net_851)
	);

	bfr new_net_853_bfr_before (
		.din(new_net_853),
		.dout(new_net_852)
	);

	bfr new_net_854_bfr_before (
		.din(new_net_854),
		.dout(new_net_853)
	);

	spl2 N102_v_fanout (
		.a(N102),
		.b(new_net_73),
		.c(new_net_854)
	);

	bfr new_net_855_bfr_before (
		.din(new_net_855),
		.dout(new_net_76)
	);

	bfr new_net_856_bfr_before (
		.din(new_net_856),
		.dout(new_net_855)
	);

	bfr new_net_857_bfr_before (
		.din(new_net_857),
		.dout(new_net_856)
	);

	bfr new_net_858_bfr_before (
		.din(new_net_858),
		.dout(new_net_857)
	);

	bfr new_net_859_bfr_before (
		.din(new_net_859),
		.dout(new_net_858)
	);

	bfr new_net_860_bfr_before (
		.din(new_net_860),
		.dout(new_net_859)
	);

	bfr new_net_861_bfr_before (
		.din(new_net_861),
		.dout(new_net_860)
	);

	bfr new_net_862_bfr_before (
		.din(new_net_862),
		.dout(new_net_861)
	);

	spl2 N37_v_fanout (
		.a(N37),
		.b(new_net_75),
		.c(new_net_862)
	);

	bfr new_net_863_bfr_before (
		.din(new_net_863),
		.dout(new_net_64)
	);

	bfr new_net_864_bfr_before (
		.din(new_net_864),
		.dout(new_net_863)
	);

	bfr new_net_865_bfr_before (
		.din(new_net_865),
		.dout(new_net_864)
	);

	bfr new_net_866_bfr_before (
		.din(new_net_866),
		.dout(new_net_865)
	);

	bfr new_net_867_bfr_before (
		.din(new_net_867),
		.dout(new_net_866)
	);

	bfr new_net_868_bfr_before (
		.din(new_net_868),
		.dout(new_net_867)
	);

	bfr new_net_869_bfr_before (
		.din(new_net_869),
		.dout(new_net_868)
	);

	bfr new_net_870_bfr_before (
		.din(new_net_870),
		.dout(new_net_869)
	);

	bfr new_net_871_bfr_before (
		.din(new_net_871),
		.dout(new_net_870)
	);

	spl2 N43_v_fanout (
		.a(N43),
		.b(new_net_63),
		.c(new_net_871)
	);

	bfr new_net_872_bfr_before (
		.din(new_net_872),
		.dout(new_net_36)
	);

	bfr new_net_873_bfr_before (
		.din(new_net_873),
		.dout(new_net_872)
	);

	bfr new_net_874_bfr_before (
		.din(new_net_874),
		.dout(new_net_873)
	);

	bfr new_net_875_bfr_before (
		.din(new_net_875),
		.dout(new_net_874)
	);

	bfr new_net_876_bfr_before (
		.din(new_net_876),
		.dout(new_net_875)
	);

	bfr new_net_877_bfr_before (
		.din(new_net_877),
		.dout(new_net_876)
	);

	bfr new_net_878_bfr_before (
		.din(new_net_878),
		.dout(new_net_877)
	);

	bfr new_net_879_bfr_before (
		.din(new_net_879),
		.dout(new_net_878)
	);

	spl2 N69_v_fanout (
		.a(N69),
		.b(new_net_35),
		.c(new_net_879)
	);

	bfr new_net_880_bfr_before (
		.din(new_net_880),
		.dout(new_net_135)
	);

	bfr new_net_881_bfr_before (
		.din(new_net_881),
		.dout(new_net_880)
	);

	bfr new_net_882_bfr_before (
		.din(new_net_882),
		.dout(new_net_881)
	);

	bfr new_net_883_bfr_before (
		.din(new_net_883),
		.dout(new_net_882)
	);

	bfr new_net_884_bfr_before (
		.din(new_net_884),
		.dout(new_net_883)
	);

	bfr new_net_885_bfr_before (
		.din(new_net_885),
		.dout(new_net_884)
	);

	bfr new_net_886_bfr_before (
		.din(new_net_886),
		.dout(new_net_885)
	);

	bfr new_net_887_bfr_before (
		.din(new_net_887),
		.dout(new_net_886)
	);

	spl2 N30_v_fanout (
		.a(N30),
		.b(new_net_134),
		.c(new_net_887)
	);

	bfr new_net_888_bfr_after (
		.din(N27),
		.dout(new_net_888)
	);

	bfr new_net_889_bfr_after (
		.din(new_net_888),
		.dout(new_net_889)
	);

	bfr new_net_890_bfr_after (
		.din(new_net_889),
		.dout(new_net_890)
	);

	bfr new_net_891_bfr_after (
		.din(new_net_890),
		.dout(new_net_891)
	);

	bfr new_net_892_bfr_after (
		.din(new_net_891),
		.dout(new_net_892)
	);

	bfr new_net_893_bfr_after (
		.din(new_net_892),
		.dout(new_net_893)
	);

	bfr new_net_894_bfr_after (
		.din(new_net_893),
		.dout(new_net_894)
	);

	bfr new_net_895_bfr_after (
		.din(new_net_894),
		.dout(new_net_895)
	);

	bfr new_net_896_bfr_after (
		.din(new_net_895),
		.dout(new_net_896)
	);

	bfr new_net_897_bfr_after (
		.din(new_net_896),
		.dout(new_net_897)
	);

	bfr new_net_898_bfr_after (
		.din(new_net_897),
		.dout(new_net_898)
	);

	bfr new_net_899_bfr_after (
		.din(new_net_898),
		.dout(new_net_899)
	);

	bfr new_net_900_bfr_after (
		.din(new_net_899),
		.dout(new_net_900)
	);

	bfr new_net_901_bfr_after (
		.din(new_net_900),
		.dout(new_net_901)
	);

	bfr new_net_902_bfr_after (
		.din(new_net_901),
		.dout(new_net_902)
	);

	bfr new_net_903_bfr_after (
		.din(new_net_902),
		.dout(new_net_903)
	);

	bfr new_net_904_bfr_after (
		.din(new_net_903),
		.dout(new_net_904)
	);

	bfr new_net_905_bfr_after (
		.din(new_net_904),
		.dout(new_net_905)
	);

	bfr new_net_906_bfr_after (
		.din(new_net_905),
		.dout(new_net_906)
	);

	bfr new_net_907_bfr_after (
		.din(new_net_906),
		.dout(new_net_907)
	);

	bfr new_net_908_bfr_after (
		.din(new_net_907),
		.dout(new_net_908)
	);

	bfr new_net_909_bfr_before (
		.din(new_net_909),
		.dout(new_net_90)
	);

	bfr new_net_910_bfr_before (
		.din(new_net_910),
		.dout(new_net_909)
	);

	bfr new_net_911_bfr_before (
		.din(new_net_911),
		.dout(new_net_910)
	);

	bfr new_net_912_bfr_before (
		.din(new_net_912),
		.dout(new_net_911)
	);

	bfr new_net_913_bfr_before (
		.din(new_net_913),
		.dout(new_net_912)
	);

	bfr new_net_914_bfr_before (
		.din(new_net_914),
		.dout(new_net_913)
	);

	bfr new_net_915_bfr_before (
		.din(new_net_915),
		.dout(new_net_914)
	);

	bfr new_net_916_bfr_before (
		.din(new_net_916),
		.dout(new_net_915)
	);

	spl2 N27_v_fanout (
		.a(new_net_908),
		.b(new_net_89),
		.c(new_net_916)
	);

	bfr new_net_169_bfr_after (
		.din(N24),
		.dout(new_net_169)
	);

	bfr new_net_172_bfr_after (
		.din(N63),
		.dout(new_net_172)
	);

	bfr new_net_917_bfr_after (
		.din(new_net_192),
		.dout(new_net_917)
	);

	bfr new_net_918_bfr_after (
		.din(new_net_917),
		.dout(new_net_918)
	);

	bfr new_net_919_bfr_after (
		.din(new_net_918),
		.dout(new_net_919)
	);

	bfr new_net_920_bfr_after (
		.din(new_net_919),
		.dout(new_net_920)
	);

	bfr new_net_921_bfr_after (
		.din(new_net_920),
		.dout(new_net_921)
	);

	bfr new_net_922_bfr_after (
		.din(new_net_921),
		.dout(new_net_922)
	);

	bfr new_net_923_bfr_after (
		.din(new_net_922),
		.dout(new_net_923)
	);

	bfr new_net_924_bfr_after (
		.din(new_net_923),
		.dout(new_net_924)
	);

	bfr new_net_925_bfr_after (
		.din(new_net_924),
		.dout(new_net_925)
	);

	bfr new_net_926_bfr_after (
		.din(new_net_925),
		.dout(new_net_926)
	);

	bfr new_net_927_bfr_after (
		.din(new_net_926),
		.dout(new_net_927)
	);

	bfr new_net_928_bfr_after (
		.din(new_net_927),
		.dout(new_net_928)
	);

	bfr new_net_929_bfr_after (
		.din(new_net_928),
		.dout(new_net_929)
	);

	bfr new_net_930_bfr_after (
		.din(new_net_929),
		.dout(new_net_930)
	);

	bfr new_net_931_bfr_after (
		.din(new_net_930),
		.dout(new_net_931)
	);

	bfr new_net_932_bfr_after (
		.din(new_net_931),
		.dout(new_net_932)
	);

	bfr new_net_933_bfr_after (
		.din(new_net_932),
		.dout(new_net_933)
	);

	bfr new_net_934_bfr_after (
		.din(new_net_933),
		.dout(new_net_934)
	);

	bfr new_net_935_bfr_after (
		.din(new_net_934),
		.dout(new_net_935)
	);

	bfr new_net_936_bfr_after (
		.din(new_net_935),
		.dout(new_net_936)
	);

	bfr new_net_937_bfr_after (
		.din(new_net_936),
		.dout(new_net_937)
	);

	bfr new_net_938_bfr_after (
		.din(new_net_937),
		.dout(new_net_938)
	);

	bfr new_net_939_bfr_after (
		.din(new_net_938),
		.dout(new_net_939)
	);

	bfr new_net_940_bfr_after (
		.din(new_net_939),
		.dout(new_net_940)
	);

	bfr new_net_941_bfr_after (
		.din(new_net_940),
		.dout(new_net_941)
	);

	bfr new_net_942_bfr_after (
		.din(new_net_941),
		.dout(new_net_942)
	);

	bfr new_net_943_bfr_after (
		.din(new_net_942),
		.dout(new_net_943)
	);

	bfr new_net_944_bfr_after (
		.din(new_net_943),
		.dout(new_net_944)
	);

	bfr N223_bfr_after (
		.din(new_net_944),
		.dout(N223)
	);

	bfr new_net_188_bfr_after (
		.din(_050_),
		.dout(new_net_188)
	);

	bfr new_net_171_bfr_after (
		.din(_064_),
		.dout(new_net_171)
	);

	bfr new_net_178_bfr_after (
		.din(_099_),
		.dout(new_net_178)
	);

	bfr new_net_179_bfr_after (
		.din(_092_),
		.dout(new_net_179)
	);

	bfr new_net_945_bfr_after (
		.din(N66),
		.dout(new_net_945)
	);

	bfr new_net_946_bfr_after (
		.din(new_net_945),
		.dout(new_net_946)
	);

	bfr new_net_947_bfr_after (
		.din(new_net_946),
		.dout(new_net_947)
	);

	bfr new_net_948_bfr_after (
		.din(new_net_947),
		.dout(new_net_948)
	);

	bfr new_net_949_bfr_after (
		.din(new_net_948),
		.dout(new_net_949)
	);

	bfr new_net_950_bfr_after (
		.din(new_net_949),
		.dout(new_net_950)
	);

	bfr new_net_951_bfr_after (
		.din(new_net_950),
		.dout(new_net_951)
	);

	bfr new_net_952_bfr_after (
		.din(new_net_951),
		.dout(new_net_952)
	);

	bfr new_net_953_bfr_after (
		.din(new_net_952),
		.dout(new_net_953)
	);

	bfr new_net_954_bfr_after (
		.din(new_net_953),
		.dout(new_net_954)
	);

	bfr new_net_955_bfr_after (
		.din(new_net_954),
		.dout(new_net_955)
	);

	bfr new_net_956_bfr_after (
		.din(new_net_955),
		.dout(new_net_956)
	);

	bfr new_net_957_bfr_after (
		.din(new_net_956),
		.dout(new_net_957)
	);

	bfr new_net_958_bfr_after (
		.din(new_net_957),
		.dout(new_net_958)
	);

	bfr new_net_959_bfr_after (
		.din(new_net_958),
		.dout(new_net_959)
	);

	bfr new_net_960_bfr_after (
		.din(new_net_959),
		.dout(new_net_960)
	);

	bfr new_net_961_bfr_after (
		.din(new_net_960),
		.dout(new_net_961)
	);

	bfr new_net_962_bfr_after (
		.din(new_net_961),
		.dout(new_net_962)
	);

	bfr new_net_963_bfr_after (
		.din(new_net_962),
		.dout(new_net_963)
	);

	bfr new_net_964_bfr_after (
		.din(new_net_963),
		.dout(new_net_964)
	);

	bfr new_net_965_bfr_after (
		.din(new_net_964),
		.dout(new_net_965)
	);

	bfr new_net_181_bfr_after (
		.din(new_net_965),
		.dout(new_net_181)
	);

	bfr new_net_183_bfr_after (
		.din(_027_),
		.dout(new_net_183)
	);

	bfr new_net_186_bfr_after (
		.din(_039_),
		.dout(new_net_186)
	);

	bfr new_net_966_bfr_after (
		.din(_013_),
		.dout(new_net_966)
	);

	bfr new_net_184_bfr_after (
		.din(new_net_966),
		.dout(new_net_184)
	);

	bfr new_net_187_bfr_after (
		.din(_049_),
		.dout(new_net_187)
	);

	bfr new_net_182_bfr_after (
		.din(_016_),
		.dout(new_net_182)
	);

	bfr new_net_967_bfr_after (
		.din(_006_),
		.dout(new_net_967)
	);

	bfr new_net_185_bfr_after (
		.din(new_net_967),
		.dout(new_net_185)
	);

	bfr new_net_180_bfr_after (
		.din(_115_),
		.dout(new_net_180)
	);

	bfr new_net_173_bfr_after (
		.din(_070_),
		.dout(new_net_173)
	);

	bfr new_net_968_bfr_after (
		.din(new_net_196),
		.dout(new_net_968)
	);

	bfr N431_bfr_after (
		.din(new_net_968),
		.dout(N431)
	);

	bfr new_net_170_bfr_after (
		.din(_062_),
		.dout(new_net_170)
	);

	bfr new_net_174_bfr_after (
		.din(_074_),
		.dout(new_net_174)
	);

	bfr new_net_175_bfr_after (
		.din(_068_),
		.dout(new_net_175)
	);

	bfr new_net_969_bfr_after (
		.din(_063_),
		.dout(new_net_969)
	);

	bfr new_net_176_bfr_after (
		.din(new_net_969),
		.dout(new_net_176)
	);

	bfr new_net_177_bfr_after (
		.din(_102_),
		.dout(new_net_177)
	);

	bfr new_net_189_bfr_after (
		.din(_051_),
		.dout(new_net_189)
	);

	bfr new_net_970_bfr_after (
		.din(_054_),
		.dout(new_net_970)
	);

	bfr new_net_971_bfr_after (
		.din(new_net_970),
		.dout(new_net_971)
	);

	bfr new_net_972_bfr_after (
		.din(new_net_971),
		.dout(new_net_972)
	);

	bfr new_net_973_bfr_after (
		.din(new_net_972),
		.dout(new_net_973)
	);

	bfr new_net_974_bfr_after (
		.din(new_net_973),
		.dout(new_net_974)
	);

	bfr new_net_190_bfr_after (
		.din(new_net_974),
		.dout(new_net_190)
	);

	bfr new_net_191_bfr_after (
		.din(_058_),
		.dout(new_net_191)
	);

	bfr new_net_975_bfr_after (
		.din(new_net_198),
		.dout(new_net_975)
	);

	bfr new_net_976_bfr_after (
		.din(new_net_975),
		.dout(new_net_976)
	);

	bfr new_net_977_bfr_after (
		.din(new_net_976),
		.dout(new_net_977)
	);

	bfr new_net_978_bfr_after (
		.din(new_net_977),
		.dout(new_net_978)
	);

	bfr new_net_979_bfr_after (
		.din(new_net_978),
		.dout(new_net_979)
	);

	bfr new_net_980_bfr_after (
		.din(new_net_979),
		.dout(new_net_980)
	);

	bfr new_net_981_bfr_after (
		.din(new_net_980),
		.dout(new_net_981)
	);

	bfr N370_bfr_after (
		.din(new_net_981),
		.dout(N370)
	);

	bfr new_net_982_bfr_after (
		.din(new_net_194),
		.dout(new_net_982)
	);

	bfr new_net_983_bfr_after (
		.din(new_net_982),
		.dout(new_net_983)
	);

	bfr new_net_984_bfr_after (
		.din(new_net_983),
		.dout(new_net_984)
	);

	bfr new_net_985_bfr_after (
		.din(new_net_984),
		.dout(new_net_985)
	);

	bfr new_net_986_bfr_after (
		.din(new_net_985),
		.dout(new_net_986)
	);

	bfr new_net_987_bfr_after (
		.din(new_net_986),
		.dout(new_net_987)
	);

	bfr new_net_988_bfr_after (
		.din(new_net_987),
		.dout(new_net_988)
	);

	bfr new_net_989_bfr_after (
		.din(new_net_988),
		.dout(new_net_989)
	);

	bfr new_net_990_bfr_after (
		.din(new_net_989),
		.dout(new_net_990)
	);

	bfr new_net_991_bfr_after (
		.din(new_net_990),
		.dout(new_net_991)
	);

	bfr new_net_992_bfr_after (
		.din(new_net_991),
		.dout(new_net_992)
	);

	bfr new_net_993_bfr_after (
		.din(new_net_992),
		.dout(new_net_993)
	);

	bfr new_net_994_bfr_after (
		.din(new_net_993),
		.dout(new_net_994)
	);

	bfr new_net_995_bfr_after (
		.din(new_net_994),
		.dout(new_net_995)
	);

	bfr new_net_996_bfr_after (
		.din(new_net_995),
		.dout(new_net_996)
	);

	bfr new_net_997_bfr_after (
		.din(new_net_996),
		.dout(new_net_997)
	);

	bfr new_net_998_bfr_after (
		.din(new_net_997),
		.dout(new_net_998)
	);

	bfr new_net_999_bfr_after (
		.din(new_net_998),
		.dout(new_net_999)
	);

	bfr N329_bfr_after (
		.din(new_net_999),
		.dout(N329)
	);

endmodule