module c6288(N426,N154,N358,N69,N18,N443,N494,N222,N171,N477,N273,N392,N52,N375,N290,N1,N103,N188,N205,N256,N409,N86,N137,N511,N307,N35,N460,N239,N324,N341,N528,N120);
    wire new_Jinkela_wire_6612;
    wire new_Jinkela_wire_20206;
    wire _0481_;
    wire new_Jinkela_wire_16010;
    wire new_Jinkela_wire_18474;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_1559;
    wire _1686_;
    wire new_Jinkela_wire_7233;
    wire new_Jinkela_wire_12649;
    wire new_Jinkela_wire_17249;
    wire new_Jinkela_wire_19210;
    wire new_Jinkela_wire_11193;
    wire new_Jinkela_wire_2733;
    wire new_Jinkela_wire_17546;
    wire new_Jinkela_wire_4695;
    wire new_Jinkela_wire_8412;
    wire _0807_;
    wire new_Jinkela_wire_8507;
    wire new_Jinkela_wire_7584;
    wire _0152_;
    wire _1666_;
    wire new_Jinkela_wire_13003;
    wire new_Jinkela_wire_13103;
    wire new_Jinkela_wire_14660;
    wire new_Jinkela_wire_17703;
    wire new_Jinkela_wire_8519;
    wire new_Jinkela_wire_13840;
    wire new_Jinkela_wire_10260;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_18042;
    wire new_Jinkela_wire_12354;
    wire new_Jinkela_wire_17377;
    wire new_Jinkela_wire_4821;
    wire new_Jinkela_wire_17113;
    wire new_Jinkela_wire_18469;
    wire new_Jinkela_wire_14155;
    wire new_Jinkela_wire_3263;
    wire new_Jinkela_wire_19501;
    wire new_Jinkela_wire_16027;
    wire new_Jinkela_wire_9403;
    wire new_Jinkela_wire_20565;
    wire new_Jinkela_wire_7952;
    wire new_Jinkela_wire_18953;
    wire new_Jinkela_wire_13159;
    wire new_Jinkela_wire_4360;
    wire new_Jinkela_wire_20229;
    wire new_Jinkela_wire_17240;
    wire new_Jinkela_wire_4328;
    wire new_Jinkela_wire_19962;
    wire new_Jinkela_wire_16994;
    wire new_Jinkela_wire_5526;
    wire new_Jinkela_wire_16125;
    wire new_Jinkela_wire_17237;
    wire new_Jinkela_wire_5703;
    wire _1239_;
    wire new_Jinkela_wire_17492;
    wire new_Jinkela_wire_19126;
    wire new_Jinkela_wire_18123;
    wire new_Jinkela_wire_10389;
    wire new_Jinkela_wire_8207;
    wire new_Jinkela_wire_5813;
    wire new_Jinkela_wire_4116;
    wire new_Jinkela_wire_3049;
    wire new_Jinkela_wire_6203;
    wire new_Jinkela_wire_17454;
    wire new_Jinkela_wire_12024;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_3419;
    wire new_Jinkela_wire_13382;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_15610;
    wire _1240_;
    wire new_Jinkela_wire_20069;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_16203;
    wire new_Jinkela_wire_2569;
    wire new_Jinkela_wire_17840;
    wire new_Jinkela_wire_6173;
    wire new_Jinkela_wire_9415;
    wire new_Jinkela_wire_8842;
    wire _1482_;
    wire new_Jinkela_wire_9998;
    wire new_Jinkela_wire_10172;
    wire new_Jinkela_wire_2340;
    wire _1530_;
    wire new_Jinkela_wire_3052;
    wire new_Jinkela_wire_20357;
    wire _0976_;
    wire new_Jinkela_wire_8474;
    wire new_Jinkela_wire_3822;
    wire new_Jinkela_wire_5312;
    wire new_Jinkela_wire_21254;
    wire new_Jinkela_wire_10905;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_13290;
    wire new_Jinkela_wire_12274;
    wire new_Jinkela_wire_9176;
    wire _0214_;
    wire new_Jinkela_wire_18517;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_14925;
    wire new_Jinkela_wire_8094;
    wire new_Jinkela_wire_7097;
    wire new_Jinkela_wire_6619;
    wire _1544_;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_11493;
    wire new_Jinkela_wire_10078;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_18858;
    wire new_Jinkela_wire_19717;
    wire _1176_;
    wire _0406_;
    wire new_Jinkela_wire_10282;
    wire new_Jinkela_wire_12986;
    wire new_Jinkela_wire_12323;
    wire new_Jinkela_wire_20401;
    wire new_Jinkela_wire_11129;
    wire new_Jinkela_wire_15876;
    wire new_Jinkela_wire_5355;
    wire new_Jinkela_wire_11481;
    wire new_Jinkela_wire_14936;
    wire new_Jinkela_wire_12149;
    wire _0979_;
    wire new_Jinkela_wire_17593;
    wire new_Jinkela_wire_9247;
    wire new_Jinkela_wire_9587;
    wire _1389_;
    wire _1086_;
    wire new_Jinkela_wire_7359;
    wire new_Jinkela_wire_6325;
    wire new_Jinkela_wire_14295;
    wire new_Jinkela_wire_19471;
    wire new_Jinkela_wire_17149;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_2527;
    wire new_Jinkela_wire_20389;
    wire new_Jinkela_wire_17099;
    wire new_Jinkela_wire_13109;
    wire new_Jinkela_wire_6672;
    wire _0763_;
    wire new_Jinkela_wire_10247;
    wire new_Jinkela_wire_17942;
    wire new_Jinkela_wire_14450;
    wire new_Jinkela_wire_4631;
    wire new_Jinkela_wire_20898;
    wire new_Jinkela_wire_12417;
    wire new_Jinkela_wire_18507;
    wire new_Jinkela_wire_5138;
    wire new_Jinkela_wire_13225;
    wire new_Jinkela_wire_6019;
    wire new_Jinkela_wire_5482;
    wire new_Jinkela_wire_4654;
    wire new_Jinkela_wire_11206;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_5010;
    wire new_Jinkela_wire_13168;
    wire new_Jinkela_wire_2300;
    wire new_Jinkela_wire_2004;
    wire new_Jinkela_wire_14405;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_4303;
    wire new_Jinkela_wire_3852;
    wire new_Jinkela_wire_5742;
    wire new_Jinkela_wire_14011;
    wire new_Jinkela_wire_15691;
    wire new_Jinkela_wire_14046;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_15488;
    wire _0564_;
    wire new_Jinkela_wire_4785;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_7499;
    wire new_Jinkela_wire_7345;
    wire new_Jinkela_wire_5948;
    wire new_Jinkela_wire_14603;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_9883;
    wire new_Jinkela_wire_17156;
    wire new_Jinkela_wire_13048;
    wire new_Jinkela_wire_16724;
    wire new_Jinkela_wire_3750;
    wire new_Jinkela_wire_9733;
    wire new_Jinkela_wire_15300;
    wire new_Jinkela_wire_3385;
    wire new_Jinkela_wire_4676;
    wire new_Jinkela_wire_6932;
    wire new_Jinkela_wire_6393;
    wire new_Jinkela_wire_10131;
    wire new_Jinkela_wire_6187;
    wire new_Jinkela_wire_15339;
    wire new_Jinkela_wire_3246;
    wire new_Jinkela_wire_2863;
    wire new_Jinkela_wire_15646;
    wire new_Jinkela_wire_9757;
    wire new_Jinkela_wire_4119;
    wire new_Jinkela_wire_8871;
    wire new_Jinkela_wire_10817;
    wire new_Jinkela_wire_7346;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_20245;
    wire new_Jinkela_wire_5556;
    wire new_Jinkela_wire_4776;
    wire new_Jinkela_wire_1893;
    wire new_Jinkela_wire_10059;
    wire new_Jinkela_wire_15460;
    wire new_Jinkela_wire_13463;
    wire new_Jinkela_wire_8385;
    wire new_Jinkela_wire_16522;
    wire new_Jinkela_wire_14710;
    wire _1398_;
    wire new_Jinkela_wire_17301;
    wire new_Jinkela_wire_15865;
    wire new_Jinkela_wire_1742;
    wire new_Jinkela_wire_13948;
    wire new_Jinkela_wire_19777;
    wire new_Jinkela_wire_19865;
    wire new_Jinkela_wire_9843;
    wire new_Jinkela_wire_21332;
    wire new_Jinkela_wire_6948;
    wire new_Jinkela_wire_21320;
    wire new_Jinkela_wire_17364;
    wire new_Jinkela_wire_15735;
    wire new_Jinkela_wire_6020;
    wire new_Jinkela_wire_16730;
    wire new_Jinkela_wire_5079;
    wire new_Jinkela_wire_6371;
    wire new_Jinkela_wire_5043;
    wire new_Jinkela_wire_16757;
    wire new_Jinkela_wire_12521;
    wire new_Jinkela_wire_19611;
    wire new_Jinkela_wire_18175;
    wire new_Jinkela_wire_16065;
    wire new_Jinkela_wire_20799;
    wire new_Jinkela_wire_5200;
    wire new_Jinkela_wire_2521;
    wire new_Jinkela_wire_9009;
    wire new_Jinkela_wire_2456;
    wire new_Jinkela_wire_8487;
    wire new_Jinkela_wire_11869;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_7470;
    wire new_Jinkela_wire_17101;
    wire new_Jinkela_wire_3040;
    wire new_Jinkela_wire_8462;
    wire new_Jinkela_wire_4687;
    wire _0700_;
    wire new_Jinkela_wire_12547;
    wire new_Jinkela_wire_19073;
    wire new_Jinkela_wire_16474;
    wire new_Jinkela_wire_12993;
    wire new_Jinkela_wire_7996;
    wire new_Jinkela_wire_20904;
    wire new_Jinkela_wire_1110;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_20685;
    wire new_Jinkela_wire_17537;
    wire new_Jinkela_wire_11907;
    wire new_Jinkela_wire_14820;
    wire new_Jinkela_wire_20714;
    wire new_Jinkela_wire_11165;
    wire _0463_;
    wire new_Jinkela_wire_17257;
    wire new_Jinkela_wire_19005;
    wire new_Jinkela_wire_13300;
    wire new_Jinkela_wire_5267;
    wire new_Jinkela_wire_12957;
    wire new_Jinkela_wire_4032;
    wire new_Jinkela_wire_12430;
    wire new_Jinkela_wire_1436;
    wire _1261_;
    wire new_Jinkela_wire_14335;
    wire new_Jinkela_wire_20973;
    wire new_Jinkela_wire_3234;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_11543;
    wire new_Jinkela_wire_20437;
    wire new_Jinkela_wire_7220;
    wire _0863_;
    wire new_Jinkela_wire_3099;
    wire new_Jinkela_wire_13778;
    wire new_Jinkela_wire_5656;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_14550;
    wire new_Jinkela_wire_18500;
    wire new_Jinkela_wire_9986;
    wire new_Jinkela_wire_1429;
    wire _0891_;
    wire new_Jinkela_wire_16918;
    wire new_Jinkela_wire_12616;
    wire new_Jinkela_wire_4285;
    wire new_Jinkela_wire_9927;
    wire new_Jinkela_wire_18010;
    wire new_Jinkela_wire_6127;
    wire new_Jinkela_wire_6163;
    wire new_Jinkela_wire_5938;
    wire new_Jinkela_wire_4721;
    wire new_Jinkela_wire_6341;
    wire new_Jinkela_wire_18267;
    wire new_Jinkela_wire_13239;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_4123;
    wire new_Jinkela_wire_13523;
    wire new_Jinkela_wire_3340;
    wire new_Jinkela_wire_10106;
    wire new_Jinkela_wire_20812;
    wire new_Jinkela_wire_14495;
    wire new_Jinkela_wire_9242;
    wire new_Jinkela_wire_9346;
    wire new_Jinkela_wire_8142;
    wire new_Jinkela_wire_18686;
    wire new_Jinkela_wire_9104;
    wire new_Jinkela_wire_15774;
    wire new_Jinkela_wire_1514;
    wire new_net_3932;
    wire new_Jinkela_wire_18823;
    wire new_Jinkela_wire_8936;
    wire new_Jinkela_wire_17180;
    wire new_Jinkela_wire_3214;
    wire new_Jinkela_wire_12688;
    wire new_Jinkela_wire_14517;
    wire new_Jinkela_wire_15917;
    wire new_Jinkela_wire_14192;
    wire new_Jinkela_wire_6160;
    wire new_Jinkela_wire_12327;
    wire new_Jinkela_wire_15353;
    wire new_Jinkela_wire_21027;
    wire new_Jinkela_wire_3039;
    wire _1199_;
    wire new_Jinkela_wire_19766;
    wire _1140_;
    wire new_Jinkela_wire_20056;
    wire _1166_;
    wire new_Jinkela_wire_2875;
    wire new_Jinkela_wire_17450;
    wire new_Jinkela_wire_3633;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_2941;
    wire new_Jinkela_wire_15773;
    wire new_Jinkela_wire_5443;
    wire new_Jinkela_wire_17708;
    wire new_Jinkela_wire_10847;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_4451;
    wire new_Jinkela_wire_6637;
    wire new_Jinkela_wire_15164;
    wire _0271_;
    wire new_Jinkela_wire_7939;
    wire new_Jinkela_wire_21142;
    wire new_Jinkela_wire_7783;
    wire new_Jinkela_wire_14416;
    wire _0018_;
    wire new_Jinkela_wire_17090;
    wire new_Jinkela_wire_13958;
    wire _0373_;
    wire _0984_;
    wire new_Jinkela_wire_11185;
    wire new_Jinkela_wire_11890;
    wire new_Jinkela_wire_2178;
    wire new_Jinkela_wire_13384;
    wire new_Jinkela_wire_17916;
    wire new_Jinkela_wire_18776;
    wire new_Jinkela_wire_15967;
    wire new_Jinkela_wire_12585;
    wire new_Jinkela_wire_7015;
    wire new_Jinkela_wire_9949;
    wire new_Jinkela_wire_2386;
    wire new_Jinkela_wire_17455;
    wire new_Jinkela_wire_13606;
    wire new_Jinkela_wire_13531;
    wire new_Jinkela_wire_5964;
    wire new_Jinkela_wire_9408;
    wire new_Jinkela_wire_9779;
    wire new_Jinkela_wire_9412;
    wire new_Jinkela_wire_2282;
    wire new_Jinkela_wire_8128;
    wire new_Jinkela_wire_15459;
    wire new_Jinkela_wire_12892;
    wire new_Jinkela_wire_20000;
    wire new_Jinkela_wire_7375;
    wire _1817_;
    wire new_Jinkela_wire_7954;
    wire _0792_;
    wire new_Jinkela_wire_3576;
    wire new_net_3940;
    wire new_Jinkela_wire_9967;
    wire new_Jinkela_wire_15254;
    wire new_Jinkela_wire_16231;
    wire new_Jinkela_wire_15429;
    wire new_Jinkela_wire_7851;
    wire _1747_;
    wire new_Jinkela_wire_19990;
    wire _0507_;
    wire new_Jinkela_wire_9205;
    wire new_Jinkela_wire_17176;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_8890;
    wire new_Jinkela_wire_4750;
    wire new_Jinkela_wire_10014;
    wire new_Jinkela_wire_12516;
    wire new_Jinkela_wire_20694;
    wire new_Jinkela_wire_11727;
    wire _1636_;
    wire new_Jinkela_wire_9648;
    wire new_Jinkela_wire_17321;
    wire new_Jinkela_wire_15584;
    wire new_Jinkela_wire_5247;
    wire new_Jinkela_wire_11182;
    wire _1678_;
    wire new_Jinkela_wire_16624;
    wire new_Jinkela_wire_18088;
    wire new_Jinkela_wire_7450;
    wire _0136_;
    wire new_Jinkela_wire_7545;
    wire new_Jinkela_wire_19765;
    wire new_Jinkela_wire_3656;
    wire new_Jinkela_wire_17891;
    wire new_Jinkela_wire_9862;
    wire new_Jinkela_wire_12485;
    wire new_Jinkela_wire_10015;
    wire new_Jinkela_wire_1036;
    wire new_Jinkela_wire_8250;
    wire new_Jinkela_wire_4446;
    wire new_Jinkela_wire_4106;
    wire new_Jinkela_wire_3830;
    wire _0248_;
    wire new_Jinkela_wire_16895;
    wire new_Jinkela_wire_16962;
    wire new_Jinkela_wire_3493;
    wire new_Jinkela_wire_8228;
    wire new_Jinkela_wire_9596;
    wire new_Jinkela_wire_10470;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_7403;
    wire new_Jinkela_wire_8132;
    wire new_Jinkela_wire_18756;
    wire new_Jinkela_wire_6292;
    wire new_Jinkela_wire_8787;
    wire new_Jinkela_wire_8537;
    wire new_Jinkela_wire_3556;
    wire _1510_;
    wire new_Jinkela_wire_6673;
    wire new_Jinkela_wire_14958;
    wire new_Jinkela_wire_17389;
    wire new_Jinkela_wire_16092;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_8712;
    wire new_Jinkela_wire_5726;
    wire new_Jinkela_wire_15822;
    wire new_Jinkela_wire_3561;
    wire new_Jinkela_wire_7614;
    wire new_Jinkela_wire_7256;
    wire new_Jinkela_wire_5349;
    wire new_Jinkela_wire_14835;
    wire new_Jinkela_wire_2865;
    wire new_Jinkela_wire_2647;
    wire new_Jinkela_wire_18939;
    wire new_Jinkela_wire_19831;
    wire new_Jinkela_wire_16168;
    wire new_Jinkela_wire_10932;
    wire new_Jinkela_wire_12965;
    wire new_Jinkela_wire_14181;
    wire _0401_;
    wire new_Jinkela_wire_7170;
    wire new_Jinkela_wire_3152;
    wire new_Jinkela_wire_19066;
    wire new_Jinkela_wire_8497;
    wire _1273_;
    wire new_Jinkela_wire_20957;
    wire new_Jinkela_wire_15271;
    wire new_Jinkela_wire_8174;
    wire new_Jinkela_wire_15156;
    wire new_Jinkela_wire_9767;
    wire new_Jinkela_wire_18141;
    wire new_Jinkela_wire_17071;
    wire new_Jinkela_wire_8370;
    wire new_Jinkela_wire_8704;
    wire _1748_;
    wire new_Jinkela_wire_10113;
    wire new_Jinkela_wire_18551;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_8103;
    wire new_Jinkela_wire_9654;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_10453;
    wire _0147_;
    wire new_Jinkela_wire_20131;
    wire new_Jinkela_wire_6550;
    wire new_Jinkela_wire_19311;
    wire _0219_;
    wire new_Jinkela_wire_8880;
    wire new_Jinkela_wire_8369;
    wire new_net_3938;
    wire new_Jinkela_wire_14256;
    wire new_Jinkela_wire_19754;
    wire new_Jinkela_wire_20668;
    wire _1531_;
    wire new_Jinkela_wire_14162;
    wire new_Jinkela_wire_13732;
    wire new_Jinkela_wire_14672;
    wire new_Jinkela_wire_19313;
    wire new_Jinkela_wire_12595;
    wire new_Jinkela_wire_12691;
    wire new_Jinkela_wire_6492;
    wire new_Jinkela_wire_9563;
    wire new_Jinkela_wire_5201;
    wire new_Jinkela_wire_11189;
    wire new_Jinkela_wire_6720;
    wire new_Jinkela_wire_9340;
    wire new_Jinkela_wire_3583;
    wire new_Jinkela_wire_12267;
    wire new_Jinkela_wire_19645;
    wire new_Jinkela_wire_16074;
    wire new_Jinkela_wire_13266;
    wire new_Jinkela_wire_15856;
    wire new_Jinkela_wire_11207;
    wire new_Jinkela_wire_9190;
    wire new_Jinkela_wire_5547;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_7252;
    wire new_Jinkela_wire_10475;
    wire new_Jinkela_wire_7948;
    wire new_Jinkela_wire_18850;
    wire new_Jinkela_wire_19340;
    wire new_Jinkela_wire_5084;
    wire new_Jinkela_wire_15642;
    wire new_Jinkela_wire_10789;
    wire new_Jinkela_wire_7940;
    wire new_Jinkela_wire_3148;
    wire new_Jinkela_wire_19286;
    wire new_Jinkela_wire_5403;
    wire new_Jinkela_wire_5143;
    wire new_Jinkela_wire_9351;
    wire new_Jinkela_wire_11996;
    wire new_Jinkela_wire_13110;
    wire new_Jinkela_wire_10710;
    wire _1783_;
    wire new_Jinkela_wire_2035;
    wire new_Jinkela_wire_9749;
    wire _0044_;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_12895;
    wire new_Jinkela_wire_9722;
    wire new_Jinkela_wire_11287;
    wire new_Jinkela_wire_10583;
    wire new_Jinkela_wire_2200;
    wire new_Jinkela_wire_14795;
    wire new_Jinkela_wire_13846;
    wire new_Jinkela_wire_8421;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_21103;
    wire new_Jinkela_wire_4302;
    wire new_Jinkela_wire_14378;
    wire new_Jinkela_wire_5558;
    wire new_Jinkela_wire_13251;
    wire new_Jinkela_wire_15641;
    wire new_Jinkela_wire_2137;
    wire new_Jinkela_wire_14120;
    wire new_Jinkela_wire_1040;
    wire new_Jinkela_wire_19753;
    wire new_Jinkela_wire_7484;
    wire new_Jinkela_wire_19525;
    wire new_Jinkela_wire_12614;
    wire new_Jinkela_wire_17877;
    wire new_Jinkela_wire_15225;
    wire new_Jinkela_wire_13627;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_9172;
    wire new_Jinkela_wire_14110;
    wire new_Jinkela_wire_4709;
    wire new_Jinkela_wire_3764;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_2451;
    wire new_Jinkela_wire_13261;
    wire new_Jinkela_wire_20158;
    wire new_Jinkela_wire_3432;
    wire new_Jinkela_wire_11846;
    wire new_Jinkela_wire_19821;
    wire new_Jinkela_wire_11300;
    wire _0982_;
    wire new_Jinkela_wire_18692;
    wire new_Jinkela_wire_3397;
    wire new_Jinkela_wire_17745;
    wire _0736_;
    wire new_Jinkela_wire_16702;
    wire new_Jinkela_wire_20280;
    wire new_Jinkela_wire_14913;
    wire new_Jinkela_wire_8937;
    wire new_Jinkela_wire_16364;
    wire new_Jinkela_wire_18413;
    wire new_Jinkela_wire_6810;
    wire new_Jinkela_wire_16477;
    wire new_Jinkela_wire_7201;
    wire new_Jinkela_wire_2874;
    wire new_Jinkela_wire_19517;
    wire new_Jinkela_wire_18005;
    wire new_Jinkela_wire_20839;
    wire new_Jinkela_wire_20563;
    wire new_Jinkela_wire_17254;
    wire new_Jinkela_wire_14246;
    wire new_Jinkela_wire_15984;
    wire new_Jinkela_wire_10142;
    wire new_Jinkela_wire_7844;
    wire new_Jinkela_wire_20109;
    wire new_Jinkela_wire_6569;
    wire new_Jinkela_wire_12446;
    wire new_Jinkela_wire_4226;
    wire new_Jinkela_wire_7119;
    wire new_Jinkela_wire_4292;
    wire new_Jinkela_wire_14153;
    wire new_Jinkela_wire_2541;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_6759;
    wire new_Jinkela_wire_11725;
    wire new_Jinkela_wire_5760;
    wire new_Jinkela_wire_19832;
    wire new_Jinkela_wire_16635;
    wire new_Jinkela_wire_19151;
    wire _1286_;
    wire new_Jinkela_wire_6164;
    wire new_Jinkela_wire_9143;
    wire _1775_;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_5212;
    wire new_Jinkela_wire_2712;
    wire _1664_;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_9214;
    wire new_Jinkela_wire_16580;
    wire _1598_;
    wire new_Jinkela_wire_6093;
    wire new_Jinkela_wire_13138;
    wire new_Jinkela_wire_11063;
    wire new_Jinkela_wire_17054;
    wire new_Jinkela_wire_18080;
    wire new_net_3972;
    wire new_Jinkela_wire_15487;
    wire new_Jinkela_wire_5649;
    wire _0116_;
    wire new_Jinkela_wire_18734;
    wire new_Jinkela_wire_12528;
    wire new_Jinkela_wire_16601;
    wire new_Jinkela_wire_20233;
    wire new_Jinkela_wire_8445;
    wire new_Jinkela_wire_14225;
    wire new_Jinkela_wire_2084;
    wire new_Jinkela_wire_19861;
    wire new_Jinkela_wire_3825;
    wire new_Jinkela_wire_5887;
    wire new_Jinkela_wire_11643;
    wire new_Jinkela_wire_2154;
    wire new_Jinkela_wire_6246;
    wire new_Jinkela_wire_11724;
    wire new_Jinkela_wire_8319;
    wire new_Jinkela_wire_12342;
    wire new_Jinkela_wire_19421;
    wire new_Jinkela_wire_5576;
    wire new_Jinkela_wire_16823;
    wire new_Jinkela_wire_12812;
    wire new_Jinkela_wire_17961;
    wire new_Jinkela_wire_6234;
    wire new_Jinkela_wire_4907;
    wire new_Jinkela_wire_2293;
    wire new_Jinkela_wire_9282;
    wire new_Jinkela_wire_12467;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_9450;
    wire new_Jinkela_wire_11552;
    wire new_Jinkela_wire_7733;
    wire new_Jinkela_wire_4157;
    wire new_Jinkela_wire_18808;
    wire new_Jinkela_wire_12636;
    wire new_Jinkela_wire_20860;
    wire new_Jinkela_wire_17141;
    wire new_Jinkela_wire_7519;
    wire new_Jinkela_wire_1698;
    wire new_Jinkela_wire_18198;
    wire new_Jinkela_wire_20700;
    wire new_Jinkela_wire_7444;
    wire new_Jinkela_wire_17138;
    wire new_Jinkela_wire_10011;
    wire new_Jinkela_wire_1691;
    wire new_Jinkela_wire_10417;
    wire new_net_3930;
    wire new_Jinkela_wire_9701;
    wire new_Jinkela_wire_19925;
    wire _1143_;
    wire new_Jinkela_wire_16202;
    wire new_Jinkela_wire_2652;
    wire new_Jinkela_wire_2103;
    wire new_Jinkela_wire_10775;
    wire _0850_;
    wire new_Jinkela_wire_18596;
    wire new_Jinkela_wire_19612;
    wire new_Jinkela_wire_9374;
    wire new_Jinkela_wire_7422;
    wire new_Jinkela_wire_3430;
    wire new_Jinkela_wire_4061;
    wire new_Jinkela_wire_19687;
    wire _1196_;
    wire new_Jinkela_wire_13333;
    wire new_Jinkela_wire_12279;
    wire new_Jinkela_wire_16217;
    wire new_Jinkela_wire_2148;
    wire new_Jinkela_wire_14498;
    wire new_Jinkela_wire_4013;
    wire new_Jinkela_wire_6349;
    wire new_Jinkela_wire_4077;
    wire new_Jinkela_wire_12641;
    wire new_Jinkela_wire_4874;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_18046;
    wire _1622_;
    wire new_Jinkela_wire_12481;
    wire new_Jinkela_wire_13461;
    wire new_Jinkela_wire_5851;
    wire new_Jinkela_wire_17387;
    wire new_Jinkela_wire_10252;
    wire new_Jinkela_wire_17573;
    wire _0834_;
    wire new_Jinkela_wire_20236;
    wire new_Jinkela_wire_3660;
    wire new_Jinkela_wire_14083;
    wire new_Jinkela_wire_5126;
    wire new_Jinkela_wire_4489;
    wire new_Jinkela_wire_8468;
    wire _1509_;
    wire new_Jinkela_wire_14076;
    wire new_Jinkela_wire_12862;
    wire new_Jinkela_wire_15332;
    wire new_Jinkela_wire_14117;
    wire new_Jinkela_wire_21076;
    wire _1046_;
    wire new_Jinkela_wire_7388;
    wire new_Jinkela_wire_17478;
    wire new_Jinkela_wire_16991;
    wire new_Jinkela_wire_20801;
    wire new_Jinkela_wire_21268;
    wire new_Jinkela_wire_4493;
    wire new_Jinkela_wire_17755;
    wire new_Jinkela_wire_3285;
    wire new_Jinkela_wire_13806;
    wire new_Jinkela_wire_13480;
    wire new_Jinkela_wire_13761;
    wire new_Jinkela_wire_5580;
    wire new_Jinkela_wire_13292;
    wire new_Jinkela_wire_15455;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_7847;
    wire new_Jinkela_wire_15014;
    wire new_Jinkela_wire_13388;
    wire _1570_;
    wire new_Jinkela_wire_2561;
    wire new_Jinkela_wire_5860;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_17606;
    wire new_Jinkela_wire_9834;
    wire new_Jinkela_wire_7853;
    wire new_Jinkela_wire_5314;
    wire new_Jinkela_wire_5412;
    wire new_Jinkela_wire_6011;
    wire new_Jinkela_wire_7894;
    wire _0162_;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_9149;
    wire _0126_;
    wire new_Jinkela_wire_3281;
    wire new_Jinkela_wire_17887;
    wire new_Jinkela_wire_16003;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_17560;
    wire new_Jinkela_wire_20702;
    wire new_Jinkela_wire_15450;
    wire new_Jinkela_wire_18660;
    wire new_Jinkela_wire_11749;
    wire _1065_;
    wire new_Jinkela_wire_4005;
    wire new_Jinkela_wire_12226;
    wire new_Jinkela_wire_5237;
    wire new_Jinkela_wire_11029;
    wire new_Jinkela_wire_6331;
    wire new_Jinkela_wire_9187;
    wire new_Jinkela_wire_3222;
    wire new_Jinkela_wire_14279;
    wire new_Jinkela_wire_8185;
    wire new_Jinkela_wire_2082;
    wire new_Jinkela_wire_14475;
    wire new_Jinkela_wire_8177;
    wire new_Jinkela_wire_20950;
    wire new_Jinkela_wire_13629;
    wire new_Jinkela_wire_5653;
    wire new_Jinkela_wire_8382;
    wire _0365_;
    wire _1592_;
    wire new_Jinkela_wire_3757;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_13817;
    wire new_Jinkela_wire_15352;
    wire new_Jinkela_wire_16788;
    wire new_Jinkela_wire_3973;
    wire new_Jinkela_wire_12277;
    wire new_Jinkela_wire_18314;
    wire new_Jinkela_wire_7524;
    wire new_Jinkela_wire_20367;
    wire _0167_;
    wire new_Jinkela_wire_19665;
    wire _0841_;
    wire new_Jinkela_wire_4964;
    wire new_Jinkela_wire_5219;
    wire new_Jinkela_wire_14644;
    wire new_Jinkela_wire_6411;
    wire new_Jinkela_wire_15495;
    wire new_Jinkela_wire_6551;
    wire new_Jinkela_wire_10755;
    wire new_Jinkela_wire_6293;
    wire new_Jinkela_wire_16193;
    wire new_Jinkela_wire_20935;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_2512;
    wire new_Jinkela_wire_16545;
    wire new_Jinkela_wire_8909;
    wire new_Jinkela_wire_2266;
    wire new_Jinkela_wire_16448;
    wire new_Jinkela_wire_15812;
    wire new_Jinkela_wire_21113;
    wire _1105_;
    wire _0183_;
    wire new_Jinkela_wire_8033;
    wire new_Jinkela_wire_16213;
    wire new_Jinkela_wire_10882;
    wire new_Jinkela_wire_13162;
    wire new_Jinkela_wire_9610;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_19949;
    wire new_Jinkela_wire_3756;
    wire new_Jinkela_wire_9691;
    wire new_Jinkela_wire_17984;
    wire _0512_;
    wire new_Jinkela_wire_10731;
    wire _0325_;
    wire new_Jinkela_wire_5006;
    wire new_Jinkela_wire_13763;
    wire new_Jinkela_wire_5152;
    wire new_Jinkela_wire_4347;
    wire new_Jinkela_wire_20541;
    wire new_Jinkela_wire_11614;
    wire new_Jinkela_wire_15358;
    wire new_Jinkela_wire_3814;
    wire new_Jinkela_wire_12900;
    wire new_Jinkela_wire_17183;
    wire new_Jinkela_wire_13434;
    wire new_Jinkela_wire_16798;
    wire new_Jinkela_wire_6326;
    wire new_Jinkela_wire_15726;
    wire new_Jinkela_wire_8384;
    wire _1299_;
    wire new_Jinkela_wire_4925;
    wire new_Jinkela_wire_16131;
    wire new_Jinkela_wire_11428;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_20761;
    wire new_Jinkela_wire_12637;
    wire new_Jinkela_wire_8425;
    wire new_Jinkela_wire_11291;
    wire new_Jinkela_wire_9369;
    wire new_Jinkela_wire_5804;
    wire new_Jinkela_wire_10484;
    wire new_Jinkela_wire_11549;
    wire new_Jinkela_wire_6994;
    wire new_Jinkela_wire_17718;
    wire new_Jinkela_wire_21182;
    wire new_Jinkela_wire_10536;
    wire new_Jinkela_wire_7696;
    wire new_Jinkela_wire_2894;
    wire new_Jinkela_wire_19329;
    wire new_Jinkela_wire_16139;
    wire new_Jinkela_wire_19529;
    wire new_Jinkela_wire_5075;
    wire new_Jinkela_wire_3934;
    wire new_Jinkela_wire_4002;
    wire new_Jinkela_wire_13246;
    wire new_Jinkela_wire_13146;
    wire new_Jinkela_wire_12543;
    wire new_Jinkela_wire_14131;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_16309;
    wire new_Jinkela_wire_2378;
    wire new_Jinkela_wire_12308;
    wire new_Jinkela_wire_5174;
    wire new_Jinkela_wire_7692;
    wire new_Jinkela_wire_20170;
    wire _1385_;
    wire new_Jinkela_wire_12723;
    wire new_Jinkela_wire_7114;
    wire new_Jinkela_wire_4400;
    wire new_Jinkela_wire_14716;
    wire new_Jinkela_wire_2578;
    wire new_Jinkela_wire_14768;
    wire new_Jinkela_wire_14129;
    wire new_Jinkela_wire_7740;
    wire new_Jinkela_wire_5907;
    wire _0113_;
    wire _1749_;
    wire new_Jinkela_wire_18024;
    wire new_Jinkela_wire_12062;
    wire new_Jinkela_wire_10683;
    wire new_Jinkela_wire_10970;
    wire new_Jinkela_wire_7746;
    wire new_Jinkela_wire_1800;
    wire new_Jinkela_wire_20383;
    wire new_Jinkela_wire_3956;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_15785;
    wire new_Jinkela_wire_4247;
    wire _0972_;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_14024;
    wire new_Jinkela_wire_15649;
    wire new_net_3970;
    wire _1361_;
    wire new_Jinkela_wire_5545;
    wire new_Jinkela_wire_16633;
    wire _0431_;
    wire new_Jinkela_wire_20561;
    wire new_Jinkela_wire_17431;
    wire new_Jinkela_wire_3412;
    wire new_Jinkela_wire_6718;
    wire new_Jinkela_wire_8116;
    wire new_Jinkela_wire_16708;
    wire new_Jinkela_wire_3684;
    wire new_Jinkela_wire_13122;
    wire new_Jinkela_wire_14185;
    wire new_Jinkela_wire_10061;
    wire new_Jinkela_wire_4475;
    wire new_Jinkela_wire_18444;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_12846;
    wire new_Jinkela_wire_2630;
    wire new_Jinkela_wire_18247;
    wire new_Jinkela_wire_16672;
    wire new_Jinkela_wire_10769;
    wire new_Jinkela_wire_9084;
    wire new_Jinkela_wire_10790;
    wire _1405_;
    wire new_Jinkela_wire_17962;
    wire new_Jinkela_wire_20036;
    wire new_Jinkela_wire_17611;
    wire new_Jinkela_wire_11950;
    wire new_Jinkela_wire_20468;
    wire new_Jinkela_wire_10020;
    wire new_Jinkela_wire_11731;
    wire new_Jinkela_wire_7126;
    wire new_Jinkela_wire_6639;
    wire new_Jinkela_wire_18483;
    wire new_Jinkela_wire_21165;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_19676;
    wire new_Jinkela_wire_10757;
    wire new_Jinkela_wire_3510;
    wire new_Jinkela_wire_14688;
    wire new_Jinkela_wire_9799;
    wire new_Jinkela_wire_8630;
    wire new_Jinkela_wire_19007;
    wire new_Jinkela_wire_9089;
    wire new_Jinkela_wire_7250;
    wire new_Jinkela_wire_10413;
    wire new_Jinkela_wire_18769;
    wire new_Jinkela_wire_12663;
    wire new_Jinkela_wire_10108;
    wire new_Jinkela_wire_3496;
    wire new_Jinkela_wire_6439;
    wire new_Jinkela_wire_13343;
    wire new_Jinkela_wire_8840;
    wire new_Jinkela_wire_12652;
    wire new_Jinkela_wire_5714;
    wire new_Jinkela_wire_9285;
    wire new_Jinkela_wire_9882;
    wire new_Jinkela_wire_10259;
    wire new_Jinkela_wire_8558;
    wire new_Jinkela_wire_18228;
    wire new_Jinkela_wire_6688;
    wire new_Jinkela_wire_10593;
    wire new_Jinkela_wire_5000;
    wire new_Jinkela_wire_6077;
    wire new_Jinkela_wire_15769;
    wire new_Jinkela_wire_8685;
    wire new_Jinkela_wire_8007;
    wire new_Jinkela_wire_2706;
    wire new_Jinkela_wire_20246;
    wire _0883_;
    wire new_Jinkela_wire_2687;
    wire new_Jinkela_wire_11299;
    wire new_Jinkela_wire_11174;
    wire new_Jinkela_wire_14519;
    wire new_Jinkela_wire_10869;
    wire new_Jinkela_wire_20789;
    wire new_Jinkela_wire_17583;
    wire new_Jinkela_wire_7206;
    wire new_Jinkela_wire_16971;
    wire new_Jinkela_wire_7160;
    wire new_Jinkela_wire_18399;
    wire new_Jinkela_wire_19499;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_14987;
    wire new_Jinkela_wire_17975;
    wire new_Jinkela_wire_6884;
    wire new_Jinkela_wire_14136;
    wire new_Jinkela_wire_13650;
    wire new_Jinkela_wire_20952;
    wire new_Jinkela_wire_15121;
    wire new_Jinkela_wire_2755;
    wire new_Jinkela_wire_3092;
    wire new_Jinkela_wire_18173;
    wire new_Jinkela_wire_17483;
    wire new_Jinkela_wire_6059;
    wire new_Jinkela_wire_5016;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_4087;
    wire new_Jinkela_wire_4095;
    wire new_Jinkela_wire_18391;
    wire new_Jinkela_wire_5790;
    wire _0633_;
    wire new_Jinkela_wire_3243;
    wire new_Jinkela_wire_6263;
    wire new_Jinkela_wire_16963;
    wire new_Jinkela_wire_4434;
    wire new_Jinkela_wire_12388;
    wire new_Jinkela_wire_10909;
    wire new_Jinkela_wire_15776;
    wire new_Jinkela_wire_7636;
    wire new_Jinkela_wire_12462;
    wire new_Jinkela_wire_12903;
    wire new_Jinkela_wire_12010;
    wire _0613_;
    wire new_Jinkela_wire_18452;
    wire new_Jinkela_wire_12538;
    wire new_Jinkela_wire_9397;
    wire new_Jinkela_wire_9791;
    wire new_Jinkela_wire_12329;
    wire new_Jinkela_wire_12078;
    wire new_Jinkela_wire_17049;
    wire new_Jinkela_wire_12330;
    wire new_Jinkela_wire_2217;
    wire new_Jinkela_wire_2143;
    wire new_Jinkela_wire_14041;
    wire new_Jinkela_wire_11709;
    wire new_Jinkela_wire_4305;
    wire _1464_;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_18725;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_10141;
    wire new_Jinkela_wire_9948;
    wire new_Jinkela_wire_20969;
    wire new_Jinkela_wire_13070;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_13598;
    wire new_Jinkela_wire_4102;
    wire _0137_;
    wire new_Jinkela_wire_17042;
    wire new_Jinkela_wire_12377;
    wire new_Jinkela_wire_13782;
    wire new_Jinkela_wire_7402;
    wire new_Jinkela_wire_13536;
    wire new_Jinkela_wire_12834;
    wire new_Jinkela_wire_18671;
    wire new_Jinkela_wire_10124;
    wire new_Jinkela_wire_12724;
    wire new_Jinkela_wire_18807;
    wire new_Jinkela_wire_16905;
    wire new_Jinkela_wire_12060;
    wire new_Jinkela_wire_3353;
    wire new_Jinkela_wire_167;
    wire _0653_;
    wire new_Jinkela_wire_6470;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_8750;
    wire new_Jinkela_wire_18357;
    wire new_Jinkela_wire_12897;
    wire new_Jinkela_wire_3521;
    wire new_Jinkela_wire_11342;
    wire new_Jinkela_wire_8464;
    wire new_Jinkela_wire_20084;
    wire new_Jinkela_wire_18126;
    wire new_Jinkela_wire_12612;
    wire new_Jinkela_wire_7024;
    wire new_Jinkela_wire_5984;
    wire new_Jinkela_wire_16828;
    wire new_Jinkela_wire_14793;
    wire new_Jinkela_wire_6511;
    wire new_Jinkela_wire_20693;
    wire new_Jinkela_wire_20376;
    wire new_Jinkela_wire_5901;
    wire new_Jinkela_wire_18626;
    wire new_Jinkela_wire_5954;
    wire new_Jinkela_wire_11661;
    wire new_Jinkela_wire_20252;
    wire new_Jinkela_wire_12904;
    wire new_Jinkela_wire_10094;
    wire new_Jinkela_wire_20458;
    wire new_Jinkela_wire_7793;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_13739;
    wire new_Jinkela_wire_10518;
    wire new_Jinkela_wire_5148;
    wire new_Jinkela_wire_21047;
    wire new_Jinkela_wire_14393;
    wire new_Jinkela_wire_18421;
    wire new_Jinkela_wire_5217;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_5236;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_3260;
    wire new_Jinkela_wire_9889;
    wire new_Jinkela_wire_14064;
    wire _0555_;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_15565;
    wire new_Jinkela_wire_12326;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_15013;
    wire new_Jinkela_wire_10205;
    wire new_Jinkela_wire_20232;
    wire new_Jinkela_wire_10169;
    wire new_Jinkela_wire_1941;
    wire new_Jinkela_wire_11490;
    wire new_Jinkela_wire_19461;
    wire new_Jinkela_wire_9000;
    wire new_Jinkela_wire_12956;
    wire new_Jinkela_wire_16440;
    wire new_Jinkela_wire_15809;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_13921;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_7612;
    wire new_Jinkela_wire_10268;
    wire new_Jinkela_wire_2167;
    wire new_Jinkela_wire_11438;
    wire new_Jinkela_wire_6228;
    wire new_Jinkela_wire_8383;
    wire new_Jinkela_wire_12391;
    wire new_Jinkela_wire_19711;
    wire new_Jinkela_wire_6733;
    wire _1380_;
    wire new_Jinkela_wire_2346;
    wire new_Jinkela_wire_10028;
    wire new_Jinkela_wire_7810;
    wire _0383_;
    wire new_Jinkela_wire_13202;
    wire new_Jinkela_wire_2516;
    wire _0058_;
    wire new_Jinkela_wire_12008;
    wire new_Jinkela_wire_7653;
    wire new_Jinkela_wire_13979;
    wire new_Jinkela_wire_12316;
    wire new_Jinkela_wire_16447;
    wire new_Jinkela_wire_17252;
    wire _0455_;
    wire new_Jinkela_wire_7627;
    wire new_Jinkela_wire_8291;
    wire new_Jinkela_wire_18900;
    wire new_Jinkela_wire_5792;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_17068;
    wire new_Jinkela_wire_4375;
    wire new_Jinkela_wire_5694;
    wire new_Jinkela_wire_15357;
    wire new_Jinkela_wire_6670;
    wire new_Jinkela_wire_6087;
    wire new_Jinkela_wire_8343;
    wire new_Jinkela_wire_15304;
    wire new_Jinkela_wire_13753;
    wire new_Jinkela_wire_3242;
    wire new_Jinkela_wire_20419;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_15606;
    wire _1222_;
    wire new_Jinkela_wire_10467;
    wire new_Jinkela_wire_18417;
    wire new_Jinkela_wire_12730;
    wire new_Jinkela_wire_5001;
    wire new_Jinkela_wire_17574;
    wire new_Jinkela_wire_2117;
    wire _1060_;
    wire new_Jinkela_wire_2639;
    wire new_Jinkela_wire_10167;
    wire new_Jinkela_wire_16051;
    wire new_Jinkela_wire_12999;
    wire new_Jinkela_wire_15435;
    wire new_Jinkela_wire_3605;
    wire new_Jinkela_wire_3137;
    wire new_Jinkela_wire_19362;
    wire new_Jinkela_wire_16880;
    wire new_Jinkela_wire_20648;
    wire new_Jinkela_wire_6625;
    wire _1357_;
    wire new_Jinkela_wire_2193;
    wire new_Jinkela_wire_20918;
    wire new_Jinkela_wire_2808;
    wire new_net_3952;
    wire _0444_;
    wire new_Jinkela_wire_18835;
    wire new_Jinkela_wire_17965;
    wire new_Jinkela_wire_9680;
    wire _0299_;
    wire new_Jinkela_wire_14383;
    wire new_Jinkela_wire_12257;
    wire _0537_;
    wire new_Jinkela_wire_9975;
    wire new_Jinkela_wire_5565;
    wire new_Jinkela_wire_20211;
    wire new_Jinkela_wire_7192;
    wire _1326_;
    wire new_Jinkela_wire_7713;
    wire new_Jinkela_wire_12596;
    wire new_Jinkela_wire_9676;
    wire new_Jinkela_wire_14754;
    wire new_Jinkela_wire_1817;
    wire new_Jinkela_wire_3248;
    wire new_Jinkela_wire_7779;
    wire new_Jinkela_wire_10442;
    wire new_Jinkela_wire_17655;
    wire new_Jinkela_wire_14282;
    wire new_Jinkela_wire_20750;
    wire new_Jinkela_wire_4339;
    wire new_Jinkela_wire_4117;
    wire new_Jinkela_wire_20451;
    wire new_Jinkela_wire_7236;
    wire new_Jinkela_wire_9650;
    wire new_Jinkela_wire_20832;
    wire new_Jinkela_wire_6606;
    wire new_Jinkela_wire_13903;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_9588;
    wire new_Jinkela_wire_2334;
    wire _1668_;
    wire new_Jinkela_wire_8179;
    wire new_Jinkela_wire_14002;
    wire new_Jinkela_wire_3032;
    wire _0795_;
    wire new_Jinkela_wire_4708;
    wire new_Jinkela_wire_3276;
    wire new_Jinkela_wire_12370;
    wire new_Jinkela_wire_17370;
    wire new_Jinkela_wire_18690;
    wire new_Jinkela_wire_4035;
    wire _0771_;
    wire _0525_;
    wire new_Jinkela_wire_11107;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_12172;
    wire new_Jinkela_wire_17973;
    wire _0852_;
    wire new_Jinkela_wire_13920;
    wire new_Jinkela_wire_13488;
    wire new_Jinkela_wire_21088;
    wire new_Jinkela_wire_10162;
    wire new_Jinkela_wire_5303;
    wire new_Jinkela_wire_10600;
    wire new_Jinkela_wire_5485;
    wire new_Jinkela_wire_10773;
    wire new_Jinkela_wire_19430;
    wire new_Jinkela_wire_3586;
    wire new_Jinkela_wire_4770;
    wire new_Jinkela_wire_13548;
    wire _0442_;
    wire new_Jinkela_wire_17229;
    wire new_Jinkela_wire_7642;
    wire new_Jinkela_wire_20331;
    wire new_Jinkela_wire_16771;
    wire _1430_;
    wire new_Jinkela_wire_3091;
    wire _0621_;
    wire new_Jinkela_wire_3007;
    wire new_Jinkela_wire_9157;
    wire new_Jinkela_wire_5560;
    wire new_Jinkela_wire_6373;
    wire new_Jinkela_wire_10588;
    wire new_Jinkela_wire_8960;
    wire new_Jinkela_wire_9331;
    wire new_Jinkela_wire_16571;
    wire _1721_;
    wire new_Jinkela_wire_6267;
    wire new_Jinkela_wire_13558;
    wire new_Jinkela_wire_3901;
    wire new_Jinkela_wire_7824;
    wire new_Jinkela_wire_19393;
    wire new_Jinkela_wire_11406;
    wire new_Jinkela_wire_10762;
    wire new_Jinkela_wire_5715;
    wire new_Jinkela_wire_11338;
    wire new_Jinkela_wire_15623;
    wire _0951_;
    wire new_Jinkela_wire_5117;
    wire new_Jinkela_wire_11199;
    wire new_Jinkela_wire_16546;
    wire new_Jinkela_wire_17400;
    wire new_Jinkela_wire_8962;
    wire _1675_;
    wire new_Jinkela_wire_18304;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_15517;
    wire new_Jinkela_wire_16275;
    wire new_Jinkela_wire_12939;
    wire new_Jinkela_wire_19326;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_12402;
    wire new_Jinkela_wire_17990;
    wire new_Jinkela_wire_15902;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_20626;
    wire new_Jinkela_wire_13884;
    wire new_Jinkela_wire_10625;
    wire new_Jinkela_wire_14311;
    wire new_Jinkela_wire_6601;
    wire new_Jinkela_wire_1152;
    wire _0786_;
    wire new_Jinkela_wire_3582;
    wire new_Jinkela_wire_5995;
    wire new_Jinkela_wire_6038;
    wire new_Jinkela_wire_2074;
    wire new_Jinkela_wire_4590;
    wire new_Jinkela_wire_10359;
    wire new_Jinkela_wire_3030;
    wire new_Jinkela_wire_18057;
    wire _1122_;
    wire new_Jinkela_wire_3067;
    wire new_Jinkela_wire_17762;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_3654;
    wire new_Jinkela_wire_6746;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_18151;
    wire new_Jinkela_wire_13366;
    wire new_Jinkela_wire_16188;
    wire new_Jinkela_wire_11511;
    wire new_Jinkela_wire_2817;
    wire new_Jinkela_wire_6977;
    wire new_Jinkela_wire_6001;
    wire new_Jinkela_wire_2371;
    wire new_Jinkela_wire_7994;
    wire _1009_;
    wire new_Jinkela_wire_18936;
    wire new_Jinkela_wire_15663;
    wire _0843_;
    wire new_Jinkela_wire_9647;
    wire new_Jinkela_wire_11233;
    wire new_Jinkela_wire_15790;
    wire new_Jinkela_wire_15361;
    wire new_Jinkela_wire_8836;
    wire new_Jinkela_wire_15534;
    wire new_Jinkela_wire_13231;
    wire new_Jinkela_wire_2983;
    wire new_Jinkela_wire_5690;
    wire new_Jinkela_wire_13779;
    wire new_Jinkela_wire_2379;
    wire new_Jinkela_wire_2374;
    wire new_Jinkela_wire_11143;
    wire new_Jinkela_wire_10992;
    wire new_Jinkela_wire_19380;
    wire new_Jinkela_wire_19423;
    wire new_Jinkela_wire_13830;
    wire new_Jinkela_wire_3972;
    wire new_Jinkela_wire_1883;
    wire new_Jinkela_wire_5345;
    wire new_Jinkela_wire_4358;
    wire new_Jinkela_wire_8941;
    wire new_Jinkela_wire_19212;
    wire new_Jinkela_wire_17979;
    wire new_Jinkela_wire_15482;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_6302;
    wire new_Jinkela_wire_21153;
    wire new_Jinkela_wire_14449;
    wire new_Jinkela_wire_8631;
    wire new_Jinkela_wire_20755;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_3640;
    wire new_Jinkela_wire_13164;
    wire new_Jinkela_wire_5302;
    wire new_Jinkela_wire_10845;
    wire new_Jinkela_wire_21239;
    wire new_Jinkela_wire_17248;
    wire new_Jinkela_wire_7949;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_5125;
    wire new_Jinkela_wire_10474;
    wire new_Jinkela_wire_8659;
    wire new_Jinkela_wire_18846;
    wire new_Jinkela_wire_17522;
    wire new_Jinkela_wire_14979;
    wire new_Jinkela_wire_14437;
    wire new_Jinkela_wire_9631;
    wire new_Jinkela_wire_4891;
    wire new_Jinkela_wire_8689;
    wire new_Jinkela_wire_11759;
    wire new_Jinkela_wire_10524;
    wire new_Jinkela_wire_4682;
    wire new_Jinkela_wire_15757;
    wire new_Jinkela_wire_14573;
    wire new_Jinkela_wire_19586;
    wire new_Jinkela_wire_9726;
    wire new_Jinkela_wire_9284;
    wire new_Jinkela_wire_19283;
    wire new_Jinkela_wire_1135;
    wire new_Jinkela_wire_19268;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_21109;
    wire new_Jinkela_wire_16544;
    wire new_Jinkela_wire_377;
    wire _0936_;
    wire new_Jinkela_wire_11371;
    wire new_Jinkela_wire_3952;
    wire new_Jinkela_wire_3336;
    wire new_Jinkela_wire_19396;
    wire new_Jinkela_wire_14467;
    wire new_Jinkela_wire_18201;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_14671;
    wire new_Jinkela_wire_11266;
    wire new_Jinkela_wire_12787;
    wire new_Jinkela_wire_6408;
    wire new_Jinkela_wire_10276;
    wire new_Jinkela_wire_17002;
    wire new_Jinkela_wire_15458;
    wire new_Jinkela_wire_20304;
    wire new_Jinkela_wire_16792;
    wire _0378_;
    wire new_Jinkela_wire_13111;
    wire new_Jinkela_wire_13929;
    wire new_Jinkela_wire_4370;
    wire _0262_;
    wire new_Jinkela_wire_14003;
    wire new_Jinkela_wire_13125;
    wire new_Jinkela_wire_17460;
    wire new_Jinkela_wire_6389;
    wire new_Jinkela_wire_7377;
    wire new_Jinkela_wire_9286;
    wire new_Jinkela_wire_1996;
    wire new_Jinkela_wire_19134;
    wire new_Jinkela_wire_9152;
    wire new_Jinkela_wire_3725;
    wire _0259_;
    wire new_Jinkela_wire_15885;
    wire new_Jinkela_wire_3452;
    wire new_Jinkela_wire_11935;
    wire _1662_;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_16831;
    wire new_Jinkela_wire_6643;
    wire new_Jinkela_wire_16423;
    wire new_Jinkela_wire_21106;
    wire _1801_;
    wire new_Jinkela_wire_12622;
    wire new_Jinkela_wire_3163;
    wire new_Jinkela_wire_14993;
    wire new_Jinkela_wire_8714;
    wire new_Jinkela_wire_16071;
    wire new_Jinkela_wire_13102;
    wire _0671_;
    wire new_Jinkela_wire_15471;
    wire new_Jinkela_wire_17200;
    wire new_Jinkela_wire_2365;
    wire new_Jinkela_wire_8229;
    wire new_Jinkela_wire_18250;
    wire new_Jinkela_wire_4773;
    wire new_Jinkela_wire_8014;
    wire new_Jinkela_wire_5363;
    wire new_Jinkela_wire_20965;
    wire new_Jinkela_wire_9095;
    wire _1604_;
    wire new_Jinkela_wire_15053;
    wire new_Jinkela_wire_2539;
    wire new_Jinkela_wire_15600;
    wire new_Jinkela_wire_20048;
    wire new_Jinkela_wire_7304;
    wire new_Jinkela_wire_3196;
    wire new_Jinkela_wire_17030;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_10312;
    wire new_Jinkela_wire_11673;
    wire new_Jinkela_wire_3445;
    wire new_Jinkela_wire_19942;
    wire new_Jinkela_wire_2982;
    wire new_Jinkela_wire_10346;
    wire new_Jinkela_wire_14877;
    wire new_Jinkela_wire_6320;
    wire new_Jinkela_wire_14445;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_14345;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_19654;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_7897;
    wire new_Jinkela_wire_14134;
    wire new_Jinkela_wire_3646;
    wire new_Jinkela_wire_5092;
    wire new_Jinkela_wire_12933;
    wire _0820_;
    wire new_Jinkela_wire_6907;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_9413;
    wire new_Jinkela_wire_10266;
    wire new_Jinkela_wire_9222;
    wire _0089_;
    wire new_Jinkela_wire_9893;
    wire new_Jinkela_wire_8847;
    wire _0140_;
    wire new_Jinkela_wire_11056;
    wire _0994_;
    wire new_Jinkela_wire_12364;
    wire new_Jinkela_wire_2198;
    wire new_Jinkela_wire_2216;
    wire new_Jinkela_wire_8556;
    wire new_Jinkela_wire_12981;
    wire new_Jinkela_wire_6063;
    wire new_Jinkela_wire_18001;
    wire new_Jinkela_wire_3068;
    wire new_Jinkela_wire_4842;
    wire new_Jinkela_wire_2237;
    wire new_Jinkela_wire_16054;
    wire new_Jinkela_wire_7973;
    wire new_Jinkela_wire_20122;
    wire new_Jinkela_wire_15764;
    wire new_Jinkela_wire_20200;
    wire new_Jinkela_wire_19763;
    wire new_Jinkela_wire_19728;
    wire new_Jinkela_wire_11369;
    wire new_Jinkela_wire_7997;
    wire new_Jinkela_wire_20101;
    wire new_Jinkela_wire_3559;
    wire new_Jinkela_wire_16602;
    wire new_Jinkela_wire_13247;
    wire new_Jinkela_wire_3895;
    wire new_Jinkela_wire_10686;
    wire new_Jinkela_wire_15454;
    wire new_Jinkela_wire_1861;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_20846;
    wire new_Jinkela_wire_5970;
    wire new_Jinkela_wire_7603;
    wire new_Jinkela_wire_13636;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_13212;
    wire new_Jinkela_wire_17563;
    wire new_Jinkela_wire_14086;
    wire _1420_;
    wire new_Jinkela_wire_20942;
    wire new_Jinkela_wire_13099;
    wire new_Jinkela_wire_5923;
    wire new_Jinkela_wire_4114;
    wire new_Jinkela_wire_21178;
    wire new_Jinkela_wire_19103;
    wire new_Jinkela_wire_8508;
    wire new_Jinkela_wire_14954;
    wire new_Jinkela_wire_10349;
    wire new_Jinkela_wire_19943;
    wire new_Jinkela_wire_7995;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_9552;
    wire new_Jinkela_wire_9355;
    wire new_Jinkela_wire_12620;
    wire new_Jinkela_wire_5097;
    wire new_Jinkela_wire_16868;
    wire new_Jinkela_wire_4166;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_21274;
    wire new_Jinkela_wire_6833;
    wire new_Jinkela_wire_19063;
    wire _0992_;
    wire new_Jinkela_wire_15549;
    wire new_Jinkela_wire_16161;
    wire new_Jinkela_wire_12117;
    wire new_Jinkela_wire_14762;
    wire new_Jinkela_wire_5571;
    wire new_Jinkela_wire_15322;
    wire new_Jinkela_wire_15029;
    wire new_Jinkela_wire_15181;
    wire new_Jinkela_wire_11622;
    wire new_Jinkela_wire_7786;
    wire new_Jinkela_wire_18611;
    wire new_Jinkela_wire_17939;
    wire _1465_;
    wire new_Jinkela_wire_3631;
    wire new_Jinkela_wire_5508;
    wire new_Jinkela_wire_4093;
    wire new_Jinkela_wire_12197;
    wire new_Jinkela_wire_20015;
    wire new_Jinkela_wire_8792;
    wire new_Jinkela_wire_4388;
    wire new_Jinkela_wire_10766;
    wire new_Jinkela_wire_7796;
    wire new_Jinkela_wire_19183;
    wire new_Jinkela_wire_21001;
    wire _1446_;
    wire new_Jinkela_wire_3499;
    wire new_Jinkela_wire_17008;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_8691;
    wire new_Jinkela_wire_21126;
    wire new_Jinkela_wire_14686;
    wire new_Jinkela_wire_11512;
    wire new_Jinkela_wire_4610;
    wire new_Jinkela_wire_14730;
    wire new_Jinkela_wire_8019;
    wire new_Jinkela_wire_19616;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_20974;
    wire new_Jinkela_wire_18195;
    wire new_Jinkela_wire_15676;
    wire new_Jinkela_wire_8581;
    wire new_Jinkela_wire_18761;
    wire new_Jinkela_wire_6749;
    wire new_Jinkela_wire_20539;
    wire new_Jinkela_wire_9370;
    wire new_Jinkela_wire_6071;
    wire new_Jinkela_wire_4367;
    wire new_Jinkela_wire_9192;
    wire new_Jinkela_wire_10186;
    wire new_Jinkela_wire_3279;
    wire new_Jinkela_wire_9350;
    wire new_Jinkela_wire_10718;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_3887;
    wire new_Jinkela_wire_18328;
    wire new_Jinkela_wire_17442;
    wire new_Jinkela_wire_12380;
    wire new_Jinkela_wire_3573;
    wire new_Jinkela_wire_18032;
    wire new_Jinkela_wire_16036;
    wire new_Jinkela_wire_6431;
    wire new_Jinkela_wire_17433;
    wire new_Jinkela_wire_7726;
    wire new_Jinkela_wire_14249;
    wire new_Jinkela_wire_15196;
    wire new_Jinkela_wire_12000;
    wire new_Jinkela_wire_13865;
    wire new_Jinkela_wire_3736;
    wire new_Jinkela_wire_4373;
    wire new_Jinkela_wire_5369;
    wire new_Jinkela_wire_11508;
    wire new_Jinkela_wire_7629;
    wire new_Jinkela_wire_20759;
    wire new_Jinkela_wire_21269;
    wire new_Jinkela_wire_3599;
    wire new_Jinkela_wire_17854;
    wire new_Jinkela_wire_4254;
    wire new_Jinkela_wire_2756;
    wire new_Jinkela_wire_11084;
    wire new_Jinkela_wire_2590;
    wire new_Jinkela_wire_12229;
    wire _1113_;
    wire new_Jinkela_wire_19378;
    wire new_Jinkela_wire_20460;
    wire new_Jinkela_wire_6073;
    wire new_Jinkela_wire_10180;
    wire new_Jinkela_wire_3053;
    wire _1557_;
    wire new_Jinkela_wire_19568;
    wire new_Jinkela_wire_13784;
    wire new_Jinkela_wire_19263;
    wire new_Jinkela_wire_8539;
    wire new_Jinkela_wire_7747;
    wire new_Jinkela_wire_14459;
    wire new_Jinkela_wire_12998;
    wire new_Jinkela_wire_4097;
    wire _1208_;
    wire new_Jinkela_wire_19189;
    wire new_Jinkela_wire_3593;
    wire new_Jinkela_wire_10930;
    wire new_Jinkela_wire_7473;
    wire new_Jinkela_wire_17425;
    wire new_Jinkela_wire_10840;
    wire new_Jinkela_wire_14825;
    wire new_Jinkela_wire_5214;
    wire new_Jinkela_wire_2978;
    wire new_Jinkela_wire_10517;
    wire new_Jinkela_wire_8419;
    wire new_Jinkela_wire_15558;
    wire new_Jinkela_wire_7637;
    wire new_Jinkela_wire_17879;
    wire new_Jinkela_wire_15449;
    wire new_Jinkela_wire_13999;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_7813;
    wire new_Jinkela_wire_2446;
    wire _0194_;
    wire new_Jinkela_wire_15685;
    wire new_Jinkela_wire_18271;
    wire _0945_;
    wire new_Jinkela_wire_10023;
    wire new_Jinkela_wire_5094;
    wire new_Jinkela_wire_6515;
    wire new_Jinkela_wire_11988;
    wire new_Jinkela_wire_9851;
    wire new_Jinkela_wire_4274;
    wire new_Jinkela_wire_9349;
    wire new_Jinkela_wire_21164;
    wire new_Jinkela_wire_4755;
    wire new_Jinkela_wire_3898;
    wire new_Jinkela_wire_9820;
    wire new_Jinkela_wire_9524;
    wire new_Jinkela_wire_18870;
    wire new_Jinkela_wire_11773;
    wire new_Jinkela_wire_19986;
    wire new_Jinkela_wire_4075;
    wire _0708_;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_16554;
    wire new_Jinkela_wire_20763;
    wire new_Jinkela_wire_16616;
    wire new_Jinkela_wire_19353;
    wire new_Jinkela_wire_18602;
    wire new_Jinkela_wire_6295;
    wire _0781_;
    wire new_Jinkela_wire_6231;
    wire new_Jinkela_wire_2965;
    wire new_Jinkela_wire_3511;
    wire new_Jinkela_wire_15965;
    wire new_Jinkela_wire_20603;
    wire new_Jinkela_wire_16950;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_7641;
    wire new_Jinkela_wire_7578;
    wire new_Jinkela_wire_13740;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_2557;
    wire new_Jinkela_wire_13597;
    wire new_Jinkela_wire_16243;
    wire new_Jinkela_wire_10425;
    wire new_Jinkela_wire_10018;
    wire new_Jinkela_wire_9434;
    wire new_Jinkela_wire_12126;
    wire new_Jinkela_wire_16445;
    wire new_Jinkela_wire_9887;
    wire new_Jinkela_wire_12160;
    wire new_Jinkela_wire_12865;
    wire new_Jinkela_wire_7540;
    wire new_Jinkela_wire_18406;
    wire new_Jinkela_wire_16978;
    wire new_Jinkela_wire_11908;
    wire new_Jinkela_wire_14355;
    wire new_Jinkela_wire_13568;
    wire new_Jinkela_wire_6929;
    wire new_Jinkela_wire_11387;
    wire new_Jinkela_wire_9923;
    wire new_Jinkela_wire_2773;
    wire new_Jinkela_wire_13069;
    wire new_Jinkela_wire_7811;
    wire new_Jinkela_wire_13950;
    wire new_Jinkela_wire_4621;
    wire new_Jinkela_wire_19705;
    wire _1476_;
    wire new_Jinkela_wire_14767;
    wire new_Jinkela_wire_13917;
    wire new_Jinkela_wire_15274;
    wire new_Jinkela_wire_20963;
    wire new_Jinkela_wire_14926;
    wire new_Jinkela_wire_12512;
    wire new_Jinkela_wire_18435;
    wire new_Jinkela_wire_15052;
    wire new_Jinkela_wire_6102;
    wire new_Jinkela_wire_13555;
    wire new_Jinkela_wire_21205;
    wire new_Jinkela_wire_19867;
    wire new_Jinkela_wire_14889;
    wire new_Jinkela_wire_16965;
    wire _0848_;
    wire new_Jinkela_wire_17731;
    wire new_Jinkela_wire_2176;
    wire _0317_;
    wire new_Jinkela_wire_8238;
    wire new_Jinkela_wire_7311;
    wire new_Jinkela_wire_10423;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_2345;
    wire new_Jinkela_wire_15492;
    wire new_Jinkela_wire_13890;
    wire new_Jinkela_wire_18560;
    wire _0337_;
    wire new_Jinkela_wire_5755;
    wire new_Jinkela_wire_13263;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_16183;
    wire _1545_;
    wire new_Jinkela_wire_8972;
    wire new_Jinkela_wire_8611;
    wire new_Jinkela_wire_13839;
    wire new_Jinkela_wire_14867;
    wire new_Jinkela_wire_14012;
    wire new_Jinkela_wire_6485;
    wire new_Jinkela_wire_14058;
    wire new_Jinkela_wire_18177;
    wire new_Jinkela_wire_5370;
    wire new_Jinkela_wire_10341;
    wire new_Jinkela_wire_18874;
    wire new_Jinkela_wire_6922;
    wire new_Jinkela_wire_5664;
    wire new_Jinkela_wire_4313;
    wire new_Jinkela_wire_6516;
    wire new_Jinkela_wire_20247;
    wire new_Jinkela_wire_7520;
    wire new_Jinkela_wire_8593;
    wire new_Jinkela_wire_9569;
    wire new_Jinkela_wire_5852;
    wire new_Jinkela_wire_11397;
    wire _1549_;
    wire new_Jinkela_wire_3563;
    wire new_Jinkela_wire_4729;
    wire new_Jinkela_wire_14812;
    wire new_Jinkela_wire_12833;
    wire new_Jinkela_wire_17946;
    wire new_Jinkela_wire_15681;
    wire new_Jinkela_wire_3897;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_20440;
    wire new_Jinkela_wire_12885;
    wire new_Jinkela_wire_2439;
    wire new_Jinkela_wire_7380;
    wire new_Jinkela_wire_17024;
    wire new_Jinkela_wire_18550;
    wire new_Jinkela_wire_3622;
    wire _1533_;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_12943;
    wire new_Jinkela_wire_7199;
    wire new_Jinkela_wire_9549;
    wire new_Jinkela_wire_4504;
    wire new_Jinkela_wire_19660;
    wire new_Jinkela_wire_2745;
    wire _1076_;
    wire new_Jinkela_wire_16399;
    wire new_Jinkela_wire_8411;
    wire new_Jinkela_wire_19318;
    wire new_Jinkela_wire_8488;
    wire new_Jinkela_wire_16200;
    wire new_Jinkela_wire_11113;
    wire new_Jinkela_wire_12005;
    wire _0760_;
    wire new_Jinkela_wire_3955;
    wire new_Jinkela_wire_7761;
    wire new_Jinkela_wire_18875;
    wire new_Jinkela_wire_16776;
    wire new_Jinkela_wire_20373;
    wire new_Jinkela_wire_7198;
    wire _1175_;
    wire new_Jinkela_wire_11515;
    wire new_Jinkela_wire_2492;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_7462;
    wire new_Jinkela_wire_15002;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_12872;
    wire new_Jinkela_wire_11586;
    wire new_Jinkela_wire_17785;
    wire new_Jinkela_wire_6255;
    wire _0575_;
    wire new_Jinkela_wire_15388;
    wire new_Jinkela_wire_5199;
    wire new_Jinkela_wire_12304;
    wire new_Jinkela_wire_11655;
    wire new_Jinkela_wire_5502;
    wire _1341_;
    wire new_Jinkela_wire_7971;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_4552;
    wire _0604_;
    wire new_Jinkela_wire_16167;
    wire _0237_;
    wire new_Jinkela_wire_2876;
    wire new_Jinkela_wire_12856;
    wire new_Jinkela_wire_13503;
    wire new_Jinkela_wire_18382;
    wire new_Jinkela_wire_16630;
    wire new_Jinkela_wire_11738;
    wire new_Jinkela_wire_11507;
    wire new_Jinkela_wire_18076;
    wire new_Jinkela_wire_8644;
    wire new_Jinkela_wire_8493;
    wire new_Jinkela_wire_21170;
    wire new_Jinkela_wire_21247;
    wire new_Jinkela_wire_19114;
    wire new_Jinkela_wire_9764;
    wire new_Jinkela_wire_4537;
    wire _0527_;
    wire new_Jinkela_wire_21141;
    wire new_Jinkela_wire_5304;
    wire new_Jinkela_wire_11305;
    wire new_Jinkela_wire_18922;
    wire new_Jinkela_wire_20718;
    wire new_Jinkela_wire_3924;
    wire new_Jinkela_wire_6351;
    wire new_Jinkela_wire_6539;
    wire new_Jinkela_wire_980;
    wire _1336_;
    wire new_Jinkela_wire_19412;
    wire new_Jinkela_wire_18116;
    wire _0875_;
    wire new_Jinkela_wire_14109;
    wire new_Jinkela_wire_18168;
    wire new_Jinkela_wire_13106;
    wire new_Jinkela_wire_20706;
    wire new_Jinkela_wire_4713;
    wire new_Jinkela_wire_2141;
    wire new_Jinkela_wire_10316;
    wire new_Jinkela_wire_15859;
    wire new_Jinkela_wire_1951;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_8133;
    wire new_Jinkela_wire_17393;
    wire new_Jinkela_wire_21060;
    wire new_Jinkela_wire_8626;
    wire new_Jinkela_wire_3641;
    wire new_Jinkela_wire_16567;
    wire new_Jinkela_wire_16178;
    wire new_Jinkela_wire_15501;
    wire new_Jinkela_wire_8551;
    wire new_Jinkela_wire_12269;
    wire new_Jinkela_wire_11545;
    wire new_Jinkela_wire_2251;
    wire new_Jinkela_wire_2467;
    wire _1681_;
    wire new_Jinkela_wire_18436;
    wire new_Jinkela_wire_1843;
    wire new_Jinkela_wire_12551;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_16896;
    wire new_Jinkela_wire_3915;
    wire new_Jinkela_wire_7387;
    wire new_Jinkela_wire_15725;
    wire new_Jinkela_wire_9321;
    wire new_Jinkela_wire_14152;
    wire new_Jinkela_wire_10152;
    wire new_Jinkela_wire_5278;
    wire _0928_;
    wire new_Jinkela_wire_17931;
    wire new_Jinkela_wire_11015;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_13955;
    wire new_Jinkela_wire_7950;
    wire new_Jinkela_wire_13435;
    wire new_Jinkela_wire_17726;
    wire new_Jinkela_wire_3106;
    wire new_Jinkela_wire_18751;
    wire new_Jinkela_wire_10708;
    wire new_Jinkela_wire_4167;
    wire new_Jinkela_wire_6317;
    wire new_Jinkela_wire_2499;
    wire new_Jinkela_wire_20856;
    wire new_Jinkela_wire_19107;
    wire new_Jinkela_wire_5635;
    wire new_Jinkela_wire_13121;
    wire new_Jinkela_wire_13637;
    wire new_Jinkela_wire_7622;
    wire _0667_;
    wire new_Jinkela_wire_20147;
    wire new_Jinkela_wire_1975;
    wire _1820_;
    wire new_Jinkela_wire_20928;
    wire new_Jinkela_wire_2926;
    wire new_Jinkela_wire_16851;
    wire new_Jinkela_wire_1906;
    wire new_Jinkela_wire_7728;
    wire new_Jinkela_wire_4337;
    wire new_Jinkela_wire_2768;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_11274;
    wire new_Jinkela_wire_6734;
    wire new_Jinkela_wire_6502;
    wire new_Jinkela_wire_8212;
    wire new_Jinkela_wire_9387;
    wire new_Jinkela_wire_5784;
    wire new_Jinkela_wire_8692;
    wire new_Jinkela_wire_19180;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_19591;
    wire new_Jinkela_wire_8135;
    wire new_Jinkela_wire_10134;
    wire new_Jinkela_wire_13295;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_17983;
    wire new_Jinkela_wire_12571;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_18655;
    wire new_Jinkela_wire_16403;
    wire new_Jinkela_wire_17207;
    wire new_Jinkela_wire_3264;
    wire new_Jinkela_wire_3268;
    wire new_Jinkela_wire_16777;
    wire new_Jinkela_wire_4178;
    wire new_Jinkela_wire_15198;
    wire new_Jinkela_wire_19987;
    wire new_Jinkela_wire_13490;
    wire new_Jinkela_wire_6284;
    wire new_Jinkela_wire_13483;
    wire new_Jinkela_wire_5254;
    wire _1762_;
    wire new_Jinkela_wire_14779;
    wire new_Jinkela_wire_4515;
    wire new_Jinkela_wire_18345;
    wire new_Jinkela_wire_4156;
    wire new_Jinkela_wire_12923;
    wire new_Jinkela_wire_3409;
    wire new_Jinkela_wire_17638;
    wire new_Jinkela_wire_14646;
    wire new_Jinkela_wire_15792;
    wire new_Jinkela_wire_20222;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_19148;
    wire new_Jinkela_wire_16987;
    wire new_Jinkela_wire_13566;
    wire new_Jinkela_wire_12186;
    wire new_Jinkela_wire_2059;
    wire new_Jinkela_wire_6084;
    wire new_Jinkela_wire_2673;
    wire new_Jinkela_wire_9260;
    wire new_Jinkela_wire_8289;
    wire new_Jinkela_wire_6845;
    wire new_Jinkela_wire_15648;
    wire new_Jinkela_wire_6145;
    wire new_Jinkela_wire_6655;
    wire new_Jinkela_wire_7904;
    wire new_Jinkela_wire_5677;
    wire new_Jinkela_wire_6607;
    wire _0381_;
    wire new_Jinkela_wire_18679;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_2174;
    wire new_Jinkela_wire_9858;
    wire new_Jinkela_wire_19041;
    wire _1524_;
    wire new_Jinkela_wire_1886;
    wire new_Jinkela_wire_6456;
    wire new_Jinkela_wire_3837;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_8629;
    wire new_Jinkela_wire_2116;
    wire new_Jinkela_wire_19192;
    wire new_Jinkela_wire_14023;
    wire new_Jinkela_wire_5787;
    wire new_Jinkela_wire_2910;
    wire new_Jinkela_wire_13133;
    wire new_Jinkela_wire_2520;
    wire new_Jinkela_wire_4147;
    wire new_Jinkela_wire_8674;
    wire new_Jinkela_wire_10046;
    wire new_Jinkela_wire_4332;
    wire new_Jinkela_wire_20406;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_11601;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_19933;
    wire new_Jinkela_wire_18872;
    wire new_Jinkela_wire_6114;
    wire new_Jinkela_wire_14398;
    wire new_Jinkela_wire_11922;
    wire new_Jinkela_wire_15135;
    wire new_Jinkela_wire_18533;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_7991;
    wire new_Jinkela_wire_7318;
    wire new_Jinkela_wire_16173;
    wire new_Jinkela_wire_13517;
    wire new_Jinkela_wire_15983;
    wire new_Jinkela_wire_5438;
    wire new_Jinkela_wire_17858;
    wire new_Jinkela_wire_19528;
    wire new_Jinkela_wire_6847;
    wire new_Jinkela_wire_20444;
    wire _1649_;
    wire new_Jinkela_wire_14420;
    wire new_Jinkela_wire_4389;
    wire new_Jinkela_wire_11059;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_12899;
    wire new_Jinkela_wire_8725;
    wire _0125_;
    wire new_Jinkela_wire_18373;
    wire new_Jinkela_wire_11211;
    wire new_Jinkela_wire_5011;
    wire new_Jinkela_wire_13259;
    wire new_Jinkela_wire_17320;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_14549;
    wire new_Jinkela_wire_20981;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_8732;
    wire new_Jinkela_wire_17224;
    wire _0360_;
    wire new_Jinkela_wire_16726;
    wire new_Jinkela_wire_3318;
    wire new_Jinkela_wire_20657;
    wire new_Jinkela_wire_19182;
    wire new_Jinkela_wire_17849;
    wire new_Jinkela_wire_18246;
    wire new_Jinkela_wire_18047;
    wire new_Jinkela_wire_7374;
    wire new_Jinkela_wire_18127;
    wire new_Jinkela_wire_12449;
    wire _1132_;
    wire _0256_;
    wire new_Jinkela_wire_13622;
    wire new_Jinkela_wire_3649;
    wire _0245_;
    wire new_Jinkela_wire_14272;
    wire new_Jinkela_wire_20730;
    wire _1819_;
    wire new_Jinkela_wire_6579;
    wire _0375_;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_6695;
    wire new_Jinkela_wire_3359;
    wire new_Jinkela_wire_11602;
    wire new_Jinkela_wire_4715;
    wire new_Jinkela_wire_10199;
    wire new_Jinkela_wire_3807;
    wire new_Jinkela_wire_14833;
    wire new_Jinkela_wire_10315;
    wire new_Jinkela_wire_20739;
    wire new_Jinkela_wire_19964;
    wire new_Jinkela_wire_17317;
    wire new_Jinkela_wire_2146;
    wire new_Jinkela_wire_16150;
    wire new_Jinkela_wire_16465;
    wire new_Jinkela_wire_14342;
    wire new_Jinkela_wire_4711;
    wire new_Jinkela_wire_3437;
    wire new_Jinkela_wire_16096;
    wire new_Jinkela_wire_5142;
    wire new_Jinkela_wire_2581;
    wire new_Jinkela_wire_1230;
    wire _1203_;
    wire new_Jinkela_wire_14862;
    wire new_Jinkela_wire_9855;
    wire new_Jinkela_wire_4396;
    wire new_Jinkela_wire_20221;
    wire new_Jinkela_wire_6866;
    wire new_Jinkela_wire_15261;
    wire new_Jinkela_wire_20704;
    wire new_Jinkela_wire_21020;
    wire new_Jinkela_wire_8194;
    wire new_Jinkela_wire_15896;
    wire new_Jinkela_wire_12974;
    wire _0388_;
    wire new_Jinkela_wire_12984;
    wire new_Jinkela_wire_11989;
    wire new_Jinkela_wire_6674;
    wire new_Jinkela_wire_11228;
    wire new_Jinkela_wire_8542;
    wire new_Jinkela_wire_9278;
    wire new_Jinkela_wire_13617;
    wire new_Jinkela_wire_8122;
    wire new_Jinkela_wire_18664;
    wire new_Jinkela_wire_20023;
    wire new_Jinkela_wire_3638;
    wire new_Jinkela_wire_13363;
    wire new_Jinkela_wire_12951;
    wire new_Jinkela_wire_19050;
    wire new_Jinkela_wire_11619;
    wire new_Jinkela_wire_8339;
    wire new_Jinkela_wire_11482;
    wire new_Jinkela_wire_12675;
    wire new_Jinkela_wire_12898;
    wire new_Jinkela_wire_13105;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_5290;
    wire new_Jinkela_wire_12783;
    wire new_Jinkela_wire_16392;
    wire new_Jinkela_wire_15982;
    wire new_Jinkela_wire_3387;
    wire new_Jinkela_wire_624;
    wire _1210_;
    wire new_Jinkela_wire_8980;
    wire new_Jinkela_wire_6685;
    wire new_Jinkela_wire_2043;
    wire new_net_3918;
    wire new_Jinkela_wire_2599;
    wire new_Jinkela_wire_4224;
    wire new_Jinkela_wire_16709;
    wire new_Jinkela_wire_7309;
    wire new_Jinkela_wire_17578;
    wire new_Jinkela_wire_20360;
    wire new_Jinkela_wire_8456;
    wire new_Jinkela_wire_15193;
    wire new_Jinkela_wire_15457;
    wire _0584_;
    wire new_Jinkela_wire_6066;
    wire new_Jinkela_wire_8022;
    wire new_Jinkela_wire_14268;
    wire new_Jinkela_wire_2206;
    wire new_Jinkela_wire_15991;
    wire _0529_;
    wire new_Jinkela_wire_12655;
    wire new_Jinkela_wire_3354;
    wire new_Jinkela_wire_14822;
    wire _1792_;
    wire new_Jinkela_wire_14614;
    wire new_Jinkela_wire_3847;
    wire new_Jinkela_wire_10225;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_5646;
    wire new_Jinkela_wire_9922;
    wire new_Jinkela_wire_14896;
    wire new_Jinkela_wire_2189;
    wire new_Jinkela_wire_20258;
    wire new_Jinkela_wire_7194;
    wire new_Jinkela_wire_5877;
    wire new_Jinkela_wire_10241;
    wire new_Jinkela_wire_2285;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_14212;
    wire new_Jinkela_wire_9283;
    wire new_Jinkela_wire_10947;
    wire new_Jinkela_wire_6214;
    wire new_Jinkela_wire_4506;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_17612;
    wire new_Jinkela_wire_14737;
    wire new_Jinkela_wire_18525;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_17693;
    wire new_Jinkela_wire_5879;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_9603;
    wire new_Jinkela_wire_12385;
    wire new_Jinkela_wire_5391;
    wire new_Jinkela_wire_13174;
    wire new_Jinkela_wire_20455;
    wire new_Jinkela_wire_14361;
    wire new_Jinkela_wire_15408;
    wire new_Jinkela_wire_11535;
    wire new_Jinkela_wire_16155;
    wire new_Jinkela_wire_8754;
    wire new_Jinkela_wire_3252;
    wire new_Jinkela_wire_20278;
    wire _0246_;
    wire new_Jinkela_wire_10035;
    wire new_Jinkela_wire_2390;
    wire new_Jinkela_wire_9776;
    wire new_Jinkela_wire_10126;
    wire new_Jinkela_wire_14736;
    wire new_Jinkela_wire_4467;
    wire new_Jinkela_wire_13229;
    wire _0233_;
    wire new_Jinkela_wire_4815;
    wire new_Jinkela_wire_16785;
    wire new_Jinkela_wire_5713;
    wire new_Jinkela_wire_12930;
    wire new_Jinkela_wire_15945;
    wire new_Jinkela_wire_18723;
    wire new_Jinkela_wire_12631;
    wire new_Jinkela_wire_6992;
    wire new_Jinkela_wire_7370;
    wire new_Jinkela_wire_17663;
    wire new_Jinkela_wire_15645;
    wire new_Jinkela_wire_13364;
    wire new_Jinkela_wire_17005;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_19403;
    wire _0566_;
    wire new_Jinkela_wire_19712;
    wire new_Jinkela_wire_13861;
    wire new_Jinkela_wire_17512;
    wire new_Jinkela_wire_21287;
    wire new_Jinkela_wire_6413;
    wire new_Jinkela_wire_15270;
    wire new_Jinkela_wire_5232;
    wire new_Jinkela_wire_14401;
    wire _0267_;
    wire new_Jinkela_wire_9045;
    wire new_Jinkela_wire_14289;
    wire new_Jinkela_wire_9810;
    wire new_Jinkela_wire_2016;
    wire new_Jinkela_wire_11437;
    wire new_Jinkela_wire_5300;
    wire new_Jinkela_wire_3133;
    wire new_Jinkela_wire_4607;
    wire new_Jinkela_wire_10903;
    wire _1016_;
    wire new_Jinkela_wire_16515;
    wire new_Jinkela_wire_15250;
    wire new_Jinkela_wire_15390;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_17044;
    wire new_Jinkela_wire_14043;
    wire new_Jinkela_wire_1309;
    wire new_Jinkela_wire_13402;
    wire new_Jinkela_wire_21055;
    wire new_Jinkela_wire_15531;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_19052;
    wire new_Jinkela_wire_13735;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_7693;
    wire _1627_;
    wire new_Jinkela_wire_21080;
    wire _0148_;
    wire new_Jinkela_wire_13682;
    wire new_Jinkela_wire_2986;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_17437;
    wire new_Jinkela_wire_12089;
    wire new_Jinkela_wire_8085;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_16126;
    wire new_Jinkela_wire_16205;
    wire new_Jinkela_wire_5099;
    wire new_Jinkela_wire_3298;
    wire new_Jinkela_wire_12471;
    wire new_Jinkela_wire_18523;
    wire new_Jinkela_wire_10880;
    wire new_Jinkela_wire_6904;
    wire new_Jinkela_wire_11847;
    wire new_Jinkela_wire_20664;
    wire new_Jinkela_wire_3062;
    wire new_Jinkela_wire_6136;
    wire new_Jinkela_wire_15037;
    wire _0929_;
    wire new_Jinkela_wire_18236;
    wire new_Jinkela_wire_7183;
    wire new_Jinkela_wire_12260;
    wire new_Jinkela_wire_14741;
    wire new_Jinkela_wire_3601;
    wire new_Jinkela_wire_19792;
    wire new_Jinkela_wire_4048;
    wire new_Jinkela_wire_7263;
    wire new_Jinkela_wire_12756;
    wire new_Jinkela_wire_16590;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_15874;
    wire new_Jinkela_wire_3004;
    wire new_Jinkela_wire_19469;
    wire new_Jinkela_wire_20477;
    wire new_Jinkela_wire_2114;
    wire new_Jinkela_wire_14248;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_7765;
    wire new_Jinkela_wire_5692;
    wire _1354_;
    wire _1640_;
    wire new_Jinkela_wire_2845;
    wire _0830_;
    wire new_Jinkela_wire_4392;
    wire new_Jinkela_wire_7806;
    wire new_Jinkela_wire_17506;
    wire new_Jinkela_wire_20082;
    wire new_Jinkela_wire_20560;
    wire new_Jinkela_wire_14252;
    wire new_Jinkela_wire_2519;
    wire new_Jinkela_wire_14242;
    wire new_Jinkela_wire_9500;
    wire new_Jinkela_wire_5999;
    wire new_Jinkela_wire_6401;
    wire new_Jinkela_wire_9175;
    wire new_Jinkela_wire_319;
    wire _0511_;
    wire new_Jinkela_wire_20708;
    wire new_Jinkela_wire_3708;
    wire new_Jinkela_wire_3377;
    wire new_Jinkela_wire_9581;
    wire new_Jinkela_wire_11924;
    wire new_Jinkela_wire_15528;
    wire new_Jinkela_wire_14535;
    wire new_Jinkela_wire_16526;
    wire new_Jinkela_wire_18911;
    wire new_Jinkela_wire_14766;
    wire new_Jinkela_wire_13474;
    wire new_Jinkela_wire_10030;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_12312;
    wire new_Jinkela_wire_17528;
    wire new_Jinkela_wire_5076;
    wire new_Jinkela_wire_10986;
    wire new_Jinkela_wire_19463;
    wire new_Jinkela_wire_12115;
    wire new_Jinkela_wire_11033;
    wire new_Jinkela_wire_5336;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_7977;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_6189;
    wire new_Jinkela_wire_15087;
    wire _0350_;
    wire new_Jinkela_wire_7686;
    wire _0748_;
    wire new_Jinkela_wire_18428;
    wire new_Jinkela_wire_20807;
    wire new_Jinkela_wire_18512;
    wire new_Jinkela_wire_3447;
    wire new_Jinkela_wire_15878;
    wire new_Jinkela_wire_15465;
    wire new_net_3974;
    wire new_Jinkela_wire_19526;
    wire new_Jinkela_wire_15954;
    wire new_Jinkela_wire_12120;
    wire new_Jinkela_wire_2681;
    wire new_Jinkela_wire_18963;
    wire new_Jinkela_wire_19099;
    wire new_Jinkela_wire_3404;
    wire new_Jinkela_wire_3993;
    wire new_Jinkela_wire_4343;
    wire new_Jinkela_wire_5499;
    wire new_Jinkela_wire_13684;
    wire new_Jinkela_wire_3316;
    wire new_Jinkela_wire_21067;
    wire new_Jinkela_wire_5086;
    wire new_Jinkela_wire_8489;
    wire new_Jinkela_wire_18052;
    wire new_Jinkela_wire_2079;
    wire new_Jinkela_wire_12332;
    wire new_Jinkela_wire_8770;
    wire new_Jinkela_wire_20624;
    wire new_Jinkela_wire_19170;
    wire new_Jinkela_wire_17987;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_19910;
    wire _1033_;
    wire new_Jinkela_wire_10262;
    wire new_Jinkela_wire_14655;
    wire _1690_;
    wire new_Jinkela_wire_5492;
    wire new_Jinkela_wire_7058;
    wire new_Jinkela_wire_6991;
    wire new_Jinkela_wire_15590;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_3041;
    wire new_Jinkela_wire_2882;
    wire new_Jinkela_wire_17322;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_9070;
    wire new_Jinkela_wire_10043;
    wire new_Jinkela_wire_9464;
    wire new_Jinkela_wire_8139;
    wire _0265_;
    wire new_Jinkela_wire_7550;
    wire _0885_;
    wire new_Jinkela_wire_12056;
    wire new_Jinkela_wire_8364;
    wire new_Jinkela_wire_12769;
    wire new_Jinkela_wire_13166;
    wire new_Jinkela_wire_2213;
    wire new_Jinkela_wire_2621;
    wire new_Jinkela_wire_11821;
    wire new_Jinkela_wire_19123;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_11597;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_18091;
    wire new_Jinkela_wire_6968;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_17140;
    wire new_Jinkela_wire_15041;
    wire new_Jinkela_wire_4840;
    wire new_Jinkela_wire_5132;
    wire new_Jinkela_wire_3699;
    wire new_Jinkela_wire_14665;
    wire new_Jinkela_wire_6666;
    wire new_Jinkela_wire_9441;
    wire new_Jinkela_wire_13565;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_19598;
    wire new_Jinkela_wire_19678;
    wire new_Jinkela_wire_10412;
    wire new_Jinkela_wire_3836;
    wire _1573_;
    wire new_Jinkela_wire_13471;
    wire _1163_;
    wire new_Jinkela_wire_12739;
    wire new_Jinkela_wire_10615;
    wire new_Jinkela_wire_8920;
    wire _0943_;
    wire new_Jinkela_wire_10074;
    wire new_Jinkela_wire_5188;
    wire new_Jinkela_wire_9671;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_3194;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_1643;
    wire new_Jinkela_wire_10054;
    wire new_Jinkela_wire_8946;
    wire new_Jinkela_wire_3787;
    wire new_Jinkela_wire_3508;
    wire new_Jinkela_wire_13581;
    wire new_Jinkela_wire_7618;
    wire new_Jinkela_wire_8215;
    wire new_Jinkela_wire_20417;
    wire _1574_;
    wire new_Jinkela_wire_16070;
    wire new_Jinkela_wire_3422;
    wire new_Jinkela_wire_16166;
    wire new_Jinkela_wire_17004;
    wire _1043_;
    wire new_Jinkela_wire_17521;
    wire new_Jinkela_wire_9951;
    wire _0132_;
    wire new_Jinkela_wire_14331;
    wire new_Jinkela_wire_18962;
    wire new_Jinkela_wire_12952;
    wire new_Jinkela_wire_4959;
    wire new_Jinkela_wire_11190;
    wire new_Jinkela_wire_9665;
    wire new_Jinkela_wire_8841;
    wire new_Jinkela_wire_7086;
    wire new_Jinkela_wire_18099;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_13734;
    wire new_Jinkela_wire_9518;
    wire new_Jinkela_wire_15160;
    wire new_Jinkela_wire_5208;
    wire new_Jinkela_wire_4728;
    wire new_Jinkela_wire_9475;
    wire new_Jinkela_wire_16059;
    wire _0138_;
    wire new_Jinkela_wire_12214;
    wire new_Jinkela_wire_3812;
    wire new_Jinkela_wire_19907;
    wire new_Jinkela_wire_17621;
    wire _1710_;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_12522;
    wire new_Jinkela_wire_20662;
    wire new_Jinkela_wire_6694;
    wire new_Jinkela_wire_10963;
    wire new_Jinkela_wire_3642;
    wire new_Jinkela_wire_17913;
    wire new_Jinkela_wire_7548;
    wire new_Jinkela_wire_20936;
    wire new_Jinkela_wire_10101;
    wire new_Jinkela_wire_18221;
    wire new_Jinkela_wire_13210;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_15082;
    wire new_Jinkela_wire_20530;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_3948;
    wire _0255_;
    wire _1572_;
    wire new_Jinkela_wire_19425;
    wire new_Jinkela_wire_16290;
    wire new_Jinkela_wire_9825;
    wire new_Jinkela_wire_11036;
    wire _1322_;
    wire new_Jinkela_wire_13838;
    wire new_Jinkela_wire_7294;
    wire new_Jinkela_wire_2836;
    wire new_Jinkela_wire_5870;
    wire new_Jinkela_wire_5604;
    wire new_Jinkela_wire_7835;
    wire new_Jinkela_wire_9510;
    wire new_Jinkela_wire_19954;
    wire _1578_;
    wire new_Jinkela_wire_8669;
    wire new_Jinkela_wire_18717;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_5931;
    wire new_Jinkela_wire_19308;
    wire new_Jinkela_wire_5783;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_20112;
    wire new_Jinkela_wire_16581;
    wire new_Jinkela_wire_3097;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_16930;
    wire new_Jinkela_wire_7121;
    wire new_Jinkela_wire_17435;
    wire new_Jinkela_wire_8003;
    wire new_Jinkela_wire_4113;
    wire new_Jinkela_wire_20115;
    wire new_Jinkela_wire_17730;
    wire new_Jinkela_wire_12713;
    wire new_Jinkela_wire_14848;
    wire new_Jinkela_wire_14752;
    wire _1832_;
    wire new_Jinkela_wire_14493;
    wire new_Jinkela_wire_16551;
    wire new_Jinkela_wire_6191;
    wire new_Jinkela_wire_11596;
    wire new_Jinkela_wire_16499;
    wire new_Jinkela_wire_17892;
    wire _0103_;
    wire new_Jinkela_wire_3171;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_9261;
    wire new_Jinkela_wire_19795;
    wire new_Jinkela_wire_5591;
    wire new_Jinkela_wire_4350;
    wire new_Jinkela_wire_7293;
    wire new_Jinkela_wire_10376;
    wire new_Jinkela_wire_9110;
    wire new_Jinkela_wire_13321;
    wire new_Jinkela_wire_18674;
    wire new_Jinkela_wire_13464;
    wire new_Jinkela_wire_18785;
    wire new_Jinkela_wire_15544;
    wire new_Jinkela_wire_6766;
    wire new_Jinkela_wire_14584;
    wire new_Jinkela_wire_15415;
    wire new_Jinkela_wire_14546;
    wire new_Jinkela_wire_11648;
    wire new_Jinkela_wire_7247;
    wire new_Jinkela_wire_21003;
    wire new_Jinkela_wire_13011;
    wire new_Jinkela_wire_5162;
    wire new_Jinkela_wire_1840;
    wire _0950_;
    wire new_Jinkela_wire_11050;
    wire new_Jinkela_wire_7361;
    wire new_Jinkela_wire_18748;
    wire new_Jinkela_wire_7938;
    wire new_Jinkela_wire_8518;
    wire new_Jinkela_wire_20556;
    wire new_Jinkela_wire_11427;
    wire new_Jinkela_wire_10291;
    wire new_Jinkela_wire_15860;
    wire new_Jinkela_wire_12941;
    wire new_Jinkela_wire_6964;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_19424;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_6753;
    wire new_Jinkela_wire_10984;
    wire new_Jinkela_wire_19345;
    wire _0180_;
    wire new_Jinkela_wire_2504;
    wire new_Jinkela_wire_13944;
    wire _0021_;
    wire new_Jinkela_wire_14813;
    wire new_Jinkela_wire_8746;
    wire new_Jinkela_wire_8338;
    wire _1254_;
    wire new_Jinkela_wire_11993;
    wire new_Jinkela_wire_18218;
    wire new_Jinkela_wire_4657;
    wire new_Jinkela_wire_7344;
    wire new_Jinkela_wire_4630;
    wire new_Jinkela_wire_20507;
    wire new_Jinkela_wire_5350;
    wire new_Jinkela_wire_15640;
    wire new_Jinkela_wire_10153;
    wire new_Jinkela_wire_11568;
    wire new_Jinkela_wire_4267;
    wire new_Jinkela_wire_7678;
    wire new_Jinkela_wire_17225;
    wire new_Jinkela_wire_4563;
    wire new_Jinkela_wire_18414;
    wire new_Jinkela_wire_15607;
    wire new_Jinkela_wire_15437;
    wire new_Jinkela_wire_19395;
    wire new_Jinkela_wire_3326;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_2225;
    wire new_Jinkela_wire_16406;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_5628;
    wire new_Jinkela_wire_11980;
    wire new_Jinkela_wire_19588;
    wire new_Jinkela_wire_20185;
    wire new_Jinkela_wire_19407;
    wire new_Jinkela_wire_6814;
    wire new_Jinkela_wire_4479;
    wire new_Jinkela_wire_19413;
    wire new_Jinkela_wire_13652;
    wire new_Jinkela_wire_20116;
    wire new_Jinkela_wire_7412;
    wire new_Jinkela_wire_18516;
    wire new_Jinkela_wire_13380;
    wire new_Jinkela_wire_14222;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_12753;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_13841;
    wire new_Jinkela_wire_3416;
    wire new_Jinkela_wire_3591;
    wire new_Jinkela_wire_18766;
    wire new_Jinkela_wire_11109;
    wire new_Jinkela_wire_2885;
    wire new_Jinkela_wire_21150;
    wire new_Jinkela_wire_15559;
    wire new_Jinkela_wire_13593;
    wire new_Jinkela_wire_15615;
    wire new_Jinkela_wire_2013;
    wire new_Jinkela_wire_10997;
    wire new_Jinkela_wire_17319;
    wire new_Jinkela_wire_15285;
    wire new_Jinkela_wire_1823;
    wire _1634_;
    wire new_Jinkela_wire_6754;
    wire new_Jinkela_wire_8162;
    wire new_Jinkela_wire_18146;
    wire new_Jinkela_wire_10328;
    wire new_Jinkela_wire_6477;
    wire new_Jinkela_wire_7118;
    wire new_Jinkela_wire_18912;
    wire new_Jinkela_wire_20996;
    wire new_Jinkela_wire_18465;
    wire new_Jinkela_wire_11346;
    wire new_Jinkela_wire_19814;
    wire new_Jinkela_wire_21310;
    wire new_Jinkela_wire_13466;
    wire new_Jinkela_wire_4500;
    wire new_Jinkela_wire_16920;
    wire _0472_;
    wire new_Jinkela_wire_18783;
    wire new_Jinkela_wire_17028;
    wire new_Jinkela_wire_5672;
    wire new_Jinkela_wire_5634;
    wire new_Jinkela_wire_3648;
    wire new_Jinkela_wire_14468;
    wire new_Jinkela_wire_17766;
    wire new_Jinkela_wire_4380;
    wire new_Jinkela_wire_8303;
    wire new_Jinkela_wire_15626;
    wire new_Jinkela_wire_14720;
    wire new_Jinkela_wire_16209;
    wire new_Jinkela_wire_15713;
    wire new_Jinkela_wire_14770;
    wire new_Jinkela_wire_9861;
    wire new_Jinkela_wire_9944;
    wire new_Jinkela_wire_10544;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_7585;
    wire new_Jinkela_wire_5642;
    wire new_Jinkela_wire_6479;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_20520;
    wire new_Jinkela_wire_13874;
    wire new_Jinkela_wire_2368;
    wire new_Jinkela_wire_19466;
    wire new_Jinkela_wire_3435;
    wire new_Jinkela_wire_2309;
    wire new_Jinkela_wire_10867;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_4206;
    wire new_Jinkela_wire_14940;
    wire new_Jinkela_wire_10726;
    wire new_Jinkela_wire_16355;
    wire new_Jinkela_wire_8837;
    wire new_Jinkela_wire_10016;
    wire new_Jinkela_wire_12086;
    wire new_Jinkela_wire_3747;
    wire new_Jinkela_wire_6381;
    wire new_Jinkela_wire_21000;
    wire new_Jinkela_wire_8337;
    wire new_Jinkela_wire_13194;
    wire new_Jinkela_wire_11917;
    wire new_Jinkela_wire_7623;
    wire new_Jinkela_wire_7273;
    wire new_Jinkela_wire_17037;
    wire new_Jinkela_wire_14321;
    wire _0610_;
    wire new_Jinkela_wire_13322;
    wire _1706_;
    wire new_Jinkela_wire_14367;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_3726;
    wire new_Jinkela_wire_3569;
    wire new_Jinkela_wire_4020;
    wire _1281_;
    wire _1109_;
    wire new_Jinkela_wire_678;
    wire _0835_;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_16306;
    wire _1228_;
    wire new_Jinkela_wire_3181;
    wire new_Jinkela_wire_10886;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_9497;
    wire new_Jinkela_wire_5789;
    wire new_Jinkela_wire_12270;
    wire new_Jinkela_wire_12349;
    wire new_Jinkela_wire_5530;
    wire new_Jinkela_wire_2577;
    wire new_Jinkela_wire_16866;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_5757;
    wire new_Jinkela_wire_8454;
    wire new_Jinkela_wire_15364;
    wire new_Jinkela_wire_4848;
    wire new_Jinkela_wire_17793;
    wire new_Jinkela_wire_12033;
    wire new_Jinkela_wire_19719;
    wire new_Jinkela_wire_13241;
    wire new_Jinkela_wire_21120;
    wire new_Jinkela_wire_7789;
    wire new_Jinkela_wire_7191;
    wire new_Jinkela_wire_15887;
    wire _0108_;
    wire new_Jinkela_wire_3745;
    wire new_Jinkela_wire_8317;
    wire new_Jinkela_wire_6442;
    wire new_Jinkela_wire_14561;
    wire new_Jinkela_wire_17260;
    wire new_Jinkela_wire_16614;
    wire new_Jinkela_wire_13616;
    wire new_Jinkela_wire_6700;
    wire new_Jinkela_wire_12542;
    wire new_Jinkela_wire_18972;
    wire new_Jinkela_wire_16636;
    wire new_Jinkela_wire_8728;
    wire _1288_;
    wire new_Jinkela_wire_17717;
    wire new_Jinkela_wire_5979;
    wire new_Jinkela_wire_16419;
    wire new_Jinkela_wire_18224;
    wire new_Jinkela_wire_3821;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_7112;
    wire new_Jinkela_wire_20810;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_3906;
    wire new_Jinkela_wire_4714;
    wire new_Jinkela_wire_12849;
    wire new_Jinkela_wire_6640;
    wire new_Jinkela_wire_10280;
    wire new_Jinkela_wire_8641;
    wire new_Jinkela_wire_7125;
    wire new_Jinkela_wire_15853;
    wire new_Jinkela_wire_8983;
    wire new_Jinkela_wire_7753;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_20496;
    wire new_Jinkela_wire_3469;
    wire _1542_;
    wire new_Jinkela_wire_5816;
    wire new_Jinkela_wire_5466;
    wire new_Jinkela_wire_18455;
    wire new_Jinkela_wire_11022;
    wire new_Jinkela_wire_20886;
    wire new_Jinkela_wire_19331;
    wire _0692_;
    wire new_Jinkela_wire_6322;
    wire new_Jinkela_wire_19059;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_8512;
    wire new_Jinkela_wire_18060;
    wire new_Jinkela_wire_19271;
    wire new_Jinkela_wire_10678;
    wire new_Jinkela_wire_2275;
    wire new_Jinkela_wire_5668;
    wire new_Jinkela_wire_1234;
    wire _0879_;
    wire new_Jinkela_wire_4570;
    wire new_Jinkela_wire_4524;
    wire new_Jinkela_wire_2542;
    wire new_Jinkela_wire_18170;
    wire new_Jinkela_wire_11976;
    wire new_Jinkela_wire_7452;
    wire new_Jinkela_wire_14444;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_17704;
    wire new_Jinkela_wire_7776;
    wire new_Jinkela_wire_6764;
    wire _1156_;
    wire new_Jinkela_wire_8473;
    wire new_Jinkela_wire_19278;
    wire new_Jinkela_wire_10335;
    wire new_Jinkela_wire_8740;
    wire new_Jinkela_wire_4653;
    wire new_Jinkela_wire_10819;
    wire new_Jinkela_wire_18916;
    wire new_Jinkela_wire_12152;
    wire new_Jinkela_wire_19744;
    wire new_Jinkela_wire_8273;
    wire new_Jinkela_wire_7626;
    wire new_Jinkela_wire_8216;
    wire new_Jinkela_wire_20992;
    wire new_Jinkela_wire_13901;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_14687;
    wire new_Jinkela_wire_4450;
    wire new_Jinkela_wire_11037;
    wire new_Jinkela_wire_20362;
    wire new_Jinkela_wire_16026;
    wire new_Jinkela_wire_10607;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_12732;
    wire new_Jinkela_wire_14359;
    wire new_Jinkela_wire_12444;
    wire _1321_;
    wire new_Jinkela_wire_11672;
    wire new_Jinkela_wire_5494;
    wire new_Jinkela_wire_18795;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_4945;
    wire new_Jinkela_wire_2956;
    wire new_Jinkela_wire_2967;
    wire new_Jinkela_wire_9868;
    wire new_Jinkela_wire_14731;
    wire new_Jinkela_wire_11723;
    wire new_Jinkela_wire_1696;
    wire _0559_;
    wire new_Jinkela_wire_2131;
    wire new_Jinkela_wire_19698;
    wire new_Jinkela_wire_14399;
    wire new_Jinkela_wire_17658;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_15527;
    wire new_Jinkela_wire_18915;
    wire new_Jinkela_wire_11879;
    wire new_Jinkela_wire_4466;
    wire new_Jinkela_wire_13485;
    wire new_Jinkela_wire_15502;
    wire new_Jinkela_wire_16927;
    wire new_Jinkela_wire_16466;
    wire new_Jinkela_wire_7609;
    wire new_Jinkela_wire_15927;
    wire new_Jinkela_wire_7392;
    wire new_Jinkela_wire_4791;
    wire new_Jinkela_wire_2220;
    wire new_Jinkela_wire_16671;
    wire new_Jinkela_wire_15346;
    wire new_Jinkela_wire_20962;
    wire new_Jinkela_wire_13793;
    wire new_Jinkela_wire_5229;
    wire new_Jinkela_wire_2458;
    wire new_Jinkela_wire_8795;
    wire new_Jinkela_wire_20703;
    wire new_Jinkela_wire_2202;
    wire new_Jinkela_wire_10462;
    wire new_Jinkela_wire_7127;
    wire new_Jinkela_wire_9881;
    wire new_Jinkela_wire_16555;
    wire new_Jinkela_wire_20610;
    wire new_Jinkela_wire_18320;
    wire new_Jinkela_wire_3162;
    wire new_Jinkela_wire_3761;
    wire new_Jinkela_wire_8918;
    wire new_Jinkela_wire_20005;
    wire new_Jinkela_wire_15260;
    wire new_Jinkela_wire_14876;
    wire _0437_;
    wire new_Jinkela_wire_6443;
    wire new_Jinkela_wire_6090;
    wire new_Jinkela_wire_9425;
    wire new_Jinkela_wire_13074;
    wire new_Jinkela_wire_9908;
    wire new_Jinkela_wire_2883;
    wire new_Jinkela_wire_2769;
    wire new_Jinkela_wire_13957;
    wire new_Jinkela_wire_2799;
    wire new_Jinkela_wire_5448;
    wire new_Jinkela_wire_12154;
    wire new_Jinkela_wire_8336;
    wire new_Jinkela_wire_8053;
    wire _0734_;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_8496;
    wire new_Jinkela_wire_20902;
    wire new_Jinkela_wire_7803;
    wire new_Jinkela_wire_17213;
    wire new_Jinkela_wire_15597;
    wire new_Jinkela_wire_13672;
    wire new_Jinkela_wire_3107;
    wire new_Jinkela_wire_14677;
    wire new_Jinkela_wire_14293;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_8236;
    wire new_Jinkela_wire_5539;
    wire new_Jinkela_wire_10495;
    wire new_Jinkela_wire_18026;
    wire new_Jinkela_wire_9910;
    wire new_Jinkela_wire_8184;
    wire new_Jinkela_wire_4459;
    wire new_Jinkela_wire_18547;
    wire new_Jinkela_wire_5533;
    wire new_Jinkela_wire_14635;
    wire new_Jinkela_wire_16437;
    wire new_Jinkela_wire_18845;
    wire new_Jinkela_wire_3543;
    wire new_Jinkela_wire_3910;
    wire new_Jinkela_wire_5926;
    wire new_Jinkela_wire_5652;
    wire new_Jinkela_wire_6276;
    wire new_Jinkela_wire_5082;
    wire new_Jinkela_wire_4517;
    wire new_Jinkela_wire_16304;
    wire new_Jinkela_wire_15899;
    wire new_Jinkela_wire_9746;
    wire new_Jinkela_wire_7416;
    wire new_Jinkela_wire_4937;
    wire new_Jinkela_wire_19436;
    wire new_Jinkela_wire_2126;
    wire new_Jinkela_wire_14101;
    wire new_Jinkela_wire_1398;
    wire new_Jinkela_wire_13314;
    wire _0798_;
    wire new_Jinkela_wire_17744;
    wire new_Jinkela_wire_16843;
    wire new_Jinkela_wire_20629;
    wire new_Jinkela_wire_20093;
    wire new_Jinkela_wire_18458;
    wire new_Jinkela_wire_9033;
    wire new_Jinkela_wire_1437;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_2942;
    wire new_Jinkela_wire_3892;
    wire new_Jinkela_wire_16287;
    wire new_Jinkela_wire_10571;
    wire new_Jinkela_wire_5081;
    wire new_Jinkela_wire_19093;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_13877;
    wire new_Jinkela_wire_2678;
    wire new_Jinkela_wire_2322;
    wire new_Jinkela_wire_18003;
    wire new_Jinkela_wire_16360;
    wire new_Jinkela_wire_4655;
    wire new_Jinkela_wire_14533;
    wire new_Jinkela_wire_9841;
    wire new_Jinkela_wire_14930;
    wire _0106_;
    wire new_Jinkela_wire_3738;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_20397;
    wire new_Jinkela_wire_2827;
    wire new_Jinkela_wire_16000;
    wire new_Jinkela_wire_8092;
    wire new_Jinkela_wire_1093;
    wire new_Jinkela_wire_19773;
    wire new_Jinkela_wire_3719;
    wire _0937_;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_3471;
    wire new_Jinkela_wire_1390;
    wire _0340_;
    wire new_Jinkela_wire_12476;
    wire new_Jinkela_wire_12301;
    wire new_Jinkela_wire_10692;
    wire new_Jinkela_wire_4898;
    wire new_Jinkela_wire_4334;
    wire _0310_;
    wire new_Jinkela_wire_17369;
    wire new_Jinkela_wire_19845;
    wire new_Jinkela_wire_3170;
    wire new_Jinkela_wire_4967;
    wire new_Jinkela_wire_9850;
    wire new_Jinkela_wire_11040;
    wire new_Jinkela_wire_18575;
    wire new_Jinkela_wire_9039;
    wire new_Jinkela_wire_12764;
    wire new_Jinkela_wire_7610;
    wire new_Jinkela_wire_14652;
    wire new_Jinkela_wire_14983;
    wire new_Jinkela_wire_12425;
    wire new_Jinkela_wire_10609;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_9827;
    wire new_Jinkela_wire_12989;
    wire new_Jinkela_wire_20328;
    wire new_Jinkela_wire_15770;
    wire new_Jinkela_wire_10112;
    wire new_Jinkela_wire_11104;
    wire new_Jinkela_wire_12340;
    wire new_Jinkela_wire_6951;
    wire new_Jinkela_wire_13442;
    wire new_Jinkela_wire_17111;
    wire new_Jinkela_wire_2797;
    wire new_Jinkela_wire_12400;
    wire new_Jinkela_wire_8738;
    wire new_Jinkela_wire_11529;
    wire new_Jinkela_wire_13387;
    wire new_Jinkela_wire_8305;
    wire new_Jinkela_wire_20640;
    wire new_Jinkela_wire_13351;
    wire new_Jinkela_wire_3476;
    wire new_Jinkela_wire_7807;
    wire new_Jinkela_wire_19609;
    wire new_Jinkela_wire_1156;
    wire _1247_;
    wire new_Jinkela_wire_14662;
    wire new_Jinkela_wire_18969;
    wire new_Jinkela_wire_8164;
    wire new_Jinkela_wire_3514;
    wire new_Jinkela_wire_10550;
    wire new_Jinkela_wire_14633;
    wire new_Jinkela_wire_11116;
    wire new_Jinkela_wire_6793;
    wire new_Jinkela_wire_4692;
    wire new_Jinkela_wire_5574;
    wire new_Jinkela_wire_8528;
    wire new_Jinkela_wire_15619;
    wire new_Jinkela_wire_6823;
    wire new_Jinkela_wire_17296;
    wire new_Jinkela_wire_21321;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_6355;
    wire new_Jinkela_wire_16234;
    wire new_Jinkela_wire_10063;
    wire _1270_;
    wire new_Jinkela_wire_13075;
    wire _0652_;
    wire new_Jinkela_wire_13534;
    wire new_Jinkela_wire_7120;
    wire new_Jinkela_wire_12835;
    wire new_Jinkela_wire_7825;
    wire new_Jinkela_wire_8210;
    wire new_Jinkela_wire_18743;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_19939;
    wire new_Jinkela_wire_18181;
    wire new_Jinkela_wire_3885;
    wire new_Jinkela_wire_16481;
    wire new_Jinkela_wire_5427;
    wire new_Jinkela_wire_12222;
    wire new_Jinkela_wire_6101;
    wire new_Jinkela_wire_15147;
    wire new_Jinkela_wire_12704;
    wire new_Jinkela_wire_14756;
    wire new_Jinkela_wire_2830;
    wire new_Jinkela_wire_11258;
    wire new_Jinkela_wire_7660;
    wire _1560_;
    wire new_Jinkela_wire_3974;
    wire new_Jinkela_wire_16016;
    wire new_Jinkela_wire_3798;
    wire new_Jinkela_wire_6130;
    wire new_Jinkela_wire_1145;
    wire new_Jinkela_wire_20574;
    wire new_Jinkela_wire_14747;
    wire new_Jinkela_wire_2690;
    wire new_Jinkela_wire_19021;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_16270;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_6687;
    wire new_Jinkela_wire_2686;
    wire new_Jinkela_wire_3415;
    wire new_Jinkela_wire_6565;
    wire new_Jinkela_wire_18303;
    wire new_Jinkela_wire_7085;
    wire new_Jinkela_wire_3441;
    wire new_Jinkela_wire_10546;
    wire new_Jinkela_wire_6473;
    wire new_Jinkela_wire_16548;
    wire new_Jinkela_wire_11968;
    wire new_Jinkela_wire_10145;
    wire new_Jinkela_wire_4723;
    wire new_Jinkela_wire_12127;
    wire new_Jinkela_wire_6109;
    wire new_Jinkela_wire_15312;
    wire new_Jinkela_wire_14413;
    wire new_Jinkela_wire_13344;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_20647;
    wire new_Jinkela_wire_19824;
    wire new_Jinkela_wire_8;
    wire _0751_;
    wire new_Jinkela_wire_2459;
    wire new_Jinkela_wire_1874;
    wire new_Jinkela_wire_5252;
    wire new_Jinkela_wire_16872;
    wire _0723_;
    wire new_Jinkela_wire_14464;
    wire new_Jinkela_wire_4560;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_11152;
    wire new_Jinkela_wire_8595;
    wire new_Jinkela_wire_6303;
    wire new_Jinkela_wire_7672;
    wire new_Jinkela_wire_14204;
    wire new_Jinkela_wire_12180;
    wire new_Jinkela_wire_19673;
    wire _0170_;
    wire new_Jinkela_wire_15655;
    wire _0453_;
    wire new_Jinkela_wire_11780;
    wire _1328_;
    wire new_Jinkela_wire_6668;
    wire new_Jinkela_wire_9225;
    wire new_Jinkela_wire_6949;
    wire new_Jinkela_wire_4932;
    wire new_Jinkela_wire_15797;
    wire new_Jinkela_wire_21121;
    wire new_Jinkela_wire_5839;
    wire new_Jinkela_wire_7710;
    wire new_Jinkela_wire_5606;
    wire new_Jinkela_wire_16274;
    wire new_Jinkela_wire_10784;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_2271;
    wire new_Jinkela_wire_10987;
    wire new_Jinkela_wire_17656;
    wire new_Jinkela_wire_4407;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_7442;
    wire new_Jinkela_wire_11776;
    wire new_Jinkela_wire_12051;
    wire new_Jinkela_wire_9766;
    wire _1148_;
    wire new_Jinkela_wire_20001;
    wire new_Jinkela_wire_15730;
    wire new_Jinkela_wire_5648;
    wire new_Jinkela_wire_10800;
    wire new_Jinkela_wire_17933;
    wire new_Jinkela_wire_17628;
    wire _0362_;
    wire new_Jinkela_wire_15941;
    wire new_Jinkela_wire_18814;
    wire new_Jinkela_wire_11769;
    wire new_Jinkela_wire_16532;
    wire new_Jinkela_wire_20713;
    wire new_Jinkela_wire_18710;
    wire new_Jinkela_wire_18588;
    wire new_Jinkela_wire_17114;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_12204;
    wire new_Jinkela_wire_11826;
    wire new_Jinkela_wire_7356;
    wire new_Jinkela_wire_12714;
    wire new_Jinkela_wire_3505;
    wire new_Jinkela_wire_13022;
    wire new_Jinkela_wire_2435;
    wire new_Jinkela_wire_6543;
    wire new_Jinkela_wire_12137;
    wire new_Jinkela_wire_14138;
    wire new_Jinkela_wire_10504;
    wire new_Jinkela_wire_13656;
    wire new_Jinkela_wire_17484;
    wire _0921_;
    wire new_Jinkela_wire_20601;
    wire new_Jinkela_wire_20521;
    wire new_Jinkela_wire_8929;
    wire new_Jinkela_wire_11112;
    wire new_Jinkela_wire_6256;
    wire new_Jinkela_wire_2579;
    wire new_Jinkela_wire_16658;
    wire new_Jinkela_wire_10834;
    wire new_Jinkela_wire_13235;
    wire new_Jinkela_wire_15009;
    wire new_Jinkela_wire_15801;
    wire new_Jinkela_wire_11147;
    wire new_Jinkela_wire_16867;
    wire new_Jinkela_wire_2075;
    wire _1568_;
    wire new_Jinkela_wire_15654;
    wire new_Jinkela_wire_4408;
    wire new_Jinkela_wire_19512;
    wire new_Jinkela_wire_20006;
    wire _0115_;
    wire new_Jinkela_wire_7775;
    wire _0687_;
    wire new_Jinkela_wire_19013;
    wire new_Jinkela_wire_18309;
    wire _0942_;
    wire new_Jinkela_wire_13826;
    wire _0176_;
    wire new_Jinkela_wire_15368;
    wire new_Jinkela_wire_5497;
    wire new_Jinkela_wire_5308;
    wire new_Jinkela_wire_9103;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_4223;
    wire new_Jinkela_wire_7040;
    wire new_Jinkela_wire_11336;
    wire _0948_;
    wire new_Jinkela_wire_17815;
    wire new_Jinkela_wire_14027;
    wire new_Jinkela_wire_17193;
    wire new_Jinkela_wire_10918;
    wire new_Jinkela_wire_18470;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_9161;
    wire new_Jinkela_wire_13047;
    wire new_Jinkela_wire_17824;
    wire new_Jinkela_wire_6081;
    wire new_Jinkela_wire_2765;
    wire new_Jinkela_wire_8430;
    wire new_Jinkela_wire_615;
    wire _0930_;
    wire new_Jinkela_wire_18464;
    wire new_Jinkela_wire_8418;
    wire new_Jinkela_wire_18606;
    wire new_Jinkela_wire_13012;
    wire new_Jinkela_wire_2349;
    wire _1507_;
    wire new_Jinkela_wire_6328;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_11567;
    wire new_Jinkela_wire_5559;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_19316;
    wire new_Jinkela_wire_5483;
    wire new_Jinkela_wire_10551;
    wire _1769_;
    wire new_Jinkela_wire_6249;
    wire new_Jinkela_wire_6537;
    wire new_Jinkela_wire_16164;
    wire new_Jinkela_wire_6421;
    wire new_Jinkela_wire_10846;
    wire _0422_;
    wire _0338_;
    wire new_Jinkela_wire_6563;
    wire new_Jinkela_wire_2532;
    wire new_Jinkela_wire_7625;
    wire new_Jinkela_wire_10924;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_7899;
    wire new_Jinkela_wire_4160;
    wire new_Jinkela_wire_20049;
    wire new_Jinkela_wire_18094;
    wire new_Jinkela_wire_4502;
    wire new_Jinkela_wire_15729;
    wire new_Jinkela_wire_7978;
    wire new_Jinkela_wire_11317;
    wire new_Jinkela_wire_12318;
    wire new_Jinkela_wire_2671;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_13021;
    wire new_Jinkela_wire_3100;
    wire new_Jinkela_wire_19993;
    wire new_Jinkela_wire_4321;
    wire new_Jinkela_wire_7931;
    wire new_Jinkela_wire_2289;
    wire new_Jinkela_wire_9932;
    wire new_Jinkela_wire_13311;
    wire new_Jinkela_wire_20947;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_9794;
    wire new_Jinkela_wire_9681;
    wire new_Jinkela_wire_16836;
    wire new_Jinkela_wire_21243;
    wire new_Jinkela_wire_3678;
    wire _0826_;
    wire new_Jinkela_wire_12665;
    wire new_Jinkela_wire_20841;
    wire new_Jinkela_wire_12502;
    wire new_Jinkela_wire_2677;
    wire new_Jinkela_wire_9546;
    wire new_Jinkela_wire_8243;
    wire new_Jinkela_wire_11745;
    wire new_Jinkela_wire_9852;
    wire new_Jinkela_wire_14802;
    wire new_Jinkela_wire_19392;
    wire new_Jinkela_wire_9992;
    wire _0447_;
    wire new_Jinkela_wire_19513;
    wire new_Jinkela_wire_8294;
    wire new_Jinkela_wire_7053;
    wire new_Jinkela_wire_13891;
    wire new_Jinkela_wire_5118;
    wire new_Jinkela_wire_3270;
    wire new_Jinkela_wire_18923;
    wire _1303_;
    wire new_Jinkela_wire_18689;
    wire new_Jinkela_wire_2513;
    wire new_Jinkela_wire_8707;
    wire new_Jinkela_wire_10021;
    wire new_Jinkela_wire_1963;
    wire new_Jinkela_wire_11067;
    wire new_Jinkela_wire_8131;
    wire _1393_;
    wire _0520_;
    wire _1498_;
    wire new_Jinkela_wire_17289;
    wire new_Jinkela_wire_11402;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_8407;
    wire new_Jinkela_wire_8874;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_14088;
    wire new_Jinkela_wire_20064;
    wire new_Jinkela_wire_7935;
    wire new_Jinkela_wire_11151;
    wire new_Jinkela_wire_3018;
    wire new_Jinkela_wire_3006;
    wire new_Jinkela_wire_16748;
    wire new_Jinkela_wire_13743;
    wire new_Jinkela_wire_15843;
    wire new_Jinkela_wire_20571;
    wire new_Jinkela_wire_16004;
    wire new_Jinkela_wire_4850;
    wire new_Jinkela_wire_16291;
    wire new_Jinkela_wire_20653;
    wire _1091_;
    wire new_Jinkela_wire_16660;
    wire new_Jinkela_wire_19691;
    wire new_Jinkela_wire_2434;
    wire new_Jinkela_wire_15301;
    wire new_Jinkela_wire_15919;
    wire new_Jinkela_wire_18685;
    wire new_Jinkela_wire_14309;
    wire new_Jinkela_wire_4365;
    wire new_Jinkela_wire_1137;
    wire new_Jinkela_wire_10426;
    wire new_Jinkela_wire_10979;
    wire new_Jinkela_wire_13726;
    wire new_Jinkela_wire_6651;
    wire new_Jinkela_wire_12087;
    wire new_Jinkela_wire_2996;
    wire new_Jinkela_wire_11737;
    wire new_Jinkela_wire_17274;
    wire new_Jinkela_wire_2326;
    wire new_Jinkela_wire_18586;
    wire new_Jinkela_wire_6332;
    wire new_Jinkela_wire_6188;
    wire new_Jinkela_wire_6804;
    wire new_Jinkela_wire_20466;
    wire new_Jinkela_wire_20837;
    wire _0030_;
    wire new_Jinkela_wire_3239;
    wire new_Jinkela_wire_4545;
    wire new_Jinkela_wire_4579;
    wire new_Jinkela_wire_12863;
    wire new_Jinkela_wire_16045;
    wire new_Jinkela_wire_4796;
    wire new_Jinkela_wire_20775;
    wire new_Jinkela_wire_6874;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_12720;
    wire new_Jinkela_wire_4511;
    wire new_Jinkela_wire_10807;
    wire new_Jinkela_wire_8987;
    wire new_Jinkela_wire_16860;
    wire new_Jinkela_wire_15257;
    wire new_Jinkela_wire_11068;
    wire new_Jinkela_wire_1478;
    wire _1130_;
    wire new_Jinkela_wire_14503;
    wire new_Jinkela_wire_15416;
    wire new_Jinkela_wire_17750;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_19040;
    wire new_Jinkela_wire_21026;
    wire new_Jinkela_wire_1806;
    wire new_Jinkela_wire_7979;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_20598;
    wire new_Jinkela_wire_5719;
    wire new_Jinkela_wire_19236;
    wire new_Jinkela_wire_6458;
    wire new_Jinkela_wire_19629;
    wire new_Jinkela_wire_1724;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_6074;
    wire new_Jinkela_wire_16910;
    wire new_Jinkela_wire_16470;
    wire new_Jinkela_wire_8090;
    wire new_Jinkela_wire_8349;
    wire new_Jinkela_wire_13869;
    wire new_Jinkela_wire_18366;
    wire new_Jinkela_wire_4127;
    wire new_Jinkela_wire_8872;
    wire new_Jinkela_wire_8017;
    wire _1798_;
    wire new_Jinkela_wire_12741;
    wire new_Jinkela_wire_16146;
    wire _1144_;
    wire new_Jinkela_wire_15775;
    wire new_Jinkela_wire_15576;
    wire _1421_;
    wire new_Jinkela_wire_9638;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_10533;
    wire new_Jinkela_wire_7539;
    wire new_Jinkela_wire_8280;
    wire new_Jinkela_wire_16089;
    wire new_Jinkela_wire_19250;
    wire new_Jinkela_wire_17368;
    wire new_Jinkela_wire_17445;
    wire new_Jinkela_wire_6013;
    wire _0900_;
    wire new_Jinkela_wire_2199;
    wire new_Jinkela_wire_2635;
    wire new_Jinkela_wire_4946;
    wire new_Jinkela_wire_17622;
    wire new_Jinkela_wire_6029;
    wire new_Jinkela_wire_12619;
    wire new_Jinkela_wire_6277;
    wire new_Jinkela_wire_12667;
    wire new_Jinkela_wire_11654;
    wire new_Jinkela_wire_11319;
    wire new_Jinkela_wire_2190;
    wire _1804_;
    wire new_Jinkela_wire_12611;
    wire new_Jinkela_wire_7841;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_19877;
    wire _1319_;
    wire new_Jinkela_wire_14107;
    wire new_Jinkela_wire_20786;
    wire new_Jinkela_wire_16992;
    wire new_Jinkela_wire_14575;
    wire new_Jinkela_wire_7324;
    wire new_Jinkela_wire_17458;
    wire new_Jinkela_wire_9396;
    wire new_Jinkela_wire_1856;
    wire new_Jinkela_wire_16959;
    wire new_Jinkela_wire_15891;
    wire _1516_;
    wire new_Jinkela_wire_6945;
    wire new_Jinkela_wire_20517;
    wire new_Jinkela_wire_8498;
    wire new_Jinkela_wire_16585;
    wire new_Jinkela_wire_6482;
    wire new_Jinkela_wire_16246;
    wire new_Jinkela_wire_14708;
    wire new_Jinkela_wire_20695;
    wire new_Jinkela_wire_12176;
    wire new_Jinkela_wire_14729;
    wire new_Jinkela_wire_10324;
    wire _1396_;
    wire new_Jinkela_wire_8973;
    wire new_Jinkela_wire_5102;
    wire new_Jinkela_wire_1627;
    wire new_Jinkela_wire_10642;
    wire new_Jinkela_wire_9573;
    wire new_Jinkela_wire_10691;
    wire new_Jinkela_wire_8957;
    wire new_Jinkela_wire_10688;
    wire new_Jinkela_wire_6419;
    wire new_Jinkela_wire_9303;
    wire new_Jinkela_wire_14214;
    wire new_Jinkela_wire_20249;
    wire new_Jinkela_wire_5109;
    wire new_Jinkela_wire_7767;
    wire new_Jinkela_wire_14481;
    wire new_Jinkela_wire_3662;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_17948;
    wire new_Jinkela_wire_11500;
    wire new_Jinkela_wire_18199;
    wire new_Jinkela_wire_7491;
    wire new_Jinkela_wire_14369;
    wire new_Jinkela_wire_21196;
    wire new_Jinkela_wire_6423;
    wire new_Jinkela_wire_12894;
    wire new_Jinkela_wire_10017;
    wire new_Jinkela_wire_9655;
    wire new_Jinkela_wire_1405;
    wire new_Jinkela_wire_5091;
    wire new_Jinkela_wire_9678;
    wire new_Jinkela_wire_11128;
    wire new_Jinkela_wire_10486;
    wire new_Jinkela_wire_21173;
    wire new_Jinkela_wire_9646;
    wire new_Jinkela_wire_15599;
    wire new_Jinkela_wire_2089;
    wire new_Jinkela_wire_4456;
    wire new_Jinkela_wire_6137;
    wire new_Jinkela_wire_18128;
    wire new_Jinkela_wire_14572;
    wire new_Jinkela_wire_5566;
    wire new_Jinkela_wire_19419;
    wire new_Jinkela_wire_10823;
    wire new_Jinkela_wire_15854;
    wire new_Jinkela_wire_19803;
    wire new_Jinkela_wire_16565;
    wire new_Jinkela_wire_20299;
    wire new_Jinkela_wire_19442;
    wire new_Jinkela_wire_20031;
    wire new_Jinkela_wire_15568;
    wire new_Jinkela_wire_15235;
    wire new_Jinkela_wire_10448;
    wire new_Jinkela_wire_20767;
    wire new_Jinkela_wire_12191;
    wire new_Jinkela_wire_11505;
    wire new_Jinkela_wire_16484;
    wire new_Jinkela_wire_7826;
    wire new_Jinkela_wire_10493;
    wire new_Jinkela_wire_9471;
    wire new_Jinkela_wire_14539;
    wire new_Jinkela_wire_12814;
    wire new_Jinkela_wire_16172;
    wire new_Jinkela_wire_13664;
    wire new_Jinkela_wire_3932;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_18715;
    wire new_Jinkela_wire_2037;
    wire new_Jinkela_wire_20914;
    wire new_Jinkela_wire_5963;
    wire new_Jinkela_wire_15311;
    wire new_Jinkela_wire_3069;
    wire new_Jinkela_wire_14829;
    wire new_Jinkela_wire_10673;
    wire new_Jinkela_wire_11014;
    wire new_Jinkela_wire_7463;
    wire new_Jinkela_wire_12800;
    wire new_Jinkela_wire_10360;
    wire new_Jinkela_wire_11254;
    wire new_Jinkela_wire_14245;
    wire new_Jinkela_wire_17994;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_16227;
    wire new_Jinkela_wire_13959;
    wire new_Jinkela_wire_8434;
    wire new_Jinkela_wire_7645;
    wire new_Jinkela_wire_6012;
    wire new_Jinkela_wire_18140;
    wire new_Jinkela_wire_20787;
    wire _1173_;
    wire new_Jinkela_wire_10895;
    wire new_Jinkela_wire_10257;
    wire new_Jinkela_wire_19232;
    wire new_Jinkela_wire_8878;
    wire new_Jinkela_wire_14037;
    wire new_Jinkela_wire_19656;
    wire new_Jinkela_wire_21218;
    wire new_Jinkela_wire_7663;
    wire new_Jinkela_wire_2904;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_12794;
    wire new_Jinkela_wire_8070;
    wire new_Jinkela_wire_16656;
    wire new_Jinkela_wire_10306;
    wire new_Jinkela_wire_16486;
    wire new_Jinkela_wire_9626;
    wire _1694_;
    wire new_Jinkela_wire_21312;
    wire _1280_;
    wire new_Jinkela_wire_9964;
    wire new_Jinkela_wire_19854;
    wire new_Jinkela_wire_3824;
    wire new_Jinkela_wire_14972;
    wire new_Jinkela_wire_17011;
    wire _0206_;
    wire new_Jinkela_wire_13648;
    wire new_Jinkela_wire_11186;
    wire new_Jinkela_wire_8680;
    wire new_Jinkela_wire_18971;
    wire new_Jinkela_wire_5039;
    wire new_Jinkela_wire_2110;
    wire new_Jinkela_wire_13204;
    wire new_Jinkela_wire_6483;
    wire new_Jinkela_wire_18677;
    wire new_Jinkela_wire_7597;
    wire new_Jinkela_wire_5573;
    wire new_Jinkela_wire_2804;
    wire new_Jinkela_wire_13812;
    wire _1422_;
    wire new_Jinkela_wire_7290;
    wire new_Jinkela_wire_9147;
    wire new_Jinkela_wire_11753;
    wire new_Jinkela_wire_5525;
    wire new_Jinkela_wire_20828;
    wire new_Jinkela_wire_15417;
    wire new_Jinkela_wire_11096;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_15243;
    wire new_Jinkela_wire_15858;
    wire new_Jinkela_wire_8323;
    wire new_Jinkela_wire_1871;
    wire new_Jinkela_wire_11713;
    wire new_Jinkela_wire_8196;
    wire _0707_;
    wire new_Jinkela_wire_4578;
    wire new_Jinkela_wire_17734;
    wire new_Jinkela_wire_14918;
    wire new_Jinkela_wire_17153;
    wire new_Jinkela_wire_6735;
    wire new_Jinkela_wire_18735;
    wire new_Jinkela_wire_3991;
    wire new_Jinkela_wire_11915;
    wire new_Jinkela_wire_10513;
    wire new_Jinkela_wire_3156;
    wire new_Jinkela_wire_16452;
    wire new_Jinkela_wire_6807;
    wire new_Jinkela_wire_15777;
    wire new_Jinkela_wire_19858;
    wire new_Jinkela_wire_4881;
    wire new_Jinkela_wire_20179;
    wire _1071_;
    wire new_Jinkela_wire_18712;
    wire new_Jinkela_wire_12988;
    wire _1676_;
    wire new_Jinkela_wire_13939;
    wire new_Jinkela_wire_7088;
    wire new_Jinkela_wire_6004;
    wire new_Jinkela_wire_5815;
    wire new_Jinkela_wire_6813;
    wire new_Jinkela_wire_20990;
    wire new_Jinkela_wire_14722;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_11899;
    wire new_Jinkela_wire_10468;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_5361;
    wire new_Jinkela_wire_7741;
    wire new_Jinkela_wire_8902;
    wire new_Jinkela_wire_10714;
    wire new_Jinkela_wire_8565;
    wire new_Jinkela_wire_2960;
    wire new_Jinkela_wire_8717;
    wire new_Jinkela_wire_3940;
    wire new_Jinkela_wire_2180;
    wire new_Jinkela_wire_13771;
    wire new_Jinkela_wire_3735;
    wire new_Jinkela_wire_13729;
    wire new_Jinkela_wire_11859;
    wire new_Jinkela_wire_15407;
    wire new_Jinkela_wire_19357;
    wire _0000_;
    wire new_Jinkela_wire_5442;
    wire new_Jinkela_wire_6282;
    wire new_Jinkela_wire_15287;
    wire new_Jinkela_wire_16763;
    wire new_Jinkela_wire_4170;
    wire new_Jinkela_wire_18446;
    wire _1579_;
    wire new_Jinkela_wire_6215;
    wire new_Jinkela_wire_15036;
    wire _0901_;
    wire new_Jinkela_wire_1897;
    wire new_Jinkela_wire_14651;
    wire new_Jinkela_wire_18383;
    wire new_Jinkela_wire_16973;
    wire new_Jinkela_wire_11409;
    wire new_Jinkela_wire_5215;
    wire new_Jinkela_wire_1878;
    wire new_Jinkela_wire_7048;
    wire new_Jinkela_wire_10874;
    wire new_Jinkela_wire_15950;
    wire new_Jinkela_wire_4989;
    wire new_Jinkela_wire_12909;
    wire _1746_;
    wire new_Jinkela_wire_17642;
    wire new_Jinkela_wire_10050;
    wire new_Jinkela_wire_5987;
    wire new_Jinkela_wire_15046;
    wire new_Jinkela_wire_13408;
    wire new_Jinkela_wire_15137;
    wire new_Jinkela_wire_8440;
    wire new_Jinkela_wire_5636;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_21307;
    wire new_Jinkela_wire_8439;
    wire new_Jinkela_wire_921;
    wire _0815_;
    wire new_Jinkela_wire_3095;
    wire new_Jinkela_wire_12420;
    wire new_Jinkela_wire_7157;
    wire new_Jinkela_wire_14587;
    wire new_Jinkela_wire_9338;
    wire new_Jinkela_wire_2784;
    wire new_Jinkela_wire_5564;
    wire _0503_;
    wire new_Jinkela_wire_12129;
    wire new_Jinkela_wire_4290;
    wire new_Jinkela_wire_19167;
    wire new_Jinkela_wire_10237;
    wire new_Jinkela_wire_11295;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_14237;
    wire _1767_;
    wire new_Jinkela_wire_15498;
    wire new_Jinkela_wire_12283;
    wire new_Jinkela_wire_9445;
    wire new_Jinkela_wire_9979;
    wire new_Jinkela_wire_16501;
    wire new_Jinkela_wire_11607;
    wire new_Jinkela_wire_6360;
    wire new_Jinkela_wire_16610;
    wire new_Jinkela_wire_8045;
    wire new_Jinkela_wire_6990;
    wire new_Jinkela_wire_3382;
    wire new_Jinkela_wire_3922;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_14700;
    wire new_Jinkela_wire_4053;
    wire new_Jinkela_wire_3848;
    wire new_Jinkela_wire_6121;
    wire new_net_3948;
    wire new_Jinkela_wire_13092;
    wire new_Jinkela_wire_14849;
    wire new_Jinkela_wire_8106;
    wire new_Jinkela_wire_6052;
    wire new_Jinkela_wire_11187;
    wire new_Jinkela_wire_9167;
    wire new_Jinkela_wire_10998;
    wire new_Jinkela_wire_16504;
    wire new_Jinkela_wire_4386;
    wire new_Jinkela_wire_11341;
    wire new_Jinkela_wire_11715;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_4423;
    wire new_Jinkela_wire_14385;
    wire new_Jinkela_wire_1657;
    wire new_Jinkela_wire_2531;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_14442;
    wire new_Jinkela_wire_9012;
    wire new_Jinkela_wire_20608;
    wire new_Jinkela_wire_7923;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_19890;
    wire new_Jinkela_wire_18594;
    wire new_Jinkela_wire_19966;
    wire new_Jinkela_wire_15995;
    wire new_Jinkela_wire_20459;
    wire new_Jinkela_wire_3358;
    wire new_Jinkela_wire_11238;
    wire new_Jinkela_wire_7707;
    wire new_Jinkela_wire_18375;
    wire _0709_;
    wire new_Jinkela_wire_16894;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_12037;
    wire new_Jinkela_wire_5913;
    wire new_Jinkela_wire_12309;
    wire new_Jinkela_wire_15098;
    wire new_Jinkela_wire_12840;
    wire new_Jinkela_wire_6475;
    wire new_Jinkela_wire_11599;
    wire new_Jinkela_wire_14266;
    wire new_Jinkela_wire_13781;
    wire new_Jinkela_wire_10950;
    wire new_Jinkela_wire_10791;
    wire new_Jinkela_wire_17010;
    wire new_Jinkela_wire_2261;
    wire new_Jinkela_wire_5738;
    wire new_Jinkela_wire_10340;
    wire new_Jinkela_wire_21270;
    wire new_Jinkela_wire_12570;
    wire new_Jinkela_wire_11793;
    wire new_Jinkela_wire_3724;
    wire new_Jinkela_wire_16498;
    wire new_Jinkela_wire_16182;
    wire new_Jinkela_wire_4108;
    wire new_Jinkela_wire_12535;
    wire new_Jinkela_wire_15855;
    wire new_Jinkela_wire_14203;
    wire _0428_;
    wire _1231_;
    wire new_Jinkela_wire_3323;
    wire new_Jinkela_wire_15994;
    wire _0714_;
    wire new_Jinkela_wire_20782;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_17045;
    wire new_Jinkela_wire_19774;
    wire new_Jinkela_wire_5154;
    wire new_Jinkela_wire_12246;
    wire new_Jinkela_wire_6107;
    wire new_Jinkela_wire_18755;
    wire new_Jinkela_wire_11259;
    wire new_Jinkela_wire_3581;
    wire new_Jinkela_wire_1097;
    wire _1274_;
    wire new_Jinkela_wire_5496;
    wire new_Jinkela_wire_12823;
    wire new_Jinkela_wire_13205;
    wire _1445_;
    wire new_Jinkela_wire_3114;
    wire new_Jinkela_wire_18187;
    wire new_Jinkela_wire_17228;
    wire new_Jinkela_wire_14933;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_20827;
    wire _1831_;
    wire new_Jinkela_wire_6435;
    wire new_Jinkela_wire_5671;
    wire new_Jinkela_wire_9700;
    wire new_Jinkela_wire_13010;
    wire _0141_;
    wire _0799_;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_2661;
    wire new_Jinkela_wire_20572;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_5786;
    wire _1084_;
    wire new_Jinkela_wire_16106;
    wire new_Jinkela_wire_8947;
    wire new_Jinkela_wire_17800;
    wire new_Jinkela_wire_17680;
    wire new_Jinkela_wire_21255;
    wire new_Jinkela_wire_16727;
    wire new_Jinkela_wire_10208;
    wire _0521_;
    wire new_Jinkela_wire_2234;
    wire new_Jinkela_wire_5605;
    wire new_Jinkela_wire_11944;
    wire new_Jinkela_wire_12573;
    wire new_Jinkela_wire_9577;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_17807;
    wire new_Jinkela_wire_16563;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_6771;
    wire new_Jinkela_wire_18851;
    wire new_Jinkela_wire_18190;
    wire new_Jinkela_wire_14592;
    wire new_Jinkela_wire_10093;
    wire new_Jinkela_wire_16627;
    wire _1711_;
    wire new_Jinkela_wire_9515;
    wire _0814_;
    wire new_Jinkela_wire_10654;
    wire new_Jinkela_wire_5758;
    wire new_Jinkela_wire_15066;
    wire new_Jinkela_wire_7960;
    wire new_Jinkela_wire_15253;
    wire _0670_;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_20930;
    wire new_Jinkela_wire_8733;
    wire new_Jinkela_wire_2871;
    wire new_Jinkela_wire_21098;
    wire new_Jinkela_wire_11566;
    wire new_Jinkela_wire_4063;
    wire new_Jinkela_wire_5422;
    wire new_Jinkela_wire_2611;
    wire new_Jinkela_wire_5144;
    wire new_Jinkela_wire_14489;
    wire new_Jinkela_wire_963;
    wire _1414_;
    wire new_Jinkela_wire_19306;
    wire new_Jinkela_wire_18289;
    wire new_Jinkela_wire_9494;
    wire new_Jinkela_wire_12563;
    wire new_Jinkela_wire_663;
    wire new_net_3950;
    wire new_Jinkela_wire_10183;
    wire new_Jinkela_wire_16133;
    wire new_Jinkela_wire_6742;
    wire new_Jinkela_wire_8982;
    wire new_Jinkela_wire_17618;
    wire new_Jinkela_wire_21124;
    wire new_Jinkela_wire_3917;
    wire new_Jinkela_wire_17686;
    wire new_Jinkela_wire_5344;
    wire new_Jinkela_wire_5464;
    wire new_Jinkela_wire_10890;
    wire new_Jinkela_wire_6498;
    wire new_Jinkela_wire_16958;
    wire _0571_;
    wire new_Jinkela_wire_5167;
    wire new_Jinkela_wire_5873;
    wire new_Jinkela_wire_8532;
    wire _1082_;
    wire new_Jinkela_wire_11294;
    wire new_Jinkela_wire_3484;
    wire new_Jinkela_wire_17826;
    wire new_Jinkela_wire_6386;
    wire new_Jinkela_wire_11765;
    wire new_Jinkela_wire_10557;
    wire new_Jinkela_wire_20113;
    wire new_Jinkela_wire_15365;
    wire _0917_;
    wire _1285_;
    wire new_Jinkela_wire_16329;
    wire new_Jinkela_wire_11501;
    wire new_Jinkela_wire_13227;
    wire new_Jinkela_wire_12574;
    wire new_Jinkela_wire_15895;
    wire new_Jinkela_wire_20559;
    wire new_Jinkela_wire_8306;
    wire new_Jinkela_wire_19493;
    wire new_Jinkela_wire_18910;
    wire new_Jinkela_wire_8831;
    wire new_Jinkela_wire_11635;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_9666;
    wire new_Jinkela_wire_13800;
    wire new_Jinkela_wire_4779;
    wire new_Jinkela_wire_1721;
    wire new_Jinkela_wire_3374;
    wire new_Jinkela_wire_8299;
    wire new_Jinkela_wire_10944;
    wire new_Jinkela_wire_14749;
    wire new_Jinkela_wire_18258;
    wire new_Jinkela_wire_20028;
    wire new_Jinkela_wire_11302;
    wire new_Jinkela_wire_3330;
    wire new_Jinkela_wire_5041;
    wire new_Jinkela_wire_16286;
    wire new_Jinkela_wire_6756;
    wire new_Jinkela_wire_15092;
    wire new_Jinkela_wire_15108;
    wire new_Jinkela_wire_21283;
    wire new_Jinkela_wire_7129;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_8265;
    wire new_Jinkela_wire_11111;
    wire new_Jinkela_wire_5258;
    wire new_Jinkela_wire_4480;
    wire new_Jinkela_wire_19820;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_17291;
    wire new_Jinkela_wire_12932;
    wire new_Jinkela_wire_19688;
    wire new_Jinkela_wire_11887;
    wire new_Jinkela_wire_3418;
    wire new_Jinkela_wire_18316;
    wire new_Jinkela_wire_18106;
    wire new_Jinkela_wire_5264;
    wire new_Jinkela_wire_19147;
    wire new_Jinkela_wire_13217;
    wire new_Jinkela_wire_6441;
    wire new_Jinkela_wire_8705;
    wire new_Jinkela_wire_11383;
    wire new_Jinkela_wire_9984;
    wire new_Jinkela_wire_10000;
    wire new_Jinkela_wire_17568;
    wire _0576_;
    wire new_Jinkela_wire_12156;
    wire new_Jinkela_wire_6997;
    wire new_Jinkela_wire_18209;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_21029;
    wire new_Jinkela_wire_5770;
    wire new_Jinkela_wire_16451;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_15894;
    wire new_Jinkela_wire_14532;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_5801;
    wire _0647_;
    wire new_Jinkela_wire_19470;
    wire new_Jinkela_wire_4199;
    wire new_Jinkela_wire_19336;
    wire new_Jinkela_wire_7819;
    wire new_Jinkela_wire_8475;
    wire new_Jinkela_wire_4996;
    wire _1324_;
    wire new_Jinkela_wire_20847;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_7967;
    wire new_Jinkela_wire_11972;
    wire new_Jinkela_wire_17488;
    wire new_Jinkela_wire_20346;
    wire new_Jinkela_wire_5141;
    wire new_Jinkela_wire_17643;
    wire new_Jinkela_wire_9594;
    wire new_Jinkela_wire_18073;
    wire new_Jinkela_wire_6045;
    wire new_Jinkela_wire_19996;
    wire new_Jinkela_wire_10218;
    wire new_Jinkela_wire_10200;
    wire new_Jinkela_wire_9273;
    wire new_Jinkela_wire_8256;
    wire new_Jinkela_wire_15370;
    wire new_Jinkela_wire_835;
    wire new_Jinkela_wire_8327;
    wire new_Jinkela_wire_8482;
    wire new_Jinkela_wire_11329;
    wire new_Jinkela_wire_13358;
    wire new_Jinkela_wire_7791;
    wire new_Jinkela_wire_7705;
    wire new_Jinkela_wire_11155;
    wire new_Jinkela_wire_17376;
    wire new_Jinkela_wire_17182;
    wire new_Jinkela_wire_5903;
    wire new_Jinkela_wire_16417;
    wire new_Jinkela_wire_8790;
    wire new_Jinkela_wire_13262;
    wire new_Jinkela_wire_9440;
    wire new_Jinkela_wire_18764;
    wire new_Jinkela_wire_13124;
    wire new_Jinkela_wire_18918;
    wire new_Jinkela_wire_16391;
    wire new_Jinkela_wire_12082;
    wire new_Jinkela_wire_13309;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_13678;
    wire new_Jinkela_wire_2744;
    wire new_Jinkela_wire_14353;
    wire _0128_;
    wire new_Jinkela_wire_16966;
    wire new_Jinkela_wire_10645;
    wire new_Jinkela_wire_4361;
    wire new_Jinkela_wire_12445;
    wire new_Jinkela_wire_18857;
    wire new_Jinkela_wire_14727;
    wire new_net_3936;
    wire new_Jinkela_wire_16439;
    wire new_Jinkela_wire_15745;
    wire new_Jinkela_wire_12886;
    wire new_Jinkela_wire_8354;
    wire new_Jinkela_wire_14049;
    wire new_Jinkela_wire_3272;
    wire new_Jinkela_wire_6005;
    wire new_Jinkela_wire_9737;
    wire new_Jinkela_wire_16976;
    wire new_Jinkela_wire_5449;
    wire new_Jinkela_wire_10272;
    wire new_Jinkela_wire_6943;
    wire _0878_;
    wire new_Jinkela_wire_5772;
    wire new_Jinkela_wire_11965;
    wire new_Jinkela_wire_7734;
    wire new_Jinkela_wire_13181;
    wire new_Jinkela_wire_2626;
    wire new_Jinkela_wire_2297;
    wire new_Jinkela_wire_516;
    wire new_Jinkela_wire_15343;
    wire new_Jinkela_wire_4732;
    wire new_Jinkela_wire_14409;
    wire new_Jinkela_wire_18728;
    wire new_Jinkela_wire_17735;
    wire new_Jinkela_wire_9474;
    wire new_Jinkela_wire_5900;
    wire new_Jinkela_wire_1904;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_6220;
    wire new_Jinkela_wire_3267;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_8503;
    wire new_Jinkela_wire_13020;
    wire new_Jinkela_wire_21007;
    wire new_Jinkela_wire_12182;
    wire new_Jinkela_wire_17923;
    wire new_Jinkela_wire_21034;
    wire new_Jinkela_wire_13871;
    wire new_Jinkela_wire_8015;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_17251;
    wire new_Jinkela_wire_4359;
    wire new_Jinkela_wire_11979;
    wire new_Jinkela_wire_15072;
    wire new_Jinkela_wire_2530;
    wire new_Jinkela_wire_8442;
    wire new_Jinkela_wire_13264;
    wire new_Jinkela_wire_17678;
    wire new_Jinkela_wire_3393;
    wire new_Jinkela_wire_14360;
    wire new_Jinkela_wire_9565;
    wire new_Jinkela_wire_2843;
    wire new_Jinkela_wire_18425;
    wire new_Jinkela_wire_13195;
    wire new_Jinkela_wire_11818;
    wire new_Jinkela_wire_4322;
    wire new_Jinkela_wire_20060;
    wire new_Jinkela_wire_8037;
    wire new_Jinkela_wire_17773;
    wire new_Jinkela_wire_2214;
    wire new_Jinkela_wire_8991;
    wire new_Jinkela_wire_15778;
    wire _0195_;
    wire new_Jinkela_wire_11137;
    wire new_Jinkela_wire_7716;
    wire new_Jinkela_wire_19238;
    wire new_Jinkela_wire_2170;
    wire new_Jinkela_wire_16177;
    wire new_Jinkela_wire_18419;
    wire new_Jinkela_wire_8044;
    wire new_Jinkela_wire_11931;
    wire new_Jinkela_wire_12227;
    wire new_Jinkela_wire_10856;
    wire new_Jinkela_wire_13269;
    wire new_Jinkela_wire_18447;
    wire new_Jinkela_wire_6055;
    wire new_Jinkela_wire_13444;
    wire new_Jinkela_wire_19385;
    wire new_Jinkela_wire_7679;
    wire new_Jinkela_wire_14161;
    wire new_Jinkela_wire_9580;
    wire new_Jinkela_wire_20058;
    wire new_Jinkela_wire_16948;
    wire new_Jinkela_wire_17921;
    wire new_Jinkela_wire_5660;
    wire new_Jinkela_wire_11985;
    wire new_Jinkela_wire_16765;
    wire _0624_;
    wire new_Jinkela_wire_7822;
    wire new_Jinkela_wire_10129;
    wire new_Jinkela_wire_21280;
    wire new_Jinkela_wire_16441;
    wire new_Jinkela_wire_6135;
    wire new_Jinkela_wire_15690;
    wire _1702_;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_15418;
    wire new_Jinkela_wire_16318;
    wire _0278_;
    wire new_Jinkela_wire_18029;
    wire new_Jinkela_wire_5752;
    wire new_Jinkela_wire_18329;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_3454;
    wire _0623_;
    wire new_Jinkela_wire_18810;
    wire new_Jinkela_wire_20845;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_4193;
    wire new_Jinkela_wire_4658;
    wire _1397_;
    wire new_Jinkela_wire_6544;
    wire new_Jinkela_wire_17630;
    wire new_Jinkela_wire_5189;
    wire new_Jinkela_wire_18576;
    wire new_Jinkela_wire_12295;
    wire new_Jinkela_wire_6025;
    wire new_Jinkela_wire_3540;
    wire new_Jinkela_wire_19176;
    wire new_Jinkela_wire_10572;
    wire new_Jinkela_wire_2522;
    wire new_Jinkela_wire_8860;
    wire new_Jinkela_wire_4968;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_6299;
    wire new_Jinkela_wire_3920;
    wire new_Jinkela_wire_7568;
    wire _1201_;
    wire new_Jinkela_wire_12496;
    wire new_Jinkela_wire_19004;
    wire new_Jinkela_wire_15582;
    wire new_Jinkela_wire_7096;
    wire new_Jinkela_wire_3494;
    wire new_Jinkela_wire_18205;
    wire new_Jinkela_wire_13978;
    wire new_Jinkela_wire_18995;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_4188;
    wire new_Jinkela_wire_5136;
    wire new_Jinkela_wire_13472;
    wire new_Jinkela_wire_3347;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_17526;
    wire new_Jinkela_wire_12973;
    wire new_Jinkela_wire_19055;
    wire new_Jinkela_wire_4647;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_8693;
    wire _1318_;
    wire new_Jinkela_wire_10753;
    wire new_Jinkela_wire_12278;
    wire new_Jinkela_wire_18318;
    wire new_Jinkela_wire_3296;
    wire new_Jinkela_wire_7551;
    wire new_Jinkela_wire_10421;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_19269;
    wire new_Jinkela_wire_3185;
    wire new_Jinkela_wire_2872;
    wire new_Jinkela_wire_18138;
    wire new_Jinkela_wire_14215;
    wire new_Jinkela_wire_5884;
    wire new_Jinkela_wire_8043;
    wire new_Jinkela_wire_10443;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_3251;
    wire new_Jinkela_wire_14223;
    wire new_Jinkela_wire_4054;
    wire new_Jinkela_wire_10500;
    wire new_Jinkela_wire_11320;
    wire new_Jinkela_wire_10358;
    wire new_Jinkela_wire_17396;
    wire new_Jinkela_wire_10803;
    wire new_Jinkela_wire_17303;
    wire new_Jinkela_wire_8720;
    wire _1508_;
    wire _0056_;
    wire new_Jinkela_wire_15483;
    wire new_Jinkela_wire_21048;
    wire new_Jinkela_wire_2903;
    wire new_Jinkela_wire_4369;
    wire new_Jinkela_wire_4081;
    wire new_Jinkela_wire_6404;
    wire new_Jinkela_wire_4897;
    wire new_Jinkela_wire_14842;
    wire new_Jinkela_wire_15617;
    wire new_Jinkela_wire_20667;
    wire new_Jinkela_wire_19477;
    wire new_Jinkela_wire_19849;
    wire new_Jinkela_wire_10492;
    wire new_Jinkela_wire_10758;
    wire new_Jinkela_wire_14233;
    wire new_Jinkela_wire_2122;
    wire new_Jinkela_wire_19750;
    wire new_Jinkela_wire_7057;
    wire new_Jinkela_wire_5622;
    wire new_Jinkela_wire_2369;
    wire new_Jinkela_wire_7209;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_8491;
    wire new_Jinkela_wire_15551;
    wire new_Jinkela_wire_8410;
    wire new_Jinkela_wire_9806;
    wire new_Jinkela_wire_13060;
    wire new_Jinkela_wire_7845;
    wire _1752_;
    wire new_Jinkela_wire_1747;
    wire new_Jinkela_wire_2655;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_20309;
    wire new_Jinkela_wire_2767;
    wire new_Jinkela_wire_19467;
    wire new_Jinkela_wire_16469;
    wire new_Jinkela_wire_8197;
    wire new_Jinkela_wire_7607;
    wire new_Jinkela_wire_15751;
    wire new_Jinkela_wire_6034;
    wire new_Jinkela_wire_19951;
    wire new_Jinkela_wire_8848;
    wire new_Jinkela_wire_16984;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_10586;
    wire new_Jinkela_wire_14033;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_6909;
    wire _0981_;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_9541;
    wire new_Jinkela_wire_9179;
    wire new_Jinkela_wire_5428;
    wire new_Jinkela_wire_19950;
    wire new_Jinkela_wire_18699;
    wire new_Jinkela_wire_16232;
    wire new_Jinkela_wire_7476;
    wire new_Jinkela_wire_15591;
    wire new_Jinkela_wire_17277;
    wire new_Jinkela_wire_2667;
    wire new_Jinkela_wire_13505;
    wire new_Jinkela_wire_10217;
    wire new_Jinkela_wire_12564;
    wire _0363_;
    wire new_Jinkela_wire_17681;
    wire new_Jinkela_wire_4892;
    wire new_Jinkela_wire_10887;
    wire new_Jinkela_wire_8026;
    wire new_Jinkela_wire_6755;
    wire new_Jinkela_wire_20796;
    wire new_Jinkela_wire_1916;
    wire new_Jinkela_wire_13596;
    wire new_Jinkela_wire_17567;
    wire new_Jinkela_wire_4518;
    wire new_Jinkela_wire_18287;
    wire new_Jinkela_wire_11513;
    wire _0274_;
    wire new_Jinkela_wire_4911;
    wire new_Jinkela_wire_14580;
    wire new_Jinkela_wire_4742;
    wire new_Jinkela_wire_20271;
    wire new_Jinkela_wire_5106;
    wire new_Jinkela_wire_21203;
    wire new_Jinkela_wire_17411;
    wire new_Jinkela_wire_100;
    wire _0414_;
    wire new_Jinkela_wire_17874;
    wire new_Jinkela_wire_11360;
    wire new_Jinkela_wire_17463;
    wire new_Jinkela_wire_15419;
    wire new_Jinkela_wire_6974;
    wire new_Jinkela_wire_12324;
    wire new_Jinkela_wire_15692;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_17121;
    wire new_Jinkela_wire_7487;
    wire new_Jinkela_wire_7918;
    wire new_Jinkela_wire_18780;
    wire new_Jinkela_wire_20882;
    wire new_Jinkela_wire_6512;
    wire new_Jinkela_wire_4864;
    wire new_Jinkela_wire_12261;
    wire new_Jinkela_wire_18557;
    wire new_Jinkela_wire_8316;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_12395;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_5431;
    wire new_Jinkela_wire_11452;
    wire new_Jinkela_wire_13790;
    wire new_Jinkela_wire_19481;
    wire new_Jinkela_wire_7242;
    wire _0518_;
    wire new_Jinkela_wire_10722;
    wire new_Jinkela_wire_16947;
    wire _1624_;
    wire _0586_;
    wire _0314_;
    wire new_Jinkela_wire_19218;
    wire new_Jinkela_wire_13708;
    wire new_Jinkela_wire_19903;
    wire new_Jinkela_wire_21202;
    wire new_Jinkela_wire_8779;
    wire new_Jinkela_wire_17648;
    wire new_Jinkela_wire_7630;
    wire new_Jinkela_wire_10929;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_4179;
    wire new_Jinkela_wire_7735;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_6548;
    wire new_Jinkela_wire_9144;
    wire new_Jinkela_wire_12041;
    wire new_Jinkela_wire_4934;
    wire new_Jinkela_wire_6525;
    wire new_Jinkela_wire_9502;
    wire new_Jinkela_wire_9457;
    wire new_Jinkela_wire_20590;
    wire new_Jinkela_wire_19410;
    wire new_Jinkela_wire_8523;
    wire new_Jinkela_wire_3159;
    wire new_Jinkela_wire_16990;
    wire new_Jinkela_wire_8856;
    wire new_Jinkela_wire_19225;
    wire _1619_;
    wire new_Jinkela_wire_11069;
    wire new_Jinkela_wire_4485;
    wire new_Jinkela_wire_15953;
    wire new_Jinkela_wire_7586;
    wire new_Jinkela_wire_19188;
    wire new_Jinkela_wire_9644;
    wire new_Jinkela_wire_19644;
    wire _1532_;
    wire new_Jinkela_wire_13416;
    wire new_Jinkela_wire_19548;
    wire new_Jinkela_wire_15318;
    wire new_Jinkela_wire_5856;
    wire new_Jinkela_wire_14251;
    wire new_Jinkela_wire_13298;
    wire _1356_;
    wire new_Jinkela_wire_7682;
    wire new_Jinkela_wire_14963;
    wire new_Jinkela_wire_6476;
    wire new_Jinkela_wire_18241;
    wire new_Jinkela_wire_9040;
    wire new_Jinkela_wire_2375;
    wire new_Jinkela_wire_18513;
    wire new_Jinkela_wire_4649;
    wire new_Jinkela_wire_15637;
    wire new_Jinkela_wire_4296;
    wire new_Jinkela_wire_6518;
    wire new_Jinkela_wire_20290;
    wire new_Jinkela_wire_6083;
    wire new_Jinkela_wire_13079;
    wire _0272_;
    wire new_Jinkela_wire_16020;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_5698;
    wire new_Jinkela_wire_10952;
    wire new_Jinkela_wire_9981;
    wire new_Jinkela_wire_6885;
    wire new_Jinkela_wire_11812;
    wire new_Jinkela_wire_3794;
    wire new_Jinkela_wire_7133;
    wire _0025_;
    wire new_Jinkela_wire_1819;
    wire new_Jinkela_wire_7837;
    wire new_Jinkela_wire_9174;
    wire new_Jinkela_wire_4656;
    wire new_Jinkela_wire_6196;
    wire new_Jinkela_wire_19924;
    wire new_Jinkela_wire_6092;
    wire new_Jinkela_wire_12871;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_1549;
    wire new_Jinkela_wire_16085;
    wire new_Jinkela_wire_6740;
    wire new_Jinkela_wire_2247;
    wire new_Jinkela_wire_12094;
    wire new_Jinkela_wire_8144;
    wire new_Jinkela_wire_16838;
    wire new_Jinkela_wire_17633;
    wire new_Jinkela_wire_3792;
    wire new_Jinkela_wire_1357;
    wire _0865_;
    wire new_Jinkela_wire_5051;
    wire new_Jinkela_wire_13514;
    wire new_Jinkela_wire_18908;
    wire _0543_;
    wire new_Jinkela_wire_11479;
    wire _0485_;
    wire new_Jinkela_wire_4830;
    wire new_Jinkela_wire_17168;
    wire new_Jinkela_wire_18775;
    wire new_Jinkela_wire_13675;
    wire new_Jinkela_wire_18048;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_9738;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_8614;
    wire new_Jinkela_wire_20842;
    wire new_Jinkela_wire_4745;
    wire new_Jinkela_wire_12077;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_14071;
    wire new_Jinkela_wire_11992;
    wire new_Jinkela_wire_20511;
    wire new_Jinkela_wire_2279;
    wire new_Jinkela_wire_10483;
    wire new_Jinkela_wire_16489;
    wire new_Jinkela_wire_12737;
    wire new_Jinkela_wire_20819;
    wire new_Jinkela_wire_10222;
    wire new_Jinkela_wire_16952;
    wire new_Jinkela_wire_15593;
    wire new_Jinkela_wire_17292;
    wire new_Jinkela_wire_6877;
    wire _1643_;
    wire new_Jinkela_wire_16593;
    wire new_Jinkela_wire_19901;
    wire new_Jinkela_wire_16753;
    wire new_Jinkela_wire_10485;
    wire new_Jinkela_wire_3140;
    wire new_Jinkela_wire_18948;
    wire new_Jinkela_wire_6942;
    wire _0873_;
    wire new_Jinkela_wire_9988;
    wire _1609_;
    wire new_Jinkela_wire_8954;
    wire new_Jinkela_wire_7695;
    wire new_Jinkela_wire_15171;
    wire new_Jinkela_wire_16863;
    wire new_Jinkela_wire_11269;
    wire new_Jinkela_wire_17355;
    wire new_Jinkela_wire_18044;
    wire new_Jinkela_wire_18017;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_18767;
    wire new_Jinkela_wire_8855;
    wire new_Jinkela_wire_2993;
    wire new_Jinkela_wire_11325;
    wire new_Jinkela_wire_17015;
    wire new_Jinkela_wire_12282;
    wire new_Jinkela_wire_11333;
    wire new_Jinkela_wire_1717;
    wire _0902_;
    wire new_Jinkela_wire_20649;
    wire _1081_;
    wire new_Jinkela_wire_18973;
    wire new_Jinkela_wire_8393;
    wire new_Jinkela_wire_17944;
    wire new_Jinkela_wire_2806;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_17764;
    wire new_Jinkela_wire_20864;
    wire new_Jinkela_wire_19553;
    wire new_Jinkela_wire_8005;
    wire new_Jinkela_wire_10859;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_14668;
    wire _0083_;
    wire new_Jinkela_wire_8332;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_2814;
    wire new_Jinkela_wire_12718;
    wire new_Jinkela_wire_7895;
    wire new_Jinkela_wire_18792;
    wire new_Jinkela_wire_13766;
    wire new_Jinkela_wire_7207;
    wire new_Jinkela_wire_20531;
    wire new_Jinkela_wire_6716;
    wire new_Jinkela_wire_8683;
    wire new_Jinkela_wire_2311;
    wire new_Jinkela_wire_6562;
    wire new_Jinkela_wire_16497;
    wire new_Jinkela_wire_4684;
    wire new_Jinkela_wire_3398;
    wire new_Jinkela_wire_11081;
    wire new_Jinkela_wire_6930;
    wire new_Jinkela_wire_17206;
    wire new_Jinkela_wire_7842;
    wire new_Jinkela_wire_10120;
    wire new_Jinkela_wire_2826;
    wire _0159_;
    wire _1305_;
    wire new_Jinkela_wire_11139;
    wire new_Jinkela_wire_21192;
    wire new_Jinkela_wire_4325;
    wire new_Jinkela_wire_13334;
    wire new_Jinkela_wire_3525;
    wire new_Jinkela_wire_6950;
    wire new_Jinkela_wire_14978;
    wire _0331_;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_16434;
    wire new_Jinkela_wire_3075;
    wire new_Jinkela_wire_3145;
    wire new_Jinkela_wire_7055;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_3080;
    wire _0215_;
    wire new_Jinkela_wire_4833;
    wire new_Jinkela_wire_13906;
    wire new_Jinkela_wire_5287;
    wire new_Jinkela_wire_17279;
    wire new_Jinkela_wire_14657;
    wire new_Jinkela_wire_3769;
    wire new_Jinkela_wire_3462;
    wire _0871_;
    wire new_Jinkela_wire_4056;
    wire new_Jinkela_wire_18975;
    wire new_Jinkela_wire_5158;
    wire new_Jinkela_wire_7090;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_9044;
    wire _1159_;
    wire new_Jinkela_wire_12415;
    wire new_Jinkela_wire_14540;
    wire new_Jinkela_wire_7599;
    wire new_Jinkela_wire_9796;
    wire new_Jinkela_wire_10772;
    wire new_Jinkela_wire_304;
    wire _1382_;
    wire new_Jinkela_wire_16902;
    wire new_Jinkela_wire_14217;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_21248;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_5684;
    wire new_Jinkela_wire_10549;
    wire new_Jinkela_wire_7534;
    wire new_Jinkela_wire_8129;
    wire _1741_;
    wire new_Jinkela_wire_12994;
    wire _1734_;
    wire _1120_;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_11771;
    wire new_Jinkela_wire_17991;
    wire new_Jinkela_wire_3722;
    wire new_Jinkela_wire_17895;
    wire new_Jinkela_wire_12852;
    wire new_Jinkela_wire_4153;
    wire _0075_;
    wire new_Jinkela_wire_6353;
    wire new_Jinkela_wire_20379;
    wire new_Jinkela_wire_12772;
    wire new_Jinkela_wire_10068;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_12561;
    wire new_Jinkela_wire_14158;
    wire new_Jinkela_wire_7743;
    wire new_Jinkela_wire_6053;
    wire new_Jinkela_wire_13971;
    wire new_Jinkela_wire_18045;
    wire new_Jinkela_wire_15327;
    wire new_Jinkela_wire_5933;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_17765;
    wire new_Jinkela_wire_12776;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_11024;
    wire new_Jinkela_wire_14534;
    wire new_Jinkela_wire_21241;
    wire new_Jinkela_wire_17707;
    wire new_Jinkela_wire_10665;
    wire new_Jinkela_wire_15341;
    wire new_Jinkela_wire_1855;
    wire _0100_;
    wire new_Jinkela_wire_4420;
    wire new_Jinkela_wire_4651;
    wire new_Jinkela_wire_2056;
    wire new_Jinkela_wire_18286;
    wire new_Jinkela_wire_2419;
    wire new_Jinkela_wire_11119;
    wire new_Jinkela_wire_18542;
    wire new_Jinkela_wire_4999;
    wire new_Jinkela_wire_2607;
    wire new_Jinkela_wire_5067;
    wire new_Jinkela_wire_7766;
    wire new_Jinkela_wire_15906;
    wire new_Jinkela_wire_17929;
    wire new_Jinkela_wire_8381;
    wire new_Jinkela_wire_16711;
    wire new_Jinkela_wire_7163;
    wire new_Jinkela_wire_3269;
    wire new_Jinkela_wire_11588;
    wire new_Jinkela_wire_15379;
    wire new_Jinkela_wire_13428;
    wire new_Jinkela_wire_19784;
    wire new_Jinkela_wire_3384;
    wire _0907_;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_7718;
    wire new_Jinkela_wire_11967;
    wire new_Jinkela_wire_19669;
    wire new_Jinkela_wire_15042;
    wire new_Jinkela_wire_19504;
    wire new_Jinkela_wire_7633;
    wire new_Jinkela_wire_19975;
    wire new_Jinkela_wire_12374;
    wire new_Jinkela_wire_5908;
    wire new_Jinkela_wire_11311;
    wire new_Jinkela_wire_9235;
    wire new_Jinkela_wire_3902;
    wire _0638_;
    wire new_Jinkela_wire_11534;
    wire new_Jinkela_wire_1709;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_17331;
    wire new_Jinkela_wire_9957;
    wire new_Jinkela_wire_17775;
    wire new_Jinkela_wire_2030;
    wire new_Jinkela_wire_19663;
    wire new_Jinkela_wire_18806;
    wire new_Jinkela_wire_5630;
    wire new_Jinkela_wire_8169;
    wire new_Jinkela_wire_12161;
    wire new_Jinkela_wire_12249;
    wire new_Jinkela_wire_13006;
    wire new_Jinkela_wire_10672;
    wire _1460_;
    wire new_Jinkela_wire_13077;
    wire new_Jinkela_wire_13799;
    wire new_Jinkela_wire_20941;
    wire new_Jinkela_wire_3618;
    wire new_Jinkela_wire_11350;
    wire new_Jinkela_wire_17264;
    wire new_Jinkela_wire_18670;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_12238;
    wire new_Jinkela_wire_9485;
    wire new_Jinkela_wire_20547;
    wire new_Jinkela_wire_14771;
    wire new_Jinkela_wire_10980;
    wire new_Jinkela_wire_17021;
    wire new_Jinkela_wire_2107;
    wire new_Jinkela_wire_10185;
    wire new_Jinkela_wire_8547;
    wire new_Jinkela_wire_8529;
    wire new_Jinkela_wire_7521;
    wire new_Jinkela_wire_5658;
    wire new_Jinkela_wire_20961;
    wire new_Jinkela_wire_13995;
    wire new_Jinkela_wire_12579;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_7658;
    wire _1744_;
    wire new_Jinkela_wire_20148;
    wire new_Jinkela_wire_21082;
    wire new_Jinkela_wire_279;
    wire new_Jinkela_wire_19085;
    wire new_Jinkela_wire_10455;
    wire new_Jinkela_wire_1746;
    wire new_Jinkela_wire_3284;
    wire new_Jinkela_wire_4807;
    wire new_Jinkela_wire_17935;
    wire new_Jinkela_wire_61;
    wire _1599_;
    wire new_Jinkela_wire_16277;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_15739;
    wire new_Jinkela_wire_10302;
    wire new_Jinkela_wire_6204;
    wire new_Jinkela_wire_9928;
    wire new_Jinkela_wire_8536;
    wire new_Jinkela_wire_11304;
    wire new_Jinkela_wire_12029;
    wire _0532_;
    wire new_Jinkela_wire_5401;
    wire new_Jinkela_wire_5943;
    wire new_Jinkela_wire_9451;
    wire new_Jinkela_wire_4172;
    wire new_Jinkela_wire_19327;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_16250;
    wire new_Jinkela_wire_18231;
    wire new_Jinkela_wire_14165;
    wire new_Jinkela_wire_14966;
    wire new_Jinkela_wire_10233;
    wire new_Jinkela_wire_14466;
    wire new_Jinkela_wire_16485;
    wire new_Jinkela_wire_18844;
    wire _0041_;
    wire new_Jinkela_wire_5699;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_16144;
    wire new_Jinkela_wire_238;
    wire _0492_;
    wire new_Jinkela_wire_11761;
    wire new_Jinkela_wire_19502;
    wire new_Jinkela_wire_12083;
    wire new_Jinkela_wire_3168;
    wire new_Jinkela_wire_12837;
    wire new_Jinkela_wire_18577;
    wire new_Jinkela_wire_15247;
    wire new_Jinkela_wire_4868;
    wire new_Jinkela_wire_19206;
    wire new_Jinkela_wire_12531;
    wire new_Jinkela_wire_10616;
    wire new_Jinkela_wire_21151;
    wire new_Jinkela_wire_3417;
    wire new_Jinkela_wire_9682;
    wire new_Jinkela_wire_8054;
    wire new_Jinkela_wire_13685;
    wire new_Jinkela_wire_3465;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_10788;
    wire new_Jinkela_wire_14333;
    wire new_Jinkela_wire_6854;
    wire new_Jinkela_wire_11453;
    wire _1756_;
    wire new_Jinkela_wire_5347;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_13186;
    wire new_Jinkela_wire_17688;
    wire new_Jinkela_wire_11194;
    wire new_Jinkela_wire_11474;
    wire new_Jinkela_wire_2902;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_14929;
    wire new_Jinkela_wire_16260;
    wire new_Jinkela_wire_3449;
    wire new_Jinkela_wire_7729;
    wire new_Jinkela_wire_9407;
    wire new_Jinkela_wire_14281;
    wire new_Jinkela_wire_14641;
    wire new_Jinkela_wire_16472;
    wire new_Jinkela_wire_2009;
    wire new_Jinkela_wire_8628;
    wire new_Jinkela_wire_4136;
    wire new_Jinkela_wire_3526;
    wire new_Jinkela_wire_2316;
    wire new_Jinkela_wire_5295;
    wire new_Jinkela_wire_20381;
    wire new_Jinkela_wire_11783;
    wire new_Jinkela_wire_8271;
    wire new_Jinkela_wire_1202;
    wire new_Jinkela_wire_5029;
    wire new_Jinkela_wire_8460;
    wire new_Jinkela_wire_5450;
    wire new_Jinkela_wire_6003;
    wire new_Jinkela_wire_9333;
    wire new_Jinkela_wire_7443;
    wire new_Jinkela_wire_17823;
    wire new_Jinkela_wire_10191;
    wire new_Jinkela_wire_16359;
    wire new_Jinkela_wire_10553;
    wire new_Jinkela_wire_8388;
    wire new_Jinkela_wire_10201;
    wire _0778_;
    wire new_Jinkela_wire_17023;
    wire new_Jinkela_wire_3172;
    wire new_Jinkela_wire_11443;
    wire new_Jinkela_wire_10055;
    wire new_Jinkela_wire_18219;
    wire new_Jinkela_wire_3225;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_8709;
    wire new_Jinkela_wire_2629;
    wire new_Jinkela_wire_19521;
    wire new_Jinkela_wire_5934;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_15900;
    wire new_Jinkela_wire_15720;
    wire new_Jinkela_wire_8224;
    wire _0562_;
    wire _1603_;
    wire new_Jinkela_wire_13152;
    wire new_Jinkela_wire_18131;
    wire _1179_;
    wire new_Jinkela_wire_4129;
    wire new_Jinkela_wire_2025;
    wire _0470_;
    wire new_Jinkela_wire_7358;
    wire new_Jinkela_wire_13032;
    wire new_Jinkela_wire_6313;
    wire new_Jinkela_wire_10310;
    wire new_Jinkela_wire_16001;
    wire new_Jinkela_wire_19017;
    wire new_Jinkela_wire_13524;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_2395;
    wire new_Jinkela_wire_2859;
    wire new_Jinkela_wire_20262;
    wire new_Jinkela_wire_10195;
    wire new_Jinkela_wire_13310;
    wire _0002_;
    wire new_Jinkela_wire_18661;
    wire new_Jinkela_wire_7546;
    wire new_Jinkela_wire_3562;
    wire _1673_;
    wire new_Jinkela_wire_1763;
    wire new_Jinkela_wire_19382;
    wire new_Jinkela_wire_14775;
    wire new_Jinkela_wire_20378;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_16362;
    wire new_Jinkela_wire_19235;
    wire new_Jinkela_wire_9406;
    wire new_Jinkela_wire_16575;
    wire new_Jinkela_wire_20984;
    wire new_Jinkela_wire_20193;
    wire _0789_;
    wire new_Jinkela_wire_5978;
    wire new_Jinkela_wire_17789;
    wire new_Jinkela_wire_19394;
    wire new_Jinkela_wire_7039;
    wire new_Jinkela_wire_2973;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_11271;
    wire new_Jinkela_wire_6402;
    wire new_Jinkela_wire_15890;
    wire new_Jinkela_wire_9589;
    wire new_Jinkela_wire_17841;
    wire new_Jinkela_wire_18813;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_9073;
    wire new_Jinkela_wire_13666;
    wire new_Jinkela_wire_9295;
    wire new_Jinkela_wire_18278;
    wire new_Jinkela_wire_11856;
    wire new_Jinkela_wire_10459;
    wire new_Jinkela_wire_2657;
    wire new_Jinkela_wire_4912;
    wire new_Jinkela_wire_11420;
    wire new_Jinkela_wire_10377;
    wire new_Jinkela_wire_11710;
    wire new_Jinkela_wire_3854;
    wire new_Jinkela_wire_7571;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_6532;
    wire new_Jinkela_wire_12401;
    wire new_Jinkela_wire_19140;
    wire new_Jinkela_wire_12883;
    wire new_Jinkela_wire_16192;
    wire new_Jinkela_wire_20298;
    wire new_Jinkela_wire_7002;
    wire new_Jinkela_wire_8375;
    wire new_Jinkela_wire_6698;
    wire new_Jinkela_wire_7492;
    wire new_Jinkela_wire_4233;
    wire new_Jinkela_wire_13253;
    wire _0500_;
    wire new_Jinkela_wire_8147;
    wire new_Jinkela_wire_3796;
    wire new_Jinkela_wire_19875;
    wire new_Jinkela_wire_15214;
    wire new_Jinkela_wire_10596;
    wire new_Jinkela_wire_5311;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_13985;
    wire _1017_;
    wire new_Jinkela_wire_6266;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_3929;
    wire new_Jinkela_wire_8782;
    wire new_Jinkela_wire_4648;
    wire new_Jinkela_wire_16688;
    wire new_Jinkela_wire_6364;
    wire new_Jinkela_wire_9537;
    wire new_Jinkela_wire_18155;
    wire new_Jinkela_wire_17079;
    wire new_Jinkela_wire_19465;
    wire new_Jinkela_wire_17938;
    wire new_Jinkela_wire_19559;
    wire new_Jinkela_wire_5151;
    wire new_Jinkela_wire_16047;
    wire new_Jinkela_wire_10627;
    wire new_Jinkela_wire_11487;
    wire new_Jinkela_wire_16162;
    wire new_Jinkela_wire_17825;
    wire new_Jinkela_wire_20721;
    wire new_Jinkela_wire_981;
    wire new_Jinkela_wire_14630;
    wire _1621_;
    wire new_Jinkela_wire_1818;
    wire _0753_;
    wire new_Jinkela_wire_13949;
    wire new_Jinkela_wire_15239;
    wire new_Jinkela_wire_16648;
    wire _0858_;
    wire new_Jinkela_wire_9363;
    wire new_Jinkela_wire_15075;
    wire new_Jinkela_wire_19226;
    wire new_Jinkela_wire_18528;
    wire new_Jinkela_wire_18214;
    wire new_Jinkela_wire_16520;
    wire new_Jinkela_wire_7401;
    wire _0161_;
    wire new_Jinkela_wire_5296;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_13924;
    wire new_Jinkela_wire_11309;
    wire new_Jinkela_wire_8563;
    wire new_Jinkela_wire_12664;
    wire new_Jinkela_wire_15971;
    wire new_Jinkela_wire_9206;
    wire new_Jinkela_wire_14118;
    wire new_Jinkela_wire_14219;
    wire new_Jinkela_wire_16848;
    wire new_Jinkela_wire_11027;
    wire new_Jinkela_wire_11609;
    wire new_Jinkela_wire_6842;
    wire new_Jinkela_wire_3742;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_10033;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_15232;
    wire new_Jinkela_wire_5570;
    wire new_Jinkela_wire_15632;
    wire new_Jinkela_wire_18691;
    wire new_Jinkela_wire_18386;
    wire new_Jinkela_wire_20899;
    wire new_Jinkela_wire_6801;
    wire new_Jinkela_wire_17555;
    wire _0202_;
    wire new_Jinkela_wire_7762;
    wire new_Jinkela_wire_3211;
    wire new_Jinkela_wire_15523;
    wire new_Jinkela_wire_2614;
    wire new_Jinkela_wire_7234;
    wire _0874_;
    wire new_Jinkela_wire_4769;
    wire new_Jinkela_wire_9914;
    wire new_Jinkela_wire_18226;
    wire new_Jinkela_wire_10507;
    wire new_Jinkela_wire_17084;
    wire new_Jinkela_wire_8235;
    wire new_Jinkela_wire_13277;
    wire new_Jinkela_wire_13660;
    wire new_Jinkela_wire_16574;
    wire new_Jinkela_wire_20868;
    wire new_Jinkela_wire_18696;
    wire new_Jinkela_wire_6553;
    wire new_Jinkela_wire_13794;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_18659;
    wire new_Jinkela_wire_8200;
    wire new_Jinkela_wire_15378;
    wire new_Jinkela_wire_7562;
    wire new_Jinkela_wire_17673;
    wire new_Jinkela_wire_19456;
    wire new_Jinkela_wire_14830;
    wire new_Jinkela_wire_4606;
    wire new_Jinkela_wire_18281;
    wire new_Jinkela_wire_9529;
    wire new_Jinkela_wire_3232;
    wire new_Jinkela_wire_11719;
    wire _1672_;
    wire new_Jinkela_wire_10159;
    wire new_Jinkela_wire_2179;
    wire new_Jinkela_wire_4184;
    wire new_Jinkela_wire_14811;
    wire new_Jinkela_wire_11798;
    wire new_Jinkela_wire_8352;
    wire new_Jinkela_wire_20794;
    wire new_Jinkela_wire_16496;
    wire new_Jinkela_wire_16082;
    wire new_Jinkela_wire_20288;
    wire new_Jinkela_wire_18016;
    wire new_Jinkela_wire_7920;
    wire new_Jinkela_wire_12096;
    wire new_Jinkela_wire_20617;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_9381;
    wire _1094_;
    wire new_Jinkela_wire_20338;
    wire new_Jinkela_wire_8234;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_8854;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_13635;
    wire new_Jinkela_wire_13715;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_15394;
    wire new_Jinkela_wire_17222;
    wire new_Jinkela_wire_20843;
    wire new_Jinkela_wire_8573;
    wire _1392_;
    wire new_Jinkela_wire_19844;
    wire new_Jinkela_wire_2534;
    wire new_Jinkela_wire_13094;
    wire new_Jinkela_wire_12258;
    wire new_Jinkela_wire_13587;
    wire new_Jinkela_wire_4533;
    wire new_Jinkela_wire_11153;
    wire new_Jinkela_wire_13056;
    wire new_Jinkela_wire_5867;
    wire new_Jinkela_wire_6597;
    wire new_Jinkela_wire_15695;
    wire new_Jinkela_wire_8259;
    wire new_Jinkela_wire_15382;
    wire new_Jinkela_wire_2507;
    wire new_Jinkela_wire_4331;
    wire new_Jinkela_wire_10808;
    wire new_Jinkela_wire_11772;
    wire new_Jinkela_wire_8664;
    wire new_Jinkela_wire_17329;
    wire new_Jinkela_wire_18862;
    wire new_Jinkela_wire_5779;
    wire new_Jinkela_wire_9266;
    wire new_Jinkela_wire_3315;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_8420;
    wire new_Jinkela_wire_8752;
    wire new_Jinkela_wire_3608;
    wire _1719_;
    wire new_Jinkela_wire_2679;
    wire _1379_;
    wire new_Jinkela_wire_8554;
    wire new_Jinkela_wire_5209;
    wire _1194_;
    wire new_Jinkela_wire_11000;
    wire new_Jinkela_wire_14384;
    wire new_Jinkela_wire_19027;
    wire new_Jinkela_wire_16564;
    wire new_Jinkela_wire_13731;
    wire new_Jinkela_wire_12233;
    wire new_Jinkela_wire_3989;
    wire new_Jinkela_wire_13396;
    wire new_Jinkela_wire_5626;
    wire new_Jinkela_wire_18364;
    wire new_Jinkela_wire_11986;
    wire _0179_;
    wire new_Jinkela_wire_19506;
    wire new_Jinkela_wire_12306;
    wire new_Jinkela_wire_16002;
    wire new_Jinkela_wire_6453;
    wire new_Jinkela_wire_15350;
    wire new_Jinkela_wire_13631;
    wire new_Jinkela_wire_19561;
    wire new_Jinkela_wire_9727;
    wire new_Jinkela_wire_1749;
    wire new_Jinkela_wire_10854;
    wire new_Jinkela_wire_2955;
    wire new_Jinkela_wire_15545;
    wire new_Jinkela_wire_5040;
    wire new_Jinkela_wire_17349;
    wire new_Jinkela_wire_20866;
    wire new_Jinkela_wire_4432;
    wire new_Jinkela_wire_11735;
    wire new_Jinkela_wire_2149;
    wire new_Jinkela_wire_18678;
    wire new_Jinkela_wire_2939;
    wire new_Jinkela_wire_7135;
    wire new_Jinkela_wire_13592;
    wire new_Jinkela_wire_21297;
    wire new_Jinkela_wire_16734;
    wire new_Jinkela_wire_18720;
    wire new_Jinkela_wire_15184;
    wire new_Jinkela_wire_12877;
    wire new_Jinkela_wire_11314;
    wire new_Jinkela_wire_10630;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_4269;
    wire new_Jinkela_wire_8953;
    wire new_Jinkela_wire_21272;
    wire new_Jinkela_wire_12653;
    wire new_Jinkela_wire_18503;
    wire _0275_;
    wire new_Jinkela_wire_2895;
    wire new_Jinkela_wire_20348;
    wire new_Jinkela_wire_17272;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_3636;
    wire new_Jinkela_wire_14801;
    wire new_Jinkela_wire_2812;
    wire new_Jinkela_wire_9942;
    wire new_Jinkela_wire_4730;
    wire new_Jinkela_wire_15179;
    wire new_Jinkela_wire_11521;
    wire _1195_;
    wire new_Jinkela_wire_11857;
    wire new_Jinkela_wire_20529;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_17601;
    wire new_Jinkela_wire_6309;
    wire new_Jinkela_wire_7301;
    wire new_Jinkela_wire_18703;
    wire new_Jinkela_wire_3463;
    wire new_Jinkela_wire_14952;
    wire new_Jinkela_wire_6816;
    wire new_Jinkela_wire_9828;
    wire _1449_;
    wire new_Jinkela_wire_21262;
    wire new_Jinkela_wire_16911;
    wire new_Jinkela_wire_16467;
    wire new_Jinkela_wire_10743;
    wire new_Jinkela_wire_12140;
    wire new_Jinkela_wire_4990;
    wire new_Jinkela_wire_12911;
    wire new_Jinkela_wire_17298;
    wire new_Jinkela_wire_10634;
    wire new_Jinkela_wire_9208;
    wire new_Jinkela_wire_20432;
    wire new_Jinkela_wire_6557;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_7436;
    wire _0660_;
    wire new_Jinkela_wire_20044;
    wire new_Jinkela_wire_6152;
    wire new_Jinkela_wire_1612;
    wire new_Jinkela_wire_10830;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_8417;
    wire new_Jinkela_wire_14844;
    wire new_Jinkela_wire_9311;
    wire new_Jinkela_wire_8646;
    wire _0358_;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_14887;
    wire new_Jinkela_wire_8452;
    wire new_Jinkela_wire_7838;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_13589;
    wire new_Jinkela_wire_5936;
    wire new_Jinkela_wire_10245;
    wire new_Jinkela_wire_19817;
    wire new_Jinkela_wire_3431;
    wire new_Jinkela_wire_4112;
    wire new_Jinkela_wire_16615;
    wire new_Jinkela_wire_10288;
    wire new_Jinkela_wire_6906;
    wire new_Jinkela_wire_19222;
    wire new_Jinkela_wire_6578;
    wire new_Jinkela_wire_3405;
    wire new_Jinkela_wire_17556;
    wire new_Jinkela_wire_5920;
    wire new_Jinkela_wire_12052;
    wire new_Jinkela_wire_7342;
    wire new_Jinkela_wire_18331;
    wire new_Jinkela_wire_15839;
    wire new_Jinkela_wire_20792;
    wire new_Jinkela_wire_7367;
    wire new_Jinkela_wire_19449;
    wire new_Jinkela_wire_17269;
    wire new_Jinkela_wire_20399;
    wire _0595_;
    wire new_Jinkela_wire_15326;
    wire new_Jinkela_wire_12018;
    wire new_Jinkela_wire_3667;
    wire _0585_;
    wire new_Jinkela_wire_20549;
    wire new_Jinkela_wire_3197;
    wire _0039_;
    wire new_Jinkela_wire_15058;
    wire new_Jinkela_wire_9673;
    wire new_Jinkela_wire_10863;
    wire new_Jinkela_wire_6388;
    wire new_Jinkela_wire_13538;
    wire new_Jinkela_wire_19980;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_11123;
    wire new_Jinkela_wire_14336;
    wire new_Jinkela_wire_20988;
    wire new_Jinkela_wire_3098;
    wire new_Jinkela_wire_10891;
    wire new_Jinkela_wire_15273;
    wire new_Jinkela_wire_5608;
    wire new_Jinkela_wire_16308;
    wire new_Jinkela_wire_1737;
    wire _1246_;
    wire new_Jinkela_wire_12656;
    wire new_Jinkela_wire_14543;
    wire new_Jinkela_wire_9871;
    wire new_Jinkela_wire_14051;
    wire new_Jinkela_wire_10894;
    wire new_Jinkela_wire_21105;
    wire new_Jinkela_wire_18585;
    wire _0704_;
    wire new_Jinkela_wire_3935;
    wire new_Jinkela_wire_13165;
    wire new_Jinkela_wire_11488;
    wire new_Jinkela_wire_11114;
    wire new_Jinkela_wire_10165;
    wire new_Jinkela_wire_16645;
    wire new_Jinkela_wire_5230;
    wire new_Jinkela_wire_10117;
    wire new_Jinkela_wire_18365;
    wire _1697_;
    wire new_Jinkela_wire_17777;
    wire new_Jinkela_wire_4804;
    wire new_Jinkela_wire_2305;
    wire new_Jinkela_wire_9006;
    wire new_Jinkela_wire_3219;
    wire new_Jinkela_wire_12843;
    wire _1594_;
    wire new_Jinkela_wire_7715;
    wire new_Jinkela_wire_14863;
    wire new_Jinkela_wire_13160;
    wire new_Jinkela_wire_17314;
    wire _0569_;
    wire new_Jinkela_wire_10342;
    wire new_Jinkela_wire_16778;
    wire new_Jinkela_wire_7644;
    wire new_Jinkela_wire_6712;
    wire new_Jinkela_wire_19242;
    wire new_Jinkela_wire_19697;
    wire new_Jinkela_wire_8662;
    wire new_Jinkela_wire_2351;
    wire new_Jinkela_wire_17829;
    wire new_Jinkela_wire_19009;
    wire new_Jinkela_wire_21009;
    wire new_Jinkela_wire_8161;
    wire new_Jinkela_wire_13718;
    wire new_Jinkela_wire_14907;
    wire new_Jinkela_wire_9288;
    wire new_Jinkela_wire_4094;
    wire new_Jinkela_wire_21025;
    wire new_Jinkela_wire_20439;
    wire new_Jinkela_wire_7968;
    wire new_Jinkela_wire_4784;
    wire new_Jinkela_wire_10681;
    wire new_Jinkela_wire_10502;
    wire _0466_;
    wire new_Jinkela_wire_12484;
    wire new_Jinkela_wire_5766;
    wire _1387_;
    wire new_Jinkela_wire_7383;
    wire new_Jinkela_wire_8642;
    wire new_Jinkela_wire_6641;
    wire new_Jinkela_wire_17300;
    wire new_Jinkela_wire_6707;
    wire new_Jinkela_wire_16543;
    wire new_Jinkela_wire_15230;
    wire new_Jinkela_wire_11845;
    wire new_Jinkela_wire_10877;
    wire new_Jinkela_wire_7265;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_18227;
    wire new_Jinkela_wire_20909;
    wire new_Jinkela_wire_21225;
    wire new_Jinkela_wire_11062;
    wire new_Jinkela_wire_4270;
    wire new_Jinkela_wire_2506;
    wire new_Jinkela_wire_2191;
    wire new_Jinkela_wire_10220;
    wire _1068_;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_10595;
    wire new_Jinkela_wire_8645;
    wire new_Jinkela_wire_20933;
    wire new_Jinkela_wire_19919;
    wire _0926_;
    wire new_Jinkela_wire_16289;
    wire new_Jinkela_wire_11536;
    wire new_Jinkela_wire_1776;
    wire _0258_;
    wire _0367_;
    wire new_Jinkela_wire_18288;
    wire new_Jinkela_wire_5356;
    wire new_Jinkela_wire_16949;
    wire new_Jinkela_wire_10662;
    wire new_Jinkela_wire_18698;
    wire new_Jinkela_wire_11669;
    wire new_Jinkela_wire_10574;
    wire new_Jinkela_wire_13630;
    wire new_Jinkela_wire_14905;
    wire new_Jinkela_wire_3360;
    wire new_Jinkela_wire_16909;
    wire new_Jinkela_wire_5059;
    wire new_Jinkela_wire_4526;
    wire new_Jinkela_wire_8597;
    wire new_Jinkela_wire_14056;
    wire _1074_;
    wire new_Jinkela_wire_16803;
    wire new_Jinkela_wire_5659;
    wire new_Jinkela_wire_11429;
    wire new_Jinkela_wire_18284;
    wire new_Jinkela_wire_14347;
    wire new_Jinkela_wire_4921;
    wire new_Jinkela_wire_2324;
    wire new_Jinkela_wire_14229;
    wire new_Jinkela_wire_15722;
    wire new_Jinkela_wire_17581;
    wire new_Jinkela_wire_18279;
    wire new_Jinkela_wire_6591;
    wire new_Jinkela_wire_11468;
    wire new_Jinkela_wire_13864;
    wire new_Jinkela_wire_12759;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_20798;
    wire new_Jinkela_wire_6269;
    wire new_Jinkela_wire_9452;
    wire new_Jinkela_wire_14092;
    wire new_Jinkela_wire_20554;
    wire new_Jinkela_wire_4364;
    wire new_Jinkela_wire_6354;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_1945;
    wire new_Jinkela_wire_12286;
    wire new_Jinkela_wire_19221;
    wire new_Jinkela_wire_6667;
    wire new_Jinkela_wire_15392;
    wire new_Jinkela_wire_3720;
    wire new_Jinkela_wire_11423;
    wire new_Jinkela_wire_10441;
    wire new_Jinkela_wire_9968;
    wire new_Jinkela_wire_4602;
    wire new_Jinkela_wire_19142;
    wire new_Jinkela_wire_18714;
    wire new_Jinkela_wire_4377;
    wire new_Jinkela_wire_7749;
    wire new_Jinkela_wire_6786;
    wire new_Jinkela_wire_3094;
    wire new_Jinkela_wire_6697;
    wire new_Jinkela_wire_10402;
    wire new_Jinkela_wire_10774;
    wire new_Jinkela_wire_6158;
    wire new_Jinkela_wire_17402;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_11525;
    wire new_Jinkela_wire_18427;
    wire new_Jinkela_wire_15732;
    wire new_Jinkela_wire_21132;
    wire new_Jinkela_wire_15697;
    wire new_Jinkela_wire_17029;
    wire new_Jinkela_wire_13513;
    wire new_Jinkela_wire_14283;
    wire new_Jinkela_wire_7700;
    wire new_Jinkela_wire_10435;
    wire new_Jinkela_wire_16749;
    wire new_Jinkela_wire_19289;
    wire new_Jinkela_wire_12875;
    wire new_Jinkela_wire_6507;
    wire new_Jinkela_wire_20654;
    wire _0439_;
    wire new_Jinkela_wire_8906;
    wire new_Jinkela_wire_3059;
    wire new_Jinkela_wire_14430;
    wire new_Jinkela_wire_6519;
    wire new_Jinkela_wire_8686;
    wire new_Jinkela_wire_11351;
    wire new_Jinkela_wire_15283;
    wire new_Jinkela_wire_4476;
    wire new_Jinkela_wire_11125;
    wire new_Jinkela_wire_19272;
    wire new_Jinkela_wire_7910;
    wire new_Jinkela_wire_19596;
    wire new_Jinkela_wire_3937;
    wire new_Jinkela_wire_19324;
    wire new_Jinkela_wire_10797;
    wire new_Jinkela_wire_8772;
    wire new_Jinkela_wire_17201;
    wire new_Jinkela_wire_3880;
    wire new_Jinkela_wire_19043;
    wire new_Jinkela_wire_20597;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_20545;
    wire new_Jinkela_wire_12972;
    wire new_Jinkela_wire_4008;
    wire new_Jinkela_wire_13131;
    wire new_Jinkela_wire_2650;
    wire new_Jinkela_wire_11073;
    wire new_Jinkela_wire_20353;
    wire new_Jinkela_wire_17039;
    wire new_Jinkela_wire_17774;
    wire new_Jinkela_wire_14147;
    wire new_Jinkela_wire_19592;
    wire new_Jinkela_wire_7190;
    wire _1648_;
    wire new_Jinkela_wire_5918;
    wire new_Jinkela_wire_3507;
    wire new_Jinkela_wire_19547;
    wire new_Jinkela_wire_15848;
    wire new_Jinkela_wire_4214;
    wire _1064_;
    wire new_Jinkela_wire_12680;
    wire new_Jinkela_wire_14742;
    wire new_Jinkela_wire_10466;
    wire new_Jinkela_wire_18636;
    wire new_Jinkela_wire_5057;
    wire new_Jinkela_wire_11345;
    wire new_Jinkela_wire_19039;
    wire new_Jinkela_wire_3921;
    wire new_Jinkela_wire_12367;
    wire new_Jinkela_wire_6993;
    wire new_Jinkela_wire_17842;
    wire new_Jinkela_wire_9702;
    wire new_Jinkela_wire_11711;
    wire new_Jinkela_wire_11118;
    wire new_Jinkela_wire_2741;
    wire new_Jinkela_wire_21097;
    wire new_Jinkela_wire_19279;
    wire new_Jinkela_wire_15423;
    wire new_Jinkela_wire_11978;
    wire new_Jinkela_wire_7434;
    wire new_Jinkela_wire_15694;
    wire new_Jinkela_wire_13510;
    wire new_Jinkela_wire_15027;
    wire new_Jinkela_wire_20283;
    wire new_Jinkela_wire_4221;
    wire new_Jinkela_wire_480;
    wire new_Jinkela_wire_17865;
    wire new_Jinkela_wire_14346;
    wire new_Jinkela_wire_17767;
    wire new_Jinkela_wire_19177;
    wire new_Jinkela_wire_2128;
    wire new_Jinkela_wire_5561;
    wire new_Jinkela_wire_7673;
    wire new_Jinkela_wire_4243;
    wire new_Jinkela_wire_16975;
    wire new_Jinkela_wire_7145;
    wire new_Jinkela_wire_12265;
    wire new_Jinkela_wire_19195;
    wire new_Jinkela_wire_4571;
    wire new_Jinkela_wire_19888;
    wire new_Jinkela_wire_15561;
    wire new_Jinkela_wire_3947;
    wire new_Jinkela_wire_7109;
    wire new_Jinkela_wire_17440;
    wire new_Jinkela_wire_17187;
    wire new_Jinkela_wire_2591;
    wire new_Jinkela_wire_20503;
    wire new_Jinkela_wire_2404;
    wire new_Jinkela_wire_13249;
    wire new_Jinkela_wire_3518;
    wire _0825_;
    wire new_Jinkela_wire_2366;
    wire new_Jinkela_wire_14286;
    wire new_Jinkela_wire_20118;
    wire new_Jinkela_wire_3337;
    wire new_Jinkela_wire_18283;
    wire new_Jinkela_wire_11808;
    wire new_Jinkela_wire_13591;
    wire new_Jinkela_wire_13141;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_18385;
    wire _1308_;
    wire new_Jinkela_wire_14269;
    wire new_Jinkela_wire_19500;
    wire new_Jinkela_wire_3596;
    wire new_Jinkela_wire_18955;
    wire new_Jinkela_wire_6175;
    wire new_Jinkela_wire_18302;
    wire new_Jinkela_wire_5393;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_14408;
    wire new_Jinkela_wire_19060;
    wire new_Jinkela_wire_7366;
    wire new_Jinkela_wire_12319;
    wire new_Jinkela_wire_1506;
    wire new_Jinkela_wire_17082;
    wire new_Jinkela_wire_3157;
    wire new_Jinkela_wire_2648;
    wire new_Jinkela_wire_4469;
    wire new_Jinkela_wire_14819;
    wire new_Jinkela_wire_12768;
    wire new_Jinkela_wire_3959;
    wire new_Jinkela_wire_12334;
    wire new_Jinkela_wire_16087;
    wire _1469_;
    wire new_Jinkela_wire_10702;
    wire new_Jinkela_wire_17406;
    wire new_Jinkela_wire_14062;
    wire new_Jinkela_wire_1224;
    wire new_Jinkela_wire_16254;
    wire new_Jinkela_wire_5168;
    wire new_Jinkela_wire_5791;
    wire new_Jinkela_wire_20161;
    wire new_Jinkela_wire_19247;
    wire new_Jinkela_wire_8997;
    wire _0738_;
    wire new_Jinkela_wire_18926;
    wire new_Jinkela_wire_13911;
    wire new_Jinkela_wire_8307;
    wire new_Jinkela_wire_6780;
    wire new_Jinkela_wire_4464;
    wire new_Jinkela_wire_13218;
    wire new_Jinkela_wire_7615;
    wire _1083_;
    wire new_Jinkela_wire_15043;
    wire new_Jinkela_wire_17075;
    wire new_Jinkela_wire_11572;
    wire new_Jinkela_wire_18944;
    wire new_Jinkela_wire_18960;
    wire new_Jinkela_wire_16330;
    wire _0909_;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_15188;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_5583;
    wire new_Jinkela_wire_12497;
    wire new_Jinkela_wire_16847;
    wire new_Jinkela_wire_9270;
    wire new_Jinkela_wire_4034;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_13327;
    wire _1287_;
    wire new_Jinkela_wire_7264;
    wire new_Jinkela_wire_13360;
    wire new_Jinkela_wire_5467;
    wire new_Jinkela_wire_5424;
    wire new_Jinkela_wire_7390;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_10942;
    wire new_Jinkela_wire_6871;
    wire new_Jinkela_wire_21014;
    wire new_Jinkela_wire_7547;
    wire new_Jinkela_wire_2719;
    wire new_Jinkela_wire_14800;
    wire _0226_;
    wire new_Jinkela_wire_15380;
    wire new_Jinkela_wire_16882;
    wire new_Jinkela_wire_16314;
    wire new_Jinkela_wire_14619;
    wire new_Jinkela_wire_19927;
    wire new_Jinkela_wire_19900;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_4073;
    wire new_Jinkela_wire_10135;
    wire new_Jinkela_wire_19285;
    wire new_Jinkela_wire_15714;
    wire new_Jinkela_wire_17917;
    wire new_Jinkela_wire_2464;
    wire new_Jinkela_wire_9022;
    wire new_Jinkela_wire_9863;
    wire _1177_;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_7621;
    wire new_Jinkela_wire_14685;
    wire new_Jinkela_wire_16302;
    wire new_Jinkela_wire_15622;
    wire new_Jinkela_wire_15605;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_6151;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_11720;
    wire new_Jinkela_wire_18866;
    wire _0410_;
    wire new_Jinkela_wire_18981;
    wire new_Jinkela_wire_16900;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_18121;
    wire new_Jinkela_wire_5633;
    wire new_Jinkela_wire_2287;
    wire new_Jinkela_wire_21259;
    wire new_Jinkela_wire_14260;
    wire new_Jinkela_wire_4811;
    wire new_Jinkela_wire_14696;
    wire new_Jinkela_wire_4774;
    wire new_Jinkela_wire_2341;
    wire new_Jinkela_wire_13383;
    wire new_Jinkela_wire_12977;
    wire new_Jinkela_wire_10652;
    wire new_Jinkela_wire_16794;
    wire new_Jinkela_wire_13575;
    wire new_Jinkela_wire_20316;
    wire new_Jinkela_wire_4901;
    wire new_Jinkela_wire_13863;
    wire new_Jinkela_wire_17499;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_14853;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_21282;
    wire _0235_;
    wire new_Jinkela_wire_5876;
    wire new_Jinkela_wire_10394;
    wire new_Jinkela_wire_7916;
    wire new_Jinkela_wire_3349;
    wire new_Jinkela_wire_4908;
    wire new_Jinkela_wire_12239;
    wire new_Jinkela_wire_6058;
    wire new_Jinkela_wire_8900;
    wire new_Jinkela_wire_2090;
    wire new_Jinkela_wire_21057;
    wire new_Jinkela_wire_16457;
    wire new_Jinkela_wire_17112;
    wire new_Jinkela_wire_8351;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_9354;
    wire new_Jinkela_wire_9467;
    wire new_Jinkela_wire_4808;
    wire new_Jinkela_wire_15369;
    wire new_Jinkela_wire_4546;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_11603;
    wire new_Jinkela_wire_2284;
    wire new_Jinkela_wire_7362;
    wire new_Jinkela_wire_12343;
    wire new_Jinkela_wire_12866;
    wire new_Jinkela_wire_16862;
    wire new_Jinkela_wire_15360;
    wire _0281_;
    wire new_Jinkela_wire_12050;
    wire new_Jinkela_wire_14679;
    wire new_Jinkela_wire_3150;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_20425;
    wire new_Jinkela_wire_3866;
    wire new_Jinkela_wire_9645;
    wire _1235_;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_10591;
    wire _0556_;
    wire new_Jinkela_wire_16062;
    wire new_Jinkela_wire_10993;
    wire new_Jinkela_wire_16034;
    wire new_Jinkela_wire_18255;
    wire new_Jinkela_wire_5764;
    wire new_Jinkela_wire_999;
    wire new_Jinkela_wire_18376;
    wire new_Jinkela_wire_1743;
    wire new_Jinkela_wire_20403;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_6184;
    wire _1044_;
    wire new_Jinkela_wire_18349;
    wire new_Jinkela_wire_2308;
    wire new_Jinkela_wire_1675;
    wire new_Jinkela_wire_2807;
    wire new_Jinkela_wire_1785;
    wire new_Jinkela_wire_13107;
    wire new_Jinkela_wire_9162;
    wire new_Jinkela_wire_6219;
    wire new_Jinkela_wire_7933;
    wire new_Jinkela_wire_19508;
    wire new_Jinkela_wire_13870;
    wire new_Jinkela_wire_3623;
    wire new_Jinkela_wire_18759;
    wire new_Jinkela_wire_8588;
    wire new_Jinkela_wire_19079;
    wire new_Jinkela_wire_14988;
    wire new_Jinkela_wire_8476;
    wire new_Jinkela_wire_12689;
    wire new_Jinkela_wire_3042;
    wire new_Jinkela_wire_17238;
    wire _0680_;
    wire new_Jinkela_wire_20239;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_7038;
    wire new_Jinkela_wire_7596;
    wire new_Jinkela_wire_4584;
    wire new_Jinkela_wire_19955;
    wire new_Jinkela_wire_7712;
    wire new_Jinkela_wire_9121;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_6070;
    wire new_Jinkela_wire_13467;
    wire new_Jinkela_wire_11690;
    wire new_Jinkela_wire_16333;
    wire new_Jinkela_wire_6971;
    wire new_Jinkela_wire_17978;
    wire _0012_;
    wire new_Jinkela_wire_8990;
    wire _1768_;
    wire new_Jinkela_wire_19479;
    wire new_Jinkela_wire_12216;
    wire new_Jinkela_wire_12355;
    wire _0517_;
    wire new_Jinkela_wire_19959;
    wire new_Jinkela_wire_17120;
    wire new_Jinkela_wire_18897;
    wire new_Jinkela_wire_11222;
    wire new_Jinkela_wire_4634;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_20576;
    wire new_Jinkela_wire_18736;
    wire new_Jinkela_wire_12281;
    wire new_Jinkela_wire_20279;
    wire new_Jinkela_wire_6447;
    wire new_Jinkela_wire_21267;
    wire new_Jinkela_wire_17797;
    wire new_Jinkela_wire_15039;
    wire new_Jinkela_wire_6258;
    wire new_Jinkela_wire_17438;
    wire new_Jinkela_wire_20385;
    wire new_Jinkela_wire_2934;
    wire new_Jinkela_wire_11955;
    wire new_Jinkela_wire_11257;
    wire new_Jinkela_wire_10230;
    wire new_Jinkela_wire_13612;
    wire new_Jinkela_wire_6887;
    wire new_Jinkela_wire_14882;
    wire new_Jinkela_wire_2666;
    wire new_Jinkela_wire_15921;
    wire new_Jinkela_wire_6851;
    wire new_Jinkela_wire_15877;
    wire new_Jinkela_wire_21265;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_7494;
    wire new_Jinkela_wire_2800;
    wire new_Jinkela_wire_5114;
    wire new_Jinkela_wire_18013;
    wire new_Jinkela_wire_10760;
    wire new_Jinkela_wire_11959;
    wire new_Jinkela_wire_8534;
    wire new_Jinkela_wire_11990;
    wire new_Jinkela_wire_17999;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_18665;
    wire new_Jinkela_wire_13634;
    wire new_Jinkela_wire_2277;
    wire _0672_;
    wire new_Jinkela_wire_6984;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_18675;
    wire new_Jinkela_wire_18225;
    wire new_Jinkela_wire_3988;
    wire new_Jinkela_wire_6467;
    wire new_Jinkela_wire_3117;
    wire new_Jinkela_wire_11374;
    wire new_Jinkela_wire_11160;
    wire new_Jinkela_wire_17083;
    wire new_Jinkela_wire_15060;
    wire new_Jinkela_wire_12864;
    wire new_Jinkela_wire_16262;
    wire new_Jinkela_wire_3061;
    wire new_Jinkela_wire_5262;
    wire new_Jinkela_wire_17165;
    wire new_Jinkela_wire_6348;
    wire new_Jinkela_wire_8986;
    wire new_Jinkela_wire_19746;
    wire new_Jinkela_wire_13352;
    wire new_Jinkela_wire_5034;
    wire new_Jinkela_wire_10084;
    wire new_Jinkela_wire_4736;
    wire new_Jinkela_wire_8531;
    wire new_Jinkela_wire_10056;
    wire new_Jinkela_wire_5864;
    wire new_Jinkela_wire_5197;
    wire new_Jinkela_wire_14591;
    wire new_Jinkela_wire_15252;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_12964;
    wire new_Jinkela_wire_7799;
    wire new_Jinkela_wire_12615;
    wire new_Jinkela_wire_12963;
    wire new_Jinkela_wire_18488;
    wire new_Jinkela_wire_7504;
    wire new_Jinkela_wire_12722;
    wire new_Jinkela_wire_10725;
    wire new_Jinkela_wire_2152;
    wire new_Jinkela_wire_8373;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_17605;
    wire new_Jinkela_wire_15908;
    wire new_Jinkela_wire_17170;
    wire new_Jinkela_wire_14055;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_7101;
    wire new_Jinkela_wire_19874;
    wire new_Jinkela_wire_11472;
    wire new_Jinkela_wire_1950;
    wire new_Jinkela_wire_2233;
    wire new_Jinkela_wire_16050;
    wire new_Jinkela_wire_11805;
    wire new_Jinkela_wire_11256;
    wire new_Jinkela_wire_20217;
    wire new_Jinkela_wire_4582;
    wire new_Jinkela_wire_15331;
    wire new_net_3942;
    wire new_Jinkela_wire_5455;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_4509;
    wire new_Jinkela_wire_10644;
    wire new_Jinkela_wire_4152;
    wire new_Jinkela_wire_12237;
    wire new_Jinkela_wire_11683;
    wire new_Jinkela_wire_10368;
    wire new_Jinkela_wire_13487;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_16369;
    wire new_Jinkela_wire_18864;
    wire new_Jinkela_wire_4535;
    wire new_Jinkela_wire_6194;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_9705;
    wire new_Jinkela_wire_16789;
    wire new_Jinkela_wire_12601;
    wire new_Jinkela_wire_19670;
    wire new_Jinkela_wire_14593;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_5187;
    wire _0944_;
    wire _0678_;
    wire new_Jinkela_wire_289;
    wire _1661_;
    wire new_Jinkela_wire_15556;
    wire new_Jinkela_wire_4950;
    wire new_Jinkela_wire_2759;
    wire _1610_;
    wire new_Jinkela_wire_14880;
    wire new_Jinkela_wire_4544;
    wire new_Jinkela_wire_19567;
    wire new_Jinkela_wire_21030;
    wire new_Jinkela_wire_13083;
    wire new_Jinkela_wire_5069;
    wire new_Jinkela_wire_2917;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_13814;
    wire new_Jinkela_wire_12387;
    wire new_Jinkela_wire_16881;
    wire new_Jinkela_wire_19042;
    wire new_Jinkela_wire_18793;
    wire new_Jinkela_wire_18344;
    wire _1432_;
    wire _1035_;
    wire new_Jinkela_wire_16805;
    wire new_Jinkela_wire_4568;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_3890;
    wire new_Jinkela_wire_4759;
    wire new_Jinkela_wire_14942;
    wire new_Jinkela_wire_9628;
    wire new_Jinkela_wire_11424;
    wire new_Jinkela_wire_10558;
    wire new_Jinkela_wire_6894;
    wire new_Jinkela_wire_16723;
    wire new_Jinkela_wire_2966;
    wire _0765_;
    wire new_Jinkela_wire_11744;
    wire new_Jinkela_wire_19211;
    wire new_Jinkela_wire_19560;
    wire new_Jinkela_wire_5131;
    wire new_Jinkela_wire_20196;
    wire new_Jinkela_wire_20953;
    wire _0212_;
    wire _0046_;
    wire new_Jinkela_wire_3565;
    wire new_Jinkela_wire_8609;
    wire new_Jinkela_wire_16008;
    wire new_Jinkela_wire_18937;
    wire new_Jinkela_wire_11461;
    wire new_Jinkela_wire_11751;
    wire new_Jinkela_wire_2715;
    wire new_Jinkela_wire_7708;
    wire new_Jinkela_wire_8089;
    wire new_Jinkela_wire_16888;
    wire new_Jinkela_wire_9915;
    wire _0545_;
    wire new_Jinkela_wire_14431;
    wire new_Jinkela_wire_21177;
    wire new_Jinkela_wire_7706;
    wire new_Jinkela_wire_16622;
    wire new_Jinkela_wire_5389;
    wire new_Jinkela_wire_13945;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_18863;
    wire new_Jinkela_wire_14315;
    wire new_Jinkela_wire_8926;
    wire new_Jinkela_wire_16946;
    wire new_Jinkela_wire_2689;
    wire new_Jinkela_wire_5014;
    wire new_Jinkela_wire_4462;
    wire new_Jinkela_wire_2381;
    wire new_Jinkela_wire_12807;
    wire new_Jinkela_wire_20305;
    wire new_Jinkela_wire_18149;
    wire new_Jinkela_wire_8470;
    wire new_Jinkela_wire_18928;
    wire new_Jinkela_wire_16165;
    wire _0424_;
    wire new_Jinkela_wire_11519;
    wire new_Jinkela_wire_16342;
    wire new_Jinkela_wire_6392;
    wire new_Jinkela_wire_12838;
    wire new_Jinkela_wire_5020;
    wire new_Jinkela_wire_12185;
    wire new_Jinkela_wire_7027;
    wire _1368_;
    wire _1425_;
    wire new_Jinkela_wire_14536;
    wire new_Jinkela_wire_13190;
    wire new_Jinkela_wire_18486;
    wire new_Jinkela_wire_18946;
    wire new_Jinkela_wire_2747;
    wire new_Jinkela_wire_9712;
    wire new_Jinkela_wire_18909;
    wire new_Jinkela_wire_12499;
    wire new_Jinkela_wire_21303;
    wire new_Jinkela_wire_15452;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_2962;
    wire new_Jinkela_wire_17199;
    wire new_Jinkela_wire_2256;
    wire new_Jinkela_wire_7357;
    wire new_Jinkela_wire_17351;
    wire new_Jinkela_wire_13862;
    wire new_Jinkela_wire_1727;
    wire new_Jinkela_wire_2801;
    wire new_Jinkela_wire_19842;
    wire new_Jinkela_wire_9290;
    wire _0969_;
    wire new_Jinkela_wire_2634;
    wire new_Jinkela_wire_7834;
    wire new_Jinkela_wire_8506;
    wire new_Jinkela_wire_9109;
    wire new_Jinkela_wire_18641;
    wire new_Jinkela_wire_19320;
    wire new_Jinkela_wire_2834;
    wire new_Jinkela_wire_1939;
    wire new_Jinkela_wire_4866;
    wire new_Jinkela_wire_3209;
    wire new_Jinkela_wire_7561;
    wire new_Jinkela_wire_12600;
    wire new_Jinkela_wire_7624;
    wire new_Jinkela_wire_3779;
    wire new_Jinkela_wire_13014;
    wire new_Jinkela_wire_4617;
    wire new_Jinkela_wire_8172;
    wire new_Jinkela_wire_5730;
    wire new_Jinkela_wire_18322;
    wire new_Jinkela_wire_16773;
    wire new_Jinkela_wire_15244;
    wire new_Jinkela_wire_1725;
    wire _1525_;
    wire new_Jinkela_wire_15660;
    wire new_Jinkela_wire_6946;
    wire new_Jinkela_wire_10384;
    wire new_Jinkela_wire_4431;
    wire new_Jinkela_wire_7501;
    wire new_Jinkela_wire_16137;
    wire new_Jinkela_wire_8287;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_4025;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_15267;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_15505;
    wire new_Jinkela_wire_9232;
    wire new_Jinkela_wire_850;
    wire new_Jinkela_wire_3643;
    wire new_Jinkela_wire_15090;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_3286;
    wire new_Jinkela_wire_17341;
    wire new_Jinkela_wire_17786;
    wire new_Jinkela_wire_16266;
    wire _0887_;
    wire new_Jinkela_wire_16224;
    wire new_Jinkela_wire_14087;
    wire new_Jinkela_wire_17932;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_11517;
    wire new_Jinkela_wire_10102;
    wire new_Jinkela_wire_15373;
    wire new_Jinkela_wire_4088;
    wire _0787_;
    wire new_Jinkela_wire_19418;
    wire _0656_;
    wire new_Jinkela_wire_17127;
    wire new_Jinkela_wire_18662;
    wire new_Jinkela_wire_8974;
    wire new_Jinkela_wire_12774;
    wire new_Jinkela_wire_21213;
    wire new_Jinkela_wire_13301;
    wire new_Jinkela_wire_2099;
    wire _0290_;
    wire new_Jinkela_wire_10210;
    wire new_Jinkela_wire_15083;
    wire _0718_;
    wire new_Jinkela_wire_9618;
    wire new_Jinkela_wire_8389;
    wire new_Jinkela_wire_20638;
    wire new_Jinkela_wire_17625;
    wire new_Jinkela_wire_7468;
    wire new_Jinkela_wire_20420;
    wire new_Jinkela_wire_20748;
    wire new_Jinkela_wire_5025;
    wire new_Jinkela_wire_11331;
    wire new_Jinkela_wire_4953;
    wire new_Jinkela_wire_20227;
    wire new_Jinkela_wire_8260;
    wire new_Jinkela_wire_16717;
    wire new_Jinkela_wire_11576;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_9193;
    wire new_Jinkela_wire_18816;
    wire new_Jinkela_wire_17845;
    wire new_Jinkela_wire_14694;
    wire new_Jinkela_wire_9633;
    wire _0793_;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_17057;
    wire new_Jinkela_wire_2564;
    wire new_Jinkela_wire_5436;
    wire new_Jinkela_wire_19818;
    wire new_Jinkela_wire_15513;
    wire new_Jinkela_wire_14969;
    wire new_Jinkela_wire_17233;
    wire new_Jinkela_wire_16169;
    wire new_Jinkela_wire_12873;
    wire new_Jinkela_wire_15461;
    wire new_Jinkela_wire_13882;
    wire new_Jinkela_wire_19100;
    wire new_Jinkela_wire_6808;
    wire new_Jinkela_wire_20509;
    wire new_Jinkela_wire_5280;
    wire new_Jinkela_wire_19022;
    wire new_Jinkela_wire_11162;
    wire new_Jinkela_wire_13054;
    wire new_Jinkela_wire_18033;
    wire new_Jinkela_wire_11777;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_20026;
    wire new_Jinkela_wire_16972;
    wire new_Jinkela_wire_2482;
    wire new_Jinkela_wire_2363;
    wire new_Jinkela_wire_8437;
    wire new_Jinkela_wire_11577;
    wire new_Jinkela_wire_15673;
    wire new_Jinkela_wire_20133;
    wire new_Jinkela_wire_2995;
    wire new_Jinkela_wire_2555;
    wire new_Jinkela_wire_5650;
    wire new_Jinkela_wire_7274;
    wire new_Jinkela_wire_16390;
    wire new_Jinkela_wire_4574;
    wire new_Jinkela_wire_12878;
    wire new_Jinkela_wire_15138;
    wire new_Jinkela_wire_16115;
    wire _1485_;
    wire _1023_;
    wire new_Jinkela_wire_20004;
    wire new_Jinkela_wire_2775;
    wire new_Jinkela_wire_18544;
    wire new_Jinkela_wire_2743;
    wire new_Jinkela_wire_10464;
    wire new_Jinkela_wire_9711;
    wire new_Jinkela_wire_19198;
    wire new_Jinkela_wire_4622;
    wire new_Jinkela_wire_8756;
    wire new_Jinkela_wire_15871;
    wire new_Jinkela_wire_15705;
    wire new_Jinkela_wire_8486;
    wire new_Jinkela_wire_19184;
    wire new_Jinkela_wire_16986;
    wire new_Jinkela_wire_20593;
    wire _0790_;
    wire new_Jinkela_wire_5002;
    wire new_Jinkela_wire_20551;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_2427;
    wire new_Jinkela_wire_17388;
    wire new_Jinkela_wire_3000;
    wire new_Jinkela_wire_20719;
    wire new_Jinkela_wire_17837;
    wire new_Jinkela_wire_10303;
    wire new_Jinkela_wire_7510;
    wire new_Jinkela_wire_15054;
    wire new_Jinkela_wire_10090;
    wire new_Jinkela_wire_6216;
    wire new_Jinkela_wire_1884;
    wire new_Jinkela_wire_12093;
    wire new_Jinkela_wire_13674;
    wire new_Jinkela_wire_14962;
    wire new_Jinkela_wire_8436;
    wire new_Jinkela_wire_14127;
    wire _1146_;
    wire new_Jinkela_wire_7373;
    wire new_Jinkela_wire_14576;
    wire _0728_;
    wire _1437_;
    wire _0927_;
    wire new_Jinkela_wire_8263;
    wire new_Jinkela_wire_13339;
    wire new_Jinkela_wire_5171;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_9775;
    wire _1466_;
    wire new_Jinkela_wire_3457;
    wire new_Jinkela_wire_11087;
    wire new_Jinkela_wire_16492;
    wire new_Jinkela_wire_15105;
    wire new_Jinkela_wire_16459;
    wire new_Jinkela_wire_4686;
    wire new_Jinkela_wire_3592;
    wire new_Jinkela_wire_6075;
    wire new_Jinkela_wire_12311;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_8767;
    wire new_Jinkela_wire_19839;
    wire new_Jinkela_wire_8495;
    wire new_Jinkela_wire_6290;
    wire new_Jinkela_wire_15817;
    wire new_Jinkela_wire_12550;
    wire _0122_;
    wire new_Jinkela_wire_6339;
    wire new_Jinkela_wire_3089;
    wire new_Jinkela_wire_13473;
    wire new_Jinkela_wire_12046;
    wire new_Jinkela_wire_18672;
    wire new_Jinkela_wire_18515;
    wire new_Jinkela_wire_3577;
    wire new_Jinkela_wire_2018;
    wire new_Jinkela_wire_18389;
    wire new_Jinkela_wire_14435;
    wire new_Jinkela_wire_16368;
    wire new_Jinkela_wire_19435;
    wire new_Jinkela_wire_18904;
    wire new_Jinkela_wire_3229;
    wire new_Jinkela_wire_7400;
    wire new_Jinkela_wire_20481;
    wire new_Jinkela_wire_2173;
    wire _1330_;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_18346;
    wire new_Jinkela_wire_16893;
    wire new_Jinkela_wire_7724;
    wire _1323_;
    wire new_Jinkela_wire_9114;
    wire new_Jinkela_wire_6671;
    wire new_Jinkela_wire_6731;
    wire new_Jinkela_wire_2452;
    wire new_Jinkela_wire_18113;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_7598;
    wire new_Jinkela_wire_16697;
    wire new_Jinkela_wire_21197;
    wire _1518_;
    wire new_Jinkela_wire_21108;
    wire new_Jinkela_wire_14934;
    wire new_Jinkela_wire_18264;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_15759;
    wire new_Jinkela_wire_5505;
    wire new_Jinkela_wire_11375;
    wire new_Jinkela_wire_11499;
    wire new_Jinkela_wire_9632;
    wire new_Jinkela_wire_6310;
    wire new_Jinkela_wire_3277;
    wire new_Jinkela_wire_7774;
    wire new_Jinkela_wire_12760;
    wire new_Jinkela_wire_4044;
    wire new_Jinkela_wire_8764;
    wire new_Jinkela_wire_11065;
    wire new_Jinkela_wire_19048;
    wire new_Jinkela_wire_20446;
    wire new_Jinkela_wire_4111;
    wire new_Jinkela_wire_6782;
    wire new_Jinkela_wire_16066;
    wire new_Jinkela_wire_7016;
    wire new_Jinkela_wire_17995;
    wire new_Jinkela_wire_10250;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_10311;
    wire new_Jinkela_wire_14901;
    wire new_Jinkela_wire_2003;
    wire new_Jinkela_wire_11657;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_20589;
    wire new_Jinkela_wire_19258;
    wire _1062_;
    wire _1665_;
    wire new_Jinkela_wire_5600;
    wire new_Jinkela_wire_17589;
    wire new_Jinkela_wire_14654;
    wire new_Jinkela_wire_14227;
    wire new_Jinkela_wire_19389;
    wire new_Jinkela_wire_10805;
    wire new_Jinkela_wire_8903;
    wire new_Jinkela_wire_6783;
    wire new_Jinkela_wire_21005;
    wire new_Jinkela_wire_10447;
    wire new_Jinkela_wire_15222;
    wire new_Jinkela_wire_8138;
    wire new_Jinkela_wire_20623;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_14207;
    wire new_Jinkela_wire_6574;
    wire new_Jinkela_wire_18629;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_9885;
    wire new_Jinkela_wire_19693;
    wire new_Jinkela_wire_11991;
    wire new_Jinkela_wire_16621;
    wire new_Jinkela_wire_3595;
    wire new_Jinkela_wire_21220;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_11995;
    wire new_Jinkela_wire_7772;
    wire new_Jinkela_wire_4441;
    wire new_Jinkela_wire_20829;
    wire _0280_;
    wire new_Jinkela_wire_5078;
    wire new_Jinkela_wire_16953;
    wire new_Jinkela_wire_6208;
    wire new_Jinkela_wire_9163;
    wire new_Jinkela_wire_5068;
    wire new_Jinkela_wire_19720;
    wire new_Jinkela_wire_15035;
    wire new_Jinkela_wire_18310;
    wire new_Jinkela_wire_8308;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_20053;
    wire new_Jinkela_wire_13824;
    wire new_Jinkela_wire_9275;
    wire _1547_;
    wire new_Jinkela_wire_17487;
    wire new_Jinkela_wire_13845;
    wire new_Jinkela_wire_2069;
    wire new_Jinkela_wire_11236;
    wire new_Jinkela_wire_14372;
    wire new_Jinkela_wire_11660;
    wire _1463_;
    wire new_Jinkela_wire_21100;
    wire _1705_;
    wire new_Jinkela_wire_12757;
    wire new_Jinkela_wire_7397;
    wire new_Jinkela_wire_7606;
    wire new_Jinkela_wire_10176;
    wire new_Jinkela_wire_11231;
    wire _0502_;
    wire new_Jinkela_wire_15028;
    wire new_Jinkela_wire_13379;
    wire new_Jinkela_wire_5015;
    wire new_Jinkela_wire_7105;
    wire new_Jinkela_wire_17846;
    wire new_Jinkela_wire_20175;
    wire new_Jinkela_wire_14205;
    wire new_Jinkela_wire_19078;
    wire new_Jinkela_wire_4076;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_20022;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_9789;
    wire _0551_;
    wire new_Jinkela_wire_15004;
    wire new_Jinkela_wire_9627;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_20436;
    wire new_Jinkela_wire_6777;
    wire _0117_;
    wire new_Jinkela_wire_20835;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_19613;
    wire new_Jinkela_wire_11348;
    wire new_Jinkela_wire_17778;
    wire new_Jinkela_wire_13371;
    wire new_Jinkela_wire_2547;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_21281;
    wire new_Jinkela_wire_20724;
    wire new_Jinkela_wire_17508;
    wire new_Jinkela_wire_13477;
    wire new_Jinkela_wire_19187;
    wire new_Jinkela_wire_14238;
    wire new_Jinkela_wire_13451;
    wire _0352_;
    wire new_Jinkela_wire_8071;
    wire new_Jinkela_wire_10734;
    wire new_Jinkela_wire_6078;
    wire new_Jinkela_wire_6747;
    wire new_Jinkela_wire_16875;
    wire new_Jinkela_wire_17059;
    wire new_Jinkela_wire_14840;
    wire new_Jinkela_wire_10967;
    wire _1602_;
    wire new_Jinkela_wire_13412;
    wire new_Jinkela_wire_9004;
    wire new_Jinkela_wire_7573;
    wire new_Jinkela_wire_11897;
    wire new_Jinkela_wire_15841;
    wire new_Jinkela_wire_12092;
    wire new_Jinkela_wire_4442;
    wire new_Jinkela_wire_263;
    wire new_Jinkela_wire_3265;
    wire _0542_;
    wire new_Jinkela_wire_7982;
    wire new_Jinkela_wire_5822;
    wire new_Jinkela_wire_17426;
    wire new_Jinkela_wire_2950;
    wire new_Jinkela_wire_2738;
    wire new_Jinkela_wire_18482;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_19582;
    wire new_Jinkela_wire_14358;
    wire new_Jinkela_wire_13889;
    wire new_Jinkela_wire_20853;
    wire new_Jinkela_wire_9344;
    wire new_Jinkela_wire_19240;
    wire new_Jinkela_wire_16834;
    wire new_Jinkela_wire_20264;
    wire new_Jinkela_wire_18826;
    wire new_Jinkela_wire_12042;
    wire new_Jinkela_wire_14395;
    wire new_Jinkela_wire_8183;
    wire new_Jinkela_wire_4918;
    wire new_Jinkela_wire_10781;
    wire new_Jinkela_wire_13394;
    wire new_Jinkela_wire_1632;
    wire _1242_;
    wire new_Jinkela_wire_4740;
    wire new_Jinkela_wire_12901;
    wire new_Jinkela_wire_10999;
    wire new_Jinkela_wire_20368;
    wire new_Jinkela_wire_19161;
    wire new_Jinkela_wire_13704;
    wire new_Jinkela_wire_13243;
    wire new_Jinkela_wire_6800;
    wire new_Jinkela_wire_6743;
    wire new_Jinkela_wire_8786;
    wire new_Jinkela_wire_3509;
    wire new_Jinkela_wire_12276;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_2860;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_10361;
    wire new_Jinkela_wire_5137;
    wire new_Jinkela_wire_21066;
    wire new_Jinkela_wire_13432;
    wire new_Jinkela_wire_4717;
    wire new_Jinkela_wire_3942;
    wire new_Jinkela_wire_9955;
    wire new_Jinkela_wire_16104;
    wire new_Jinkela_wire_15049;
    wire new_Jinkela_wire_13677;
    wire new_Jinkela_wire_4238;
    wire new_Jinkela_wire_14406;
    wire new_Jinkela_wire_9473;
    wire new_Jinkela_wire_7169;
    wire new_Jinkela_wire_4605;
    wire new_Jinkela_wire_14314;
    wire new_Jinkela_wire_19427;
    wire new_Jinkela_wire_2705;
    wire new_Jinkela_wire_6050;
    wire new_Jinkela_wire_2402;
    wire new_Jinkela_wire_11010;
    wire new_Jinkela_wire_9833;
    wire new_Jinkela_wire_17533;
    wire _0370_;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_4210;
    wire new_Jinkela_wire_1828;
    wire new_Jinkela_wire_14778;
    wire new_Jinkela_wire_5581;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_21300;
    wire new_Jinkela_wire_20182;
    wire new_Jinkela_wire_13896;
    wire _0213_;
    wire new_Jinkela_wire_7146;
    wire new_Jinkela_wire_8817;
    wire new_Jinkela_wire_4733;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_1816;
    wire new_Jinkela_wire_16679;
    wire new_Jinkela_wire_20741;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_11282;
    wire new_Jinkela_wire_11144;
    wire new_Jinkela_wire_85;
    wire _0184_;
    wire new_Jinkela_wire_16410;
    wire new_Jinkela_wire_12820;
    wire new_Jinkela_wire_14482;
    wire _0776_;
    wire new_Jinkela_wire_20785;
    wire new_Jinkela_wire_5733;
    wire new_Jinkela_wire_9423;
    wire new_Jinkela_wire_17184;
    wire new_Jinkela_wire_3843;
    wire new_Jinkela_wire_16925;
    wire new_Jinkela_wire_17966;
    wire new_Jinkela_wire_15961;
    wire new_Jinkela_wire_8149;
    wire new_Jinkela_wire_9315;
    wire new_Jinkela_wire_1853;
    wire new_Jinkela_wire_6289;
    wire new_Jinkela_wire_16572;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_10386;
    wire _1202_;
    wire new_Jinkela_wire_21159;
    wire _1289_;
    wire new_Jinkela_wire_4149;
    wire new_Jinkela_wire_2385;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_14308;
    wire new_Jinkela_wire_13926;
    wire new_Jinkela_wire_16121;
    wire new_Jinkela_wire_14924;
    wire new_Jinkela_wire_20416;
    wire _0611_;
    wire new_Jinkela_wire_13197;
    wire new_Jinkela_wire_11851;
    wire new_Jinkela_wire_2396;
    wire new_Jinkela_wire_14725;
    wire new_Jinkela_wire_18103;
    wire new_Jinkela_wire_12927;
    wire new_Jinkela_wire_10745;
    wire new_Jinkela_wire_14786;
    wire new_Jinkela_wire_15256;
    wire new_Jinkela_wire_6928;
    wire new_Jinkela_wire_4813;
    wire new_Jinkela_wire_7087;
    wire new_Jinkela_wire_13389;
    wire new_Jinkela_wire_19841;
    wire new_Jinkela_wire_19249;
    wire new_Jinkela_wire_7617;
    wire _0635_;
    wire new_Jinkela_wire_5975;
    wire new_Jinkela_wire_10226;
    wire new_Jinkela_wire_13495;
    wire new_Jinkela_wire_4522;
    wire new_Jinkela_wire_20888;
    wire new_Jinkela_wire_6522;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_13792;
    wire new_Jinkela_wire_21119;
    wire new_Jinkela_wire_9758;
    wire _0567_;
    wire new_Jinkela_wire_12501;
    wire new_Jinkela_wire_3438;
    wire new_Jinkela_wire_17347;
    wire new_Jinkela_wire_9472;
    wire new_Jinkela_wire_6921;
    wire new_Jinkela_wire_5439;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_12975;
    wire new_Jinkela_wire_4282;
    wire new_Jinkela_wire_10527;
    wire new_Jinkela_wire_3727;
    wire new_Jinkela_wire_19348;
    wire new_Jinkela_wire_18791;
    wire new_Jinkela_wire_7333;
    wire new_Jinkela_wire_9449;
    wire _0007_;
    wire new_Jinkela_wire_17109;
    wire new_Jinkela_wire_14928;
    wire new_Jinkela_wire_16179;
    wire new_Jinkela_wire_16055;
    wire new_Jinkela_wire_17087;
    wire new_Jinkela_wire_18156;
    wire new_Jinkela_wire_21110;
    wire new_Jinkela_wire_7103;
    wire new_Jinkela_wire_5453;
    wire new_Jinkela_wire_21087;
    wire _1696_;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_3367;
    wire new_Jinkela_wire_17928;
    wire new_Jinkela_wire_15202;
    wire new_Jinkela_wire_9513;
    wire new_Jinkela_wire_2481;
    wire new_Jinkela_wire_14410;
    wire new_Jinkela_wire_280;
    wire _1157_;
    wire new_Jinkela_wire_8524;
    wire new_Jinkela_wire_18825;
    wire new_Jinkela_wire_4219;
    wire _0693_;
    wire new_Jinkela_wire_2932;
    wire new_Jinkela_wire_9368;
    wire new_Jinkela_wire_14496;
    wire new_Jinkela_wire_10115;
    wire new_Jinkela_wire_2410;
    wire new_Jinkela_wire_18805;
    wire new_Jinkela_wire_10907;
    wire new_Jinkela_wire_5071;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_10680;
    wire new_Jinkela_wire_2109;
    wire new_Jinkela_wire_12028;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_16084;
    wire new_Jinkela_wire_16694;
    wire _1315_;
    wire _0074_;
    wire new_Jinkela_wire_17838;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_1929;
    wire _0173_;
    wire new_Jinkela_wire_2707;
    wire new_Jinkela_wire_3343;
    wire new_Jinkela_wire_16375;
    wire new_Jinkela_wire_15062;
    wire new_Jinkela_wire_4177;
    wire new_Jinkela_wire_3026;
    wire _1047_;
    wire new_Jinkela_wire_11820;
    wire new_Jinkela_wire_21308;
    wire new_Jinkela_wire_8873;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_6715;
    wire new_Jinkela_wire_7000;
    wire new_Jinkela_wire_5324;
    wire new_Jinkela_wire_2058;
    wire new_Jinkela_wire_13308;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_1908;
    wire new_Jinkela_wire_6678;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_5139;
    wire new_Jinkela_wire_12313;
    wire new_Jinkela_wire_3063;
    wire new_Jinkela_wire_17756;
    wire new_Jinkela_wire_18891;
    wire new_Jinkela_wire_10215;
    wire new_Jinkela_wire_10709;
    wire new_Jinkela_wire_13081;
    wire new_Jinkela_wire_13433;
    wire new_Jinkela_wire_12934;
    wire new_Jinkela_wire_9148;
    wire new_Jinkela_wire_1947;
    wire new_Jinkela_wire_9436;
    wire new_Jinkela_wire_4228;
    wire new_Jinkela_wire_4130;
    wire new_Jinkela_wire_10254;
    wire new_Jinkela_wire_11009;
    wire new_Jinkela_wire_5289;
    wire new_Jinkela_wire_15870;
    wire new_Jinkela_wire_5378;
    wire new_Jinkela_wire_8441;
    wire new_Jinkela_wire_20213;
    wire new_Jinkela_wire_19782;
    wire new_Jinkela_wire_4461;
    wire new_Jinkela_wire_16935;
    wire new_Jinkela_wire_11316;
    wire new_Jinkela_wire_7541;
    wire new_Jinkela_wire_15409;
    wire new_Jinkela_wire_3482;
    wire new_Jinkela_wire_18879;
    wire new_Jinkela_wire_1617;
    wire _1588_;
    wire new_Jinkela_wire_5476;
    wire new_Jinkela_wire_16138;
    wire new_Jinkela_wire_3420;
    wire new_Jinkela_wire_12785;
    wire new_Jinkela_wire_14045;
    wire new_Jinkela_wire_16685;
    wire new_Jinkela_wire_15236;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_9189;
    wire new_Jinkela_wire_16781;
    wire new_Jinkela_wire_18860;
    wire new_Jinkela_wire_7270;
    wire new_Jinkela_wire_19761;
    wire new_Jinkela_wire_19648;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_6675;
    wire new_Jinkela_wire_19406;
    wire new_Jinkela_wire_15920;
    wire new_Jinkela_wire_5932;
    wire new_Jinkela_wire_11328;
    wire new_Jinkela_wire_15949;
    wire new_Jinkela_wire_15016;
    wire _1227_;
    wire new_Jinkela_wire_20612;
    wire new_Jinkela_wire_2260;
    wire new_Jinkela_wire_18760;
    wire new_Jinkela_wire_14115;
    wire new_Jinkela_wire_4086;
    wire new_Jinkela_wire_10086;
    wire new_Jinkela_wire_12409;
    wire new_Jinkela_wire_9086;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_66;
    wire _1687_;
    wire new_Jinkela_wire_4963;
    wire new_Jinkela_wire_4896;
    wire new_Jinkela_wire_18337;
    wire new_Jinkela_wire_9057;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_4507;
    wire new_Jinkela_wire_6830;
    wire new_Jinkela_wire_5563;
    wire new_Jinkela_wire_2432;
    wire new_Jinkela_wire_11615;
    wire new_Jinkela_wire_14163;
    wire new_Jinkela_wire_12945;
    wire _0216_;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_10263;
    wire new_Jinkela_wire_14271;
    wire new_Jinkela_wire_4889;
    wire _1164_;
    wire new_Jinkela_wire_1252;
    wire new_Jinkela_wire_11334;
    wire _1283_;
    wire new_Jinkela_wire_5233;
    wire _1423_;
    wire _1731_;
    wire new_Jinkela_wire_13860;
    wire new_Jinkela_wire_18369;
    wire new_Jinkela_wire_10885;
    wire new_Jinkela_wire_19790;
    wire new_Jinkela_wire_7662;
    wire _0821_;
    wire new_Jinkela_wire_4698;
    wire new_Jinkela_wire_10248;
    wire new_Jinkela_wire_8889;
    wire new_Jinkela_wire_15671;
    wire new_Jinkela_wire_20797;
    wire new_Jinkela_wire_9366;
    wire _1139_;
    wire new_Jinkela_wire_12860;
    wire new_Jinkela_wire_11676;
    wire new_Jinkela_wire_14826;
    wire new_Jinkela_wire_20194;
    wire new_Jinkela_wire_7993;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_15143;
    wire new_Jinkela_wire_5841;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_189;
    wire _0407_;
    wire new_Jinkela_wire_16405;
    wire new_Jinkela_wire_8293;
    wire new_Jinkela_wire_6911;
    wire new_Jinkela_wire_19153;
    wire new_Jinkela_wire_19280;
    wire new_Jinkela_wire_19262;
    wire new_Jinkela_wire_14964;
    wire new_Jinkela_wire_8561;
    wire new_Jinkela_wire_9574;
    wire new_Jinkela_wire_9438;
    wire new_Jinkela_wire_7284;
    wire new_Jinkela_wire_14072;
    wire new_Jinkela_wire_9685;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_14363;
    wire new_Jinkela_wire_9226;
    wire new_Jinkela_wire_10219;
    wire new_Jinkela_wire_16598;
    wire new_Jinkela_wire_9380;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_2717;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_20803;
    wire new_Jinkela_wire_16662;
    wire new_Jinkela_wire_17853;
    wire _1190_;
    wire new_Jinkela_wire_2572;
    wire new_Jinkela_wire_8310;
    wire new_Jinkela_wire_14228;
    wire new_Jinkela_wire_12676;
    wire new_Jinkela_wire_11270;
    wire new_Jinkela_wire_16387;
    wire new_Jinkela_wire_11358;
    wire new_Jinkela_wire_10283;
    wire new_Jinkela_wire_5177;
    wire _0662_;
    wire new_Jinkela_wire_5909;
    wire new_Jinkela_wire_16216;
    wire new_Jinkela_wire_15432;
    wire new_Jinkela_wire_5826;
    wire new_Jinkela_wire_6115;
    wire new_Jinkela_wire_6464;
    wire new_net_3956;
    wire new_Jinkela_wire_11928;
    wire new_Jinkela_wire_17018;
    wire new_Jinkela_wire_21285;
    wire new_Jinkela_wire_16704;
    wire new_Jinkela_wire_2332;
    wire _0209_;
    wire new_Jinkela_wire_10535;
    wire new_Jinkela_wire_18549;
    wire new_Jinkela_wire_14588;
    wire new_Jinkela_wire_7536;
    wire new_Jinkela_wire_2477;
    wire new_Jinkela_wire_13057;
    wire new_Jinkela_wire_19948;
    wire _1499_;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_13489;
    wire new_Jinkela_wire_13843;
    wire new_Jinkela_wire_10977;
    wire new_Jinkela_wire_6590;
    wire _1087_;
    wire new_Jinkela_wire_2393;
    wire new_Jinkela_wire_12625;
    wire new_Jinkela_wire_12012;
    wire new_Jinkela_wire_15299;
    wire _0896_;
    wire new_Jinkela_wire_10633;
    wire new_Jinkela_wire_4942;
    wire new_Jinkela_wire_16509;
    wire new_Jinkela_wire_15630;
    wire new_Jinkela_wire_5575;
    wire new_Jinkela_wire_10066;
    wire new_Jinkela_wire_5294;
    wire new_Jinkela_wire_12213;
    wire new_Jinkela_wire_10747;
    wire new_Jinkela_wire_2515;
    wire new_Jinkela_wire_3723;
    wire new_Jinkela_wire_8275;
    wire new_Jinkela_wire_3945;
    wire new_Jinkela_wire_14411;
    wire new_Jinkela_wire_17710;
    wire new_Jinkela_wire_20078;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_14798;
    wire new_Jinkela_wire_11064;
    wire new_Jinkela_wire_10347;
    wire new_Jinkela_wire_18367;
    wire _0578_;
    wire new_Jinkela_wire_16281;
    wire new_Jinkela_wire_19710;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_7588;
    wire new_Jinkela_wire_3440;
    wire _0908_;
    wire new_Jinkela_wire_11285;
    wire new_Jinkela_wire_20939;
    wire new_Jinkela_wire_15007;
    wire new_Jinkela_wire_12157;
    wire new_Jinkela_wire_7654;
    wire new_Jinkela_wire_7472;
    wire new_Jinkela_wire_2897;
    wire new_Jinkela_wire_11889;
    wire new_Jinkela_wire_18213;
    wire new_Jinkela_wire_9884;
    wire new_Jinkela_wire_4405;
    wire new_Jinkela_wire_2183;
    wire new_Jinkela_wire_4935;
    wire new_Jinkela_wire_10034;
    wire new_Jinkela_wire_16450;
    wire new_Jinkela_wire_3002;
    wire new_Jinkela_wire_12546;
    wire new_Jinkela_wire_1048;
    wire _0541_;
    wire new_Jinkela_wire_18615;
    wire new_Jinkela_wire_7059;
    wire new_Jinkela_wire_12075;
    wire new_Jinkela_wire_12816;
    wire new_Jinkela_wire_14032;
    wire new_Jinkela_wire_19165;
    wire _0654_;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_16657;
    wire new_Jinkela_wire_12341;
    wire new_Jinkela_wire_13607;
    wire new_Jinkela_wire_18445;
    wire new_Jinkela_wire_18847;
    wire _1011_;
    wire new_Jinkela_wire_11884;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_2165;
    wire new_Jinkela_wire_9469;
    wire new_Jinkela_wire_8594;
    wire new_Jinkela_wire_11570;
    wire new_Jinkela_wire_18307;
    wire new_Jinkela_wire_7795;
    wire new_Jinkela_wire_11245;
    wire _0010_;
    wire new_Jinkela_wire_6352;
    wire new_Jinkela_wire_4006;
    wire new_Jinkela_wire_2273;
    wire new_Jinkela_wire_20102;
    wire new_Jinkela_wire_19388;
    wire new_Jinkela_wire_7885;
    wire new_Jinkela_wire_12091;
    wire new_Jinkela_wire_18739;
    wire new_Jinkela_wire_14324;
    wire new_Jinkela_wire_10025;
    wire new_Jinkela_wire_13221;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_12116;
    wire new_Jinkela_wire_11938;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_16876;
    wire new_Jinkela_wire_12043;
    wire new_Jinkela_wire_16225;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_21107;
    wire _1215_;
    wire new_Jinkela_wire_2938;
    wire new_Jinkela_wire_8570;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_20065;
    wire new_Jinkela_wire_15485;
    wire new_Jinkela_wire_15133;
    wire new_Jinkela_wire_13937;
    wire new_Jinkela_wire_5352;
    wire new_Jinkela_wire_11275;
    wire new_Jinkela_wire_3780;
    wire new_Jinkela_wire_6426;
    wire new_Jinkela_wire_17639;
    wire new_Jinkela_wire_16244;
    wire _1793_;
    wire new_Jinkela_wire_12593;
    wire new_Jinkela_wire_2150;
    wire new_Jinkela_wire_6281;
    wire new_Jinkela_wire_14586;
    wire new_Jinkela_wire_17645;
    wire new_Jinkela_wire_9383;
    wire new_Jinkela_wire_12404;
    wire new_Jinkela_wire_13711;
    wire new_Jinkela_wire_18762;
    wire new_Jinkela_wire_5976;
    wire new_Jinkela_wire_20728;
    wire new_Jinkela_wire_9249;
    wire new_Jinkela_wire_15985;
    wire new_Jinkela_wire_4181;
    wire new_Jinkela_wire_2480;
    wire _1401_;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_16682;
    wire new_Jinkela_wire_15868;
    wire new_Jinkela_wire_10825;
    wire new_Jinkela_wire_20971;
    wire new_Jinkela_wire_19960;
    wire new_Jinkela_wire_8424;
    wire new_Jinkela_wire_10012;
    wire new_Jinkela_wire_19299;
    wire new_Jinkela_wire_9291;
    wire new_Jinkela_wire_19797;
    wire new_Jinkela_wire_16201;
    wire new_Jinkela_wire_20365;
    wire new_Jinkela_wire_6859;
    wire new_Jinkela_wire_2034;
    wire new_Jinkela_wire_9201;
    wire _0580_;
    wire new_Jinkela_wire_3570;
    wire new_Jinkela_wire_19397;
    wire new_Jinkela_wire_8600;
    wire new_Jinkela_wire_3655;
    wire new_Jinkela_wire_19144;
    wire _1225_;
    wire new_Jinkela_wire_19404;
    wire new_Jinkela_wire_14297;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_19605;
    wire new_Jinkela_wire_17361;
    wire new_Jinkela_wire_13671;
    wire new_Jinkela_wire_12533;
    wire new_Jinkela_wire_1931;
    wire new_Jinkela_wire_10214;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_4272;
    wire new_Jinkela_wire_15911;
    wire new_Jinkela_wire_2096;
    wire new_Jinkela_wire_13724;
    wire new_Jinkela_wire_9160;
    wire new_Jinkela_wire_5644;
    wire new_Jinkela_wire_3620;
    wire new_Jinkela_wire_6652;
    wire new_Jinkela_wire_12604;
    wire new_Jinkela_wire_15228;
    wire new_Jinkela_wire_11318;
    wire new_Jinkela_wire_11072;
    wire new_Jinkela_wire_5761;
    wire new_Jinkela_wire_13426;
    wire new_Jinkela_wire_15550;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_17174;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_13341;
    wire new_Jinkela_wire_13960;
    wire _0129_;
    wire new_Jinkela_wire_16547;
    wire new_Jinkela_wire_19379;
    wire _1671_;
    wire _1167_;
    wire new_Jinkela_wire_1801;
    wire new_Jinkela_wire_8963;
    wire new_Jinkela_wire_16899;
    wire new_Jinkela_wire_11426;
    wire new_Jinkela_wire_12068;
    wire new_Jinkela_wire_9695;
    wire new_Jinkela_wire_18407;
    wire new_Jinkela_wire_11766;
    wire new_Jinkela_wire_15926;
    wire new_Jinkela_wire_7407;
    wire new_Jinkela_wire_20467;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_5416;
    wire new_Jinkela_wire_10326;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_7421;
    wire new_Jinkela_wire_10715;
    wire new_Jinkela_wire_5310;
    wire new_Jinkela_wire_20410;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_7391;
    wire new_Jinkela_wire_16716;
    wire new_Jinkela_wire_2968;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_6900;
    wire _0218_;
    wire new_Jinkela_wire_17711;
    wire new_Jinkela_wire_16680;
    wire _1583_;
    wire new_Jinkela_wire_17741;
    wire new_Jinkela_wire_3410;
    wire new_Jinkela_wire_6935;
    wire new_Jinkela_wire_12966;
    wire new_Jinkela_wire_4490;
    wire new_Jinkela_wire_21012;
    wire new_Jinkela_wire_3965;
    wire new_Jinkela_wire_14695;
    wire new_Jinkela_wire_5516;
    wire _0893_;
    wire new_Jinkela_wire_10767;
    wire new_Jinkela_wire_3190;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_12369;
    wire new_Jinkela_wire_8367;
    wire new_Jinkela_wire_10278;
    wire new_Jinkela_wire_7656;
    wire new_Jinkela_wire_20471;
    wire new_Jinkela_wire_4175;
    wire new_Jinkela_wire_13372;
    wire new_Jinkela_wire_320;
    wire _1220_;
    wire new_Jinkela_wire_14703;
    wire new_Jinkela_wire_4856;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_4520;
    wire new_Jinkela_wire_6611;
    wire new_Jinkela_wire_17759;
    wire new_Jinkela_wire_8055;
    wire new_Jinkela_wire_10826;
    wire new_Jinkela_wire_13232;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_19051;
    wire new_Jinkela_wire_9909;
    wire new_Jinkela_wire_14480;
    wire new_Jinkela_wire_2984;
    wire new_Jinkela_wire_15433;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_10910;
    wire new_Jinkela_wire_2535;
    wire new_Jinkela_wire_17691;
    wire new_Jinkela_wire_6860;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_19806;
    wire new_Jinkela_wire_19958;
    wire new_Jinkela_wire_7852;
    wire _1500_;
    wire new_Jinkela_wire_7175;
    wire new_Jinkela_wire_13785;
    wire new_Jinkela_wire_21289;
    wire new_Jinkela_wire_10921;
    wire new_Jinkela_wire_1782;
    wire new_Jinkela_wire_16379;
    wire new_Jinkela_wire_19702;
    wire new_Jinkela_wire_7846;
    wire new_Jinkela_wire_7310;
    wire new_Jinkela_wire_6869;
    wire new_Jinkela_wire_7306;
    wire _1443_;
    wire new_Jinkela_wire_14938;
    wire new_Jinkela_wire_14226;
    wire new_Jinkela_wire_14661;
    wire new_Jinkela_wire_18627;
    wire new_Jinkela_wire_9198;
    wire new_Jinkela_wire_8397;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_12460;
    wire new_Jinkela_wire_20550;
    wire new_Jinkela_wire_14991;
    wire new_Jinkela_wire_16578;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_16326;
    wire new_Jinkela_wire_17372;
    wire new_Jinkela_wire_2625;
    wire new_Jinkela_wire_5594;
    wire new_Jinkela_wire_12179;
    wire new_Jinkela_wire_16652;
    wire new_Jinkela_wire_8852;
    wire new_Jinkela_wire_11778;
    wire new_Jinkela_wire_9297;
    wire new_Jinkela_wire_12597;
    wire new_Jinkela_wire_15289;
    wire new_Jinkela_wire_11850;
    wire new_Jinkela_wire_18580;
    wire new_Jinkela_wire_19971;
    wire new_Jinkela_wire_19640;
    wire new_Jinkela_wire_2356;
    wire new_Jinkela_wire_20524;
    wire new_Jinkela_wire_4514;
    wire new_Jinkela_wire_12733;
    wire new_Jinkela_wire_6452;
    wire new_Jinkela_wire_19627;
    wire new_Jinkela_wire_3555;
    wire new_Jinkela_wire_19780;
    wire new_Jinkela_wire_2665;
    wire new_Jinkela_wire_15308;
    wire new_Jinkela_wire_3697;
    wire _0890_;
    wire new_Jinkela_wire_12202;
    wire new_Jinkela_wire_14617;
    wire _1268_;
    wire new_Jinkela_wire_5366;
    wire new_Jinkela_wire_3283;
    wire new_Jinkela_wire_15504;
    wire new_Jinkela_wire_8803;
    wire new_Jinkela_wire_14196;
    wire new_Jinkela_wire_16755;
    wire new_Jinkela_wire_3109;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_19794;
    wire new_Jinkela_wire_19879;
    wire new_Jinkela_wire_8608;
    wire new_Jinkela_wire_9517;
    wire _0731_;
    wire new_Jinkela_wire_17013;
    wire new_Jinkela_wire_7964;
    wire new_Jinkela_wire_8072;
    wire new_Jinkela_wire_387;
    wire _1456_;
    wire new_Jinkela_wire_5410;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_13931;
    wire new_Jinkela_wire_8617;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_4404;
    wire new_Jinkela_wire_6882;
    wire new_Jinkela_wire_5473;
    wire new_Jinkela_wire_6745;
    wire new_Jinkela_wire_11911;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_13758;
    wire new_Jinkela_wire_12861;
    wire new_Jinkela_wire_10409;
    wire _0721_;
    wire new_Jinkela_wire_7661;
    wire new_Jinkela_wire_15097;
    wire new_Jinkela_wire_16037;
    wire new_Jinkela_wire_5120;
    wire new_Jinkela_wire_17674;
    wire new_Jinkela_wire_10211;
    wire new_Jinkela_wire_18333;
    wire new_Jinkela_wire_11942;
    wire new_Jinkela_wire_1948;
    wire new_Jinkela_wire_3498;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_11178;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_12815;
    wire new_Jinkela_wire_5398;
    wire new_Jinkela_wire_19003;
    wire _1730_;
    wire new_Jinkela_wire_2355;
    wire new_Jinkela_wire_20628;
    wire new_Jinkela_wire_15085;
    wire new_Jinkela_wire_9687;
    wire new_Jinkela_wire_8910;
    wire new_Jinkela_wire_16154;
    wire _0711_;
    wire new_Jinkela_wire_18833;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_12854;
    wire new_Jinkela_wire_18651;
    wire new_Jinkela_wire_21291;
    wire new_Jinkela_wire_15869;
    wire new_Jinkela_wire_12916;
    wire new_Jinkela_wire_4314;
    wire new_Jinkela_wire_18582;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_10948;
    wire new_Jinkela_wire_18790;
    wire new_Jinkela_wire_8721;
    wire _1645_;
    wire new_Jinkela_wire_8771;
    wire new_Jinkela_wire_5848;
    wire new_Jinkela_wire_4548;
    wire new_Jinkela_wire_19823;
    wire new_Jinkela_wire_6523;
    wire new_Jinkela_wire_13577;
    wire new_Jinkela_wire_19230;
    wire new_Jinkela_wire_17338;
    wire new_Jinkela_wire_20753;
    wire new_Jinkela_wire_19191;
    wire new_Jinkela_wire_5159;
    wire _0283_;
    wire new_Jinkela_wire_7864;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_18943;
    wire new_Jinkela_wire_15497;
    wire new_Jinkela_wire_12428;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_8853;
    wire new_Jinkela_wire_4696;
    wire _1782_;
    wire new_Jinkela_wire_6761;
    wire new_Jinkela_wire_10746;
    wire new_Jinkela_wire_9066;
    wire new_Jinkela_wire_17603;
    wire _0169_;
    wire _0646_;
    wire _0151_;
    wire new_Jinkela_wire_14472;
    wire new_Jinkela_wire_8603;
    wire new_Jinkela_wire_12384;
    wire new_Jinkela_wire_4173;
    wire new_Jinkela_wire_16941;
    wire new_Jinkela_wire_9512;
    wire new_Jinkela_wire_19248;
    wire new_Jinkela_wire_11337;
    wire new_Jinkela_wire_14382;
    wire new_Jinkela_wire_16347;
    wire _0570_;
    wire new_Jinkela_wire_14294;
    wire new_Jinkela_wire_13519;
    wire new_Jinkela_wire_13320;
    wire new_Jinkela_wire_11548;
    wire new_Jinkela_wire_8458;
    wire new_Jinkela_wire_13287;
    wire new_Jinkela_wire_10828;
    wire new_Jinkela_wire_6811;
    wire new_Jinkela_wire_10285;
    wire new_Jinkela_wire_16752;
    wire new_Jinkela_wire_18508;
    wire new_Jinkela_wire_8344;
    wire new_Jinkela_wire_20772;
    wire new_Jinkela_wire_18252;
    wire new_Jinkela_wire_9660;
    wire new_Jinkela_wire_9238;
    wire new_Jinkela_wire_20285;
    wire new_Jinkela_wire_3104;
    wire new_Jinkela_wire_6633;
    wire new_Jinkela_wire_19655;
    wire new_Jinkela_wire_13385;
    wire new_Jinkela_wire_10330;
    wire new_Jinkela_wire_4435;
    wire new_Jinkela_wire_18188;
    wire new_Jinkela_wire_21176;
    wire new_Jinkela_wire_9248;
    wire new_Jinkela_wire_11363;
    wire new_Jinkela_wire_15824;
    wire new_Jinkela_wire_3017;
    wire new_Jinkela_wire_7961;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_17288;
    wire new_Jinkela_wire_8402;
    wire new_Jinkela_wire_20350;
    wire new_Jinkela_wire_16954;
    wire new_Jinkela_wire_18120;
    wire new_Jinkela_wire_16491;
    wire new_Jinkela_wire_14381;
    wire _1200_;
    wire new_Jinkela_wire_10104;
    wire new_Jinkela_wire_13034;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_11471;
    wire new_Jinkela_wire_14376;
    wire new_Jinkela_wire_13440;
    wire new_Jinkela_wire_9800;
    wire new_Jinkela_wire_5234;
    wire new_Jinkela_wire_3048;
    wire new_Jinkela_wire_9320;
    wire _1134_;
    wire new_Jinkela_wire_18539;
    wire new_Jinkela_wire_20448;
    wire new_Jinkela_wire_3302;
    wire new_Jinkela_wire_9435;
    wire new_Jinkela_wire_6636;
    wire _0353_;
    wire new_Jinkela_wire_3481;
    wire new_Jinkela_wire_7647;
    wire new_Jinkela_wire_19199;
    wire new_Jinkela_wire_20643;
    wire new_Jinkela_wire_21324;
    wire new_Jinkela_wire_10506;
    wire new_Jinkela_wire_7365;
    wire _1506_;
    wire new_Jinkela_wire_17210;
    wire new_Jinkela_wire_4394;
    wire new_Jinkela_wire_4877;
    wire new_Jinkela_wire_16715;
    wire new_Jinkela_wire_10829;
    wire new_Jinkela_wire_10292;
    wire new_Jinkela_wire_19064;
    wire new_Jinkela_wire_17699;
    wire _0250_;
    wire new_Jinkela_wire_2219;
    wire new_Jinkela_wire_7262;
    wire new_Jinkela_wire_6427;
    wire new_Jinkela_wire_12114;
    wire new_Jinkela_wire_17804;
    wire new_Jinkela_wire_3539;
    wire new_Jinkela_wire_8279;
    wire new_Jinkela_wire_6981;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_15200;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_16854;
    wire new_Jinkela_wire_10452;
    wire new_Jinkela_wire_17421;
    wire _1442_;
    wire new_Jinkela_wire_6270;
    wire new_Jinkela_wire_4281;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_9182;
    wire new_Jinkela_wire_8366;
    wire _0471_;
    wire _1584_;
    wire new_Jinkela_wire_9253;
    wire new_Jinkela_wire_13104;
    wire new_Jinkela_wire_9343;
    wire new_Jinkela_wire_9798;
    wire new_Jinkela_wire_13858;
    wire new_Jinkela_wire_10737;
    wire new_Jinkela_wire_3651;
    wire new_Jinkela_wire_4820;
    wire new_Jinkela_wire_15721;
    wire new_Jinkela_wire_21221;
    wire new_Jinkela_wire_12255;
    wire new_Jinkela_wire_6944;
    wire _0620_;
    wire new_Jinkela_wire_19708;
    wire new_Jinkela_wire_13033;
    wire new_Jinkela_wire_4635;
    wire new_Jinkela_wire_13145;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_9892;
    wire new_Jinkela_wire_4583;
    wire new_Jinkela_wire_2055;
    wire new_Jinkela_wire_3031;
    wire new_Jinkela_wire_18161;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_11544;
    wire new_Jinkela_wire_2964;
    wire new_Jinkela_wire_6144;
    wire new_Jinkela_wire_10378;
    wire new_Jinkela_wire_3259;
    wire new_Jinkela_wire_3192;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_7643;
    wire new_Jinkela_wire_15386;
    wire _1781_;
    wire new_Jinkela_wire_13750;
    wire new_Jinkela_wire_17232;
    wire new_Jinkela_wire_18754;
    wire new_Jinkela_wire_16507;
    wire new_Jinkela_wire_20201;
    wire new_Jinkela_wire_10111;
    wire new_Jinkela_wire_9516;
    wire new_Jinkela_wire_8827;
    wire _1654_;
    wire new_Jinkela_wire_15248;
    wire new_Jinkela_wire_9530;
    wire new_Jinkela_wire_5411;
    wire new_Jinkela_wire_5568;
    wire new_Jinkela_wire_16582;
    wire new_Jinkela_wire_15514;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_12218;
    wire new_Jinkela_wire_19829;
    wire new_Jinkela_wire_8653;
    wire new_Jinkela_wire_16531;
    wire new_Jinkela_wire_16721;
    wire _1511_;
    wire new_Jinkela_wire_18104;
    wire new_Jinkela_wire_13281;
    wire new_Jinkela_wire_4691;
    wire new_Jinkela_wire_15753;
    wire new_Jinkela_wire_17805;
    wire new_Jinkela_wire_13430;
    wire new_Jinkela_wire_13780;
    wire new_Jinkela_wire_11166;
    wire new_Jinkela_wire_9240;
    wire new_Jinkela_wire_11854;
    wire new_Jinkela_wire_7657;
    wire new_Jinkela_wire_14975;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_5329;
    wire new_Jinkela_wire_19498;
    wire new_Jinkela_wire_18196;
    wire new_Jinkela_wire_9561;
    wire new_Jinkela_wire_8774;
    wire new_Jinkela_wire_2320;
    wire new_Jinkela_wire_19667;
    wire new_Jinkela_wire_11188;
    wire new_Jinkela_wire_18931;
    wire new_Jinkela_wire_16799;
    wire new_Jinkela_wire_16420;
    wire new_Jinkela_wire_2891;
    wire new_Jinkela_wire_8916;
    wire _1213_;
    wire new_Jinkela_wire_7010;
    wire new_Jinkela_wire_4944;
    wire new_Jinkela_wire_2957;
    wire new_Jinkela_wire_18920;
    wire new_Jinkela_wire_7181;
    wire new_Jinkela_wire_12177;
    wire new_Jinkela_wire_4354;
    wire new_Jinkela_wire_8865;
    wire new_Jinkela_wire_14221;
    wire _0387_;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_14341;
    wire new_Jinkela_wire_2846;
    wire new_Jinkela_wire_8451;
    wire _0857_;
    wire new_Jinkela_wire_12949;
    wire new_Jinkela_wire_18041;
    wire new_Jinkela_wire_15489;
    wire new_Jinkela_wire_19386;
    wire new_Jinkela_wire_13541;
    wire _0302_;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_13378;
    wire new_Jinkela_wire_3123;
    wire new_Jinkela_wire_8502;
    wire _0087_;
    wire new_Jinkela_wire_10628;
    wire new_Jinkela_wire_150;
    wire new_Jinkela_wire_11705;
    wire new_Jinkela_wire_6369;
    wire new_Jinkela_wire_17033;
    wire new_Jinkela_wire_10375;
    wire new_Jinkela_wire_19282;
    wire new_Jinkela_wire_4257;
    wire new_Jinkela_wire_5326;
    wire new_Jinkela_wire_1603;
    wire _0612_;
    wire new_Jinkela_wire_6770;
    wire new_Jinkela_wire_17903;
    wire new_Jinkela_wire_16740;
    wire new_Jinkela_wire_19476;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_13481;
    wire new_Jinkela_wire_8358;
    wire new_Jinkela_wire_19011;
    wire new_Jinkela_wire_18087;
    wire new_Jinkela_wire_6368;
    wire new_Jinkela_wire_13560;
    wire new_Jinkela_wire_16427;
    wire new_Jinkela_wire_2027;
    wire _1760_;
    wire new_Jinkela_wire_8763;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_15015;
    wire new_Jinkela_wire_21089;
    wire new_Jinkela_wire_1994;
    wire new_Jinkela_wire_3531;
    wire new_Jinkela_wire_2821;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_8955;
    wire new_Jinkela_wire_20154;
    wire new_Jinkela_wire_8992;
    wire new_Jinkela_wire_2151;
    wire new_Jinkela_wire_15277;
    wire new_Jinkela_wire_12474;
    wire new_Jinkela_wire_10173;
    wire new_Jinkela_wire_4956;
    wire new_Jinkela_wire_11702;
    wire new_Jinkela_wire_13497;
    wire new_Jinkela_wire_13420;
    wire new_Jinkela_wire_15000;
    wire new_Jinkela_wire_2094;
    wire new_Jinkela_wire_11454;
    wire new_Jinkela_wire_20209;
    wire new_Jinkela_wire_5098;
    wire new_Jinkela_wire_18185;
    wire new_Jinkela_wire_18668;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_9203;
    wire new_Jinkela_wire_13737;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_14681;
    wire new_Jinkela_wire_2304;
    wire new_Jinkela_wire_2181;
    wire new_Jinkela_wire_2780;
    wire new_Jinkela_wire_14581;
    wire new_Jinkela_wire_5950;
    wire new_Jinkela_wire_16795;
    wire new_Jinkela_wire_20596;
    wire _0966_;
    wire new_Jinkela_wire_3023;
    wire new_Jinkela_wire_20490;
    wire new_Jinkela_wire_18623;
    wire new_Jinkela_wire_17551;
    wire new_Jinkela_wire_20166;
    wire new_Jinkela_wire_13167;
    wire new_Jinkela_wire_14394;
    wire new_Jinkela_wire_19563;
    wire new_Jinkela_wire_8241;
    wire new_Jinkela_wire_4816;
    wire new_Jinkela_wire_7902;
    wire new_Jinkela_wire_13448;
    wire new_Jinkela_wire_13499;
    wire new_Jinkela_wire_7934;
    wire new_Jinkela_wire_15157;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_801;
    wire _1753_;
    wire new_Jinkela_wire_16012;
    wire _1346_;
    wire new_Jinkela_wire_17500;
    wire new_Jinkela_wire_18093;
    wire new_Jinkela_wire_16093;
    wire new_Jinkela_wire_14967;
    wire new_Jinkela_wire_6044;
    wire new_Jinkela_wire_20949;
    wire new_Jinkela_wire_17868;
    wire _1390_;
    wire new_Jinkela_wire_10179;
    wire new_Jinkela_wire_18940;
    wire new_Jinkela_wire_6490;
    wire new_Jinkela_wire_18251;
    wire new_Jinkela_wire_15391;
    wire new_Jinkela_wire_4639;
    wire new_Jinkela_wire_3650;
    wire new_Jinkela_wire_13113;
    wire new_Jinkela_wire_20293;
    wire new_Jinkela_wire_13409;
    wire new_Jinkela_wire_13940;
    wire new_Jinkela_wire_9918;
    wire new_Jinkela_wire_13935;
    wire new_Jinkela_wire_13180;
    wire new_Jinkela_wire_12178;
    wire new_Jinkela_wire_3846;
    wire new_Jinkela_wire_16348;
    wire new_Jinkela_wire_8084;
    wire new_Jinkela_wire_17883;
    wire new_Jinkela_wire_12241;
    wire new_Jinkela_wire_12416;
    wire new_Jinkela_wire_4283;
    wire new_Jinkela_wire_14075;
    wire new_Jinkela_wire_19341;
    wire new_Jinkela_wire_20594;
    wire new_Jinkela_wire_6744;
    wire new_Jinkela_wire_5609;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_19531;
    wire _1020_;
    wire new_Jinkela_wire_19364;
    wire new_Jinkela_wire_10003;
    wire _1452_;
    wire new_Jinkela_wire_8671;
    wire new_Jinkela_wire_4665;
    wire new_Jinkela_wire_18280;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_5123;
    wire new_Jinkela_wire_5935;
    wire new_Jinkela_wire_16815;
    wire new_Jinkela_wire_9752;
    wire _1644_;
    wire new_Jinkela_wire_19207;
    wire new_Jinkela_wire_12839;
    wire new_Jinkela_wire_17209;
    wire new_Jinkela_wire_14391;
    wire new_Jinkela_wire_20872;
    wire new_Jinkela_wire_14362;
    wire new_Jinkela_wire_12285;
    wire new_Jinkela_wire_9713;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_7433;
    wire new_Jinkela_wire_8654;
    wire new_Jinkela_wire_13455;
    wire new_Jinkela_wire_5190;
    wire new_Jinkela_wire_15674;
    wire new_Jinkela_wire_5874;
    wire new_Jinkela_wire_10676;
    wire _0940_;
    wire new_Jinkela_wire_20614;
    wire new_Jinkela_wire_13932;
    wire new_Jinkela_wire_6988;
    wire new_Jinkela_wire_20934;
    wire _0761_;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_15126;
    wire new_Jinkela_wire_16508;
    wire _0894_;
    wire _1034_;
    wire new_Jinkela_wire_19789;
    wire new_Jinkela_wire_7065;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_18115;
    wire _1207_;
    wire new_Jinkela_wire_5203;
    wire new_Jinkela_wire_13522;
    wire new_Jinkela_wire_15662;
    wire new_Jinkela_wire_6496;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_16525;
    wire new_Jinkela_wire_8863;
    wire new_Jinkela_wire_13988;
    wire new_Jinkela_wire_16673;
    wire new_Jinkela_wire_12858;
    wire new_Jinkela_wire_15766;
    wire new_Jinkela_wire_20670;
    wire new_Jinkela_wire_14879;
    wire new_Jinkela_wire_16739;
    wire new_Jinkela_wire_15178;
    wire new_Jinkela_wire_13283;
    wire new_Jinkela_wire_2062;
    wire new_Jinkela_wire_10424;
    wire new_Jinkela_wire_10351;
    wire new_Jinkela_wire_4555;
    wire new_Jinkela_wire_13876;
    wire new_Jinkela_wire_1967;
    wire new_Jinkela_wire_2752;
    wire new_Jinkela_wire_10236;
    wire new_Jinkela_wire_8347;
    wire new_Jinkela_wire_20242;
    wire new_Jinkela_wire_13375;
    wire new_Jinkela_wire_4010;
    wire new_Jinkela_wire_7288;
    wire new_Jinkela_wire_17342;
    wire new_Jinkela_wire_1591;
    wire new_Jinkela_wire_12166;
    wire new_Jinkela_wire_3855;
    wire new_Jinkela_wire_6273;
    wire new_Jinkela_wire_17203;
    wire new_Jinkela_wire_20744;
    wire new_Jinkela_wire_9938;
    wire new_Jinkela_wire_11631;
    wire new_Jinkela_wire_12162;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_15520;
    wire new_Jinkela_wire_11048;
    wire new_Jinkela_wire_18424;
    wire new_Jinkela_wire_3003;
    wire new_Jinkela_wire_1486;
    wire _1058_;
    wire new_Jinkela_wire_15453;
    wire new_Jinkela_wire_20701;
    wire new_Jinkela_wire_5206;
    wire _0627_;
    wire new_Jinkela_wire_14697;
    wire new_Jinkela_wire_12248;
    wire new_Jinkela_wire_19384;
    wire new_Jinkela_wire_19503;
    wire _1488_;
    wire new_Jinkela_wire_4970;
    wire new_Jinkela_wire_11214;
    wire new_Jinkela_wire_17262;
    wire new_Jinkela_wire_5104;
    wire new_Jinkela_wire_2562;
    wire new_Jinkela_wire_5952;
    wire new_Jinkela_wire_21010;
    wire new_Jinkela_wire_20635;
    wire new_Jinkela_wire_10748;
    wire new_Jinkela_wire_20076;
    wire new_Jinkela_wire_5829;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_13093;
    wire new_Jinkela_wire_7246;
    wire new_Jinkela_wire_8165;
    wire new_Jinkela_wire_6635;
    wire _0064_;
    wire new_Jinkela_wire_1993;
    wire new_Jinkela_wire_18152;
    wire new_Jinkela_wire_18396;
    wire new_Jinkela_wire_20874;
    wire new_Jinkela_wire_17404;
    wire new_Jinkela_wire_16163;
    wire new_Jinkela_wire_5632;
    wire new_Jinkela_wire_12801;
    wire new_Jinkela_wire_5396;
    wire new_Jinkela_wire_12450;
    wire _1350_;
    wire _0876_;
    wire new_Jinkela_wire_5681;
    wire new_Jinkela_wire_20407;
    wire _0794_;
    wire new_Jinkela_wire_9462;
    wire new_Jinkela_wire_2585;
    wire _1803_;
    wire new_Jinkela_wire_10655;
    wire new_Jinkela_wire_2140;
    wire new_Jinkela_wire_13887;
    wire new_Jinkela_wire_3908;
    wire new_Jinkela_wire_17214;
    wire _0334_;
    wire new_Jinkela_wire_12315;
    wire new_Jinkela_wire_3050;
    wire new_Jinkela_wire_17378;
    wire new_Jinkela_wire_2209;
    wire new_Jinkela_wire_5921;
    wire new_Jinkela_wire_8999;
    wire new_Jinkela_wire_19923;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_13018;
    wire new_Jinkela_wire_12541;
    wire new_Jinkela_wire_7448;
    wire new_Jinkela_wire_7512;
    wire new_Jinkela_wire_17897;
    wire _1607_;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_18077;
    wire new_Jinkela_wire_5781;
    wire new_Jinkela_wire_4536;
    wire new_Jinkela_wire_14320;
    wire new_Jinkela_wire_8819;
    wire new_Jinkela_wire_3681;
    wire new_Jinkela_wire_9625;
    wire new_Jinkela_wire_20199;
    wire new_Jinkela_wire_20462;
    wire new_Jinkela_wire_11828;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_19088;
    wire new_Jinkela_wire_19411;
    wire new_Jinkela_wire_12346;
    wire new_Jinkela_wire_15835;
    wire _1689_;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_15131;
    wire new_Jinkela_wire_4417;
    wire new_Jinkela_wire_20896;
    wire new_Jinkela_wire_7893;
    wire _1014_;
    wire new_Jinkela_wire_17302;
    wire _0204_;
    wire new_Jinkela_wire_9437;
    wire new_Jinkela_wire_19662;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_20068;
    wire new_Jinkela_wire_18062;
    wire new_Jinkela_wire_20077;
    wire new_Jinkela_wire_19201;
    wire new_Jinkela_wire_14452;
    wire new_Jinkela_wire_19869;
    wire new_Jinkela_wire_15661;
    wire new_Jinkela_wire_15981;
    wire new_Jinkela_wire_18730;
    wire new_Jinkela_wire_15297;
    wire new_Jinkela_wire_13017;
    wire new_Jinkela_wire_9689;
    wire new_Jinkela_wire_7187;
    wire new_Jinkela_wire_7887;
    wire new_Jinkela_wire_4318;
    wire new_Jinkela_wire_9972;
    wire new_Jinkela_wire_14784;
    wire new_Jinkela_wire_15038;
    wire new_Jinkela_wire_10109;
    wire new_Jinkela_wire_5555;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_9555;
    wire new_Jinkela_wire_6451;
    wire new_Jinkela_wire_14091;
    wire new_Jinkela_wire_18381;
    wire new_Jinkela_wire_18078;
    wire new_Jinkela_wire_14013;
    wire new_Jinkela_wire_12701;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_9690;
    wire new_Jinkela_wire_6629;
    wire new_Jinkela_wire_16418;
    wire new_Jinkela_wire_20611;
    wire new_Jinkela_wire_21317;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_13994;
    wire new_Jinkela_wire_10150;
    wire new_Jinkela_wire_15736;
    wire new_Jinkela_wire_17770;
    wire new_Jinkela_wire_2916;
    wire new_Jinkela_wire_5737;
    wire new_Jinkela_wire_2448;
    wire new_Jinkela_wire_7502;
    wire new_Jinkela_wire_20606;
    wire new_Jinkela_wire_16148;
    wire new_Jinkela_wire_4268;
    wire new_Jinkela_wire_19569;
    wire new_Jinkela_wire_19455;
    wire new_Jinkela_wire_15677;
    wire new_Jinkela_wire_16446;
    wire _0669_;
    wire new_Jinkela_wire_7489;
    wire new_Jinkela_wire_3355;
    wire new_Jinkela_wire_3851;
    wire new_Jinkela_wire_17273;
    wire new_Jinkela_wire_10983;
    wire new_Jinkela_wire_8387;
    wire new_Jinkela_wire_17676;
    wire new_Jinkela_wire_9329;
    wire new_Jinkela_wire_17787;
    wire new_Jinkela_wire_13410;
    wire new_Jinkela_wire_12268;
    wire new_Jinkela_wire_17884;
    wire new_Jinkela_wire_14689;
    wire new_Jinkela_wire_19307;
    wire new_Jinkela_wire_7073;
    wire new_Jinkela_wire_10476;
    wire new_Jinkela_wire_14323;
    wire new_Jinkela_wire_8907;
    wire new_Jinkela_wire_14673;
    wire new_Jinkela_wire_5823;
    wire new_Jinkela_wire_8858;
    wire new_Jinkela_wire_8822;
    wire new_Jinkela_wire_19723;
    wire new_Jinkela_wire_9082;
    wire new_Jinkela_wire_13203;
    wire new_Jinkela_wire_7737;
    wire new_Jinkela_wire_5661;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_7430;
    wire new_Jinkela_wire_19130;
    wire new_Jinkela_wire_3610;
    wire new_Jinkela_wire_10575;
    wire new_Jinkela_wire_18064;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_8378;
    wire new_Jinkela_wire_5968;
    wire new_Jinkela_wire_15099;
    wire new_Jinkela_wire_9154;
    wire _1439_;
    wire new_Jinkela_wire_16649;
    wire new_Jinkela_wire_14128;
    wire _0150_;
    wire new_Jinkela_wire_20867;
    wire new_Jinkela_wire_16011;
    wire new_Jinkela_wire_3087;
    wire new_Jinkela_wire_14712;
    wire _1795_;
    wire new_Jinkela_wire_3338;
    wire new_Jinkela_wire_10638;
    wire _1187_;
    wire new_Jinkela_wire_17318;
    wire new_Jinkela_wire_10411;
    wire new_Jinkela_wire_6999;
    wire new_Jinkela_wire_19671;
    wire new_Jinkela_wire_7204;
    wire _0230_;
    wire new_Jinkela_wire_13848;
    wire _1054_;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_11659;
    wire new_Jinkela_wire_3548;
    wire new_Jinkela_wire_14636;
    wire new_Jinkela_wire_1258;
    wire _0522_;
    wire new_Jinkela_wire_9258;
    wire new_Jinkela_wire_3466;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_20525;
    wire new_Jinkela_wire_6471;
    wire new_Jinkela_wire_7702;
    wire new_Jinkela_wire_16228;
    wire new_Jinkela_wire_10457;
    wire new_Jinkela_wire_12922;
    wire new_Jinkela_wire_9501;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_20526;
    wire new_Jinkela_wire_10541;
    wire new_Jinkela_wire_15578;
    wire new_Jinkela_wire_13947;
    wire new_Jinkela_wire_2994;
    wire new_Jinkela_wire_13553;
    wire new_Jinkela_wire_15749;
    wire new_Jinkela_wire_12562;
    wire new_Jinkela_wire_3587;
    wire new_Jinkela_wire_8113;
    wire new_Jinkela_wire_8124;
    wire new_Jinkela_wire_2575;
    wire new_Jinkela_wire_9804;
    wire new_Jinkela_wire_2954;
    wire new_Jinkela_wire_19256;
    wire new_Jinkela_wire_8112;
    wire new_Jinkela_wire_18988;
    wire new_Jinkela_wire_13055;
    wire _0131_;
    wire new_Jinkela_wire_13829;
    wire new_Jinkela_wire_3715;
    wire _1257_;
    wire new_Jinkela_wire_5488;
    wire new_Jinkela_wire_12473;
    wire new_Jinkela_wire_17137;
    wire new_Jinkela_wire_20811;
    wire new_Jinkela_wire_2348;
    wire new_Jinkela_wire_12697;
    wire new_Jinkela_wire_19636;
    wire new_Jinkela_wire_10238;
    wire new_Jinkela_wire_10640;
    wire new_Jinkela_wire_3635;
    wire _0730_;
    wire new_Jinkela_wire_6920;
    wire new_Jinkela_wire_12530;
    wire new_Jinkela_wire_2907;
    wire new_Jinkela_wire_19527;
    wire new_Jinkela_wire_17186;
    wire _1234_;
    wire new_Jinkela_wire_18774;
    wire new_Jinkela_wire_1144;
    wire _0557_;
    wire new_Jinkela_wire_7215;
    wire new_Jinkela_wire_7326;
    wire new_Jinkela_wire_14276;
    wire new_Jinkela_wire_17752;
    wire new_Jinkela_wire_14605;
    wire new_Jinkela_wire_4503;
    wire new_Jinkela_wire_7449;
    wire new_Jinkela_wire_11667;
    wire new_Jinkela_wire_4905;
    wire new_Jinkela_wire_11762;
    wire new_Jinkela_wire_9931;
    wire new_Jinkela_wire_14518;
    wire new_Jinkela_wire_20268;
    wire new_Jinkela_wire_10811;
    wire new_Jinkela_wire_16021;
    wire new_Jinkela_wire_10463;
    wire new_Jinkela_wire_12479;
    wire new_Jinkela_wire_4974;
    wire new_Jinkela_wire_3470;
    wire new_Jinkela_wire_14951;
    wire _0552_;
    wire _1276_;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_10445;
    wire new_Jinkela_wire_4007;
    wire new_Jinkela_wire_15828;
    wire _1049_;
    wire new_Jinkela_wire_14970;
    wire new_Jinkela_wire_5481;
    wire new_Jinkela_wire_18978;
    wire _0752_;
    wire new_Jinkela_wire_19695;
    wire new_Jinkela_wire_20319;
    wire new_Jinkela_wire_4561;
    wire _0082_;
    wire new_Jinkela_wire_6201;
    wire new_Jinkela_wire_8625;
    wire new_Jinkela_wire_13714;
    wire new_Jinkela_wire_3850;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_15468;
    wire new_Jinkela_wire_13776;
    wire new_Jinkela_wire_13579;
    wire new_Jinkela_wire_7681;
    wire _1709_;
    wire new_Jinkela_wire_20375;
    wire new_Jinkela_wire_13330;
    wire new_Jinkela_wire_20479;
    wire new_Jinkela_wire_16430;
    wire new_Jinkela_wire_16463;
    wire new_Jinkela_wire_11787;
    wire new_Jinkela_wire_14469;
    wire new_Jinkela_wire_17725;
    wire new_Jinkela_wire_20679;
    wire new_Jinkela_wire_8002;
    wire new_Jinkela_wire_4125;
    wire _0364_;
    wire new_Jinkela_wire_10080;
    wire new_Jinkela_wire_10331;
    wire new_Jinkela_wire_4725;
    wire new_Jinkela_wire_2228;
    wire _1311_;
    wire new_Jinkela_wire_13936;
    wire new_Jinkela_wire_19224;
    wire new_Jinkela_wire_3503;
    wire new_Jinkela_wire_9309;
    wire _1495_;
    wire new_Jinkela_wire_3782;
    wire new_Jinkela_wire_20519;
    wire new_Jinkela_wire_3305;
    wire new_Jinkela_wire_18568;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_5288;
    wire new_Jinkela_wire_8466;
    wire _0808_;
    wire new_Jinkela_wire_5871;
    wire _0084_;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_2508;
    wire new_Jinkela_wire_5180;
    wire new_Jinkela_wire_6996;
    wire new_Jinkela_wire_5012;
    wire new_Jinkela_wire_18681;
    wire new_Jinkela_wire_15321;
    wire new_Jinkela_wire_8869;
    wire new_Jinkela_wire_5321;
    wire new_Jinkela_wire_14417;
    wire new_Jinkela_wire_15328;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_15245;
    wire new_Jinkela_wire_5688;
    wire new_Jinkela_wire_19112;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_20063;
    wire new_Jinkela_wire_15793;
    wire new_Jinkela_wire_5383;
    wire new_Jinkela_wire_5706;
    wire new_Jinkela_wire_8249;
    wire _1724_;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_19621;
    wire new_Jinkela_wire_20769;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_2344;
    wire new_Jinkela_wire_1847;
    wire new_Jinkela_wire_2609;
    wire new_Jinkela_wire_16273;
    wire new_Jinkela_wire_12136;
    wire new_Jinkela_wire_17977;
    wire new_Jinkela_wire_19730;
    wire new_Jinkela_wire_8887;
    wire new_Jinkela_wire_7179;
    wire new_Jinkela_wire_15425;
    wire new_Jinkela_wire_20321;
    wire new_Jinkela_wire_18282;
    wire new_Jinkela_wire_5578;
    wire new_Jinkela_wire_6649;
    wire new_Jinkela_wire_11412;
    wire new_Jinkela_wire_7405;
    wire new_Jinkela_wire_20123;
    wire new_Jinkela_wire_10099;
    wire new_Jinkela_wire_4180;
    wire new_Jinkela_wire_5892;
    wire new_Jinkela_wire_20292;
    wire new_Jinkela_wire_20029;
    wire new_Jinkela_wire_11754;
    wire new_Jinkela_wire_5728;
    wire new_Jinkela_wire_7947;
    wire new_Jinkela_wire_11449;
    wire new_Jinkela_wire_16764;
    wire new_Jinkela_wire_20255;
    wire new_Jinkela_wire_18566;
    wire _0303_;
    wire _1416_;
    wire new_Jinkela_wire_855;
    wire _0031_;
    wire new_Jinkela_wire_11671;
    wire new_Jinkela_wire_13076;
    wire new_Jinkela_wire_10639;
    wire new_Jinkela_wire_12432;
    wire new_Jinkela_wire_9393;
    wire new_Jinkela_wire_15169;
    wire new_Jinkela_wire_8099;
    wire new_Jinkela_wire_5678;
    wire new_Jinkela_wire_15152;
    wire new_Jinkela_wire_19855;
    wire new_Jinkela_wire_15208;
    wire new_Jinkela_wire_14794;
    wire new_Jinkela_wire_8610;
    wire new_Jinkela_wire_12348;
    wire new_Jinkela_wire_7542;
    wire _1095_;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_18370;
    wire new_Jinkela_wire_1913;
    wire new_Jinkela_wire_19458;
    wire new_Jinkela_wire_3984;
    wire new_Jinkela_wire_20684;
    wire new_Jinkela_wire_1753;
    wire _1067_;
    wire new_Jinkela_wire_18030;
    wire new_Jinkela_wire_11094;
    wire new_Jinkela_wire_10296;
    wire new_Jinkela_wire_2080;
    wire new_Jinkela_wire_17619;
    wire _0827_;
    wire new_Jinkela_wire_8739;
    wire new_Jinkela_wire_8073;
    wire new_Jinkela_wire_8285;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_15439;
    wire _1520_;
    wire new_Jinkela_wire_11002;
    wire new_Jinkela_wire_16933;
    wire new_Jinkela_wire_19911;
    wire _1670_;
    wire new_Jinkela_wire_8513;
    wire new_Jinkela_wire_5268;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_5341;
    wire new_Jinkela_wire_17103;
    wire new_Jinkela_wire_15929;
    wire new_Jinkela_wire_19944;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_3186;
    wire new_Jinkela_wire_4393;
    wire new_Jinkela_wire_12906;
    wire new_Jinkela_wire_8800;
    wire new_Jinkela_wire_7506;
    wire _1745_;
    wire new_Jinkela_wire_18293;
    wire new_Jinkela_wire_5364;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_3492;
    wire new_Jinkela_wire_11297;
    wire new_Jinkela_wire_17510;
    wire new_Jinkela_wire_4333;
    wire _1805_;
    wire new_Jinkela_wire_11229;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_16407;
    wire new_Jinkela_wire_18634;
    wire new_Jinkela_wire_15145;
    wire new_Jinkela_wire_12915;
    wire new_Jinkela_wire_5983;
    wire _0768_;
    wire new_Jinkela_wire_13268;
    wire new_Jinkela_wire_18100;
    wire new_Jinkela_wire_19264;
    wire new_Jinkela_wire_2969;
    wire new_Jinkela_wire_3490;
    wire new_Jinkela_wire_12378;
    wire new_Jinkela_wire_11477;
    wire new_Jinkela_wire_2197;
    wire new_Jinkela_wire_19330;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_4703;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_6361;
    wire _1815_;
    wire new_Jinkela_wire_18277;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_14904;
    wire new_Jinkela_wire_12076;
    wire _0514_;
    wire _1723_;
    wire new_Jinkela_wire_6763;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_13540;
    wire new_Jinkela_wire_7640;
    wire _1115_;
    wire new_Jinkela_wire_14318;
    wire new_Jinkela_wire_2215;
    wire new_Jinkela_wire_7467;
    wire new_Jinkela_wire_4688;
    wire new_Jinkela_wire_18462;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_8998;
    wire new_Jinkela_wire_18266;
    wire new_Jinkela_wire_10780;
    wire new_Jinkela_wire_6159;
    wire new_Jinkela_wire_12874;
    wire new_Jinkela_wire_14746;
    wire new_Jinkela_wire_13602;
    wire new_Jinkela_wire_9730;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_9540;
    wire new_Jinkela_wire_20850;
    wire new_Jinkela_wire_16906;
    wire _0780_;
    wire new_Jinkela_wire_14558;
    wire new_Jinkela_wire_8137;
    wire new_Jinkela_wire_2113;
    wire new_Jinkela_wire_5720;
    wire new_Jinkela_wire_19337;
    wire new_Jinkela_wire_19998;
    wire new_Jinkela_wire_4413;
    wire new_Jinkela_wire_19014;
    wire new_Jinkela_wire_20734;
    wire new_Jinkela_wire_9468;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_18297;
    wire new_Jinkela_wire_20924;
    wire new_Jinkela_wire_18220;
    wire new_Jinkela_wire_17543;
    wire new_Jinkela_wire_14939;
    wire new_Jinkela_wire_3158;
    wire new_Jinkela_wire_15371;
    wire new_Jinkela_wire_11998;
    wire new_Jinkela_wire_17538;
    wire new_Jinkela_wire_17412;
    wire new_Jinkela_wire_18781;
    wire new_Jinkela_wire_16400;
    wire new_Jinkela_wire_15587;
    wire new_Jinkela_wire_8716;
    wire new_Jinkela_wire_6955;
    wire new_Jinkela_wire_108;
    wire _1552_;
    wire new_Jinkela_wire_18701;
    wire new_Jinkela_wire_20546;
    wire new_Jinkela_wire_11946;
    wire new_Jinkela_wire_10319;
    wire new_Jinkela_wire_10069;
    wire new_Jinkela_wire_19400;
    wire new_Jinkela_wire_16080;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_18753;
    wire new_Jinkela_wire_8056;
    wire new_Jinkela_wire_11307;
    wire new_Jinkela_wire_1541;
    wire _0217_;
    wire new_Jinkela_wire_18932;
    wire new_Jinkela_wire_18467;
    wire new_Jinkela_wire_19787;
    wire new_Jinkela_wire_10027;
    wire new_Jinkela_wire_20688;
    wire new_Jinkela_wire_3816;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_20192;
    wire new_Jinkela_wire_12634;
    wire new_Jinkela_wire_15737;
    wire new_Jinkela_wire_3280;
    wire new_Jinkela_wire_21175;
    wire new_Jinkela_wire_2196;
    wire new_Jinkela_wire_20225;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_19202;
    wire new_Jinkela_wire_2606;
    wire new_Jinkela_wire_6333;
    wire new_Jinkela_wire_4786;
    wire new_Jinkela_wire_9741;
    wire new_Jinkela_wire_4185;
    wire new_Jinkela_wire_9125;
    wire new_Jinkela_wire_11038;
    wire _0963_;
    wire new_Jinkela_wire_3290;
    wire new_Jinkela_wire_6627;
    wire new_Jinkela_wire_16367;
    wire new_Jinkela_wire_13914;
    wire new_Jinkela_wire_8648;
    wire _1121_;
    wire new_Jinkela_wire_6238;
    wire _1475_;
    wire new_Jinkela_wire_20808;
    wire new_Jinkela_wire_3923;
    wire new_Jinkela_wire_6251;
    wire new_Jinkela_wire_17192;
    wire new_Jinkela_wire_3534;
    wire new_Jinkela_wire_8446;
    wire new_Jinkela_wire_9421;
    wire new_Jinkela_wire_12294;
    wire new_Jinkela_wire_11034;
    wire new_Jinkela_wire_19862;
    wire new_Jinkela_wire_17014;
    wire new_Jinkela_wire_3495;
    wire new_Jinkela_wire_9622;
    wire new_Jinkela_wire_11860;
    wire new_Jinkela_wire_6154;
    wire _0596_;
    wire new_Jinkela_wire_11634;
    wire new_Jinkela_wire_5625;
    wire new_Jinkela_wire_17571;
    wire new_Jinkela_wire_10460;
    wire new_Jinkela_wire_7009;
    wire new_Jinkela_wire_10597;
    wire new_Jinkela_wire_8191;
    wire new_Jinkela_wire_8218;
    wire new_Jinkela_wire_20770;
    wire new_Jinkela_wire_11717;
    wire _0785_;
    wire new_Jinkela_wire_16461;
    wire new_Jinkela_wire_19703;
    wire new_Jinkela_wire_5265;
    wire new_Jinkela_wire_2389;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_16112;
    wire new_Jinkela_wire_4340;
    wire new_Jinkela_wire_12806;
    wire new_Jinkela_wire_19872;
    wire new_Jinkela_wire_11172;
    wire new_Jinkela_wire_11941;
    wire new_Jinkela_wire_17629;
    wire new_Jinkela_wire_21305;
    wire new_Jinkela_wire_14365;
    wire new_Jinkela_wire_19543;
    wire new_Jinkela_wire_11013;
    wire new_Jinkela_wire_15100;
    wire new_Jinkela_wire_18838;
    wire new_Jinkela_wire_9809;
    wire new_Jinkela_wire_4513;
    wire new_Jinkela_wire_13404;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_11806;
    wire new_Jinkela_wire_11216;
    wire new_Jinkela_wire_8217;
    wire new_Jinkela_wire_16808;
    wire new_Jinkela_wire_17575;
    wire new_Jinkela_wire_15530;
    wire new_Jinkela_wire_20488;
    wire new_Jinkela_wire_11347;
    wire _0024_;
    wire new_Jinkela_wire_5773;
    wire new_Jinkela_wire_1984;
    wire new_Jinkela_wire_3637;
    wire _1032_;
    wire _1455_;
    wire new_Jinkela_wire_12587;
    wire new_Jinkela_wire_21071;
    wire new_Jinkela_wire_20518;
    wire _0196_;
    wire new_Jinkela_wire_3426;
    wire new_Jinkela_wire_20998;
    wire new_Jinkela_wire_1294;
    wire _1223_;
    wire new_Jinkela_wire_7879;
    wire new_Jinkela_wire_19607;
    wire new_Jinkela_wire_7275;
    wire _0777_;
    wire new_Jinkela_wire_15670;
    wire new_Jinkela_wire_10305;
    wire new_Jinkela_wire_9080;
    wire new_Jinkela_wire_11684;
    wire _1394_;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_3297;
    wire new_Jinkela_wire_13543;
    wire new_Jinkela_wire_11393;
    wire new_Jinkela_wire_11598;
    wire new_Jinkela_wire_6067;
    wire new_Jinkela_wire_6463;
    wire new_Jinkela_wire_16957;
    wire new_Jinkela_wire_2779;
    wire new_Jinkela_wire_9999;
    wire new_Jinkela_wire_6002;
    wire new_Jinkela_wire_8844;
    wire new_Jinkela_wire_8181;
    wire new_Jinkela_wire_17496;
    wire new_Jinkela_wire_5716;
    wire new_Jinkela_wire_8876;
    wire new_Jinkela_wire_13445;
    wire new_Jinkela_wire_8223;
    wire new_Jinkela_wire_15444;
    wire new_Jinkela_wire_9572;
    wire new_Jinkela_wire_17640;
    wire new_Jinkela_wire_10327;
    wire _0597_;
    wire new_Jinkela_wire_5544;
    wire new_Jinkela_wire_4588;
    wire _0919_;
    wire new_Jinkela_wire_12131;
    wire new_Jinkela_wire_19074;
    wire new_Jinkela_wire_19480;
    wire new_Jinkela_wire_1745;
    wire new_Jinkela_wire_12291;
    wire new_Jinkela_wire_7229;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_15367;
    wire new_Jinkela_wire_6455;
    wire new_Jinkela_wire_1829;
    wire new_Jinkela_wire_17885;
    wire new_Jinkela_wire_9818;
    wire new_Jinkela_wire_14760;
    wire new_Jinkela_wire_15614;
    wire new_Jinkela_wire_16099;
    wire new_Jinkela_wire_6472;
    wire new_Jinkela_wire_11173;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_11936;
    wire new_Jinkela_wire_10422;
    wire new_Jinkela_wire_20978;
    wire new_Jinkela_wire_15863;
    wire _0134_;
    wire new_Jinkela_wire_20569;
    wire new_Jinkela_wire_9420;
    wire new_Jinkela_wire_12802;
    wire new_Jinkela_wire_12128;
    wire new_Jinkela_wire_2159;
    wire _0764_;
    wire new_Jinkela_wire_1073;
    wire new_Jinkela_wire_18509;
    wire new_Jinkela_wire_19749;
    wire new_Jinkela_wire_2158;
    wire new_Jinkela_wire_2763;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_20238;
    wire new_Jinkela_wire_14824;
    wire new_Jinkela_wire_20287;
    wire new_Jinkela_wire_17729;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_1935;
    wire new_Jinkela_wire_4165;
    wire new_Jinkela_wire_11538;
    wire new_Jinkela_wire_17988;
    wire new_Jinkela_wire_12196;
    wire new_Jinkela_wire_3998;
    wire new_Jinkela_wire_19065;
    wire new_Jinkela_wire_13818;
    wire new_Jinkela_wire_2725;
    wire new_Jinkela_wire_4614;
    wire new_Jinkela_wire_16013;
    wire new_Jinkela_wire_3983;
    wire new_Jinkela_wire_7052;
    wire new_Jinkela_wire_2292;
    wire new_Jinkela_wire_4739;
    wire new_Jinkela_wire_17834;
    wire new_Jinkela_wire_19551;
    wire new_Jinkela_wire_19738;
    wire new_Jinkela_wire_9029;
    wire new_Jinkela_wire_14955;
    wire new_Jinkela_wire_20256;
    wire new_Jinkela_wire_16058;
    wire new_Jinkela_wire_10621;
    wire new_Jinkela_wire_11098;
    wire new_Jinkela_wire_3797;
    wire new_Jinkela_wire_9170;
    wire _1555_;
    wire new_Jinkela_wire_19589;
    wire new_Jinkela_wire_17242;
    wire new_Jinkela_wire_13046;
    wire new_Jinkela_wire_17398;
    wire new_Jinkela_wire_11868;
    wire new_Jinkela_wire_16840;
    wire new_Jinkela_wire_15999;
    wire new_Jinkela_wire_2576;
    wire new_Jinkela_wire_17304;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_5796;
    wire new_Jinkela_wire_12576;
    wire new_Jinkela_wire_18986;
    wire new_Jinkela_wire_9342;
    wire _1491_;
    wire new_Jinkela_wire_11520;
    wire new_Jinkela_wire_3663;
    wire new_Jinkela_wire_16135;
    wire new_Jinkela_wire_4875;
    wire new_Jinkela_wire_3571;
    wire new_Jinkela_wire_18608;
    wire new_Jinkela_wire_3876;
    wire new_Jinkela_wire_8938;
    wire new_Jinkela_wire_9388;
    wire new_Jinkela_wire_3831;
    wire new_Jinkela_wire_8189;
    wire new_Jinkela_wire_18794;
    wire new_Jinkela_wire_5418;
    wire new_Jinkela_wire_13304;
    wire new_Jinkela_wire_13112;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_21002;
    wire new_Jinkela_wire_5056;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_6892;
    wire new_Jinkela_wire_18643;
    wire new_Jinkela_wire_9001;
    wire new_Jinkela_wire_8993;
    wire new_Jinkela_wire_4788;
    wire new_Jinkela_wire_8703;
    wire _1794_;
    wire _1262_;
    wire new_Jinkela_wire_4829;
    wire new_Jinkela_wire_12090;
    wire new_Jinkela_wire_4382;
    wire _0257_;
    wire new_Jinkela_wire_6167;
    wire new_Jinkela_wire_2372;
    wire new_Jinkela_wire_6605;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_2145;
    wire new_Jinkela_wire_6583;
    wire new_Jinkela_wire_14739;
    wire new_Jinkela_wire_3990;
    wire new_Jinkela_wire_19473;
    wire new_Jinkela_wire_3845;
    wire new_Jinkela_wire_12368;
    wire new_Jinkela_wire_9717;
    wire new_Jinkela_wire_14724;
    wire _0615_;
    wire new_Jinkela_wire_9880;
    wire new_Jinkela_wire_20038;
    wire new_Jinkela_wire_3291;
    wire new_Jinkela_wire_7164;
    wire new_Jinkela_wire_20366;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_5768;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_17278;
    wire new_Jinkela_wire_18326;
    wire _0872_;
    wire new_Jinkela_wire_18837;
    wire new_Jinkela_wire_9335;
    wire new_Jinkela_wire_19205;
    wire new_Jinkela_wire_8471;
    wire new_Jinkela_wire_18498;
    wire _1630_;
    wire new_Jinkela_wire_11718;
    wire new_Jinkela_wire_17920;
    wire new_Jinkela_wire_6308;
    wire new_Jinkela_wire_16664;
    wire new_Jinkela_wire_3249;
    wire new_Jinkela_wire_13030;
    wire new_Jinkela_wire_6879;
    wire new_Jinkela_wire_10884;
    wire new_Jinkela_wire_10166;
    wire new_Jinkela_wire_18966;
    wire new_Jinkela_wire_6796;
    wire new_Jinkela_wire_17791;
    wire new_Jinkela_wire_17429;
    wire _0124_;
    wire new_Jinkela_wire_5335;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_10232;
    wire new_Jinkela_wire_7856;
    wire new_Jinkela_wire_14669;
    wire new_Jinkela_wire_13582;
    wire new_Jinkela_wire_11903;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_18441;
    wire new_Jinkela_wire_16855;
    wire new_Jinkela_wire_12061;
    wire new_Jinkela_wire_17065;
    wire new_Jinkela_wire_20661;
    wire new_Jinkela_wire_7140;
    wire _0824_;
    wire new_Jinkela_wire_4496;
    wire new_Jinkela_wire_5676;
    wire new_Jinkela_wire_4550;
    wire new_Jinkela_wire_2360;
    wire new_Jinkela_wire_17722;
    wire new_Jinkela_wire_3733;
    wire new_Jinkela_wire_6941;
    wire new_Jinkela_wire_5313;
    wire _0423_;
    wire new_Jinkela_wire_2086;
    wire _0844_;
    wire new_Jinkela_wire_21212;
    wire new_Jinkela_wire_2280;
    wire new_Jinkela_wire_7649;
    wire _0957_;
    wire new_Jinkela_wire_10194;
    wire new_Jinkela_wire_16283;
    wire new_Jinkela_wire_4650;
    wire new_Jinkela_wire_14559;
    wire new_Jinkela_wire_10777;
    wire new_Jinkela_wire_12275;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_7176;
    wire new_Jinkela_wire_11327;
    wire new_Jinkela_wire_5362;
    wire new_Jinkela_wire_17221;
    wire new_Jinkela_wire_9859;
    wire new_Jinkela_wire_18599;
    wire new_Jinkela_wire_10552;
    wire new_Jinkela_wire_16014;
    wire new_Jinkela_wire_18256;
    wire new_Jinkela_wire_17599;
    wire new_Jinkela_wire_19490;
    wire _0093_;
    wire _0494_;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_5103;
    wire new_Jinkela_wire_3161;
    wire new_Jinkela_wire_7567;
    wire new_Jinkela_wire_18721;
    wire new_Jinkela_wire_21215;
    wire new_Jinkela_wire_4900;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_2357;
    wire new_Jinkela_wire_18069;
    wire new_Jinkela_wire_20267;
    wire new_Jinkela_wire_7017;
    wire new_Jinkela_wire_5753;
    wire new_Jinkela_wire_7701;
    wire new_Jinkela_wire_8074;
    wire new_Jinkela_wire_17397;
    wire new_Jinkela_wire_2012;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_7128;
    wire new_Jinkela_wire_13052;
    wire new_Jinkela_wire_4825;
    wire new_Jinkela_wire_17096;
    wire new_Jinkela_wire_12193;
    wire new_Jinkela_wire_20486;
    wire new_Jinkela_wire_18821;
    wire _1653_;
    wire new_Jinkela_wire_18656;
    wire new_Jinkela_wire_4978;
    wire new_Jinkela_wire_16668;
    wire new_Jinkela_wire_16607;
    wire new_Jinkela_wire_12410;
    wire new_Jinkela_wire_9465;
    wire new_Jinkela_wire_20428;
    wire new_Jinkela_wire_4443;
    wire new_Jinkela_wire_16141;
    wire new_Jinkela_wire_12441;
    wire new_Jinkela_wire_5776;
    wire new_Jinkela_wire_16692;
    wire new_Jinkela_wire_4961;
    wire new_Jinkela_wire_18694;
    wire new_Jinkela_wire_4327;
    wire new_Jinkela_wire_5592;
    wire new_Jinkela_wire_19317;
    wire _1048_;
    wire new_Jinkela_wire_13200;
    wire new_Jinkela_wire_17945;
    wire new_Jinkela_wire_12559;
    wire new_Jinkela_wire_7092;
    wire _0211_;
    wire new_Jinkela_wire_21227;
    wire new_Jinkela_wire_11283;
    wire new_Jinkela_wire_3598;
    wire new_Jinkela_wire_15334;
    wire new_Jinkela_wire_4899;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_15159;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_11101;
    wire new_Jinkela_wire_18265;
    wire new_Jinkela_wire_19335;
    wire new_Jinkela_wire_15080;
    wire new_Jinkela_wire_3758;
    wire new_Jinkela_wire_19215;
    wire new_Jinkela_wire_19186;
    wire new_Jinkela_wire_4460;
    wire new_Jinkela_wire_18824;
    wire new_Jinkela_wire_6632;
    wire new_Jinkela_wire_12510;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_7455;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_14755;
    wire new_Jinkela_wire_16839;
    wire new_Jinkela_wire_16282;
    wire new_Jinkela_wire_19468;
    wire new_Jinkela_wire_2849;
    wire _0080_;
    wire new_Jinkela_wire_14837;
    wire new_Jinkela_wire_20583;
    wire new_Jinkela_wire_5048;
    wire new_Jinkela_wire_5298;
    wire new_Jinkela_wire_12890;
    wire _0175_;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_20751;
    wire new_Jinkela_wire_4134;
    wire new_Jinkela_wire_16960;
    wire new_Jinkela_wire_13496;
    wire new_Jinkela_wire_20302;
    wire new_Jinkela_wire_10279;
    wire new_Jinkela_wire_20831;
    wire new_Jinkela_wire_4834;
    wire new_Jinkela_wire_14999;
    wire new_Jinkela_wire_3379;
    wire new_Jinkela_wire_5541;
    wire new_Jinkela_wire_21013;
    wire new_Jinkela_wire_17763;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_12219;
    wire new_Jinkela_wire_8406;
    wire new_Jinkela_wire_7351;
    wire new_Jinkela_wire_18705;
    wire new_Jinkela_wire_7907;
    wire new_Jinkela_wire_17453;
    wire new_Jinkela_wire_9112;
    wire new_Jinkela_wire_7413;
    wire new_Jinkela_wire_19373;
    wire new_Jinkela_wire_5833;
    wire new_Jinkela_wire_10103;
    wire new_Jinkela_wire_16594;
    wire new_Jinkela_wire_13736;
    wire new_Jinkela_wire_5181;
    wire new_Jinkela_wire_17855;
    wire new_Jinkela_wire_3386;
    wire new_Jinkela_wire_8086;
    wire new_Jinkela_wire_2813;
    wire new_Jinkela_wire_19478;
    wire new_Jinkela_wire_17143;
    wire new_Jinkela_wire_9158;
    wire new_Jinkela_wire_5817;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_18216;
    wire new_Jinkela_wire_3729;
    wire new_Jinkela_wire_5357;
    wire new_Jinkela_wire_18403;
    wire new_Jinkela_wire_15172;
    wire new_Jinkela_wire_8710;
    wire new_Jinkela_wire_8356;
    wire _1788_;
    wire new_Jinkela_wire_20104;
    wire new_Jinkela_wire_4402;
    wire new_Jinkela_wire_14304;
    wire new_Jinkela_wire_19431;
    wire new_Jinkela_wire_15466;
    wire new_Jinkela_wire_19213;
    wire new_Jinkela_wire_8001;
    wire new_Jinkela_wire_20698;
    wire new_Jinkela_wire_9966;
    wire new_Jinkela_wire_3120;
    wire new_Jinkela_wire_13478;
    wire new_Jinkela_wire_4827;
    wire new_Jinkela_wire_7254;
    wire new_Jinkela_wire_21236;
    wire new_Jinkela_wire_2554;
    wire new_Jinkela_wire_11767;
    wire new_Jinkela_wire_3453;
    wire new_Jinkela_wire_18174;
    wire new_Jinkela_wire_8193;
    wire new_Jinkela_wire_4594;
    wire new_Jinkela_wire_4448;
    wire new_Jinkela_wire_2399;
    wire new_Jinkela_wire_20958;
    wire new_Jinkela_wire_2153;
    wire new_Jinkela_wire_7577;
    wire new_Jinkela_wire_17261;
    wire new_Jinkela_wire_12016;
    wire new_Jinkela_wire_3795;
    wire new_Jinkela_wire_6741;
    wire new_Jinkela_wire_5498;
    wire new_Jinkela_wire_11213;
    wire new_Jinkela_wire_16110;
    wire new_Jinkela_wire_9919;
    wire new_Jinkela_wire_20475;
    wire new_Jinkela_wire_3871;
    wire new_Jinkela_wire_8190;
    wire new_Jinkela_wire_18359;
    wire new_Jinkela_wire_19132;
    wire new_Jinkela_wire_20735;
    wire new_Jinkela_wire_19056;
    wire new_Jinkela_wire_1689;
    wire _1028_;
    wire new_Jinkela_wire_13641;
    wire new_Jinkela_wire_20895;
    wire new_Jinkela_wire_6110;
    wire new_Jinkela_wire_20482;
    wire new_Jinkela_wire_19843;
    wire new_Jinkela_wire_13139;
    wire new_Jinkela_wire_6592;
    wire new_Jinkela_wire_6334;
    wire new_Jinkela_wire_9856;
    wire new_Jinkela_wire_20137;
    wire new_Jinkela_wire_3804;
    wire new_Jinkela_wire_16111;
    wire new_Jinkela_wire_18490;
    wire new_Jinkela_wire_5807;
    wire new_Jinkela_wire_3028;
    wire new_Jinkela_wire_17972;
    wire new_Jinkela_wire_21155;
    wire new_Jinkela_wire_14715;
    wire new_Jinkela_wire_2864;
    wire _1784_;
    wire new_Jinkela_wire_1899;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_7763;
    wire new_Jinkela_wire_10146;
    wire new_Jinkela_wire_8943;
    wire new_Jinkela_wire_8403;
    wire new_Jinkela_wire_19110;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_10290;
    wire new_Jinkela_wire_11425;
    wire new_Jinkela_wire_3918;
    wire _0886_;
    wire new_Jinkela_wire_11467;
    wire new_Jinkela_wire_8649;
    wire new_Jinkela_wire_8010;
    wire new_Jinkela_wire_13819;
    wire new_Jinkela_wire_13423;
    wire new_Jinkela_wire_9848;
    wire new_Jinkela_wire_6567;
    wire _0460_;
    wire new_Jinkela_wire_16579;
    wire new_Jinkela_wire_18804;
    wire new_Jinkela_wire_10635;
    wire new_Jinkela_wire_8970;
    wire new_Jinkela_wire_14932;
    wire new_Jinkela_wire_10601;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_7006;
    wire new_Jinkela_wire_20164;
    wire new_Jinkela_wire_895;
    wire new_Jinkela_wire_6926;
    wire new_Jinkela_wire_6918;
    wire new_Jinkela_wire_16877;
    wire new_Jinkela_wire_8557;
    wire new_Jinkela_wire_3446;
    wire new_Jinkela_wire_4576;
    wire new_Jinkela_wire_9003;
    wire new_Jinkela_wire_18072;
    wire new_Jinkela_wire_8843;
    wire new_Jinkela_wire_4914;
    wire new_Jinkela_wire_5373;
    wire _1772_;
    wire _0912_;
    wire new_Jinkela_wire_8353;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_4700;
    wire _0078_;
    wire new_Jinkela_wire_4818;
    wire new_Jinkela_wire_13662;
    wire new_Jinkela_wire_20527;
    wire new_Jinkela_wire_7295;
    wire _1037_;
    wire new_Jinkela_wire_14285;
    wire new_Jinkela_wire_12321;
    wire new_Jinkela_wire_17482;
    wire new_Jinkela_wire_15832;
    wire new_Jinkela_wire_2238;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_6982;
    wire new_Jinkela_wire_9489;
    wire new_Jinkela_wire_5360;
    wire new_Jinkela_wire_11132;
    wire new_Jinkela_wire_19514;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_15712;
    wire new_Jinkela_wire_15467;
    wire new_Jinkela_wire_9177;
    wire new_Jinkela_wire_4525;
    wire new_Jinkela_wire_3224;
    wire new_Jinkela_wire_19487;
    wire new_Jinkela_wire_2135;
    wire new_Jinkela_wire_16383;
    wire new_Jinkela_wire_11262;
    wire new_Jinkela_wire_13626;
    wire new_Jinkela_wire_4019;
    wire new_Jinkela_wire_13661;
    wire new_Jinkela_wire_7719;
    wire _1785_;
    wire new_Jinkela_wire_19536;
    wire new_Jinkela_wire_17784;
    wire new_Jinkela_wire_19146;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_8295;
    wire new_Jinkela_wire_16068;
    wire new_Jinkela_wire_16312;
    wire new_Jinkela_wire_17687;
    wire new_Jinkela_wire_10617;
    wire new_Jinkela_wire_3861;
    wire new_Jinkela_wire_14478;
    wire new_Jinkela_wire_14329;
    wire new_Jinkela_wire_8759;
    wire new_Jinkela_wire_9891;
    wire new_Jinkela_wire_4190;
    wire new_Jinkela_wire_2691;
    wire new_Jinkela_wire_4294;
    wire new_Jinkela_wire_9506;
    wire new_Jinkela_wire_12074;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_11894;
    wire new_Jinkela_wire_10022;
    wire new_Jinkela_wire_19058;
    wire new_Jinkela_wire_8632;
    wire new_Jinkela_wire_19154;
    wire new_Jinkela_wire_6888;
    wire _0415_;
    wire _1136_;
    wire new_Jinkela_wire_7669;
    wire new_Jinkela_wire_19253;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_10091;
    wire new_Jinkela_wire_9216;
    wire new_Jinkela_wire_10540;
    wire new_Jinkela_wire_3179;
    wire new_Jinkela_wire_8034;
    wire new_Jinkela_wire_14850;
    wire new_Jinkela_wire_17000;
    wire new_Jinkela_wire_19530;
    wire _1055_;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_6162;
    wire new_Jinkela_wire_3938;
    wire new_Jinkela_wire_12626;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_20659;
    wire new_Jinkela_wire_15484;
    wire new_Jinkela_wire_3306;
    wire new_Jinkela_wire_16032;
    wire new_Jinkela_wire_20190;
    wire new_Jinkela_wire_6306;
    wire new_Jinkela_wire_10965;
    wire new_Jinkela_wire_19102;
    wire new_Jinkela_wire_13447;
    wire new_Jinkela_wire_1178;
    wire new_Jinkela_wire_20625;
    wire new_Jinkela_wire_12847;
    wire new_Jinkela_wire_4883;
    wire _0305_;
    wire new_Jinkela_wire_6165;
    wire new_Jinkela_wire_18453;
    wire new_Jinkela_wire_3309;
    wire new_Jinkela_wire_4186;
    wire new_Jinkela_wire_15324;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_18493;
    wire new_Jinkela_wire_4980;
    wire new_Jinkela_wire_11083;
    wire new_Jinkela_wire_2303;
    wire new_Jinkela_wire_12659;
    wire new_Jinkela_wire_9188;
    wire new_Jinkela_wire_12284;
    wire new_Jinkela_wire_13050;
    wire new_Jinkela_wire_18229;
    wire new_Jinkela_wire_13041;
    wire new_Jinkela_wire_9559;
    wire new_Jinkela_wire_16710;
    wire _1258_;
    wire _0616_;
    wire new_Jinkela_wire_13576;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_10835;
    wire new_Jinkela_wire_6376;
    wire new_Jinkela_wire_18083;
    wire new_Jinkela_wire_20322;
    wire new_Jinkela_wire_18249;
    wire new_Jinkela_wire_18448;
    wire new_Jinkela_wire_17814;
    wire new_Jinkela_wire_2401;
    wire _0097_;
    wire new_Jinkela_wire_5111;
    wire new_Jinkela_wire_12155;
    wire new_Jinkela_wire_11473;
    wire _0391_;
    wire new_Jinkela_wire_14270;
    wire _0837_;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_10079;
    wire new_Jinkela_wire_6028;
    wire new_Jinkela_wire_19899;
    wire new_Jinkela_wire_17308;
    wire new_Jinkela_wire_7488;
    wire new_Jinkela_wire_21140;
    wire new_Jinkela_wire_5129;
    wire new_Jinkela_wire_3072;
    wire new_Jinkela_wire_12350;
    wire new_Jinkela_wire_2714;
    wire new_Jinkela_wire_16819;
    wire new_Jinkela_wire_7915;
    wire new_Jinkela_wire_12520;
    wire new_Jinkela_wire_6340;
    wire new_Jinkela_wire_20341;
    wire new_Jinkela_wire_14538;
    wire new_Jinkela_wire_7074;
    wire new_Jinkela_wire_14977;
    wire new_Jinkela_wire_5461;
    wire new_Jinkela_wire_12991;
    wire new_Jinkela_wire_11858;
    wire new_Jinkela_wire_9037;
    wire new_Jinkela_wire_9223;
    wire new_Jinkela_wire_8897;
    wire new_Jinkela_wire_20871;
    wire new_Jinkela_wire_9334;
    wire new_Jinkela_wire_15825;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_4747;
    wire new_Jinkela_wire_6422;
    wire new_Jinkela_wire_16928;
    wire new_Jinkela_wire_4447;
    wire new_Jinkela_wire_8988;
    wire new_Jinkela_wire_18999;
    wire new_Jinkela_wire_7184;
    wire new_Jinkela_wire_18067;
    wire new_Jinkela_wire_16586;
    wire new_Jinkela_wire_10964;
    wire _0822_;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_2210;
    wire new_Jinkela_wire_15543;
    wire new_Jinkela_wire_8075;
    wire new_Jinkela_wire_19936;
    wire new_Jinkela_wire_7634;
    wire _0440_;
    wire new_Jinkela_wire_4449;
    wire new_Jinkela_wire_5235;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_13867;
    wire _1351_;
    wire _1013_;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_15313;
    wire new_Jinkela_wire_14412;
    wire new_Jinkela_wire_19277;
    wire new_Jinkela_wire_4398;
    wire new_Jinkela_wire_15293;
    wire _0630_;
    wire new_Jinkela_wire_3071;
    wire new_Jinkela_wire_5859;
    wire new_Jinkela_wire_11616;
    wire new_Jinkela_wire_15963;
    wire new_Jinkela_wire_2856;
    wire new_Jinkela_wire_9670;
    wire new_Jinkela_wire_11085;
    wire new_Jinkela_wire_10547;
    wire new_Jinkela_wire_17863;
    wire new_Jinkela_wire_20297;
    wire new_Jinkela_wire_3105;
    wire new_Jinkela_wire_6989;
    wire new_Jinkela_wire_19072;
    wire new_Jinkela_wire_10223;
    wire new_Jinkela_wire_10899;
    wire new_Jinkela_wire_9697;
    wire new_Jinkela_wire_2132;
    wire new_Jinkela_wire_11940;
    wire new_Jinkela_wire_17468;
    wire new_Jinkela_wire_11381;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_13907;
    wire new_Jinkela_wire_6047;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_13673;
    wire new_Jinkela_wire_18722;
    wire new_Jinkela_wire_3927;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_8727;
    wire new_Jinkela_wire_2426;
    wire new_Jinkela_wire_9050;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_19185;
    wire new_Jinkela_wire_4083;
    wire new_Jinkela_wire_7244;
    wire new_Jinkela_wire_4933;
    wire new_Jinkela_wire_9470;
    wire _1012_;
    wire new_Jinkela_wire_14451;
    wire new_Jinkela_wire_16829;
    wire new_Jinkela_wire_7227;
    wire new_Jinkela_wire_4951;
    wire new_Jinkela_wire_1166;
    wire new_Jinkela_wire_2353;
    wire new_Jinkela_wire_14068;
    wire new_Jinkela_wire_15942;
    wire new_Jinkela_wire_15699;
    wire new_Jinkela_wire_7781;
    wire new_Jinkela_wire_10297;
    wire new_Jinkela_wire_11608;
    wire new_Jinkela_wire_9879;
    wire new_Jinkela_wire_15581;
    wire new_Jinkela_wire_15084;
    wire new_Jinkela_wire_16968;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_15986;
    wire new_Jinkela_wire_11827;
    wire new_Jinkela_wire_6300;
    wire new_Jinkela_wire_5886;
    wire new_Jinkela_wire_14142;
    wire new_Jinkela_wire_8564;
    wire new_Jinkela_wire_12383;
    wire new_Jinkela_wire_10966;
    wire new_Jinkela_wire_9075;
    wire new_Jinkela_wire_16830;
    wire new_Jinkela_wire_6068;
    wire new_Jinkela_wire_16932;
    wire new_Jinkela_wire_11496;
    wire new_Jinkela_wire_9583;
    wire new_Jinkela_wire_20578;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_2184;
    wire new_Jinkela_wire_19518;
    wire new_Jinkela_wire_18056;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_20705;
    wire new_Jinkela_wire_19904;
    wire new_Jinkela_wire_12280;
    wire new_Jinkela_wire_6794;
    wire new_Jinkela_wire_13915;
    wire new_Jinkela_wire_21092;
    wire new_Jinkela_wire_3450;
    wire new_Jinkela_wire_7936;
    wire new_Jinkela_wire_2701;
    wire new_Jinkela_wire_6099;
    wire new_Jinkela_wire_19546;
    wire new_Jinkela_wire_10140;
    wire _1409_;
    wire new_Jinkela_wire_12719;
    wire new_Jinkela_wire_17107;
    wire new_Jinkela_wire_3460;
    wire new_Jinkela_wire_2742;
    wire new_Jinkela_wire_15448;
    wire new_net_3964;
    wire new_Jinkela_wire_16850;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_13719;
    wire new_Jinkela_wire_20764;
    wire new_Jinkela_wire_21035;
    wire new_Jinkela_wire_16741;
    wire new_Jinkela_wire_15795;
    wire new_Jinkela_wire_2853;
    wire new_Jinkela_wire_3838;
    wire new_Jinkela_wire_4852;
    wire new_Jinkela_wire_5800;
    wire new_Jinkela_wire_10427;
    wire new_Jinkela_wire_16267;
    wire new_Jinkela_wire_18901;
    wire new_Jinkela_wire_6449;
    wire new_Jinkela_wire_4260;
    wire new_Jinkela_wire_16425;
    wire new_Jinkela_wire_7297;
    wire new_Jinkela_wire_20141;
    wire new_Jinkela_wire_11249;
    wire new_Jinkela_wire_2125;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_7330;
    wire new_Jinkela_wire_16223;
    wire new_Jinkela_wire_8833;
    wire new_Jinkela_wire_20676;
    wire new_Jinkela_wire_19541;
    wire new_Jinkela_wire_19614;
    wire new_Jinkela_wire_4308;
    wire _1597_;
    wire new_Jinkela_wire_2592;
    wire new_Jinkela_wire_4217;
    wire new_Jinkela_wire_13136;
    wire new_Jinkela_wire_5930;
    wire new_Jinkela_wire_11960;
    wire new_Jinkela_wire_20931;
    wire new_Jinkela_wire_2548;
    wire new_Jinkela_wire_8478;
    wire new_Jinkela_wire_6682;
    wire new_Jinkela_wire_12690;
    wire new_Jinkela_wire_7291;
    wire new_Jinkela_wire_20181;
    wire new_Jinkela_wire_20449;
    wire new_Jinkela_wire_11547;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_10761;
    wire new_Jinkela_wire_12418;
    wire new_Jinkela_wire_5746;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_13398;
    wire new_Jinkela_wire_16435;
    wire new_Jinkela_wire_412;
    wire _1774_;
    wire new_Jinkela_wire_8575;
    wire new_Jinkela_wire_3255;
    wire new_Jinkela_wire_5095;
    wire new_Jinkela_wire_19597;
    wire new_Jinkela_wire_16464;
    wire new_Jinkela_wire_11235;
    wire new_Jinkela_wire_6374;
    wire new_Jinkela_wire_15012;
    wire new_Jinkela_wire_6072;
    wire new_Jinkela_wire_20052;
    wire new_Jinkela_wire_5325;
    wire new_Jinkela_wire_15447;
    wire new_Jinkela_wire_5891;
    wire new_Jinkela_wire_13885;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_15183;
    wire new_Jinkela_wire_1957;
    wire new_Jinkela_wire_5883;
    wire new_Jinkela_wire_6963;
    wire new_Jinkela_wire_16901;
    wire new_Jinkela_wire_21032;
    wire new_Jinkela_wire_20879;
    wire new_Jinkela_wire_12007;
    wire new_Jinkela_wire_2602;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_6278;
    wire new_Jinkela_wire_19729;
    wire new_Jinkela_wire_16818;
    wire new_Jinkela_wire_19641;
    wire new_Jinkela_wire_3680;
    wire new_Jinkela_wire_9138;
    wire new_Jinkela_wire_10915;
    wire new_Jinkela_wire_2644;
    wire new_Jinkela_wire_8698;
    wire new_Jinkela_wire_12171;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_21038;
    wire new_Jinkela_wire_9482;
    wire new_Jinkela_wire_3131;
    wire new_Jinkela_wire_4849;
    wire _1461_;
    wire _1165_;
    wire new_Jinkela_wire_3981;
    wire _1329_;
    wire new_Jinkela_wire_17539;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_2367;
    wire new_Jinkela_wire_8264;
    wire new_Jinkela_wire_5501;
    wire new_Jinkela_wire_9386;
    wire new_Jinkela_wire_18037;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_20289;
    wire new_Jinkela_wire_12668;
    wire new_Jinkela_wire_10689;
    wire new_Jinkela_wire_10534;
    wire new_Jinkela_wire_15852;
    wire new_Jinkela_wire_13315;
    wire new_Jinkela_wire_3818;
    wire new_Jinkela_wire_19562;
    wire new_Jinkela_wire_5146;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_18361;
    wire new_Jinkela_wire_9164;
    wire new_Jinkela_wire_13741;
    wire new_Jinkela_wire_16591;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_20854;
    wire new_Jinkela_wire_16806;
    wire new_Jinkela_wire_7258;
    wire new_Jinkela_wire_12151;
    wire _0050_;
    wire new_Jinkela_wire_15424;
    wire _1088_;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_5331;
    wire new_Jinkela_wire_16747;
    wire new_Jinkela_wire_8724;
    wire new_Jinkela_wire_14244;
    wire new_Jinkela_wire_10875;
    wire new_Jinkela_wire_12524;
    wire new_Jinkela_wire_7011;
    wire new_Jinkela_wire_5960;
    wire new_Jinkela_wire_5420;
    wire new_Jinkela_wire_11774;
    wire new_Jinkela_wire_7151;
    wire new_Jinkela_wire_18693;
    wire new_Jinkela_wire_16372;
    wire new_Jinkela_wire_9836;
    wire new_Jinkela_wire_3549;
    wire new_Jinkela_wire_8825;
    wire new_Jinkela_wire_21325;
    wire new_Jinkela_wire_14332;
    wire new_Jinkela_wire_17259;
    wire new_Jinkela_wire_15130;
    wire new_Jinkela_wire_9762;
    wire new_Jinkela_wire_3274;
    wire new_Jinkela_wire_7580;
    wire new_Jinkela_wire_21200;
    wire new_Jinkela_wire_15420;
    wire new_Jinkela_wire_20210;
    wire new_Jinkela_wire_12947;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_13356;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_12422;
    wire new_Jinkela_wire_2754;
    wire new_Jinkela_wire_6080;
    wire new_Jinkela_wire_14090;
    wire new_Jinkela_wire_14616;
    wire new_Jinkela_wire_19031;
    wire new_Jinkela_wire_1797;
    wire new_Jinkela_wire_14615;
    wire new_Jinkela_wire_7493;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_7316;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_11882;
    wire new_Jinkela_wire_20542;
    wire new_Jinkela_wire_18009;
    wire new_Jinkela_wire_12211;
    wire new_Jinkela_wire_9166;
    wire new_Jinkela_wire_21163;
    wire new_Jinkela_wire_12797;
    wire new_Jinkela_wire_3213;
    wire new_Jinkela_wire_4844;
    wire new_Jinkela_wire_4235;
    wire new_Jinkela_wire_17244;
    wire new_Jinkela_wire_20983;
    wire new_Jinkela_wire_2155;
    wire new_Jinkela_wire_16606;
    wire _0242_;
    wire new_Jinkela_wire_5147;
    wire new_Jinkela_wire_16631;
    wire _1010_;
    wire new_Jinkela_wire_18352;
    wire new_Jinkela_wire_12399;
    wire new_Jinkela_wire_14845;
    wire new_Jinkela_wire_10151;
    wire new_Jinkela_wire_9657;
    wire _1541_;
    wire _0036_;
    wire new_Jinkela_wire_18876;
    wire new_Jinkela_wire_20027;
    wire _1692_;
    wire _0853_;
    wire new_Jinkela_wire_15511;
    wire new_Jinkela_wire_5767;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_8885;
    wire new_Jinkela_wire_21040;
    wire new_Jinkela_wire_4146;
    wire new_Jinkela_wire_10479;
    wire new_Jinkela_wire_16530;
    wire _1008_;
    wire new_Jinkela_wire_5108;
    wire new_Jinkela_wire_18260;
    wire new_Jinkela_wire_20034;
    wire new_Jinkela_wire_15067;
    wire new_Jinkela_wire_5819;
    wire new_Jinkela_wire_21295;
    wire new_Jinkela_wire_12210;
    wire new_Jinkela_wire_6223;
    wire new_Jinkela_wire_9566;
    wire new_Jinkela_wire_5774;
    wire new_Jinkela_wire_10754;
    wire new_Jinkela_wire_20573;
    wire new_Jinkela_wire_9231;
    wire _0298_;
    wire new_Jinkela_wire_11197;
    wire new_Jinkela_wire_2971;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_15633;
    wire new_Jinkela_wire_6513;
    wire new_Jinkela_wire_15362;
    wire new_Jinkela_wire_121;
    wire new_Jinkela_wire_4593;
    wire new_Jinkela_wire_11949;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_12553;
    wire new_Jinkela_wire_9209;
    wire new_Jinkela_wire_3128;
    wire new_Jinkela_wire_11243;
    wire new_Jinkela_wire_5793;
    wire new_Jinkela_wire_8527;
    wire new_Jinkela_wire_6040;
    wire new_Jinkela_wire_3096;
    wire new_Jinkela_wire_5087;
    wire new_Jinkela_wire_16025;
    wire new_Jinkela_wire_12850;
    wire new_Jinkela_wire_12953;
    wire new_Jinkela_wire_8046;
    wire new_Jinkela_wire_12023;
    wire new_Jinkela_wire_20749;
    wire new_Jinkela_wire_17284;
    wire new_Jinkela_wire_2918;
    wire new_Jinkela_wire_4604;
    wire _0519_;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_18861;
    wire new_Jinkela_wire_14102;
    wire new_Jinkela_wire_5953;
    wire _0533_;
    wire new_Jinkela_wire_11591;
    wire _0011_;
    wire new_Jinkela_wire_14957;
    wire new_Jinkela_wire_1802;
    wire new_Jinkela_wire_12066;
    wire _0094_;
    wire new_Jinkela_wire_20317;
    wire _0057_;
    wire _0964_;
    wire new_Jinkela_wire_11987;
    wire _0665_;
    wire new_Jinkela_wire_16160;
    wire new_Jinkela_wire_4263;
    wire new_Jinkela_wire_3743;
    wire new_Jinkela_wire_18603;
    wire new_Jinkela_wire_12201;
    wire new_Jinkela_wire_18313;
    wire new_Jinkela_wire_6889;
    wire new_Jinkela_wire_5971;
    wire new_Jinkela_wire_8969;
    wire new_Jinkela_wire_11445;
    wire new_Jinkela_wire_3545;
    wire new_Jinkela_wire_10937;
    wire new_Jinkela_wire_4039;
    wire new_Jinkela_wire_12781;
    wire new_Jinkela_wire_11658;
    wire new_Jinkela_wire_13798;
    wire new_Jinkela_wire_4801;
    wire new_Jinkela_wire_20208;
    wire new_Jinkela_wire_11785;
    wire new_Jinkela_wire_9060;
    wire new_Jinkela_wire_19649;
    wire new_Jinkela_wire_6529;
    wire new_Jinkela_wire_8325;
    wire new_Jinkela_wire_20940;
    wire new_Jinkela_wire_7659;
    wire new_Jinkela_wire_7870;
    wire new_Jinkela_wire_2255;
    wire new_Jinkela_wire_14421;
    wire new_Jinkela_wire_10081;
    wire new_Jinkela_wire_843;
    wire _0454_;
    wire new_Jinkela_wire_1249;
    wire _0146_;
    wire new_Jinkela_wire_20604;
    wire new_Jinkela_wire_15348;
    wire new_Jinkela_wire_8995;
    wire new_Jinkela_wire_14797;
    wire new_Jinkela_wire_8018;
    wire new_Jinkela_wire_17724;
    wire new_Jinkela_wire_14759;
    wire new_Jinkela_wire_11902;
    wire new_Jinkela_wire_3467;
    wire new_Jinkela_wire_6785;
    wire new_Jinkela_wire_10133;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_10538;
    wire new_Jinkela_wire_9824;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_8591;
    wire new_Jinkela_wire_4326;
    wire new_Jinkela_wire_11623;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_4923;
    wire new_Jinkela_wire_17727;
    wire new_Jinkela_wire_1723;
    wire new_Jinkela_wire_3399;
    wire new_Jinkela_wire_18724;
    wire new_Jinkela_wire_13873;
    wire new_Jinkela_wire_9422;
    wire new_Jinkela_wire_17894;
    wire new_Jinkela_wire_15477;
    wire new_Jinkela_wire_10370;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_18832;
    wire new_Jinkela_wire_5088;
    wire new_Jinkela_wire_20752;
    wire new_Jinkela_wire_14390;
    wire new_Jinkela_wire_6602;
    wire new_Jinkela_wire_4286;
    wire new_Jinkela_wire_14832;
    wire new_Jinkela_wire_3090;
    wire new_Jinkela_wire_3879;
    wire new_Jinkela_wire_5249;
    wire new_Jinkela_wire_5163;
    wire new_Jinkela_wire_18803;
    wire new_Jinkela_wire_9990;
    wire new_Jinkela_wire_19319;
    wire new_Jinkela_wire_9788;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_15592;
    wire new_Jinkela_wire_3791;
    wire new_Jinkela_wire_8743;
    wire new_Jinkela_wire_2980;
    wire new_Jinkela_wire_18363;
    wire new_Jinkela_wire_4862;
    wire new_Jinkela_wire_17830;
    wire new_Jinkela_wire_16878;
    wire new_Jinkela_wire_12250;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_21149;
    wire new_Jinkela_wire_19633;
    wire new_Jinkela_wire_4985;
    wire new_Jinkela_wire_2748;
    wire new_Jinkela_wire_15073;
    wire new_Jinkela_wire_21070;
    wire new_Jinkela_wire_21129;
    wire new_Jinkela_wire_10611;
    wire new_Jinkela_wire_1114;
    wire new_Jinkela_wire_4902;
    wire new_Jinkela_wire_13669;
    wire _0243_;
    wire new_Jinkela_wire_15335;
    wire new_Jinkela_wire_7805;
    wire new_Jinkela_wire_1995;
    wire new_Jinkela_wire_16559;
    wire new_Jinkela_wire_19485;
    wire new_Jinkela_wire_12212;
    wire new_Jinkela_wire_10679;
    wire _1244_;
    wire _0573_;
    wire new_Jinkela_wire_15070;
    wire new_Jinkela_wire_3873;
    wire new_Jinkela_wire_10348;
    wire new_Jinkela_wire_10075;
    wire new_Jinkela_wire_9663;
    wire new_Jinkela_wire_5178;
    wire new_Jinkela_wire_12640;
    wire new_Jinkela_wire_17886;
    wire new_Jinkela_wire_10872;
    wire _1809_;
    wire new_Jinkela_wire_13810;
    wire new_Jinkela_wire_10207;
    wire new_Jinkela_wire_21223;
    wire _1617_;
    wire new_Jinkela_wire_7959;
    wire new_Jinkela_wire_11223;
    wire _1714_;
    wire new_Jinkela_wire_17982;
    wire new_Jinkela_wire_2888;
    wire new_Jinkela_wire_3996;
    wire new_Jinkela_wire_20677;
    wire new_Jinkela_wire_6148;
    wire new_Jinkela_wire_18881;
    wire new_Jinkela_wire_17702;
    wire new_Jinkela_wire_12931;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_21210;
    wire new_Jinkela_wire_14389;
    wire new_Jinkela_wire_2416;
    wire new_Jinkela_wire_18607;
    wire new_Jinkela_wire_5080;
    wire new_Jinkela_wire_2015;
    wire new_Jinkela_wire_8233;
    wire new_Jinkela_wire_18031;
    wire new_Jinkela_wire_21143;
    wire new_Jinkela_wire_6722;
    wire new_Jinkela_wire_7014;
    wire new_Jinkela_wire_2364;
    wire new_Jinkela_wire_14789;
    wire new_Jinkela_wire_9902;
    wire new_Jinkela_wire_10398;
    wire new_Jinkela_wire_17626;
    wire new_Jinkela_wire_17074;
    wire new_Jinkela_wire_15653;
    wire new_Jinkela_wire_2490;
    wire new_Jinkela_wire_14176;
    wire new_Jinkela_wire_15748;
    wire new_Jinkela_wire_17159;
    wire new_Jinkela_wire_15115;
    wire new_Jinkela_wire_6719;
    wire new_Jinkela_wire_2258;
    wire new_Jinkela_wire_13313;
    wire new_Jinkela_wire_14732;
    wire new_Jinkela_wire_20746;
    wire new_Jinkela_wire_20144;
    wire new_Jinkela_wire_8939;
    wire new_Jinkela_wire_16924;
    wire new_Jinkela_wire_16079;
    wire new_Jinkela_wire_11356;
    wire new_Jinkela_wire_10273;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_18097;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_14065;
    wire new_Jinkela_wire_14216;
    wire new_Jinkela_wire_19399;
    wire new_Jinkela_wire_7581;
    wire new_Jinkela_wire_18887;
    wire new_Jinkela_wire_9706;
    wire new_Jinkela_wire_21184;
    wire new_Jinkela_wire_17811;
    wire new_Jinkela_wire_20398;
    wire _0802_;
    wire new_Jinkela_wire_14050;
    wire new_Jinkela_wire_9021;
    wire new_Jinkela_wire_8477;
    wire new_Jinkela_wire_6799;
    wire new_Jinkela_wire_11556;
    wire new_Jinkela_wire_6023;
    wire new_Jinkela_wire_12902;
    wire new_Jinkela_wire_3371;
    wire new_Jinkela_wire_5840;
    wire new_Jinkela_wire_20276;
    wire new_Jinkela_wire_6315;
    wire new_Jinkela_wire_20177;
    wire new_Jinkela_wire_9200;
    wire new_Jinkela_wire_11370;
    wire new_Jinkela_wire_6653;
    wire new_Jinkela_wire_8757;
    wire new_Jinkela_wire_12758;
    wire new_Jinkela_wire_9970;
    wire new_Jinkela_wire_12483;
    wire new_Jinkela_wire_16429;
    wire new_Jinkela_wire_18746;
    wire new_Jinkela_wire_17523;
    wire new_Jinkela_wire_6819;
    wire new_Jinkela_wire_19089;
    wire new_Jinkela_wire_5495;
    wire new_Jinkela_wire_13902;
    wire new_Jinkela_wire_17275;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_7384;
    wire new_Jinkela_wire_7723;
    wire _0055_;
    wire new_Jinkela_wire_18892;
    wire new_Jinkela_wire_4074;
    wire new_Jinkela_wire_17131;
    wire new_Jinkela_wire_7289;
    wire new_Jinkela_wire_11573;
    wire new_Jinkela_wire_17918;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_4793;
    wire new_Jinkela_wire_10325;
    wire new_Jinkela_wire_4557;
    wire _0228_;
    wire new_Jinkela_wire_7987;
    wire new_Jinkela_wire_7440;
    wire new_Jinkela_wire_11108;
    wire new_Jinkela_wire_4465;
    wire new_Jinkela_wire_13067;
    wire new_Jinkela_wire_16871;
    wire new_Jinkela_wire_6546;
    wire new_Jinkela_wire_12245;
    wire new_Jinkela_wire_18147;
    wire new_Jinkela_wire_14164;
    wire new_Jinkela_wire_3012;
    wire new_Jinkela_wire_14774;
    wire new_Jinkela_wire_9585;
    wire new_Jinkela_wire_10352;
    wire new_Jinkela_wire_20454;
    wire new_Jinkela_wire_15966;
    wire new_Jinkela_wire_3705;
    wire new_Jinkela_wire_16514;
    wire new_Jinkela_wire_20426;
    wire new_Jinkela_wire_14006;
    wire new_Jinkela_wire_7218;
    wire new_Jinkela_wire_8687;
    wire new_Jinkela_wire_15150;
    wire new_Jinkela_wire_5286;
    wire new_Jinkela_wire_13391;
    wire _1277_;
    wire new_Jinkela_wire_18002;
    wire _1282_;
    wire new_Jinkela_wire_13196;
    wire new_Jinkela_wire_13436;
    wire new_Jinkela_wire_15688;
    wire new_Jinkela_wire_18752;
    wire new_Jinkela_wire_9952;
    wire new_Jinkela_wire_18315;
    wire new_Jinkela_wire_14184;
    wire new_Jinkela_wire_5798;
    wire new_Jinkela_wire_3941;
    wire new_Jinkela_wire_3037;
    wire new_Jinkela_wire_14460;
    wire new_Jinkela_wire_17960;
    wire new_Jinkela_wire_5532;
    wire _1001_;
    wire _1063_;
    wire new_Jinkela_wire_6037;
    wire _0190_;
    wire new_Jinkela_wire_7020;
    wire new_Jinkela_wire_9608;
    wire new_Jinkela_wire_6379;
    wire new_Jinkela_wire_18461;
    wire new_Jinkela_wire_11378;
    wire new_Jinkela_wire_6648;
    wire new_Jinkela_wire_2335;
    wire _0838_;
    wire new_Jinkela_wire_2726;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_7594;
    wire new_Jinkela_wire_8151;
    wire _0052_;
    wire new_Jinkela_wire_4615;
    wire new_Jinkela_wire_18796;
    wire new_Jinkela_wire_8247;
    wire new_Jinkela_wire_12494;
    wire new_Jinkela_wire_8076;
    wire new_Jinkela_wire_18773;
    wire new_Jinkela_wire_15629;
    wire _1450_;
    wire new_Jinkela_wire_5552;
    wire new_Jinkela_wire_12003;
    wire new_Jinkela_wire_4015;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_9052;
    wire new_Jinkela_wire_3250;
    wire new_Jinkela_wire_10981;
    wire new_Jinkela_wire_19915;
    wire _1812_;
    wire new_Jinkela_wire_18663;
    wire new_Jinkela_wire_13764;
    wire new_Jinkela_wire_4189;
    wire new_Jinkela_wire_15314;
    wire new_Jinkela_wire_12987;
    wire new_Jinkela_wire_19098;
    wire new_Jinkela_wire_6508;
    wire new_Jinkela_wire_5426;
    wire new_Jinkela_wire_17218;
    wire new_Jinkela_wire_2423;
    wire new_Jinkela_wire_10836;
    wire new_Jinkela_wire_3765;
    wire new_Jinkela_wire_2930;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_6526;
    wire new_Jinkela_wire_6457;
    wire new_Jinkela_wire_17760;
    wire new_Jinkela_wire_8945;
    wire new_Jinkela_wire_3683;
    wire new_Jinkela_wire_1862;
    wire new_Jinkela_wire_14875;
    wire new_Jinkela_wire_4541;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_15011;
    wire new_Jinkela_wire_16883;
    wire new_Jinkela_wire_16756;
    wire new_Jinkela_wire_13462;
    wire new_Jinkela_wire_11799;
    wire new_Jinkela_wire_8178;
    wire new_Jinkela_wire_7394;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_11357;
    wire _1172_;
    wire new_Jinkela_wire_7874;
    wire new_Jinkela_wire_4445;
    wire new_Jinkela_wire_19284;
    wire _1102_;
    wire new_Jinkela_wire_3025;
    wire new_Jinkela_wire_8530;
    wire new_Jinkela_wire_3262;
    wire _1057_;
    wire new_Jinkela_wire_14148;
    wire new_Jinkela_wire_3707;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_2636;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_15201;
    wire new_Jinkela_wire_6865;
    wire new_Jinkela_wire_17385;
    wire new_Jinkela_wire_14230;
    wire new_Jinkela_wire_14267;
    wire new_Jinkela_wire_17608;
    wire new_Jinkela_wire_13091;
    wire new_Jinkela_wire_15443;
    wire new_Jinkela_wire_15680;
    wire new_Jinkela_wire_6225;
    wire new_Jinkela_wire_20461;
    wire new_Jinkela_wire_19565;
    wire new_Jinkela_wire_14531;
    wire new_Jinkela_wire_10883;
    wire new_Jinkela_wire_19932;
    wire new_Jinkela_wire_11290;
    wire new_Jinkela_wire_6975;
    wire new_Jinkela_wire_6938;
    wire new_Jinkela_wire_3202;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_10482;
    wire new_Jinkela_wire_4046;
    wire new_Jinkela_wire_2631;
    wire _0142_;
    wire new_Jinkela_wire_2358;
    wire new_Jinkela_wire_20402;
    wire new_Jinkela_wire_6663;
    wire new_Jinkela_wire_5582;
    wire new_Jinkela_wire_17142;
    wire new_Jinkela_wire_16319;
    wire new_Jinkela_wire_1865;
    wire new_Jinkela_wire_17819;
    wire new_Jinkela_wire_15711;
    wire new_Jinkela_wire_14429;
    wire new_Jinkela_wire_10049;
    wire new_Jinkela_wire_14343;
    wire new_Jinkela_wire_8638;
    wire new_Jinkela_wire_2595;
    wire new_Jinkela_wire_16929;
    wire new_Jinkela_wire_7867;
    wire new_Jinkela_wire_1832;
    wire new_Jinkela_wire_6288;
    wire new_Jinkela_wire_18967;
    wire new_Jinkela_wire_13044;
    wire new_Jinkela_wire_19124;
    wire new_Jinkela_wire_10406;
    wire new_Jinkela_wire_16687;
    wire _1632_;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_14053;
    wire new_Jinkela_wire_12958;
    wire new_Jinkela_wire_19338;
    wire new_Jinkela_wire_13427;
    wire new_Jinkela_wire_18384;
    wire new_Jinkela_wire_9105;
    wire new_Jinkela_wire_8722;
    wire new_Jinkela_wire_4195;
    wire new_Jinkela_wire_13962;
    wire new_Jinkela_wire_6367;
    wire new_Jinkela_wire_16700;
    wire new_Jinkela_wire_13399;
    wire _0158_;
    wire new_Jinkela_wire_17150;
    wire new_Jinkela_wire_20599;
    wire new_Jinkela_wire_5334;
    wire new_Jinkela_wire_10010;
    wire new_Jinkela_wire_2067;
    wire new_Jinkela_wire_17172;
    wire new_Jinkela_wire_10132;
    wire new_Jinkela_wire_19033;
    wire new_Jinkela_wire_12599;
    wire new_Jinkela_wire_14748;
    wire new_Jinkela_wire_11872;
    wire new_Jinkela_wire_17461;
    wire new_Jinkela_wire_8940;
    wire new_Jinkela_wire_8623;
    wire new_Jinkela_wire_5227;
    wire new_Jinkela_wire_6382;
    wire _1481_;
    wire new_Jinkela_wire_9014;
    wire new_Jinkela_wire_20655;
    wire new_Jinkela_wire_13150;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_19873;
    wire _1529_;
    wire new_Jinkela_wire_7554;
    wire new_Jinkela_wire_9793;
    wire new_Jinkela_wire_13787;
    wire new_Jinkela_wire_4527;
    wire _1684_;
    wire new_Jinkela_wire_3806;
    wire new_Jinkela_wire_16124;
    wire new_Jinkela_wire_16108;
    wire new_Jinkela_wire_11323;
    wire new_Jinkela_wire_9076;
    wire new_Jinkela_wire_13912;
    wire new_Jinkela_wire_12328;
    wire new_Jinkela_wire_739;
    wire new_Jinkela_wire_11531;
    wire new_Jinkela_wire_15575;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_1924;
    wire new_Jinkela_wire_6262;
    wire new_Jinkela_wire_1015;
    wire _1537_;
    wire new_Jinkela_wire_18716;
    wire new_Jinkela_wire_12976;
    wire new_Jinkela_wire_10701;
    wire new_Jinkela_wire_16921;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_11066;
    wire new_Jinkela_wire_19632;
    wire new_Jinkela_wire_16401;
    wire new_Jinkela_wire_15019;
    wire new_Jinkela_wire_6345;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_8666;
    wire new_Jinkela_wire_4169;
    wire new_Jinkela_wire_5645;
    wire new_Jinkela_wire_14577;
    wire new_Jinkela_wire_7286;
    wire new_Jinkela_wire_21174;
    wire new_Jinkela_wire_3464;
    wire new_Jinkela_wire_8514;
    wire new_Jinkela_wire_15101;
    wire new_Jinkela_wire_21081;
    wire new_Jinkela_wire_3027;
    wire new_Jinkela_wire_17457;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_6182;
    wire new_Jinkela_wire_16214;
    wire new_Jinkela_wire_11480;
    wire new_Jinkela_wire_14020;
    wire new_Jinkela_wire_6280;
    wire new_Jinkela_wire_7255;
    wire new_Jinkela_wire_14085;
    wire new_Jinkela_wire_3054;
    wire new_Jinkela_wire_17330;
    wire new_Jinkela_wire_5248;
    wire _0312_;
    wire new_Jinkela_wire_18647;
    wire new_Jinkela_wire_19946;
    wire new_Jinkela_wire_23;
    wire new_Jinkela_wire_13213;
    wire _0955_;
    wire new_Jinkela_wire_17227;
    wire new_Jinkela_wire_8394;
    wire new_Jinkela_wire_7911;
    wire new_Jinkela_wire_11192;
    wire _1383_;
    wire new_Jinkela_wire_5902;
    wire new_Jinkela_wire_8039;
    wire new_Jinkela_wire_21293;
    wire new_Jinkela_wire_12088;
    wire new_Jinkela_wire_4091;
    wire new_Jinkela_wire_5122;
    wire new_Jinkela_wire_2130;
    wire new_Jinkela_wire_6849;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_16171;
    wire new_Jinkela_wire_7280;
    wire new_Jinkela_wire_18321;
    wire new_Jinkela_wire_5858;
    wire _1090_;
    wire _1271_;
    wire new_Jinkela_wire_2352;
    wire new_Jinkela_wire_11729;
    wire new_Jinkela_wire_20094;
    wire new_Jinkela_wire_6547;
    wire new_Jinkela_wire_16384;
    wire new_Jinkela_wire_15562;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_6594;
    wire new_Jinkela_wire_4790;
    wire new_Jinkela_wire_2276;
    wire new_Jinkela_wire_8061;
    wire new_Jinkela_wire_16796;
    wire new_Jinkela_wire_20815;
    wire new_Jinkela_wire_13171;
    wire new_Jinkela_wire_8672;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_14594;
    wire _0540_;
    wire new_Jinkela_wire_21260;
    wire new_Jinkela_wire_5651;
    wire new_Jinkela_wire_19579;
    wire new_Jinkela_wire_5925;
    wire new_Jinkela_wire_7089;
    wire new_Jinkela_wire_20543;
    wire new_Jinkela_wire_9433;
    wire new_Jinkela_wire_10353;
    wire new_Jinkela_wire_12696;
    wire new_Jinkela_wire_14906;
    wire new_Jinkela_wire_10857;
    wire _1150_;
    wire new_Jinkela_wire_16389;
    wire new_Jinkela_wire_18924;
    wire new_Jinkela_wire_8274;
    wire _0425_;
    wire new_Jinkela_wire_18416;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_20327;
    wire new_Jinkela_wire_13400;
    wire new_Jinkela_wire_8574;
    wire new_Jinkela_wire_17584;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_11041;
    wire new_Jinkela_wire_16573;
    wire new_Jinkela_wire_11664;
    wire new_Jinkela_wire_3240;
    wire new_Jinkela_wire_5590;
    wire new_Jinkela_wire_21264;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_18119;
    wire new_Jinkela_wire_6774;
    wire _1814_;
    wire new_Jinkela_wire_10707;
    wire new_Jinkela_wire_17245;
    wire new_Jinkela_wire_18687;
    wire new_Jinkela_wire_16705;
    wire new_Jinkela_wire_19809;
    wire new_Jinkela_wire_14047;
    wire new_Jinkela_wire_19760;
    wire new_Jinkela_wire_20484;
    wire new_Jinkela_wire_7108;
    wire new_Jinkela_wire_1889;
    wire new_Jinkela_wire_7720;
    wire new_Jinkela_wire_17586;
    wire new_Jinkela_wire_9128;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_18300;
    wire new_Jinkela_wire_6279;
    wire new_Jinkela_wire_12979;
    wire new_Jinkela_wire_18535;
    wire new_Jinkela_wire_10619;
    wire new_Jinkela_wire_12465;
    wire new_Jinkela_wire_20105;
    wire new_Jinkela_wire_7349;
    wire new_Jinkela_wire_18979;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_20483;
    wire new_Jinkela_wire_3479;
    wire new_Jinkela_wire_8052;
    wire new_Jinkela_wire_13040;
    wire new_Jinkela_wire_14126;
    wire new_Jinkela_wire_18485;
    wire new_Jinkela_wire_9959;
    wire new_Jinkela_wire_4497;
    wire new_Jinkela_wire_17902;
    wire new_Jinkela_wire_6791;
    wire _0430_;
    wire new_Jinkela_wire_14100;
    wire new_Jinkela_wire_2066;
    wire new_Jinkela_wire_15474;
    wire new_Jinkela_wire_10570;
    wire new_Jinkela_wire_10510;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_5447;
    wire _0583_;
    wire new_Jinkela_wire_3717;
    wire new_Jinkela_wire_5241;
    wire new_Jinkela_wire_13938;
    wire new_Jinkela_wire_10076;
    wire new_Jinkela_wire_5474;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_7797;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_6108;
    wire new_Jinkela_wire_20707;
    wire new_Jinkela_wire_6122;
    wire new_Jinkela_wire_14807;
    wire new_Jinkela_wire_5468;
    wire new_Jinkela_wire_9593;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_16344;
    wire _1691_;
    wire new_Jinkela_wire_5562;
    wire new_Jinkela_wire_15625;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_13813;
    wire new_Jinkela_wire_19700;
    wire new_Jinkela_wire_5231;
    wire new_Jinkela_wire_8248;
    wire new_Jinkela_wire_6705;
    wire new_Jinkela_wire_1037;
    wire new_Jinkela_wire_10841;
    wire new_Jinkela_wire_19762;
    wire new_Jinkela_wire_7985;
    wire new_Jinkela_wire_20758;
    wire new_Jinkela_wire_19002;
    wire new_Jinkela_wire_6363;
    wire new_Jinkela_wire_7889;
    wire new_Jinkela_wire_6178;
    wire new_Jinkela_wire_4612;
    wire new_Jinkela_wire_19273;
    wire new_Jinkela_wire_3706;
    wire new_Jinkela_wire_19231;
    wire new_Jinkela_wire_19981;
    wire _0177_;
    wire new_Jinkela_wire_11626;
    wire new_Jinkela_wire_16780;
    wire new_Jinkela_wire_13176;
    wire new_Jinkela_wire_14213;
    wire new_Jinkela_wire_3160;
    wire new_Jinkela_wire_17562;
    wire new_Jinkela_wire_9371;
    wire new_Jinkela_wire_18719;
    wire new_Jinkela_wire_16376;
    wire new_Jinkela_wire_18019;
    wire new_Jinkela_wire_7372;
    wire new_Jinkela_wire_6646;
    wire new_Jinkela_wire_15494;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_18883;
    wire new_Jinkela_wire_20273;
    wire new_Jinkela_wire_17147;
    wire _0047_;
    wire new_Jinkela_wire_20678;
    wire _1307_;
    wire new_Jinkela_wire_1530;
    wire new_Jinkela_wire_5617;
    wire new_Jinkela_wire_14872;
    wire new_Jinkela_wire_13026;
    wire new_Jinkela_wire_8220;
    wire new_Jinkela_wire_9098;
    wire new_Jinkela_wire_18132;
    wire _0251_;
    wire new_Jinkela_wire_19756;
    wire new_Jinkela_wire_6226;
    wire new_Jinkela_wire_9185;
    wire new_Jinkela_wire_5693;
    wire new_Jinkela_wire_2914;
    wire new_Jinkela_wire_18521;
    wire new_Jinkela_wire_7158;
    wire new_Jinkela_wire_9430;
    wire new_Jinkela_wire_9754;
    wire new_Jinkela_wire_2972;
    wire new_Jinkela_wire_2919;
    wire new_Jinkela_wire_19815;
    wire new_Jinkela_wire_20473;
    wire new_Jinkela_wire_3378;
    wire new_Jinkela_wire_7552;
    wire new_Jinkela_wire_9136;
    wire new_Jinkela_wire_7460;
    wire new_Jinkela_wire_19038;
    wire new_Jinkela_wire_19555;
    wire new_Jinkela_wire_12687;
    wire new_Jinkela_wire_7787;
    wire new_Jinkela_wire_16198;
    wire new_Jinkela_wire_6157;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_5522;
    wire new_Jinkela_wire_5408;
    wire new_Jinkela_wire_9709;
    wire new_Jinkela_wire_18090;
    wire new_Jinkela_wire_2670;
    wire new_Jinkela_wire_15573;
    wire new_Jinkela_wire_14005;
    wire new_Jinkela_wire_3746;
    wire new_Jinkela_wire_13413;
    wire new_Jinkela_wire_4922;
    wire _1410_;
    wire new_Jinkela_wire_3394;
    wire new_Jinkela_wire_7875;
    wire new_Jinkela_wire_9864;
    wire new_Jinkela_wire_20014;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_11653;
    wire new_Jinkela_wire_3665;
    wire new_Jinkela_wire_3864;
    wire new_Jinkela_wire_17077;
    wire new_Jinkela_wire_5866;
    wire new_Jinkela_wire_5881;
    wire _1551_;
    wire new_Jinkela_wire_8775;
    wire new_Jinkela_wire_3657;
    wire new_Jinkela_wire_8134;
    wire new_Jinkela_wire_20908;
    wire new_Jinkela_wire_19781;
    wire new_Jinkela_wire_13425;
    wire new_Jinkela_wire_6732;
    wire new_Jinkela_wire_15166;
    wire new_Jinkela_wire_14018;
    wire new_Jinkela_wire_21288;
    wire new_Jinkela_wire_13668;
    wire new_Jinkela_wire_11076;
    wire new_Jinkela_wire_40;
    wire new_Jinkela_wire_15957;
    wire new_Jinkela_wire_2408;
    wire new_Jinkela_wire_18392;
    wire _0961_;
    wire new_Jinkela_wire_11364;
    wire new_Jinkela_wire_10301;
    wire new_Jinkela_wire_11246;
    wire _0450_;
    wire new_Jinkela_wire_12594;
    wire _1808_;
    wire new_Jinkela_wire_5150;
    wire new_Jinkela_wire_5058;
    wire new_Jinkela_wire_16248;
    wire new_Jinkela_wire_12299;
    wire new_Jinkela_wire_2628;
    wire new_Jinkela_wire_11796;
    wire new_Jinkela_wire_4444;
    wire new_Jinkela_wire_2633;
    wire _0607_;
    wire new_Jinkela_wire_15089;
    wire new_Jinkela_wire_17495;
    wire new_Jinkela_wire_2314;
    wire new_Jinkela_wire_10329;
    wire new_Jinkela_wire_15892;
    wire new_Jinkela_wire_19474;
    wire new_Jinkela_wire_11742;
    wire new_Jinkela_wire_2098;
    wire new_Jinkela_wire_12290;
    wire new_Jinkela_wire_20171;
    wire new_Jinkela_wire_7482;
    wire new_Jinkela_wire_18217;
    wire _0523_;
    wire new_Jinkela_wire_12995;
    wire new_Jinkela_wire_12456;
    wire new_Jinkela_wire_8148;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_10381;
    wire new_Jinkela_wire_13659;
    wire new_Jinkela_wire_8966;
    wire new_Jinkela_wire_13922;
    wire new_Jinkela_wire_10739;
    wire new_Jinkela_wire_16444;
    wire new_Jinkela_wire_14758;
    wire new_Jinkela_wire_1262;
    wire _0221_;
    wire new_Jinkela_wire_6056;
    wire new_Jinkela_wire_5435;
    wire new_Jinkela_wire_20447;
    wire new_Jinkela_wire_3009;
    wire new_Jinkela_wire_17344;
    wire new_Jinkela_wire_7514;
    wire new_Jinkela_wire_19714;
    wire new_Jinkela_wire_7941;
    wire new_Jinkela_wire_4754;
    wire new_Jinkela_wire_18548;
    wire new_Jinkela_wire_13512;
    wire new_Jinkela_wire_15667;
    wire new_Jinkela_wire_9156;
    wire new_Jinkela_wire_6664;
    wire _1005_;
    wire new_Jinkela_wire_12379;
    wire new_Jinkela_wire_20540;
    wire new_Jinkela_wire_9071;
    wire new_Jinkela_wire_10228;
    wire new_Jinkela_wire_9018;
    wire new_Jinkela_wire_9961;
    wire _1586_;
    wire new_Jinkela_wire_8107;
    wire new_Jinkela_wire_2398;
    wire new_Jinkela_wire_16643;
    wire new_Jinkela_wire_13493;
    wire new_Jinkela_wire_2819;
    wire new_Jinkela_wire_9904;
    wire _1739_;
    wire new_Jinkela_wire_20294;
    wire _1526_;
    wire new_Jinkela_wire_925;
    wire new_Jinkela_wire_16053;
    wire new_Jinkela_wire_20642;
    wire new_Jinkela_wire_12113;
    wire new_Jinkela_wire_2468;
    wire new_Jinkela_wire_20157;
    wire new_Jinkela_wire_19391;
    wire new_Jinkela_wire_17660;
    wire new_Jinkela_wire_12373;
    wire new_Jinkela_wire_9958;
    wire new_Jinkela_wire_13049;
    wire new_Jinkela_wire_12209;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_15162;
    wire new_Jinkela_wire_20009;
    wire new_Jinkela_wire_12666;
    wire new_Jinkela_wire_9568;
    wire new_Jinkela_wire_3329;
    wire new_Jinkela_wire_19520;
    wire new_Jinkela_wire_5211;
    wire new_Jinkela_wire_16285;
    wire new_Jinkela_wire_16024;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_15702;
    wire new_Jinkela_wire_5717;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_18902;
    wire new_Jinkela_wire_10585;
    wire new_Jinkela_wire_20139;
    wire new_Jinkela_wire_9974;
    wire new_Jinkela_wire_11149;
    wire new_Jinkela_wire_6357;
    wire _1080_;
    wire new_Jinkela_wire_8596;
    wire new_Jinkela_wire_9980;
    wire new_Jinkela_wire_11298;
    wire _1407_;
    wire new_Jinkela_wire_20645;
    wire new_Jinkela_wire_11865;
    wire new_Jinkela_wire_16884;
    wire new_Jinkela_wire_8742;
    wire new_Jinkela_wire_14462;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_9651;
    wire new_Jinkela_wire_11833;
    wire new_Jinkela_wire_6576;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_13730;
    wire new_Jinkela_wire_2693;
    wire new_Jinkela_wire_4858;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_9778;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_17055;
    wire new_Jinkela_wire_17155;
    wire new_Jinkela_wire_8096;
    wire new_Jinkela_wire_20881;
    wire new_Jinkela_wire_7143;
    wire new_Jinkela_wire_20800;
    wire new_Jinkela_wire_15249;
    wire new_Jinkela_wire_7591;
    wire new_Jinkela_wire_16462;
    wire _0757_;
    wire new_Jinkela_wire_7167;
    wire new_Jinkela_wire_20062;
    wire new_Jinkela_wire_10660;
    wire _1447_;
    wire _1112_;
    wire new_Jinkela_wire_21160;
    wire new_Jinkela_wire_2558;
    wire new_Jinkela_wire_15176;
    wire new_Jinkela_wire_11232;
    wire _1304_;
    wire _0501_;
    wire new_Jinkela_wire_19356;
    wire new_Jinkela_wire_9377;
    wire new_Jinkela_wire_11158;
    wire new_Jinkela_wire_18680;
    wire new_Jinkela_wire_15786;
    wire new_Jinkela_wire_8095;
    wire _0164_;
    wire new_Jinkela_wire_18232;
    wire new_Jinkela_wire_19298;
    wire new_Jinkela_wire_12896;
    wire new_Jinkela_wire_11250;
    wire new_Jinkela_wire_5463;
    wire new_Jinkela_wire_7453;
    wire new_Jinkela_wire_7432;
    wire new_Jinkela_wire_7574;
    wire new_Jinkela_wire_20045;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_12466;
    wire new_Jinkela_wire_12777;
    wire new_Jinkela_wire_17544;
    wire new_Jinkela_wire_10951;
    wire new_Jinkela_wire_6030;
    wire new_Jinkela_wire_11691;
    wire new_Jinkela_wire_14639;
    wire new_Jinkela_wire_11470;
    wire new_Jinkela_wire_16613;
    wire new_Jinkela_wire_9486;
    wire new_Jinkela_wire_19886;
    wire new_Jinkela_wire_9250;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_12163;
    wire new_Jinkela_wire_20128;
    wire new_Jinkela_wire_14008;
    wire new_Jinkela_wire_6531;
    wire new_Jinkela_wire_6209;
    wire new_Jinkela_wire_5780;
    wire new_Jinkela_wire_19037;
    wire new_Jinkela_wire_17267;
    wire new_Jinkela_wire_8706;
    wire new_Jinkela_wire_10873;
    wire new_Jinkela_wire_13900;
    wire new_Jinkela_wire_11248;
    wire new_Jinkela_wire_12408;
    wire new_Jinkela_wire_14548;
    wire new_Jinkela_wire_11832;
    wire new_Jinkela_wire_18682;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_6915;
    wire new_Jinkela_wire_15186;
    wire _1024_;
    wire _1359_;
    wire new_Jinkela_wire_5831;
    wire new_Jinkela_wire_18194;
    wire new_Jinkela_wire_9787;
    wire new_Jinkela_wire_20618;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_10581;
    wire new_Jinkela_wire_16814;
    wire new_Jinkela_wire_9304;
    wire new_Jinkela_wire_4569;
    wire new_Jinkela_wire_14172;
    wire new_Jinkela_wire_15146;
    wire new_Jinkela_wire_5927;
    wire new_Jinkela_wire_16982;
    wire new_Jinkela_wire_6462;
    wire new_Jinkela_wire_1089;
    wire new_Jinkela_wire_17964;
    wire new_Jinkela_wire_7543;
    wire new_Jinkela_wire_4798;
    wire new_Jinkela_wire_3324;
    wire new_Jinkela_wire_19892;
    wire new_Jinkela_wire_20138;
    wire new_Jinkela_wire_15403;
    wire new_Jinkela_wire_17476;
    wire new_Jinkela_wire_18084;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_6430;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_19866;
    wire new_Jinkela_wire_5405;
    wire _1441_;
    wire new_Jinkela_wire_8702;
    wire new_Jinkela_wire_4284;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_9399;
    wire new_Jinkela_wire_13005;
    wire new_Jinkela_wire_18504;
    wire new_Jinkela_wire_8266;
    wire new_Jinkela_wire_6510;
    wire _0121_;
    wire _0210_;
    wire new_Jinkela_wire_6174;
    wire new_Jinkela_wire_21207;
    wire new_Jinkela_wire_7069;
    wire _0888_;
    wire _0750_;
    wire new_Jinkela_wire_2615;
    wire new_Jinkela_wire_20956;
    wire new_Jinkela_wire_4390;
    wire new_Jinkela_wire_18843;
    wire new_Jinkela_wire_8230;
    wire new_Jinkela_wire_2543;
    wire _0104_;
    wire new_Jinkela_wire_7576;
    wire new_Jinkela_wire_18350;
    wire new_Jinkela_wire_16561;
    wire new_Jinkela_wire_4399;
    wire new_Jinkela_wire_11947;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_17217;
    wire new_Jinkela_wire_4523;
    wire new_Jinkela_wire_20180;
    wire _0882_;
    wire new_Jinkela_wire_12371;
    wire new_Jinkela_wire_17701;
    wire _1224_;
    wire new_Jinkela_wire_2139;
    wire _0205_;
    wire _1056_;
    wire new_Jinkela_wire_9398;
    wire new_Jinkela_wire_4018;
    wire new_Jinkela_wire_12014;
    wire new_Jinkela_wire_13355;
    wire new_Jinkela_wire_3882;
    wire new_Jinkela_wire_8639;
    wire new_Jinkela_wire_11920;
    wire _0293_;
    wire new_Jinkela_wire_6736;
    wire new_Jinkela_wire_9612;
    wire new_Jinkela_wire_7698;
    wire new_Jinkela_wire_15538;
    wire _1364_;
    wire new_Jinkela_wire_3064;
    wire new_Jinkela_wire_13101;
    wire new_Jinkela_wire_20228;
    wire new_Jinkela_wire_11242;
    wire new_Jinkela_wire_11555;
    wire new_Jinkela_wire_6478;
    wire new_Jinkela_wire_20699;
    wire new_Jinkela_wire_15910;
    wire new_Jinkela_wire_14642;
    wire new_Jinkela_wire_2051;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_13633;
    wire new_Jinkela_wire_3714;
    wire _0342_;
    wire new_Jinkela_wire_7197;
    wire new_Jinkela_wire_5155;
    wire new_Jinkela_wire_20970;
    wire _0605_;
    wire new_Jinkela_wire_20226;
    wire new_Jinkela_wire_7750;
    wire new_Jinkela_wire_19143;
    wire new_Jinkela_wire_6850;
    wire new_Jinkela_wire_3485;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_15818;
    wire _1209_;
    wire new_Jinkela_wire_20343;
    wire new_Jinkela_wire_18869;
    wire new_Jinkela_wire_3842;
    wire new_Jinkela_wire_9924;
    wire new_Jinkela_wire_10505;
    wire _0402_;
    wire new_Jinkela_wire_6213;
    wire new_Jinkela_wire_11221;
    wire new_Jinkela_wire_20795;
    wire _1370_;
    wire new_Jinkela_wire_18411;
    wire new_Jinkela_wire_15703;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_4872;
    wire new_Jinkela_wire_11196;
    wire new_Jinkela_wire_8892;
    wire new_Jinkela_wire_3774;
    wire new_Jinkela_wire_20880;
    wire new_Jinkela_wire_4171;
    wire new_Jinkela_wire_13788;
    wire new_Jinkela_wire_15672;
    wire new_Jinkela_wire_4100;
    wire new_Jinkela_wire_18942;
    wire new_Jinkela_wire_15760;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_19440;
    wire new_Jinkela_wire_430;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_21069;
    wire new_Jinkela_wire_6211;
    wire new_Jinkela_wire_8562;
    wire new_Jinkela_wire_18063;
    wire new_Jinkela_wire_2257;
    wire new_Jinkela_wire_4416;
    wire new_Jinkela_wire_16363;
    wire new_Jinkela_wire_13981;
    wire new_Jinkela_wire_11265;
    wire new_Jinkela_wire_7177;
    wire new_Jinkela_wire_6980;
    wire new_Jinkela_wire_7142;
    wire new_Jinkela_wire_20388;
    wire new_Jinkela_wire_12234;
    wire new_Jinkela_wire_7210;
    wire new_Jinkela_wire_14574;
    wire _0828_;
    wire new_Jinkela_wire_8433;
    wire new_Jinkela_wire_9531;
    wire new_Jinkela_wire_11953;
    wire new_Jinkela_wire_3803;
    wire new_Jinkela_wire_6584;
    wire new_Jinkela_wire_13494;
    wire new_Jinkela_wire_2751;
    wire new_Jinkela_wire_17202;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_11977;
    wire new_Jinkela_wire_19332;
    wire new_Jinkela_wire_5471;
    wire new_Jinkela_wire_10525;
    wire new_Jinkela_wire_9769;
    wire new_Jinkela_wire_15756;
    wire _1553_;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_18499;
    wire new_Jinkela_wire_3732;
    wire _1467_;
    wire new_Jinkela_wire_14815;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_16865;
    wire new_Jinkela_wire_17714;
    wire new_net_3954;
    wire new_Jinkela_wire_8082;
    wire new_Jinkela_wire_21049;
    wire new_Jinkela_wire_10516;
    wire _0111_;
    wire new_Jinkela_wire_11362;
    wire new_Jinkela_wire_15837;
    wire new_Jinkela_wire_18856;
    wire new_Jinkela_wire_2909;
    wire new_Jinkela_wire_14599;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_5348;
    wire new_Jinkela_wire_16549;
    wire new_Jinkela_wire_12967;
    wire new_Jinkela_wire_6862;
    wire new_Jinkela_wire_16240;
    wire new_Jinkela_wire_17405;
    wire new_Jinkela_wire_11674;
    wire new_Jinkela_wire_12532;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_20607;
    wire new_Jinkela_wire_20318;
    wire new_Jinkela_wire_10958;
    wire new_Jinkela_wire_8545;
    wire new_Jinkela_wire_10812;
    wire _0069_;
    wire new_Jinkela_wire_6358;
    wire new_Jinkela_wire_3195;
    wire new_Jinkela_wire_9995;
    wire new_Jinkela_wire_14239;
    wire new_Jinkela_wire_11126;
    wire new_Jinkela_wire_3033;
    wire new_Jinkela_wire_4424;
    wire new_Jinkela_wire_17996;
    wire new_Jinkela_wire_12990;
    wire new_Jinkela_wire_15656;
    wire new_Jinkela_wire_8292;
    wire _1226_;
    wire new_Jinkela_wire_17579;
    wire _0716_;
    wire new_Jinkela_wire_6394;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_5598;
    wire new_Jinkela_wire_10184;
    wire new_Jinkela_wire_9602;
    wire new_Jinkela_wire_16381;
    wire new_Jinkela_wire_12580;
    wire new_Jinkela_wire_5301;
    wire new_Jinkela_wire_15363;
    wire new_Jinkela_wire_11146;
    wire new_Jinkela_wire_4230;
    wire new_Jinkela_wire_5135;
    wire new_Jinkela_wire_5518;
    wire new_Jinkela_wire_19328;
    wire new_Jinkela_wire_8363;
    wire new_Jinkela_wire_12264;
    wire new_Jinkela_wire_7045;
    wire _0451_;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_7107;
    wire new_Jinkela_wire_11663;
    wire new_Jinkela_wire_11209;
    wire new_Jinkela_wire_13823;
    wire new_Jinkela_wire_14099;
    wire new_Jinkela_wire_16073;
    wire new_Jinkela_wire_14084;
    wire new_Jinkela_wire_8504;
    wire new_Jinkela_wire_19047;
    wire new_Jinkela_wire_15650;
    wire new_Jinkela_wire_5343;
    wire new_Jinkela_wire_3169;
    wire new_Jinkela_wire_18907;
    wire new_Jinkela_wire_13086;
    wire new_Jinkela_wire_14714;
    wire _1348_;
    wire new_Jinkela_wire_15263;
    wire new_Jinkela_wire_5795;
    wire new_Jinkela_wire_16997;
    wire _1763_;
    wire new_Jinkela_wire_16196;
    wire new_Jinkela_wire_12672;
    wire new_Jinkela_wire_9079;
    wire new_Jinkela_wire_5023;
    wire new_Jinkela_wire_15627;
    wire new_Jinkela_wire_7798;
    wire new_Jinkela_wire_7863;
    wire new_Jinkela_wire_6724;
    wire new_Jinkela_wire_6533;
    wire new_Jinkela_wire_2083;
    wire new_Jinkela_wire_16596;
    wire new_Jinkela_wire_16479;
    wire _0895_;
    wire new_Jinkela_wire_3227;
    wire new_Jinkela_wire_4693;
    wire new_Jinkela_wire_7411;
    wire new_Jinkela_wire_7230;
    wire _0812_;
    wire new_Jinkela_wire_10472;
    wire new_Jinkela_wire_14218;
    wire new_Jinkela_wire_13941;
    wire new_Jinkela_wire_11413;
    wire new_Jinkela_wire_16599;
    wire new_Jinkela_wire_17690;
    wire new_Jinkela_wire_17997;
    wire new_Jinkela_wire_21292;
    wire new_Jinkela_wire_9802;
    wire new_Jinkela_wire_17502;
    wire new_Jinkela_wire_4315;
    wire new_Jinkela_wire_15351;
    wire new_Jinkela_wire_14151;
    wire new_Jinkela_wire_12307;
    wire new_Jinkela_wire_16937;
    wire new_Jinkela_wire_17035;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_6252;
    wire new_Jinkela_wire_12411;
    wire new_Jinkela_wire_12482;
    wire new_Jinkela_wire_5846;
    wire new_Jinkela_wire_18947;
    wire new_Jinkela_wire_12039;
    wire new_Jinkela_wire_14368;
    wire new_Jinkela_wire_12940;
    wire new_Jinkela_wire_4917;
    wire new_Jinkela_wire_8793;
    wire new_Jinkela_wire_8886;
    wire new_Jinkela_wire_11914;
    wire new_Jinkela_wire_18644;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_5491;
    wire new_Jinkela_wire_2208;
    wire new_Jinkela_wire_17326;
    wire new_Jinkela_wire_11679;
    wire new_Jinkela_wire_10687;
    wire new_Jinkela_wire_3233;
    wire new_Jinkela_wire_13326;
    wire new_Jinkela_wire_13584;
    wire new_Jinkela_wire_8814;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_5548;
    wire new_Jinkela_wire_8921;
    wire new_Jinkela_wire_20910;
    wire new_Jinkela_wire_5957;
    wire new_Jinkela_wire_13144;
    wire new_Jinkela_wire_19788;
    wire new_Jinkela_wire_17036;
    wire new_Jinkela_wire_8635;
    wire new_Jinkela_wire_7691;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_12036;
    wire new_Jinkela_wire_4572;
    wire new_Jinkela_wire_13098;
    wire new_Jinkela_wire_16783;
    wire new_Jinkela_wire_18137;
    wire new_Jinkela_wire_3474;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_17771;
    wire new_Jinkela_wire_12079;
    wire new_Jinkela_wire_12848;
    wire new_Jinkela_wire_8578;
    wire new_Jinkela_wire_6880;
    wire _0066_;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_16912;
    wire new_Jinkela_wire_13728;
    wire new_Jinkela_wire_12644;
    wire new_Jinkela_wire_1439;
    wire new_Jinkela_wire_5735;
    wire _0524_;
    wire _1618_;
    wire new_Jinkela_wire_14914;
    wire new_Jinkela_wire_2144;
    wire new_Jinkela_wire_18182;
    wire new_Jinkela_wire_9444;
    wire new_Jinkela_wire_6852;
    wire new_Jinkela_wire_13748;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_2731;
    wire new_Jinkela_wire_2553;
    wire new_Jinkela_wire_5788;
    wire new_Jinkela_wire_6616;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_15020;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_4510;
    wire new_Jinkela_wire_19164;
    wire new_Jinkela_wire_2892;
    wire new_Jinkela_wire_7969;
    wire new_Jinkela_wire_13786;
    wire new_Jinkela_wire_14284;
    wire new_Jinkela_wire_9656;
    wire new_Jinkela_wire_16655;
    wire new_Jinkela_wire_8931;
    wire new_Jinkela_wire_14502;
    wire new_Jinkela_wire_2077;
    wire new_Jinkela_wire_5421;
    wire new_Jinkela_wire_8834;
    wire new_Jinkela_wire_15522;
    wire new_Jinkela_wire_13770;
    wire new_Jinkela_wire_5192;
    wire _0715_;
    wire new_Jinkela_wire_2226;
    wire new_Jinkela_wire_6831;
    wire new_Jinkela_wire_11335;
    wire new_Jinkela_wire_11366;
    wire new_Jinkela_wire_17235;
    wire new_Jinkela_wire_17060;
    wire new_Jinkela_wire_12654;
    wire new_Jinkela_wire_8219;
    wire new_Jinkela_wire_6703;
    wire new_Jinkela_wire_21096;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_3589;
    wire _1344_;
    wire new_Jinkela_wire_4957;
    wire new_Jinkela_wire_14499;
    wire new_Jinkela_wire_7061;
    wire new_Jinkela_wire_16681;
    wire new_Jinkela_wire_10414;
    wire new_Jinkela_wire_18502;
    wire new_Jinkela_wire_11281;
    wire new_Jinkela_wire_4913;
    wire new_Jinkela_wire_9312;
    wire new_Jinkela_wire_3546;
    wire new_Jinkela_wire_18420;
    wire new_Jinkela_wire_2816;
    wire new_Jinkela_wire_11523;
    wire new_Jinkela_wire_8697;
    wire new_Jinkela_wire_6661;
    wire new_Jinkela_wire_9184;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_4782;
    wire new_Jinkela_wire_18584;
    wire new_Jinkela_wire_12296;
    wire new_Jinkela_wire_8153;
    wire new_Jinkela_wire_10989;
    wire new_Jinkela_wire_18848;
    wire new_Jinkela_wire_5243;
    wire new_Jinkela_wire_15924;
    wire new_Jinkela_wire_17346;
    wire new_Jinkela_wire_14718;
    wire new_Jinkela_wire_4661;
    wire new_Jinkela_wire_10039;
    wire new_Jinkela_wire_12134;
    wire new_Jinkela_wire_1687;
    wire new_Jinkela_wire_7998;
    wire new_Jinkela_wire_8807;
    wire new_Jinkela_wire_4828;
    wire new_Jinkela_wire_2559;
    wire new_Jinkela_wire_7032;
    wire new_Jinkela_wire_3486;
    wire new_Jinkela_wire_10355;
    wire _1417_;
    wire new_Jinkela_wire_9721;
    wire new_Jinkela_wire_20442;
    wire new_Jinkela_wire_1750;
    wire new_Jinkela_wire_7240;
    wire new_Jinkela_wire_3763;
    wire _0990_;
    wire new_Jinkela_wire_20224;
    wire _0497_;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_9597;
    wire new_Jinkela_wire_4718;
    wire new_Jinkela_wire_5072;
    wire new_Jinkela_wire_5305;
    wire new_Jinkela_wire_13698;
    wire new_Jinkela_wire_8541;
    wire _1657_;
    wire new_Jinkela_wire_12198;
    wire new_Jinkela_wire_13406;
    wire new_Jinkela_wire_8784;
    wire new_Jinkela_wire_6497;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_8589;
    wire new_Jinkela_wire_15354;
    wire new_Jinkela_wire_522;
    wire _0866_;
    wire new_Jinkela_wire_11893;
    wire new_Jinkela_wire_3253;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_8533;
    wire new_Jinkela_wire_13923;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_14675;
    wire _1833_;
    wire _0746_;
    wire new_Jinkela_wire_8422;
    wire new_Jinkela_wire_14143;
    wire new_Jinkela_wire_21123;
    wire new_Jinkela_wire_7437;
    wire new_Jinkela_wire_7441;
    wire new_Jinkela_wire_13275;
    wire new_Jinkela_wire_19069;
    wire new_Jinkela_wire_13946;
    wire new_Jinkela_wire_19550;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_21244;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_5089;
    wire new_Jinkela_wire_15333;
    wire new_Jinkela_wire_12633;
    wire new_Jinkela_wire_15746;
    wire _0294_;
    wire new_Jinkela_wire_18591;
    wire new_Jinkela_wire_5696;
    wire new_Jinkela_wire_11934;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_7099;
    wire new_Jinkela_wire_16666;
    wire new_Jinkela_wire_13280;
    wire new_Jinkela_wire_20663;
    wire _0698_;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_12101;
    wire _0658_;
    wire new_Jinkela_wire_18919;
    wire new_Jinkela_wire_10270;
    wire new_Jinkela_wire_15218;
    wire new_Jinkela_wire_5917;
    wire new_Jinkela_wire_2437;
    wire new_Jinkela_wire_14861;
    wire new_Jinkela_wire_11016;
    wire new_Jinkela_wire_4099;
    wire new_Jinkela_wire_2946;
    wire new_Jinkela_wire_7927;
    wire new_Jinkela_wire_5512;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_3206;
    wire new_Jinkela_wire_16844;
    wire new_Jinkela_wire_14485;
    wire new_Jinkela_wire_15372;
    wire new_Jinkela_wire_5133;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_21183;
    wire new_Jinkela_wire_5351;
    wire new_Jinkela_wire_13234;
    wire new_Jinkela_wire_19524;
    wire new_Jinkela_wire_19870;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_14638;
    wire new_Jinkela_wire_10171;
    wire new_Jinkela_wire_21073;
    wire new_Jinkela_wire_9710;
    wire new_Jinkela_wire_8736;
    wire new_Jinkela_wire_3517;
    wire new_Jinkela_wire_5047;
    wire new_Jinkela_wire_14263;
    wire new_Jinkela_wire_15317;
    wire new_Jinkela_wire_17616;
    wire new_Jinkela_wire_15922;
    wire new_Jinkela_wire_13713;
    wire new_Jinkela_wire_18925;
    wire new_Jinkela_wire_2906;
    wire new_Jinkela_wire_16653;
    wire new_Jinkela_wire_19061;
    wire new_Jinkela_wire_11638;
    wire new_Jinkela_wire_6015;
    wire new_Jinkela_wire_3781;
    wire new_Jinkela_wire_12591;
    wire new_Jinkela_wire_13705;
    wire _0043_;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_11442;
    wire new_Jinkela_wire_14761;
    wire _1022_;
    wire new_Jinkela_wire_12518;
    wire new_Jinkela_wire_13289;
    wire new_Jinkela_wire_19827;
    wire new_Jinkela_wire_4161;
    wire new_Jinkela_wire_9550;
    wire new_Jinkela_wire_8820;
    wire new_Jinkela_wire_16156;
    wire new_Jinkela_wire_3519;
    wire new_Jinkela_wire_2177;
    wire new_Jinkela_wire_8777;
    wire new_Jinkela_wire_14301;
    wire new_Jinkela_wire_11043;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_16455;
    wire new_Jinkela_wire_8100;
    wire new_Jinkela_wire_15946;
    wire new_Jinkela_wire_9293;
    wire new_Jinkela_wire_11202;
    wire new_Jinkela_wire_7287;
    wire new_Jinkela_wire_20972;
    wire new_Jinkela_wire_20344;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_16042;
    wire new_Jinkela_wire_17850;
    wire new_Jinkela_wire_16812;
    wire new_Jinkela_wire_8188;
    wire new_Jinkela_wire_16603;
    wire new_Jinkela_wire_12453;
    wire new_Jinkela_wire_10973;
    wire new_Jinkela_wire_16743;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_20012;
    wire new_Jinkela_wire_7757;
    wire new_Jinkela_wire_9409;
    wire new_Jinkela_wire_13395;
    wire new_Jinkela_wire_17491;
    wire new_Jinkela_wire_20577;
    wire new_Jinkela_wire_14740;
    wire new_Jinkela_wire_4843;
    wire new_Jinkela_wire_13996;
    wire new_Jinkela_wire_9962;
    wire new_Jinkela_wire_19880;
    wire new_Jinkela_wire_2106;
    wire new_Jinkela_wire_9271;
    wire new_Jinkela_wire_21138;
    wire _0232_;
    wire new_Jinkela_wire_20937;
    wire new_Jinkela_wire_19704;
    wire new_Jinkela_wire_19303;
    wire new_Jinkela_wire_10577;
    wire new_Jinkela_wire_12035;
    wire new_Jinkela_wire_17211;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_8024;
    wire new_Jinkela_wire_20487;
    wire new_Jinkela_wire_8298;
    wire new_Jinkela_wire_4802;
    wire new_Jinkela_wire_7898;
    wire new_Jinkela_wire_20400;
    wire new_Jinkela_wire_16568;
    wire new_Jinkela_wire_21230;
    wire _0554_;
    wire _1260_;
    wire new_Jinkela_wire_17747;
    wire new_Jinkela_wire_2134;
    wire new_Jinkela_wire_2899;
    wire new_Jinkela_wire_17511;
    wire new_Jinkela_wire_9244;
    wire new_Jinkela_wire_19010;
    wire new_Jinkela_wire_16382;
    wire new_Jinkela_wire_4335;
    wire new_Jinkela_wire_6699;
    wire new_Jinkela_wire_7760;
    wire new_Jinkela_wire_11218;
    wire new_Jinkela_wire_14923;
    wire new_Jinkela_wire_18573;
    wire new_Jinkela_wire_3771;
    wire new_Jinkela_wire_15762;
    wire new_Jinkela_wire_12893;
    wire new_Jinkela_wire_5589;
    wire new_Jinkela_wire_4241;
    wire new_Jinkela_wire_14265;
    wire new_Jinkela_wire_18733;
    wire new_Jinkela_wire_16219;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_11057;
    wire new_Jinkela_wire_5674;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_11685;
    wire new_Jinkela_wire_18290;
    wire new_Jinkela_wire_10629;
    wire new_Jinkela_wire_4455;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_7159;
    wire new_Jinkela_wire_18574;
    wire new_Jinkela_wire_18653;
    wire new_Jinkela_wire_2900;
    wire new_Jinkela_wire_13397;
    wire new_Jinkela_wire_8576;
    wire _1695_;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_17515;
    wire new_Jinkela_wire_4383;
    wire new_Jinkela_wire_17299;
    wire new_Jinkela_wire_4055;
    wire new_Jinkela_wire_8111;
    wire _1515_;
    wire new_Jinkela_wire_19533;
    wire new_Jinkela_wire_18336;
    wire new_Jinkela_wire_15241;
    wire new_Jinkela_wire_20723;
    wire new_Jinkela_wire_17580;
    wire new_Jinkela_wire_10308;
    wire new_Jinkela_wire_8520;
    wire new_Jinkela_wire_10338;
    wire _0513_;
    wire new_Jinkela_wire_11574;
    wire new_Jinkela_wire_20085;
    wire new_Jinkela_wire_12427;
    wire new_Jinkela_wire_4135;
    wire new_Jinkela_wire_13639;
    wire new_Jinkela_wire_3904;
    wire new_Jinkela_wire_20788;
    wire new_Jinkela_wire_7134;
    wire new_Jinkela_wire_11813;
    wire _0269_;
    wire new_Jinkela_wire_12454;
    wire new_Jinkela_wire_19334;
    wire new_Jinkela_wire_9929;
    wire new_Jinkela_wire_6265;
    wire new_Jinkela_wire_15412;
    wire new_Jinkela_wire_15830;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_14232;
    wire new_Jinkela_wire_15303;
    wire new_Jinkela_wire_7565;
    wire new_Jinkela_wire_14325;
    wire _0729_;
    wire new_Jinkela_wire_4419;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_19414;
    wire new_Jinkela_wire_3528;
    wire new_Jinkela_wire_4421;
    wire _0426_;
    wire new_Jinkela_wire_15096;
    wire new_Jinkela_wire_20072;
    wire new_Jinkela_wire_17981;
    wire new_Jinkela_wire_5638;
    wire new_Jinkela_wire_12413;
    wire new_Jinkela_wire_4001;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_11733;
    wire new_Jinkela_wire_3713;
    wire new_Jinkela_wire_2221;
    wire new_Jinkela_wire_3174;
    wire new_Jinkela_wire_15005;
    wire new_Jinkela_wire_2318;
    wire new_Jinkela_wire_15330;
    wire new_Jinkela_wire_8619;
    wire new_Jinkela_wire_8368;
    wire new_Jinkela_wire_6031;
    wire new_Jinkela_wire_8362;
    wire new_Jinkela_wire_15603;
    wire new_Jinkela_wire_9877;
    wire new_Jinkela_wire_18081;
    wire new_Jinkela_wire_19046;
    wire new_Jinkela_wire_13697;
    wire new_Jinkela_wire_8009;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_19747;
    wire new_Jinkela_wire_20580;
    wire new_Jinkela_wire_12011;
    wire new_Jinkela_wire_14620;
    wire new_Jinkela_wire_12926;
    wire new_Jinkela_wire_1869;
    wire new_Jinkela_wire_9869;
    wire new_Jinkela_wire_21099;
    wire new_Jinkela_wire_20370;
    wire new_Jinkela_wire_1315;
    wire new_Jinkela_wire_15395;
    wire new_Jinkela_wire_11138;
    wire new_Jinkela_wire_8510;
    wire new_Jinkela_wire_2710;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_3217;
    wire new_Jinkela_wire_12819;
    wire new_Jinkela_wire_12648;
    wire new_Jinkela_wire_8525;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_13183;
    wire new_Jinkela_wire_21191;
    wire new_Jinkela_wire_6210;
    wire new_Jinkela_wire_10855;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_9668;
    wire new_Jinkela_wire_15727;
    wire new_Jinkela_wire_15438;
    wire new_Jinkela_wire_7921;
    wire new_Jinkela_wire_15808;
    wire new_Jinkela_wire_19141;
    wire new_Jinkela_wire_21043;
    wire new_Jinkela_wire_21226;
    wire new_Jinkela_wire_4070;
    wire new_Jinkela_wire_19510;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_14792;
    wire new_Jinkela_wire_21279;
    wire new_Jinkela_wire_13278;
    wire new_Jinkela_wire_17666;
    wire new_Jinkela_wire_20176;
    wire new_Jinkela_wire_19305;
    wire new_Jinkela_wire_16642;
    wire new_Jinkela_wire_8136;
    wire new_Jinkela_wire_17667;
    wire new_Jinkela_wire_12603;
    wire new_Jinkela_wire_1846;
    wire new_Jinkela_wire_14623;
    wire new_Jinkela_wire_13881;
    wire new_Jinkela_wire_16341;
    wire new_Jinkela_wire_20465;
    wire new_Jinkela_wire_6199;
    wire new_Jinkela_wire_18468;
    wire new_Jinkela_wire_7364;
    wire new_Jinkela_wire_9336;
    wire new_Jinkela_wire_11416;
    wire new_Jinkela_wire_16114;
    wire new_Jinkela_wire_5394;
    wire new_Jinkela_wire_5319;
    wire new_Jinkela_wire_11100;
    wire new_Jinkela_wire_19483;
    wire new_Jinkela_wire_245;
    wire _0473_;
    wire new_Jinkela_wire_13989;
    wire _1448_;
    wire new_Jinkela_wire_13527;
    wire new_Jinkela_wire_19371;
    wire new_Jinkela_wire_15796;
    wire new_Jinkela_wire_11730;
    wire _0118_;
    wire new_Jinkela_wire_15658;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_7884;
    wire new_Jinkela_wire_3334;
    wire new_Jinkela_wire_11103;
    wire new_Jinkela_wire_3428;
    wire new_Jinkela_wire_13980;
    wire new_Jinkela_wire_18164;
    wire new_Jinkela_wire_4981;
    wire new_Jinkela_wire_18886;
    wire new_Jinkela_wire_10941;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_5727;
    wire new_Jinkela_wire_14602;
    wire new_Jinkela_wire_19811;
    wire new_Jinkela_wire_3078;
    wire new_Jinkela_wire_3221;
    wire new_Jinkela_wire_20240;
    wire new_Jinkela_wire_3187;
    wire new_Jinkela_wire_9553;
    wire new_Jinkela_wire_2406;
    wire new_Jinkela_wire_5708;
    wire new_Jinkela_wire_17871;
    wire new_Jinkela_wire_5799;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_2659;
    wire _1236_;
    wire _0829_;
    wire new_Jinkela_wire_5110;
    wire new_Jinkela_wire_9736;
    wire new_Jinkela_wire_13913;
    wire new_Jinkela_wire_4559;
    wire new_Jinkela_wire_7873;
    wire new_Jinkela_wire_2302;
    wire new_Jinkela_wire_16701;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_2093;
    wire new_Jinkela_wire_12457;
    wire new_Jinkela_wire_2596;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_14169;
    wire new_Jinkela_wire_3045;
    wire new_Jinkela_wire_7193;
    wire new_Jinkela_wire_3844;
    wire _1306_;
    wire _0380_;
    wire new_Jinkela_wire_20844;
    wire new_Jinkela_wire_8324;
    wire new_Jinkela_wire_19884;
    wire new_Jinkela_wire_12107;
    wire new_Jinkela_wire_14319;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_9171;
    wire new_Jinkela_wire_18012;
    wire new_Jinkela_wire_9424;
    wire new_Jinkela_wire_18501;
    wire _0435_;
    wire new_Jinkela_wire_11559;
    wire new_Jinkela_wire_11463;
    wire new_Jinkela_wire_12057;
    wire new_Jinkela_wire_17250;
    wire new_Jinkela_wire_2783;
    wire new_Jinkela_wire_6857;
    wire new_Jinkela_wire_6235;
    wire new_Jinkela_wire_5207;
    wire new_Jinkela_wire_9011;
    wire new_Jinkela_wire_13073;
    wire _0918_;
    wire new_Jinkela_wire_2987;
    wire new_Jinkela_wire_13621;
    wire new_Jinkela_wire_1773;
    wire new_Jinkela_wire_15329;
    wire new_Jinkela_wire_19175;
    wire new_Jinkela_wire_6076;
    wire new_Jinkela_wire_18089;
    wire new_Jinkela_wire_9448;
    wire new_Jinkela_wire_14330;
    wire _0033_;
    wire new_Jinkela_wire_15451;
    wire new_Jinkela_wire_10724;
    wire new_Jinkela_wire_12436;
    wire new_Jinkela_wire_14094;
    wire new_Jinkela_wire_5765;
    wire new_Jinkela_wire_14149;
    wire new_Jinkela_wire_14702;
    wire new_Jinkela_wire_6217;
    wire new_Jinkela_wire_3914;
    wire new_Jinkela_wire_15814;
    wire new_Jinkela_wire_1285;
    wire _0774_;
    wire new_Jinkela_wire_9582;
    wire new_Jinkela_wire_3677;
    wire new_Jinkela_wire_19819;
    wire new_Jinkela_wire_8490;
    wire new_Jinkela_wire_15211;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_13468;
    wire new_Jinkela_wire_2722;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_7958;
    wire new_Jinkela_wire_11792;
    wire new_Jinkela_wire_8959;
    wire new_Jinkela_wire_10461;
    wire new_Jinkela_wire_9458;
    wire new_Jinkela_wire_5967;
    wire new_Jinkela_wire_8828;
    wire new_Jinkela_wire_16663;
    wire new_Jinkela_wire_7639;
    wire new_Jinkela_wire_19495;
    wire new_Jinkela_wire_7447;
    wire new_Jinkela_wire_7100;
    wire new_Jinkela_wire_7532;
    wire new_Jinkela_wire_15074;
    wire new_Jinkela_wire_12577;
    wire new_Jinkela_wire_5919;
    wire new_Jinkela_wire_9926;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_8914;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_12322;
    wire new_Jinkela_wire_19401;
    wire new_Jinkela_wire_15836;
    wire new_Jinkela_wire_2809;
    wire new_Jinkela_wire_16775;
    wire new_Jinkela_wire_13486;
    wire new_Jinkela_wire_20071;
    wire new_Jinkela_wire_3348;
    wire new_Jinkela_wire_18394;
    wire _0619_;
    wire new_Jinkela_wire_9823;
    wire new_Jinkela_wire_13530;
    wire new_Jinkela_wire_5038;
    wire new_Jinkela_wire_8205;
    wire new_Jinkela_wire_2061;
    wire new_Jinkela_wire_2887;
    wire new_Jinkela_wire_12681;
    wire new_Jinkela_wire_15635;
    wire new_Jinkela_wire_4107;
    wire new_Jinkela_wire_13338;
    wire new_Jinkela_wire_13207;
    wire new_Jinkela_wire_20913;
    wire new_Jinkela_wire_3500;
    wire new_Jinkela_wire_17576;
    wire new_Jinkela_wire_5096;
    wire new_Jinkela_wire_16510;
    wire new_Jinkela_wire_14589;
    wire new_Jinkela_wire_5675;
    wire new_Jinkela_wire_5330;
    wire new_Jinkela_wire_2049;
    wire new_Jinkela_wire_9686;
    wire new_Jinkela_wire_20405;
    wire new_Jinkela_wire_3558;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_21042;
    wire new_Jinkela_wire_11405;
    wire _0328_;
    wire new_Jinkela_wire_6035;
    wire _0959_;
    wire new_Jinkela_wire_14823;
    wire new_Jinkela_wire_16325;
    wire new_Jinkela_wire_21084;
    wire new_Jinkela_wire_3661;
    wire _0160_;
    wire new_Jinkela_wire_10659;
    wire new_Jinkela_wire_9265;
    wire new_Jinkela_wire_13254;
    wire new_Jinkela_wire_9658;
    wire new_Jinkela_wire_11451;
    wire new_Jinkela_wire_10919;
    wire new_Jinkela_wire_11849;
    wire new_Jinkela_wire_9106;
    wire new_Jinkela_wire_9115;
    wire new_Jinkela_wire_8140;
    wire new_Jinkela_wire_11131;
    wire new_Jinkela_wire_10923;
    wire new_Jinkela_wire_13791;
    wire new_Jinkela_wire_16475;
    wire new_Jinkela_wire_3074;
    wire new_Jinkela_wire_15733;
    wire new_Jinkela_wire_2832;
    wire new_Jinkela_wire_10032;
    wire new_Jinkela_wire_10242;
    wire _1036_;
    wire new_Jinkela_wire_8405;
    wire new_Jinkela_wire_7974;
    wire new_Jinkela_wire_4471;
    wire new_Jinkela_wire_10178;
    wire new_Jinkela_wire_14231;
    wire new_Jinkela_wire_8549;
    wire new_Jinkela_wire_2162;
    wire new_Jinkela_wire_15059;
    wire new_Jinkela_wire_5175;
    wire new_Jinkela_wire_18597;
    wire new_Jinkela_wire_19019;
    wire new_Jinkela_wire_15918;
    wire new_Jinkela_wire_20720;
    wire new_Jinkela_wire_11790;
    wire new_Jinkela_wire_9669;
    wire new_Jinkela_wire_3542;
    wire new_Jinkela_wire_9579;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_4667;
    wire new_Jinkela_wire_4258;
    wire new_Jinkela_wire_14692;
    wire new_Jinkela_wire_9126;
    wire new_Jinkela_wire_11921;
    wire new_Jinkela_wire_7522;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_12523;
    wire _0589_;
    wire new_Jinkela_wire_11708;
    wire new_Jinkela_wire_12734;
    wire new_Jinkela_wire_20639;
    wire new_Jinkela_wire_12709;
    wire new_Jinkela_wire_11755;
    wire new_Jinkela_wire_11047;
    wire new_Jinkela_wire_17181;
    wire new_Jinkela_wire_3628;
    wire new_Jinkela_wire_13676;
    wire new_Jinkela_wire_5018;
    wire new_Jinkela_wire_14313;
    wire new_Jinkela_wire_9460;
    wire new_Jinkela_wire_3314;
    wire _1290_;
    wire new_Jinkela_wire_14463;
    wire new_Jinkela_wire_7277;
    wire new_Jinkela_wire_7836;
    wire new_Jinkela_wire_11825;
    wire new_Jinkela_wire_10911;
    wire new_Jinkela_wire_17532;
    wire new_Jinkela_wire_20938;
    wire new_Jinkela_wire_17204;
    wire new_Jinkela_wire_11130;
    wire new_Jinkela_wire_19963;
    wire new_Jinkela_wire_4058;
    wire new_Jinkela_wire_16122;
    wire new_Jinkela_wire_4549;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_16123;
    wire new_Jinkela_wire_6858;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_11741;
    wire new_Jinkela_wire_11693;
    wire new_Jinkela_wire_16190;
    wire _0608_;
    wire new_Jinkela_wire_2790;
    wire _1125_;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_5878;
    wire new_Jinkela_wire_21053;
    wire new_Jinkela_wire_5191;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_20337;
    wire new_Jinkela_wire_16476;
    wire new_Jinkela_wire_9829;
    wire new_Jinkela_wire_18933;
    wire new_Jinkela_wire_6318;
    wire new_Jinkela_wire_16473;
    wire new_Jinkela_wire_6026;
    wire _0260_;
    wire new_Jinkela_wire_6505;
    wire new_Jinkela_wire_7302;
    wire new_Jinkela_wire_2129;
    wire new_Jinkela_wire_16904;
    wire new_Jinkela_wire_11183;
    wire new_Jinkela_wire_16695;
    wire new_Jinkela_wire_16366;
    wire _0459_;
    wire new_Jinkela_wire_18204;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_5452;
    wire _0252_;
    wire new_Jinkela_wire_5061;
    wire _0110_;
    wire _1123_;
    wire new_Jinkela_wire_16513;
    wire new_Jinkela_wire_18192;
    wire new_Jinkela_wire_1570;
    wire _1253_;
    wire new_Jinkela_wire_3391;
    wire new_Jinkela_wire_5946;
    wire _0983_;
    wire new_Jinkela_wire_16907;
    wire new_Jinkela_wire_14145;
    wire new_Jinkela_wire_19838;
    wire new_Jinkela_wire_9906;
    wire new_Jinkela_wire_14528;
    wire new_Jinkela_wire_5196;
    wire _0960_;
    wire new_Jinkela_wire_19496;
    wire new_Jinkela_wire_15838;
    wire new_Jinkela_wire_12081;
    wire new_Jinkela_wire_18167;
    wire new_Jinkela_wire_3674;
    wire new_Jinkela_wire_12557;
    wire new_Jinkela_wire_8572;
    wire new_Jinkela_wire_7689;
    wire new_Jinkela_wire_8186;
    wire new_Jinkela_wire_10192;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_2091;
    wire new_Jinkela_wire_16967;
    wire new_Jinkela_wire_10914;
    wire new_Jinkela_wire_16737;
    wire new_Jinkela_wire_20079;
    wire new_Jinkela_wire_2787;
    wire new_Jinkela_wire_10508;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_17220;
    wire new_Jinkela_wire_4749;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_12960;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_10936;
    wire new_Jinkela_wire_7595;
    wire new_Jinkela_wire_9023;
    wire new_Jinkela_wire_6307;
    wire new_Jinkela_wire_3487;
    wire new_Jinkela_wire_3132;
    wire _0788_;
    wire new_Jinkela_wire_2925;
    wire new_Jinkela_wire_10221;
    wire new_Jinkela_wire_17280;
    wire new_Jinkela_wire_8255;
    wire new_Jinkela_wire_17550;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_10608;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_20119;
    wire new_Jinkela_wire_5985;
    wire new_Jinkela_wire_15284;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_9592;
    wire new_Jinkela_wire_19057;
    wire new_Jinkela_wire_17954;
    wire new_Jinkela_wire_7155;
    wire new_Jinkela_wire_1751;
    wire new_Jinkela_wire_21063;
    wire new_Jinkela_wire_14364;
    wire new_Jinkela_wire_2195;
    wire new_Jinkela_wire_10653;
    wire new_Jinkela_wire_7575;
    wire new_Jinkela_wire_16620;
    wire new_Jinkela_wire_9913;
    wire new_Jinkela_wire_12168;
    wire new_Jinkela_wire_3273;
    wire new_Jinkela_wire_18274;
    wire new_Jinkela_wire_19511;
    wire new_Jinkela_wire_19229;
    wire new_Jinkela_wire_2772;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_21021;
    wire new_Jinkela_wire_4232;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_16048;
    wire new_Jinkela_wire_5454;
    wire new_Jinkela_wire_10189;
    wire new_Jinkela_wire_8949;
    wire new_Jinkela_wire_20384;
    wire new_Jinkela_wire_8301;
    wire new_Jinkela_wire_4938;
    wire new_Jinkela_wire_2796;
    wire new_Jinkela_wire_19044;
    wire new_Jinkela_wire_3212;
    wire new_Jinkela_wire_5134;
    wire new_Jinkela_wire_20691;
    wire _0722_;
    wire new_Jinkela_wire_19441;
    wire new_Jinkela_wire_14070;
    wire new_Jinkela_wire_20875;
    wire _0574_;
    wire new_Jinkela_wire_13796;
    wire new_Jinkela_wire_19237;
    wire new_Jinkela_wire_15537;
    wire _0102_;
    wire new_Jinkela_wire_21166;
    wire new_Jinkela_wire_6654;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_10429;
    wire new_Jinkela_wire_15103;
    wire new_Jinkela_wire_9389;
    wire new_Jinkela_wire_9181;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_20129;
    wire new_Jinkela_wire_7224;
    wire new_Jinkela_wire_17243;
    wire new_Jinkela_wire_4279;
    wire new_Jinkela_wire_11692;
    wire new_Jinkela_wire_19023;
    wire new_Jinkela_wire_18211;
    wire new_Jinkela_wire_7635;
    wire new_Jinkela_wire_17145;
    wire new_Jinkela_wire_2940;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_5273;
    wire new_Jinkela_wire_10733;
    wire new_Jinkela_wire_10451;
    wire new_Jinkela_wire_15031;
    wire _0239_;
    wire new_Jinkela_wire_9996;
    wire new_Jinkela_wire_19405;
    wire new_Jinkela_wire_17401;
    wire _0993_;
    wire new_Jinkela_wire_3961;
    wire new_Jinkela_wire_19139;
    wire new_Jinkela_wire_3057;
    wire new_Jinkela_wire_21294;
    wire new_Jinkela_wire_19736;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_14492;
    wire new_Jinkela_wire_2528;
    wire new_Jinkela_wire_14133;
    wire new_Jinkela_wire_18676;
    wire new_Jinkela_wire_19770;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_5585;
    wire new_Jinkela_wire_17234;
    wire new_Jinkela_wire_19658;
    wire new_Jinkela_wire_16864;
    wire new_Jinkela_wire_10969;
    wire new_Jinkela_wire_13297;
    wire new_Jinkela_wire_20433;
    wire new_Jinkela_wire_15909;
    wire new_Jinkela_wire_5712;
    wire new_Jinkela_wire_19214;
    wire new_Jinkela_wire_12027;
    wire new_Jinkela_wire_11645;
    wire new_Jinkela_wire_14945;
    wire new_Jinkela_wire_1942;
    wire new_Jinkela_wire_20393;
    wire _1567_;
    wire _1169_;
    wire new_Jinkela_wire_10750;
    wire _0696_;
    wire new_Jinkela_wire_3191;
    wire new_Jinkela_wire_12365;
    wire new_Jinkela_wire_8912;
    wire new_Jinkela_wire_19917;
    wire new_Jinkela_wire_19935;
    wire new_Jinkela_wire_13088;
    wire new_Jinkela_wire_16833;
    wire new_Jinkela_wire_19791;
    wire _1184_;
    wire new_Jinkela_wire_16433;
    wire new_Jinkela_wire_2070;
    wire new_Jinkela_wire_17253;
    wire new_Jinkela_wire_15886;
    wire new_Jinkela_wire_9191;
    wire new_Jinkela_wire_20915;
    wire new_Jinkela_wire_9872;
    wire new_Jinkela_wire_14081;
    wire new_Jinkela_wire_9899;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_3121;
    wire new_Jinkela_wire_9803;
    wire new_Jinkela_wire_19833;
    wire new_Jinkela_wire_9455;
    wire new_Jinkela_wire_15217;
    wire _1613_;
    wire new_Jinkela_wire_18817;
    wire new_Jinkela_wire_3155;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_11204;
    wire new_Jinkela_wire_7560;
    wire new_Jinkela_wire_8780;
    wire new_Jinkela_wire_16377;
    wire new_Jinkela_wire_18553;
    wire new_Jinkela_wire_20780;
    wire _0641_;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_8845;
    wire new_Jinkela_wire_8668;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_10831;
    wire new_Jinkela_wire_9941;
    wire new_Jinkela_wire_11642;
    wire new_Jinkela_wire_7646;
    wire new_Jinkela_wire_15109;
    wire new_Jinkela_wire_14897;
    wire new_Jinkela_wire_6954;
    wire new_Jinkela_wire_12230;
    wire new_Jinkela_wire_9985;
    wire new_Jinkela_wire_20622;
    wire new_Jinkela_wire_16735;
    wire new_Jinkela_wire_6762;
    wire new_Jinkela_wire_2653;
    wire new_Jinkela_wire_4287;
    wire new_Jinkela_wire_11585;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_15406;
    wire new_Jinkela_wire_6683;
    wire new_Jinkela_wire_9394;
    wire new_Jinkela_wire_4556;
    wire new_Jinkela_wire_14649;
    wire new_Jinkela_wire_8522;
    wire new_Jinkela_wire_12767;
    wire new_Jinkela_wire_5506;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_7538;
    wire new_Jinkela_wire_2818;
    wire new_Jinkela_wire_15127;
    wire new_Jinkela_wire_7694;
    wire new_Jinkela_wire_3760;
    wire new_Jinkela_wire_4242;
    wire new_Jinkela_wire_5665;
    wire new_Jinkela_wire_2438;
    wire new_Jinkela_wire_9694;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_13305;
    wire new_Jinkela_wire_2774;
    wire new_Jinkela_wire_6750;
    wire new_Jinkela_wire_18049;
    wire new_Jinkela_wire_18410;
    wire new_Jinkela_wire_18654;
    wire new_Jinkela_wire_12980;
    wire _0374_;
    wire new_Jinkela_wire_18562;
    wire new_Jinkela_wire_13599;
    wire new_Jinkela_wire_15768;
    wire new_Jinkela_wire_20903;
    wire new_Jinkela_wire_8365;
    wire new_Jinkela_wire_14690;
    wire new_Jinkela_wire_15512;
    wire new_Jinkela_wire_18913;
    wire new_Jinkela_wire_7267;
    wire new_Jinkela_wire_12671;
    wire new_Jinkela_wire_4962;
    wire new_Jinkela_wire_15309;
    wire new_Jinkela_wire_16346;
    wire new_Jinkela_wire_15077;
    wire new_Jinkela_wire_9277;
    wire new_Jinkela_wire_9551;
    wire new_Jinkela_wire_6410;
    wire new_Jinkela_wire_11434;
    wire new_Jinkela_wire_6554;
    wire new_Jinkela_wire_7903;
    wire new_Jinkela_wire_14191;
    wire new_Jinkela_wire_2549;
    wire new_Jinkela_wire_6434;
    wire new_Jinkela_wire_7611;
    wire new_Jinkela_wire_5579;
    wire new_Jinkela_wire_6312;
    wire new_Jinkela_wire_17715;
    wire new_Jinkela_wire_14902;
    wire new_Jinkela_wire_1775;
    wire new_Jinkela_wire_17820;
    wire new_Jinkela_wire_12791;
    wire _0096_;
    wire new_Jinkela_wire_21296;
    wire new_Jinkela_wire_14704;
    wire new_Jinkela_wire_10404;
    wire new_Jinkela_wire_8057;
    wire _1674_;
    wire new_Jinkela_wire_20443;
    wire new_Jinkela_wire_8975;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_15431;
    wire new_Jinkela_wire_16035;
    wire new_Jinkela_wire_9243;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_7395;
    wire new_Jinkela_wire_3778;
    wire new_Jinkela_wire_10770;
    wire new_Jinkela_wire_8606;
    wire new_Jinkela_wire_16185;
    wire new_Jinkela_wire_2005;
    wire new_Jinkela_wire_20261;
    wire new_Jinkela_wire_10309;
    wire new_Jinkela_wire_4038;
    wire new_Jinkela_wire_15272;
    wire new_Jinkela_wire_21301;
    wire _1211_;
    wire new_Jinkela_wire_17524;
    wire new_Jinkela_wire_7339;
    wire new_Jinkela_wire_20266;
    wire new_Jinkela_wire_16889;
    wire new_Jinkela_wire_8796;
    wire new_Jinkela_wire_6016;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_19594;
    wire _1114_;
    wire new_Jinkela_wire_8755;
    wire new_Jinkela_wire_19893;
    wire new_Jinkela_wire_18433;
    wire new_Jinkela_wire_18884;
    wire new_Jinkela_wire_1892;
    wire new_Jinkela_wire_20906;
    wire new_Jinkela_wire_4227;
    wire _1259_;
    wire new_Jinkela_wire_19343;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_8098;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_4673;
    wire new_Jinkela_wire_20173;
    wire new_Jinkela_wire_11469;
    wire new_Jinkela_wire_2259;
    wire new_Jinkela_wire_9352;
    wire new_Jinkela_wire_17353;
    wire new_Jinkela_wire_4886;
    wire new_Jinkela_wire_14022;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_8416;
    wire new_Jinkela_wire_19116;
    wire new_Jinkela_wire_14998;
    wire _0744_;
    wire new_Jinkela_wire_6480;
    wire new_Jinkela_wire_4638;
    wire new_Jinkela_wire_6665;
    wire new_Jinkela_wire_9087;
    wire new_Jinkela_wire_12031;
    wire new_Jinkela_wire_7420;
    wire new_Jinkela_wire_19429;
    wire new_Jinkela_wire_12534;
    wire new_Jinkela_wire_9276;
    wire new_Jinkela_wire_5710;
    wire new_Jinkela_wire_17163;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_20890;
    wire new_Jinkela_wire_4832;
    wire new_Jinkela_wire_15508;
    wire new_Jinkela_wire_20387;
    wire new_Jinkela_wire_3832;
    wire new_Jinkela_wire_2493;
    wire new_Jinkela_wire_12684;
    wire new_Jinkela_wire_12638;
    wire _1474_;
    wire new_Jinkela_wire_11422;
    wire new_Jinkela_wire_9708;
    wire new_Jinkela_wire_10105;
    wire new_Jinkela_wire_6346;
    wire new_Jinkela_wire_17905;
    wire new_Jinkela_wire_20911;
    wire new_Jinkela_wire_4758;
    wire new_Jinkela_wire_13476;
    wire new_Jinkela_wire_3189;
    wire new_Jinkela_wire_18815;
    wire new_Jinkela_wire_12743;
    wire new_Jinkela_wire_16892;
    wire new_Jinkela_wire_14490;
    wire new_Jinkela_wire_20932;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_13572;
    wire new_Jinkela_wire_7785;
    wire _0939_;
    wire new_Jinkela_wire_5470;
    wire new_Jinkela_wire_4250;
    wire new_Jinkela_wire_4458;
    wire new_Jinkela_wire_5205;
    wire new_Jinkela_wire_4836;
    wire new_Jinkela_wire_7814;
    wire new_Jinkela_wire_19984;
    wire new_Jinkela_wire_13306;
    wire new_Jinkela_wire_8933;
    wire new_Jinkela_wire_20374;
    wire new_Jinkela_wire_15977;
    wire new_Jinkela_wire_13717;
    wire new_Jinkela_wire_19570;
    wire new_Jinkela_wire_6024;
    wire new_Jinkela_wire_19301;
    wire new_Jinkela_wire_13964;
    wire new_Jinkela_wire_19913;
    wire new_Jinkela_wire_2694;
    wire new_Jinkela_wire_6552;
    wire new_Jinkela_wire_18802;
    wire new_Jinkela_wire_14892;
    wire new_Jinkela_wire_16300;
    wire new_Jinkela_wire_15204;
    wire _0810_;
    wire new_Jinkela_wire_14402;
    wire _0931_;
    wire new_Jinkela_wire_10087;
    wire new_Jinkela_wire_10246;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_2598;
    wire new_Jinkela_wire_13665;
    wire new_Jinkela_wire_17737;
    wire _0433_;
    wire new_Jinkela_wire_17661;
    wire new_Jinkela_wire_12431;
    wire new_Jinkela_wire_17672;
    wire new_Jinkela_wire_4349;
    wire new_Jinkela_wire_18338;
    wire new_Jinkela_wire_17739;
    wire new_Jinkela_wire_13368;
    wire new_Jinkela_wire_18294;
    wire new_Jinkela_wire_15389;
    wire new_Jinkela_wire_2889;
    wire new_Jinkela_wire_16353;
    wire new_Jinkela_wire_19096;
    wire new_Jinkela_wire_6000;
    wire new_Jinkela_wire_19351;
    wire new_Jinkela_wire_20710;
    wire new_Jinkela_wire_8160;
    wire new_Jinkela_wire_12491;
    wire new_Jinkela_wire_9599;
    wire new_Jinkela_wire_5353;
    wire new_Jinkela_wire_19930;
    wire new_Jinkela_wire_3624;
    wire new_Jinkela_wire_1765;
    wire _1564_;
    wire _1496_;
    wire new_Jinkela_wire_19600;
    wire new_Jinkela_wire_2815;
    wire new_Jinkela_wire_18669;
    wire new_Jinkela_wire_10065;
    wire new_Jinkela_wire_9725;
    wire _0884_;
    wire new_Jinkela_wire_17062;
    wire new_Jinkela_wire_19290;
    wire new_Jinkela_wire_9215;
    wire new_Jinkela_wire_6927;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_15563;
    wire new_Jinkela_wire_3013;
    wire new_Jinkela_wire_8981;
    wire new_Jinkela_wire_5425;
    wire new_Jinkela_wire_20043;
    wire new_Jinkela_wire_7613;
    wire new_Jinkela_wire_13772;
    wire new_Jinkela_wire_8040;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_19459;
    wire new_Jinkela_wire_6335;
    wire new_Jinkela_wire_17659;
    wire new_Jinkela_wire_4104;
    wire new_Jinkela_wire_6613;
    wire new_Jinkela_wire_1955;
    wire new_Jinkela_wire_15349;
    wire new_Jinkela_wire_12412;
    wire new_Jinkela_wire_16057;
    wire new_Jinkela_wire_17270;
    wire new_Jinkela_wire_3022;
    wire new_Jinkela_wire_1360;
    wire _0277_;
    wire _1637_;
    wire new_Jinkela_wire_16480;
    wire new_Jinkela_wire_6329;
    wire new_Jinkela_wire_5049;
    wire _1248_;
    wire new_Jinkela_wire_8505;
    wire new_Jinkela_wire_12394;
    wire new_Jinkela_wire_20650;
    wire new_Jinkela_wire_10728;
    wire new_Jinkela_wire_5317;
    wire new_Jinkela_wire_6126;
    wire new_Jinkela_wire_7041;
    wire new_Jinkela_wire_19383;
    wire _0468_;
    wire new_Jinkela_wire_13072;
    wire new_Jinkela_wire_18885;
    wire new_Jinkela_wire_2873;
    wire _0452_;
    wire new_Jinkela_wire_13966;
    wire new_Jinkela_wire_9400;
    wire new_Jinkela_wire_12613;
    wire new_Jinkela_wire_15955;
    wire _1039_;
    wire _1093_;
    wire new_Jinkela_wire_14349;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_8195;
    wire new_Jinkela_wire_9479;
    wire new_Jinkela_wire_12717;
    wire new_Jinkela_wire_11636;
    wire new_Jinkela_wire_6128;
    wire new_Jinkela_wire_10943;
    wire new_Jinkela_wire_5503;
    wire new_Jinkela_wire_16964;
    wire new_Jinkela_wire_21023;
    wire new_Jinkela_wire_10175;
    wire _1238_;
    wire new_Jinkela_wire_5744;
    wire new_Jinkela_wire_8214;
    wire new_Jinkela_wire_20587;
    wire new_Jinkela_wire_18457;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_8182;
    wire new_Jinkela_wire_21134;
    wire new_Jinkela_wire_19976;
    wire new_Jinkela_wire_3698;
    wire new_Jinkela_wire_6387;
    wire new_Jinkela_wire_11595;
    wire new_Jinkela_wire_14438;
    wire new_Jinkela_wire_11841;
    wire new_Jinkela_wire_15006;
    wire new_Jinkela_wire_13236;
    wire _0457_;
    wire new_Jinkela_wire_9888;
    wire new_Jinkela_wire_17779;
    wire _0565_;
    wire new_Jinkela_wire_7980;
    wire new_Jinkela_wire_4666;
    wire new_Jinkela_wire_14827;
    wire new_Jinkela_wire_20533;
    wire new_Jinkela_wire_8435;
    wire new_Jinkela_wire_13983;
    wire new_Jinkela_wire_9492;
    wire new_Jinkela_wire_10070;
    wire new_Jinkela_wire_13571;
    wire new_Jinkela_wire_18257;
    wire new_Jinkela_wire_11589;
    wire new_Jinkela_wire_6338;
    wire _1181_;
    wire new_Jinkela_wire_9348;
    wire new_Jinkela_wire_7860;
    wire new_Jinkela_wire_12711;
    wire new_Jinkela_wire_11918;
    wire new_Jinkela_wire_15763;
    wire new_Jinkela_wire_6344;
    wire new_Jinkela_wire_10295;
    wire new_Jinkela_wire_13804;
    wire new_Jinkela_wire_20329;
    wire _0877_;
    wire new_Jinkela_wire_17641;
    wire new_Jinkela_wire_6959;
    wire new_Jinkela_wire_11875;
    wire new_Jinkela_wire_18865;
    wire new_Jinkela_wire_15195;
    wire new_Jinkela_wire_12194;
    wire new_Jinkela_wire_4079;
    wire new_Jinkela_wire_17452;
    wire new_Jinkela_wire_12970;
    wire new_Jinkela_wire_3676;
    wire new_Jinkela_wire_18212;
    wire new_Jinkela_wire_9376;
    wire new_Jinkela_wire_11973;
    wire new_Jinkela_wire_8245;
    wire new_Jinkela_wire_15010;
    wire new_Jinkela_wire_8201;
    wire new_Jinkela_wire_2182;
    wire new_Jinkela_wire_14871;
    wire new_Jinkela_wire_1792;
    wire new_Jinkela_wire_7062;
    wire new_Jinkela_wire_17439;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_5924;
    wire new_Jinkela_wire_11584;
    wire new_Jinkela_wire_12320;
    wire _0977_;
    wire new_Jinkela_wire_11855;
    wire new_Jinkela_wire_14611;
    wire new_Jinkela_wire_18158;
    wire new_Jinkela_wire_11227;
    wire new_Jinkela_wire_20120;
    wire new_Jinkela_wire_17081;
    wire new_Jinkela_wire_10704;
    wire new_Jinkela_wire_1567;
    wire new_Jinkela_wire_16095;
    wire new_Jinkela_wire_17624;
    wire new_Jinkela_wire_15095;
    wire new_Jinkela_wire_10765;
    wire new_Jinkela_wire_12084;
    wire new_Jinkela_wire_6934;
    wire _1002_;
    wire _1777_;
    wire new_Jinkela_wire_5008;
    wire new_Jinkela_wire_12558;
    wire new_Jinkela_wire_12173;
    wire new_Jinkela_wire_6079;
    wire new_Jinkela_wire_18368;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_3639;
    wire new_Jinkela_wire_21130;
    wire new_Jinkela_wire_9664;
    wire new_Jinkela_wire_7269;
    wire new_Jinkela_wire_14865;
    wire new_Jinkela_wire_3436;
    wire new_Jinkela_wire_5276;
    wire new_Jinkela_wire_13140;
    wire new_Jinkela_wire_10369;
    wire new_Jinkela_wire_9840;
    wire _0009_;
    wire new_Jinkela_wire_16629;
    wire new_Jinkela_wire_6767;
    wire new_Jinkela_wire_5802;
    wire new_Jinkela_wire_13312;
    wire new_Jinkela_wire_3578;
    wire new_Jinkela_wire_5382;
    wire new_Jinkela_wire_18673;
    wire new_Jinkela_wire_21172;
    wire new_Jinkela_wire_13100;
    wire new_Jinkela_wire_15567;
    wire new_Jinkela_wire_4636;
    wire new_Jinkela_wire_10100;
    wire new_Jinkela_wire_19982;
    wire new_Jinkela_wire_16891;
    wire new_Jinkela_wire_3102;
    wire new_Jinkela_wire_11475;
    wire _0284_;
    wire new_Jinkela_wire_14029;
    wire new_Jinkela_wire_21077;
    wire new_Jinkela_wire_6296;
    wire _1333_;
    wire new_Jinkela_wire_1312;
    wire _1111_;
    wire new_Jinkela_wire_2288;
    wire new_Jinkela_wire_6702;
    wire _0105_;
    wire new_Jinkela_wire_2568;
    wire new_Jinkela_wire_10399;
    wire new_Jinkela_wire_3670;
    wire _0297_;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_13252;
    wire new_Jinkela_wire_11051;
    wire new_Jinkela_wire_10787;
    wire new_Jinkela_wire_13564;
    wire new_Jinkela_wire_3066;
    wire new_Jinkela_wire_10564;
    wire new_Jinkela_wire_6129;
    wire new_Jinkela_wire_14888;
    wire new_Jinkela_wire_11528;
    wire new_Jinkela_wire_12187;
    wire new_Jinkela_wire_10881;
    wire new_Jinkela_wire_15170;
    wire new_Jinkela_wire_8048;
    wire new_Jinkela_wire_8864;
    wire new_Jinkela_wire_15979;
    wire new_Jinkela_wire_2307;
    wire new_Jinkela_wire_4819;
    wire _0345_;
    wire new_Jinkela_wire_10197;
    wire new_Jinkela_wire_2620;
    wire new_Jinkela_wire_10332;
    wire new_Jinkela_wire_17809;
    wire new_Jinkela_wire_18727;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_4675;
    wire new_Jinkela_wire_11665;
    wire new_Jinkela_wire_9199;
    wire _0413_;
    wire new_Jinkela_wire_7699;
    wire new_Jinkela_wire_19735;
    wire _0682_;
    wire new_Jinkela_wire_9213;
    wire new_Jinkela_wire_9616;
    wire new_Jinkela_wire_15547;
    wire new_Jinkela_wire_10590;
    wire new_Jinkela_wire_10764;
    wire new_Jinkela_wire_3744;
    wire new_Jinkela_wire_8069;
    wire new_Jinkela_wire_21125;
    wire new_Jinkela_wire_13156;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_1286;
    wire new_Jinkela_wire_12698;
    wire new_Jinkela_wire_6960;
    wire new_Jinkela_wire_15376;
    wire new_Jinkela_wire_3976;
    wire new_Jinkela_wire_7601;
    wire new_Jinkela_wire_10396;
    wire new_Jinkela_wire_10304;
    wire new_Jinkela_wire_15767;
    wire new_Jinkela_wire_7036;
    wire new_Jinkela_wire_13299;
    wire new_Jinkela_wire_15515;
    wire new_Jinkela_wire_16810;
    wire new_Jinkela_wire_8708;
    wire new_Jinkela_wire_8311;
    wire new_Jinkela_wire_6429;
    wire new_Jinkela_wire_12813;
    wire _0266_;
    wire new_Jinkela_wire_11278;
    wire new_Jinkela_wire_7283;
    wire new_Jinkela_wire_15844;
    wire new_Jinkela_wire_4863;
    wire new_Jinkela_wire_17613;
    wire new_Jinkela_wire_4426;
    wire new_Jinkela_wire_7976;
    wire new_Jinkela_wire_14017;
    wire new_Jinkela_wire_11697;
    wire new_Jinkela_wire_9729;
    wire new_Jinkela_wire_16103;
    wire new_Jinkela_wire_18066;
    wire new_Jinkela_wire_13702;
    wire new_Jinkela_wire_13303;
    wire new_Jinkela_wire_3712;
    wire new_Jinkela_wire_18763;
    wire new_Jinkela_wire_3863;
    wire new_Jinkela_wire_12169;
    wire _0897_;
    wire new_Jinkela_wire_13169;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_3321;
    wire new_Jinkela_wire_9674;
    wire new_Jinkela_wire_5861;
    wire new_Jinkela_wire_15904;
    wire new_Jinkela_wire_4995;
    wire new_Jinkela_wire_4927;
    wire new_Jinkela_wire_17926;
    wire new_Jinkela_wire_10264;
    wire new_Jinkela_wire_19908;
    wire new_Jinkela_wire_10656;
    wire new_Jinkela_wire_20160;
    wire new_Jinkela_wire_3044;
    wire new_Jinkela_wire_16245;
    wire new_Jinkela_wire_11161;
    wire new_Jinkela_wire_13738;
    wire new_Jinkela_wire_16845;
    wire new_Jinkela_wire_12254;
    wire new_Jinkela_wire_10666;
    wire new_Jinkela_wire_20146;
    wire new_Jinkela_wire_4065;
    wire new_Jinkela_wire_7034;
    wire new_Jinkela_wire_7399;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_6009;
    wire new_Jinkela_wire_13811;
    wire new_Jinkela_wire_19208;
    wire new_Jinkela_wire_8908;
    wire _1314_;
    wire new_Jinkela_wire_17196;
    wire new_Jinkela_wire_19928;
    wire new_Jinkela_wire_1977;
    wire new_Jinkela_wire_10584;
    wire new_Jinkela_wire_3834;
    wire new_Jinkela_wire_6179;
    wire new_Jinkela_wire_4059;
    wire new_Jinkela_wire_11768;
    wire new_Jinkela_wire_7832;
    wire new_Jinkela_wire_15040;
    wire new_Jinkela_wire_9845;
    wire new_Jinkela_wire_6010;
    wire new_Jinkela_wire_15323;
    wire new_Jinkela_wire_6912;
    wire new_Jinkela_wire_9447;
    wire _1272_;
    wire new_Jinkela_wire_14274;
    wire new_Jinkela_wire_17295;
    wire new_Jinkela_wire_6843;
    wire new_Jinkela_wire_3685;
    wire new_Jinkela_wire_13492;
    wire new_Jinkela_wire_6205;
    wire new_Jinkela_wire_18162;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_5959;
    wire new_Jinkela_wire_18484;
    wire new_Jinkela_wire_9264;
    wire new_Jinkela_wire_18129;
    wire new_Jinkela_wire_6298;
    wire new_Jinkela_wire_14019;
    wire new_Jinkela_wire_12192;
    wire new_Jinkela_wire_3256;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_15521;
    wire new_Jinkela_wire_15469;
    wire new_Jinkela_wire_16258;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_8928;
    wire new_Jinkela_wire_10821;
    wire new_Jinkela_wire_15715;
    wire new_Jinkela_wire_8879;
    wire new_Jinkela_wire_15948;
    wire new_Jinkela_wire_14520;
    wire new_Jinkela_wire_12809;
    wire new_Jinkela_wire_6321;
    wire new_Jinkela_wire_3501;
    wire _1585_;
    wire new_Jinkela_wire_9116;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_5657;
    wire new_Jinkela_wire_15784;
    wire new_Jinkela_wire_3380;
    wire new_Jinkela_wire_17053;
    wire _0015_;
    wire new_Jinkela_wire_18442;
    wire _0842_;
    wire new_Jinkela_wire_5845;
    wire new_Jinkela_wire_4192;
    wire new_Jinkela_wire_3950;
    wire new_Jinkela_wire_3459;
    wire new_Jinkela_wire_5731;
    wire new_Jinkela_wire_17415;
    wire _0591_;
    wire new_Jinkela_wire_9847;
    wire new_Jinkela_wire_8898;
    wire new_Jinkela_wire_9544;
    wire new_Jinkela_wire_14174;
    wire _1118_;
    wire new_Jinkela_wire_3886;
    wire _1628_;
    wire new_Jinkela_wire_8340;
    wire new_Jinkela_wire_21144;
    wire _1589_;
    wire new_Jinkela_wire_9484;
    wire new_Jinkela_wire_10902;
    wire new_Jinkela_wire_12867;
    wire new_Jinkela_wire_15393;
    wire new_Jinkela_wire_18374;
    wire new_Jinkela_wire_15710;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_9740;
    wire new_Jinkela_wire_19940;
    wire new_Jinkela_wire_16393;
    wire new_Jinkela_wire_17595;
    wire new_Jinkela_wire_19111;
    wire new_Jinkela_wire_15519;
    wire new_Jinkela_wire_10779;
    wire new_Jinkela_wire_4633;
    wire new_Jinkela_wire_13258;
    wire new_Jinkela_wire_11478;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_2231;
    wire new_Jinkela_wire_9591;
    wire new_Jinkela_wire_13605;
    wire new_Jinkela_wire_19297;
    wire new_Jinkela_wire_2290;
    wire new_Jinkela_wire_15167;
    wire new_Jinkela_wire_4702;
    wire new_Jinkela_wire_4202;
    wire new_Jinkela_wire_11418;
    wire new_Jinkela_wire_17290;
    wire new_Jinkela_wire_7926;
    wire new_Jinkela_wire_17919;
    wire new_Jinkela_wire_9488;
    wire new_Jinkela_wire_15185;
    wire new_Jinkela_wire_20011;
    wire new_Jinkela_wire_2327;
    wire new_Jinkela_wire_8390;
    wire _1367_;
    wire _0022_;
    wire new_Jinkela_wire_14943;
    wire new_Jinkela_wire_20474;
    wire new_Jinkela_wire_10229;
    wire new_Jinkela_wire_20212;
    wire new_Jinkela_wire_18616;
    wire new_Jinkela_wire_12141;
    wire new_Jinkela_wire_8213;
    wire new_Jinkela_wire_20821;
    wire new_Jinkela_wire_3247;
    wire _0816_;
    wire new_Jinkela_wire_7970;
    wire new_Jinkela_wire_16238;
    wire new_Jinkela_wire_2164;
    wire new_Jinkela_wire_9805;
    wire new_Jinkela_wire_16256;
    wire new_Jinkela_wire_10450;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_8735;
    wire new_Jinkela_wire_19934;
    wire _1735_;
    wire new_Jinkela_wire_13393;
    wire new_Jinkela_wire_13757;
    wire new_Jinkela_wire_19887;
    wire new_Jinkela_wire_16822;
    wire new_Jinkela_wire_1630;
    wire new_Jinkela_wire_20396;
    wire new_Jinkela_wire_3356;
    wire new_Jinkela_wire_20848;
    wire new_Jinkela_wire_13335;
    wire new_Jinkela_wire_3139;
    wire new_Jinkela_wire_4972;
    wire new_Jinkela_wire_10824;
    wire new_Jinkela_wire_20214;
    wire new_Jinkela_wire_7675;
    wire new_Jinkela_wire_14976;
    wire new_Jinkela_wire_2795;
    wire new_Jinkela_wire_16159;
    wire new_Jinkela_wire_11621;
    wire new_Jinkela_wire_4457;
    wire new_Jinkela_wire_10515;
    wire new_Jinkela_wire_4814;
    wire new_Jinkela_wire_8942;
    wire new_Jinkela_wire_12175;
    wire _0330_;
    wire new_Jinkela_wire_2323;
    wire new_Jinkela_wire_17952;
    wire new_Jinkela_wire_8804;
    wire new_Jinkela_wire_6739;
    wire new_Jinkela_wire_16265;
    wire new_Jinkela_wire_15913;
    wire _0188_;
    wire new_Jinkela_wire_9797;
    wire new_Jinkela_wire_20423;
    wire new_Jinkela_wire_2339;
    wire new_Jinkela_wire_13990;
    wire new_Jinkela_wire_12588;
    wire new_Jinkela_wire_18519;
    wire new_Jinkela_wire_12938;
    wire new_Jinkela_wire_20108;
    wire new_Jinkela_wire_538;
    wire _0675_;
    wire new_Jinkela_wire_4538;
    wire new_Jinkela_wire_3101;
    wire new_Jinkela_wire_6356;
    wire _1365_;
    wire new_Jinkela_wire_6086;
    wire new_Jinkela_wire_9940;
    wire new_Jinkela_wire_17514;
    wire _0060_;
    wire new_Jinkela_wire_11951;
    wire new_Jinkela_wire_2068;
    wire new_Jinkela_wire_16782;
    wire new_Jinkela_wire_15227;
    wire new_Jinkela_wire_14621;
    wire new_Jinkela_wire_3809;
    wire new_Jinkela_wire_629;
    wire _1189_;
    wire new_Jinkela_wire_18332;
    wire new_Jinkela_wire_10307;
    wire new_Jinkela_wire_20680;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_20153;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_10684;
    wire _0988_;
    wire new_Jinkela_wire_5156;
    wire new_Jinkela_wire_18439;
    wire new_Jinkela_wire_15683;
    wire new_Jinkela_wire_13457;
    wire new_Jinkela_wire_12357;
    wire new_Jinkela_wire_3308;
    wire new_Jinkela_wire_14523;
    wire _0702_;
    wire new_Jinkela_wire_17104;
    wire new_Jinkela_wire_5543;
    wire new_Jinkela_wire_6757;
    wire new_Jinkela_wire_12289;
    wire new_Jinkela_wire_4174;
    wire new_Jinkela_wire_14711;
    wire new_Jinkela_wire_8170;
    wire new_Jinkela_wire_18700;
    wire new_Jinkela_wire_16733;
    wire new_Jinkela_wire_8081;
    wire new_Jinkela_wire_18578;
    wire new_Jinkela_wire_2124;
    wire _1629_;
    wire new_Jinkela_wire_17525;
    wire new_Jinkela_wire_12305;
    wire new_Jinkela_wire_4581;
    wire new_Jinkela_wire_10982;
    wire new_Jinkela_wire_9478;
    wire _1403_;
    wire new_Jinkela_wire_2664;
    wire new_Jinkela_wire_14057;
    wire new_Jinkela_wire_5121;
    wire new_Jinkela_wire_10471;
    wire new_Jinkela_wire_6141;
    wire new_Jinkela_wire_2709;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_19450;
    wire new_Jinkela_wire_19758;
    wire new_Jinkela_wire_8409;
    wire new_Jinkela_wire_6286;
    wire new_Jinkela_wire_9401;
    wire new_Jinkela_wire_16784;
    wire new_Jinkela_wire_14487;
    wire new_Jinkela_wire_5623;
    wire _0436_;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_3047;
    wire new_Jinkela_wire_3894;
    wire new_Jinkela_wire_14791;
    wire new_Jinkela_wire_15506;
    wire new_Jinkela_wire_8984;
    wire new_Jinkela_wire_2253;
    wire new_Jinkela_wire_7684;
    wire new_Jinkela_wire_9830;
    wire new_Jinkela_wire_7456;
    wire new_Jinkela_wire_19281;
    wire new_Jinkela_wire_13120;
    wire new_Jinkela_wire_13332;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_17893;
    wire new_Jinkela_wire_2218;
    wire new_Jinkela_wire_20055;
    wire new_Jinkela_wire_7418;
    wire new_Jinkela_wire_6171;
    wire new_Jinkela_wire_17748;
    wire new_Jinkela_wire_13294;
    wire new_Jinkela_wire_11829;
    wire new_Jinkela_wire_19119;
    wire new_Jinkela_wire_6418;
    wire new_Jinkela_wire_2739;
    wire _0144_;
    wire new_Jinkela_wire_13805;
    wire new_Jinkela_wire_20681;
    wire new_Jinkela_wire_17783;
    wire new_Jinkela_wire_7378;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_5220;
    wire new_Jinkela_wire_14114;
    wire _0393_;
    wire new_Jinkela_wire_12135;
    wire new_Jinkela_wire_15740;
    wire new_Jinkela_wire_12829;
    wire new_Jinkela_wire_7185;
    wire _1312_;
    wire new_Jinkela_wire_4256;
    wire new_Jinkela_wire_11870;
    wire new_Jinkela_wire_11349;
    wire new_Jinkela_wire_9507;
    wire new_Jinkela_wire_8413;
    wire new_Jinkela_wire_13803;
    wire new_Jinkela_wire_19810;
    wire new_Jinkela_wire_9564;
    wire new_Jinkela_wire_5523;
    wire new_Jinkela_wire_2112;
    wire new_Jinkela_wire_4585;
    wire new_Jinkela_wire_11618;
    wire new_Jinkela_wire_19978;
    wire new_Jinkela_wire_8762;
    wire new_Jinkela_wire_12339;
    wire new_Jinkela_wire_12434;
    wire new_Jinkela_wire_16989;
    wire new_Jinkela_wire_14625;
    wire new_Jinkela_wire_11625;
    wire new_Jinkela_wire_19979;
    wire new_Jinkela_wire_10796;
    wire new_Jinkela_wire_4324;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_9946;
    wire new_Jinkela_wire_19558;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_2566;
    wire new_Jinkela_wire_3930;
    wire new_Jinkela_wire_18011;
    wire new_Jinkela_wire_5599;
    wire new_Jinkela_wire_4182;
    wire new_Jinkela_wire_12545;
    wire new_Jinkela_wire_8580;
    wire new_Jinkela_wire_19860;
    wire new_Jinkela_wire_16523;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_13542;
    wire new_Jinkela_wire_11180;
    wire new_Jinkela_wire_3204;
    wire new_Jinkela_wire_15281;
    wire new_Jinkela_wire_11095;
    wire new_Jinkela_wire_18039;
    wire new_Jinkela_wire_5748;
    wire new_Jinkela_wire_20033;
    wire new_Jinkela_wire_13053;
    wire new_Jinkela_wire_16890;
    wire new_Jinkela_wire_20361;
    wire new_Jinkela_wire_10161;
    wire new_Jinkela_wire_3868;
    wire new_Jinkela_wire_15761;
    wire new_Jinkela_wire_15187;
    wire new_Jinkela_wire_14453;
    wire _1751_;
    wire new_Jinkela_wire_20007;
    wire new_Jinkela_wire_17198;
    wire new_Jinkela_wire_4880;
    wire new_Jinkela_wire_15107;
    wire new_Jinkela_wire_7999;
    wire new_Jinkela_wire_13951;
    wire new_Jinkela_wire_5662;
    wire new_Jinkela_wire_15734;
    wire new_Jinkela_wire_19929;
    wire new_Jinkela_wire_10798;
    wire new_Jinkela_wire_17950;
    wire new_Jinkela_wire_7890;
    wire new_Jinkela_wire_20987;
    wire new_Jinkela_wire_9296;
    wire new_Jinkela_wire_2188;
    wire new_Jinkela_wire_20754;
    wire new_Jinkela_wire_15158;
    wire new_Jinkela_wire_5610;
    wire new_Jinkela_wire_2700;
    wire new_Jinkela_wire_9459;
    wire new_Jinkela_wire_15741;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_15993;
    wire new_Jinkela_wire_18522;
    wire new_Jinkela_wire_1809;
    wire new_Jinkela_wire_7505;
    wire _1216_;
    wire new_Jinkela_wire_11359;
    wire _1789_;
    wire new_Jinkela_wire_15305;
    wire _0509_;
    wire new_Jinkela_wire_12426;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_12910;
    wire new_Jinkela_wire_4669;
    wire new_Jinkela_wire_10449;
    wire new_Jinkela_wire_8665;
    wire _0767_;
    wire new_Jinkela_wire_11873;
    wire new_Jinkela_wire_5045;
    wire new_Jinkela_wire_16625;
    wire new_Jinkela_wire_12529;
    wire new_Jinkela_wire_20303;
    wire _1650_;
    wire new_Jinkela_wire_4767;
    wire new_Jinkela_wire_16040;
    wire new_Jinkela_wire_5272;
    wire new_Jinkela_wire_9326;
    wire new_Jinkela_wire_11361;
    wire _0403_;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_10503;
    wire new_Jinkela_wire_17366;
    wire _1658_;
    wire new_Jinkela_wire_18614;
    wire new_Jinkela_wire_12236;
    wire new_Jinkela_wire_7379;
    wire new_Jinkela_wire_2777;
    wire new_Jinkela_wire_14893;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_17161;
    wire new_Jinkela_wire_7722;
    wire new_Jinkela_wire_8548;
    wire new_Jinkela_wire_6207;
    wire new_Jinkela_wire_18272;
    wire new_Jinkela_wire_7030;
    wire new_Jinkela_wire_13147;
    wire new_Jinkela_wire_14063;
    wire new_Jinkela_wire_20089;
    wire new_Jinkela_wire_10956;
    wire new_Jinkela_wire_8171;
    wire new_Jinkela_wire_10667;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_7253;
    wire new_Jinkela_wire_8538;
    wire new_Jinkela_wire_20538;
    wire new_Jinkela_wire_13390;
    wire new_Jinkela_wire_13551;
    wire new_Jinkela_wire_20535;
    wire new_Jinkela_wire_11581;
    wire _0172_;
    wire new_Jinkela_wire_12712;
    wire new_Jinkela_wire_6765;
    wire new_Jinkela_wire_14015;
    wire new_Jinkela_wire_3547;
    wire new_Jinkela_wire_17017;
    wire new_Jinkela_wire_15611;
    wire new_Jinkela_wire_8881;
    wire new_Jinkela_wire_3768;
    wire new_Jinkela_wire_11533;
    wire _1683_;
    wire new_Jinkela_wire_6446;
    wire new_Jinkela_wire_19032;
    wire new_Jinkela_wire_14645;
    wire new_Jinkela_wire_10898;
    wire new_Jinkela_wire_7515;
    wire new_Jinkela_wire_2461;
    wire new_Jinkela_wire_11541;
    wire new_Jinkela_wire_2884;
    wire new_Jinkela_wire_9127;
    wire new_Jinkela_wire_18638;
    wire new_Jinkela_wire_3143;
    wire new_Jinkela_wire_16706;
    wire new_Jinkela_wire_10042;
    wire new_Jinkela_wire_8913;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_20066;
    wire new_Jinkela_wire_19197;
    wire new_Jinkela_wire_13153;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_6120;
    wire new_Jinkela_wire_3134;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_8809;
    wire new_Jinkela_wire_20051;
    wire new_Jinkela_wire_4014;
    wire new_Jinkela_wire_3552;
    wire _0705_;
    wire new_Jinkela_wire_9719;
    wire new_Jinkela_wire_20620;
    wire _1659_;
    wire new_Jinkela_wire_6375;
    wire new_Jinkela_wire_10554;
    wire new_Jinkela_wire_2252;
    wire new_Jinkela_wire_6039;
    wire new_Jinkela_wire_10231;
    wire new_Jinkela_wire_21277;
    wire new_Jinkela_wire_8958;
    wire new_Jinkela_wire_12643;
    wire new_Jinkela_wire_2654;
    wire new_Jinkela_wire_15988;
    wire new_Jinkela_wire_13535;
    wire new_Jinkela_wire_7500;
    wire new_Jinkela_wire_4276;
    wire new_Jinkela_wire_16031;
    wire _0506_;
    wire new_Jinkela_wire_5641;
    wire new_Jinkela_wire_18934;
    wire new_Jinkela_wire_7188;
    wire new_Jinkela_wire_11390;
    wire new_Jinkela_wire_4273;
    wire new_Jinkela_wire_5775;
    wire new_Jinkela_wire_3986;
    wire _0341_;
    wire new_Jinkela_wire_3381;
    wire new_Jinkela_wire_7840;
    wire _0417_;
    wire new_Jinkela_wire_4619;
    wire new_Jinkela_wire_9483;
    wire new_Jinkela_wire_16577;
    wire new_Jinkela_wire_10501;
    wire new_Jinkela_wire_8329;
    wire new_Jinkela_wire_6370;
    wire new_Jinkela_wire_15034;
    wire new_Jinkela_wire_11925;
    wire new_Jinkela_wire_15336;
    wire new_Jinkela_wire_5998;
    wire new_Jinkela_wire_20135;
    wire new_Jinkela_wire_16421;
    wire _0923_;
    wire new_Jinkela_wire_19852;
    wire new_Jinkela_wire_4677;
    wire new_Jinkela_wire_19171;
    wire new_Jinkela_wire_11647;
    wire new_Jinkela_wire_17798;
    wire new_Jinkela_wire_10735;
    wire new_Jinkela_wire_20356;
    wire new_Jinkela_wire_14884;
    wire new_Jinkela_wire_3288;
    wire _0664_;
    wire new_Jinkela_wire_2121;
    wire new_Jinkela_wire_6111;
    wire new_Jinkela_wire_20669;
    wire _0599_;
    wire new_Jinkela_wire_19309;
    wire new_Jinkela_wire_17339;
    wire _0244_;
    wire new_Jinkela_wire_8978;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_10202;
    wire new_Jinkela_wire_7056;
    wire new_Jinkela_wire_18621;
    wire new_Jinkela_wire_8526;
    wire new_Jinkela_wire_19593;
    wire new_Jinkela_wire_10158;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_11212;
    wire new_Jinkela_wire_7924;
    wire new_Jinkela_wire_1358;
    wire new_Jinkela_wire_9410;
    wire new_Jinkela_wire_6474;
    wire new_Jinkela_wire_1403;
    wire new_Jinkela_wire_2168;
    wire _0677_;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_8155;
    wire new_Jinkela_wire_3805;
    wire new_Jinkela_wire_15958;
    wire new_Jinkela_wire_6324;
    wire new_Jinkela_wire_3613;
    wire new_Jinkela_wire_2893;
    wire new_Jinkela_wire_16033;
    wire new_Jinkela_wire_4683;
    wire new_Jinkela_wire_20092;
    wire new_Jinkela_wire_20687;
    wire new_Jinkela_wire_19601;
    wire new_Jinkela_wire_6630;
    wire new_Jinkela_wire_3860;
    wire new_Jinkela_wire_21238;
    wire new_Jinkela_wire_15265;
    wire new_Jinkela_wire_12300;
    wire new_Jinkela_wire_7408;
    wire _0222_;
    wire _0932_;
    wire new_Jinkela_wire_6319;
    wire new_Jinkela_wire_13199;
    wire new_Jinkela_wire_5333;
    wire new_Jinkela_wire_3949;
    wire _1580_;
    wire new_Jinkela_wire_15698;
    wire new_Jinkela_wire_18145;
    wire _0037_;
    wire new_Jinkela_wire_8423;
    wire new_Jinkela_wire_19062;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_14721;
    wire new_Jinkela_wire_18704;
    wire new_Jinkela_wire_8459;
    wire _1606_;
    wire new_Jinkela_wire_17980;
    wire new_Jinkela_wire_9279;
    wire new_Jinkela_wire_8296;
    wire new_Jinkela_wire_6730;
    wire new_Jinkela_wire_18443;
    wire new_Jinkela_wire_3504;
    wire new_Jinkela_wire_12729;
    wire new_Jinkela_wire_18270;
    wire new_Jinkela_wire_9365;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_1807;
    wire new_Jinkela_wire_11537;
    wire new_Jinkela_wire_4916;
    wire new_Jinkela_wire_1759;
    wire new_Jinkela_wire_3339;
    wire new_Jinkela_wire_6896;
    wire new_Jinkela_wire_19315;
    wire new_Jinkela_wire_9813;
    wire new_Jinkela_wire_15215;
    wire new_Jinkela_wire_3118;
    wire new_Jinkela_wire_11604;
    wire new_Jinkela_wire_5955;
    wire new_Jinkela_wire_11651;
    wire new_Jinkela_wire_17094;
    wire new_Jinkela_wire_7988;
    wire new_Jinkela_wire_10138;
    wire new_Jinkela_wire_5504;
    wire new_Jinkela_wire_4057;
    wire new_Jinkela_wire_2071;
    wire new_Jinkela_wire_8571;
    wire new_Jinkela_wire_10045;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_13608;
    wire new_Jinkela_wire_11219;
    wire new_net_3920;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_4225;
    wire new_Jinkela_wire_4022;
    wire new_Jinkela_wire_5164;
    wire new_Jinkela_wire_12345;
    wire new_Jinkela_wire_2048;
    wire new_Jinkela_wire_20003;
    wire new_Jinkela_wire_6304;
    wire new_Jinkela_wire_3153;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_2589;
    wire new_Jinkela_wire_18105;
    wire new_Jinkela_wire_4757;
    wire new_Jinkela_wire_6260;
    wire new_Jinkela_wire_13526;
    wire new_Jinkela_wire_15589;
    wire new_Jinkela_wire_20046;
    wire new_Jinkela_wire_4414;
    wire new_Jinkela_wire_15944;
    wire new_Jinkela_wire_17768;
    wire new_Jinkela_wire_19168;
    wire new_Jinkela_wire_15867;
    wire _1575_;
    wire new_Jinkela_wire_3226;
    wire new_Jinkela_wire_13001;
    wire new_Jinkela_wire_14985;
    wire _0659_;
    wire new_Jinkela_wire_15601;
    wire new_Jinkela_wire_17097;
    wire new_Jinkela_wire_4712;
    wire new_Jinkela_wire_11848;
    wire new_Jinkela_wire_3964;
    wire _0769_;
    wire new_Jinkela_wire_19376;
    wire new_Jinkela_wire_14255;
    wire new_Jinkela_wire_17078;
    wire _0952_;
    wire new_Jinkela_wire_10478;
    wire _1626_;
    wire new_Jinkela_wire_4857;
    wire new_Jinkela_wire_7850;
    wire new_Jinkela_wire_12044;
    wire new_Jinkela_wire_13859;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_13658;
    wire _1077_;
    wire new_Jinkela_wire_17594;
    wire new_Jinkela_wire_11055;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_20414;
    wire new_Jinkela_wire_3468;
    wire new_Jinkela_wire_17178;
    wire new_Jinkela_wire_18025;
    wire new_Jinkela_wire_12519;
    wire new_Jinkela_wire_11867;
    wire new_Jinkela_wire_16576;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_15608;
    wire new_Jinkela_wire_14980;
    wire new_Jinkela_wire_15916;
    wire new_Jinkela_wire_13769;
    wire new_Jinkela_wire_8414;
    wire new_Jinkela_wire_16067;
    wire new_Jinkela_wire_12971;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_6704;
    wire new_Jinkela_wire_18625;
    wire _1727_;
    wire new_Jinkela_wire_4531;
    wire new_Jinkela_wire_3926;
    wire new_Jinkela_wire_19349;
    wire new_Jinkela_wire_8130;
    wire _1656_;
    wire new_Jinkela_wire_7725;
    wire new_Jinkela_wire_4092;
    wire new_Jinkela_wire_16416;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_15199;
    wire new_Jinkela_wire_5173;
    wire new_Jinkela_wire_1636;
    wire new_net_0;
    wire new_Jinkela_wire_14014;
    wire new_Jinkela_wire_8816;
    wire new_Jinkela_wire_16288;
    wire new_Jinkela_wire_9617;
    wire new_Jinkela_wire_8350;
    wire new_Jinkela_wire_19162;
    wire _1269_;
    wire new_Jinkela_wire_14277;
    wire new_Jinkela_wire_14201;
    wire new_Jinkela_wire_13066;
    wire new_Jinkela_wire_15596;
    wire new_Jinkela_wire_16858;
    wire _0355_;
    wire new_Jinkela_wire_4764;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_17408;
    wire new_Jinkela_wire_13610;
    wire new_Jinkela_wire_18545;
    wire new_Jinkela_wire_5685;
    wire new_Jinkela_wire_18991;
    wire new_Jinkela_wire_10568;
    wire _0546_;
    wire new_Jinkela_wire_18180;
    wire new_Jinkela_wire_17654;
    wire new_Jinkela_wire_13916;
    wire new_Jinkela_wire_7054;
    wire new_Jinkela_wire_1854;
    wire new_Jinkela_wire_6065;
    wire new_Jinkela_wire_3322;
    wire new_Jinkela_wire_6202;
    wire new_Jinkela_wire_3154;
    wire _1454_;
    wire new_Jinkela_wire_19274;
    wire new_Jinkela_wire_6686;
    wire new_Jinkela_wire_9442;
    wire new_Jinkela_wire_13570;
    wire new_Jinkela_wire_17384;
    wire new_Jinkela_wire_3113;
    wire new_Jinkela_wire_7427;
    wire new_Jinkela_wire_5444;
    wire new_Jinkela_wire_4748;
    wire new_Jinkela_wire_6337;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_10542;
    wire _1154_;
    wire new_Jinkela_wire_17048;
    wire new_Jinkela_wire_3008;
    wire new_Jinkela_wire_14247;
    wire new_Jinkela_wire_6890;
    wire new_Jinkela_wire_13756;
    wire new_Jinkela_wire_11385;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_4998;
    wire new_Jinkela_wire_8083;
    wire new_Jinkela_wire_9456;
    wire new_Jinkela_wire_16556;
    wire new_Jinkela_wire_10490;
    wire new_Jinkela_wire_2463;
    wire new_Jinkela_wire_7360;
    wire new_Jinkela_wire_13998;
    wire new_Jinkela_wire_15102;
    wire new_Jinkela_wire_6580;
    wire new_Jinkela_wire_13027;
    wire new_Jinkela_wire_11822;
    wire new_Jinkela_wire_18440;
    wire new_Jinkela_wire_6787;
    wire new_Jinkela_wire_15842;
    wire new_Jinkela_wire_20733;
    wire new_Jinkela_wire_21189;
    wire new_Jinkela_wire_18982;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_9642;
    wire _0356_;
    wire new_Jinkela_wire_9821;
    wire new_Jinkela_wire_3425;
    wire new_Jinkela_wire_13544;
    wire new_Jinkela_wire_8239;
    wire new_Jinkela_wire_6962;
    wire new_Jinkela_wire_21072;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_8607;
    wire new_Jinkela_wire_1702;
    wire new_Jinkela_wire_12954;
    wire new_Jinkela_wire_3175;
    wire new_Jinkela_wire_19350;
    wire new_Jinkela_wire_11810;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_10548;
    wire _0803_;
    wire new_Jinkela_wire_5534;
    wire new_Jinkela_wire_3810;
    wire new_Jinkela_wire_3083;
    wire new_Jinkela_wire_14031;
    wire new_Jinkela_wire_5456;
    wire new_Jinkela_wire_5906;
    wire _0013_;
    wire new_Jinkela_wire_5910;
    wire new_Jinkela_wire_4351;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_19482;
    wire new_Jinkela_wire_17394;
    wire new_Jinkela_wire_16931;
    wire new_Jinkela_wire_5193;
    wire new_Jinkela_wire_3913;
    wire new_Jinkela_wire_16207;
    wire new_Jinkela_wire_15718;
    wire new_Jinkela_wire_10036;
    wire new_Jinkela_wire_17873;
    wire new_Jinkela_wire_11962;
    wire new_Jinkela_wire_3369;
    wire new_Jinkela_wire_17475;
    wire new_Jinkela_wire_15259;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_17236;
    wire new_Jinkela_wire_17772;
    wire new_Jinkela_wire_4121;
    wire new_Jinkela_wire_14522;
    wire new_Jinkela_wire_20954;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_17125;
    wire _0017_;
    wire new_Jinkela_wire_20178;
    wire new_Jinkela_wire_3891;
    wire new_Jinkela_wire_15686;
    wire new_Jinkela_wire_10239;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_9816;
    wire new_Jinkela_wire_4126;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_10968;
    wire new_Jinkela_wire_3817;
    wire new_Jinkela_wire_1063;
    wire _0163_;
    wire new_Jinkela_wire_20124;
    wire new_Jinkela_wire_15687;
    wire new_Jinkela_wire_12703;
    wire new_Jinkela_wire_4384;
    wire new_Jinkela_wire_16252;
    wire new_Jinkela_wire_16247;
    wire new_Jinkela_wire_2831;
    wire new_Jinkela_wire_5371;
    wire new_Jinkela_wire_11874;
    wire new_Jinkela_wire_17231;
    wire new_Jinkela_wire_9953;
    wire new_Jinkela_wire_4903;
    wire new_Jinkela_wire_4491;
    wire new_Jinkela_wire_11208;
    wire new_Jinkela_wire_2838;
    wire new_Jinkela_wire_20320;
    wire new_Jinkela_wire_6528;
    wire new_Jinkela_wire_3295;
    wire new_Jinkela_wire_18899;
    wire new_Jinkela_wire_14744;
    wire new_Jinkela_wire_15294;
    wire _1363_;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_11368;
    wire new_Jinkela_wire_18839;
    wire new_Jinkela_wire_6454;
    wire new_Jinkela_wire_2638;
    wire new_Jinkela_wire_10408;
    wire new_Jinkela_wire_2235;
    wire new_Jinkela_wire_14287;
    wire _1623_;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_5958;
    wire new_Jinkela_wire_5165;
    wire new_Jinkela_wire_10637;
    wire new_Jinkela_wire_6751;
    wire new_Jinkela_wire_12583;
    wire new_Jinkela_wire_3551;
    wire new_Jinkela_wire_5847;
    wire new_Jinkela_wire_17751;
    wire new_Jinkela_wire_6342;
    wire new_Jinkela_wire_5725;
    wire new_Jinkela_wire_1427;
    wire _0199_;
    wire new_Jinkela_wire_15893;
    wire new_Jinkela_wire_20421;
    wire new_Jinkela_wire_8227;
    wire new_Jinkela_wire_17064;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_9048;
    wire new_Jinkela_wire_12495;
    wire new_Jinkela_wire_11952;
    wire new_Jinkela_wire_2462;
    wire new_Jinkela_wire_4965;
    wire new_Jinkela_wire_19544;
    wire new_Jinkela_wire_8276;
    wire _1317_;
    wire new_Jinkela_wire_18343;
    wire new_Jinkela_wire_2428;
    wire new_Jinkela_wire_5989;
    wire new_Jinkela_wire_16816;
    wire new_Jinkela_wire_14322;
    wire new_Jinkela_wire_17796;
    wire new_Jinkela_wire_15493;
    wire new_Jinkela_wire_15175;
    wire new_Jinkela_wire_12817;
    wire new_Jinkela_wire_13096;
    wire new_Jinkela_wire_5667;
    wire new_Jinkela_wire_17646;
    wire new_Jinkela_wire_19772;
    wire new_Jinkela_wire_8682;
    wire new_Jinkela_wire_14757;
    wire new_Jinkela_wire_20191;
    wire new_Jinkela_wire_7322;
    wire new_Jinkela_wire_7717;
    wire new_Jinkela_wire_20121;
    wire new_Jinkela_wire_4762;
    wire new_Jinkela_wire_12790;
    wire new_Jinkela_wire_14965;
    wire new_Jinkela_wire_12567;
    wire new_Jinkela_wire_12771;
    wire new_Jinkela_wire_8467;
    wire new_Jinkela_wire_8163;
    wire new_Jinkela_wire_17728;
    wire new_Jinkela_wire_11605;
    wire new_Jinkela_wire_20429;
    wire new_Jinkela_wire_10168;
    wire new_Jinkela_wire_6709;
    wire new_Jinkela_wire_12099;
    wire new_Jinkela_wire_3421;
    wire new_Jinkela_wire_14190;
    wire new_Jinkela_wire_18589;
    wire _0495_;
    wire new_Jinkela_wire_8067;
    wire new_Jinkela_wire_14682;
    wire new_Jinkela_wire_2224;
    wire new_Jinkela_wire_9379;
    wire new_Jinkela_wire_10300;
    wire new_Jinkela_wire_17354;
    wire new_Jinkela_wire_9083;
    wire new_Jinkela_wire_15827;
    wire new_Jinkela_wire_8658;
    wire new_Jinkela_wire_14392;
    wire _1720_;
    wire new_Jinkela_wire_15541;
    wire new_Jinkela_wire_7549;
    wire new_Jinkela_wire_15149;
    wire new_Jinkela_wire_16628;
    wire new_Jinkela_wire_16604;
    wire new_Jinkela_wire_17040;
    wire new_Jinkela_wire_16349;
    wire new_Jinkela_wire_13119;
    wire new_Jinkela_wire_6835;
    wire new_Jinkela_wire_17116;
    wire new_Jinkela_wire_10732;
    wire new_Jinkela_wire_3235;
    wire new_Jinkela_wire_8108;
    wire new_Jinkela_wire_708;
    wire _0208_;
    wire new_Jinkela_wire_10698;
    wire new_Jinkela_wire_16617;
    wire new_Jinkela_wire_10700;
    wire new_Jinkela_wire_12002;
    wire new_Jinkela_wire_7535;
    wire new_Jinkela_wire_4947;
    wire new_Jinkela_wire_18393;
    wire new_Jinkela_wire_17345;
    wire new_Jinkela_wire_8893;
    wire new_Jinkela_wire_16639;
    wire new_Jinkela_wire_12513;
    wire new_Jinkela_wire_10759;
    wire new_Jinkela_wire_7830;
    wire new_Jinkela_wire_14512;
    wire new_Jinkela_wire_13142;
    wire new_Jinkela_wire_7962;
    wire new_Jinkela_wire_4139;
    wire new_Jinkela_wire_3146;
    wire new_Jinkela_wire_746;
    wire _0467_;
    wire new_Jinkela_wire_10473;
    wire _0549_;
    wire _0588_;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_9817;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_17861;
    wire new_Jinkela_wire_19439;
    wire _0965_;
    wire new_Jinkela_wire_12181;
    wire new_Jinkela_wire_6192;
    wire new_Jinkela_wire_20742;
    wire new_Jinkela_wire_11629;
    wire new_Jinkela_wire_7029;
    wire new_Jinkela_wire_20172;
    wire new_Jinkela_wire_6362;
    wire new_Jinkela_wire_17479;
    wire new_Jinkela_wire_3138;
    wire new_Jinkela_wire_18269;
    wire new_Jinkela_wire_6917;
    wire new_Jinkela_wire_21275;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_10354;
    wire new_Jinkela_wire_5990;
    wire new_Jinkela_wire_10926;
    wire new_Jinkela_wire_20690;
    wire new_Jinkela_wire_9053;
    wire new_Jinkela_wire_19602;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_16028;
    wire new_Jinkela_wire_17889;
    wire new_Jinkela_wire_10599;
    wire new_Jinkela_wire_1655;
    wire new_Jinkela_wire_17706;
    wire new_Jinkela_wire_78;
    wire _1440_;
    wire new_Jinkela_wire_21284;
    wire new_Jinkela_wire_4345;
    wire new_Jinkela_wire_7186;
    wire new_Jinkela_wire_11075;
    wire new_Jinkela_wire_12111;
    wire new_Jinkela_wire_4222;
    wire new_Jinkela_wire_13386;
    wire new_Jinkela_wire_15997;
    wire new_Jinkela_wire_6778;
    wire new_Jinkela_wire_20220;
    wire new_Jinkela_wire_5031;
    wire new_Jinkela_wire_12085;
    wire new_Jinkela_wire_19545;
    wire new_Jinkela_wire_18118;
    wire new_Jinkela_wire_2612;
    wire new_Jinkela_wire_15970;
    wire new_Jinkela_wire_7223;
    wire new_Jinkela_wire_8068;
    wire new_Jinkela_wire_16370;
    wire new_Jinkela_wire_10866;
    wire new_Jinkela_wire_16774;
    wire new_Jinkela_wire_528;
    wire _1161_;
    wire new_Jinkela_wire_12818;
    wire new_Jinkela_wire_20358;
    wire new_Jinkela_wire_20485;
    wire new_Jinkela_wire_19255;
    wire _0683_;
    wire new_Jinkela_wire_6558;
    wire new_Jinkela_wire_13624;
    wire new_Jinkela_wire_10865;
    wire new_Jinkela_wire_12310;
    wire new_Jinkela_wire_7004;
    wire new_Jinkela_wire_9621;
    wire _1755_;
    wire new_Jinkela_wire_15613;
    wire new_Jinkela_wire_6836;
    wire new_Jinkela_wire_20372;
    wire new_Jinkela_wire_4437;
    wire _0703_;
    wire new_Jinkela_wire_6150;
    wire new_Jinkela_wire_17740;
    wire new_Jinkela_wire_3082;
    wire new_Jinkela_wire_18612;
    wire new_Jinkela_wire_14734;
    wire new_Jinkela_wire_11023;
    wire new_Jinkela_wire_7942;
    wire new_Jinkela_wire_20243;
    wire new_Jinkela_wire_12375;
    wire new_Jinkela_wire_9765;
    wire new_Jinkela_wire_7314;
    wire new_Jinkela_wire_5186;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_5763;
    wire new_Jinkela_wire_12352;
    wire new_Jinkela_wire_6147;
    wire _1459_;
    wire new_Jinkela_wire_5724;
    wire new_Jinkela_wire_15552;
    wire new_Jinkela_wire_7106;
    wire new_Jinkela_wire_8699;
    wire new_Jinkela_wire_14307;
    wire new_Jinkela_wire_10650;
    wire new_Jinkela_wire_12876;
    wire new_Jinkela_wire_21188;
    wire new_Jinkela_wire_16955;
    wire new_Jinkela_wire_1086;
    wire new_Jinkela_wire_21059;
    wire new_Jinkela_wire_17827;
    wire new_Jinkela_wire_15665;
    wire new_Jinkela_wire_3388;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_3632;
    wire new_Jinkela_wire_16511;
    wire new_Jinkela_wire_14396;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_18237;
    wire new_Jinkela_wire_18273;
    wire new_Jinkela_wire_3395;
    wire _0166_;
    wire new_Jinkela_wire_577;
    wire _1562_;
    wire new_Jinkela_wire_19204;
    wire new_Jinkela_wire_15932;
    wire new_Jinkela_wire_21133;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_4231;
    wire new_Jinkela_wire_10776;
    wire new_Jinkela_wire_18193;
    wire new_Jinkela_wire_3331;
    wire new_Jinkela_wire_14769;
    wire new_Jinkela_wire_5553;
    wire new_Jinkela_wire_16988;
    wire new_Jinkela_wire_2651;
    wire new_Jinkela_wire_9229;
    wire new_Jinkela_wire_4787;
    wire new_Jinkela_wire_16332;
    wire new_Jinkela_wire_3515;
    wire new_Jinkela_wire_19580;
    wire new_Jinkela_wire_14292;
    wire new_Jinkela_wire_20900;
    wire new_Jinkela_wire_259;
    wire _0071_;
    wire new_Jinkela_wire_3177;
    wire new_Jinkela_wire_3604;
    wire new_Jinkela_wire_11840;
    wire new_Jinkela_wire_8605;
    wire new_Jinkela_wire_19909;
    wire new_Jinkela_wire_20818;
    wire new_Jinkela_wire_13392;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_12677;
    wire new_Jinkela_wire_10661;
    wire new_Jinkela_wire_19683;
    wire new_Jinkela_wire_2388;
    wire new_Jinkela_wire_19433;
    wire new_Jinkela_wire_13905;
    wire new_Jinkela_wire_19995;
    wire new_Jinkela_wire_3566;
    wire new_Jinkela_wire_2913;
    wire new_Jinkela_wire_3184;
    wire new_Jinkela_wire_20359;
    wire _1427_;
    wire new_Jinkela_wire_4805;
    wire new_Jinkela_wire_3084;
    wire new_Jinkela_wire_19537;
    wire new_Jinkela_wire_6383;
    wire new_Jinkela_wire_15144;
    wire _1737_;
    wire new_Jinkela_wire_6297;
    wire new_Jinkela_wire_11136;
    wire new_Jinkela_wire_13354;
    wire new_Jinkela_wire_7871;
    wire new_Jinkela_wire_18990;
    wire new_Jinkela_wire_3793;
    wire new_Jinkela_wire_11784;
    wire new_Jinkela_wire_8553;
    wire new_Jinkela_wire_7928;
    wire new_Jinkela_wire_7983;
    wire new_Jinkela_wire_13879;
    wire new_Jinkela_wire_5309;
    wire new_Jinkela_wire_13135;
    wire new_Jinkela_wire_19725;
    wire new_Jinkela_wire_5242;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_19581;
    wire new_Jinkela_wire_20944;
    wire new_Jinkela_wire_12138;
    wire new_Jinkela_wire_4929;
    wire _1415_;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_10646;
    wire new_Jinkela_wire_9417;
    wire new_Jinkela_wire_5337;
    wire _0234_;
    wire new_Jinkela_wire_21051;
    wire _0867_;
    wire new_Jinkela_wire_20923;
    wire new_Jinkela_wire_17657;
    wire new_Jinkela_wire_19685;
    wire new_Jinkela_wire_11045;
    wire new_Jinkela_wire_20269;
    wire new_Jinkela_wire_3969;
    wire _1069_;
    wire new_Jinkela_wire_2820;
    wire new_Jinkela_wire_18489;
    wire new_Jinkela_wire_5107;
    wire new_Jinkela_wire_7098;
    wire new_Jinkela_wire_16132;
    wire new_Jinkela_wire_11086;
    wire new_Jinkela_wire_21015;
    wire new_Jinkela_wire_2514;
    wire new_Jinkela_wire_12493;
    wire new_Jinkela_wire_5577;
    wire new_Jinkela_wire_17417;
    wire new_Jinkela_wire_8904;
    wire new_Jinkela_wire_15499;
    wire new_Jinkela_wire_14497;
    wire _1462_;
    wire new_Jinkela_wire_14328;
    wire new_Jinkela_wire_2753;
    wire new_Jinkela_wire_17465;
    wire new_Jinkela_wire_10163;
    wire new_Jinkela_wire_4355;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_7080;
    wire new_Jinkela_wire_8715;
    wire new_Jinkela_wire_6540;
    wire new_Jinkela_wire_5009;
    wire new_Jinkela_wire_12144;
    wire _1601_;
    wire new_Jinkela_wire_6582;
    wire _1362_;
    wire _0626_;
    wire new_Jinkela_wire_2660;
    wire new_Jinkela_wire_8996;
    wire new_Jinkela_wire_19999;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_20765;
    wire new_Jinkela_wire_9027;
    wire new_Jinkela_wire_5179;
    wire new_Jinkela_wire_19646;
    wire new_Jinkela_wire_13115;
    wire new_Jinkela_wire_7312;
    wire new_Jinkela_wire_14179;
    wire new_Jinkela_wire_3282;
    wire new_Jinkela_wire_20098;
    wire new_Jinkela_wire_14168;
    wire new_Jinkela_wire_14683;
    wire new_Jinkela_wire_20696;
    wire new_Jinkela_wire_2803;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_10960;
    wire new_Jinkela_wire_14052;
    wire new_Jinkela_wire_20219;
    wire new_Jinkela_wire_2104;
    wire new_Jinkela_wire_21198;
    wire new_Jinkela_wire_3046;
    wire _0958_;
    wire new_Jinkela_wire_8808;
    wire new_Jinkela_wire_20820;
    wire new_Jinkela_wire_6713;
    wire _0727_;
    wire new_Jinkela_wire_15381;
    wire new_Jinkela_wire_2473;
    wire new_Jinkela_wire_2911;
    wire new_Jinkela_wire_2494;
    wire new_Jinkela_wire_13623;
    wire new_Jinkela_wire_16241;
    wire new_Jinkela_wire_10961;
    wire new_Jinkela_wire_16742;
    wire new_Jinkela_wire_16707;
    wire new_Jinkela_wire_10920;
    wire new_Jinkela_wire_17806;
    wire new_Jinkela_wire_2454;
    wire new_Jinkela_wire_8209;
    wire _1335_;
    wire new_Jinkela_wire_10265;
    wire new_Jinkela_wire_11526;
    wire new_Jinkela_wire_14424;
    wire new_Jinkela_wire_4936;
    wire _1813_;
    wire new_Jinkela_wire_8058;
    wire new_Jinkela_wire_11540;
    wire new_Jinkela_wire_10605;
    wire new_Jinkela_wire_11876;
    wire new_Jinkela_wire_6706;
    wire new_Jinkela_wire_9426;
    wire new_Jinkela_wire_7688;
    wire new_Jinkela_wire_11964;
    wire new_Jinkela_wire_9624;
    wire new_Jinkela_wire_1141;
    wire new_Jinkela_wire_7180;
    wire _1302_;
    wire new_Jinkela_wire_15969;
    wire new_Jinkela_wire_14981;
    wire new_Jinkela_wire_11261;
    wire new_Jinkela_wire_6853;
    wire new_Jinkela_wire_3609;
    wire new_Jinkela_wire_4734;
    wire new_Jinkela_wire_6391;
    wire new_Jinkela_wire_12628;
    wire new_Jinkela_wire_3011;
    wire new_Jinkela_wire_20686;
    wire new_Jinkela_wire_9743;
    wire new_Jinkela_wire_10321;
    wire new_Jinkela_wire_21232;
    wire new_Jinkela_wire_4244;
    wire new_Jinkela_wire_7272;
    wire new_Jinkela_wire_4756;
    wire _0182_;
    wire new_Jinkela_wire_3516;
    wire _0282_;
    wire new_Jinkela_wire_5895;
    wire new_Jinkela_wire_3541;
    wire new_Jinkela_wire_2272;
    wire _1773_;
    wire new_Jinkela_wire_3238;
    wire new_Jinkela_wire_13815;
    wire new_Jinkela_wire_16669;
    wire new_Jinkela_wire_2782;
    wire new_Jinkela_wire_20926;
    wire new_Jinkela_wire_5618;
    wire new_Jinkela_wire_15399;
    wire new_Jinkela_wire_13065;
    wire new_Jinkela_wire_10560;
    wire new_Jinkela_wire_5624;
    wire new_Jinkela_wire_2485;
    wire new_Jinkela_wire_10334;
    wire new_Jinkela_wire_14604;
    wire new_Jinkela_wire_580;
    wire _1018_;
    wire new_Jinkela_wire_10988;
    wire new_Jinkela_wire_11811;
    wire new_Jinkela_wire_20207;
    wire new_Jinkela_wire_3777;
    wire new_Jinkela_wire_3967;
    wire new_Jinkela_wire_11971;
    wire new_Jinkela_wire_11025;
    wire new_Jinkela_wire_2898;
    wire new_Jinkela_wire_10148;
    wire new_Jinkela_wire_11007;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_18819;
    wire new_Jinkela_wire_3827;
    wire new_Jinkela_wire_14116;
    wire new_Jinkela_wire_17305;
    wire new_Jinkela_wire_10026;
    wire new_Jinkela_wire_8483;
    wire new_Jinkela_wire_17167;
    wire new_Jinkela_wire_15134;
    wire new_Jinkela_wire_3522;
    wire new_Jinkela_wire_3480;
    wire _1790_;
    wire new_Jinkela_wire_16914;
    wire new_Jinkela_wire_19882;
    wire _0032_;
    wire new_Jinkela_wire_4879;
    wire new_Jinkela_wire_7901;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_13501;
    wire new_Jinkela_wire_17130;
    wire new_Jinkela_wire_9732;
    wire new_Jinkela_wire_7465;
    wire new_Jinkela_wire_3659;
    wire new_Jinkela_wire_11932;
    wire new_Jinkela_wire_4436;
    wire new_Jinkela_wire_18108;
    wire new_Jinkela_wire_19974;
    wire _0920_;
    wire new_Jinkela_wire_4652;
    wire new_Jinkela_wire_5257;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_13825;
    wire new_Jinkela_wire_12884;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_21085;
    wire new_Jinkela_wire_14828;
    wire new_Jinkela_wire_6817;
    wire new_Jinkela_wire_13827;
    wire new_Jinkela_wire_13208;
    wire new_Jinkela_wire_9228;
    wire new_Jinkela_wire_4084;
    wire new_Jinkela_wire_2407;
    wire new_Jinkela_wire_3122;
    wire new_Jinkela_wire_6622;
    wire new_Jinkela_wire_16939;
    wire new_Jinkela_wire_20757;
    wire new_Jinkela_wire_4752;
    wire new_Jinkela_wire_5584;
    wire new_Jinkela_wire_7922;
    wire new_Jinkela_wire_10579;
    wire new_Jinkela_wire_5718;
    wire new_Jinkela_wire_5385;
    wire _1186_;
    wire new_Jinkela_wire_12749;
    wire new_Jinkela_wire_3931;
    wire new_Jinkela_wire_14698;
    wire new_Jinkela_wire_6568;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_10582;
    wire new_Jinkela_wire_8121;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_1755;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_19152;
    wire new_Jinkela_wire_2431;
    wire _0399_;
    wire new_Jinkela_wire_11696;
    wire new_Jinkela_wire_2491;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_18592;
    wire new_Jinkela_wire_7888;
    wire new_Jinkela_wire_8110;
    wire _0379_;
    wire new_Jinkela_wire_9299;
    wire new_Jinkela_wire_18487;
    wire new_Jinkela_wire_18538;
    wire new_Jinkela_wire_13899;
    wire new_Jinkela_wire_20760;
    wire new_Jinkela_wire_20107;
    wire new_Jinkela_wire_7508;
    wire new_Jinkela_wire_18828;
    wire _1538_;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_7883;
    wire new_Jinkela_wire_8300;
    wire new_Jinkela_wire_3533;
    wire new_Jinkela_wire_5228;
    wire new_Jinkela_wire_16787;
    wire new_Jinkela_wire_12882;
    wire new_Jinkela_wire_12726;
    wire new_Jinkela_wire_20682;
    wire new_Jinkela_wire_6781;
    wire new_Jinkela_wire_20989;
    wire new_Jinkela_wire_17367;
    wire new_Jinkela_wire_12608;
    wire new_Jinkela_wire_15882;
    wire new_Jinkela_wire_14426;
    wire new_Jinkela_wire_13316;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_13722;
    wire new_Jinkela_wire_17590;
    wire new_Jinkela_wire_13742;
    wire new_Jinkela_wire_2445;
    wire new_Jinkela_wire_10730;
    wire new_Jinkela_wire_14693;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_4532;
    wire new_Jinkela_wire_18018;
    wire _1395_;
    wire new_Jinkela_wire_3829;
    wire new_Jinkela_wire_10251;
    wire _1492_;
    wire new_Jinkela_wire_9763;
    wire _1453_;
    wire new_Jinkela_wire_11447;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_17443;
    wire new_Jinkela_wire_12256;
    wire new_Jinkela_wire_17878;
    wire new_Jinkela_wire_3005;
    wire new_Jinkela_wire_12145;
    wire new_Jinkela_wire_2953;
    wire new_Jinkela_wire_8627;
    wire new_Jinkela_wire_17381;
    wire new_Jinkela_wire_17106;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_15288;
    wire new_Jinkela_wire_15139;
    wire new_Jinkela_wire_18914;
    wire new_Jinkela_wire_16832;
    wire new_Jinkela_wire_2663;
    wire new_Jinkela_wire_20284;
    wire new_Jinkela_wire_8577;
    wire new_Jinkela_wire_17553;
    wire new_Jinkela_wire_20697;
    wire new_Jinkela_wire_10052;
    wire new_Jinkela_wire_7858;
    wire new_Jinkela_wire_18646;
    wire _1639_;
    wire new_Jinkela_wire_13954;
    wire new_Jinkela_wire_21273;
    wire new_Jinkela_wire_7113;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_2977;
    wire new_Jinkela_wire_5654;
    wire new_Jinkela_wire_9197;
    wire new_Jinkela_wire_10456;
    wire new_Jinkela_wire_5981;
    wire new_Jinkela_wire_17614;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_19826;
    wire new_Jinkela_wire_10;
    wire _0155_;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_8924;
    wire new_Jinkela_wire_13886;
    wire new_Jinkela_wire_21276;
    wire new_Jinkela_wire_14511;
    wire new_Jinkela_wire_20804;
    wire new_Jinkela_wire_19733;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_8964;
    wire new_Jinkela_wire_13282;
    wire new_Jinkela_wire_12118;
    wire new_Jinkela_wire_3574;
    wire new_Jinkela_wire_19160;
    wire new_Jinkela_wire_7579;
    wire new_Jinkela_wire_21157;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_6657;
    wire new_Jinkela_wire_15723;
    wire _1512_;
    wire new_Jinkela_wire_2696;
    wire _0091_;
    wire _1400_;
    wire new_Jinkela_wire_14461;
    wire new_Jinkela_wire_2033;
    wire new_Jinkela_wire_20441;
    wire new_Jinkela_wire_16849;
    wire new_Jinkela_wire_5479;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_3311;
    wire new_Jinkela_wire_10092;
    wire new_Jinkela_wire_5850;
    wire new_Jinkela_wire_17462;
    wire new_Jinkela_wire_18579;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_870;
    wire _0409_;
    wire new_Jinkela_wire_18732;
    wire new_Jinkela_wire_15428;
    wire new_Jinkela_wire_8321;
    wire new_Jinkela_wire_13547;
    wire new_Jinkela_wire_15174;
    wire new_Jinkela_wire_17348;
    wire new_Jinkela_wire_16779;
    wire new_Jinkela_wire_7376;
    wire new_Jinkela_wire_18771;
    wire _0480_;
    wire new_Jinkela_wire_16253;
    wire _0092_;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_9461;
    wire new_Jinkela_wire_15794;
    wire new_Jinkela_wire_20087;
    wire new_Jinkela_wire_17473;
    wire new_Jinkela_wire_15120;
    wire _0869_;
    wire new_Jinkela_wire_2850;
    wire new_Jinkela_wire_12997;
    wire _1212_;
    wire new_Jinkela_wire_9119;
    wire new_Jinkela_wire_17833;
    wire new_Jinkela_wire_13374;
    wire new_Jinkela_wire_2567;
    wire new_Jinkela_wire_19006;
    wire new_Jinkela_wire_20351;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_13245;
    wire new_Jinkela_wire_18230;
    wire new_Jinkela_wire_10044;
    wire new_Jinkela_wire_2239;
    wire new_Jinkela_wire_2556;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_3266;
    wire new_Jinkela_wire_4409;
    wire new_Jinkela_wire_9774;
    wire new_Jinkela_wire_13850;
    wire new_Jinkela_wire_14653;
    wire new_Jinkela_wire_19755;
    wire new_Jinkela_wire_13557;
    wire new_Jinkela_wire_20111;
    wire new_Jinkela_wire_6806;
    wire new_Jinkela_wire_5507;
    wire new_Jinkela_wire_12338;
    wire new_Jinkela_wire_18437;
    wire new_Jinkela_wire_5736;
    wire new_Jinkela_wire_10416;
    wire new_Jinkela_wire_12055;
    wire new_Jinkela_wire_4357;
    wire new_Jinkela_wire_14846;
    wire new_Jinkela_wire_8643;
    wire new_Jinkela_wire_10041;
    wire new_Jinkela_wire_15275;
    wire new_Jinkela_wire_16677;
    wire new_Jinkela_wire_10736;
    wire new_Jinkela_wire_9604;
    wire new_Jinkela_wire_9362;
    wire new_Jinkela_wire_17520;
    wire new_Jinkela_wire_4554;
    wire new_Jinkela_wire_20218;
    wire new_Jinkela_wire_12924;
    wire new_Jinkela_wire_21302;
    wire new_Jinkela_wire_13437;
    wire new_Jinkela_wire_16284;
    wire new_Jinkela_wire_19125;
    wire new_Jinkela_wire_12143;
    wire new_Jinkela_wire_15445;
    wire new_Jinkela_wire_8146;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_16956;
    wire _1124_;
    wire new_Jinkela_wire_17157;
    wire new_Jinkela_wire_2222;
    wire new_Jinkela_wire_9310;
    wire new_Jinkela_wire_3230;
    wire new_Jinkela_wire_8948;
    wire new_Jinkela_wire_2623;
    wire new_Jinkela_wire_18160;
    wire new_Jinkela_wire_1180;
    wire _0171_;
    wire new_Jinkela_wire_19707;
    wire new_Jinkela_wire_9072;
    wire new_Jinkela_wire_3896;
    wire new_Jinkela_wire_8811;
    wire new_Jinkela_wire_19275;
    wire new_Jinkela_wire_4356;
    wire new_Jinkela_wire_7064;
    wire new_Jinkela_wire_4144;
    wire new_Jinkela_wire_6176;
    wire new_Jinkela_wire_1985;
    wire new_Jinkela_wire_7861;
    wire new_Jinkela_wire_5603;
    wire new_Jinkela_wire_14036;
    wire _1264_;
    wire new_Jinkela_wire_15422;
    wire new_Jinkela_wire_17309;
    wire new_Jinkela_wire_15975;
    wire new_Jinkela_wire_9997;
    wire new_Jinkela_wire_13833;
    wire new_Jinkela_wire_6495;
    wire new_Jinkela_wire_16490;
    wire new_Jinkela_wire_9753;
    wire new_Jinkela_wire_6229;
    wire new_Jinkela_wire_19359;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_14743;
    wire new_Jinkela_wire_2580;
    wire new_Jinkela_wire_15881;
    wire new_Jinkela_wire_19991;
    wire new_Jinkela_wire_6903;
    wire new_Jinkela_wire_11590;
    wire new_Jinkela_wire_6390;
    wire _0112_;
    wire _0038_;
    wire new_Jinkela_wire_10971;
    wire new_Jinkela_wire_7353;
    wire new_Jinkela_wire_16915;
    wire _0085_;
    wire new_Jinkela_wire_14483;
    wire new_Jinkela_wire_17540;
    wire new_Jinkela_wire_9099;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_16516;
    wire new_Jinkela_wire_5993;
    wire new_Jinkela_wire_14912;
    wire _0640_;
    wire new_Jinkela_wire_6134;
    wire new_Jinkela_wire_12766;
    wire new_Jinkela_wire_4150;
    wire new_Jinkela_wire_19259;
    wire new_Jinkela_wire_17311;
    wire _1554_;
    wire new_Jinkela_wire_17164;
    wire new_Jinkela_wire_13419;
    wire _1663_;
    wire new_Jinkela_wire_9814;
    wire new_Jinkela_wire_14857;
    wire new_Jinkela_wire_8815;
    wire new_Jinkela_wire_17151;
    wire new_Jinkela_wire_7070;
    wire new_net_3944;
    wire new_Jinkela_wire_9613;
    wire new_Jinkela_wire_10392;
    wire new_Jinkela_wire_2674;
    wire new_Jinkela_wire_18688;
    wire new_Jinkela_wire_14643;
    wire new_Jinkela_wire_21128;
    wire new_Jinkela_wire_11758;
    wire new_Jinkela_wire_12406;
    wire new_Jinkela_wire_8252;
    wire _1646_;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_6933;
    wire new_Jinkela_wire_4207;
    wire new_Jinkela_wire_4495;
    wire _1468_;
    wire new_Jinkela_wire_18929;
    wire new_Jinkela_wire_2232;
    wire new_Jinkela_wire_18176;
    wire new_Jinkela_wire_8297;
    wire new_Jinkela_wire_11284;
    wire new_Jinkela_wire_20450;
    wire new_Jinkela_wire_9269;
    wire new_Jinkela_wire_10833;
    wire new_Jinkela_wire_9327;
    wire new_Jinkela_wire_20633;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_15978;
    wire new_Jinkela_wire_2858;
    wire new_Jinkela_wire_3400;
    wire new_Jinkela_wire_18778;
    wire new_Jinkela_wire_6573;
    wire new_Jinkela_wire_20711;
    wire new_Jinkela_wire_5973;
    wire _1191_;
    wire new_Jinkela_wire_4411;
    wire new_Jinkela_wire_4248;
    wire new_Jinkela_wire_19121;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_12660;
    wire new_Jinkela_wire_17337;
    wire new_Jinkela_wire_9008;
    wire new_Jinkela_wire_10006;
    wire new_Jinkela_wire_6272;
    wire new_Jinkela_wire_9611;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_15569;
    wire _0859_;
    wire new_Jinkela_wire_6514;
    wire new_Jinkela_wire_20126;
    wire new_Jinkela_wire_14629;
    wire _0224_;
    wire new_Jinkela_wire_16651;
    wire new_Jinkela_wire_19090;
    wire _0295_;
    wire new_Jinkela_wire_13965;
    wire new_Jinkela_wire_17357;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_18827;
    wire new_Jinkela_wire_9786;
    wire new_Jinkela_wire_14434;
    wire new_Jinkela_wire_20968;
    wire new_Jinkela_wire_18071;
    wire new_Jinkela_wire_13908;
    wire new_Jinkela_wire_15401;
    wire new_Jinkela_wire_6486;
    wire new_Jinkela_wire_16824;
    wire _1480_;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_9844;
    wire new_Jinkela_wire_16251;
    wire new_Jinkela_wire_11028;
    wire new_Jinkela_wire_7604;
    wire new_Jinkela_wire_5915;
    wire new_Jinkela_wire_13751;
    wire new_Jinkela_wire_2185;
    wire new_Jinkela_wire_9108;
    wire new_Jinkela_wire_7593;
    wire new_Jinkela_wire_20025;
    wire _0836_;
    wire new_Jinkela_wire_4789;
    wire new_Jinkela_wire_18492;
    wire _1434_;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_18020;
    wire new_Jinkela_wire_14858;
    wire new_Jinkela_wire_16720;
    wire new_Jinkela_wire_4155;
    wire _0528_;
    wire new_Jinkela_wire_15110;
    wire new_Jinkela_wire_7525;
    wire new_Jinkela_wire_7131;
    wire new_Jinkela_wire_12742;
    wire new_Jinkela_wire_12682;
    wire new_Jinkela_wire_681;
    wire _0114_;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_9061;
    wire new_Jinkela_wire_16194;
    wire new_Jinkela_wire_2866;
    wire new_Jinkela_wire_5554;
    wire new_Jinkela_wire_9255;
    wire new_Jinkela_wire_10274;
    wire new_Jinkela_wire_4726;
    wire new_Jinkela_wire_21316;
    wire new_Jinkela_wire_14590;
    wire new_Jinkela_wire_17173;
    wire new_Jinkela_wire_4853;
    wire new_Jinkela_wire_13211;
    wire new_Jinkela_wire_9937;
    wire new_Jinkela_wire_10154;
    wire new_Jinkela_wire_15216;
    wire new_Jinkela_wire_8093;
    wire new_Jinkela_wire_20312;
    wire new_Jinkela_wire_20658;
    wire new_Jinkela_wire_4089;
    wire new_Jinkela_wire_7245;
    wire new_Jinkela_wire_6861;
    wire new_Jinkela_wire_15182;
    wire new_Jinkela_wire_3210;
    wire new_Jinkela_wire_21330;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_3813;
    wire new_Jinkela_wire_4026;
    wire new_Jinkela_wire_4694;
    wire new_Jinkela_wire_17328;
    wire new_Jinkela_wire_16397;
    wire new_Jinkela_wire_4004;
    wire new_Jinkela_wire_14160;
    wire new_Jinkela_wire_18050;
    wire new_Jinkela_wire_19822;
    wire new_Jinkela_wire_17447;
    wire new_Jinkela_wire_13429;
    wire new_Jinkela_wire_6714;
    wire _1729_;
    wire new_Jinkela_wire_8036;
    wire new_Jinkela_wire_14971;
    wire new_net_3934;
    wire new_Jinkela_wire_17947;
    wire new_Jinkela_wire_18340;
    wire new_Jinkela_wire_15163;
    wire new_Jinkela_wire_4427;
    wire new_Jinkela_wire_12921;
    wire new_Jinkela_wire_19484;
    wire new_Jinkela_wire_6535;
    wire new_Jinkela_wire_19223;
    wire _0026_;
    wire new_Jinkela_wire_20254;
    wire new_Jinkela_wire_5486;
    wire new_Jinkela_wire_19694;
    wire new_Jinkela_wire_4674;
    wire new_Jinkela_wire_11726;
    wire new_Jinkela_wire_4041;
    wire new_Jinkela_wire_18702;
    wire _0240_;
    wire _0061_;
    wire new_Jinkela_wire_12065;
    wire new_Jinkela_wire_4440;
    wire new_Jinkela_wire_13619;
    wire new_Jinkela_wire_2102;
    wire new_Jinkela_wire_8620;
    wire new_Jinkela_wire_21116;
    wire new_Jinkela_wire_3376;
    wire new_Jinkela_wire_6459;
    wire new_Jinkela_wire_11678;
    wire new_Jinkela_wire_3625;
    wire new_Jinkela_wire_7620;
    wire _0446_;
    wire new_Jinkela_wire_17822;
    wire _0643_;
    wire new_Jinkela_wire_5384;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_8753;
    wire new_Jinkela_wire_18558;
    wire new_Jinkela_wire_14144;
    wire new_Jinkela_wire_6396;
    wire new_Jinkela_wire_15738;
    wire new_Jinkela_wire_11823;
    wire new_Jinkela_wire_11617;
    wire new_Jinkela_wire_17799;
    wire new_Jinkela_wire_4158;
    wire new_Jinkela_wire_2582;
    wire new_Jinkela_wire_6969;
    wire _0394_;
    wire new_Jinkela_wire_4551;
    wire new_Jinkela_wire_11779;
    wire new_Jinkela_wire_13127;
    wire new_Jinkela_wire_11606;
    wire new_Jinkela_wire_2861;
    wire new_Jinkela_wire_13470;
    wire new_Jinkela_wire_16063;
    wire new_Jinkela_wire_15155;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_9090;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_19764;
    wire new_Jinkela_wire_4952;
    wire _0268_;
    wire new_Jinkela_wire_19699;
    wire new_Jinkela_wire_2823;
    wire new_Jinkela_wire_15542;
    wire new_Jinkela_wire_15302;
    wire new_Jinkela_wire_6168;
    wire new_Jinkela_wire_11881;
    wire new_Jinkela_wire_20809;
    wire new_Jinkela_wire_20106;
    wire new_Jinkela_wire_17694;
    wire new_Jinkela_wire_13349;
    wire new_Jinkela_wire_17332;
    wire new_Jinkela_wire_5803;
    wire new_Jinkela_wire_5613;
    wire _0531_;
    wire new_Jinkela_wire_7321;
    wire new_Jinkela_wire_18191;
    wire new_Jinkela_wire_15684;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_7892;
    wire new_Jinkela_wire_9130;
    wire new_Jinkela_wire_8472;
    wire new_Jinkela_wire_12203;
    wire new_Jinkela_wire_15209;
    wire new_Jinkela_wire_18537;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_17263;
    wire new_Jinkela_wire_12451;
    wire new_Jinkela_wire_5751;
    wire new_Jinkela_wire_16853;
    wire new_Jinkela_wire_17547;
    wire new_Jinkela_wire_9077;
    wire new_Jinkela_wire_19347;
    wire new_Jinkela_wire_6060;
    wire new_Jinkela_wire_18065;
    wire new_Jinkela_wire_18952;
    wire new_Jinkela_wire_11032;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_8994;
    wire new_Jinkela_wire_11791;
    wire new_Jinkela_wire_7486;
    wire new_Jinkela_wire_1971;
    wire new_Jinkela_wire_3176;
    wire new_Jinkela_wire_7260;
    wire new_Jinkela_wire_11106;
    wire new_Jinkela_wire_16117;
    wire new_Jinkela_wire_6822;
    wire new_Jinkela_wire_19997;
    wire new_Jinkela_wire_15820;
    wire new_Jinkela_wire_5332;
    wire new_Jinkela_wire_21018;
    wire new_Jinkela_wire_17671;
    wire new_Jinkela_wire_12064;
    wire new_Jinkela_wire_17958;
    wire new_Jinkela_wire_7756;
    wire new_Jinkela_wire_10901;
    wire new_Jinkela_wire_17423;
    wire new_Jinkela_wire_4628;
    wire new_Jinkela_wire_10896;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_13479;
    wire new_Jinkela_wire_19689;
    wire new_Jinkela_wire_9067;
    wire new_Jinkela_wire_17572;
    wire _0343_;
    wire new_Jinkela_wire_2063;
    wire new_Jinkela_wire_18540;
    wire new_Jinkela_wire_18206;
    wire new_Jinkela_wire_10636;
    wire new_Jinkela_wire_6902;
    wire new_Jinkela_wire_13749;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_9960;
    wire new_Jinkela_wire_2584;
    wire new_Jinkela_wire_18317;
    wire new_Jinkela_wire_1425;
    wire _1178_;
    wire new_Jinkela_wire_14316;
    wire _0238_;
    wire new_Jinkela_wire_19233;
    wire _0408_;
    wire new_Jinkela_wire_17585;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_20523;
    wire new_Jinkela_wire_5460;
    wire new_Jinkela_wire_6832;
    wire new_Jinkela_wire_8944;
    wire new_Jinkela_wire_5962;
    wire new_Jinkela_wire_5100;
    wire new_Jinkela_wire_16078;
    wire new_Jinkela_wire_11127;
    wire new_Jinkela_wire_16380;
    wire new_Jinkela_wire_9662;
    wire new_Jinkela_wire_2724;
    wire new_Jinkela_wire_15387;
    wire new_Jinkela_wire_8062;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_18812;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_13573;
    wire _1006_;
    wire new_Jinkela_wire_10871;
    wire new_Jinkela_wire_13821;
    wire new_Jinkela_wire_11279;
    wire new_Jinkela_wire_12789;
    wire new_Jinkela_wire_3560;
    wire new_Jinkela_wire_16691;
    wire new_Jinkela_wire_10317;
    wire new_Jinkela_wire_20773;
    wire new_Jinkela_wire_19300;
    wire new_Jinkela_wire_2240;
    wire new_Jinkela_wire_21252;
    wire new_Jinkela_wire_14122;
    wire new_Jinkela_wire_20008;
    wire new_Jinkela_wire_7425;
    wire new_Jinkela_wire_12725;
    wire _1424_;
    wire new_Jinkela_wire_1722;
    wire new_Jinkela_wire_20415;
    wire new_Jinkela_wire_9195;
    wire new_Jinkela_wire_5342;
    wire new_Jinkela_wire_7474;
    wire new_Jinkela_wire_18163;
    wire new_Jinkela_wire_17668;
    wire new_Jinkela_wire_21044;
    wire _0186_;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_7139;
    wire new_Jinkela_wire_21039;
    wire new_Jinkela_wire_10430;
    wire _0538_;
    wire new_Jinkela_wire_2166;
    wire new_Jinkela_wire_17379;
    wire new_Jinkela_wire_9781;
    wire new_Jinkela_wire_17683;
    wire new_Jinkela_wire_7817;
    wire new_Jinkela_wire_18561;
    wire new_Jinkela_wire_16487;
    wire new_Jinkela_wire_13670;
    wire new_Jinkela_wire_3669;
    wire new_Jinkela_wire_15414;
    wire new_Jinkela_wire_12071;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_11524;
    wire new_Jinkela_wire_19497;
    wire new_Jinkela_wire_7093;
    wire _0048_;
    wire new_Jinkela_wire_11379;
    wire new_Jinkela_wire_15048;
    wire new_Jinkela_wire_9867;
    wire new_Jinkela_wire_11026;
    wire new_Jinkela_wire_11600;
    wire new_Jinkela_wire_20125;
    wire new_Jinkela_wire_17001;
    wire new_Jinkela_wire_3458;
    wire new_Jinkela_wire_9298;
    wire new_Jinkela_wire_17743;
    wire new_Jinkela_wire_18867;
    wire new_Jinkela_wire_8979;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_20080;
    wire new_Jinkela_wire_15003;
    wire _0855_;
    wire new_Jinkela_wire_20783;
    wire new_Jinkela_wire_20737;
    wire new_Jinkela_wire_15571;
    wire new_Jinkela_wire_6125;
    wire _0724_;
    wire new_Jinkela_wire_4251;
    wire new_Jinkela_wire_12642;
    wire new_Jinkela_wire_5210;
    wire new_Jinkela_wire_7102;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_13655;
    wire new_Jinkela_wire_20548;
    wire new_Jinkela_wire_16979;
    wire new_Jinkela_wire_15063;
    wire new_Jinkela_wire_21146;
    wire new_Jinkela_wire_5655;
    wire new_Jinkela_wire_12423;
    wire new_Jinkela_wire_19864;
    wire new_Jinkela_wire_5074;
    wire new_Jinkela_wire_4637;
    wire new_Jinkela_wire_11184;
    wire new_Jinkela_wire_5627;
    wire new_Jinkela_wire_7203;
    wire new_Jinkela_wire_19488;
    wire new_Jinkela_wire_18495;
    wire new_Jinkela_wire_4954;
    wire new_Jinkela_wire_16297;
    wire new_Jinkela_wire_15116;
    wire new_Jinkela_wire_12438;
    wire new_Jinkela_wire_15295;
    wire new_Jinkela_wire_12252;
    wire new_Jinkela_wire_10051;
    wire new_Jinkela_wire_16077;
    wire new_Jinkela_wire_6956;
    wire new_Jinkela_wire_19742;
    wire new_Jinkela_wire_5487;
    wire new_Jinkela_wire_10603;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_8967;
    wire new_Jinkela_wire_10096;
    wire new_Jinkela_wire_14473;
    wire new_Jinkela_wire_15310;
    wire new_Jinkela_wire_9118;
    wire new_Jinkela_wire_1987;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_20018;
    wire new_Jinkela_wire_9521;
    wire new_Jinkela_wire_14878;
    wire new_Jinkela_wire_5318;
    wire new_Jinkela_wire_21195;
    wire new_Jinkela_wire_16130;
    wire new_Jinkela_wire_7332;
    wire new_Jinkela_wire_12200;
    wire new_Jinkela_wire_2470;
    wire new_Jinkela_wire_5514;
    wire new_Jinkela_wire_10531;
    wire new_Jinkela_wire_6711;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_19008;
    wire new_Jinkela_wire_18085;
    wire new_Jinkela_wire_12868;
    wire new_Jinkela_wire_11983;
    wire new_Jinkela_wire_8258;
    wire _0755_;
    wire new_Jinkela_wire_15636;
    wire new_Jinkela_wire_12130;
    wire new_Jinkela_wire_3840;
    wire new_Jinkela_wire_11909;
    wire new_Jinkela_wire_13691;
    wire new_Jinkela_wire_8156;
    wire new_Jinkela_wire_17162;
    wire new_Jinkela_wire_14039;
    wire new_Jinkela_wire_6690;
    wire new_Jinkela_wire_13755;
    wire new_Jinkela_wire_12224;
    wire new_Jinkela_wire_16944;
    wire new_Jinkela_wire_5244;
    wire _0695_;
    wire new_Jinkela_wire_21313;
    wire new_Jinkela_wire_17689;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_9576;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_2127;
    wire new_Jinkela_wire_7697;
    wire new_Jinkela_wire_20513;
    wire new_Jinkela_wire_13663;
    wire new_Jinkela_wire_20575;
    wire new_Jinkela_wire_6680;
    wire new_Jinkela_wire_7770;
    wire new_Jinkela_wire_4895;
    wire new_Jinkela_wire_17675;
    wire _0593_;
    wire new_Jinkela_wire_10957;
    wire new_Jinkela_wire_10521;
    wire new_Jinkela_wire_13716;
    wire new_Jinkela_wire_18527;
    wire new_Jinkela_wire_1485;
    wire new_Jinkela_wire_18112;
    wire new_Jinkela_wire_15805;
    wire new_Jinkela_wire_21036;
    wire _1536_;
    wire new_Jinkela_wire_13563;
    wire new_Jinkela_wire_11641;
    wire _0766_;
    wire new_Jinkela_wire_21199;
    wire new_Jinkela_wire_9912;
    wire _1377_;
    wire new_Jinkela_wire_17297;
    wire new_Jinkela_wire_436;
    wire _1126_;
    wire new_Jinkela_wire_17899;
    wire new_Jinkela_wire_1895;
    wire new_Jinkela_wire_7925;
    wire new_Jinkela_wire_5004;
    wire new_Jinkela_wire_6242;
    wire new_Jinkela_wire_17561;
    wire new_Jinkela_wire_10939;
    wire _0308_;
    wire new_Jinkela_wire_4103;
    wire new_Jinkela_wire_6166;
    wire new_Jinkela_wire_2974;
    wire _0420_;
    wire new_Jinkela_wire_8835;
    wire new_Jinkela_wire_5266;
    wire new_Jinkela_wire_13201;
    wire new_Jinkela_wire_19883;
    wire new_Jinkela_wire_14407;
    wire new_Jinkela_wire_18035;
    wire new_Jinkela_wire_18992;
    wire new_Jinkela_wire_15826;
    wire new_Jinkela_wire_15221;
    wire new_Jinkela_wire_14814;
    wire new_Jinkela_wire_20464;
    wire new_Jinkela_wire_17043;
    wire new_Jinkela_wire_10286;
    wire new_Jinkela_wire_19775;
    wire new_Jinkela_wire_4031;
    wire new_Jinkela_wire_13883;
    wire new_Jinkela_wire_13765;
    wire new_Jinkela_wire_6905;
    wire _0292_;
    wire new_Jinkela_wire_13025;
    wire new_Jinkela_wire_3319;
    wire new_Jinkela_wire_1786;
    wire new_Jinkela_wire_11530;
    wire new_Jinkela_wire_4955;
    wire new_Jinkela_wire_9378;
    wire new_Jinkela_wire_6414;
    wire new_Jinkela_wire_19460;
    wire new_Jinkela_wire_18238;
    wire new_Jinkela_wire_18964;
    wire new_Jinkela_wire_10062;
    wire new_Jinkela_wire_10019;
    wire new_Jinkela_wire_17089;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_6784;
    wire new_Jinkela_wire_11326;
    wire new_Jinkela_wire_17817;
    wire new_Jinkela_wire_16197;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_7343;
    wire new_Jinkela_wire_19635;
    wire new_Jinkela_wire_20747;
    wire new_Jinkela_wire_2486;
    wire new_Jinkela_wire_20168;
    wire _1426_;
    wire new_Jinkela_wire_12552;
    wire new_Jinkela_wire_6970;
    wire new_Jinkela_wire_10838;
    wire new_Jinkela_wire_6913;
    wire new_Jinkela_wire_4422;
    wire new_Jinkela_wire_6772;
    wire new_Jinkela_wire_18111;
    wire new_Jinkela_wire_20865;
    wire new_Jinkela_wire_14986;
    wire _0079_;
    wire new_Jinkela_wire_3704;
    wire new_Jinkela_wire_13974;
    wire new_Jinkela_wire_19590;
    wire new_Jinkela_wire_8730;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_9120;
    wire new_Jinkela_wire_13837;
    wire _1770_;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_21104;
    wire new_Jinkela_wire_2870;
    wire new_Jinkela_wire_11497;
    wire new_Jinkela_wire_11054;
    wire new_Jinkela_wire_9784;
    wire new_Jinkela_wire_14995;
    wire new_Jinkela_wire_4724;
    wire new_Jinkela_wire_17776;
    wire new_Jinkela_wire_8481;
    wire new_Jinkela_wire_19577;
    wire new_Jinkela_wire_9921;
    wire new_Jinkela_wire_7513;
    wire new_Jinkela_wire_12826;
    wire new_Jinkela_wire_6409;
    wire new_Jinkela_wire_4045;
    wire new_Jinkela_wire_3766;
    wire new_Jinkela_wire_5170;
    wire new_Jinkela_wire_16365;
    wire new_Jinkela_wire_19523;
    wire new_Jinkela_wire_4403;
    wire new_Jinkela_wire_14881;
    wire new_Jinkela_wire_8535;
    wire new_Jinkela_wire_2829;
    wire new_Jinkela_wire_2476;
    wire new_Jinkela_wire_13035;
    wire new_Jinkela_wire_15298;
    wire new_Jinkela_wire_18830;
    wire new_Jinkela_wire_17086;
    wire new_Jinkela_wire_20282;
    wire new_Jinkela_wire_6621;
    wire new_Jinkela_wire_4573;
    wire new_Jinkela_wire_7990;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_11583;
    wire new_Jinkela_wire_7174;
    wire new_Jinkela_wire_2613;
    wire new_Jinkela_wire_16120;
    wire new_Jinkela_wire_19454;
    wire new_Jinkela_wire_16670;
    wire new_Jinkela_wire_19276;
    wire new_Jinkela_wire_16044;
    wire new_Jinkela_wire_11927;
    wire new_Jinkela_wire_14000;
    wire new_Jinkela_wire_15462;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_15280;
    wire new_Jinkela_wire_11008;
    wire new_Jinkela_wire_5392;
    wire _0699_;
    wire new_Jinkela_wire_4870;
    wire new_Jinkela_wire_2478;
    wire new_Jinkela_wire_12397;
    wire new_Jinkela_wire_14530;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_3936;
    wire new_Jinkela_wire_21145;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_9359;
    wire _0819_;
    wire new_Jinkela_wire_10437;
    wire new_Jinkela_wire_21058;
    wire new_Jinkela_wire_7528;
    wire new_Jinkela_wire_9812;
    wire new_Jinkela_wire_6488;
    wire new_Jinkela_wire_6153;
    wire new_Jinkela_wire_13649;
    wire new_Jinkela_wire_5021;
    wire new_Jinkela_wire_8376;
    wire new_Jinkela_wire_11142;
    wire new_Jinkela_wire_4539;
    wire _1128_;
    wire new_Jinkela_wire_16041;
    wire new_Jinkela_wire_11957;
    wire new_Jinkela_wire_3299;
    wire new_Jinkela_wire_6428;
    wire _0558_;
    wire _0285_;
    wire new_Jinkela_wire_12205;
    wire new_Jinkela_wire_20725;
    wire new_Jinkela_wire_14596;
    wire new_Jinkela_wire_10174;
    wire new_Jinkela_wire_14182;
    wire new_Jinkela_wire_8253;
    wire new_Jinkela_wire_20660;
    wire _0127_;
    wire new_Jinkela_wire_17283;
    wire new_Jinkela_wire_16339;
    wire new_Jinkela_wire_15709;
    wire new_Jinkela_wire_13927;
    wire new_Jinkela_wire_4293;
    wire new_Jinkela_wire_4812;
    wire new_Jinkela_wire_8154;
    wire new_Jinkela_wire_16837;
    wire new_Jinkela_wire_17148;
    wire new_Jinkela_wire_7886;
    wire _0049_;
    wire new_Jinkela_wire_12639;
    wire new_Jinkela_wire_6867;
    wire new_Jinkela_wire_3856;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_10539;
    wire new_Jinkela_wire_6559;
    wire new_Jinkela_wire_17662;
    wire new_Jinkela_wire_5754;
    wire new_Jinkela_wire_17063;
    wire new_Jinkela_wire_13302;
    wire new_Jinkela_wire_11167;
    wire _1642_;
    wire new_Jinkela_wire_2922;
    wire new_Jinkela_wire_2484;
    wire _0003_;
    wire _1550_;
    wire new_Jinkela_wire_18355;
    wire new_Jinkela_wire_20386;
    wire new_Jinkela_wire_19239;
    wire new_Jinkela_wire_3928;
    wire new_Jinkela_wire_11797;
    wire new_Jinkela_wire_9239;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_16558;
    wire new_Jinkela_wire_19905;
    wire new_Jinkela_wire_10372;
    wire new_Jinkela_wire_11561;
    wire new_Jinkela_wire_12165;
    wire new_Jinkela_wire_13520;
    wire new_Jinkela_wire_5896;
    wire new_Jinkela_wire_18404;
    wire new_Jinkela_wire_11682;
    wire new_Jinkela_wire_4940;
    wire new_Jinkela_wire_17749;
    wire new_Jinkela_wire_13373;
    wire new_Jinkela_wire_14040;
    wire new_Jinkela_wire_16215;
    wire new_Jinkela_wire_18432;
    wire new_Jinkela_wire_10494;
    wire new_Jinkela_wire_4598;
    wire new_Jinkela_wire_12208;
    wire new_Jinkela_wire_15951;
    wire new_Jinkela_wire_16804;
    wire new_Jinkela_wire_5747;
    wire new_Jinkela_wire_12405;
    wire new_Jinkela_wire_19522;
    wire new_Jinkela_wire_12034;
    wire new_Jinkela_wire_2502;
    wire new_Jinkela_wire_10395;
    wire new_Jinkela_wire_5535;
    wire new_Jinkela_wire_11042;
    wire new_Jinkela_wire_14960;
    wire new_Jinkela_wire_10711;
    wire _1243_;
    wire _1802_;
    wire new_Jinkela_wire_12754;
    wire new_Jinkela_wire_18976;
    wire new_Jinkela_wire_16076;
    wire new_Jinkela_wire_20132;
    wire new_Jinkela_wire_13644;
    wire new_Jinkela_wire_4391;
    wire new_Jinkela_wire_17647;
    wire new_Jinkela_wire_9748;
    wire new_Jinkela_wire_18893;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_16038;
    wire new_Jinkela_wire_7424;
    wire new_Jinkela_wire_13588;
    wire new_Jinkela_wire_16006;
    wire new_Jinkela_wire_10945;
    wire new_Jinkela_wire_14457;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_4540;
    wire new_Jinkela_wire_12351;
    wire new_Jinkela_wire_6503;
    wire new_Jinkela_wire_15612;
    wire new_Jinkela_wire_12452;
    wire new_Jinkela_wire_6014;
    wire new_Jinkela_wire_3411;
    wire new_Jinkela_wire_13878;
    wire new_Jinkela_wire_3953;
    wire _1040_;
    wire new_Jinkela_wire_13898;
    wire new_Jinkela_wire_310;
    wire new_Jinkela_wire_9140;
    wire new_Jinkela_wire_14098;
    wire _0508_;
    wire _0648_;
    wire new_Jinkela_wire_10465;
    wire new_Jinkela_wire_19106;
    wire new_Jinkela_wire_9543;
    wire new_Jinkela_wire_10543;
    wire new_Jinkela_wire_20434;
    wire new_Jinkela_wire_14458;
    wire new_Jinkela_wire_12955;
    wire new_Jinkela_wire_19573;
    wire new_Jinkela_wire_13401;
    wire new_Jinkela_wire_2291;
    wire new_Jinkela_wire_19402;
    wire new_Jinkela_wire_6274;
    wire new_Jinkela_wire_17880;
    wire new_Jinkela_wire_2095;
    wire new_Jinkela_wire_5085;
    wire new_Jinkela_wire_9759;
    wire new_Jinkela_wire_5027;
    wire new_Jinkela_wire_16052;
    wire new_Jinkela_wire_18451;
    wire new_Jinkela_wire_1880;
    wire new_Jinkela_wire_13058;
    wire _1503_;
    wire new_Jinkela_wire_14198;
    wire new_Jinkela_wire_4183;
    wire new_Jinkela_wire_6725;
    wire _0690_;
    wire new_Jinkela_wire_6301;
    wire new_Jinkela_wire_15142;
    wire new_Jinkela_wire_4330;
    wire new_Jinkela_wire_8677;
    wire new_Jinkela_wire_7068;
    wire new_Jinkela_wire_5855;
    wire new_Jinkela_wire_3182;
    wire new_Jinkela_wire_11630;
    wire new_Jinkela_wire_19486;
    wire new_Jinkela_wire_5511;
    wire new_Jinkela_wire_13450;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_16638;
    wire new_Jinkela_wire_18970;
    wire _1004_;
    wire new_Jinkela_wire_19519;
    wire new_Jinkela_wire_14541;
    wire new_Jinkela_wire_13842;
    wire new_Jinkela_wire_16151;
    wire new_Jinkela_wire_14910;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_7216;
    wire _1611_;
    wire new_Jinkela_wire_8850;
    wire new_Jinkela_wire_18058;
    wire new_Jinkela_wire_3341;
    wire new_Jinkela_wire_11560;
    wire new_Jinkela_wire_19834;
    wire _0996_;
    wire new_Jinkela_wire_8560;
    wire new_Jinkela_wire_3653;
    wire new_Jinkela_wire_2201;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_21266;
    wire new_Jinkela_wire_8829;
    wire _0676_;
    wire new_Jinkela_wire_3772;
    wire _0628_;
    wire new_Jinkela_wire_4220;
    wire new_Jinkela_wire_13747;
    wire new_Jinkela_wire_10432;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_12982;
    wire new_Jinkela_wire_9605;
    wire new_Jinkela_wire_3536;
    wire new_Jinkela_wire_12073;
    wire new_Jinkela_wire_6738;
    wire new_Jinkela_wire_4671;
    wire new_Jinkela_wire_12618;
    wire new_Jinkela_wire_2497;
    wire new_Jinkela_wire_14627;
    wire new_Jinkela_wire_19049;
    wire new_Jinkela_wire_11458;
    wire new_Jinkela_wire_17012;
    wire new_Jinkela_wire_9677;
    wire new_Jinkela_wire_19179;
    wire new_Jinkela_wire_13177;
    wire new_Jinkela_wire_3442;
    wire new_Jinkela_wire_11863;
    wire new_Jinkela_wire_9446;
    wire new_Jinkela_wire_17095;
    wire new_Jinkela_wire_7667;
    wire new_Jinkela_wire_11226;
    wire new_Jinkela_wire_11666;
    wire new_Jinkela_wire_14275;
    wire new_Jinkela_wire_5619;
    wire new_Jinkela_wire_15153;
    wire new_Jinkela_wire_11237;
    wire new_Jinkela_wire_7063;
    wire new_Jinkela_wire_17696;
    wire new_Jinkela_wire_19741;
    wire new_Jinkela_wire_21253;
    wire new_Jinkela_wire_10738;
    wire new_Jinkela_wire_7060;
    wire new_Jinkela_wire_16536;
    wire new_Jinkela_wire_18086;
    wire new_Jinkela_wire_4613;
    wire new_Jinkela_wire_5947;
    wire new_Jinkela_wire_12360;
    wire new_Jinkela_wire_12335;
    wire new_Jinkela_wire_2469;
    wire new_Jinkela_wire_19387;
    wire new_Jinkela_wire_9062;
    wire new_Jinkela_wire_10614;
    wire new_Jinkela_wire_16619;
    wire new_Jinkela_wire_9339;
    wire new_Jinkela_wire_2792;
    wire new_Jinkela_wire_9707;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_18640;
    wire new_Jinkela_wire_6873;
    wire new_Jinkela_wire_8934;
    wire new_Jinkela_wire_18023;
    wire new_Jinkela_wire_10719;
    wire _0632_;
    wire _1180_;
    wire new_Jinkela_wire_5184;
    wire new_Jinkela_wire_12870;
    wire new_Jinkela_wire_13013;
    wire new_Jinkela_wire_3216;
    wire new_Jinkela_wire_10511;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_9300;
    wire new_Jinkela_wire_7516;
    wire _0309_;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_11652;
    wire new_Jinkela_wire_12560;
    wire new_Jinkela_wire_13325;
    wire new_Jinkela_wire_14334;
    wire new_Jinkela_wire_15148;
    wire _0568_;
    wire new_Jinkela_wire_12692;
    wire new_Jinkela_wire_18268;
    wire new_Jinkela_wire_14113;
    wire new_Jinkela_wire_2571;
    wire new_Jinkela_wire_18648;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_12830;
    wire new_Jinkela_wire_4387;
    wire new_Jinkela_wire_10038;
    wire new_Jinkela_wire_7148;
    wire new_Jinkela_wire_8453;
    wire new_Jinkela_wire_13744;
    wire new_Jinkela_wire_18935;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_13291;
    wire new_Jinkela_wire_17812;
    wire new_Jinkela_wire_5322;
    wire new_Jinkela_wire_13028;
    wire new_Jinkela_wire_8690;
    wire new_Jinkela_wire_16738;
    wire new_Jinkela_wire_18179;
    wire new_Jinkela_wire_17286;
    wire new_Jinkela_wire_5832;
    wire new_Jinkela_wire_10439;
    wire new_Jinkela_wire_11352;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_20506;
    wire new_Jinkela_wire_15872;
    wire new_Jinkela_wire_18871;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_6726;
    wire new_Jinkela_wire_1671;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_1507;
    wire _1490_;
    wire new_Jinkela_wire_6007;
    wire new_Jinkela_wire_17875;
    wire new_Jinkela_wire_18415;
    wire new_Jinkela_wire_20579;
    wire new_Jinkela_wire_6538;
    wire new_Jinkela_wire_12581;
    wire new_Jinkela_wire_2001;
    wire new_Jinkela_wire_11714;
    wire new_Jinkela_wire_12702;
    wire new_Jinkela_wire_18263;
    wire new_Jinkela_wire_4137;
    wire new_Jinkela_wire_8652;
    wire new_Jinkela_wire_18285;
    wire new_Jinkela_wire_8765;
    wire new_Jinkela_wire_10996;
    wire new_Jinkela_wire_12825;
    wire new_Jinkela_wire_16307;
    wire new_Jinkela_wire_2601;
    wire new_Jinkela_wire_3088;
    wire new_Jinkela_wire_8011;
    wire _1539_;
    wire new_Jinkela_wire_11800;
    wire new_Jinkela_wire_5749;
    wire new_Jinkela_wire_14917;
    wire new_Jinkela_wire_14508;
    wire new_Jinkela_wire_18096;
    wire new_Jinkela_wire_3320;
    wire new_Jinkela_wire_19108;
    wire _1596_;
    wire new_Jinkela_wire_18787;
    wire _0181_;
    wire new_Jinkela_wire_16560;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_18740;
    wire new_Jinkela_wire_5794;
    wire new_Jinkela_wire_14016;
    wire new_Jinkela_wire_12488;
    wire new_Jinkela_wire_6634;
    wire new_Jinkela_wire_6729;
    wire new_Jinkela_wire_17808;
    wire new_Jinkela_wire_12366;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_17554;
    wire new_Jinkela_wire_2632;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_3709;
    wire new_Jinkela_wire_6450;
    wire new_Jinkela_wire_6033;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_3289;
    wire new_Jinkela_wire_2915;
    wire new_Jinkela_wire_9347;
    wire new_Jinkela_wire_19083;
    wire new_Jinkela_wire_4562;
    wire new_Jinkela_wire_2078;
    wire new_Jinkela_wire_16335;
    wire new_Jinkela_wire_14563;
    wire new_Jinkela_wire_12549;
    wire new_Jinkela_wire_12054;
    wire new_Jinkela_wire_16807;
    wire new_Jinkela_wire_16157;
    wire new_Jinkela_wire_12240;
    wire new_Jinkela_wire_20382;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_7165;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_11135;
    wire new_Jinkela_wire_15344;
    wire new_Jinkela_wire_6248;
    wire new_Jinkela_wire_2786;
    wire new_Jinkela_wire_13693;
    wire new_Jinkela_wire_4299;
    wire new_Jinkela_wire_6604;
    wire new_Jinkela_wire_12880;
    wire new_Jinkela_wire_14146;
    wire new_Jinkela_wire_10763;
    wire new_Jinkela_wire_20671;
    wire new_Jinkela_wire_4000;
    wire _0307_;
    wire new_Jinkela_wire_15510;
    wire new_Jinkela_wire_19428;
    wire new_Jinkela_wire_9890;
    wire new_Jinkela_wire_10658;
    wire new_Jinkela_wire_15533;
    wire new_Jinkela_wire_17591;
    wire _1376_;
    wire new_Jinkela_wire_4966;
    wire new_Jinkela_wire_6239;
    wire new_Jinkela_wire_9385;
    wire new_Jinkela_wire_4304;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_16271;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_21219;
    wire new_Jinkela_wire_14765;
    wire new_Jinkela_wire_20291;
    wire new_Jinkela_wire_20457;
    wire new_Jinkela_wire_11252;
    wire new_Jinkela_wire_6161;
    wire new_Jinkela_wire_4312;
    wire new_Jinkela_wire_9636;
    wire new_Jinkela_wire_9054;
    wire _1444_;
    wire new_Jinkela_wire_3672;
    wire new_Jinkela_wire_3433;
    wire new_Jinkela_wire_13760;
    wire new_Jinkela_wire_16846;
    wire new_Jinkela_wire_17529;
    wire new_Jinkela_wire_9491;
    wire new_Jinkela_wire_7426;
    wire new_Jinkela_wire_19217;
    wire _0490_;
    wire new_Jinkela_wire_8794;
    wire new_Jinkela_wire_14803;
    wire new_Jinkela_wire_9911;
    wire new_Jinkela_wire_17466;
    wire new_Jinkela_wire_9525;
    wire new_Jinkela_wire_8455;
    wire new_Jinkela_wire_8849;
    wire new_Jinkela_wire_2989;
    wire new_Jinkela_wire_14189;
    wire new_Jinkela_wire_11039;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_3762;
    wire new_Jinkela_wire_5250;
    wire new_Jinkela_wire_19054;
    wire new_Jinkela_wire_13963;
    wire new_Jinkela_wire_8277;
    wire new_Jinkela_wire_7406;
    wire new_Jinkela_wire_3151;
    wire new_Jinkela_wire_2373;
    wire new_Jinkela_wire_19937;
    wire new_Jinkela_wire_13007;
    wire _0915_;
    wire _0949_;
    wire new_Jinkela_wire_13816;
    wire new_Jinkela_wire_12302;
    wire new_Jinkela_wire_3767;
    wire new_Jinkela_wire_13002;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_8544;
    wire new_Jinkela_wire_4201;
    wire new_Jinkela_wire_19918;
    wire new_Jinkela_wire_6417;
    wire new_Jinkela_wire_11448;
    wire _0332_;
    wire new_Jinkela_wire_20552;
    wire new_Jinkela_wire_16699;
    wire new_Jinkela_wire_16449;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_16129;
    wire _1293_;
    wire new_Jinkela_wire_3111;
    wire new_Jinkela_wire_13969;
    wire new_Jinkela_wire_13370;
    wire new_Jinkela_wire_14264;
    wire new_Jinkela_wire_4707;
    wire new_Jinkela_wire_16689;
    wire new_Jinkela_wire_15823;
    wire new_Jinkela_wire_16538;
    wire new_Jinkela_wire_20582;
    wire new_Jinkela_wire_13707;
    wire new_Jinkela_wire_6760;
    wire new_Jinkela_wire_2361;
    wire new_Jinkela_wire_17665;
    wire new_Jinkela_wire_15093;
    wire new_Jinkela_wire_12100;
    wire new_Jinkela_wire_17403;
    wire new_Jinkela_wire_17867;
    wire new_Jinkela_wire_3035;
    wire new_Jinkela_wire_14949;
    wire new_Jinkela_wire_6638;
    wire new_Jinkela_wire_3889;
    wire new_Jinkela_wire_2728;
    wire new_Jinkela_wire_1989;
    wire new_Jinkela_wire_15246;
    wire new_Jinkela_wire_2948;
    wire new_Jinkela_wire_11775;
    wire new_Jinkela_wire_19786;
    wire new_Jinkela_wire_14719;
    wire new_Jinkela_wire_11575;
    wire new_Jinkela_wire_19200;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_17444;
    wire new_Jinkela_wire_12715;
    wire new_Jinkela_wire_18520;
    wire _0636_;
    wire new_Jinkela_wire_13224;
    wire new_Jinkela_wire_15226;
    wire _1375_;
    wire new_Jinkela_wire_9194;
    wire _0899_;
    wire new_Jinkela_wire_16091;
    wire new_Jinkela_wire_14578;
    wire _0461_;
    wire new_Jinkela_wire_13220;
    wire new_Jinkela_wire_3621;
    wire new_Jinkela_wire_1844;
    wire new_Jinkela_wire_14375;
    wire new_Jinkela_wire_1661;
    wire new_Jinkela_wire_9723;
    wire new_Jinkela_wire_16760;
    wire new_Jinkela_wire_17009;
    wire new_Jinkela_wire_77;
    wire _1388_;
    wire new_Jinkela_wire_13453;
    wire _0606_;
    wire new_Jinkela_wire_14900;
    wire new_Jinkela_wire_18581;
    wire new_Jinkela_wire_19163;
    wire new_Jinkela_wire_14726;
    wire new_Jinkela_wire_9322;
    wire new_Jinkela_wire_12795;
    wire new_Jinkela_wire_10720;
    wire new_Jinkela_wire_7742;
    wire new_Jinkela_wire_19799;
    wire new_Jinkela_wire_6985;
    wire new_Jinkela_wire_3686;
    wire new_Jinkela_wire_6008;
    wire new_Jinkela_wire_13273;
    wire new_Jinkela_wire_11593;
    wire new_Jinkela_wire_19016;
    wire new_Jinkela_wire_1815;
    wire new_Jinkela_wire_13331;
    wire new_Jinkela_wire_8221;
    wire _0809_;
    wire _0839_;
    wire new_Jinkela_wire_11546;
    wire new_Jinkela_wire_2319;
    wire new_Jinkela_wire_3557;
    wire new_Jinkela_wire_21237;
    wire new_Jinkela_wire_11444;
    wire new_Jinkela_wire_4705;
    wire new_Jinkela_wire_9204;
    wire new_Jinkela_wire_10339;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_12139;
    wire new_Jinkela_wire_4033;
    wire new_Jinkela_wire_9527;
    wire new_Jinkela_wire_1774;
    wire _1778_;
    wire new_Jinkela_wire_12710;
    wire new_Jinkela_wire_9292;
    wire new_Jinkela_wire_4101;
    wire new_Jinkela_wire_7066;
    wire new_Jinkela_wire_14241;
    wire new_Jinkela_wire_5854;
    wire new_Jinkela_wire_16386;
    wire new_Jinkela_wire_16413;
    wire new_Jinkela_wire_16600;
    wire new_Jinkela_wire_7005;
    wire new_Jinkela_wire_9623;
    wire new_Jinkela_wire_20495;
    wire new_Jinkela_wire_11558;
    wire new_Jinkela_wire_18301;
    wire _0449_;
    wire new_Jinkela_wire_8157;
    wire new_Jinkela_wire_15104;
    wire new_Jinkela_wire_8372;
    wire new_Jinkela_wire_15507;
    wire new_Jinkela_wire_18510;
    wire new_Jinkela_wire_4348;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_16398;
    wire new_Jinkela_wire_14137;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_14089;
    wire new_Jinkela_wire_10815;
    wire new_Jinkela_wire_18122;
    wire new_Jinkela_wire_17557;
    wire new_Jinkela_wire_14299;
    wire new_Jinkela_wire_19664;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_14066;
    wire new_Jinkela_wire_21083;
    wire new_Jinkela_wire_5354;
    wire _1655_;
    wire new_Jinkela_wire_17219;
    wire new_Jinkela_wire_11191;
    wire new_Jinkela_wire_11794;
    wire new_Jinkela_wire_15113;
    wire new_Jinkela_wire_14121;
    wire new_Jinkela_wire_9698;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_3119;
    wire new_Jinkela_wire_15755;
    wire new_Jinkela_wire_8077;
    wire new_Jinkela_wire_18784;
    wire new_Jinkela_wire_19322;
    wire new_Jinkela_wire_16046;
    wire new_Jinkela_wire_16299;
    wire new_Jinkela_wire_12763;
    wire new_Jinkela_wire_18135;
    wire new_Jinkela_wire_20979;
    wire new_Jinkela_wire_16746;
    wire new_Jinkela_wire_5750;
    wire new_Jinkela_wire_16140;
    wire new_Jinkela_wire_7251;
    wire new_Jinkela_wire_19535;
    wire new_Jinkela_wire_11292;
    wire new_Jinkela_wire_12517;
    wire _0270_;
    wire new_Jinkela_wire_1741;
    wire new_Jinkela_wire_4824;
    wire new_Jinkela_wire_3036;
    wire new_Jinkela_wire_5042;
    wire new_Jinkela_wire_7075;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_14254;
    wire new_Jinkela_wire_5060;
    wire new_Jinkela_wire_19585;
    wire new_Jinkela_wire_20354;
    wire new_Jinkela_wire_12232;
    wire new_Jinkela_wire_2243;
    wire new_Jinkela_wire_8386;
    wire new_Jinkela_wire_9375;
    wire _1107_;
    wire new_Jinkela_wire_18695;
    wire new_Jinkela_wire_12303;
    wire new_Jinkela_wire_12469;
    wire new_Jinkela_wire_14648;
    wire new_Jinkela_wire_12621;
    wire new_Jinkela_wire_17472;
    wire new_Jinkela_wire_4082;
    wire new_Jinkela_wire_16852;
    wire new_Jinkela_wire_3919;
    wire new_Jinkela_wire_10119;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_19615;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_7409;
    wire _1811_;
    wire new_Jinkela_wire_14583;
    wire new_Jinkela_wire_15069;
    wire new_Jinkela_wire_21201;
    wire new_Jinkela_wire_7355;
    wire new_Jinkela_wire_8158;
    wire new_Jinkela_wire_11943;
    wire new_Jinkela_wire_16343;
    wire _0854_;
    wire new_Jinkela_wire_12617;
    wire _0770_;
    wire new_Jinkela_wire_10401;
    wire new_Jinkela_wire_19104;
    wire new_Jinkela_wire_5299;
    wire new_Jinkela_wire_3363;
    wire new_Jinkela_wire_6064;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_17653;
    wire _1301_;
    wire new_Jinkela_wire_16977;
    wire new_Jinkela_wire_9950;
    wire _0477_;
    wire new_Jinkela_wire_19532;
    wire new_Jinkela_wire_11701;
    wire new_Jinkela_wire_3567;
    wire _0304_;
    wire new_Jinkela_wire_17898;
    wire new_Jinkela_wire_13042;
    wire new_Jinkela_wire_19105;
    wire new_Jinkela_wire_2264;
    wire new_Jinkela_wire_10320;
    wire new_Jinkela_wire_7352;
    wire new_Jinkela_wire_6898;
    wire _0287_;
    wire new_Jinkela_wire_18254;
    wire new_Jinkela_wire_5519;
    wire new_Jinkela_wire_9391;
    wire new_Jinkela_wire_13459;
    wire new_Jinkela_wire_6855;
    wire new_Jinkela_wire_15516;
    wire new_Jinkela_wire_18409;
    wire new_Jinkela_wire_14296;
    wire new_Jinkela_wire_5868;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_18894;
    wire new_Jinkela_wire_7957;
    wire new_Jinkela_wire_11001;
    wire new_Jinkela_wire_6659;
    wire new_Jinkela_wire_10356;
    wire _0510_;
    wire new_Jinkela_wire_6571;
    wire new_Jinkela_wire_12735;
    wire new_Jinkela_wire_7951;
    wire new_Jinkela_wire_15079;
    wire new_Jinkela_wire_5567;
    wire _0191_;
    wire new_Jinkela_wire_8208;
    wire new_Jinkela_wire_17610;
    wire new_Jinkela_wire_15707;
    wire new_Jinkela_wire_8985;
    wire new_Jinkela_wire_12568;
    wire new_Jinkela_wire_13347;
    wire new_Jinkela_wire_7116;
    wire new_Jinkela_wire_4887;
    wire new_Jinkela_wire_7268;
    wire _0088_;
    wire new_Jinkela_wire_3997;
    wire new_Jinkela_wire_18305;
    wire _0099_;
    wire _1038_;
    wire new_Jinkela_wire_8448;
    wire new_Jinkela_wire_14433;
    wire new_Jinkela_wire_17900;
    wire new_Jinkela_wire_17212;
    wire new_Jinkela_wire_2449;
    wire new_Jinkela_wire_2959;
    wire new_Jinkela_wire_11628;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_8333;
    wire new_Jinkela_wire_16623;
    wire new_Jinkela_wire_7714;
    wire new_Jinkela_wire_19973;
    wire new_Jinkela_wire_10089;
    wire new_Jinkela_wire_9994;
    wire new_Jinkela_wire_7257;
    wire new_Jinkela_wire_18068;
    wire new_Jinkela_wire_17414;
    wire new_Jinkela_wire_2802;
    wire new_Jinkela_wire_21117;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_11377;
    wire new_Jinkela_wire_11376;
    wire new_Jinkela_wire_7674;
    wire new_Jinkela_wire_11853;
    wire new_Jinkela_wire_3634;
    wire new_Jinkela_wire_8760;
    wire new_Jinkela_wire_6737;
    wire new_Jinkela_wire_12925;
    wire _0934_;
    wire new_Jinkela_wire_6193;
    wire new_Jinkela_wire_20997;
    wire new_Jinkela_wire_17016;
    wire new_Jinkela_wire_10367;
    wire new_Jinkela_wire_7919;
    wire new_Jinkela_wire_6170;
    wire new_Jinkela_wire_8269;
    wire new_Jinkela_wire_17430;
    wire new_Jinkela_wire_10851;
    wire new_Jinkela_wire_9696;
    wire new_Jinkela_wire_12627;
    wire new_Jinkela_wire_15047;
    wire new_Jinkela_wire_17441;
    wire new_Jinkela_wire_18749;
    wire new_Jinkela_wire_10322;
    wire new_Jinkela_wire_9402;
    wire new_Jinkela_wire_6116;
    wire new_Jinkela_wire_14180;
    wire new_Jinkela_wire_19802;
    wire new_Jinkela_wire_17340;
    wire new_Jinkela_wire_18747;
    wire new_Jinkela_wire_7189;
    wire new_Jinkela_wire_11748;
    wire _0254_;
    wire new_Jinkela_wire_11391;
    wire new_Jinkela_wire_8120;
    wire new_Jinkela_wire_19128;
    wire new_Jinkela_wire_7130;
    wire new_Jinkela_wire_21258;
    wire new_Jinkela_wire_10861;
    wire new_Jinkela_wire_5053;
    wire new_Jinkela_wire_4381;
    wire new_Jinkela_wire_8008;
    wire new_Jinkela_wire_2169;
    wire new_Jinkela_wire_19566;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_14678;
    wire new_Jinkela_wire_5307;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_16226;
    wire new_Jinkela_wire_10752;
    wire new_Jinkela_wire_19086;
    wire new_Jinkela_wire_17956;
    wire new_Jinkela_wire_10380;
    wire new_Jinkela_wire_9230;
    wire new_Jinkela_wire_20392;
    wire new_Jinkela_wire_15400;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_5065;
    wire new_Jinkela_wire_2574;
    wire new_Jinkela_wire_11888;
    wire new_Jinkela_wire_16999;
    wire _0498_;
    wire new_Jinkela_wire_6380;
    wire new_Jinkela_wire_20480;
    wire new_Jinkela_wire_15045;
    wire new_Jinkela_wire_9026;
    wire new_Jinkela_wire_2294;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_3368;
    wire _1821_;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_15783;
    wire new_Jinkela_wire_19026;
    wire new_Jinkela_wire_11308;
    wire new_Jinkela_wire_6656;
    wire new_Jinkela_wire_10771;
    wire new_Jinkela_wire_16533;
    wire new_Jinkela_wire_19261;
    wire new_Jinkela_wire_11170;
    wire new_Jinkela_wire_15237;
    wire new_Jinkela_wire_15964;
    wire _1546_;
    wire new_Jinkela_wire_4049;
    wire new_Jinkela_wire_2867;
    wire new_Jinkela_wire_11485;
    wire new_Jinkela_wire_20470;
    wire _1830_;
    wire new_Jinkela_wire_9173;
    wire new_Jinkela_wire_14095;
    wire new_Jinkela_wire_7816;
    wire new_Jinkela_wire_3584;
    wire new_Jinkela_wire_8379;
    wire new_Jinkela_wire_11105;
    wire new_Jinkela_wire_6117;
    wire new_Jinkela_wire_15668;
    wire new_Jinkela_wire_18737;
    wire new_Jinkela_wire_1911;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_7876;
    wire new_Jinkela_wire_10433;
    wire new_Jinkela_wire_19957;
    wire new_Jinkela_wire_13795;
    wire new_Jinkela_wire_20666;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_20286;
    wire new_Jinkela_wire_19117;
    wire new_Jinkela_wire_4198;
    wire new_Jinkela_wire_6995;
    wire new_Jinkela_wire_12125;
    wire new_Jinkela_wire_14843;
    wire new_Jinkela_wire_2038;
    wire new_Jinkela_wire_6006;
    wire new_Jinkela_wire_6527;
    wire new_Jinkela_wire_13336;
    wire new_Jinkela_wire_9659;
    wire new_Jinkela_wire_13561;
    wire new_Jinkela_wire_21190;
    wire new_Jinkela_wire_10697;
    wire new_Jinkela_wire_4062;
    wire new_Jinkela_wire_12537;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_17914;
    wire new_Jinkela_wire_9607;
    wire new_Jinkela_wire_18600;
    wire new_Jinkela_wire_19120;
    wire new_Jinkela_wire_14177;
    wire new_Jinkela_wire_5929;
    wire new_Jinkela_wire_13288;
    wire new_Jinkela_wire_16518;
    wire new_Jinkela_wire_20894;
    wire new_Jinkela_wire_8494;
    wire _0995_;
    wire new_Jinkela_wire_15782;
    wire new_Jinkela_wire_18472;
    wire new_Jinkela_wire_17504;
    wire _0286_;
    wire _0178_;
    wire new_Jinkela_wire_10127;
    wire _0740_;
    wire new_Jinkela_wire_11839;
    wire new_Jinkela_wire_12536;
    wire new_Jinkela_wire_9699;
    wire new_Jinkela_wire_9314;
    wire new_Jinkela_wire_13975;
    wire new_Jinkela_wire_2087;
    wire new_Jinkela_wire_21298;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_13377;
    wire new_Jinkela_wire_9477;
    wire new_Jinkela_wire_15976;
    wire new_Jinkela_wire_19895;
    wire new_Jinkela_wire_9693;
    wire new_Jinkela_wire_7566;
    wire new_Jinkela_wire_6560;
    wire new_Jinkela_wire_13828;
    wire new_Jinkela_wire_3786;
    wire _0489_;
    wire new_Jinkela_wire_14125;
    wire new_Jinkela_wire_16841;
    wire new_Jinkela_wire_9895;
    wire new_Jinkela_wire_6305;
    wire new_Jinkela_wire_3228;
    wire new_Jinkela_wire_15088;
    wire new_Jinkela_wire_5358;
    wire new_Jinkela_wire_11721;
    wire new_Jinkela_wire_15161;
    wire new_Jinkela_wire_18434;
    wire new_Jinkela_wire_12699;
    wire new_Jinkela_wire_9755;
    wire new_Jinkela_wire_12475;
    wire new_Jinkela_wire_12913;
    wire new_Jinkela_wire_15861;
    wire new_Jinkela_wire_11435;
    wire new_Jinkela_wire_20665;
    wire new_Jinkela_wire_3423;
    wire new_Jinkela_wire_14356;
    wire new_Jinkela_wire_20537;
    wire new_Jinkela_wire_9443;
    wire new_Jinkela_wire_14566;
    wire new_Jinkela_wire_11686;
    wire new_Jinkela_wire_12624;
    wire new_Jinkela_wire_10849;
    wire new_Jinkela_wire_18930;
    wire new_Jinkela_wire_12761;
    wire new_Jinkela_wire_5054;
    wire new_Jinkela_wire_18945;
    wire new_Jinkela_wire_8719;
    wire new_Jinkela_wire_3647;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_8832;
    wire new_Jinkela_wire_9854;
    wire new_Jinkela_wire_2587;
    wire new_Jinkela_wire_10024;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_20793;
    wire new_Jinkela_wire_21322;
    wire new_Jinkela_wire_18598;
    wire _1796_;
    wire new_Jinkela_wire_14167;
    wire new_Jinkela_wire_2642;
    wire new_Jinkela_wire_11198;
    wire new_Jinkela_wire_5376;
    wire new_Jinkela_wire_4412;
    wire new_Jinkela_wire_20994;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_10839;
    wire new_Jinkela_wire_17255;
    wire new_Jinkela_wire_4575;
    wire new_Jinkela_wire_4196;
    wire new_Jinkela_wire_19166;
    wire new_Jinkela_wire_14306;
    wire new_Jinkela_wire_7503;
    wire new_Jinkela_wire_18043;
    wire new_Jinkela_wire_14634;
    wire new_Jinkela_wire_2347;
    wire new_Jinkela_wire_5239;
    wire new_Jinkela_wire_14551;
    wire new_Jinkela_wire_4401;
    wire new_Jinkela_wire_16772;
    wire new_Jinkela_wire_4266;
    wire new_Jinkela_wire_10545;
    wire new_Jinkela_wire_5269;
    wire new_Jinkela_wire_15864;
    wire new_Jinkela_wire_21065;
    wire new_Jinkela_wire_14916;
    wire new_Jinkela_wire_20097;
    wire new_Jinkela_wire_20075;
    wire new_Jinkela_wire_6347;
    wire new_Jinkela_wire_7553;
    wire _0679_;
    wire new_Jinkela_wire_19745;
    wire new_Jinkela_wire_12437;
    wire new_Jinkela_wire_8501;
    wire new_Jinkela_wire_12153;
    wire new_Jinkela_wire_10888;
    wire new_Jinkela_wire_18098;
    wire new_Jinkela_wire_8114;
    wire new_Jinkela_wire_3841;
    wire _0681_;
    wire new_Jinkela_wire_16587;
    wire new_Jinkela_wire_13956;
    wire new_Jinkela_wire_20151;
    wire new_Jinkela_wire_10721;
    wire _1245_;
    wire new_Jinkela_wire_10580;
    wire new_Jinkela_wire_19448;
    wire new_Jinkela_wire_11689;
    wire new_Jinkela_wire_2281;
    wire new_Jinkela_wire_3530;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_7908;
    wire new_Jinkela_wire_19752;
    wire new_Jinkela_wire_13694;
    wire new_Jinkela_wire_5586;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_7563;
    wire _0614_;
    wire new_Jinkela_wire_9405;
    wire new_Jinkela_wire_3711;
    wire new_Jinkela_wire_4664;
    wire new_Jinkela_wire_2890;
    wire new_Jinkela_wire_16767;
    wire new_Jinkela_wire_6384;
    wire new_Jinkela_wire_5857;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_6253;
    wire new_Jinkela_wire_17373;
    wire new_Jinkela_wire_11205;
    wire new_Jinkela_wire_6327;
    wire new_Jinkela_wire_18718;
    wire new_Jinkela_wire_12032;
    wire new_Jinkela_wire_6556;
    wire new_Jinkela_wire_14199;
    wire _1502_;
    wire new_Jinkela_wire_19639;
    wire new_Jinkela_wire_5430;
    wire new_Jinkela_wire_13089;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_20514;
    wire _0397_;
    wire new_Jinkela_wire_6285;
    wire new_Jinkela_wire_13746;
    wire new_Jinkela_wire_16535;
    wire _0023_;
    wire new_Jinkela_wire_18524;
    wire new_Jinkela_wire_14290;
    wire new_Jinkela_wire_20270;
    wire new_Jinkela_wire_11933;
    wire new_Jinkela_wire_19216;
    wire new_Jinkela_wire_14170;
    wire new_Jinkela_wire_19785;
    wire new_Jinkela_wire_5404;
    wire new_Jinkela_wire_13158;
    wire new_Jinkela_wire_10058;
    wire new_Jinkela_wire_18729;
    wire new_Jinkela_wire_14869;
    wire new_Jinkela_wire_18325;
    wire _1296_;
    wire new_Jinkela_wire_17906;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_7091;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_15165;
    wire new_Jinkela_wire_12526;
    wire _1015_;
    wire new_Jinkela_wire_19254;
    wire new_Jinkela_wire_7282;
    wire new_Jinkela_wire_19304;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_16083;
    wire new_Jinkela_wire_19793;
    wire new_Jinkela_wire_2766;
    wire new_Jinkela_wire_9528;
    wire new_Jinkela_wire_11557;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_20921;
    wire new_Jinkela_wire_20505;
    wire new_Jinkela_wire_7478;
    wire new_Jinkela_wire_10690;
    wire new_Jinkela_wire_3365;
    wire new_Jinkela_wire_9305;
    wire new_Jinkela_wire_15750;
    wire new_Jinkela_wire_19267;
    wire new_Jinkela_wire_6432;
    wire new_Jinkela_wire_18261;
    wire new_Jinkela_wire_17313;
    wire new_Jinkela_wire_5130;
    wire new_Jinkela_wire_9936;
    wire new_Jinkela_wire_15366;
    wire _0550_;
    wire _1141_;
    wire new_Jinkela_wire_9159;
    wire new_Jinkela_wire_5721;
    wire new_Jinkela_wire_8989;
    wire new_Jinkela_wire_5083;
    wire _0737_;
    wire new_Jinkela_wire_15051;
    wire new_Jinkela_wire_8797;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_18054;
    wire new_Jinkela_wire_17831;
    wire new_Jinkela_wire_13475;
    wire new_Jinkela_wire_11703;
    wire new_Jinkela_wire_6224;
    wire new_Jinkela_wire_1384;
    wire _1182_;
    wire new_Jinkela_wire_20504;
    wire new_Jinkela_wire_13161;
    wire new_Jinkela_wire_6669;
    wire new_Jinkela_wire_6244;
    wire new_Jinkela_wire_17632;
    wire new_Jinkela_wire_19643;
    wire new_Jinkela_wire_6186;
    wire new_Jinkela_wire_13620;
    wire new_Jinkela_wire_2583;
    wire new_Jinkela_wire_7590;
    wire new_Jinkela_wire_8592;
    wire new_Jinkela_wire_19053;
    wire new_Jinkela_wire_8318;
    wire new_Jinkela_wire_7428;
    wire new_Jinkela_wire_2429;
    wire new_Jinkela_wire_8028;
    wire _0385_;
    wire new_Jinkela_wire_6658;
    wire new_Jinkela_wire_9117;
    wire new_Jinkela_wire_11681;
    wire new_Jinkela_wire_16315;
    wire new_Jinkela_wire_19339;
    wire new_Jinkela_wire_15875;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_11587;
    wire new_Jinkela_wire_17723;
    wire new_Jinkela_wire_13525;
    wire _0797_;
    wire new_Jinkela_wire_3783;
    wire new_Jinkela_wire_11052;
    wire new_Jinkela_wire_15402;
    wire new_Jinkela_wire_19837;
    wire _1411_;
    wire _1162_;
    wire new_Jinkela_wire_19599;
    wire new_Jinkela_wire_17602;
    wire new_Jinkela_wire_5238;
    wire new_Jinkela_wire_5640;
    wire _1170_;
    wire new_Jinkela_wire_17124;
    wire new_Jinkela_wire_18950;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_3414;
    wire _0198_;
    wire _1807_;
    wire new_Jinkela_wire_20858;
    wire _0359_;
    wire new_Jinkela_wire_13405;
    wire new_Jinkela_wire_698;
    wire _0077_;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_2299;
    wire _0987_;
    wire new_Jinkela_wire_5259;
    wire new_Jinkela_wire_4486;
    wire _0713_;
    wire new_Jinkela_wire_5777;
    wire new_Jinkela_wire_12985;
    wire new_Jinkela_wire_19145;
    wire new_Jinkela_wire_8328;
    wire new_net_3966;
    wire new_Jinkela_wire_13230;
    wire new_Jinkela_wire_7454;
    wire new_net_3962;
    wire _1757_;
    wire new_Jinkela_wire_17870;
    wire new_Jinkela_wire_18595;
    wire new_Jinkela_wire_20030;
    wire new_Jinkela_wire_9761;
    wire _0758_;
    wire new_Jinkela_wire_10077;
    wire new_Jinkela_wire_16276;
    wire new_Jinkela_wire_15898;
    wire new_Jinkela_wire_18061;
    wire new_Jinkela_wire_2998;
    wire new_Jinkela_wire_7732;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_3978;
    wire new_Jinkela_wire_21214;
    wire new_Jinkela_wire_19294;
    wire new_Jinkela_wire_10519;
    wire new_Jinkela_wire_13242;
    wire new_Jinkela_wire_11431;
    wire new_Jinkela_wire_17241;
    wire new_Jinkela_wire_17565;
    wire new_Jinkela_wire_18248;
    wire new_Jinkela_wire_21135;
    wire new_Jinkela_wire_12443;
    wire new_Jinkela_wire_2538;
    wire new_Jinkela_wire_15574;
    wire new_Jinkela_wire_16528;
    wire new_Jinkela_wire_16136;
    wire new_Jinkela_wire_6596;
    wire new_Jinkela_wire_2540;
    wire new_Jinkela_wire_19084;
    wire new_Jinkela_wire_8663;
    wire _0400_;
    wire new_Jinkela_wire_14571;
    wire new_Jinkela_wire_14183;
    wire new_Jinkela_wire_19715;
    wire _1497_;
    wire new_Jinkela_wire_15180;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_6818;
    wire new_Jinkela_wire_4809;
    wire _1214_;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_10668;
    wire new_Jinkela_wire_15564;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_18015;
    wire new_Jinkela_wire_7217;
    wire new_Jinkela_wire_12001;
    wire _1217_;
    wire new_Jinkela_wire_15935;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_2708;
    wire new_Jinkela_wire_7790;
    wire new_Jinkela_wire_3506;
    wire _0421_;
    wire new_Jinkela_wire_18854;
    wire new_Jinkela_wire_13059;
    wire new_Jinkela_wire_4151;
    wire new_Jinkela_wire_11455;
    wire new_Jinkela_wire_10879;
    wire new_Jinkela_wire_19661;
    wire new_Jinkela_wire_8839;
    wire _0368_;
    wire new_Jinkela_wire_6979;
    wire new_Jinkela_wire_16769;
    wire new_Jinkela_wire_13720;
    wire new_Jinkela_wire_6521;
    wire new_Jinkela_wire_3679;
    wire new_Jinkela_wire_5536;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_19863;
    wire new_Jinkela_wire_3188;
    wire new_Jinkela_wire_3081;
    wire new_Jinkela_wire_18873;
    wire _0465_;
    wire new_Jinkela_wire_3456;
    wire new_Jinkela_wire_11974;
    wire new_Jinkela_wire_18034;
    wire new_Jinkela_wire_11750;
    wire new_Jinkela_wire_13296;
    wire new_Jinkela_wire_16712;
    wire new_Jinkela_wire_12700;
    wire new_Jinkela_wire_19556;
    wire new_Jinkela_wire_5844;
    wire new_Jinkela_wire_4376;
    wire new_Jinkela_wire_7117;
    wire new_Jinkela_wire_9714;
    wire new_Jinkela_wire_14994;
    wire new_Jinkela_wire_2645;
    wire new_Jinkela_wire_16644;
    wire new_Jinkela_wire_8272;
    wire new_Jinkela_wire_20422;
    wire new_Jinkela_wire_16718;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_20277;
    wire new_Jinkela_wire_16713;
    wire new_Jinkela_wire_12225;
    wire new_Jinkela_wire_13270;
    wire new_Jinkela_wire_19916;
    wire new_Jinkela_wire_16943;
    wire new_Jinkela_wire_2879;
    wire new_Jinkela_wire_6042;
    wire new_Jinkela_wire_14817;
    wire new_Jinkela_wire_18133;
    wire new_Jinkela_wire_2359;
    wire new_Jinkela_wire_4777;
    wire new_Jinkela_wire_21078;
    wire new_Jinkela_wire_9476;
    wire new_Jinkela_wire_4265;
    wire new_Jinkela_wire_7651;
    wire new_Jinkela_wire_2065;
    wire new_Jinkela_wire_14600;
    wire new_Jinkela_wire_8251;
    wire new_Jinkela_wire_20083;
    wire new_Jinkela_wire_5194;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_20364;
    wire _0967_;
    wire new_Jinkela_wire_4885;
    wire new_Jinkela_wire_12440;
    wire new_Jinkela_wire_12968;
    wire new_Jinkela_wire_17066;
    wire new_Jinkela_wire_19095;
    wire new_Jinkela_wire_21217;
    wire new_Jinkela_wire_19731;
    wire new_Jinkela_wire_6377;
    wire new_Jinkela_wire_11460;
    wire new_Jinkela_wire_8313;
    wire new_Jinkela_wire_4309;
    wire _1291_;
    wire new_Jinkela_wire_20230;
    wire new_Jinkela_wire_3513;
    wire new_Jinkela_wire_16094;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_19080;
    wire new_Jinkela_wire_20438;
    wire new_Jinkela_wire_8701;
    wire new_Jinkela_wire_11610;
    wire new_Jinkela_wire_12490;
    wire new_Jinkela_wire_12063;
    wire _1740_;
    wire new_Jinkela_wire_18613;
    wire new_Jinkela_wire_17705;
    wire new_Jinkela_wire_2680;
    wire new_Jinkela_wire_6821;
    wire new_Jinkela_wire_13286;
    wire new_Jinkela_wire_9074;
    wire new_Jinkela_wire_13567;
    wire new_Jinkela_wire_12013;
    wire new_Jinkela_wire_9584;
    wire _0456_;
    wire new_Jinkela_wire_16974;
    wire new_Jinkela_wire_20528;
    wire new_Jinkela_wire_7619;
    wire new_Jinkela_wire_12566;
    wire new_Jinkela_wire_14931;
    wire new_Jinkela_wire_8773;
    wire new_Jinkela_wire_19897;
    wire new_Jinkela_wire_17399;
    wire _1494_;
    wire new_Jinkela_wire_4591;
    wire new_Jinkela_wire_14178;
    wire _1278_;
    wire new_Jinkela_wire_15866;
    wire new_Jinkela_wire_3275;
    wire new_Jinkela_wire_7137;
    wire new_Jinkela_wire_13759;
    wire new_Jinkela_wire_19131;
    wire new_Jinkela_wire_12514;
    wire new_Jinkela_wire_14982;
    wire new_Jinkela_wire_2698;
    wire _0617_;
    wire new_Jinkela_wire_4213;
    wire new_Jinkela_wire_6779;
    wire new_Jinkela_wire_9718;
    wire new_Jinkela_wire_13897;
    wire new_Jinkela_wire_13228;
    wire new_Jinkela_wire_7335;
    wire new_Jinkela_wire_9064;
    wire new_Jinkela_wire_19390;
    wire new_Jinkela_wire_5945;
    wire new_Jinkela_wire_20325;
    wire new_Jinkela_wire_17371;
    wire new_Jinkela_wire_8604;
    wire new_Jinkela_wire_18642;
    wire new_Jinkela_wire_15933;
    wire new_Jinkela_wire_9294;
    wire new_Jinkela_wire_3943;
    wire new_Jinkela_wire_17498;
    wire new_Jinkela_wire_3721;
    wire new_Jinkela_wire_15124;
    wire new_Jinkela_wire_19922;
    wire new_Jinkela_wire_17052;
    wire new_Jinkela_wire_9241;
    wire new_Jinkela_wire_1788;
    wire new_Jinkela_wire_16698;
    wire new_Jinkela_wire_8167;
    wire new_Jinkela_wire_13276;
    wire new_Jinkela_wire_2444;
    wire new_Jinkela_wire_5291;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_2441;
    wire new_Jinkela_wire_7464;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_14206;
    wire new_Jinkela_wire_5986;
    wire new_Jinkela_wire_12609;
    wire new_Jinkela_wire_7007;
    wire new_Jinkela_wire_12929;
    wire new_Jinkela_wire_6644;
    wire new_Jinkela_wire_20020;
    wire new_Jinkela_wire_11816;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_9280;
    wire new_Jinkela_wire_20259;
    wire new_Jinkela_wire_19491;
    wire new_Jinkela_wire_2518;
    wire new_Jinkela_wire_8428;
    wire _1682_;
    wire new_Jinkela_wire_7232;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_8246;
    wire new_Jinkela_wire_13844;
    wire new_Jinkela_wire_15141;
    wire new_Jinkela_wire_20195;
    wire new_Jinkela_wire_6491;
    wire _1406_;
    wire _1470_;
    wire new_Jinkela_wire_19603;
    wire new_Jinkela_wire_10407;
    wire new_Jinkela_wire_6227;
    wire new_Jinkela_wire_15566;
    wire new_Jinkela_wire_4565;
    wire new_Jinkela_wire_4218;
    wire new_Jinkela_wire_20731;
    wire new_Jinkela_wire_10249;
    wire new_Jinkela_wire_1072;
    wire _0577_;
    wire _0849_;
    wire new_Jinkela_wire_14764;
    wire new_Jinkela_wire_9165;
    wire new_Jinkela_wire_15539;
    wire new_Jinkela_wire_4919;
    wire new_Jinkela_wire_5631;
    wire new_Jinkela_wire_16097;
    wire new_Jinkela_wire_19489;
    wire new_Jinkela_wire_11439;
    wire new_Jinkela_wire_15602;
    wire new_Jinkela_wire_2412;
    wire new_Jinkela_wire_10994;
    wire new_Jinkela_wire_8768;
    wire new_Jinkela_wire_15136;
    wire new_Jinkela_wire_19342;
    wire new_Jinkela_wire_10212;
    wire new_Jinkela_wire_17651;
    wire new_Jinkela_wire_20849;
    wire _0143_;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_1771;
    wire new_Jinkela_wire_19576;
    wire new_Jinkela_wire_16023;
    wire new_Jinkela_wire_2338;
    wire new_Jinkela_wire_2604;
    wire new_Jinkela_wire_8027;
    wire new_Jinkela_wire_20857;
    wire new_Jinkela_wire_11704;
    wire new_Jinkela_wire_11578;
    wire new_Jinkela_wire_17135;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_3987;
    wire new_Jinkela_wire_13851;
    wire _0536_;
    wire new_Jinkela_wire_16269;
    wire new_Jinkela_wire_9411;
    wire new_Jinkela_wire_2937;
    wire new_Jinkela_wire_17380;
    wire new_Jinkela_wire_11384;
    wire new_Jinkela_wire_19606;
    wire new_Jinkela_wire_14570;
    wire new_Jinkela_wire_5261;
    wire new_Jinkela_wire_14156;
    wire _1829_;
    wire new_Jinkela_wire_10906;
    wire new_Jinkela_wire_17069;
    wire new_Jinkela_wire_9947;
    wire new_Jinkela_wire_12808;
    wire new_Jinkela_wire_19156;
    wire new_Jinkela_wire_20313;
    wire new_Jinkela_wire_19994;
    wire _0493_;
    wire new_Jinkela_wire_9030;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_2274;
    wire new_Jinkela_wire_5490;
    wire new_Jinkela_wire_7730;
    wire new_Jinkela_wire_18358;
    wire new_Jinkela_wire_12266;
    wire new_Jinkela_wire_13580;
    wire _0618_;
    wire new_Jinkela_wire_5732;
    wire new_Jinkela_wire_18095;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_5827;
    wire new_Jinkela_wire_14868;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_6089;
    wire new_Jinkela_wire_17025;
    wire new_Jinkela_wire_1872;
    wire new_Jinkela_wire_18859;
    wire new_Jinkela_wire_21185;
    wire new_Jinkela_wire_16903;
    wire new_Jinkela_wire_1969;
    wire _0073_;
    wire new_Jinkela_wire_16293;
    wire new_Jinkela_wire_18339;
    wire new_Jinkela_wire_11504;
    wire new_Jinkela_wire_6222;
    wire new_Jinkela_wire_10170;
    wire new_Jinkela_wire_15291;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_6494;
    wire new_Jinkela_wire_10649;
    wire new_Jinkela_wire_17836;
    wire new_Jinkela_wire_16428;
    wire new_Jinkela_wire_21158;
    wire _0443_;
    wire new_Jinkela_wire_14525;
    wire new_Jinkela_wire_20634;
    wire new_Jinkela_wire_6172;
    wire new_Jinkela_wire_15518;
    wire new_Jinkela_wire_15631;
    wire new_Jinkela_wire_11550;
    wire new_Jinkela_wire_10428;
    wire new_Jinkela_wire_14852;
    wire new_Jinkela_wire_5003;
    wire new_Jinkela_wire_9724;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_4492;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_21194;
    wire new_Jinkela_wire_2776;
    wire new_Jinkela_wire_19734;
    wire new_Jinkela_wire_17713;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_3970;
    wire new_Jinkela_wire_17985;
    wire new_Jinkela_wire_7498;
    wire new_Jinkela_wire_13680;
    wire new_Jinkela_wire_5388;
    wire new_Jinkela_wire_19952;
    wire new_Jinkela_wire_2600;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_7212;
    wire _1171_;
    wire new_Jinkela_wire_21136;
    wire new_Jinkela_wire_18895;
    wire new_Jinkela_wire_7334;
    wire new_Jinkela_wire_3903;
    wire new_Jinkela_wire_13182;
    wire new_Jinkela_wire_9068;
    wire new_Jinkela_wire_5462;
    wire new_Jinkela_wire_7855;
    wire new_Jinkela_wire_6875;
    wire new_Jinkela_wire_5400;
    wire new_Jinkela_wire_16072;
    wire new_Jinkela_wire_5549;
    wire new_Jinkela_wire_7023;
    wire new_Jinkela_wire_8758;
    wire new_Jinkela_wire_16064;
    wire new_Jinkela_wire_7231;
    wire new_Jinkela_wire_8431;
    wire new_Jinkela_wire_9100;
    wire new_Jinkela_wire_1867;
    wire new_Jinkela_wire_15704;
    wire new_Jinkela_wire_3327;
    wire new_Jinkela_wire_20114;
    wire new_Jinkela_wire_17794;
    wire new_Jinkela_wire_17501;
    wire new_Jinkela_wire_11179;
    wire new_Jinkela_wire_17179;
    wire _0323_;
    wire new_Jinkela_wire_6937;
    wire new_Jinkela_wire_10624;
    wire new_Jinkela_wire_16280;
    wire new_Jinkela_wire_20907;
    wire new_Jinkela_wire_20986;
    wire new_Jinkela_wire_11656;
    wire _1168_;
    wire new_Jinkela_wire_5115;
    wire new_Jinkela_wire_14891;
    wire new_Jinkela_wire_20002;
    wire new_Jinkela_wire_6803;
    wire new_Jinkela_wire_19549;
    wire new_Jinkela_wire_20644;
    wire new_Jinkela_wire_19983;
    wire new_Jinkela_wire_12602;
    wire new_Jinkela_wire_20982;
    wire new_Jinkela_wire_15936;
    wire new_Jinkela_wire_10526;
    wire new_Jinkela_wire_8569;
    wire new_Jinkela_wire_4580;
    wire new_Jinkela_wire_13603;
    wire new_Jinkela_wire_18473;
    wire new_Jinkela_wire_13484;
    wire new_Jinkela_wire_17746;
    wire new_Jinkela_wire_6614;
    wire new_Jinkela_wire_6953;
    wire new_Jinkela_wire_8599;
    wire new_Jinkela_wire_6870;
    wire new_Jinkela_wire_14488;
    wire new_Jinkela_wire_4425;
    wire new_Jinkela_wire_4765;
    wire new_Jinkela_wire_9672;
    wire new_Jinkela_wire_7396;
    wire new_Jinkela_wire_10530;
    wire new_Jinkela_wire_3448;
    wire new_Jinkela_wire_14025;
    wire new_Jinkela_wire_5898;
    wire new_Jinkela_wire_3572;
    wire new_Jinkela_wire_18262;
    wire new_Jinkela_wire_20186;
    wire new_Jinkela_wire_20946;
    wire new_Jinkela_wire_2791;
    wire _1089_;
    wire new_Jinkela_wire_17118;
    wire new_Jinkela_wire_4920;
    wire _0747_;
    wire new_Jinkela_wire_14856;
    wire new_Jinkela_wire_8097;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_10454;
    wire new_net_3958;
    wire new_Jinkela_wire_10602;
    wire new_Jinkela_wire_9785;
    wire new_Jinkela_wire_17951;
    wire new_Jinkela_wire_13362;
    wire new_net_3924;
    wire new_Jinkela_wire_2855;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_7042;
    wire new_Jinkela_wire_7077;
    wire new_Jinkela_wire_6124;
    wire new_Jinkela_wire_18620;
    wire new_Jinkela_wire_2160;
    wire new_Jinkela_wire_18341;
    wire new_Jinkela_wire_16259;
    wire new_Jinkela_wire_8211;
    wire new_Jinkela_wire_19847;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_9056;
    wire new_Jinkela_wire_8199;
    wire new_Jinkela_wire_6586;
    wire new_Jinkela_wire_5974;
    wire new_Jinkela_wire_19325;
    wire new_Jinkela_wire_13421;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_7398;
    wire new_Jinkela_wire_20736;
    wire new_Jinkela_wire_3362;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_3907;
    wire new_Jinkela_wire_10744;
    wire new_Jinkela_wire_8479;
    wire new_Jinkela_wire_21315;
    wire new_Jinkela_wire_9390;
    wire new_Jinkela_wire_2545;
    wire new_Jinkela_wire_9046;
    wire new_Jinkela_wire_21162;
    wire new_Jinkela_wire_9982;
    wire _0223_;
    wire new_Jinkela_wire_19540;
    wire new_Jinkela_wire_12386;
    wire new_Jinkela_wire_9832;
    wire new_Jinkela_wire_7385;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_15572;
    wire new_Jinkela_wire_7764;
    wire new_Jinkela_wire_6924;
    wire new_Jinkela_wire_12661;
    wire new_Jinkela_wire_7168;
    wire new_Jinkela_wire_21180;
    wire new_Jinkela_wire_5647;
    wire new_Jinkela_wire_3874;
    wire new_Jinkela_wire_19878;
    wire new_Jinkela_wire_20260;
    wire new_net_3960;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_10110;
    wire new_Jinkela_wire_19776;
    wire new_Jinkela_wire_11140;
    wire new_Jinkela_wire_3905;
    wire new_Jinkela_wire_14038;
    wire new_Jinkela_wire_14921;
    wire new_Jinkela_wire_13703;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_3739;
    wire new_Jinkela_wire_15931;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_7857;
    wire new_Jinkela_wire_18559;
    wire new_Jinkela_wire_14124;
    wire new_Jinkela_wire_3483;
    wire new_Jinkela_wire_3867;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_18820;
    wire new_Jinkela_wire_14717;
    wire new_Jinkela_wire_11154;
    wire new_Jinkela_wire_1445;
    wire _0553_;
    wire new_Jinkela_wire_8341;
    wire new_Jinkela_wire_12112;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_20544;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_15496;
    wire new_Jinkela_wire_10842;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_6588;
    wire new_Jinkela_wire_16552;
    wire new_Jinkela_wire_18842;
    wire new_Jinkela_wire_5381;
    wire new_Jinkela_wire_19686;
    wire new_Jinkela_wire_13854;
    wire new_Jinkela_wire_3853;
    wire new_Jinkela_wire_9306;
    wire _1408_;
    wire new_Jinkela_wire_12770;
    wire new_Jinkela_wire_12686;
    wire new_Jinkela_wire_2550;
    wire new_Jinkela_wire_12098;
    wire new_Jinkela_wire_7628;
    wire new_Jinkela_wire_20136;
    wire new_Jinkela_wire_8357;
    wire new_Jinkela_wire_8810;
    wire _1399_;
    wire new_Jinkela_wire_6856;
    wire new_Jinkela_wire_3313;
    wire _0296_;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_7555;
    wire new_Jinkela_wire_12022;
    wire new_Jinkela_wire_11097;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_17993;
    wire new_Jinkela_wire_12435;
    wire new_Jinkela_wire_14505;
    wire new_Jinkela_wire_9151;
    wire new_Jinkela_wire_12853;
    wire new_Jinkela_wire_8655;
    wire new_Jinkela_wire_17327;
    wire new_Jinkela_wire_4252;
    wire new_Jinkela_wire_18117;
    wire new_Jinkela_wire_13961;
    wire new_Jinkela_wire_6895;
    wire new_Jinkela_wire_14339;
    wire new_Jinkela_wire_18253;
    wire new_Jinkela_wire_5166;
    wire new_Jinkela_wire_17436;
    wire new_Jinkela_wire_3079;
    wire _0686_;
    wire new_Jinkela_wire_8202;
    wire new_Jinkela_wire_14400;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_20673;
    wire new_Jinkela_wire_2788;
    wire _1625_;
    wire new_Jinkela_wire_13446;
    wire new_Jinkela_wire_8650;
    wire new_Jinkela_wire_6802;
    wire new_Jinkela_wire_3828;
    wire new_Jinkela_wire_3958;
    wire new_Jinkela_wire_18494;
    wire new_Jinkela_wire_7531;
    wire new_Jinkela_wire_3294;
    wire new_Jinkela_wire_18526;
    wire new_Jinkela_wire_20016;
    wire new_Jinkela_wire_13460;
    wire new_Jinkela_wire_20234;
    wire new_Jinkela_wire_6530;
    wire new_Jinkela_wire_19115;
    wire new_Jinkela_wire_4600;
    wire new_Jinkela_wire_6466;
    wire new_Jinkela_wire_17194;
    wire new_Jinkela_wire_17552;
    wire new_Jinkela_wire_372;
    wire new_Jinkela_wire_5070;
    wire _0329_;
    wire new_Jinkela_wire_11904;
    wire new_Jinkela_wire_6983;
    wire new_Jinkela_wire_2295;
    wire new_Jinkela_wire_3859;
    wire new_Jinkela_wire_8023;
    wire new_Jinkela_wire_4452;
    wire new_Jinkela_wire_5225;
    wire new_Jinkela_wire_7815;
    wire new_Jinkela_wire_7008;
    wire new_Jinkela_wire_6931;
    wire new_Jinkela_wire_13178;
    wire new_Jinkela_wire_7200;
    wire new_Jinkela_wire_2588;
    wire new_Jinkela_wire_5904;
    wire new_Jinkela_wire_7490;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_18604;
    wire new_Jinkela_wire_13880;
    wire new_Jinkela_wire_2597;
    wire new_Jinkela_wire_1233;
    wire _1103_;
    wire new_Jinkela_wire_10827;
    wire new_Jinkela_wire_9036;
    wire new_Jinkela_wire_12424;
    wire new_Jinkela_wire_3304;
    wire new_Jinkela_wire_8616;
    wire new_Jinkela_wire_16675;
    wire new_Jinkela_wire_4884;
    wire new_Jinkela_wire_4731;
    wire new_Jinkela_wire_6826;
    wire new_Jinkela_wire_4067;
    wire new_Jinkela_wire_2697;
    wire new_Jinkela_wire_5434;
    wire new_Jinkela_wire_2313;
    wire new_Jinkela_wire_2979;
    wire _1797_;
    wire new_Jinkela_wire_10509;
    wire new_Jinkela_wire_10844;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_10157;
    wire new_Jinkela_wire_7386;
    wire new_Jinkela_wire_15509;
    wire new_Jinkela_wire_3166;
    wire new_Jinkela_wire_13061;
    wire new_Jinkela_wire_7049;
    wire new_Jinkela_wire_5161;
    wire _0389_;
    wire new_Jinkela_wire_4835;
    wire new_Jinkela_wire_21242;
    wire new_Jinkela_wire_2688;
    wire new_Jinkela_wire_5705;
    wire new_Jinkela_wire_9323;
    wire new_Jinkela_wire_11169;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_12123;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_9257;
    wire new_Jinkela_wire_12447;
    wire new_Jinkela_wire_11624;
    wire new_Jinkela_wire_8315;
    wire new_Jinkela_wire_4410;
    wire new_Jinkela_wire_2298;
    wire new_Jinkela_wire_3443;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_13265;
    wire new_Jinkela_wire_5940;
    wire new_Jinkela_wire_12891;
    wire new_Jinkela_wire_15001;
    wire new_Jinkela_wire_6524;
    wire _0101_;
    wire new_Jinkela_wire_16313;
    wire new_Jinkela_wire_12164;
    wire new_Jinkela_wire_18210;
    wire new_Jinkela_wire_7225;
    wire new_Jinkela_wire_3776;
    wire new_Jinkela_wire_17769;
    wire new_Jinkela_wire_16175;
    wire new_Jinkela_wire_18959;
    wire new_Jinkela_wire_14240;
    wire new_Jinkela_wire_18961;
    wire new_Jinkela_wire_18965;
    wire new_Jinkela_wire_5073;
    wire new_Jinkela_wire_17650;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_8823;
    wire new_Jinkela_wire_4689;
    wire new_Jinkela_wire_3748;
    wire new_Jinkela_wire_20636;
    wire new_Jinkela_wire_9490;
    wire new_Jinkela_wire_9360;
    wire new_Jinkela_wire_19462;
    wire new_Jinkela_wire_13710;
    wire new_Jinkela_wire_20873;
    wire new_Jinkela_wire_13318;
    wire _1384_;
    wire new_Jinkela_wire_13458;
    wire new_Jinkela_wire_20512;
    wire new_Jinkela_wire_6868;
    wire new_Jinkela_wire_8404;
    wire new_Jinkela_wire_20774;
    wire new_Jinkela_wire_10985;
    wire new_Jinkela_wire_19409;
    wire new_Jinkela_wire_5064;
    wire new_Jinkela_wire_21090;
    wire new_Jinkela_wire_21181;
    wire new_Jinkela_wire_18222;
    wire new_Jinkela_wire_19848;
    wire new_Jinkela_wire_12645;
    wire new_Jinkela_wire_16641;
    wire new_Jinkela_wire_16357;
    wire new_Jinkela_wire_4264;
    wire new_Jinkela_wire_9770;
    wire new_Jinkela_wire_8380;
    wire new_Jinkela_wire_18711;
    wire new_Jinkela_wire_17597;
    wire new_Jinkela_wire_4433;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_16218;
    wire new_Jinkela_wire_7235;
    wire new_Jinkela_wire_7156;
    wire new_Jinkela_wire_19938;
    wire new_Jinkela_wire_14262;
    wire _0922_;
    wire new_Jinkela_wire_15956;
    wire new_Jinkela_wire_13345;
    wire new_Jinkela_wire_18239;
    wire new_Jinkela_wire_8262;
    wire new_Jinkela_wire_17635;
    wire new_Jinkela_wire_13148;
    wire new_Jinkela_wire_19732;
    wire new_Jinkela_wire_18878;
    wire _0027_;
    wire new_Jinkela_wire_8449;
    wire new_Jinkela_wire_14516;
    wire new_Jinkela_wire_13000;
    wire new_Jinkela_wire_21229;
    wire new_Jinkela_wire_11417;
    wire new_Jinkela_wire_12752;
    wire _0910_;
    wire new_Jinkela_wire_7671;
    wire new_Jinkela_wire_7981;
    wire _0991_;
    wire new_Jinkela_wire_12133;
    wire new_Jinkela_wire_12344;
    wire new_Jinkela_wire_3617;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_20205;
    wire new_Jinkela_wire_20017;
    wire _0892_;
    wire new_Jinkela_wire_5828;
    wire new_Jinkela_wire_8602;
    wire new_Jinkela_wire_19727;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_20380;
    wire new_Jinkela_wire_16502;
    wire new_Jinkela_wire_3819;
    wire new_Jinkela_wire_10810;
    wire new_Jinkela_wire_14809;
    wire new_Jinkela_wire_14078;
    wire new_Jinkela_wire_7459;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_10576;
    wire new_Jinkela_wire_11770;
    wire new_Jinkela_wire_16212;
    wire new_Jinkela_wire_10889;
    wire new_Jinkela_wire_10858;
    wire new_Jinkela_wire_11061;
    wire new_Jinkela_wire_10444;
    wire new_Jinkela_wire_8398;
    wire new_Jinkela_wire_18027;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_9860;
    wire new_Jinkela_wire_16017;
    wire new_Jinkela_wire_21261;
    wire new_Jinkela_wire_11122;
    wire new_Jinkela_wire_13930;
    wire new_Jinkela_wire_4255;
    wire new_Jinkela_wire_12881;
    wire new_Jinkela_wire_17976;
    wire new_Jinkela_wire_10675;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_17940;
    wire new_Jinkela_wire_2156;
    wire new_Jinkela_wire_17391;
    wire new_Jinkela_wire_7171;
    wire new_Jinkela_wire_3236;
    wire new_Jinkela_wire_1822;
    wire new_Jinkela_wire_8261;
    wire new_Jinkela_wire_13216;
    wire new_Jinkela_wire_927;
    wire _0505_;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_17644;
    wire new_Jinkela_wire_6564;
    wire new_Jinkela_wire_13209;
    wire new_Jinkela_wire_14154;
    wire new_Jinkela_wire_14425;
    wire new_Jinkela_wire_5365;
    wire new_Jinkela_wire_15960;
    wire new_Jinkela_wire_7305;
    wire new_Jinkela_wire_20265;
    wire new_Jinkela_wire_14337;
    wire new_Jinkela_wire_805;
    wire _0139_;
    wire new_Jinkela_wire_11296;
    wire _1473_;
    wire _1713_;
    wire new_Jinkela_wire_10848;
    wire new_Jinkela_wire_20993;
    wire new_Jinkela_wire_3389;
    wire new_Jinkela_wire_21206;
    wire new_Jinkela_wire_19659;
    wire new_Jinkela_wire_6824;
    wire _0484_;
    wire _0157_;
    wire new_Jinkela_wire_16431;
    wire new_Jinkela_wire_16316;
    wire new_Jinkela_wire_6425;
    wire new_Jinkela_wire_17851;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_1779;
    wire new_Jinkela_wire_6254;
    wire new_Jinkela_wire_3403;
    wire new_Jinkela_wire_17418;
    wire new_Jinkela_wire_7328;
    wire new_Jinkela_wire_10664;
    wire new_Jinkela_wire_20489;
    wire new_Jinkela_wire_9317;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_14194;
    wire new_Jinkela_wire_2440;
    wire new_Jinkela_wire_4943;
    wire new_Jinkela_wire_19150;
    wire new_Jinkela_wire_13894;
    wire new_Jinkela_wire_6776;
    wire new_Jinkela_wire_13657;
    wire new_Jinkela_wire_20037;
    wire new_Jinkela_wire_11817;
    wire new_Jinkela_wire_4319;
    wire new_Jinkela_wire_2045;
    wire new_Jinkela_wire_14838;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_8798;
    wire new_Jinkela_wire_16842;
    wire new_Jinkela_wire_6095;
    wire new_Jinkela_wire_16608;
    wire new_Jinkela_wire_8484;
    wire new_Jinkela_wire_16683;
    wire new_Jinkela_wire_16378;
    wire new_Jinkela_wire_3350;
    wire new_Jinkela_wire_4771;
    wire new_Jinkela_wire_2161;
    wire new_Jinkela_wire_10594;
    wire new_Jinkela_wire_12657;
    wire new_Jinkela_wire_13518;
    wire new_Jinkela_wire_9963;
    wire new_Jinkela_wire_21323;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_7248;
    wire new_Jinkela_wire_18426;
    wire new_Jinkela_wire_16233;
    wire new_Jinkela_wire_7881;
    wire new_Jinkela_wire_7083;
    wire new_Jinkela_wire_10604;
    wire new_Jinkela_wire_11110;
    wire new_Jinkela_wire_20727;
    wire new_Jinkela_wire_18505;
    wire new_Jinkela_wire_18635;
    wire new_Jinkela_wire_14474;
    wire new_Jinkela_wire_12347;
    wire new_Jinkela_wire_16142;
    wire new_Jinkela_wire_9837;
    wire new_Jinkela_wire_20019;
    wire new_Jinkela_wire_20251;
    wire new_Jinkela_wire_19028;
    wire new_Jinkela_wire_20824;
    wire _0823_;
    wire new_Jinkela_wire_11486;
    wire new_Jinkela_wire_18530;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_1949;
    wire new_Jinkela_wire_6183;
    wire new_Jinkela_wire_6696;
    wire new_Jinkela_wire_4209;
    wire new_Jinkela_wire_20435;
    wire new_Jinkela_wire_19515;
    wire new_Jinkela_wire_7317;
    wire new_Jinkela_wire_11163;
    wire new_Jinkela_wire_17285;
    wire new_Jinkela_wire_6245;
    wire new_Jinkela_wire_5977;
    wire new_Jinkela_wire_19538;
    wire new_Jinkela_wire_19647;
    wire new_Jinkela_wire_4679;
    wire new_Jinkela_wire_16793;
    wire new_Jinkela_wire_5615;
    wire new_Jinkela_wire_4543;
    wire _1250_;
    wire new_Jinkela_wire_5033;
    wire new_Jinkela_wire_14317;
    wire new_Jinkela_wire_12356;
    wire new_Jinkela_wire_13653;
    wire new_Jinkela_wire_9210;
    wire new_Jinkela_wire_16562;
    wire _1451_;
    wire new_Jinkela_wire_14477;
    wire new_Jinkela_wire_16605;
    wire new_Jinkela_wire_4859;
    wire new_Jinkela_wire_8429;
    wire new_Jinkela_wire_13062;
    wire new_Jinkela_wire_9971;
    wire new_Jinkela_wire_4851;
    wire new_Jinkela_wire_21208;
    wire new_Jinkela_wire_17712;
    wire new_Jinkela_wire_11432;
    wire new_Jinkela_wire_8013;
    wire new_Jinkela_wire_11522;
    wire new_Jinkela_wire_11975;
    wire new_Jinkela_wire_17070;
    wire new_Jinkela_wire_5916;
    wire new_Jinkela_wire_14707;
    wire new_Jinkela_wire_5637;
    wire new_Jinkela_wire_14479;
    wire new_Jinkela_wire_2546;
    wire new_Jinkela_wire_3346;
    wire new_Jinkela_wire_16665;
    wire new_Jinkela_wire_17007;
    wire new_Jinkela_wire_2054;
    wire new_Jinkela_wire_4867;
    wire new_Jinkela_wire_9954;
    wire new_Jinkela_wire_10258;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_9002;
    wire new_Jinkela_wire_19716;
    wire new_Jinkela_wire_4353;
    wire new_Jinkela_wire_7466;
    wire new_Jinkela_wire_2370;
    wire new_Jinkela_wire_5202;
    wire new_Jinkela_wire_8783;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_21086;
    wire _0622_;
    wire new_Jinkela_wire_9337;
    wire new_Jinkela_wire_14042;
    wire new_Jinkela_wire_12592;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_19158;
    wire new_Jinkela_wire_6049;
    wire new_Jinkela_wire_17649;
    wire new_Jinkela_wire_6433;
    wire _1543_;
    wire new_Jinkela_wire_2981;
    wire new_Jinkela_wire_2387;
    wire new_Jinkela_wire_15535;
    wire new_Jinkela_wire_13802;
    wire new_Jinkela_wire_1151;
    wire _0603_;
    wire new_Jinkela_wire_4837;
    wire new_Jinkela_wire_19209;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_7211;
    wire _1110_;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_7237;
    wire new_Jinkela_wire_8582;
    wire new_Jinkela_wire_21045;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_19889;
    wire new_Jinkela_wire_9256;
    wire new_Jinkela_wire_19416;
    wire new_Jinkela_wire_20369;
    wire new_Jinkela_wire_7371;
    wire new_Jinkela_wire_14386;
    wire new_Jinkela_wire_2734;
    wire new_Jinkela_wire_6650;
    wire new_Jinkela_wire_10705;
    wire new_Jinkela_wire_19988;
    wire new_Jinkela_wire_10048;
    wire new_Jinkela_wire_2442;
    wire new_Jinkela_wire_7564;
    wire new_Jinkela_wire_16879;
    wire new_Jinkela_wire_15803;
    wire new_Jinkela_wire_7266;
    wire new_Jinkela_wire_15128;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_7751;
    wire new_Jinkela_wire_6461;
    wire new_Jinkela_wire_20203;
    wire new_Jinkela_wire_19437;
    wire new_Jinkela_wire_9302;
    wire new_Jinkela_wire_3293;
    wire new_Jinkela_wire_6976;
    wire new_Jinkela_wire_8747;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_10606;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_15952;
    wire new_Jinkela_wire_4291;
    wire new_Jinkela_wire_21204;
    wire new_Jinkela_wire_7587;
    wire new_Jinkela_wire_10949;
    wire new_Jinkela_wire_10498;
    wire new_Jinkela_wire_2115;
    wire new_Jinkela_wire_16612;
    wire new_Jinkela_wire_7445;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_3129;
    wire new_Jinkela_wire_13498;
    wire new_Jinkela_wire_13835;
    wire new_Jinkela_wire_18402;
    wire new_Jinkela_wire_14529;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_20476;
    wire new_Jinkela_wire_2746;
    wire _0076_;
    wire new_Jinkela_wire_12146;
    wire new_Jinkela_wire_19155;
    wire _1372_;
    wire new_Jinkela_wire_2483;
    wire new_Jinkela_wire_16686;
    wire new_Jinkela_wire_17123;
    wire new_Jinkela_wire_19251;
    wire _0486_;
    wire new_Jinkela_wire_7393;
    wire _0868_;
    wire new_Jinkela_wire_6899;
    wire new_Jinkela_wire_4138;
    wire new_Jinkela_wire_9025;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_10155;
    wire new_Jinkela_wire_20566;
    wire _1221_;
    wire new_Jinkela_wire_2662;
    wire new_Jinkela_wire_9973;
    wire new_Jinkela_wire_17872;
    wire new_Jinkela_wire_5116;
    wire new_Jinkela_wire_2619;
    wire new_Jinkela_wire_16029;
    wire new_Jinkela_wire_14447;
    wire new_Jinkela_wire_4704;
    wire new_Jinkela_wire_19970;
    wire new_Jinkela_wire_10573;
    wire new_Jinkela_wire_6598;
    wire new_Jinkela_wire_18536;
    wire _0273_;
    wire new_Jinkela_wire_1757;
    wire new_Jinkela_wire_10626;
    wire new_Jinkela_wire_15880;
    wire new_Jinkela_wire_16667;
    wire new_Jinkela_wire_13189;
    wire new_Jinkela_wire_3966;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_7414;
    wire new_Jinkela_wire_10480;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_4194;
    wire new_Jinkela_wire_9487;
    wire new_Jinkela_wire_7589;
    wire new_Jinkela_wire_2637;
    wire new_Jinkela_wire_7173;
    wire new_Jinkela_wire_13272;
    wire new_Jinkela_wire_17258;
    wire new_Jinkela_wire_3010;
    wire new_Jinkela_wire_3401;
    wire new_Jinkela_wire_7794;
    wire new_Jinkela_wire_1833;
    wire new_Jinkela_wire_10648;
    wire new_Jinkela_wire_13721;
    wire new_Jinkela_wire_17828;
    wire new_Jinkela_wire_16069;
    wire new_Jinkela_wire_2616;
    wire new_Jinkela_wire_3103;
    wire new_Jinkela_wire_16898;
    wire new_Jinkela_wire_10785;
    wire new_Jinkela_wire_2991;
    wire new_Jinkela_wire_18223;
    wire new_Jinkela_wire_9601;
    wire _0072_;
    wire new_Jinkela_wire_16527;
    wire new_Jinkela_wire_16005;
    wire new_Jinkela_wire_14557;
    wire new_Jinkela_wire_9567;
    wire new_Jinkela_wire_18745;
    wire new_Jinkela_wire_21331;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_11117;
    wire new_Jinkela_wire_4941;
    wire _1147_;
    wire new_Jinkela_wire_4987;
    wire new_Jinkela_wire_9272;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_9575;
    wire new_Jinkela_wire_19816;
    wire new_Jinkela_wire_9414;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_13875;
    wire new_Jinkela_wire_7329;
    wire new_Jinkela_wire_19137;
    wire new_Jinkela_wire_20889;
    wire new_Jinkela_wire_2384;
    wire new_Jinkela_wire_10243;
    wire new_Jinkela_wire_20863;
    wire new_Jinkela_wire_4948;
    wire new_Jinkela_wire_9049;
    wire new_Jinkela_wire_18454;
    wire new_Jinkela_wire_9866;
    wire new_Jinkela_wire_12263;
    wire new_Jinkela_wire_17310;
    wire new_Jinkela_wire_2088;
    wire new_Jinkela_wire_15320;
    wire new_Jinkela_wire_6412;
    wire new_Jinkela_wire_15915;
    wire _0068_;
    wire new_Jinkela_wire_19857;
    wire new_Jinkela_wire_14436;
    wire new_Jinkela_wire_15377;
    wire new_Jinkela_wire_8745;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_18831;
    wire new_Jinkela_wire_6106;
    wire new_Jinkela_wire_19293;
    wire new_Jinkela_wire_15831;
    wire _1340_;
    wire _0416_;
    wire new_Jinkela_wire_16732;
    wire new_Jinkela_wire_12905;
    wire new_Jinkela_wire_16443;
    wire new_Jinkela_wire_9930;
    wire new_Jinkela_wire_19030;
    wire new_Jinkela_wire_20074;
    wire new_Jinkela_wire_16646;
    wire new_Jinkela_wire_8064;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_8288;
    wire new_Jinkela_wire_8331;
    wire new_Jinkela_wire_21193;
    wire new_Jinkela_wire_12679;
    wire new_Jinkela_wire_8088;
    wire new_Jinkela_wire_14009;
    wire new_Jinkela_wire_10685;
    wire new_Jinkela_wire_18388;
    wire new_Jinkela_wire_18125;
    wire new_Jinkela_wire_5090;
    wire new_Jinkela_wire_10589;
    wire new_Jinkela_wire_15669;
    wire new_Jinkela_wire_14624;
    wire new_Jinkela_wire_4547;
    wire new_Jinkela_wire_17620;
    wire new_Jinkela_wire_3835;
    wire new_Jinkela_wire_11386;
    wire new_Jinkela_wire_9728;
    wire new_Jinkela_wire_9917;
    wire new_Jinkela_wire_12662;
    wire new_Jinkela_wire_7136;
    wire new_Jinkela_wire_2010;
    wire new_Jinkela_wire_20272;
    wire new_Jinkela_wire_11310;
    wire new_Jinkela_wire_3538;
    wire new_Jinkela_wire_11011;
    wire new_Jinkela_wire_2999;
    wire new_Jinkela_wire_6812;
    wire new_Jinkela_wire_20553;
    wire new_Jinkela_wire_19941;
    wire new_Jinkela_wire_13888;
    wire new_Jinkela_wire_21326;
    wire new_Jinkela_wire_19856;
    wire new_Jinkela_wire_8348;
    wire new_Jinkela_wire_15220;
    wire new_Jinkela_wire_13188;
    wire new_Jinkela_wire_13783;
    wire new_Jinkela_wire_11734;
    wire new_Jinkela_wire_3716;
    wire new_Jinkela_wire_2418;
    wire new_Jinkela_wire_16303;
    wire new_Jinkela_wire_11929;
    wire new_Jinkela_wire_4128;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_9155;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_21314;
    wire new_Jinkela_wire_7780;
    wire new_Jinkela_wire_16874;
    wire new_Jinkela_wire_8029;
    wire new_Jinkela_wire_20925;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_2778;
    wire new_Jinkela_wire_8021;
    wire new_Jinkela_wire_5052;
    wire new_Jinkela_wire_16236;
    wire new_Jinkela_wire_12748;
    wire new_Jinkela_wire_10695;
    wire new_Jinkela_wire_10928;
    wire new_Jinkela_wire_18379;
    wire _1030_;
    wire new_Jinkela_wire_15802;
    wire new_Jinkela_wire_10415;
    wire new_Jinkela_wire_14257;
    wire new_Jinkela_wire_18987;
    wire new_Jinkela_wire_7154;
    wire new_Jinkela_wire_18055;
    wire new_Jinkela_wire_11220;
    wire _0674_;
    wire new_Jinkela_wire_9281;
    wire new_Jinkela_wire_12414;
    wire new_Jinkela_wire_12744;
    wire new_Jinkela_wire_5500;
    wire new_Jinkela_wire_19805;
    wire _1824_;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_7769;
    wire new_Jinkela_wire_13337;
    wire new_Jinkela_wire_14501;
    wire _1521_;
    wire new_Jinkela_wire_10529;
    wire new_Jinkela_wire_12407;
    wire new_Jinkela_wire_15659;
    wire new_Jinkela_wire_11159;
    wire new_Jinkela_wire_12841;
    wire new_Jinkela_wire_2207;
    wire new_Jinkela_wire_8805;
    wire new_Jinkela_wire_6043;
    wire new_Jinkela_wire_18683;
    wire new_Jinkela_wire_16222;
    wire _0742_;
    wire new_Jinkela_wire_19740;
    wire new_Jinkela_wire_8145;
    wire new_Jinkela_wire_2254;
    wire new_Jinkela_wire_5415;
    wire new_Jinkela_wire_3254;
    wire new_Jinkela_wire_11414;
    wire new_Jinkela_wire_18570;
    wire new_Jinkela_wire_5797;
    wire new_Jinkela_wire_15765;
    wire new_Jinkela_wire_20948;
    wire new_Jinkela_wire_9237;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_11781;
    wire new_Jinkela_wire_11018;
    wire new_Jinkela_wire_12058;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_12105;
    wire new_Jinkela_wire_11542;
    wire new_Jinkela_wire_9132;
    wire new_Jinkela_wire_16409;
    wire new_Jinkela_wire_20165;
    wire new_Jinkela_wire_10287;
    wire new_Jinkela_wire_17265;
    wire new_Jinkela_wire_15526;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_4876;
    wire new_Jinkela_wire_4261;
    wire new_Jinkela_wire_5966;
    wire new_Jinkela_wire_15251;
    wire new_Jinkela_wire_2382;
    wire new_Jinkela_wire_6520;
    wire new_Jinkela_wire_9792;
    wire new_Jinkela_wire_15478;
    wire new_Jinkela_wire_12855;
    wire new_Jinkela_wire_3167;
    wire new_Jinkela_wire_12433;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_9139;
    wire new_Jinkela_wire_4894;
    wire new_Jinkela_wire_17577;
    wire new_Jinkela_wire_16468;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_2138;
    wire new_Jinkela_wire_4766;
    wire new_Jinkela_wire_13654;
    wire new_Jinkela_wire_4310;
    wire new_Jinkela_wire_15044;
    wire _1316_;
    wire new_Jinkela_wire_17818;
    wire new_Jinkela_wire_16719;
    wire new_Jinkela_wire_5537;
    wire new_Jinkela_wire_15689;
    wire new_Jinkela_wire_2430;
    wire new_Jinkela_wire_20715;
    wire _0395_;
    wire new_Jinkela_wire_18348;
    wire new_Jinkela_wire_19438;
    wire new_Jinkela_wire_12762;
    wire new_Jinkela_wire_18840;
    wire new_Jinkela_wire_13482;
    wire new_Jinkela_wire_20339;
    wire new_Jinkela_wire_2560;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_11234;
    wire new_Jinkela_wire_8500;
    wire _0999_;
    wire new_Jinkela_wire_14310;
    wire new_Jinkela_wire_11141;
    wire new_Jinkela_wire_19015;
    wire new_Jinkela_wire_1896;
    wire new_Jinkela_wire_9318;
    wire new_Jinkela_wire_8951;
    wire new_Jinkela_wire_9168;
    wire new_Jinkela_wire_12419;
    wire new_Jinkela_wire_2403;
    wire new_Jinkela_wire_11286;
    wire new_Jinkela_wire_17493;
    wire new_Jinkela_wire_8166;
    wire new_Jinkela_wire_8330;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_16352;
    wire new_Jinkela_wire_14454;
    wire new_Jinkela_wire_5387;
    wire new_Jinkela_wire_20892;
    wire new_Jinkela_wire_4792;
    wire new_Jinkela_wire_10712;
    wire new_Jinkela_wire_17312;
    wire new_Jinkela_wire_3971;
    wire new_Jinkela_wire_9392;
    wire new_Jinkela_wire_11824;
    wire new_Jinkela_wire_8618;
    wire new_Jinkela_wire_6131;
    wire new_Jinkela_wire_7279;
    wire new_Jinkela_wire_4060;
    wire new_Jinkela_wire_14235;
    wire new_Jinkela_wire_9511;
    wire new_Jinkela_wire_12231;
    wire new_Jinkela_wire_9113;
    wire new_Jinkela_wire_7882;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_3512;
    wire new_Jinkela_wire_18342;
    wire new_Jinkela_wire_19070;
    wire new_Jinkela_wire_7144;
    wire new_Jinkela_wire_7569;
    wire new_Jinkela_wire_14565;
    wire new_Jinkela_wire_14560;
    wire new_Jinkela_wire_7533;
    wire new_Jinkela_wire_21122;
    wire new_Jinkela_wire_10955;
    wire new_Jinkela_wire_15554;
    wire new_Jinkela_wire_9353;
    wire new_Jinkela_wire_9815;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_12646;
    wire new_Jinkela_wire_21299;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_20130;
    wire new_Jinkela_wire_5285;
    wire new_Jinkela_wire_17088;
    wire new_Jinkela_wire_20349;
    wire new_Jinkela_wire_4280;
    wire new_Jinkela_wire_16134;
    wire _0904_;
    wire new_Jinkela_wire_3630;
    wire _1185_;
    wire new_Jinkela_wire_16235;
    wire new_Jinkela_wire_21139;
    wire new_Jinkela_wire_14804;
    wire new_Jinkela_wire_5517;
    wire new_Jinkela_wire_16761;
    wire new_Jinkela_wire_4761;
    wire new_Jinkela_wire_9969;
    wire new_Jinkela_wire_5513;
    wire _0997_;
    wire new_Jinkela_wire_9499;
    wire new_Jinkela_wire_5691;
    wire new_Jinkela_wire_1266;
    wire new_Jinkela_wire_4047;
    wire new_Jinkela_wire_3366;
    wire new_Jinkela_wire_11491;
    wire new_Jinkela_wire_20042;
    wire _0042_;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_4009;
    wire _1458_;
    wire new_Jinkela_wire_6085;
    wire new_Jinkela_wire_9795;
    wire new_Jinkela_wire_19881;
    wire _0625_;
    wire new_Jinkela_wire_11592;
    wire new_Jinkela_wire_4372;
    wire new_Jinkela_wire_14500;
    wire new_Jinkela_wire_6987;
    wire new_Jinkela_wire_5890;
    wire _0735_;
    wire new_Jinkela_wire_11241;
    wire new_Jinkela_wire_7340;
    wire new_Jinkela_wire_2342;
    wire new_Jinkela_wire_11404;
    wire new_Jinkela_wire_18609;
    wire new_Jinkela_wire_16328;
    wire new_Jinkela_wire_13712;
    wire new_Jinkela_wire_16305;
    wire new_Jinkela_wire_5066;
    wire _0279_;
    wire new_Jinkela_wire_5951;
    wire new_Jinkela_wire_6489;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_17802;
    wire new_Jinkela_wire_9653;
    wire new_Jinkela_wire_20100;
    wire new_Jinkela_wire_17757;
    wire new_Jinkela_wire_4311;
    wire new_Jinkela_wire_2935;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_15491;
    wire new_Jinkela_wire_16018;
    wire new_Jinkela_wire_13539;
    wire _1249_;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_14504;
    wire new_Jinkela_wire_19173;
    wire new_Jinkela_wire_18506;
    wire new_Jinkela_wire_16820;
    wire new_Jinkela_wire_8041;
    wire new_Jinkela_wire_15620;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_1860;
    wire _1349_;
    wire new_Jinkela_wire_13508;
    wire new_Jinkela_wire_4751;
    wire new_Jinkela_wire_12779;
    wire new_Jinkela_wire_6062;
    wire new_Jinkela_wire_11895;
    wire new_Jinkela_wire_12959;
    wire new_Jinkela_wire_1972;
    wire new_Jinkela_wire_12273;
    wire new_Jinkela_wire_18534;
    wire new_Jinkela_wire_13942;
    wire new_Jinkela_wire_15426;
    wire new_Jinkela_wire_4960;
    wire new_Jinkela_wire_11344;
    wire new_Jinkela_wire_3946;
    wire new_Jinkela_wire_933;
    wire _1310_;
    wire new_Jinkela_wire_17623;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_4021;
    wire new_Jinkela_wire_5529;
    wire new_Jinkela_wire_17925;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_16411;
    wire new_Jinkela_wire_14908;
    wire new_Jinkela_wire_16827;
    wire new_Jinkela_wire_15094;
    wire new_Jinkela_wire_14387;
    wire new_Jinkela_wire_7115;
    wire new_Jinkela_wire_4346;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_4906;
    wire new_Jinkela_wire_13009;
    wire new_Jinkela_wire_2750;
    wire new_Jinkela_wire_13640;
    wire new_Jinkela_wire_13454;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_20314;
    wire new_Jinkela_wire_11862;
    wire _0333_;
    wire _1616_;
    wire new_Jinkela_wire_19630;
    wire new_Jinkela_wire_20204;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_21115;
    wire new_Jinkela_wire_19398;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_20651;
    wire new_Jinkela_wire_14123;
    wire new_Jinkela_wire_8391;
    wire new_Jinkela_wire_14048;
    wire new_Jinkela_wire_20418;
    wire new_Jinkela_wire_9811;
    wire new_Jinkela_wire_11551;
    wire _0685_;
    wire new_Jinkela_wire_2306;
    wire _1556_;
    wire new_Jinkela_wire_16334;
    wire new_Jinkela_wire_14186;
    wire new_Jinkela_wire_10694;
    wire new_Jinkela_wire_21114;
    wire new_Jinkela_wire_20955;
    wire new_Jinkela_wire_15647;
    wire _1127_;
    wire new_Jinkela_wire_3058;
    wire new_Jinkela_wire_13895;
    wire new_Jinkela_wire_11157;
    wire new_Jinkela_wire_21028;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_8443;
    wire _0201_;
    wire new_Jinkela_wire_12119;
    wire new_Jinkela_wire_8438;
    wire new_Jinkela_wire_15791;
    wire _0261_;
    wire new_Jinkela_wire_7788;
    wire new_Jinkela_wire_10458;
    wire new_Jinkela_wire_12796;
    wire new_Jinkela_wire_15475;
    wire new_Jinkela_wire_6972;
    wire new_Jinkela_wire_12907;
    wire new_Jinkela_wire_6190;
    wire new_Jinkela_wire_14996;
    wire new_Jinkela_wire_3056;
    wire new_Jinkela_wire_15524;
    wire new_Jinkela_wire_13260;
    wire new_Jinkela_wire_3178;
    wire new_Jinkela_wire_12026;
    wire new_Jinkela_wire_8415;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_7446;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_9364;
    wire new_Jinkela_wire_14348;
    wire new_Jinkela_wire_18233;
    wire new_Jinkela_wire_12589;
    wire new_Jinkela_wire_10001;
    wire new_Jinkela_wire_568;
    wire _0372_;
    wire new_Jinkela_wire_9404;
    wire new_Jinkela_wire_14150;
    wire new_Jinkela_wire_15996;
    wire new_Jinkela_wire_9590;
    wire new_Jinkela_wire_15888;
    wire new_Jinkela_wire_19368;
    wire _1355_;
    wire new_Jinkela_wire_14628;
    wire new_Jinkela_wire_12509;
    wire _1188_;
    wire new_Jinkela_wire_5127;
    wire new_Jinkela_wire_5991;
    wire new_Jinkela_wire_16337;
    wire new_Jinkela_wire_9259;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_17559;
    wire new_Jinkela_wire_11613;
    wire new_Jinkela_wire_7865;
    wire new_Jinkela_wire_10144;
    wire new_Jinkela_wire_1729;
    wire new_Jinkela_wire_7517;
    wire _0207_;
    wire new_Jinkela_wire_197;
    wire _0720_;
    wire new_Jinkela_wire_13554;
    wire new_Jinkela_wire_17847;
    wire new_Jinkela_wire_20110;
    wire _1600_;
    wire new_Jinkela_wire_5475;
    wire new_Jinkela_wire_16995;
    wire new_Jinkela_wire_2901;
    wire new_Jinkela_wire_9876;
    wire new_Jinkela_wire_10496;
    wire new_Jinkela_wire_10362;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_11866;
    wire new_Jinkela_wire_17427;
    wire _1369_;
    wire new_Jinkela_wire_15071;
    wire new_Jinkela_wire_8660;
    wire new_Jinkela_wire_10136;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_3271;
    wire new_Jinkela_wire_17375;
    wire new_Jinkela_wire_5689;
    wire new_Jinkela_wire_11716;
    wire _0818_;
    wire new_Jinkela_wire_12879;
    wire new_Jinkela_wire_13645;
    wire new_Jinkela_wire_8187;
    wire new_Jinkela_wire_9505;
    wire new_Jinkela_wire_3502;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_19024;
    wire new_Jinkela_wire_5939;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_19682;
    wire new_Jinkela_wire_20631;
    wire new_Jinkela_wire_6323;
    wire new_Jinkela_wire_20627;
    wire _1025_;
    wire new_Jinkela_wire_14494;
    wire new_Jinkela_wire_8729;
    wire new_Jinkela_wire_17816;
    wire new_Jinkela_wire_10613;
    wire new_Jinkela_wire_11102;
    wire new_Jinkela_wire_17395;
    wire new_Jinkela_wire_16206;
    wire new_Jinkela_wire_18124;
    wire new_Jinkela_wire_17072;
    wire new_Jinkela_wire_9679;
    wire new_Jinkela_wire_2990;
    wire new_Jinkela_wire_4888;
    wire new_Jinkela_wire_7479;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_7891;
    wire new_Jinkela_wire_5808;
    wire new_Jinkela_wire_8615;
    wire new_Jinkela_wire_20591;
    wire new_Jinkela_wire_19624;
    wire new_Jinkela_wire_19534;
    wire new_Jinkela_wire_6677;
    wire new_Jinkela_wire_14351;
    wire new_Jinkela_wire_16320;
    wire new_Jinkela_wire_4861;
    wire new_Jinkela_wire_5607;
    wire new_Jinkela_wire_10007;
    wire new_Jinkela_wire_18408;
    wire new_Jinkela_wire_9065;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_5260;
    wire new_Jinkela_wire_19507;
    wire new_Jinkela_wire_1697;
    wire new_Jinkela_wire_19444;
    wire new_Jinkela_wire_3755;
    wire new_Jinkela_wire_3142;
    wire new_Jinkela_wire_5695;
    wire new_Jinkela_wire_17205;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_2852;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_4597;
    wire _0860_;
    wire new_Jinkela_wire_6275;
    wire new_Jinkela_wire_20355;
    wire new_Jinkela_wire_12293;
    wire new_Jinkela_wire_4722;
    wire new_Jinkela_wire_14944;
    wire new_Jinkela_wire_6775;
    wire new_Jinkela_wire_13701;
    wire new_Jinkela_wire_13151;
    wire new_Jinkela_wire_9131;
    wire new_Jinkela_wire_9453;
    wire _1232_;
    wire new_Jinkela_wire_5253;
    wire new_Jinkela_wire_12167;
    wire new_Jinkela_wire_10181;
    wire new_Jinkela_wire_5524;
    wire new_Jinkela_wire_2880;
    wire new_Jinkela_wire_18330;
    wire new_Jinkela_wire_5458;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_9047;
    wire new_Jinkela_wire_12470;
    wire new_Jinkela_wire_7219;
    wire new_Jinkela_wire_5271;
    wire new_Jinkela_wire_15375;
    wire new_Jinkela_wire_8198;
    wire _0817_;
    wire new_Jinkela_wire_14733;
    wire new_Jinkela_wire_7336;
    wire new_Jinkela_wire_19344;
    wire new_Jinkela_wire_15585;
    wire _0149_;
    wire new_Jinkela_wire_17158;
    wire new_Jinkela_wire_21304;
    wire _1743_;
    wire new_Jinkela_wire_14631;
    wire new_Jinkela_wire_7809;
    wire _0563_;
    wire new_Jinkela_wire_11502;
    wire new_Jinkela_wire_8585;
    wire new_Jinkela_wire_4632;
    wire new_Jinkela_wire_18334;
    wire new_Jinkela_wire_11399;
    wire new_Jinkela_wire_16279;
    wire new_Jinkela_wire_2927;
    wire new_Jinkela_wire_11747;
    wire new_Jinkela_wire_9137;
    wire new_Jinkela_wire_4072;
    wire new_Jinkela_wire_13511;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_16790;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_14509;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_4204;
    wire new_Jinkela_wire_6620;
    wire new_Jinkela_wire_9308;
    wire new_Jinkela_wire_9773;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_11801;
    wire new_Jinkela_wire_16471;
    wire new_Jinkela_wire_16632;
    wire new_Jinkela_wire_3909;
    wire new_Jinkela_wire_7932;
    wire new_Jinkela_wire_15140;
    wire new_Jinkela_wire_2811;
    wire new_Jinkela_wire_16345;
    wire new_Jinkela_wire_20964;
    wire new_Jinkela_wire_18276;
    wire new_Jinkela_wire_4071;
    wire new_Jinkela_wire_10657;
    wire new_Jinkela_wire_11627;
    wire new_Jinkela_wire_11632;
    wire new_Jinkela_wire_3629;
    wire new_Jinkela_wire_11071;
    wire new_Jinkela_wire_6487;
    wire new_Jinkela_wire_2716;
    wire new_Jinkela_wire_6662;
    wire new_Jinkela_wire_10520;
    wire new_Jinkela_wire_14300;
    wire new_Jinkela_wire_16800;
    wire new_Jinkela_wire_7132;
    wire new_Jinkela_wire_20966;
    wire _1079_;
    wire new_Jinkela_wire_6893;
    wire new_Jinkela_wire_2057;
    wire new_Jinkela_wire_3823;
    wire new_Jinkela_wire_21318;
    wire new_Jinkela_wire_3916;
    wire new_Jinkela_wire_20061;
    wire new_Jinkela_wire_2669;
    wire new_Jinkela_wire_11150;
    wire new_Jinkela_wire_10778;
    wire new_Jinkela_wire_19505;
    wire new_Jinkela_wire_16722;
    wire new_Jinkela_wire_14728;
    wire new_Jinkela_wire_19977;
    wire _0581_;
    wire new_Jinkela_wire_10382;
    wire new_Jinkela_wire_18327;
    wire new_Jinkela_wire_14476;
    wire new_Jinkela_wire_16170;
    wire _0602_;
    wire new_Jinkela_wire_14173;
    wire new_Jinkela_wire_20117;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_18829;
    wire _0326_;
    wire new_Jinkela_wire_19310;
    wire new_Jinkela_wire_16009;
    wire new_Jinkela_wire_12650;
    wire new_Jinkela_wire_10860;
    wire new_Jinkela_wire_12389;
    wire _0469_;
    wire new_Jinkela_wire_17336;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_2944;
    wire new_Jinkela_wire_2869;
    wire new_Jinkela_wire_15651;
    wire new_Jinkela_wire_7221;
    wire new_Jinkela_wire_15206;
    wire new_Jinkela_wire_18567;
    wire new_Jinkela_wire_3888;
    wire new_Jinkela_wire_8676;
    wire new_Jinkela_wire_10224;
    wire new_Jinkela_wire_15212;
    wire new_Jinkela_wire_11177;
    wire new_Jinkela_wire_16187;
    wire new_Jinkela_wire_14132;
    wire new_Jinkela_wire_20816;
    wire new_Jinkela_wire_15595;
    wire new_Jinkela_wire_8875;
    wire new_Jinkela_wire_8400;
    wire new_Jinkela_wire_13762;
    wire new_Jinkela_wire_11164;
    wire new_Jinkela_wire_9886;
    wire new_Jinkela_wire_9933;
    wire new_Jinkela_wire_9560;
    wire new_Jinkela_wire_12486;
    wire new_Jinkela_wire_2970;
    wire new_Jinkela_wire_10418;
    wire new_Jinkela_wire_4701;
    wire new_Jinkela_wire_2622;
    wire new_Jinkela_wire_13578;
    wire new_Jinkela_wire_14613;
    wire new_Jinkela_wire_13910;
    wire new_Jinkela_wire_8901;
    wire new_Jinkela_wire_13690;
    wire new_Jinkela_wire_11743;
    wire _1540_;
    wire new_Jinkela_wire_14885;
    wire new_Jinkela_wire_20557;
    wire new_Jinkela_wire_595;
    wire _1823_;
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_17534;
    wire new_Jinkela_wire_4040;
    wire new_Jinkela_wire_6218;
    wire new_Jinkela_wire_11301;
    wire new_Jinkela_wire_13039;
    wire new_Jinkela_wire_19846;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_4783;
    wire _1726_;
    wire new_Jinkela_wire_4660;
    wire new_Jinkela_wire_14782;
    wire new_Jinkela_wire_12292;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_7202;
    wire new_Jinkela_wire_3893;
    wire new_Jinkela_wire_16637;
    wire new_Jinkela_wire_18556;
    wire new_Jinkela_wire_19956;
    wire _1667_;
    wire new_Jinkela_wire_17073;
    wire new_Jinkela_wire_20689;
    wire new_Jinkela_wire_8695;
    wire new_Jinkela_wire_19082;
    wire new_Jinkela_wire_7709;
    wire new_Jinkela_wire_14111;
    wire new_Jinkela_wire_15851;
    wire new_Jinkela_wire_18306;
    wire new_Jinkela_wire_3451;
    wire new_Jinkela_wire_21256;
    wire new_Jinkela_wire_11877;
    wire new_Jinkela_wire_14079;
    wire new_Jinkela_wire_17505;
    wire new_Jinkela_wire_6100;
    wire new_Jinkela_wire_14886;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_12548;
    wire _1142_;
    wire new_Jinkela_wire_5872;
    wire new_Jinkela_wire_1915;
    wire new_Jinkela_wire_17422;
    wire new_Jinkela_wire_19415;
    wire new_Jinkela_wire_3333;
    wire _0544_;
    wire new_Jinkela_wire_2835;
    wire new_Jinkela_wire_4710;
    wire new_Jinkela_wire_17470;
    wire new_Jinkela_wire_11565;
    wire new_Jinkela_wire_1881;
    wire new_Jinkela_wire_5980;
    wire new_Jinkela_wire_6139;
    wire new_Jinkela_wire_3789;
    wire new_Jinkela_wire_2424;
    wire new_Jinkela_wire_7955;
    wire _0411_;
    wire new_Jinkela_wire_12978;
    wire new_Jinkela_wire_2881;
    wire new_Jinkela_wire_12912;
    wire new_Jinkela_wire_2781;
    wire new_Jinkela_wire_2310;
    wire new_Jinkela_wire_11489;
    wire new_Jinkela_wire_6681;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_10098;
    wire new_Jinkela_wire_14253;
    wire new_Jinkela_wire_13357;
    wire new_Jinkela_wire_12928;
    wire new_Jinkela_wire_20945;
    wire new_Jinkela_wire_20377;
    wire new_Jinkela_wire_18395;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_9251;
    wire new_Jinkela_wire_3244;
    wire new_Jinkela_wire_20412;
    wire _0445_;
    wire new_Jinkela_wire_5956;
    wire new_Jinkela_wire_2704;
    wire new_Jinkela_wire_16817;
    wire new_Jinkela_wire_15529;
    wire new_Jinkela_wire_5593;
    wire new_Jinkela_wire_16729;
    wire new_Jinkela_wire_17795;
    wire new_Jinkela_wire_12731;
    wire new_Jinkela_wire_9875;
    wire new_Jinkela_wire_2643;
    wire new_Jinkela_wire_4564;
    wire new_Jinkela_wire_3029;
    wire _0419_;
    wire new_Jinkela_wire_5055;
    wire _0998_;
    wire new_Jinkela_wire_1130;
    wire _1799_;
    wire new_Jinkela_wire_9545;
    wire new_Jinkela_wire_15266;
    wire new_Jinkela_wire_6403;
    wire new_Jinkela_wire_7461;
    wire new_Jinkela_wire_4122;
    wire new_Jinkela_wire_8395;
    wire new_Jinkela_wire_11498;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_11373;
    wire new_Jinkela_wire_18075;
    wire new_Jinkela_wire_21068;
    wire new_Jinkela_wire_14209;
    wire new_Jinkela_wire_15962;
    wire new_Jinkela_wire_4197;
    wire new_Jinkela_wire_14607;
    wire new_Jinkela_wire_3124;
    wire new_Jinkela_wire_4915;
    wire _1487_;
    wire new_Jinkela_wire_11764;
    wire new_Jinkela_wire_10082;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_16961;
    wire new_Jinkela_wire_16684;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_5843;
    wire new_Jinkela_wire_16835;
    wire new_Jinkela_wire_10256;
    wire new_Jinkela_wire_2943;
    wire new_Jinkela_wire_14919;
    wire new_Jinkela_wire_6311;
    wire _0947_;
    wire new_Jinkela_wire_18244;
    wire new_Jinkela_wire_5182;
    wire new_Jinkela_wire_19931;
    wire new_Jinkela_wire_10209;
    wire new_Jinkela_wire_18657;
    wire new_Jinkela_wire_5477;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_10814;
    wire new_Jinkela_wire_7755;
    wire new_Jinkela_wire_11276;
    wire new_Jinkela_wire_4234;
    wire new_Jinkela_wire_15989;
    wire _1402_;
    wire new_Jinkela_wire_4037;
    wire new_Jinkela_wire_6399;
    wire new_Jinkela_wire_17634;
    wire new_Jinkela_wire_16049;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_6198;
    wire new_Jinkela_wire_5172;
    wire new_Jinkela_wire_18632;
    wire new_Jinkela_wire_13173;
    wire new_Jinkela_wire_8242;
    wire new_Jinkela_wire_14354;
    wire new_Jinkela_wire_12206;
    wire new_Jinkela_wire_11400;
    wire new_Jinkela_wire_8935;
    wire new_Jinkela_wire_10008;
    wire _1548_;
    wire new_Jinkela_wire_17419;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_11756;
    wire new_Jinkela_wire_20883;
    wire new_Jinkela_wire_2509;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_9038;
    wire new_Jinkela_wire_19475;
    wire new_Jinkela_wire_1900;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_18707;
    wire new_Jinkela_wire_12472;
    wire new_Jinkela_wire_8312;
    wire _0743_;
    wire new_Jinkela_wire_16261;
    wire new_Jinkela_wire_19595;
    wire new_Jinkela_wire_4277;
    wire new_Jinkela_wire_5679;
    wire new_Jinkela_wire_20159;
    wire new_Jinkela_wire_17294;
    wire new_Jinkela_wire_11355;
    wire new_Jinkela_wire_13909;
    wire new_Jinkela_wire_19133;
    wire new_Jinkela_wire_4690;
    wire new_Jinkela_wire_7912;
    wire new_Jinkela_wire_10487;
    wire new_Jinkela_wire_2397;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_15024;
    wire new_Jinkela_wire_20307;
    wire new_Jinkela_wire_4775;
    wire new_Jinkela_wire_19539;
    wire new_Jinkela_wire_8173;
    wire new_Jinkela_wire_6805;
    wire new_Jinkela_wire_15278;
    wire new_Jinkela_wire_8335;
    wire new_Jinkela_wire_56;
    wire _0733_;
    wire new_Jinkela_wire_15928;
    wire new_Jinkela_wire_8304;
    wire new_Jinkela_wire_11803;
    wire new_Jinkela_wire_7804;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_16351;
    wire new_Jinkela_wire_13118;
    wire new_Jinkela_wire_10275;
    wire _0035_;
    wire new_Jinkela_wire_19241;
    wire new_Jinkela_wire_2052;
    wire new_Jinkela_wire_8281;
    wire new_Jinkela_wire_5639;
    wire _1229_;
    wire new_Jinkela_wire_8401;
    wire new_Jinkela_wire_1408;
    wire new_Jinkela_wire_18898;
    wire new_Jinkela_wire_18463;
    wire new_Jinkela_wire_18770;
    wire _0706_;
    wire new_Jinkela_wire_10440;
    wire _1205_;
    wire new_Jinkela_wire_14873;
    wire new_Jinkela_wire_603;
    wire _1360_;
    wire new_Jinkela_wire_10623;
    wire new_Jinkela_wire_19554;
    wire new_net_3926;
    wire new_Jinkela_wire_20905;
    wire new_Jinkela_wire_6769;
    wire new_Jinkela_wire_17862;
    wire _0253_;
    wire _1750_;
    wire new_Jinkela_wire_9619;
    wire new_Jinkela_wire_8679;
    wire new_Jinkela_wire_18401;
    wire new_Jinkela_wire_4133;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_343;
    wire _0095_;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_8203;
    wire new_Jinkela_wire_9015;
    wire new_Jinkela_wire_9007;
    wire new_Jinkela_wire_10206;
    wire new_Jinkela_wire_9267;
    wire new_Jinkela_wire_18779;
    wire new_Jinkela_wire_6027;
    wire new_Jinkela_wire_16693;
    wire new_Jinkela_wire_3664;
    wire new_Jinkela_wire_3524;
    wire _1736_;
    wire _1641_;
    wire new_Jinkela_wire_4753;
    wire new_Jinkela_wire_4976;
    wire _1728_;
    wire new_Jinkela_wire_6710;
    wire new_Jinkela_wire_5834;
    wire new_Jinkela_wire_9870;
    wire new_Jinkela_wire_2920;
    wire new_Jinkela_wire_4215;
    wire new_Jinkela_wire_11092;
    wire new_Jinkela_wire_6032;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_17692;
    wire new_Jinkela_wire_20877;
    wire new_Jinkela_wire_13257;
    wire new_Jinkela_wire_4706;
    wire new_Jinkela_wire_18397;
    wire new_Jinkela_wire_9807;
    wire new_Jinkela_wire_12845;
    wire new_Jinkela_wire_6828;
    wire new_Jinkela_wire_15728;
    wire new_Jinkela_wire_5478;
    wire new_Jinkela_wire_2573;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_4831;
    wire new_Jinkela_wire_15666;
    wire new_Jinkela_wire_13866;
    wire new_Jinkela_wire_4379;
    wire _0081_;
    wire new_Jinkela_wire_20169;
    wire new_Jinkela_wire_9853;
    wire new_Jinkela_wire_2263;
    wire new_Jinkela_wire_3065;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_16482;
    wire new_Jinkela_wire_12244;
    wire new_Jinkela_wire_10522;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_14061;
    wire new_Jinkela_wire_10298;
    wire new_Jinkela_wire_7497;
    wire new_Jinkela_wire_18202;
    wire new_Jinkela_wire_20500;
    wire new_Jinkela_wire_16191;
    wire new_Jinkela_wire_20501;
    wire _1765_;
    wire new_Jinkela_wire_12504;
    wire new_Jinkela_wire_15621;
    wire new_Jinkela_wire_7205;
    wire new_Jinkela_wire_11802;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_19825;
    wire new_Jinkela_wire_17382;
    wire new_Jinkela_wire_17588;
    wire new_Jinkela_wire_19181;
    wire new_Jinkela_wire_16056;
    wire new_Jinkela_wire_10107;
    wire new_Jinkela_wire_4601;
    wire new_Jinkela_wire_2498;
    wire new_Jinkela_wire_12708;
    wire new_Jinkela_wire_17821;
    wire new_Jinkela_wire_15873;
    wire new_Jinkela_wire_3218;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_6541;
    wire _1806_;
    wire new_Jinkela_wire_18697;
    wire new_Jinkela_wire_18022;
    wire new_Jinkela_wire_3951;
    wire new_Jinkela_wire_20326;
    wire new_Jinkela_wire_10403;
    wire _0801_;
    wire new_Jinkela_wire_20652;
    wire new_Jinkela_wire_13185;
    wire new_Jinkela_wire_7298;
    wire new_Jinkela_wire_3710;
    wire new_Jinkela_wire_17790;
    wire new_Jinkela_wire_9123;
    wire new_Jinkela_wire_4470;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_17684;
    wire new_Jinkela_wire_5367;
    wire new_Jinkela_wire_18789;
    wire new_Jinkela_wire_7259;
    wire new_Jinkela_wire_2060;
    wire new_Jinkela_wire_14159;
    wire new_Jinkela_wire_8125;
    wire new_Jinkela_wire_5756;
    wire new_Jinkela_wire_12716;
    wire new_Jinkela_wire_16264;
    wire new_Jinkela_wire_2413;
    wire new_Jinkela_wire_7153;
    wire new_Jinkela_wire_5222;
    wire _0986_;
    wire new_Jinkela_wire_13982;
    wire new_Jinkela_wire_4275;
    wire new_Jinkela_wire_1870;
    wire new_Jinkela_wire_20869;
    wire new_Jinkela_wire_11913;
    wire new_Jinkela_wire_12038;
    wire new_Jinkela_wire_6156;
    wire new_Jinkela_wire_7820;
    wire new_Jinkela_wire_8656;
    wire new_Jinkela_wire_8870;
    wire new_Jinkela_wire_2736;
    wire new_Jinkela_wire_19244;
    wire new_Jinkela_wire_15553;
    wire new_Jinkela_wire_3112;
    wire new_Jinkela_wire_13808;
    wire new_Jinkela_wire_16301;
    wire new_Jinkela_wire_16592;
    wire new_Jinkela_wire_18362;
    wire new_Jinkela_wire_8821;
    wire new_Jinkela_wire_9498;
    wire new_Jinkela_wire_2857;
    wire new_Jinkela_wire_6185;
    wire new_Jinkela_wire_20805;
    wire new_Jinkela_wire_8006;
    wire new_Jinkela_wire_21257;
    wire new_Jinkela_wire_5423;
    wire new_Jinkela_wire_16456;
    wire new_Jinkela_wire_5101;
    wire new_Jinkela_wire_8038;
    wire new_Jinkela_wire_3345;
    wire _1021_;
    wire new_Jinkela_wire_7348;
    wire _1571_;
    wire new_Jinkela_wire_21250;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_4958;
    wire new_Jinkela_wire_15056;
    wire new_Jinkela_wire_11005;
    wire new_Jinkela_wire_16015;
    wire new_Jinkela_wire_15296;
    wire new_Jinkela_wire_20768;
    wire _0034_;
    wire new_Jinkela_wire_6123;
    wire new_Jinkela_wire_12059;
    wire new_Jinkela_wire_10064;
    wire new_Jinkela_wire_3357;
    wire new_Jinkela_wire_1626;
    wire new_Jinkela_wire_17910;
    wire new_Jinkela_wire_4670;
    wire new_Jinkela_wire_9925;
    wire new_Jinkela_wire_7410;
    wire new_Jinkela_wire_10756;
    wire new_Jinkela_wire_20155;
    wire new_Jinkela_wire_3985;
    wire new_Jinkela_wire_7341;
    wire new_Jinkela_wire_11984;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_20390;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_16371;
    wire new_Jinkela_wire_8346;
    wire new_Jinkela_wire_7784;
    wire new_Jinkela_wire_10071;
    wire new_Jinkela_wire_21037;
    wire new_Jinkela_wire_2605;
    wire new_Jinkela_wire_11176;
    wire new_Jinkela_wire_10388;
    wire new_Jinkela_wire_11883;
    wire new_Jinkela_wire_8977;
    wire _0832_;
    wire new_Jinkela_wire_14874;
    wire new_Jinkela_wire_9542;
    wire new_Jinkela_wire_15486;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_19118;
    wire _0775_;
    wire new_Jinkela_wire_7986;
    wire new_Jinkela_wire_5723;
    wire new_Jinkela_wire_15061;
    wire new_Jinkela_wire_1239;
    wire _0650_;
    wire new_Jinkela_wire_10900;
    wire new_Jinkela_wire_20674;
    wire _0247_;
    wire new_Jinkela_wire_8051;
    wire new_Jinkela_wire_10234;
    wire new_Jinkela_wire_4910;
    wire new_Jinkela_wire_17953;
    wire new_Jinkela_wire_7946;
    wire new_Jinkela_wire_8826;
    wire new_Jinkela_wire_12053;
    wire new_Jinkela_wire_20745;
    wire new_Jinkela_wire_8152;
    wire _0759_;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_3673;
    wire new_Jinkela_wire_12799;
    wire new_Jinkela_wire_5292;
    wire new_Jinkela_wire_17535;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_3491;
    wire new_Jinkela_wire_5409;
    wire _0377_;
    wire new_Jinkela_wire_7748;
    wire new_Jinkela_wire_11450;
    wire new_Jinkela_wire_6054;
    wire _0187_;
    wire new_Jinkela_wire_3687;
    wire new_Jinkela_wire_17350;
    wire new_Jinkela_wire_20522;
    wire new_Jinkela_wire_17542;
    wire new_Jinkela_wire_9991;
    wire new_Jinkela_wire_20250;
    wire new_Jinkela_wire_20897;
    wire new_Jinkela_wire_2354;
    wire new_Jinkela_wire_16569;
    wire new_Jinkela_wire_9373;
    wire new_Jinkela_wire_19178;
    wire new_Jinkela_wire_9536;
    wire new_Jinkela_wire_11539;
    wire new_Jinkela_wire_13132;
    wire _0448_;
    wire new_Jinkela_wire_5270;
    wire _1652_;
    wire new_Jinkela_wire_15798;
    wire new_Jinkela_wire_14139;
    wire new_Jinkela_wire_17721;
    wire new_Jinkela_wire_5669;
    wire new_Jinkela_wire_21022;
    wire new_Jinkela_wire_8694;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_19220;
    wire new_Jinkela_wire_11440;
    wire _1138_;
    wire new_Jinkela_wire_8932;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_18130;
    wire new_Jinkela_wire_16128;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_8499;
    wire new_Jinkela_wire_3361;
    wire new_Jinkela_wire_11582;
    wire new_Jinkela_wire_12827;
    wire new_Jinkela_wire_14258;
    wire new_Jinkela_wire_17592;
    wire new_Jinkela_wire_14021;
    wire new_Jinkela_wire_5402;
    wire new_Jinkela_wire_12683;
    wire new_Jinkela_wire_13532;
    wire new_Jinkela_wire_2825;
    wire new_Jinkela_wire_5621;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_3550;
    wire new_Jinkela_wire_8661;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_15980;
    wire new_Jinkela_wire_3939;
    wire new_Jinkela_wire_2718;
    wire new_Jinkela_wire_17175;
    wire new_Jinkela_wire_17986;
    wire new_Jinkela_wire_4810;
    wire new_Jinkela_wire_8861;
    wire new_Jinkela_wire_21152;
    wire new_Jinkela_wire_10975;
    wire new_Jinkela_wire_17144;
    wire new_Jinkela_wire_2848;
    wire new_Jinkela_wire_4478;
    wire _0745_;
    wire new_Jinkela_wire_4982;
    wire new_Jinkela_wire_6820;
    wire new_Jinkela_wire_1990;
    wire new_Jinkela_wire_10512;
    wire new_Jinkela_wire_12859;
    wire new_Jinkela_wire_1656;
    wire new_Jinkela_wire_12398;
    wire new_Jinkela_wire_15342;
    wire new_Jinkela_wire_9901;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_12887;
    wire new_Jinkela_wire_3590;
    wire new_Jinkela_wire_8587;
    wire new_Jinkela_wire_4200;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_12804;
    wire new_Jinkela_wire_5914;
    wire new_Jinkela_wire_2337;
    wire new_Jinkela_wire_11510;
    wire new_Jinkela_wire_15213;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_9945;
    wire new_Jinkela_wire_12575;
    wire new_Jinkela_wire_14074;
    wire new_Jinkela_wire_13175;
    wire new_Jinkela_wire_18531;
    wire new_Jinkela_wire_4288;
    wire new_Jinkela_wire_6839;
    wire new_Jinkela_wire_3737;
    wire new_Jinkela_wire_5806;
    wire new_Jinkela_wire_6400;
    wire _0327_;
    wire new_Jinkela_wire_8270;
    wire new_Jinkela_wire_16786;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_17569;
    wire new_Jinkela_wire_12740;
    wire new_Jinkela_wire_6848;
    wire new_Jinkela_wire_3960;
    wire _0913_;
    wire new_Jinkela_wire_14839;
    wire new_Jinkela_wire_2211;
    wire _1701_;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_6536;
    wire new_Jinkela_wire_9790;
    wire _1075_;
    wire new_Jinkela_wire_13456;
    wire new_Jinkela_wire_12359;
    wire new_Jinkela_wire_4794;
    wire new_Jinkela_wire_14443;
    wire new_Jinkela_wire_21008;
    wire new_Jinkela_wire_4854;
    wire new_Jinkela_wire_5820;
    wire new_Jinkela_wire_19288;
    wire new_Jinkela_wire_9016;
    wire new_Jinkela_wire_4297;
    wire new_Jinkela_wire_10469;
    wire new_Jinkela_wire_4994;
    wire new_Jinkela_wire_18110;
    wire new_Jinkela_wire_12745;
    wire new_Jinkela_wire_14701;
    wire new_Jinkela_wire_4839;
    wire new_Jinkela_wire_17909;
    wire new_Jinkela_wire_3954;
    wire new_Jinkela_wire_15675;
    wire new_Jinkela_wire_16373;
    wire new_Jinkela_wire_6230;
    wire new_Jinkela_wire_14471;
    wire new_Jinkela_wire_12464;
    wire new_Jinkela_wire_3594;
    wire new_Jinkela_wire_7859;
    wire _1576_;
    wire _0107_;
    wire _1595_;
    wire new_Jinkela_wire_3086;
    wire new_Jinkela_wire_17230;
    wire new_Jinkela_wire_20257;
    wire _0534_;
    wire new_Jinkela_wire_14666;
    wire new_Jinkela_wire_20826;
    wire new_Jinkela_wire_5128;
    wire new_Jinkela_wire_10431;
    wire new_Jinkela_wire_18036;
    wire _1428_;
    wire new_Jinkela_wire_6314;
    wire new_Jinkela_wire_17390;
    wire new_Jinkela_wire_19018;
    wire new_Jinkela_wire_12095;
    wire new_Jinkela_wire_17835;
    wire new_Jinkela_wire_9129;
    wire new_Jinkela_wire_9620;
    wire new_Jinkela_wire_11436;
    wire new_Jinkela_wire_19620;
    wire new_Jinkela_wire_9819;
    wire new_Jinkela_wire_2608;
    wire new_Jinkela_wire_5320;
    wire new_Jinkela_wire_6957;
    wire new_Jinkela_wire_17091;
    wire new_Jinkela_wire_14780;
    wire new_Jinkela_wire_4368;
    wire new_Jinkela_wire_10125;
    wire _0482_;
    wire new_Jinkela_wire_11046;
    wire new_Jinkela_wire_12331;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_10446;
    wire new_Jinkela_wire_5093;
    wire new_Jinkela_wire_11115;
    wire new_Jinkela_wire_4627;
    wire new_Jinkela_wire_4611;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_4487;
    wire new_Jinkela_wire_4050;
    wire _0185_;
    wire new_Jinkela_wire_11465;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_20621;
    wire _1677_;
    wire new_Jinkela_wire_2171;
    wire _0663_;
    wire new_Jinkela_wire_17031;
    wire new_Jinkela_wire_16310;
    wire new_Jinkela_wire_20637;
    wire new_Jinkela_wire_3444;
    wire new_Jinkela_wire_12448;
    wire new_Jinkela_wire_8302;
    wire new_Jinkela_wire_13346;
    wire new_Jinkela_wire_7325;
    wire _1137_;
    wire new_Jinkela_wire_8781;
    wire new_Jinkela_wire_11354;
    wire new_Jinkela_wire_9939;
    wire new_Jinkela_wire_4847;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_11070;
    wire new_Jinkela_wire_15845;
    wire new_Jinkela_wire_15598;
    wire new_Jinkela_wire_15441;
    wire new_Jinkela_wire_13613;
    wire new_Jinkela_wire_5830;
    wire _1582_;
    wire new_Jinkela_wire_10481;
    wire new_Jinkela_wire_17282;
    wire new_Jinkela_wire_1938;
    wire new_Jinkela_wire_12317;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_16934;
    wire new_Jinkela_wire_14585;
    wire new_Jinkela_wire_20463;
    wire new_Jinkela_wire_8444;
    wire new_Jinkela_wire_20184;
    wire new_Jinkela_wire_2563;
    wire new_Jinkela_wire_13411;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_1326;
    wire new_Jinkela_wire_12556;
    wire new_Jinkela_wire_7438;
    wire new_Jinkela_wire_4012;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_6645;
    wire _1522_;
    wire new_Jinkela_wire_5386;
    wire new_Jinkela_wire_19296;
    wire new_Jinkela_wire_12705;
    wire new_Jinkela_wire_3603;
    wire new_Jinkela_wire_21161;
    wire new_Jinkela_wire_8624;
    wire new_Jinkela_wire_8320;
    wire _0398_;
    wire new_Jinkela_wire_6878;
    wire new_Jinkela_wire_3606;
    wire new_Jinkela_wire_16980;
    wire new_Jinkela_wire_8621;
    wire _1565_;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_7369;
    wire new_Jinkela_wire_6717;
    wire new_Jinkela_wire_11958;
    wire new_Jinkela_wire_21222;
    wire new_Jinkela_wire_6626;
    wire new_Jinkela_wire_9989;
    wire _0040_;
    wire new_Jinkela_wire_4931;
    wire new_Jinkela_wire_3310;
    wire new_Jinkela_wire_3021;
    wire new_Jinkela_wire_5153;
    wire new_Jinkela_wire_9134;
    wire new_Jinkela_wire_8079;
    wire new_Jinkela_wire_19076;
    wire new_Jinkela_wire_3554;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_8485;
    wire _1766_;
    wire new_Jinkela_wire_4930;
    wire _0005_;
    wire new_Jinkela_wire_2333;
    wire new_Jinkela_wire_12184;
    wire new_Jinkela_wire_14595;
    wire new_Jinkela_wire_9432;
    wire new_Jinkela_wire_3568;
    wire new_Jinkela_wire_20167;
    wire new_Jinkela_wire_13625;
    wire new_Jinkela_wire_13134;
    wire new_Jinkela_wire_7914;
    wire new_Jinkela_wire_19157;
    wire new_Jinkela_wire_12610;
    wire new_Jinkela_wire_17882;
    wire new_Jinkela_wire_19709;
    wire new_Jinkela_wire_2028;
    wire new_Jinkela_wire_14899;
    wire new_Jinkela_wire_19295;
    wire new_Jinkela_wire_6838;
    wire new_Jinkela_wire_9356;
    wire new_Jinkela_wire_6689;
    wire new_Jinkela_wire_12917;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_13831;
    wire new_Jinkela_wire_18235;
    wire _0090_;
    wire new_Jinkela_wire_12942;
    wire new_Jinkela_wire_15771;
    wire new_Jinkela_wire_13632;
    wire new_Jinkela_wire_5509;
    wire new_Jinkela_wire_5140;
    wire new_Jinkela_wire_10390;
    wire new_Jinkela_wire_10820;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_7703;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_5811;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_5221;
    wire new_Jinkela_wire_4289;
    wire _0804_;
    wire new_Jinkela_wire_3472;
    wire new_Jinkela_wire_15123;
    wire _0384_;
    wire new_Jinkela_wire_17856;
    wire new_Jinkela_wire_4298;
    wire new_Jinkela_wire_2301;
    wire new_Jinkela_wire_13853;
    wire new_Jinkela_wire_18203;
    wire _0008_;
    wire new_Jinkela_wire_7570;
    wire new_Jinkela_wire_16714;
    wire new_Jinkela_wire_6233;
    wire new_Jinkela_wire_11019;
    wire new_Jinkela_wire_2471;
    wire new_Jinkela_wire_8511;
    wire new_Jinkela_wire_10912;
    wire new_Jinkela_wire_19451;
    wire new_Jinkela_wire_2223;
    wire new_Jinkela_wire_18532;
    wire new_Jinkela_wire_20096;
    wire new_Jinkela_wire_20562;
    wire new_Jinkela_wire_14298;
    wire new_Jinkela_wire_6057;
    wire new_Jinkela_wire_7110;
    wire new_Jinkela_wire_11060;
    wire new_Jinkela_wire_5707;
    wire new_Jinkela_wire_11640;
    wire new_Jinkela_wire_13063;
    wire _1309_;
    wire new_Jinkela_wire_12272;
    wire new_Jinkela_wire_17315;
    wire new_Jinkela_wire_12511;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_7937;
    wire new_Jinkela_wire_14327;
    wire new_Jinkela_wire_2496;
    wire _1160_;
    wire new_Jinkela_wire_12831;
    wire new_Jinkela_wire_5882;
    wire new_Jinkela_wire_13369;
    wire new_Jinkela_wire_9153;
    wire new_Jinkela_wire_4141;
    wire new_Jinkela_wire_20740;
    wire new_Jinkela_wire_12851;
    wire new_Jinkela_wire_6940;
    wire new_Jinkela_wire_18466;
    wire new_Jinkela_wire_11831;
    wire new_Jinkela_wire_16873;
    wire new_Jinkela_wire_15829;
    wire new_Jinkela_wire_13847;
    wire new_Jinkela_wire_18583;
    wire new_Jinkela_wire_5395;
    wire new_Jinkela_wire_17844;
    wire new_Jinkela_wire_11133;
    wire new_Jinkela_wire_9978;
    wire new_Jinkela_wire_11926;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_6212;
    wire new_Jinkela_wire_4068;
    wire new_Jinkela_wire_12586;
    wire new_Jinkela_wire_4240;
    wire new_Jinkela_wire_3034;
    wire new_Jinkela_wire_16731;
    wire new_Jinkela_wire_18917;
    wire new_Jinkela_wire_20308;
    wire new_Jinkela_wire_13681;
    wire new_Jinkela_wire_13849;
    wire new_Jinkela_wire_13797;
    wire new_Jinkela_wire_20762;
    wire new_Jinkela_wire_20912;
    wire new_Jinkela_wire_21240;
    wire new_Jinkela_wire_3878;
    wire new_Jinkela_wire_15479;
    wire new_Jinkela_wire_19542;
    wire new_Jinkela_wire_6149;
    wire new_Jinkela_wire_12174;
    wire new_Jinkela_wire_4017;
    wire new_Jinkela_wire_14428;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_13651;
    wire new_Jinkela_wire_19265;
    wire new_Jinkela_wire_6684;
    wire new_Jinkela_wire_11464;
    wire new_Jinkela_wire_5875;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_12584;
    wire new_Jinkela_wire_14776;
    wire new_Jinkela_wire_11372;
    wire _0165_;
    wire new_Jinkela_wire_5223;
    wire new_Jinkela_wire_9081;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_4795;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_19291;
    wire new_Jinkela_wire_3881;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_11611;
    wire new_Jinkela_wire_3611;
    wire new_Jinkela_wire_9316;
    wire new_Jinkela_wire_2656;
    wire new_Jinkela_wire_14200;
    wire new_Jinkela_wire_16791;
    wire new_Jinkela_wire_4642;
    wire _1438_;
    wire new_Jinkela_wire_6407;
    wire new_Jinkela_wire_12358;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_19127;
    wire new_Jinkela_wire_19743;
    wire new_Jinkela_wire_17020;
    wire new_Jinkela_wire_7831;
    wire new_Jinkela_wire_8101;
    wire new_Jinkela_wire_10804;
    wire new_Jinkela_wire_6901;
    wire new_Jinkela_wire_5771;
    wire new_Jinkela_wire_17955;
    wire new_Jinkela_wire_20253;
    wire new_Jinkela_wire_5379;
    wire new_Jinkela_wire_19346;
    wire new_Jinkela_wire_18460;
    wire new_Jinkela_wire_12651;
    wire new_Jinkela_wire_20342;
    wire new_Jinkela_wire_18114;
    wire new_Jinkela_wire_4029;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_15934;
    wire new_Jinkela_wire_12948;
    wire new_Jinkela_wire_9093;
    wire new_Jinkela_wire_5740;
    wire new_Jinkela_wire_18497;
    wire new_Jinkela_wire_9801;
    wire new_Jinkela_wire_19257;
    wire new_Jinkela_wire_15210;
    wire new_Jinkela_wire_20967;
    wire new_Jinkela_wire_9372;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_16242;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_18004;
    wire new_Jinkela_wire_6593;
    wire new_Jinkela_wire_13064;
    wire new_Jinkela_wire_8857;
    wire new_Jinkela_wire_11514;
    wire new_Jinkela_wire_5433;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_18372;
    wire new_Jinkela_wire_3619;
    wire new_Jinkela_wire_3372;
    wire new_Jinkela_wire_7848;
    wire new_Jinkela_wire_5869;
    wire new_Jinkela_wire_10782;
    wire new_Jinkela_wire_16869;
    wire new_Jinkela_wire_18543;
    wire _1027_;
    wire new_Jinkela_wire_3690;
    wire new_Jinkela_wire_9031;
    wire new_Jinkela_wire_17570;
    wire new_Jinkela_wire_6595;
    wire new_Jinkela_wire_2249;
    wire _0133_;
    wire new_Jinkela_wire_4623;
    wire new_Jinkela_wire_12097;
    wire new_Jinkela_wire_16061;
    wire new_Jinkela_wire_19287;
    wire new_Jinkela_wire_16385;
    wire new_Jinkela_wire_9606;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_12605;
    wire new_Jinkela_wire_17677;
    wire new_Jinkela_wire_18143;
    wire new_Jinkela_wire_6398;
    wire new_Jinkela_wire_16436;
    wire new_Jinkela_wire_9059;
    wire new_Jinkela_wire_18165;
    wire new_Jinkela_wire_4142;
    wire new_Jinkela_wire_4203;
    wire new_Jinkela_wire_10387;
    wire _1145_;
    wire new_Jinkela_wire_13706;
    wire new_Jinkela_wire_18888;
    wire new_Jinkela_wire_14371;
    wire new_Jinkela_wire_4098;
    wire new_Jinkela_wire_6420;
    wire new_Jinkela_wire_14647;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_9865;
    wire new_Jinkela_wire_4778;
    wire new_Jinkela_wire_20876;
    wire new_Jinkela_wire_17936;
    wire new_Jinkela_wire_7943;
    wire new_Jinkela_wire_7992;
    wire new_Jinkela_wire_15025;
    wire new_Jinkela_wire_2175;
    wire new_Jinkela_wire_6177;
    wire new_Jinkela_wire_14491;
    wire new_Jinkela_wire_18797;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_4148;
    wire new_Jinkela_wire_2414;
    wire new_Jinkela_wire_12009;
    wire new_Jinkela_wire_13238;
    wire new_Jinkela_wire_4746;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_2536;
    wire new_Jinkela_wire_20395;
    wire new_Jinkela_wire_2046;
    wire _0504_;
    wire new_Jinkela_wire_15234;
    wire new_Jinkela_wire_17839;
    wire new_Jinkela_wire_7469;
    wire new_Jinkela_wire_15337;
    wire new_Jinkela_wire_5821;
    wire new_Jinkela_wire_8222;
    wire new_Jinkela_wire_12040;
    wire new_Jinkela_wire_3682;
    wire new_Jinkela_wire_18622;
    wire new_Jinkela_wire_16454;
    wire new_Jinkela_wire_5472;
    wire new_Jinkela_wire_16414;
    wire new_Jinkela_wire_6986;
    wire new_Jinkela_wire_10933;
    wire new_Jinkela_wire_14836;
    wire new_Jinkela_wire_19101;
    wire new_Jinkela_wire_11353;
    wire _1563_;
    wire new_Jinkela_wire_8791;
    wire new_Jinkela_wire_4939;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_7638;
    wire new_Jinkela_wire_14338;
    wire new_Jinkela_wire_2250;
    wire new_Jinkela_wire_14622;
    wire new_Jinkela_wire_7773;
    wire new_Jinkela_wire_11324;
    wire _0197_;
    wire new_Jinkela_wire_11861;
    wire new_Jinkela_wire_18610;
    wire new_Jinkela_wire_4838;
    wire new_Jinkela_wire_10374;
    wire new_Jinkela_wire_13008;
    wire new_Jinkela_wire_19377;
    wire new_Jinkela_wire_16278;
    wire new_Jinkela_wire_11315;
    wire new_Jinkela_wire_4418;
    wire new_Jinkela_wire_20959;
    wire new_Jinkela_wire_20189;
    wire new_Jinkela_wire_4366;
    wire new_Jinkela_wire_7079;
    wire new_Jinkela_wire_10703;
    wire new_Jinkela_wire_4530;
    wire new_Jinkela_wire_19912;
    wire new_Jinkela_wire_10037;
    wire new_Jinkela_wire_2526;
    wire new_Jinkela_wire_10598;
    wire new_Jinkela_wire_14656;
    wire new_Jinkela_wire_5169;
    wire new_Jinkela_wire_12148;
    wire _1725_;
    wire new_Jinkela_wire_19622;
    wire new_Jinkela_wire_5437;
    wire new_Jinkela_wire_20901;
    wire _1391_;
    wire new_Jinkela_wire_12362;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_17171;
    wire new_Jinkela_wire_9739;
    wire new_Jinkela_wire_2594;
    wire new_Jinkela_wire_9782;
    wire new_Jinkela_wire_11367;
    wire new_Jinkela_wire_4969;
    wire new_Jinkela_wire_16030;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_13465;
    wire new_Jinkela_wire_16985;
    wire new_Jinkela_wire_8066;
    wire new_Jinkela_wire_6841;
    wire new_Jinkela_wire_13240;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_16923;
    wire new_Jinkela_wire_10822;
    wire new_Jinkela_wire_9768;
    wire new_Jinkela_wire_18429;
    wire new_Jinkela_wire_5419;
    wire new_Jinkela_wire_17908;
    wire new_Jinkela_wire_17652;
    wire new_Jinkela_wire_16109;
    wire new_Jinkela_wire_19628;
    wire new_Jinkela_wire_17679;
    wire new_Jinkela_wire_5837;
    wire new_Jinkela_wire_14562;
    wire new_Jinkela_wire_19494;
    wire _1501_;
    wire new_Jinkela_wire_17188;
    wire new_Jinkela_wire_9091;
    wire new_Jinkela_wire_12390;
    wire new_Jinkela_wire_12215;
    wire new_Jinkela_wire_3193;
    wire new_Jinkela_wire_15616;
    wire new_Jinkela_wire_16257;
    wire _1707_;
    wire new_Jinkela_wire_6570;
    wire new_Jinkela_wire_12019;
    wire new_Jinkela_wire_4501;
    wire new_Jinkela_wire_1918;
    wire new_Jinkela_wire_13248;
    wire new_Jinkela_wire_6385;
    wire new_Jinkela_wire_7071;
    wire _0020_;
    wire new_Jinkela_wire_8911;
    wire new_Jinkela_wire_8426;
    wire new_Jinkela_wire_19706;
    wire new_Jinkela_wire_16744;
    wire new_Jinkela_wire_13754;
    wire new_Jinkela_wire_4317;
    wire new_Jinkela_wire_2411;
    wire new_Jinkela_wire_19804;
    wire new_Jinkela_wire_14799;
    wire _1085_;
    wire _0880_;
    wire new_Jinkela_wire_4124;
    wire new_Jinkela_wire_15555;
    wire new_Jinkela_wire_5176;
    wire new_Jinkela_wire_1705;
    wire _1699_;
    wire new_Jinkela_wire_6517;
    wire new_Jinkela_wire_17530;
    wire new_Jinkela_wire_14423;
    wire new_Jinkela_wire_16220;
    wire new_Jinkela_wire_1693;
    wire new_Jinkela_wire_4301;
    wire new_Jinkela_wire_20424;
    wire new_Jinkela_wire_20609;
    wire new_Jinkela_wire_2248;
    wire new_Jinkela_wire_17970;
    wire new_Jinkela_wire_11880;
    wire new_Jinkela_wire_20413;
    wire new_Jinkela_wire_8102;
    wire new_Jinkela_wire_17637;
    wire new_Jinkela_wire_2511;
    wire new_Jinkela_wire_7243;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_19657;
    wire new_Jinkela_wire_11244;
    wire new_Jinkela_wire_7777;
    wire new_Jinkela_wire_19767;
    wire new_Jinkela_wire_1666;
    wire new_Jinkela_wire_4741;
    wire new_Jinkela_wire_9688;
    wire new_Jinkela_wire_20515;
    wire new_Jinkela_wire_21235;
    wire new_Jinkela_wire_7003;
    wire new_Jinkela_wire_17896;
    wire _0120_;
    wire new_Jinkela_wire_8521;
    wire new_Jinkela_wire_9643;
    wire new_Jinkela_wire_19443;
    wire new_Jinkela_wire_13997;
    wire new_Jinkela_wire_13036;
    wire new_Jinkela_wire_4176;
    wire _1153_;
    wire new_Jinkela_wire_3125;
    wire new_Jinkela_wire_18319;
    wire new_Jinkela_wire_1907;
    wire new_Jinkela_wire_17080;
    wire new_Jinkela_wire_7382;
    wire new_Jinkela_wire_3307;
    wire new_Jinkela_wire_4975;
    wire new_Jinkela_wire_17428;
    wire new_Jinkela_wire_9586;
    wire new_Jinkela_wire_3373;
    wire new_Jinkela_wire_10566;
    wire new_Jinkela_wire_9704;
    wire new_Jinkela_wire_4336;
    wire new_Jinkela_wire_7323;
    wire new_Jinkela_wire_16503;
    wire new_Jinkela_wire_14851;
    wire new_Jinkela_wire_11120;
    wire new_Jinkela_wire_14059;
    wire new_Jinkela_wire_6221;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_9088;
    wire new_Jinkela_wire_5019;
    wire new_Jinkela_wire_8718;
    wire new_Jinkela_wire_6448;
    wire new_Jinkela_wire_958;
    wire _0156_;
    wire new_Jinkela_wire_10927;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_17410;
    wire new_Jinkela_wire_1777;
    wire new_Jinkela_wire_3149;
    wire new_Jinkela_wire_18601;
    wire new_Jinkela_wire_16152;
    wire new_Jinkela_wire_18658;
    wire new_Jinkela_wire_12006;
    wire new_Jinkela_wire_2798;
    wire new_Jinkela_wire_11633;
    wire new_Jinkela_wire_7124;
    wire new_Jinkela_wire_15947;
    wire new_Jinkela_wire_1780;
    wire new_Jinkela_wire_10410;
    wire new_Jinkela_wire_13550;
    wire new_Jinkela_wire_15815;
    wire new_Jinkela_wire_2186;
    wire _1358_;
    wire new_Jinkela_wire_4030;
    wire new_Jinkela_wire_17507;
    wire new_Jinkela_wire_15207;
    wire new_Jinkela_wire_11954;
    wire new_Jinkela_wire_16993;
    wire _1581_;
    wire new_Jinkela_wire_11408;
    wire new_Jinkela_wire_16204;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_4680;
    wire new_Jinkela_wire_5251;
    wire new_Jinkela_wire_3872;
    wire _1477_;
    wire new_Jinkela_wire_5204;
    wire new_Jinkela_wire_13574;
    wire new_Jinkela_wire_19985;
    wire new_Jinkela_wire_21052;
    wire new_Jinkela_wire_8930;
    wire _0968_;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_19652;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_18243;
    wire new_Jinkela_wire_17139;
    wire new_Jinkela_wire_7162;
    wire new_Jinkela_wire_15223;
    wire new_Jinkela_wire_13943;
    wire new_Jinkela_wire_7483;
    wire new_Jinkela_wire_2092;
    wire new_Jinkela_wire_12190;
    wire new_Jinkela_wire_8601;
    wire new_Jinkela_wire_10555;
    wire new_Jinkela_wire_6113;
    wire new_Jinkela_wire_11273;
    wire new_Jinkela_wire_1852;
    wire new_Jinkela_wire_4973;
    wire new_Jinkela_wire_16813;
    wire new_Jinkela_wire_15503;
    wire new_Jinkela_wire_5185;
    wire new_Jinkela_wire_10029;
    wire new_Jinkela_wire_11906;
    wire new_Jinkela_wire_20951;
    wire new_Jinkela_wire_16553;
    wire new_Jinkela_wire_21127;
    wire new_Jinkela_wire_14816;
    wire new_Jinkela_wire_17324;
    wire new_Jinkela_wire_14556;
    wire new_Jinkela_wire_19136;
    wire new_Jinkela_wire_10156;
    wire new_Jinkela_wire_4618;
    wire new_Jinkela_wire_8408;
    wire new_Jinkela_wire_10393;
    wire new_Jinkela_wire_16098;
    wire _1294_;
    wire _1587_;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_7509;
    wire new_Jinkela_wire_11871;
    wire new_Jinkela_wire_19227;
    wire new_Jinkela_wire_10837;
    wire new_Jinkela_wire_18449;
    wire new_Jinkela_wire_9562;
    wire _0980_;
    wire new_Jinkela_wire_14866;
    wire new_Jinkela_wire_2618;
    wire new_Jinkela_wire_9822;
    wire new_Jinkela_wire_16022;
    wire new_Jinkela_wire_13082;
    wire new_Jinkela_wire_12243;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_4668;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_13403;
    wire new_net_3968;
    wire new_Jinkela_wire_4542;
    wire new_Jinkela_wire_13752;
    wire new_Jinkela_wire_17915;
    wire new_Jinkela_wire_2692;
    wire new_Jinkela_wire_20632;
    wire new_Jinkela_wire_11021;
    wire _0462_;
    wire new_Jinkela_wire_14326;
    wire _1700_;
    wire new_Jinkela_wire_18008;
    wire new_Jinkela_wire_19989;
    wire new_Jinkela_wire_6294;
    wire new_Jinkela_wire_8713;
    wire new_Jinkela_wire_7872;
    wire new_Jinkela_wire_7745;
    wire _0347_;
    wire _1669_;
    wire new_Jinkela_wire_3429;
    wire new_Jinkela_wire_2793;
    wire new_Jinkela_wire_20851;
    wire new_Jinkela_wire_16897;
    wire new_Jinkela_wire_17801;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_5663;
    wire new_Jinkela_wire_9013;
    wire _0322_;
    wire new_Jinkela_wire_12786;
    wire new_Jinkela_wire_5224;
    wire new_Jinkela_wire_20567;
    wire new_Jinkela_wire_18650;
    wire new_Jinkela_wire_21246;
    wire new_Jinkela_wire_4768;
    wire new_Jinkela_wire_18801;
    wire new_Jinkela_wire_17129;
    wire new_Jinkela_wire_9983;
    wire _0339_;
    wire new_Jinkela_wire_21233;
    wire new_Jinkela_wire_20183;
    wire new_Jinkela_wire_6965;
    wire new_Jinkela_wire_4928;
    wire new_Jinkela_wire_20568;
    wire new_Jinkela_wire_3692;
    wire new_Jinkela_wire_18882;
    wire new_Jinkela_wire_8392;
    wire new_Jinkela_wire_7768;
    wire new_Jinkela_wire_5022;
    wire new_Jinkela_wire_11739;
    wire new_Jinkela_wire_19270;
    wire new_Jinkela_wire_11506;
    wire _1072_;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_10870;
    wire new_Jinkela_wire_3695;
    wire new_Jinkela_wire_8647;
    wire new_Jinkela_wire_16294;
    wire _0029_;
    wire new_Jinkela_wire_7802;
    wire new_Jinkela_wire_8634;
    wire _1457_;
    wire new_Jinkela_wire_4118;
    wire new_Jinkela_wire_16127;
    wire new_Jinkela_wire_2672;
    wire new_Jinkela_wire_15580;
    wire new_Jinkela_wire_4168;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_8016;
    wire new_Jinkela_wire_6397;
    wire new_Jinkela_wire_12554;
    wire _1680_;
    wire new_Jinkela_wire_3434;
    wire new_Jinkela_wire_17110;
    wire _0935_;
    wire new_Jinkela_wire_2147;
    wire new_Jinkela_wire_14808;
    wire new_Jinkela_wire_13095;
    wire new_Jinkela_wire_3912;
    wire new_Jinkela_wire_18684;
    wire new_Jinkela_wire_4236;
    wire new_Jinkela_wire_19851;
    wire new_Jinkela_wire_5853;
    wire _1313_;
    wire new_Jinkela_wire_19564;
    wire new_Jinkela_wire_13004;
    wire new_Jinkela_wire_8888;
    wire new_Jinkela_wire_10563;
    wire new_Jinkela_wire_4629;
    wire new_Jinkela_wire_6727;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_7900;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_19068;
    wire new_Jinkela_wire_6642;
    wire new_Jinkela_wire_9220;
    wire new_Jinkela_wire_4362;
    wire new_Jinkela_wire_3801;
    wire _0973_;
    wire new_Jinkela_wire_19668;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_15356;
    wire new_Jinkela_wire_17293;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_3877;
    wire new_Jinkela_wire_15811;
    wire new_Jinkela_wire_12242;
    wire new_Jinkela_wire_12069;
    wire new_Jinkela_wire_9107;
    wire new_Jinkela_wire_10740;
    wire new_Jinkela_wire_20729;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_19045;
    wire new_Jinkela_wire_16394;
    wire new_Jinkela_wire_13934;
    wire new_Jinkela_wire_7668;
    wire new_Jinkela_wire_20478;
    wire new_Jinkela_wire_4878;
    wire new_Jinkela_wire_11121;
    wire new_Jinkela_wire_12569;
    wire new_Jinkela_wire_13820;
    wire new_Jinkela_wire_17758;
    wire new_Jinkela_wire_19830;
    wire _1620_;
    wire new_Jinkela_wire_12382;
    wire new_Jinkela_wire_3627;
    wire new_Jinkela_wire_13725;
    wire new_Jinkela_wire_17792;
    wire new_Jinkela_wire_10768;
    wire new_Jinkela_wire_14650;
    wire new_Jinkela_wire_9649;
    wire new_Jinkela_wire_20510;
    wire new_Jinkela_wire_7652;
    wire new_Jinkela_wire_10806;
    wire new_Jinkela_wire_10556;
    wire _1325_;
    wire new_Jinkela_wire_15604;
    wire new_Jinkela_wire_11516;
    wire new_Jinkela_wire_18139;
    wire new_Jinkela_wire_6958;
    wire new_Jinkela_wire_16674;
    wire new_Jinkela_wire_2947;
    wire new_Jinkela_wire_13367;
    wire new_Jinkela_wire_20862;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_11982;
    wire new_Jinkela_wire_13733;
    wire new_Jinkela_wire_10587;
    wire new_Jinkela_wire_17881;
    wire new_Jinkela_wire_11441;
    wire _1764_;
    wire new_Jinkela_wire_1055;
    wire new_Jinkela_wire_7677;
    wire new_Jinkela_wire_13191;
    wire new_Jinkela_wire_4481;
    wire new_Jinkela_wire_7711;
    wire new_Jinkela_wire_7862;
    wire new_Jinkela_wire_14903;
    wire new_Jinkela_wire_13504;
    wire new_Jinkela_wire_5256;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_16184;
    wire new_Jinkela_wire_12920;
    wire new_Jinkela_wire_7754;
    wire _0289_;
    wire new_Jinkela_wire_11509;
    wire new_Jinkela_wire_9783;
    wire new_Jinkela_wire_9069;
    wire new_Jinkela_wire_19737;
    wire new_Jinkela_wire_14777;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_19374;
    wire new_Jinkela_wire_1057;
    wire new_Jinkela_wire_15905;
    wire new_Jinkela_wire_7792;
    wire new_Jinkela_wire_5965;
    wire _0762_;
    wire new_Jinkela_wire_2101;
    wire new_Jinkela_wire_7319;
    wire new_Jinkela_wire_17061;
    wire new_Jinkela_wire_15731;
    wire new_Jinkela_wire_5216;
    wire new_Jinkela_wire_15189;
    wire new_Jinkela_wire_14555;
    wire new_Jinkela_wire_15315;
    wire _0864_;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_8004;
    wire new_Jinkela_wire_11896;
    wire new_Jinkela_wire_5036;
    wire new_Jinkela_wire_8463;
    wire new_Jinkela_wire_14427;
    wire new_Jinkela_wire_11077;
    wire new_Jinkela_wire_13438;
    wire new_Jinkela_wire_14403;
    wire new_Jinkela_wire_3200;
    wire new_Jinkela_wire_5572;
    wire new_Jinkela_wire_6908;
    wire new_Jinkela_wire_21328;
    wire new_Jinkela_wire_6048;
    wire new_Jinkela_wire_20833;
    wire new_Jinkela_wire_19420;
    wire new_Jinkela_wire_2961;
    wire new_Jinkela_wire_6676;
    wire new_Jinkela_wire_2017;
    wire new_Jinkela_wire_12778;
    wire new_Jinkela_wire_3215;
    wire new_Jinkela_wire_9395;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_20855;
    wire new_Jinkela_wire_18169;
    wire new_Jinkela_wire_10177;
    wire new_Jinkela_wire_11263;
    wire new_Jinkela_wire_9641;
    wire new_Jinkela_wire_8919;
    wire new_Jinkela_wire_8894;
    wire new_Jinkela_wire_13967;
    wire new_Jinkela_wire_5368;
    wire new_Jinkela_wire_8812;
    wire new_Jinkela_wire_3741;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_4344;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_1245;
    wire _1834_;
    wire new_Jinkela_wire_1719;
    wire _0645_;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_11662;
    wire new_Jinkela_wire_13692;
    wire _0889_;
    wire new_Jinkela_wire_7975;
    wire new_Jinkela_wire_2822;
    wire new_Jinkela_wire_9771;
    wire new_Jinkela_wire_9094;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_14579;
    wire new_Jinkela_wire_15286;
    wire _0539_;
    wire new_Jinkela_wire_8192;
    wire new_Jinkela_wire_19871;
    wire _1704_;
    wire new_Jinkela_wire_14637;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_13595;
    wire new_Jinkela_wire_4697;
    wire new_Jinkela_wire_14465;
    wire new_Jinkela_wire_4323;
    wire new_Jinkela_wire_18028;
    wire new_Jinkela_wire_15816;
    wire new_Jinkela_wire_4663;
    wire new_Jinkela_wire_5551;
    wire new_Jinkela_wire_4890;
    wire new_Jinkela_wire_9234;
    wire new_Jinkela_wire_13615;
    wire new_Jinkela_wire_5255;
    wire _0189_;
    wire new_Jinkela_wire_2317;
    wire new_Jinkela_wire_5124;
    wire new_Jinkela_wire_13323;
    wire new_Jinkela_wire_15992;
    wire new_Jinkela_wire_19571;
    wire new_Jinkela_wire_6155;
    wire _1404_;
    wire new_Jinkela_wire_9934;
    wire new_Jinkela_wire_20716;
    wire new_Jinkela_wire_9332;
    wire new_Jinkela_wire_9903;
    wire new_Jinkela_wire_13279;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_9533;
    wire new_Jinkela_wire_15940;
    wire new_Jinkela_wire_13206;
    wire new_Jinkela_wire_16759;
    wire new_Jinkela_wire_6241;
    wire new_Jinkela_wire_14608;
    wire new_Jinkela_wire_12235;
    wire new_Jinkela_wire_2841;
    wire new_Jinkela_wire_13516;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_14166;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_13233;
    wire _0014_;
    wire new_Jinkela_wire_14937;
    wire new_Jinkela_wire_19894;
    wire new_Jinkela_wire_3925;
    wire new_Jinkela_wire_10299;
    wire new_Jinkela_wire_6350;
    wire new_Jinkela_wire_20198;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_6336;
    wire new_Jinkela_wire_6617;
    wire new_Jinkela_wire_11240;
    wire new_Jinkela_wire_6572;
    wire new_Jinkela_wire_13157;
    wire new_Jinkela_wire_2133;
    wire new_Jinkela_wire_10137;
    wire new_Jinkela_wire_11809;
    wire new_Jinkela_wire_9274;
    wire new_Jinkela_wire_18799;
    wire new_Jinkela_wire_14545;
    wire new_Jinkela_wire_9640;
    wire new_Jinkela_wire_8838;
    wire _1633_;
    wire new_Jinkela_wire_8899;
    wire new_Jinkela_wire_17604;
    wire new_Jinkela_wire_12297;
    wire new_Jinkela_wire_21101;
    wire new_Jinkela_wire_5375;
    wire new_Jinkela_wire_12353;
    wire new_Jinkela_wire_12889;
    wire new_Jinkela_wire_12381;
    wire new_Jinkela_wire_18295;
    wire new_Jinkela_wire_16758;
    wire new_Jinkela_wire_7655;
    wire new_Jinkela_wire_1866;
    wire new_Jinkela_wire_10005;
    wire new_Jinkela_wire_19604;
    wire _0288_;
    wire new_Jinkela_wire_17177;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_17536;
    wire new_Jinkela_wire_15008;
    wire new_Jinkela_wire_1726;
    wire new_Jinkela_wire_20929;
    wire new_Jinkela_wire_18477;
    wire _0366_;
    wire _1252_;
    wire new_Jinkela_wire_6041;
    wire new_Jinkela_wire_9835;
    wire new_Jinkela_wire_19813;
    wire new_Jinkela_wire_3602;
    wire new_Jinkela_wire_9252;
    wire new_Jinkela_wire_17860;
    wire new_Jinkela_wire_1767;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_14713;
    wire new_Jinkela_wire_3301;
    wire new_Jinkela_wire_6679;
    wire new_Jinkela_wire_5683;
    wire new_Jinkela_wire_7868;
    wire new_Jinkela_wire_11997;
    wire new_Jinkela_wire_19896;
    wire new_Jinkela_wire_6966;
    wire new_Jinkela_wire_12477;
    wire new_Jinkela_wire_19666;
    wire _0975_;
    wire new_Jinkela_wire_16100;
    wire new_Jinkela_wire_13319;
    wire new_Jinkela_wire_2740;
    wire new_Jinkela_wire_5377;
    wire new_Jinkela_wire_19149;
    wire new_Jinkela_wire_18565;
    wire new_Jinkela_wire_17924;
    wire new_Jinkela_wire_16870;
    wire new_Jinkela_wire_8118;
    wire new_Jinkela_wire_20127;
    wire new_Jinkela_wire_6798;
    wire new_Jinkela_wire_15883;
    wire new_Jinkela_wire_11430;
    wire new_Jinkela_wire_7821;
    wire new_Jinkela_wire_13970;
    wire new_Jinkela_wire_5397;
    wire new_Jinkela_wire_18853;
    wire new_Jinkela_wire_6504;
    wire new_Jinkela_wire_20306;
    wire new_Jinkela_wire_2405;
    wire new_Jinkela_wire_15398;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_15846;
    wire new_Jinkela_wire_2267;
    wire new_Jinkela_wire_19992;
    wire new_Jinkela_wire_12189;
    wire new_Jinkela_wire_18954;
    wire new_Jinkela_wire_9010;
    wire new_Jinkela_wire_6947;
    wire _1771_;
    wire new_Jinkela_wire_17362;
    wire new_Jinkela_wire_5407;
    wire new_Jinkela_wire_4599;
    wire new_Jinkela_wire_5810;
    wire new_Jinkela_wire_19798;
    wire new_Jinkela_wire_6660;
    wire new_Jinkela_wire_17058;
    wire new_Jinkela_wire_13179;
    wire new_Jinkela_wire_13679;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_15813;
    wire new_Jinkela_wire_20985;
    wire new_Jinkela_wire_15570;
    wire new_Jinkela_wire_7182;
    wire new_Jinkela_wire_18868;
    wire new_Jinkela_wire_15800;
    wire new_Jinkela_wire_14073;
    wire new_Jinkela_wire_9496;
    wire new_Jinkela_wire_6133;
    wire new_Jinkela_wire_13953;
    wire new_Jinkela_wire_20301;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_10995;
    wire _1331_;
    wire _0006_;
    wire new_Jinkela_wire_16263;
    wire _1373_;
    wire new_Jinkela_wire_5899;
    wire new_Jinkela_wire_9307;
    wire new_Jinkela_wire_21019;
    wire new_Jinkela_wire_21079;
    wire new_Jinkela_wire_3424;
    wire new_Jinkela_wire_4143;
    wire new_Jinkela_wire_2958;
    wire new_Jinkela_wire_2730;
    wire new_Jinkela_wire_17516;
    wire new_Jinkela_wire_15472;
    wire new_Jinkela_wire_18713;
    wire new_Jinkela_wire_4991;
    wire new_Jinkela_wire_15901;
    wire new_Jinkela_wire_19333;
    wire new_Jinkela_wire_14202;
    wire new_Jinkela_wire_13353;
    wire new_Jinkela_wire_9916;
    wire new_Jinkela_wire_18849;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_14606;
    wire new_Jinkela_wire_15987;
    wire new_Jinkela_wire_13359;
    wire _1284_;
    wire new_Jinkela_wire_4096;
    wire new_Jinkela_wire_13984;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_8123;
    wire new_Jinkela_wire_12992;
    wire new_Jinkela_wire_18347;
    wire new_Jinkela_wire_17564;
    wire new_Jinkela_wire_20145;
    wire new_Jinkela_wire_10793;
    wire new_Jinkela_wire_6692;
    wire new_Jinkela_wire_12935;
    wire new_Jinkela_wire_4586;
    wire new_Jinkela_wire_14141;
    wire new_Jinkela_wire_17474;
    wire _1717_;
    wire new_Jinkela_wire_8204;
    wire new_Jinkela_wire_5596;
    wire new_Jinkela_wire_15021;
    wire new_Jinkela_wire_16395;
    wire new_Jinkela_wire_4140;
    wire new_Jinkela_wire_18079;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_3658;
    wire new_Jinkela_wire_9382;
    wire new_Jinkela_wire_2868;
    wire new_Jinkela_wire_14388;
    wire new_Jinkela_wire_2466;
    wire new_Jinkela_wire_8961;
    wire _1267_;
    wire new_Jinkela_wire_15374;
    wire new_Jinkela_wire_21251;
    wire new_Jinkela_wire_8078;
    wire new_Jinkela_wire_3165;
    wire new_Jinkela_wire_9367;
    wire new_Jinkela_wire_19372;
    wire new_Jinkela_wire_18552;
    wire new_Jinkela_wire_8360;
    wire new_Jinkela_wire_3231;
    wire new_Jinkela_wire_16916;
    wire new_Jinkela_wire_3691;
    wire new_Jinkela_wire_7828;
    wire new_Jinkela_wire_19087;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_7558;
    wire _1098_;
    wire new_Jinkela_wire_4760;
    wire new_Jinkela_wire_7537;
    wire new_Jinkela_wire_7313;
    wire new_Jinkela_wire_12540;
    wire new_Jinkela_wire_16821;
    wire new_Jinkela_wire_7930;
    wire new_Jinkela_wire_8150;
    wire new_Jinkela_wire_2501;
    wire new_Jinkela_wire_3675;
    wire new_Jinkela_wire_11484;
    wire new_Jinkela_wire_10128;
    wire new_Jinkela_wire_13376;
    wire new_Jinkela_wire_19748;
    wire new_Jinkela_wire_9703;
    wire new_Jinkela_wire_17901;
    wire new_Jinkela_wire_10204;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_18189;
    wire new_Jinkela_wire_18822;
    wire new_Jinkela_wire_12376;
    wire new_Jinkela_wire_15018;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_13646;
    wire new_Jinkela_wire_8673;
    wire _1561_;
    wire new_Jinkela_wire_14953;
    wire new_Jinkela_wire_2204;
    wire new_Jinkela_wire_12525;
    wire new_Jinkela_wire_15500;
    wire new_Jinkela_wire_3616;
    wire _1436_;
    wire new_Jinkela_wire_14735;
    wire new_Jinkela_wire_9842;
    wire _0291_;
    wire new_Jinkela_wire_10713;
    wire new_Jinkela_wire_4641;
    wire new_Jinkela_wire_18354;
    wire new_Jinkela_wire_12500;
    wire new_Jinkela_wire_5743;
    wire new_Jinkela_wire_9570;
    wire new_Jinkela_wire_9102;
    wire new_Jinkela_wire_3911;
    wire new_Jinkela_wire_1651;
    wire _0227_;
    wire new_Jinkela_wire_1317;
    wire _1019_;
    wire new_Jinkela_wire_11264;
    wire new_Jinkela_wire_8586;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_15847;
    wire new_Jinkela_wire_4662;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_17700;
    wire new_Jinkela_wire_10671;
    wire new_Jinkela_wire_2421;
    wire new_Jinkela_wire_15639;
    wire new_Jinkela_wire_18554;
    wire new_Jinkela_wire_8684;
    wire _0756_;
    wire new_Jinkela_wire_10727;
    wire new_Jinkela_wire_15122;
    wire new_Jinkela_wire_14280;
    wire new_Jinkela_wire_3696;
    wire new_Jinkela_wire_9439;
    wire new_Jinkela_wire_5569;
    wire new_Jinkela_wire_8922;
    wire new_Jinkela_wire_13601;
    wire new_Jinkela_wire_8741;
    wire new_Jinkela_wire_19464;
    wire new_Jinkela_wire_20766;
    wire new_Jinkela_wire_11239;
    wire new_Jinkela_wire_20099;
    wire new_Jinkela_wire_2878;
    wire new_Jinkela_wire_2278;
    wire new_Jinkela_wire_11807;
    wire new_Jinkela_wire_3808;
    wire new_Jinkela_wire_15903;
    wire new_Jinkela_wire_7526;
    wire new_Jinkela_wire_2794;
    wire new_Jinkela_wire_20532;
    wire new_Jinkela_wire_2265;
    wire new_Jinkela_wire_4587;
    wire new_Jinkela_wire_18563;
    wire new_Jinkela_wire_7530;
    wire _1826_;
    wire new_Jinkela_wire_17485;
    wire new_Jinkela_wire_17486;
    wire new_Jinkela_wire_19492;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_19552;
    wire new_Jinkela_wire_3615;
    wire new_Jinkela_wire_12805;
    wire new_Jinkela_wire_9571;
    wire new_Jinkela_wire_11963;
    wire new_Jinkela_wire_6097;
    wire _0657_;
    wire new_Jinkela_wire_3141;
    wire new_Jinkela_wire_10716;
    wire new_Jinkela_wire_8334;
    wire new_Jinkela_wire_21016;
    wire new_Jinkela_wire_4595;
    wire new_Jinkela_wire_17051;
    wire new_Jinkela_wire_11457;
    wire new_Jinkela_wire_17859;
    wire new_Jinkela_wire_7739;
    wire new_Jinkela_wire_6795;
    wire new_Jinkela_wire_13031;
    wire new_Jinkela_wire_11842;
    wire new_Jinkela_wire_20336;
    wire new_Jinkela_wire_7315;
    wire new_Jinkela_wire_19000;
    wire new_Jinkela_wire_21154;
    wire new_Jinkela_wire_19457;
    wire _0054_;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_2244;
    wire new_Jinkela_wire_19969;
    wire new_Jinkela_wire_16690;
    wire new_Jinkela_wire_16186;
    wire new_Jinkela_wire_20927;
    wire new_Jinkela_wire_6261;
    wire new_Jinkela_wire_19885;
    wire _1371_;
    wire new_Jinkela_wire_14197;
    wire new_Jinkela_wire_3024;
    wire new_Jinkela_wire_12632;
    wire new_Jinkela_wire_2524;
    wire new_Jinkela_wire_5032;
    wire new_Jinkela_wire_20581;
    wire new_Jinkela_wire_11003;
    wire new_Jinkela_wire_8927;
    wire new_Jinkela_wire_6104;
    wire new_Jinkela_wire_16408;
    wire new_Jinkela_wire_20813;
    wire new_Jinkela_wire_11999;
    wire new_Jinkela_wire_10792;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_13123;
    wire new_Jinkela_wire_19196;
    wire new_Jinkela_wire_14553;
    wire new_Jinkela_wire_1715;
    wire new_Jinkela_wire_4720;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_16229;
    wire new_Jinkela_wire_18400;
    wire new_Jinkela_wire_19891;
    wire new_Jinkela_wire_14259;
    wire new_Jinkela_wire_18387;
    wire new_Jinkela_wire_18398;
    wire _1693_;
    wire new_Jinkela_wire_21231;
    wire new_Jinkela_wire_8583;
    wire new_Jinkela_wire_5759;
    wire new_Jinkela_wire_17467;
    wire new_Jinkela_wire_20295;
    wire new_Jinkela_wire_7676;
    wire new_Jinkela_wire_9874;
    wire new_Jinkela_wire_2422;
    wire new_Jinkela_wire_7033;
    wire new_Jinkela_wire_20216;
    wire new_Jinkela_wire_16081;
    wire new_Jinkela_wire_8240;
    wire new_Jinkela_wire_10067;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_14432;
    wire new_Jinkela_wire_18142;
    wire new_Jinkela_wire_16336;
    wire new_Jinkela_wire_1943;
    wire new_Jinkela_wire_5390;
    wire new_Jinkela_wire_8355;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_4320;
    wire new_Jinkela_wire_16356;
    wire new_Jinkela_wire_12228;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_19252;
    wire new_Jinkela_wire_16512;
    wire new_Jinkela_wire_17992;
    wire new_Jinkela_wire_6484;
    wire new_Jinkela_wire_2203;
    wire new_Jinkela_wire_10314;
    wire new_Jinkela_wire_17117;
    wire new_Jinkela_wire_19219;
    wire _1251_;
    wire new_Jinkela_wire_13695;
    wire new_Jinkela_wire_17497;
    wire new_Jinkela_wire_18323;
    wire new_Jinkela_wire_18197;
    wire new_Jinkela_wire_11247;
    wire new_Jinkela_wire_10277;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_12188;
    wire new_Jinkela_wire_2721;
    wire new_Jinkela_wire_10795;
    wire new_Jinkela_wire_5062;
    wire new_Jinkela_wire_19071;
    wire new_Jinkela_wire_4066;
    wire new_Jinkela_wire_3198;
    wire new_Jinkela_wire_15268;
    wire new_Jinkela_wire_4893;
    wire new_Jinkela_wire_17941;
    wire _1638_;
    wire new_Jinkela_wire_12080;
    wire new_Jinkela_wire_13600;
    wire new_Jinkela_wire_12170;
    wire new_Jinkela_wire_16640;
    wire new_Jinkela_wire_20215;
    wire new_Jinkela_wire_14344;
    wire new_Jinkela_wire_8237;
    wire new_Jinkela_wire_14922;
    wire new_Jinkela_wire_20050;
    wire new_Jinkela_wire_18974;
    wire new_Jinkela_wire_15652;
    wire new_Jinkela_wire_2111;
    wire new_Jinkela_wire_4797;
    wire new_Jinkela_wire_7084;
    wire new_Jinkela_wire_7419;
    wire new_Jinkela_wire_9634;
    wire new_Jinkela_wire_19618;
    wire new_Jinkela_wire_10651;
    wire new_Jinkela_wire_19193;
    wire new_Jinkela_wire_11203;
    wire new_Jinkela_wire_5937;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_5195;
    wire new_Jinkela_wire_8268;
    wire new_Jinkela_wire_16797;
    wire _1493_;
    wire new_Jinkela_wire_11171;
    wire new_Jinkela_wire_19769;
    wire new_Jinkela_wire_18890;
    wire new_Jinkela_wire_12869;
    wire _1218_;
    wire new_Jinkela_wire_10565;
    wire new_Jinkela_wire_17957;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_15758;
    wire new_Jinkela_wire_12635;
    wire new_Jinkela_wire_3688;
    wire _0301_;
    wire new_Jinkela_wire_20039;
    wire new_Jinkela_wire_20324;
    wire new_Jinkela_wire_18880;
    wire new_Jinkela_wire_2362;
    wire _0053_;
    wire new_Jinkela_wire_2050;
    wire new_Jinkela_wire_3497;
    wire _1800_;
    wire new_Jinkela_wire_14790;
    wire new_Jinkela_wire_13348;
    wire new_Jinkela_wire_12004;
    wire new_Jinkela_wire_17333;
    wire new_Jinkela_wire_7404;
    wire new_Jinkela_wire_19246;
    wire new_Jinkela_wire_17132;
    wire new_Jinkela_wire_5459;
    wire _0572_;
    wire new_Jinkela_wire_1672;
    wire new_Jinkela_wire_10853;
    wire _0941_;
    wire _1266_;
    wire new_Jinkela_wire_10031;
    wire new_Jinkela_wire_3718;
    wire new_Jinkela_wire_16327;
    wire _1155_;
    wire new_Jinkela_wire_20275;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_16678;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_8651;
    wire _0311_;
    wire new_Jinkela_wire_17360;
    wire new_Jinkela_wire_16540;
    wire _0434_;
    wire new_Jinkela_wire_153;
    wire _1158_;
    wire new_Jinkela_wire_7690;
    wire _1366_;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_4699;
    wire new_Jinkela_wire_9245;
    wire new_Jinkela_wire_12810;
    wire new_Jinkela_wire_2330;
    wire new_Jinkela_wire_11293;
    wire new_Jinkela_wire_7214;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_19800;
    wire new_Jinkela_wire_12996;
    wire _1197_;
    wire new_Jinkela_wire_15560;
    wire new_Jinkela_wire_4979;
    wire new_Jinkela_wire_3770;
    wire new_Jinkela_wire_11494;
    wire new_Jinkela_wire_6623;
    wire new_Jinkela_wire_6506;
    wire new_Jinkela_wire_13507;
    wire new_Jinkela_wire_9463;
    wire new_Jinkela_wire_8891;
    wire new_Jinkela_wire_5414;
    wire new_Jinkela_wire_9063;
    wire _0059_;
    wire new_Jinkela_wire_15255;
    wire new_Jinkela_wire_13414;
    wire _1559_;
    wire _1031_;
    wire new_Jinkela_wire_15106;
    wire new_Jinkela_wire_20315;
    wire new_Jinkela_wire_12669;
    wire new_Jinkela_wire_13559;
    wire new_Jinkela_wire_17720;
    wire new_Jinkela_wire_7829;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_11446;
    wire new_Jinkela_wire_3703;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_9745;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_2425;
    wire new_Jinkela_wire_14291;
    wire new_Jinkela_wire_5157;
    wire new_Jinkela_wire_16611;
    wire new_Jinkela_wire_15421;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_2270;
    wire _0488_;
    wire new_Jinkela_wire_5620;
    wire new_Jinkela_wire_17223;
    wire new_Jinkela_wire_15129;
    wire new_Jinkela_wire_14547;
    wire new_Jinkela_wire_18768;
    wire new_Jinkela_wire_9750;
    wire new_Jinkela_wire_10088;
    wire new_Jinkela_wire_18852;
    wire new_Jinkela_wire_7475;
    wire new_Jinkela_wire_19012;
    wire new_Jinkela_wire_5037;
    wire new_Jinkela_wire_476;
    wire _0560_;
    wire new_Jinkela_wire_18518;
    wire new_Jinkela_wire_21093;
    wire new_Jinkela_wire_1140;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_18479;
    wire new_Jinkela_wire_15229;
    wire new_Jinkela_wire_4841;
    wire new_Jinkela_wire_7833;
    wire new_Jinkela_wire_20452;
    wire new_Jinkela_wire_19587;
    wire _0028_;
    wire new_Jinkela_wire_15023;
    wire new_Jinkela_wire_9169;
    wire new_Jinkela_wire_7480;
    wire new_Jinkela_wire_18605;
    wire new_Jinkela_wire_6259;
    wire new_Jinkela_wire_8830;
    wire new_Jinkela_wire_3110;
    wire new_Jinkela_wire_14220;
    wire _1152_;
    wire new_Jinkela_wire_19637;
    wire new_Jinkela_wire_12539;
    wire new_Jinkela_wire_5785;
    wire new_Jinkela_wire_9224;
    wire new_Jinkela_wire_7423;
    wire _1608_;
    wire new_Jinkela_wire_5245;
    wire new_Jinkela_wire_12765;
    wire new_Jinkela_wire_9744;
    wire new_Jinkela_wire_10813;
    wire new_Jinkela_wire_11343;
    wire new_Jinkela_wire_7152;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_13767;
    wire new_Jinkela_wire_8104;
    wire new_Jinkela_wire_19653;
    wire new_Jinkela_wire_9493;
    wire new_Jinkela_wire_12544;
    wire new_Jinkela_wire_17781;
    wire new_Jinkela_wire_17246;
    wire new_Jinkela_wire_8867;
    wire new_Jinkela_wire_9735;
    wire new_Jinkela_wire_14841;
    wire new_Jinkela_wire_17489;
    wire new_Jinkela_wire_8091;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_3564;
    wire new_Jinkela_wire_2842;
    wire new_Jinkela_wire_13114;
    wire new_Jinkela_wire_9429;
    wire new_Jinkela_wire_10047;
    wire new_Jinkela_wire_18877;
    wire new_Jinkela_wire_13418;
    wire _0701_;
    wire new_Jinkela_wire_13775;
    wire new_Jinkela_wire_5440;
    wire new_Jinkela_wire_11746;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_10013;
    wire new_Jinkela_wire_8031;
    wire new_Jinkela_wire_11554;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_15806;
    wire new_Jinkela_wire_1284;
    wire new_Jinkela_wire_10198;
    wire new_Jinkela_wire_20021;
    wire new_Jinkela_wire_20975;
    wire new_Jinkela_wire_18977;
    wire new_Jinkela_wire_13745;
    wire new_Jinkela_wire_18207;
    wire new_Jinkela_wire_20823;
    wire new_Jinkela_wire_14898;
    wire new_Jinkela_wire_7843;
    wire new_Jinkela_wire_11646;
    wire new_Jinkela_wire_19354;
    wire new_Jinkela_wire_7650;
    wire new_Jinkela_wire_2720;
    wire new_Jinkela_wire_16453;
    wire new_Jinkela_wire_5944;
    wire new_Jinkela_wire_3136;
    wire new_Jinkela_wire_8846;
    wire new_Jinkela_wire_20726;
    wire new_Jinkela_wire_12072;
    wire new_Jinkela_wire_21095;
    wire new_Jinkela_wire_2945;
    wire new_Jinkela_wire_16483;
    wire _0906_;
    wire new_Jinkela_wire_13537;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_16199;
    wire new_Jinkela_wire_11789;
    wire new_Jinkela_wire_17503;
    wire new_Jinkela_wire_7435;
    wire new_Jinkela_wire_7338;
    wire new_Jinkela_wire_3982;
    wire new_Jinkela_wire_315;
    wire _0741_;
    wire new_Jinkela_wire_13029;
    wire new_Jinkela_wire_9839;
    wire new_Jinkela_wire_14787;
    wire _1050_;
    wire new_Jinkela_wire_5119;
    wire new_Jinkela_wire_6916;
    wire new_Jinkela_wire_9993;
    wire new_Jinkela_wire_9019;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_11224;
    wire new_Jinkela_wire_13868;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_11410;
    wire new_Jinkela_wire_7278;
    wire new_Jinkela_wire_5338;
    wire new_Jinkela_wire_12793;
    wire new_Jinkela_wire_18765;
    wire new_Jinkela_wire_12121;
    wire new_Jinkela_wire_14864;
    wire new_Jinkela_wire_12828;
    wire new_Jinkela_wire_15939;
    wire new_Jinkela_wire_9849;
    wire new_Jinkela_wire_11782;
    wire new_Jinkela_wire_10647;
    wire new_Jinkela_wire_17732;
    wire new_Jinkela_wire_17549;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_11380;
    wire new_Jinkela_wire_2949;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_13528;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_20345;
    wire new_Jinkela_wire_6748;
    wire new_Jinkela_wire_5213;
    wire new_Jinkela_wire_15540;
    wire new_Jinkela_wire_15480;
    wire new_Jinkela_wire_18637;
    wire new_Jinkela_wire_14984;
    wire _0344_;
    wire new_Jinkela_wire_2529;
    wire new_Jinkela_wire_9124;
    wire new_Jinkela_wire_14542;
    wire new_Jinkela_wire_10438;
    wire new_Jinkela_wire_1712;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_13667;
    wire new_Jinkela_wire_2735;
    wire new_Jinkela_wire_3751;
    wire new_Jinkela_wire_5835;
    wire new_Jinkela_wire_13822;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_8286;
    wire new_Jinkela_wire_21249;
    wire new_Jinkela_wire_10488;
    wire _0601_;
    wire new_Jinkela_wire_2729;
    wire new_Jinkela_wire_9935;
    wire new_Jinkela_wire_5880;
    wire new_Jinkela_wire_12598;
    wire new_Jinkela_wire_18471;
    wire new_Jinkela_wire_13723;
    wire new_Jinkela_wire_17307;
    wire new_Jinkela_wire_10434;
    wire _0719_;
    wire new_Jinkela_wire_14288;
    wire new_Jinkela_wire_8895;
    wire new_Jinkela_wire_20534;
    wire new_Jinkela_wire_15192;
    wire new_Jinkela_wire_3478;
    wire new_Jinkela_wire_13777;
    wire new_Jinkela_wire_21046;
    wire new_Jinkela_wire_8700;
    wire new_Jinkela_wire_7556;
    wire new_Jinkela_wire_6481;
    wire new_Jinkela_wire_19445;
    wire new_Jinkela_wire_8568;
    wire new_Jinkela_wire_11994;
    wire _0483_;
    wire new_Jinkela_wire_11819;
    wire new_Jinkela_wire_3527;
    wire new_Jinkela_wire_11093;
    wire new_Jinkela_wire_5702;
    wire new_Jinkela_wire_8761;
    wire _0313_;
    wire new_Jinkela_wire_4685;
    wire new_Jinkela_wire_15678;
    wire _0732_;
    wire new_Jinkela_wire_11210;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_8731;
    wire new_Jinkela_wire_20427;
    wire new_Jinkela_wire_11814;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_18841;
    wire new_Jinkela_wire_17545;
    wire new_Jinkela_wire_18021;
    wire new_Jinkela_wire_4865;
    wire new_Jinkela_wire_8047;
    wire _1101_;
    wire new_Jinkela_wire_2525;
    wire new_Jinkela_wire_20103;
    wire new_Jinkela_wire_8976;
    wire new_Jinkela_wire_20347;
    wire new_Jinkela_wire_11707;
    wire new_Jinkela_wire_6691;
    wire new_Jinkela_wire_7984;
    wire new_Jinkela_wire_1804;
    wire _1116_;
    wire new_Jinkela_wire_8032;
    wire _1117_;
    wire new_Jinkela_wire_4262;
    wire new_Jinkela_wire_20781;
    wire new_Jinkela_wire_9287;
    wire new_Jinkela_wire_14106;
    wire new_Jinkela_wire_19696;
    wire new_Jinkela_wire_11365;
    wire new_Jinkela_wire_13683;
    wire new_Jinkela_wire_8866;
    wire _1119_;
    wire new_Jinkela_wire_15065;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_4306;
    wire new_Jinkela_wire_14103;
    wire new_Jinkela_wire_15693;
    wire new_Jinkela_wire_6967;
    wire new_Jinkela_wire_15264;
    wire _0938_;
    wire new_Jinkela_wire_12962;
    wire new_Jinkela_wire_3303;
    wire new_Jinkela_wire_9227;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_14890;
    wire _1577_;
    wire new_Jinkela_wire_4016;
    wire new_Jinkela_wire_11398;
    wire new_Jinkela_wire_18172;
    wire new_Jinkela_wire_18630;
    wire new_Jinkela_wire_8675;
    wire new_Jinkela_wire_15579;
    wire new_Jinkela_wire_6789;
    wire new_Jinkela_wire_13618;
    wire new_Jinkela_wire_5413;
    wire new_Jinkela_wire_8785;
    wire _0946_;
    wire new_Jinkela_wire_4064;
    wire new_Jinkela_wire_11698;
    wire new_Jinkela_wire_9873;
    wire new_Jinkela_wire_9466;
    wire new_Jinkela_wire_4205;
    wire new_Jinkela_wire_11433;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_15205;
    wire new_Jinkela_wire_15154;
    wire _0710_;
    wire new_Jinkela_wire_11700;
    wire new_Jinkela_wire_20595;
    wire new_Jinkela_wire_5992;
    wire new_Jinkela_wire_13502;
    wire new_Jinkela_wire_13080;
    wire new_Jinkela_wire_14753;
    wire new_Jinkela_wire_11268;
    wire new_Jinkela_wire_10562;
    wire new_Jinkela_wire_6501;
    wire new_Jinkela_wire_4439;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_4529;
    wire _1780_;
    wire new_Jinkela_wire_2854;
    wire new_Jinkela_wire_9142;
    wire new_Jinkela_wire_14211;
    wire new_Jinkela_wire_5451;
    wire new_Jinkela_wire_4904;
    wire new_Jinkela_wire_9777;
    wire new_Jinkela_wire_19626;
    wire new_Jinkela_wire_5406;
    wire new_Jinkela_wire_15125;
    wire new_Jinkela_wire_17738;
    wire new_Jinkela_wire_6091;
    wire new_Jinkela_wire_16088;
    wire new_Jinkela_wire_11786;
    wire new_Jinkela_wire_4983;
    wire new_Jinkela_wire_19367;
    wire new_Jinkela_wire_13223;
    wire new_Jinkela_wire_15634;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_9831;
    wire new_Jinkela_wire_11415;
    wire new_Jinkela_wire_19672;
    wire _0063_;
    wire new_Jinkela_wire_1960;
    wire new_Jinkela_wire_5849;
    wire new_Jinkela_wire_7078;
    wire new_Jinkela_wire_10405;
    wire new_Jinkela_wire_14377;
    wire _1339_;
    wire new_Jinkela_wire_11834;
    wire new_Jinkela_wire_7072;
    wire new_Jinkela_wire_18983;
    wire new_Jinkela_wire_8737;
    wire new_Jinkela_wire_20311;
    wire new_Jinkela_wire_160;
    wire _0264_;
    wire new_Jinkela_wire_1560;
    wire _1320_;
    wire new_Jinkela_wire_10499;
    wire new_Jinkela_wire_4624;
    wire new_Jinkela_wire_9920;
    wire new_Jinkela_wire_16249;
    wire new_Jinkela_wire_18985;
    wire new_Jinkela_wire_18618;
    wire new_Jinkela_wire_2757;
    wire new_Jinkela_wire_3402;
    wire new_Jinkela_wire_2123;
    wire new_Jinkela_wire_9183;
    wire new_Jinkela_wire_12104;
    wire new_Jinkela_wire_3700;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_3857;
    wire new_Jinkela_wire_20394;
    wire _0405_;
    wire new_Jinkela_wire_8778;
    wire new_Jinkela_wire_930;
    wire new_Jinkela_wire_3455;
    wire new_Jinkela_wire_8688;
    wire new_Jinkela_wire_3899;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_12784;
    wire new_Jinkela_wire_7285;
    wire new_Jinkela_wire_14564;
    wire new_Jinkela_wire_2771;
    wire new_Jinkela_wire_16650;
    wire new_Jinkela_wire_7241;
    wire new_Jinkela_wire_18956;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_18275;
    wire new_Jinkela_wire_10925;
    wire new_Jinkela_wire_19036;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_12606;
    wire new_Jinkela_wire_17027;
    wire new_Jinkela_wire_10751;
    wire new_Jinkela_wire_12857;
    wire new_Jinkela_wire_7281;
    wire new_Jinkela_wire_5762;
    wire _1352_;
    wire new_Jinkela_wire_6169;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_2931;
    wire new_Jinkela_wire_14763;
    wire new_Jinkela_wire_12030;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_3038;
    wire new_Jinkela_wire_3652;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_14597;
    wire new_Jinkela_wire_1882;
    wire new_Jinkela_wire_17128;
    wire new_Jinkela_wire_18511;
    wire new_Jinkela_wire_1820;
    wire new_Jinkela_wire_12919;
    wire new_Jinkela_wire_14456;
    wire new_Jinkela_wire_20493;
    wire new_Jinkela_wire_12630;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_4483;
    wire new_Jinkela_wire_4085;
    wire new_Jinkela_wire_19906;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_13987;
    wire new_Jinkela_wire_19266;
    wire new_Jinkela_wire_14340;
    wire new_Jinkela_wire_21094;
    wire new_Jinkela_wire_13307;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_21311;
    wire new_Jinkela_wire_15440;
    wire new_Jinkela_wire_5105;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_6925;
    wire _0229_;
    wire new_Jinkela_wire_14950;
    wire new_Jinkela_wire_15190;
    wire new_Jinkela_wire_2702;
    wire _1708_;
    wire new_Jinkela_wire_9058;
    wire new_Jinkela_wire_5160;
    wire new_Jinkela_wire_18572;
    wire new_Jinkela_wire_2683;
    wire new_Jinkela_wire_18541;
    wire new_Jinkela_wire_15464;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_11804;
    wire new_Jinkela_wire_14035;
    wire new_Jinkela_wire_9481;
    wire new_Jinkela_wire_178;
    wire _0354_;
    wire new_Jinkela_wire_18744;
    wire new_Jinkela_wire_4737;
    wire new_Jinkela_wire_11969;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_4499;
    wire new_Jinkela_wire_4341;
    wire new_Jinkela_wire_19432;
    wire new_Jinkela_wire_6834;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_15118;
    wire new_Jinkela_wire_19920;
    wire _0592_;
    wire new_Jinkela_wire_15943;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_9034;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_8326;
    wire new_Jinkela_wire_17963;
    wire _0547_;
    wire new_Jinkela_wire_17076;
    wire new_Jinkela_wire_4823;
    wire _0691_;
    wire new_Jinkela_wire_14860;
    wire new_Jinkela_wire_5734;
    wire new_Jinkela_wire_12045;
    wire new_Jinkela_wire_542;
    wire _0418_;
    wire _1591_;
    wire new_Jinkela_wire_13284;
    wire new_Jinkela_wire_9826;
    wire new_Jinkela_wire_20453;
    wire new_Jinkela_wire_11563;
    wire new_Jinkela_wire_8748;
    wire new_Jinkela_wire_12780;
    wire new_Jinkela_wire_2905;
    wire new_Jinkela_wire_7337;
    wire new_Jinkela_wire_15679;
    wire new_Jinkela_wire_13521;
    wire new_Jinkela_wire_4187;
    wire new_Jinkela_wire_19610;
    wire new_Jinkela_wire_11181;
    wire new_Jinkela_wire_9519;
    wire new_Jinkela_wire_11966;
    wire new_Jinkela_wire_17152;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_12392;
    wire new_Jinkela_wire_21186;
    wire new_Jinkela_wire_10116;
    wire new_Jinkela_wire_6046;
    wire new_Jinkela_wire_8359;
    wire new_Jinkela_wire_1637;
    wire _1297_;
    wire new_Jinkela_wire_2837;
    wire new_Jinkela_wire_3644;
    wire new_Jinkela_wire_2537;
    wire new_Jinkela_wire_16618;
    wire new_Jinkela_wire_2380;
    wire new_Jinkela_wire_18478;
    wire new_Jinkela_wire_18905;
    wire new_Jinkela_wire_4512;
    wire new_Jinkela_wire_6415;
    wire new_Jinkela_wire_7778;
    wire new_Jinkela_wire_6872;
    wire new_Jinkela_wire_1966;
    wire _0845_;
    wire new_Jinkela_wire_745;
    wire _1230_;
    wire new_Jinkela_wire_15972;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_5024;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_9652;
    wire new_Jinkela_wire_6257;
    wire new_Jinkela_wire_2649;
    wire new_Jinkela_wire_16019;
    wire new_Jinkela_wire_10400;
    wire new_Jinkela_wire_5812;
    wire new_Jinkela_wire_7559;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_10868;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_14989;
    wire new_Jinkela_wire_12937;
    wire new_Jinkela_wire_3278;
    wire new_Jinkela_wire_1282;
    wire _1374_;
    wire new_Jinkela_wire_5741;
    wire new_Jinkela_wire_20779;
    wire new_Jinkela_wire_8884;
    wire new_Jinkela_wire_9020;
    wire new_Jinkela_wire_534;
    wire _0655_;
    wire new_Jinkela_wire_12811;
    wire new_Jinkela_wire_2699;
    wire new_Jinkela_wire_18324;
    wire new_Jinkela_wire_7327;
    wire new_Jinkela_wire_17464;
    wire new_Jinkela_wire_7001;
    wire new_Jinkela_wire_17323;
    wire new_Jinkela_wire_16442;
    wire new_Jinkela_wire_20616;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_12361;
    wire new_Jinkela_wire_10622;
    wire new_Jinkela_wire_3883;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_19853;
    wire new_Jinkela_wire_10935;
    wire new_Jinkela_wire_8461;
    wire new_Jinkela_wire_3300;
    wire new_Jinkela_wire_15557;
    wire new_Jinkela_wire_6440;
    wire new_Jinkela_wire_4744;
    wire _0561_;
    wire _0782_;
    wire new_Jinkela_wire_15628;
    wire new_Jinkela_wire_11253;
    wire new_Jinkela_wire_9180;
    wire new_Jinkela_wire_21187;
    wire new_Jinkela_wire_16153;
    wire new_Jinkela_wire_9907;
    wire new_Jinkela_wire_6647;
    wire new_Jinkela_wire_5528;
    wire new_Jinkela_wire_20430;
    wire new_Jinkela_wire_10818;
    wire new_Jinkela_wire_14514;
    wire new_Jinkela_wire_9898;
    wire new_Jinkela_wire_2192;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_4036;
    wire new_Jinkela_wire_10620;
    wire new_Jinkela_wire_15787;
    wire new_Jinkela_wire_8971;
    wire new_Jinkela_wire_15624;
    wire new_Jinkela_wire_16230;
    wire new_Jinkela_wire_4806;
    wire new_Jinkela_wire_9454;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_19801;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_8509;
    wire new_Jinkela_wire_10121;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_8579;
    wire new_Jinkela_wire_16541;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_8801;
    wire new_Jinkela_wire_15276;
    wire new_Jinkela_wire_6250;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_9520;
    wire new_Jinkela_wire_20411;
    wire new_Jinkela_wire_3994;
    wire new_Jinkela_wire_7839;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_7457;
    wire new_Jinkela_wire_2758;
    wire new_Jinkela_wire_6618;
    wire new_Jinkela_wire_11695;
    wire new_Jinkela_wire_5274;
    wire new_Jinkela_wire_18649;
    wire _0516_;
    wire new_Jinkela_wire_14537;
    wire _1174_;
    wire new_Jinkela_wire_14667;
    wire new_Jinkela_wire_3833;
    wire new_Jinkela_wire_14080;
    wire new_Jinkela_wire_483;
    wire _0689_;
    wire new_Jinkela_wire_10419;
    wire new_Jinkela_wire_16550;
    wire new_Jinkela_wire_3752;
    wire new_Jinkela_wire_8633;
    wire new_Jinkela_wire_19453;
    wire new_Jinkela_wire_10893;
    wire new_Jinkela_wire_6910;
    wire _1412_;
    wire new_Jinkela_wire_11079;
    wire new_Jinkela_wire_15068;
    wire _1679_;
    wire new_Jinkela_wire_6549;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_16354;
    wire new_Jinkela_wire_13856;
    wire new_Jinkela_wire_18438;
    wire new_Jinkela_wire_8226;
    wire new_Jinkela_wire_6788;
    wire new_Jinkela_wire_11836;
    wire new_Jinkela_wire_2764;
    wire new_Jinkela_wire_17788;
    wire new_Jinkela_wire_18311;
    wire new_Jinkela_wire_7035;
    wire new_Jinkela_wire_3865;
    wire new_Jinkela_wire_8283;
    wire _0045_;
    wire new_Jinkela_wire_12220;
    wire new_Jinkela_wire_6405;
    wire new_Jinkela_wire_16322;
    wire new_Jinkela_wire_5457;
    wire new_Jinkela_wire_13807;
    wire new_Jinkela_wire_13809;
    wire new_Jinkela_wire_10345;
    wire new_Jinkela_wire_14810;
    wire new_Jinkela_wire_12746;
    wire new_Jinkela_wire_17848;
    wire new_Jinkela_wire_2436;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_11401;
    wire new_Jinkela_wire_15290;
    wire new_Jinkela_wire_2997;
    wire new_Jinkela_wire_15788;
    wire new_Jinkela_wire_15410;
    wire _0971_;
    wire new_Jinkela_wire_4249;
    wire new_Jinkela_wire_16524;
    wire new_Jinkela_wire_7471;
    wire _0515_;
    wire new_Jinkela_wire_9358;
    wire new_Jinkela_wire_15427;
    wire new_Jinkela_wire_11503;
    wire new_Jinkela_wire_11670;
    wire new_Jinkela_wire_19234;
    wire new_Jinkela_wire_13973;
    wire new_Jinkela_wire_11035;
    wire new_Jinkela_wire_15397;
    wire new_Jinkela_wire_14515;
    wire new_Jinkela_wire_15224;
    wire new_Jinkela_wire_4646;
    wire new_Jinkela_wire_2227;
    wire new_Jinkela_wire_5339;
    wire new_Jinkela_wire_18144;
    wire new_Jinkela_wire_2912;
    wire new_Jinkela_wire_7665;
    wire new_Jinkela_wire_18667;
    wire new_Jinkela_wire_5026;
    wire new_Jinkela_wire_4080;
    wire new_Jinkela_wire_20830;
    wire new_Jinkela_wire_13614;
    wire new_Jinkela_wire_14956;
    wire _0846_;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_1391;
    wire new_Jinkela_wire_16725;
    wire new_Jinkela_wire_19608;
    wire new_Jinkela_wire_10561;
    wire new_Jinkela_wire_7307;
    wire new_Jinkela_wire_17719;
    wire new_Jinkela_wire_17247;
    wire new_Jinkela_wire_7347;
    wire new_Jinkela_wire_7331;
    wire new_Jinkela_wire_17695;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_6232;
    wire new_Jinkela_wire_12736;
    wire new_Jinkela_wire_2229;
    wire new_Jinkela_wire_9614;
    wire new_Jinkela_wire_4589;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_14067;
    wire new_Jinkela_wire_5805;
    wire new_Jinkela_wire_12480;
    wire new_Jinkela_wire_11340;
    wire new_Jinkela_wire_17967;
    wire new_Jinkela_wire_8284;
    wire new_Jinkela_wire_6600;
    wire new_Jinkela_wire_10004;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_20040;
    wire new_net_3922;
    wire new_Jinkela_wire_2770;
    wire new_Jinkela_wire_11886;
    wire new_Jinkela_wire_7043;
    wire new_Jinkela_wire_2617;
    wire new_Jinkela_wire_18896;
    wire new_Jinkela_wire_9384;
    wire _0749_;
    wire new_Jinkela_wire_9976;
    wire new_Jinkela_wire_15279;
    wire _0382_;
    wire new_Jinkela_wire_9097;
    wire _1517_;
    wire new_Jinkela_wire_19692;
    wire new_Jinkela_wire_12792;
    wire new_Jinkela_wire_21041;
    wire new_Jinkela_wire_17742;
    wire new_Jinkela_wire_9246;
    wire new_Jinkela_wire_9896;
    wire new_Jinkela_wire_6493;
    wire new_Jinkela_wire_20333;
    wire new_Jinkela_wire_14380;
    wire _1836_;
    wire new_Jinkela_wire_8105;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_1734;
    wire new_Jinkela_wire_15696;
    wire new_Jinkela_wire_10293;
    wire new_Jinkela_wire_18958;
    wire new_Jinkela_wire_16597;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_21319;
    wire new_Jinkela_wire_5729;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_11594;
    wire new_Jinkela_wire_16426;
    wire new_Jinkela_wire_5997;
    wire new_Jinkela_wire_5700;
    wire _0791_;
    wire new_Jinkela_wire_11961;
    wire new_Jinkela_wire_19094;
    wire new_Jinkela_wire_3933;
    wire _1431_;
    wire new_Jinkela_wire_9897;
    wire new_Jinkela_wire_12693;
    wire new_Jinkela_wire_10931;
    wire new_Jinkela_wire_2328;
    wire new_Jinkela_wire_15055;
    wire new_Jinkela_wire_11795;
    wire new_Jinkela_wire_8175;
    wire _0369_;
    wire new_Jinkela_wire_11044;
    wire new_Jinkela_wire_4438;
    wire _1059_;
    wire new_Jinkela_wire_5949;
    wire new_Jinkela_wire_11466;
    wire new_Jinkela_wire_16340;
    wire new_Jinkela_wire_2205;
    wire new_Jinkela_wire_13172;
    wire new_Jinkela_wire_16908;
    wire new_Jinkela_wire_11579;
    wire new_Jinkela_wire_2675;
    wire new_Jinkela_wire_4329;
    wire new_Jinkela_wire_5588;
    wire new_Jinkela_wire_21327;
    wire new_Jinkela_wire_21102;
    wire new_Jinkela_wire_3734;
    wire new_Jinkela_wire_20134;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_9051;
    wire new_Jinkela_wire_1787;
    wire new_Jinkela_wire_10816;
    wire _0153_;
    wire _1472_;
    wire new_Jinkela_wire_7178;
    wire new_Jinkela_wire_15168;
    wire new_Jinkela_wire_13137;
    wire new_Jinkela_wire_10532;
    wire new_Jinkela_wire_9289;
    wire _1825_;
    wire new_Jinkela_wire_8399;
    wire new_Jinkela_wire_12738;
    wire new_Jinkela_wire_4603;
    wire new_Jinkela_wire_15930;
    wire new_Jinkela_wire_16537;
    wire new_Jinkela_wire_9055;
    wire new_Jinkela_wire_7631;
    wire new_Jinkela_wire_9734;
    wire new_Jinkela_wire_10897;
    wire new_Jinkela_wire_14373;
    wire new_Jinkela_wire_19321;
    wire new_Jinkela_wire_17407;
    wire new_Jinkela_wire_20712;
    wire new_Jinkela_wire_12685;
    wire new_Jinkela_wire_19092;
    wire new_Jinkela_wire_2533;
    wire new_Jinkela_wire_8109;
    wire new_Jinkela_wire_18750;
    wire new_Jinkela_wire_7300;
    wire new_Jinkela_wire_17670;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_6195;
    wire new_Jinkela_wire_10892;
    wire new_Jinkela_wire_3607;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_8267;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_18726;
    wire new_Jinkela_wire_16661;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_14818;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_11637;
    wire new_Jinkela_wire_17191;
    wire new_Jinkela_wire_9357;
    wire new_Jinkela_wire_18360;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_7511;
    wire new_Jinkela_wire_18291;
    wire new_Jinkela_wire_19375;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_2488;
    wire new_Jinkela_wire_19516;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_16143;
    wire new_Jinkela_wire_8000;
    wire new_Jinkela_wire_2212;
    wire new_Jinkela_wire_6444;
    wire new_Jinkela_wire_9122;
    wire new_Jinkela_wire_7481;
    wire new_Jinkela_wire_18587;
    wire new_Jinkela_wire_19674;
    wire new_Jinkela_wire_14990;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_3077;
    wire _1837_;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_3992;
    wire new_Jinkela_wire_8080;
    wire new_Jinkela_wire_1848;
    wire new_Jinkela_wire_20391;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_16149;
    wire new_Jinkela_wire_21006;
    wire new_Jinkela_wire_15078;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_12103;
    wire new_Jinkela_wire_1647;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_16801;
    wire new_Jinkela_wire_14997;
    wire new_Jinkela_wire_7592;
    wire new_Jinkela_wire_5686;
    wire new_Jinkela_wire_3977;
    wire new_Jinkela_wire_15436;
    wire new_Jinkela_wire_14705;
    wire new_Jinkela_wire_19228;
    wire new_Jinkela_wire_17359;
    wire new_Jinkela_wire_6886;
    wire new_Jinkela_wire_12647;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_14171;
    wire new_Jinkela_wire_20497;
    wire new_Jinkela_wire_17531;
    wire new_Jinkela_wire_20790;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_4115;
    wire new_Jinkela_wire_9150;
    wire _1151_;
    wire _1483_;
    wire new_Jinkela_wire_5602;
    wire new_Jinkela_wire_7303;
    wire new_Jinkela_wire_3597;
    wire new_Jinkela_wire_17056;
    wire new_Jinkela_wire_9427;
    wire new_Jinkela_wire_21211;
    wire new_Jinkela_wire_6118;
    wire new_Jinkela_wire_15974;
    wire new_Jinkela_wire_4871;
    wire new_Jinkela_wire_13108;
    wire new_Jinkela_wire_3342;
    wire new_Jinkela_wire_20499;
    wire new_Jinkela_wire_11492;
    wire new_Jinkela_wire_6460;
    wire new_Jinkela_wire_9675;
    wire new_Jinkela_wire_1720;
    wire new_Jinkela_wire_7047;
    wire new_Jinkela_wire_79;
    wire new_Jinkela_wire_4338;
    wire new_Jinkela_wire_15194;
    wire new_Jinkela_wire_9600;
    wire new_Jinkela_wire_2824;
    wire _1828_;
    wire new_Jinkela_wire_16412;
    wire new_Jinkela_wire_13214;
    wire new_Jinkela_wire_7818;
    wire new_Jinkela_wire_6728;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_5035;
    wire new_Jinkela_wire_5814;
    wire new_Jinkela_wire_5316;
    wire _1106_;
    wire new_Jinkela_wire_17558;
    wire new_Jinkela_wire_20836;
    wire new_Jinkela_wire_6881;
    wire new_Jinkela_wire_10940;
    wire new_Jinkela_wire_13643;
    wire new_Jinkela_wire_6197;
    wire new_Jinkela_wire_19355;
    wire new_Jinkela_wire_7417;
    wire new_Jinkela_wire_15340;
    wire new_Jinkela_wire_4738;
    wire new_Jinkela_wire_2928;
    wire new_Jinkela_wire_11939;
    wire new_Jinkela_wire_10281;
    wire new_Jinkela_wire_5112;
    wire new_Jinkela_wire_8968;
    wire new_Jinkela_wire_20771;
    wire new_Jinkela_wire_16396;
    wire new_Jinkela_wire_13852;
    wire new_Jinkela_wire_8813;
    wire new_Jinkela_wire_6587;
    wire new_Jinkela_wire_15456;
    wire new_Jinkela_wire_6575;
    wire new_Jinkela_wire_18234;
    wire new_Jinkela_wire_2624;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_14366;
    wire new_Jinkela_wire_18514;
    wire new_Jinkela_wire_3392;
    wire new_Jinkela_wire_16609;
    wire _1489_;
    wire new_Jinkela_wire_6142;
    wire new_Jinkela_wire_3344;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_17582;
    wire new_Jinkela_wire_14973;
    wire new_Jinkela_wire_7051;
    wire new_Jinkela_wire_20878;
    wire new_Jinkela_wire_4558;
    wire new_Jinkela_wire_9212;
    wire new_Jinkela_wire_2455;
    wire new_Jinkela_wire_7989;
    wire new_Jinkela_wire_10632;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_15548;
    wire new_Jinkela_wire_14847;
    wire new_Jinkela_wire_7296;
    wire _0587_;
    wire new_Jinkela_wire_11612;
    wire new_Jinkela_wire_9523;
    wire new_Jinkela_wire_19701;
    wire new_Jinkela_wire_11124;
    wire new_Jinkela_wire_4484;
    wire new_Jinkela_wire_3352;
    wire new_Jinkela_wire_18412;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_18292;
    wire new_Jinkela_wire_15643;
    wire new_Jinkela_wire_6978;
    wire new_Jinkela_wire_379;
    wire _1237_;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_18758;
    wire new_Jinkela_wire_3580;
    wire _0862_;
    wire new_Jinkela_wire_20059;
    wire new_Jinkela_wire_10592;
    wire new_Jinkela_wire_1930;
    wire new_Jinkela_wire_9635;
    wire new_Jinkela_wire_5540;
    wire new_Jinkela_wire_1859;
    wire _0956_;
    wire new_Jinkela_wire_12515;
    wire _0429_;
    wire new_Jinkela_wire_7195;
    wire new_Jinkela_wire_19067;
    wire new_Jinkela_wire_17093;
    wire new_Jinkela_wire_14946;
    wire new_Jinkela_wire_10976;
    wire new_Jinkela_wire_13415;
    wire new_Jinkela_wire_21024;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_2085;
    wire new_Jinkela_wire_4772;
    wire new_Jinkela_wire_11650;
    wire new_Jinkela_wire_12110;
    wire new_Jinkela_wire_20352;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_20088;
    wire _0600_;
    wire new_Jinkela_wire_5542;
    wire _0349_;
    wire new_Jinkela_wire_17105;
    wire new_Jinkela_wire_18107;
    wire new_Jinkela_wire_18772;
    wire new_Jinkela_wire_6330;
    wire new_Jinkela_wire_2450;
    wire new_Jinkela_wire_16926;
    wire new_Jinkela_wire_5889;
    wire new_Jinkela_wire_1973;
    wire new_Jinkela_wire_19680;
    wire new_Jinkela_wire_20162;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_13686;
    wire new_Jinkela_wire_15383;
    wire new_Jinkela_wire_8377;
    wire new_Jinkela_wire_1197;
    wire _0499_;
    wire new_Jinkela_wire_18208;
    wire new_Jinkela_wire_19638;
    wire new_Jinkela_wire_11564;
    wire new_Jinkela_wire_16237;
    wire new_Jinkela_wire_17432;
    wire new_Jinkela_wire_3995;
    wire new_Jinkela_wire_19574;
    wire new_Jinkela_wire_15925;
    wire new_Jinkela_wire_2921;
    wire new_Jinkela_wire_2187;
    wire new_Jinkela_wire_17003;
    wire new_Jinkela_wire_21054;
    wire new_Jinkela_wire_6973;
    wire new_Jinkela_wire_9328;
    wire new_Jinkela_wire_3668;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_20692;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_16174;
    wire new_Jinkela_wire_11322;
    wire new_Jinkela_wire_9846;
    wire new_Jinkela_wire_2805;
    wire new_Jinkela_wire_11175;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_1091;
    wire _1822_;
    wire _0831_;
    wire new_Jinkela_wire_14706;
    wire new_Jinkela_wire_15546;
    wire new_Jinkela_wire_6603;
    wire new_Jinkela_wire_11411;
    wire new_Jinkela_wire_19926;
    wire _1612_;
    wire new_Jinkela_wire_5612;
    wire new_Jinkela_wire_7680;
    wire new_Jinkela_wire_14422;
    wire new_Jinkela_wire_12788;
    wire new_Jinkela_wire_10294;
    wire new_Jinkela_wire_13546;
    wire new_Jinkela_wire_11864;
    wire new_Jinkela_wire_5809;
    wire new_Jinkela_wire_8059;
    wire new_Jinkela_wire_9538;
    wire new_Jinkela_wire_9637;
    wire new_Jinkela_wire_3666;
    wire new_Jinkela_wire_12674;
    wire _0933_;
    wire new_Jinkela_wire_4949;
    wire new_Jinkela_wire_2785;
    wire new_Jinkela_wire_19778;
    wire new_Jinkela_wire_12590;
    wire new_Jinkela_wire_11303;
    wire new_Jinkela_wire_10962;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_1917;
    wire new_Jinkela_wire_4845;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_16500;
    wire new_Jinkela_wire_11788;
    wire new_Jinkela_wire_11225;
    wire new_Jinkela_wire_3740;
    wire _1635_;
    wire new_Jinkela_wire_16415;
    wire new_Jinkela_wire_10631;
    wire new_Jinkela_wire_5007;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_1761;
    wire new_Jinkela_wire_181;
    wire _1716_;
    wire new_Jinkela_wire_8789;
    wire new_Jinkela_wire_6143;
    wire new_Jinkela_wire_6343;
    wire new_Jinkela_wire_7271;
    wire new_Jinkela_wire_17761;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_4616;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_18546;
    wire _1688_;
    wire new_Jinkela_wire_1744;
    wire new_Jinkela_wire_10578;
    wire new_Jinkela_wire_10741;
    wire _0649_;
    wire new_Jinkela_wire_20244;
    wire new_Jinkela_wire_14781;
    wire new_Jinkela_wire_7963;
    wire new_Jinkela_wire_17215;
    wire new_Jinkela_wire_18006;
    wire new_Jinkela_wire_2985;
    wire new_Jinkela_wire_20404;
    wire new_Jinkela_wire_10213;
    wire new_Jinkela_wire_16970;
    wire _0220_;
    wire new_Jinkela_wire_18299;
    wire new_Jinkela_wire_13768;
    wire new_Jinkela_wire_3693;
    wire new_Jinkela_wire_6438;
    wire new_Jinkela_wire_21031;
    wire new_Jinkela_wire_16181;
    wire new_Jinkela_wire_3875;
    wire new_Jinkela_wire_7028;
    wire new_Jinkela_wire_17598;
    wire new_Jinkela_wire_9943;
    wire new_Jinkela_wire_14640;
    wire new_Jinkela_wire_7896;
    wire new_Jinkela_wire_3199;
    wire new_Jinkela_wire_18353;
    wire new_Jinkela_wire_9035;
    wire new_Jinkela_wire_17281;
    wire _1332_;
    wire new_Jinkela_wire_2668;
    wire new_Jinkela_wire_7261;
    wire new_Jinkela_wire_2862;
    wire new_Jinkela_wire_14004;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_6372;
    wire new_Jinkela_wire_10060;
    wire new_Jinkela_wire_17509;
    wire new_Jinkela_wire_7906;
    wire new_Jinkela_wire_11090;
    wire new_Jinkela_wire_14250;
    wire new_Jinkela_wire_13933;
    wire new_Jinkela_wire_16996;
    wire new_Jinkela_wire_16542;
    wire new_Jinkela_wire_11562;
    wire new_Jinkela_wire_20588;
    wire new_Jinkela_wire_14440;
    wire new_Jinkela_wire_14524;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_10904;
    wire new_Jinkela_wire_16696;
    wire _1534_;
    wire new_Jinkela_wire_6609;
    wire new_Jinkela_wire_16195;
    wire new_Jinkela_wire_9145;
    wire new_Jinkela_wire_11722;
    wire new_Jinkela_wire_9133;
    wire new_Jinkela_wire_2886;
    wire new_Jinkela_wire_2245;
    wire _1590_;
    wire new_Jinkela_wire_14941;
    wire new_Jinkela_wire_19972;
    wire _0119_;
    wire new_Jinkela_wire_9186;
    wire new_Jinkela_wire_18921;
    wire new_Jinkela_wire_10139;
    wire new_Jinkela_wire_4909;
    wire new_Jinkela_wire_2732;
    wire new_Jinkela_wire_18074;
    wire new_Jinkela_wire_15030;
    wire _1685_;
    wire new_Jinkela_wire_15682;
    wire new_Jinkela_wire_1921;
    wire new_Jinkela_wire_20976;
    wire new_Jinkela_wire_11835;
    wire new_Jinkela_wire_8925;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_6036;
    wire new_Jinkela_wire_8087;
    wire _0629_;
    wire new_Jinkela_wire_5275;
    wire new_Jinkela_wire_8141;
    wire new_Jinkela_wire_1713;
    wire new_Jinkela_wire_7013;
    wire new_Jinkela_wire_18631;
    wire new_Jinkela_wire_3884;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_17813;
    wire new_Jinkela_wire_9509;
    wire new_Jinkela_wire_6615;
    wire new_Jinkela_wire_15050;
    wire new_Jinkela_wire_14854;
    wire new_Jinkela_wire_19034;
    wire new_Jinkela_wire_17600;
    wire new_Jinkela_wire_10612;
    wire new_Jinkela_wire_10862;
    wire new_Jinkela_wire_18529;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_16402;
    wire new_Jinkela_wire_2500;
    wire new_Jinkela_wire_7458;
    wire new_Jinkela_wire_15789;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_8371;
    wire new_Jinkela_wire_7759;
    wire _1816_;
    wire new_Jinkela_wire_12439;
    wire new_Jinkela_wire_12842;
    wire new_Jinkela_wire_17046;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_14350;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_11495;
    wire new_Jinkela_wire_2377;
    wire new_Jinkela_wire_18927;
    wire new_Jinkela_wire_14261;
    wire new_Jinkela_wire_10916;
    wire new_Jinkela_wire_11419;
    wire new_Jinkela_wire_16493;
    wire new_Jinkela_wire_20408;
    wire new_Jinkela_wire_1888;
    wire _0174_;
    wire new_Jinkela_wire_11483;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_5680;
    wire new_Jinkela_wire_19967;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_7731;
    wire new_Jinkela_wire_9319;
    wire new_Jinkela_wire_15064;
    wire new_Jinkela_wire_17448;
    wire new_Jinkela_wire_15316;
    wire new_Jinkela_wire_18053;
    wire new_Jinkela_wire_16478;
    wire new_Jinkela_wire_4846;
    wire new_Jinkela_wire_3520;
    wire new_Jinkela_wire_10477;
    wire new_Jinkela_wire_86;
    wire new_Jinkela_wire_11017;
    wire new_Jinkela_wire_13569;
    wire new_Jinkela_wire_12124;
    wire new_Jinkela_wire_6287;
    wire new_Jinkela_wire_15325;
    wire new_Jinkela_wire_7094;
    wire new_Jinkela_wire_17907;
    wire new_Jinkela_wire_20722;
    wire new_Jinkela_wire_14948;
    wire new_Jinkela_wire_12983;
    wire new_Jinkela_wire_20090;
    wire new_Jinkela_wire_16770;
    wire new_Jinkela_wire_14448;
    wire new_Jinkela_wire_15821;
    wire new_Jinkela_wire_16458;
    wire _0924_;
    wire new_Jinkela_wire_14959;
    wire new_Jinkela_wire_4608;
    wire new_Jinkela_wire_17146;
    wire new_Jinkela_wire_4926;
    wire new_Jinkela_wire_21209;
    wire new_Jinkela_wire_3261;
    wire new_Jinkela_wire_4727;
    wire new_Jinkela_wire_11518;
    wire new_Jinkela_wire_13500;
    wire new_Jinkela_wire_2523;
    wire _0231_;
    wire new_Jinkela_wire_3962;
    wire new_Jinkela_wire_6998;
    wire new_Jinkela_wire_18092;
    wire new_Jinkela_wire_19968;
    wire new_Jinkela_wire_14374;
    wire new_Jinkela_wire_13193;
    wire new_Jinkela_wire_2242;
    wire new_Jinkela_wire_4855;
    wire new_Jinkela_wire_4163;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_13361;
    wire _1810_;
    wire new_Jinkela_wire_13117;
    wire new_Jinkela_wire_19713;
    wire _0386_;
    wire new_Jinkela_wire_6200;
    wire new_Jinkela_wire_12721;
    wire new_Jinkela_wire_7704;
    wire new_Jinkela_wire_10610;
    wire new_Jinkela_wire_7222;
    wire new_Jinkela_wire_9041;
    wire new_Jinkela_wire_21224;
    wire new_Jinkela_wire_20508;
    wire new_Jinkela_wire_17609;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_9539;
    wire new_Jinkela_wire_14119;
    wire new_Jinkela_wire_10669;
    wire new_Jinkela_wire_20041;
    wire new_Jinkela_wire_10618;
    wire new_Jinkela_wire_4211;
    wire new_Jinkela_wire_13491;
    wire new_Jinkela_wire_15724;
    wire new_Jinkela_wire_17306;
    wire new_Jinkela_wire_18259;
    wire new_Jinkela_wire_3773;
    wire new_Jinkela_wire_1953;
    wire new_Jinkela_wire_20409;
    wire new_Jinkela_wire_5587;
    wire _0530_;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_15385;
    wire new_Jinkela_wire_6555;
    wire new_Jinkela_wire_20156;
    wire _0725_;
    wire new_Jinkela_wire_11699;
    wire new_Jinkela_wire_9595;
    wire new_Jinkela_wire_3461;
    wire new_Jinkela_wire_4043;
    wire new_Jinkela_wire_17810;
    wire new_Jinkela_wire_15752;
    wire _0661_;
    wire new_Jinkela_wire_15879;
    wire new_Jinkela_wire_17424;
    wire new_Jinkela_wire_11712;
    wire new_Jinkela_wire_14658;
    wire new_Jinkela_wire_14796;
    wire new_Jinkela_wire_18430;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_8776;
    wire new_Jinkela_wire_14484;
    wire new_Jinkela_wire_6424;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_16438;
    wire new_Jinkela_wire_11620;
    wire new_Jinkela_wire_7350;
    wire new_Jinkela_wire_12461;
    wire new_Jinkela_wire_6378;
    wire new_Jinkela_wire_18491;
    wire new_Jinkela_wire_9558;
    wire new_Jinkela_wire_2136;
    wire new_Jinkela_wire_11644;
    wire new_Jinkela_wire_2457;
    wire new_Jinkela_wire_14104;
    wire new_Jinkela_wire_21075;
    wire new_Jinkela_wire_8744;
    wire new_Jinkela_wire_20472;
    wire new_Jinkela_wire_9207;
    wire new_Jinkela_wire_7046;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_11981;
    wire new_Jinkela_wire_13149;
    wire new_Jinkela_wire_6577;
    wire _0784_;
    wire new_Jinkela_wire_15779;
    wire new_Jinkela_wire_11339;
    wire new_Jinkela_wire_17358;
    wire new_Jinkela_wire_9480;
    wire new_Jinkela_wire_21329;
    wire new_Jinkela_wire_2487;
    wire new_Jinkela_wire_13043;
    wire new_Jinkela_wire_14632;
    wire new_Jinkela_wire_20605;
    wire new_Jinkela_wire_10261;
    wire new_Jinkela_wire_12337;
    wire new_Jinkela_wire_16221;
    wire new_Jinkela_wire_10313;
    wire new_Jinkela_wire_16118;
    wire new_Jinkela_wire_19159;
    wire new_Jinkela_wire_13126;
    wire new_Jinkela_wire_14568;
    wire new_Jinkela_wire_2749;
    wire new_Jinkela_wire_19722;
    wire new_Jinkela_wire_12946;
    wire new_Jinkela_wire_6181;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_12459;
    wire new_Jinkela_wire_21061;
    wire new_Jinkela_wire_7149;
    wire new_Jinkela_wire_8917;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_18951;
    wire new_Jinkela_wire_5601;
    wire new_Jinkela_wire_13696;
    wire new_Jinkela_wire_20919;
    wire new_Jinkela_wire_15618;
    wire new_Jinkela_wire_17596;
    wire new_Jinkela_wire_8788;
    wire new_Jinkela_wire_4352;
    wire _1722_;
    wire new_Jinkela_wire_15664;
    wire new_Jinkela_wire_19169;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_7354;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_12782;
    wire new_Jinkela_wire_370;
    wire _1219_;
    wire new_Jinkela_wire_11088;
    wire new_Jinkela_wire_10240;
    wire new_Jinkela_wire_2392;
    wire new_Jinkela_wire_17490;
    wire new_Jinkela_wire_14552;
    wire new_Jinkela_wire_18380;
    wire new_Jinkela_wire_2044;
    wire new_Jinkela_wire_15973;
    wire new_Jinkela_wire_16268;
    wire new_Jinkela_wire_13545;
    wire new_Jinkela_wire_3702;
    wire new_Jinkela_wire_10706;
    wire new_Jinkela_wire_7451;
    wire new_Jinkela_wire_6864;
    wire new_Jinkela_wire_11706;
    wire new_Jinkela_wire_2417;
    wire new_Jinkela_wire_7025;
    wire _1275_;
    wire new_Jinkela_wire_17869;
    wire new_Jinkela_wire_12287;
    wire new_Jinkela_wire_15463;
    wire new_Jinkela_wire_12555;
    wire new_Jinkela_wire_7878;
    wire new_Jinkela_wire_17189;
    wire new_Jinkela_wire_16626;
    wire new_Jinkela_wire_4051;
    wire new_Jinkela_wire_20491;
    wire new_Jinkela_wire_10182;
    wire new_Jinkela_wire_4229;
    wire new_Jinkela_wire_16374;
    wire _1514_;
    wire new_Jinkela_wire_20095;
    wire new_Jinkela_wire_18215;
    wire new_Jinkela_wire_19783;
    wire _1647_;
    wire new_Jinkela_wire_9987;
    wire _1026_;
    wire new_Jinkela_wire_2603;
    wire new_Jinkela_wire_2505;
    wire new_Jinkela_wire_14609;
    wire new_Jinkela_wire_3900;
    wire new_Jinkela_wire_17420;
    wire new_Jinkela_wire_12247;
    wire new_Jinkela_wire_7827;
    wire new_Jinkela_wire_15242;
    wire new_Jinkela_wire_8806;
    wire new_Jinkela_wire_13267;
    wire new_Jinkela_wire_11923;
    wire new_Jinkela_wire_20086;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_1444;
    wire _1193_;
    wire new_Jinkela_wire_4109;
    wire new_Jinkela_wire_15923;
    wire new_Jinkela_wire_13271;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_14772;
    wire new_Jinkela_wire_4498;
    wire new_Jinkela_wire_3612;
    wire new_Jinkela_wire_15857;
    wire new_Jinkela_wire_7021;
    wire new_Jinkela_wire_11878;
    wire new_Jinkela_wire_7966;
    wire new_Jinkela_wire_2325;
    wire new_Jinkela_wire_94;
    wire _0306_;
    wire new_Jinkela_wire_12298;
    wire new_Jinkela_wire_2230;
    wire new_Jinkela_wire_5380;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_15490;
    wire new_Jinkela_wire_17930;
    wire new_Jinkela_wire_1475;
    wire new_Jinkela_wire_19363;
    wire new_Jinkela_wire_8025;
    wire new_Jinkela_wire_5673;
    wire new_Jinkela_wire_19113;
    wire new_Jinkela_wire_18564;
    wire new_Jinkela_wire_14010;
    wire new_Jinkela_wire_2851;
    wire new_Jinkela_wire_19739;
    wire new_Jinkela_wire_2844;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_11058;
    wire new_Jinkela_wire_9556;
    wire new_Jinkela_wire_4216;
    wire new_Jinkela_wire_7972;
    wire new_Jinkela_wire_14544;
    wire new_Jinkela_wire_20091;
    wire new_Jinkela_wire_3325;
    wire new_Jinkela_wire_16189;
    wire new_Jinkela_wire_6094;
    wire new_Jinkela_wire_18377;
    wire new_Jinkela_wire_4278;
    wire new_Jinkela_wire_7523;
    wire new_Jinkela_wire_6534;
    wire new_Jinkela_wire_17852;
    wire _0474_;
    wire _0870_;
    wire new_Jinkela_wire_16969;
    wire new_Jinkela_wire_2517;
    wire new_Jinkela_wire_17716;
    wire new_Jinkela_wire_7608;
    wire new_Jinkela_wire_10227;
    wire new_Jinkela_wire_3475;
    wire new_Jinkela_wire_1803;
    wire new_Jinkela_wire_3127;
    wire new_Jinkela_wire_13611;
    wire new_Jinkela_wire_11687;
    wire new_Jinkela_wire_5701;
    wire new_Jinkela_wire_8696;
    wire new_Jinkela_wire_7744;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_5183;
    wire new_Jinkela_wire_14439;
    wire new_Jinkela_wire_6051;
    wire new_Jinkela_wire_12372;
    wire new_Jinkela_wire_5996;
    wire new_Jinkela_wire_2472;
    wire new_Jinkela_wire_19718;
    wire _1715_;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_3408;
    wire new_Jinkela_wire_4212;
    wire new_Jinkela_wire_10366;
    wire new_Jinkela_wire_11332;
    wire new_Jinkela_wire_5709;
    wire new_Jinkela_wire_19312;
    wire new_Jinkela_wire_19836;
    wire new_Jinkela_wire_14961;
    wire new_Jinkela_wire_5028;
    wire new_Jinkela_wire_16557;
    wire new_Jinkela_wire_16113;
    wire new_Jinkela_wire_20592;
    wire new_Jinkela_wire_3701;
    wire new_Jinkela_wire_10364;
    wire _0644_;
    wire _0249_;
    wire new_Jinkela_wire_4378;
    wire _0694_;
    wire new_Jinkela_wire_17541;
    wire new_Jinkela_wire_12673;
    wire new_Jinkela_wire_8802;
    wire new_Jinkela_wire_20469;
    wire new_Jinkela_wire_18245;
    wire new_Jinkela_wire_3862;
    wire new_Jinkela_wire_2924;
    wire new_Jinkela_wire_21033;
    wire new_Jinkela_wire_15481;
    wire new_Jinkela_wire_6809;
    wire new_Jinkela_wire_7909;
    wire new_Jinkela_wire_16505;
    wire new_Jinkela_wire_19651;
    wire _0978_;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_17451;
    wire new_Jinkela_wire_21171;
    wire new_Jinkela_wire_18777;
    wire new_Jinkela_wire_14610;
    wire new_Jinkela_wire_6237;
    wire new_Jinkela_wire_7238;
    wire new_Jinkela_wire_14723;
    wire new_Jinkela_wire_20142;
    wire _1818_;
    wire new_Jinkela_wire_4924;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_6721;
    wire new_Jinkela_wire_12262;
    wire _0911_;
    wire new_Jinkela_wire_7812;
    wire _0319_;
    wire new_Jinkela_wire_19360;
    wire new_Jinkela_wire_21148;
    wire new_Jinkela_wire_2343;
    wire new_Jinkela_wire_2479;
    wire new_Jinkela_wire_13834;
    wire new_Jinkela_wire_11148;
    wire new_Jinkela_wire_5546;
    wire new_Jinkela_wire_16272;
    wire new_Jinkela_wire_5044;
    wire new_Jinkela_wire_5306;
    wire new_Jinkela_wire_19868;
    wire new_Jinkela_wire_12492;
    wire new_Jinkela_wire_16350;
    wire new_Jinkela_wire_7495;
    wire new_Jinkela_wire_4164;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_3237;
    wire new_Jinkela_wire_18652;
    wire new_Jinkela_wire_14077;
    wire new_Jinkela_wire_21286;
    wire _1338_;
    wire new_Jinkela_wire_15807;
    wire new_Jinkela_wire_16338;
    wire new_Jinkela_wire_17471;
    wire new_Jinkela_wire_10363;
    wire new_Jinkela_wire_4592;
    wire new_Jinkela_wire_14441;
    wire new_Jinkela_wire_17133;
    wire new_Jinkela_wire_2409;
    wire new_Jinkela_wire_10489;
    wire new_Jinkela_wire_18741;
    wire new_Jinkela_wire_10118;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_20274;
    wire new_Jinkela_wire_11580;
    wire new_Jinkela_wire_10794;
    wire new_Jinkela_wire_15914;
    wire new_Jinkela_wire_17477;
    wire new_Jinkela_wire_6936;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_3001;
    wire _1758_;
    wire new_Jinkela_wire_5928;
    wire new_Jinkela_wire_4415;
    wire new_Jinkela_wire_17876;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_4120;
    wire new_Jinkela_wire_12821;
    wire new_Jinkela_wire_7602;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_4681;
    wire new_Jinkela_wire_6863;
    wire new_Jinkela_wire_14093;
    wire new_Jinkela_wire_6708;
    wire new_Jinkela_wire_9268;
    wire _1486_;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_19876;
    wire new_Jinkela_wire_11321;
    wire new_Jinkela_wire_14026;
    wire new_Jinkela_wire_3183;
    wire _0974_;
    wire new_Jinkela_wire_8168;
    wire new_Jinkela_wire_7605;
    wire new_Jinkela_wire_20917;
    wire new_Jinkela_wire_7050;
    wire new_Jinkela_wire_13256;
    wire new_Jinkela_wire_10147;
    wire new_Jinkela_wire_19417;
    wire _1096_;
    wire new_Jinkela_wire_13219;
    wire new_Jinkela_wire_21234;
    wire _0109_;
    wire new_Jinkela_wire_14968;
    wire new_Jinkela_wire_16007;
    wire new_Jinkela_wire_17890;
    wire new_Jinkela_wire_9495;
    wire new_Jinkela_wire_3115;
    wire new_Jinkela_wire_10537;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_7138;
    wire new_Jinkela_wire_14028;
    wire new_Jinkela_wire_16998;
    wire new_Jinkela_wire_11677;
    wire new_Jinkela_wire_5597;
    wire new_Jinkela_wire_1066;
    wire _0579_;
    wire new_Jinkela_wire_17195;
    wire new_Jinkela_wire_15532;
    wire new_Jinkela_wire_17911;
    wire new_Jinkela_wire_18109;
    wire _0318_;
    wire new_Jinkela_wire_3413;
    wire new_Jinkela_wire_3785;
    wire new_Jinkela_wire_19724;
    wire new_Jinkela_wire_3944;
    wire new_Jinkela_wire_7721;
    wire new_Jinkela_wire_8862;
    wire new_Jinkela_wire_14855;
    wire new_Jinkela_wire_8905;
    wire _0800_;
    wire new_Jinkela_wire_18968;
    wire new_Jinkela_wire_10190;
    wire new_Jinkela_wire_20630;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_12487;
    wire new_Jinkela_wire_4385;
    wire new_Jinkela_wire_3535;
    wire new_Jinkela_wire_18757;
    wire new_Jinkela_wire_17832;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_9667;
    wire _0412_;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_9233;
    wire new_Jinkela_wire_2002;
    wire new_Jinkela_wire_4494;
    wire _0851_;
    wire new_Jinkela_wire_8465;
    wire new_Jinkela_wire_10095;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_2014;
    wire new_Jinkela_wire_11288;
    wire new_Jinkela_wire_20187;
    wire new_Jinkela_wire_17268;
    wire new_Jinkela_wire_13727;
    wire new_Jinkela_wire_2761;
    wire new_Jinkela_wire_10073;
    wire new_Jinkela_wire_8206;
    wire new_Jinkela_wire_6752;
    wire _0390_;
    wire new_Jinkela_wire_10235;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_8030;
    wire new_Jinkela_wire_16766;
    wire new_Jinkela_wire_8115;
    wire new_Jinkela_wire_14097;
    wire new_Jinkela_wire_9780;
    wire new_Jinkela_wire_15804;
    wire new_Jinkela_wire_15772;
    wire new_Jinkela_wire_16323;
    wire new_Jinkela_wire_20010;
    wire new_Jinkela_wire_21011;
    wire new_Jinkela_wire_3790;
    wire new_Jinkela_wire_10333;
    wire new_Jinkela_wire_7031;
    wire new_Jinkela_wire_11476;
    wire new_Jinkela_wire_16751;
    wire _0805_;
    wire new_Jinkela_wire_13991;
    wire _0192_;
    wire new_Jinkela_wire_6840;
    wire new_Jinkela_wire_5670;
    wire new_Jinkela_wire_5484;
    wire new_Jinkela_wire_5432;
    wire new_Jinkela_wire_16317;
    wire new_Jinkela_wire_14357;
    wire new_Jinkela_wire_15081;
    wire new_Jinkela_wire_12747;
    wire new_Jinkela_wire_3015;
    wire _0335_;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_4553;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_17709;
    wire new_Jinkela_wire_21245;
    wire new_Jinkela_wire_18475;
    wire new_Jinkela_wire_11078;
    wire new_Jinkela_wire_10164;
    wire new_Jinkela_wire_6268;
    wire new_Jinkela_wire_19584;
    wire new_Jinkela_wire_5469;
    wire new_Jinkela_wire_4577;
    wire new_Jinkela_wire_13255;
    wire new_Jinkela_wire_11395;
    wire new_Jinkela_wire_13215;
    wire new_Jinkela_wire_3537;
    wire new_Jinkela_wire_10559;
    wire new_Jinkela_wire_3144;
    wire new_Jinkela_wire_14806;
    wire new_Jinkela_wire_17803;
    wire new_Jinkela_wire_19029;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_5515;
    wire new_Jinkela_wire_1997;
    wire new_Jinkela_wire_10318;
    wire _1133_;
    wire new_Jinkela_wire_17685;
    wire new_Jinkela_wire_17335;
    wire new_Jinkela_wire_17607;
    wire new_Jinkela_wire_5017;
    wire new_Jinkela_wire_8012;
    wire new_Jinkela_wire_6876;
    wire new_Jinkela_wire_17494;
    wire new_Jinkela_wire_4519;
    wire new_Jinkela_wire_7161;
    wire new_Jinkela_wire_10567;
    wire new_Jinkela_wire_8637;
    wire new_Jinkela_wire_9330;
    wire _1738_;
    wire new_Jinkela_wire_6919;
    wire new_Jinkela_wire_19245;
    wire new_Jinkela_wire_13688;
    wire new_Jinkela_wire_10913;
    wire new_Jinkela_wire_12132;
    wire new_Jinkela_wire_5359;
    wire new_Jinkela_wire_8915;
    wire new_Jinkela_wire_20777;
    wire new_Jinkela_wire_6082;
    wire new_Jinkela_wire_17904;
    wire new_Jinkela_wire_20081;
    wire new_Jinkela_wire_14676;
    wire new_Jinkela_wire_9716;
    wire new_Jinkela_wire_14082;
    wire new_Jinkela_wire_5865;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_13952;
    wire new_Jinkela_wire_12403;
    wire new_Jinkela_wire_17098;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_1678;
    wire _1413_;
    wire new_Jinkela_wire_14234;
    wire new_Jinkela_wire_7683;
    wire _1593_;
    wire new_Jinkela_wire_4997;
    wire new_Jinkela_wire_18571;
    wire _0905_;
    wire new_Jinkela_wire_10682;
    wire new_Jinkela_wire_7208;
    wire new_Jinkela_wire_18619;
    wire new_Jinkela_wire_7018;
    wire new_Jinkela_wire_20656;
    wire new_Jinkela_wire_17169;
    wire new_Jinkela_wire_7439;
    wire new_Jinkela_wire_3370;
    wire new_Jinkela_wire_8883;
    wire _1519_;
    wire new_Jinkela_wire_13928;
    wire new_Jinkela_wire_2172;
    wire new_Jinkela_wire_7600;
    wire _0236_;
    wire new_Jinkela_wire_18371;
    wire _0712_;
    wire new_Jinkela_wire_17334;
    wire new_Jinkela_wire_17434;
    wire new_Jinkela_wire_12888;
    wire new_Jinkela_wire_17352;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_8049;
    wire new_Jinkela_wire_2976;
    wire new_Jinkela_wire_13452;
    wire new_Jinkela_wire_15057;
    wire new_Jinkela_wire_9503;
    wire new_Jinkela_wire_19314;
    wire new_Jinkela_wire_13904;
    wire new_Jinkela_wire_17374;
    wire new_Jinkela_wire_9416;
    wire new_Jinkela_wire_5030;
    wire new_Jinkela_wire_5521;
    wire new_Jinkela_wire_10365;
    wire new_Jinkela_wire_20330;
    wire new_Jinkela_wire_19675;
    wire new_Jinkela_wire_20991;
    wire new_Jinkela_wire_3332;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_5697;
    wire _0535_;
    wire new_Jinkela_wire_1420;
    wire new_Jinkela_wire_14598;
    wire new_Jinkela_wire_4986;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_16311;
    wire new_Jinkela_wire_17780;
    wire _1070_;
    wire _0051_;
    wire new_Jinkela_wire_14030;
    wire _0016_;
    wire new_Jinkela_wire_3788;
    wire new_Jinkela_wire_13198;
    wire new_Jinkela_wire_16887;
    wire new_Jinkela_wire_5885;
    wire new_Jinkela_wire_19965;
    wire new_Jinkela_wire_6243;
    wire new_Jinkela_wire_13789;
    wire new_Jinkela_wire_15240;
    wire new_Jinkela_wire_14419;
    wire new_Jinkela_wire_10284;
    wire new_Jinkela_wire_12844;
    wire new_Jinkela_wire_21064;
    wire new_Jinkela_wire_10383;
    wire new_Jinkela_wire_12944;
    wire new_Jinkela_wire_8469;
    wire new_Jinkela_wire_16116;
    wire new_Jinkela_wire_5905;
    wire new_Jinkela_wire_634;
    wire _0739_;
    wire new_Jinkela_wire_14664;
    wire new_Jinkela_wire_7572;
    wire new_Jinkela_wire_12728;
    wire new_Jinkela_wire_11053;
    wire new_Jinkela_wire_3600;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_10323;
    wire new_Jinkela_wire_12017;
    wire new_Jinkela_wire_5005;
    wire new_Jinkela_wire_21137;
    wire new_Jinkela_wire_10271;
    wire _1104_;
    wire _1051_;
    wire new_Jinkela_wire_17627;
    wire new_Jinkela_wire_6566;
    wire new_Jinkela_wire_15442;
    wire new_Jinkela_wire_19751;
    wire new_Jinkela_wire_20143;
    wire new_Jinkela_wire_2713;
    wire new_Jinkela_wire_13977;
    wire new_Jinkela_wire_2321;
    wire new_Jinkela_wire_2443;
    wire new_Jinkela_wire_5346;
    wire new_Jinkela_wire_14470;
    wire _0098_;
    wire _0479_;
    wire _1334_;
    wire new_Jinkela_wire_17733;
    wire new_Jinkela_wire_6585;
    wire new_Jinkela_wire_18593;
    wire new_Jinkela_wire_3093;
    wire new_Jinkela_wire_9615;
    wire _0464_;
    wire new_Jinkela_wire_6138;
    wire new_Jinkela_wire_15345;
    wire new_Jinkela_wire_14927;
    wire new_Jinkela_wire_17969;
    wire new_Jinkela_wire_5994;
    wire new_Jinkela_wire_18996;
    wire new_Jinkela_wire_13015;
    wire new_Jinkela_wire_17266;
    wire new_Jinkela_wire_13441;
    wire new_Jinkela_wire_5629;
    wire new_Jinkela_wire_18738;
    wire new_Jinkela_wire_9751;
    wire new_Jinkela_wire_13509;
    wire new_Jinkela_wire_19631;
    wire new_Jinkela_wire_9028;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_20995;
    wire new_Jinkela_wire_2142;
    wire new_Jinkela_wire_14193;
    wire _0813_;
    wire new_Jinkela_wire_17456;
    wire new_Jinkela_wire_20602;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_3051;
    wire new_Jinkela_wire_10187;
    wire new_Jinkela_wire_5372;
    wire new_Jinkela_wire_13773;
    wire new_Jinkela_wire_8282;
    wire new_Jinkela_wire_3014;
    wire new_Jinkela_wire_18903;
    wire new_Jinkela_wire_15884;
    wire new_Jinkela_wire_15292;
    wire new_Jinkela_wire_2828;
    wire new_Jinkela_wire_19447;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_20852;
    wire new_Jinkela_wire_2789;
    wire new_Jinkela_wire_2727;
    wire new_Jinkela_wire_18356;
    wire new_Jinkela_wire_16913;
    wire new_Jinkela_wire_3292;
    wire new_Jinkela_wire_11388;
    wire new_Jinkela_wire_2433;
    wire new_Jinkela_wire_7944;
    wire new_Jinkela_wire_16296;
    wire _0346_;
    wire new_Jinkela_wire_3312;
    wire new_Jinkela_wire_13832;
    wire new_Jinkela_wire_20558;
    wire new_Jinkela_wire_9345;
    wire new_Jinkela_wire_8799;
    wire new_Jinkela_wire_8657;
    wire new_Jinkela_wire_5063;
    wire new_Jinkela_wire_19091;
    wire _1569_;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_14911;
    wire new_Jinkela_wire_6827;
    wire new_Jinkela_wire_3754;
    wire new_Jinkela_wire_11031;
    wire new_Jinkela_wire_6693;
    wire new_Jinkela_wire_7196;
    wire new_Jinkela_wire_17022;
    wire new_Jinkela_wire_16750;
    wire _0847_;
    wire new_Jinkela_wire_20335;
    wire new_Jinkela_wire_16211;
    wire new_Jinkela_wire_12015;
    wire new_Jinkela_wire_5293;
    wire new_Jinkela_wire_7582;
    wire new_Jinkela_wire_19422;
    wire new_Jinkela_wire_469;
    wire _1827_;
    wire new_Jinkela_wire_12314;
    wire new_Jinkela_wire_6468;
    wire new_Jinkela_wire_15717;
    wire new_Jinkela_wire_16762;
    wire _1479_;
    wire new_Jinkela_wire_10832;
    wire new_Jinkela_wire_20332;
    wire new_Jinkela_wire_3016;
    wire _0491_;
    wire new_Jinkela_wire_11916;
    wire new_Jinkela_wire_2737;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_14404;
    wire new_Jinkela_wire_1219;
    wire _1528_;
    wire new_Jinkela_wire_3245;
    wire new_Jinkela_wire_2923;
    wire new_Jinkela_wire_12463;
    wire new_Jinkela_wire_14935;
    wire new_Jinkela_wire_10934;
    wire new_Jinkela_wire_4799;
    wire new_Jinkela_wire_20431;
    wire new_Jinkela_wire_9508;
    wire new_Jinkela_wire_5077;
    wire new_Jinkela_wire_13892;
    wire new_Jinkela_wire_12102;
    wire new_Jinkela_wire_10053;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_11970;
    wire new_Jinkela_wire_6792;
    wire new_Jinkela_wire_13038;
    wire new_Jinkela_wire_6022;
    wire new_Jinkela_wire_1483;
    wire _1099_;
    wire new_Jinkela_wire_9218;
    wire new_Jinkela_wire_1978;
    wire new_Jinkela_wire_10114;
    wire new_Jinkela_wire_2640;
    wire new_Jinkela_wire_3180;
    wire _1435_;
    wire new_Jinkela_wire_17316;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_15583;
    wire _1378_;
    wire new_Jinkela_wire_5824;
    wire new_Jinkela_wire_11844;
    wire new_Jinkela_wire_3811;
    wire new_Jinkela_wire_11688;
    wire new_Jinkela_wire_6469;
    wire new_Jinkela_wire_20502;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_4566;
    wire new_Jinkela_wire_16060;
    wire new_Jinkela_wire_9254;
    wire new_Jinkela_wire_20498;
    wire _0438_;
    wire new_Jinkela_wire_7012;
    wire new_Jinkela_wire_13556;
    wire new_Jinkela_wire_7527;
    wire new_Jinkela_wire_3957;
    wire new_Jinkela_wire_17513;
    wire new_Jinkela_wire_5961;
    wire new_Jinkela_wire_21131;
    wire new_Jinkela_wire_2120;
    wire _0914_;
    wire new_Jinkela_wire_5429;
    wire new_Jinkela_wire_12199;
    wire new_Jinkela_wire_4521;
    wire new_Jinkela_wire_12106;
    wire _0193_;
    wire new_Jinkela_wire_4295;
    wire new_Jinkela_wire_16826;
    wire new_Jinkela_wire_4625;
    wire new_Jinkela_wire_20032;
    wire new_Jinkela_wire_20231;
    wire new_Jinkela_wire_1016;
    wire _1779_;
    wire new_Jinkela_wire_10337;
    wire new_Jinkela_wire_4363;
    wire new_Jinkela_wire_13893;
    wire new_Jinkela_wire_14446;
    wire new_Jinkela_wire_3073;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_11919;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_7616;
    wire new_Jinkela_wire_15834;
    wire new_Jinkela_wire_8670;
    wire new_Jinkela_wire_7213;
    wire new_Jinkela_wire_10922;
    wire new_Jinkela_wire_15022;
    wire new_Jinkela_wire_13986;
    wire new_Jinkela_wire_20791;
    wire new_Jinkela_wire_20619;
    wire new_Jinkela_wire_7496;
    wire new_Jinkela_wire_5315;
    wire new_Jinkela_wire_11230;
    wire new_Jinkela_wire_11251;
    wire new_Jinkela_wire_8590;
    wire _0070_;
    wire new_Jinkela_wire_3575;
    wire new_Jinkela_wire_16208;
    wire new_Jinkela_wire_20281;
    wire new_Jinkela_wire_16488;
    wire new_Jinkela_wire_9431;
    wire new_Jinkela_wire_12678;
    wire new_Jinkela_wire_21050;
    wire new_Jinkela_wire_15907;
    wire new_Jinkela_wire_19828;
    wire new_Jinkela_wire_11004;
    wire new_Jinkela_wire_5327;
    wire new_Jinkela_wire_19572;
    wire new_Jinkela_wire_9361;
    wire new_Jinkela_wire_4374;
    wire new_Jinkela_wire_6961;
    wire new_Jinkela_wire_5013;
    wire new_Jinkela_wire_17041;
    wire new_Jinkela_wire_17548;
    wire new_Jinkela_wire_17615;
    wire new_Jinkela_wire_8492;
    wire new_Jinkela_wire_15032;
    wire new_net_3928;
    wire new_Jinkela_wire_5911;
    wire new_Jinkela_wire_2684;
    wire _0953_;
    wire new_Jinkela_wire_13604;
    wire new_Jinkela_wire_11462;
    wire _0754_;
    wire new_Jinkela_wire_5531;
    wire new_Jinkela_wire_20806;
    wire new_Jinkela_wire_19097;
    wire new_Jinkela_wire_12217;
    wire new_Jinkela_wire_16728;
    wire new_Jinkela_wire_18298;
    wire new_Jinkela_wire_6465;
    wire new_Jinkela_wire_13431;
    wire new_Jinkela_wire_19859;
    wire new_Jinkela_wire_18351;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_3815;
    wire new_Jinkela_wire_20675;
    wire new_Jinkela_wire_5297;
    wire new_Jinkela_wire_12288;
    wire new_Jinkela_wire_12049;
    wire _0811_;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_8859;
    wire new_Jinkela_wire_18459;
    wire new_Jinkela_wire_11910;
    wire new_Jinkela_wire_17888;
    wire new_Jinkela_wire_8769;
    wire new_Jinkela_wire_12259;
    wire new_Jinkela_wire_11912;
    wire new_Jinkela_wire_17019;
    wire new_Jinkela_wire_7022;
    wire new_Jinkela_wire_10420;
    wire _1527_;
    wire new_Jinkela_wire_18242;
    wire new_Jinkela_wire_18818;
    wire new_Jinkela_wire_5281;
    wire new_Jinkela_wire_18994;
    wire new_Jinkela_wire_11217;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_18555;
    wire new_Jinkela_wire_2447;
    wire new_Jinkela_wire_3775;
    wire new_Jinkela_wire_6914;
    wire new_Jinkela_wire_12775;
    wire _0684_;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_3968;
    wire new_Jinkela_wire_5527;
    wire new_Jinkela_wire_4817;
    wire new_Jinkela_wire_16809;
    wire new_Jinkela_wire_8824;
    wire _0598_;
    wire _1135_;
    wire new_Jinkela_wire_17006;
    wire new_Jinkela_wire_20738;
    wire new_Jinkela_wire_17226;
    wire new_Jinkela_wire_13774;
    wire new_Jinkela_wire_8374;
    wire new_Jinkela_wire_14618;
    wire new_Jinkela_wire_17085;
    wire _1698_;
    wire new_Jinkela_wire_10397;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_17518;
    wire new_Jinkela_wire_15282;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_12333;
    wire new_Jinkela_wire_13857;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_15111;
    wire new_Jinkela_wire_14486;
    wire new_Jinkela_wire_13449;
    wire new_Jinkela_wire_13515;
    wire _1419_;
    wire new_Jinkela_wire_13586;
    wire new_Jinkela_wire_11891;
    wire new_Jinkela_wire_11763;
    wire new_Jinkela_wire_6017;
    wire new_Jinkela_wire_13609;
    wire new_Jinkela_wire_7913;
    wire new_Jinkela_wire_16981;
    wire _0062_;
    wire new_Jinkela_wire_16158;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_4246;
    wire new_Jinkela_wire_10959;
    wire new_Jinkela_wire_5894;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_4474;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_7477;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_17239;
    wire _1206_;
    wire new_Jinkela_wire_16145;
    wire new_Jinkela_wire_18855;
    wire new_Jinkela_wire_9101;
    wire _1754_;
    wire new_Jinkela_wire_14894;
    wire new_Jinkela_wire_17527;
    wire new_Jinkela_wire_19681;
    wire _0476_;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_3351;
    wire new_Jinkela_wire_15233;
    wire _1052_;
    wire _1192_;
    wire new_Jinkela_wire_16043;
    wire new_Jinkela_wire_17631;
    wire new_Jinkela_wire_20564;
    wire new_Jinkela_wire_9341;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_1740;
    wire new_Jinkela_wire_16107;
    wire new_Jinkela_wire_4977;
    wire new_Jinkela_wire_7752;
    wire new_Jinkela_wire_4300;
    wire new_Jinkela_wire_9532;
    wire new_Jinkela_wire_10336;
    wire new_Jinkela_wire_10663;
    wire new_Jinkela_wire_7368;
    wire new_Jinkela_wire_4716;
    wire new_Jinkela_wire_8396;
    wire new_Jinkela_wire_9905;
    wire new_Jinkela_wire_15203;
    wire new_Jinkela_wire_7557;
    wire new_Jinkela_wire_7292;
    wire new_Jinkela_wire_2081;
    wire new_Jinkela_wire_20067;
    wire _0432_;
    wire new_Jinkela_wire_2336;
    wire new_Jinkela_wire_10786;
    wire _1183_;
    wire new_Jinkela_wire_11553;
    wire new_Jinkela_wire_3407;
    wire new_Jinkela_wire_12969;
    wire new_Jinkela_wire_13250;
    wire new_Jinkela_wire_5417;
    wire new_Jinkela_wire_16506;
    wire new_Jinkela_wire_3671;
    wire _1614_;
    wire new_Jinkela_wire_3728;
    wire new_Jinkela_wire_18184;
    wire _0898_;
    wire new_Jinkela_wire_8457;
    wire new_Jinkela_wire_14745;
    wire new_Jinkela_wire_11277;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_1631;
    wire _0135_;
    wire new_Jinkela_wire_5745;
    wire _1759_;
    wire new_Jinkela_wire_16886;
    wire new_Jinkela_wire_3802;
    wire new_Jinkela_wire_10843;
    wire new_Jinkela_wire_18998;
    wire _0925_;
    wire new_Jinkela_wire_9211;
    wire new_Jinkela_wire_19625;
    wire _1478_;
    wire new_Jinkela_wire_3523;
    wire new_Jinkela_wire_8950;
    wire new_Jinkela_wire_15937;
    wire new_Jinkela_wire_14915;
    wire _1295_;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_8345;
    wire new_Jinkela_wire_15588;
    wire new_Jinkela_wire_9772;
    wire new_Jinkela_wire_5441;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_4873;
    wire new_Jinkela_wire_17446;
    wire new_Jinkela_wire_20202;
    wire new_Jinkela_wire_10357;
    wire _1041_;
    wire new_Jinkela_wire_21156;
    wire new_Jinkela_wire_15347;
    wire new_Jinkela_wire_18186;
    wire new_Jinkela_wire_18418;
    wire new_Jinkela_wire_12150;
    wire new_Jinkela_wire_16570;
    wire new_Jinkela_wire_16588;
    wire new_Jinkela_wire_18000;
    wire new_Jinkela_wire_12458;
    wire new_Jinkela_wire_19759;
    wire new_Jinkela_wire_2551;
    wire new_Jinkela_wire_12271;
    wire new_Jinkela_wire_6291;
    wire new_Jinkela_wire_15076;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_17698;
    wire new_Jinkela_wire_4735;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_10344;
    wire new_Jinkela_wire_19138;
    wire new_Jinkela_wire_17216;
    wire _0241_;
    wire new_Jinkela_wire_17343;
    wire new_Jinkela_wire_8868;
    wire new_Jinkela_wire_4640;
    wire new_Jinkela_wire_17459;
    wire new_Jinkela_wire_18102;
    wire new_Jinkela_wire_12336;
    wire new_Jinkela_wire_7104;
    wire new_Jinkela_wire_6264;
    wire new_Jinkela_wire_17115;
    wire new_Jinkela_wire_20977;
    wire new_Jinkela_wire_16634;
    wire new_Jinkela_wire_5145;
    wire new_Jinkela_wire_4482;
    wire new_Jinkela_wire_12207;
    wire new_Jinkela_wire_14567;
    wire new_Jinkela_wire_838;
    wire _1787_;
    wire new_Jinkela_wire_2283;
    wire new_Jinkela_wire_3220;
    wire new_Jinkela_wire_7299;
    wire new_Jinkela_wire_17047;
    wire new_Jinkela_wire_12607;
    wire new_Jinkela_wire_13085;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_6561;
    wire new_Jinkela_wire_21017;
    wire new_Jinkela_wire_21004;
    wire new_Jinkela_wire_8622;
    wire _0651_;
    wire new_Jinkela_wire_7771;
    wire new_Jinkela_wire_14105;
    wire new_Jinkela_wire_15197;
    wire new_Jinkela_wire_14135;
    wire _0371_;
    wire new_Jinkela_wire_20646;
    wire new_Jinkela_wire_8552;
    wire new_Jinkela_wire_11843;
    wire new_Jinkela_wire_18423;
    wire new_Jinkela_wire_13130;
    wire new_Jinkela_wire_4596;
    wire new_Jinkela_wire_12221;
    wire new_Jinkela_wire_17864;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_6132;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_16321;
    wire new_Jinkela_wire_2565;
    wire new_Jinkela_wire_21167;
    wire new_Jinkela_wire_18456;
    wire new_Jinkela_wire_2711;
    wire new_Jinkela_wire_10749;
    wire new_Jinkela_wire_11760;
    wire new_Jinkela_wire_11900;
    wire new_Jinkela_wire_15742;
    wire new_Jinkela_wire_6846;
    wire new_Jinkela_wire_4239;
    wire new_Jinkela_wire_19408;
    wire new_Jinkela_wire_14506;
    wire new_Jinkela_wire_4472;
    wire new_Jinkela_wire_8278;
    wire new_Jinkela_wire_6589;
    wire new_Jinkela_wire_19961;
    wire new_Jinkela_wire_19369;
    wire new_Jinkela_wire_4463;
    wire new_Jinkela_wire_16802;
    wire new_Jinkela_wire_5113;
    wire _1029_;
    wire new_Jinkela_wire_6112;
    wire new_Jinkela_wire_7276;
    wire new_Jinkela_wire_11675;
    wire new_Jinkela_wire_6624;
    wire new_Jinkela_wire_12021;
    wire new_Jinkela_wire_14108;
    wire new_Jinkela_wire_8517;
    wire new_Jinkela_wire_4154;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_18159;
    wire new_Jinkela_wire_18624;
    wire new_Jinkela_wire_9522;
    wire new_Jinkela_wire_2453;
    wire new_Jinkela_wire_6105;
    wire new_Jinkela_wire_7172;
    wire new_Jinkela_wire_14224;
    wire _0315_;
    wire new_Jinkela_wire_18431;
    wire new_Jinkela_wire_6545;
    wire new_Jinkela_wire_7685;
    wire new_Jinkela_wire_2908;
    wire new_Jinkela_wire_13976;
    wire new_Jinkela_wire_20743;
    wire new_Jinkela_wire_16885;
    wire new_Jinkela_wire_14526;
    wire new_Jinkela_wire_527;
    wire _1092_;
    wire _0779_;
    wire new_Jinkela_wire_17287;
    wire new_Jinkela_wire_19835;
    wire new_Jinkela_wire_17968;
    wire new_Jinkela_wire_20570;
    wire new_Jinkela_wire_19634;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_477;
    wire new_Jinkela_wire_19953;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_13365;
    wire new_Jinkela_wire_20834;
    wire new_Jinkela_wire_16659;
    wire new_Jinkela_wire_13925;
    wire new_Jinkela_wire_9747;
    wire new_Jinkela_wire_16324;
    wire new_Jinkela_wire_18390;
    wire new_Jinkela_wire_6236;
    wire new_Jinkela_wire_5912;
    wire new_Jinkela_wire_3839;
    wire new_Jinkela_wire_2936;
    wire new_Jinkela_wire_11330;
    wire new_Jinkela_wire_10809;
    wire new_Jinkela_wire_10391;
    wire new_Jinkela_wire_14751;
    wire new_Jinkela_wire_8896;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_15413;
    wire new_Jinkela_wire_20840;
    wire new_Jinkela_wire_15114;
    wire new_Jinkela_wire_17256;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_5149;
    wire new_Jinkela_wire_3477;
    wire new_Jinkela_wire_7736;
    wire new_Jinkela_wire_13700;
    wire new_Jinkela_wire_7507;
    wire new_Jinkela_wire_8923;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_5465;
    wire _1651_;
    wire new_Jinkela_wire_12503;
    wire new_Jinkela_wire_17843;
    wire new_Jinkela_wire_12629;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_7869;
    wire new_Jinkela_wire_19292;
    wire _1298_;
    wire new_Jinkela_wire_13071;
    wire new_Jinkela_wire_12670;
    wire new_Jinkela_wire_13642;
    wire new_Jinkela_wire_15091;
    wire new_Jinkela_wire_9547;
    wire new_Jinkela_wire_14674;
    wire new_Jinkela_wire_15747;
    wire new_Jinkela_wire_17185;
    wire new_Jinkela_wire_3173;
    wire _1241_;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_8566;
    wire new_Jinkela_wire_18178;
    wire new_Jinkela_wire_2312;
    wire new_Jinkela_wire_5711;
    wire new_Jinkela_wire_6103;
    wire new_Jinkela_wire_8065;
    wire new_Jinkela_wire_8342;
    wire new_Jinkela_wire_8427;
    wire new_Jinkela_wire_8965;
    wire _1733_;
    wire new_Jinkela_wire_8851;
    wire new_Jinkela_wire_15586;
    wire new_Jinkela_wire_13226;
    wire new_Jinkela_wire_14601;
    wire new_Jinkela_wire_18136;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_19190;
    wire new_Jinkela_wire_8678;
    wire new_Jinkela_wire_3043;
    wire new_Jinkela_wire_19075;
    wire new_Jinkela_wire_9085;
    wire new_Jinkela_wire_15033;
    wire new_Jinkela_wire_19921;
    wire new_Jinkela_wire_6395;
    wire new_Jinkela_wire_12505;
    wire new_Jinkela_wire_6883;
    wire new_Jinkela_wire_20188;
    wire new_Jinkela_wire_10569;
    wire new_Jinkela_wire_6891;
    wire new_Jinkela_wire_6146;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_19194;
    wire new_Jinkela_wire_10123;
    wire new_Jinkela_wire_11649;
    wire _0526_;
    wire new_Jinkela_wire_11815;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_11313;
    wire new_Jinkela_wire_4042;
    wire _1353_;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_7485;
    wire new_Jinkela_wire_14096;
    wire new_Jinkela_wire_17959;
    wire new_Jinkela_wire_7945;
    wire _0441_;
    wire new_Jinkela_wire_16039;
    wire new_Jinkela_wire_11049;
    wire new_Jinkela_wire_11948;
    wire new_Jinkela_wire_12707;
    wire new_Jinkela_wire_20363;
    wire new_Jinkela_wire_2723;
    wire new_Jinkela_wire_15840;
    wire new_Jinkela_wire_2296;
    wire new_Jinkela_wire_12694;
    wire new_Jinkela_wire_14188;
    wire new_Jinkela_wire_14303;
    wire new_Jinkela_wire_5614;
    wire _1256_;
    wire new_Jinkela_wire_10742;
    wire new_Jinkela_wire_2489;
    wire new_Jinkela_wire_2975;
    wire new_Jinkela_wire_15719;
    wire new_Jinkela_wire_18200;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_3753;
    wire new_Jinkela_wire_4800;
    wire _0145_;
    wire new_Jinkela_wire_16583;
    wire new_Jinkela_wire_16075;
    wire new_Jinkela_wire_17392;
    wire new_Jinkela_wire_10371;
    wire new_Jinkela_wire_18082;
    wire new_Jinkela_wire_8361;
    wire new_Jinkela_wire_10723;
    wire new_Jinkela_wire_16210;
    wire new_Jinkela_wire_17664;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_8257;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_7320;
    wire new_Jinkela_wire_9609;
    wire new_Jinkela_wire_15889;
    wire new_Jinkela_wire_1781;
    wire new_Jinkela_wire_4024;
    wire new_Jinkela_wire_13285;
    wire new_Jinkela_wire_19509;
    wire new_Jinkela_wire_9534;
    wire new_Jinkela_wire_19472;
    wire new_Jinkela_wire_12836;
    wire new_Jinkela_wire_18786;
    wire new_Jinkela_wire_13583;
    wire new_Jinkela_wire_10946;
    wire new_Jinkela_wire_20884;
    wire new_Jinkela_wire_10196;
    wire new_Jinkela_wire_13992;
    wire new_Jinkela_wire_1498;
    wire _0376_;
    wire new_Jinkela_wire_17753;
    wire new_Jinkela_wire_2810;
    wire new_Jinkela_wire_20150;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_5942;
    wire new_Jinkela_wire_5838;
    wire new_Jinkela_wire_6271;
    wire new_Jinkela_wire_17669;
    wire new_Jinkela_wire_10244;
    wire new_Jinkela_wire_15258;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_12429;
    wire new_Jinkela_wire_9557;
    wire new_Jinkela_wire_2236;
    wire _0642_;
    wire new_Jinkela_wire_7529;
    wire new_Jinkela_wire_7782;
    wire _1097_;
    wire new_Jinkela_wire_20861;
    wire new_Jinkela_wire_9042;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_2246;
    wire new_Jinkela_wire_7147;
    wire new_Jinkela_wire_14684;
    wire new_Jinkela_wire_18788;
    wire new_Jinkela_wire_7758;
    wire new_Jinkela_wire_10876;
    wire new_Jinkela_wire_4429;
    wire new_Jinkela_wire_15609;
    wire new_Jinkela_wire_19025;
    wire new_Jinkela_wire_13129;
    wire new_Jinkela_wire_19358;
    wire new_Jinkela_wire_15754;
    wire _0225_;
    wire new_Jinkela_wire_9324;
    wire new_Jinkela_wire_19122;
    wire _0861_;
    wire _0594_;
    wire _1053_;
    wire new_Jinkela_wire_5682;
    wire new_Jinkela_wire_11852;
    wire new_Jinkela_wire_13993;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_10253;
    wire new_Jinkela_wire_12936;
    wire new_Jinkela_wire_10379;
    wire new_Jinkela_wire_18148;
    wire new_Jinkela_wire_7431;
    wire new_Jinkela_wire_7141;
    wire new_Jinkela_wire_15706;
    wire new_Jinkela_wire_4678;
    wire new_Jinkela_wire_14208;
    wire new_Jinkela_wire_7150;
    wire new_Jinkela_wire_14680;
    wire _1007_;
    wire new_Jinkela_wire_19721;
    wire new_Jinkela_wire_11752;
    wire new_Jinkela_wire_21062;
    wire new_Jinkela_wire_17736;
    wire new_Jinkela_wire_20248;
    wire new_Jinkela_wire_21112;
    wire _0548_;
    wire new_Jinkela_wire_5520;
    wire new_Jinkela_wire_14626;
    wire new_Jinkela_wire_9262;
    wire new_Jinkela_wire_8231;
    wire new_Jinkela_wire_18007;
    wire new_Jinkela_wire_6283;
    wire new_Jinkela_wire_10801;
    wire new_Jinkela_wire_5922;
    wire new_Jinkela_wire_14175;
    wire new_Jinkela_wire_11312;
    wire new_Jinkela_wire_15177;
    wire new_Jinkela_wire_18040;
    wire new_Jinkela_wire_9146;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_15306;
    wire new_Jinkela_wire_5778;
    wire new_Jinkela_wire_15810;
    wire new_Jinkela_wire_9629;
    wire new_Jinkela_wire_20922;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_7727;
    wire new_Jinkela_wire_11459;
    wire new_Jinkela_wire_10799;
    wire new_Jinkela_wire_7544;
    wire new_Jinkela_wire_12421;
    wire new_Jinkela_wire_7849;
    wire new_Jinkela_wire_16859;
    wire _1073_;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_6610;
    wire new_Jinkela_wire_17409;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_13381;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_110;
    wire _1327_;
    wire new_Jinkela_wire_5283;
    wire new_Jinkela_wire_9598;
    wire new_Jinkela_wire_16519;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_8555;
    wire new_Jinkela_wire_3553;
    wire new_Jinkela_wire_7415;
    wire new_Jinkela_wire_3406;
    wire new_Jinkela_wire_12109;
    wire new_Jinkela_wire_4882;
    wire new_Jinkela_wire_21074;
    wire new_Jinkela_wire_12506;
    wire new_Jinkela_wire_3784;
    wire new_Jinkela_wire_6366;
    wire new_Jinkela_wire_6021;
    wire new_Jinkela_wire_10255;
    wire new_Jinkela_wire_9032;
    wire new_Jinkela_wire_5328;
    wire new_Jinkela_wire_3108;
    wire new_Jinkela_wire_6509;
    wire new_Jinkela_wire_11403;
    wire new_Jinkela_wire_11892;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_12158;
    wire new_Jinkela_wire_3820;
    wire new_Jinkela_wire_4307;
    wire new_Jinkela_wire_16529;
    wire new_Jinkela_wire_12183;
    wire new_Jinkela_wire_2163;
    wire new_Jinkela_wire_2269;
    wire new_Jinkela_wire_8516;
    wire new_Jinkela_wire_17271;
    wire new_Jinkela_wire_17469;
    wire new_Jinkela_wire_15897;
    wire new_Jinkela_wire_10130;
    wire new_Jinkela_wire_13533;
    wire new_Jinkela_wire_8882;
    wire new_Jinkela_wire_16102;
    wire new_Jinkela_wire_11215;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_3019;
    wire new_Jinkela_wire_1748;
    wire new_Jinkela_wire_7929;
    wire new_Jinkela_wire_20152;
    wire new_Jinkela_wire_5687;
    wire new_Jinkela_wire_20584;
    wire new_Jinkela_wire_12578;
    wire new_Jinkela_wire_5825;
    wire new_Jinkela_wire_6098;
    wire new_Jinkela_wire_19898;
    wire new_Jinkela_wire_15701;
    wire new_Jinkela_wire_5550;
    wire new_Jinkela_wire_12950;
    wire new_Jinkela_wire_3585;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_16861;
    wire new_Jinkela_wire_6316;
    wire _0962_;
    wire new_Jinkela_wire_4672;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_16534;
    wire new_Jinkela_wire_18731;
    wire new_Jinkela_wire_12070;
    wire new_Jinkela_wire_18308;
    wire new_Jinkela_wire_3980;
    wire new_Jinkela_wire_18706;
    wire new_Jinkela_wire_4371;
    wire new_Jinkela_wire_14709;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_20555;
    wire new_Jinkela_wire_1934;
    wire new_Jinkela_wire_20263;
    wire new_Jinkela_wire_6608;
    wire new_Jinkela_wire_20859;
    wire new_Jinkela_wire_9043;
    wire new_Jinkela_wire_5897;
    wire new_Jinkela_wire_8546;
    wire new_Jinkela_wire_12572;
    wire new_Jinkela_wire_4826;
    wire new_Jinkela_wire_2105;
    wire new_Jinkela_wire_1991;
    wire _1131_;
    wire new_Jinkela_wire_15833;
    wire new_Jinkela_wire_12020;
    wire _1343_;
    wire new_Jinkela_wire_13443;
    wire new_Jinkela_wire_17365;
    wire new_Jinkela_wire_3730;
    wire new_Jinkela_wire_19578;
    wire new_Jinkela_wire_3241;
    wire new_Jinkela_wire_2682;
    wire new_Jinkela_wire_2072;
    wire new_Jinkela_wire_15849;
    wire new_Jinkela_wire_7687;
    wire new_Jinkela_wire_15017;
    wire new_Jinkela_wire_15191;
    wire new_Jinkela_wire_2896;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_16745;
    wire new_Jinkela_wire_11885;
    wire new_Jinkela_wire_8117;
    wire new_Jinkela_wire_21309;
    wire new_Jinkela_wire_14920;
    wire new_Jinkela_wire_18798;
    wire _0478_;
    wire new_Jinkela_wire_4803;
    wire new_Jinkela_wire_6437;
    wire new_Jinkela_wire_10385;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_17974;
    wire _0004_;
    wire new_Jinkela_wire_17971;
    wire new_Jinkela_wire_3201;
    wire new_Jinkela_wire_20887;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_8143;
    wire new_Jinkela_wire_19557;
    wire _1386_;
    wire new_Jinkela_wire_19446;
    wire new_Jinkela_wire_11091;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_16595;
    wire new_Jinkela_wire_2833;
    wire new_Jinkela_wire_16494;
    wire new_Jinkela_wire_6599;
    wire new_Jinkela_wire_13407;
    wire new_Jinkela_wire_8751;
    wire new_Jinkela_wire_14788;
    wire _1255_;
    wire new_Jinkela_wire_15716;
    wire new_Jinkela_wire_17682;
    wire new_Jinkela_wire_9683;
    wire new_Jinkela_wire_9900;
    wire new_Jinkela_wire_17481;
    wire new_Jinkela_wire_12455;
    wire new_Jinkela_wire_20778;
    wire new_Jinkela_wire_13087;
    wire new_Jinkela_wire_18481;
    wire new_Jinkela_wire_6406;
    wire new_Jinkela_wire_9096;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_20241;
    wire new_Jinkela_wire_5046;
    wire new_Jinkela_wire_12067;
    wire new_Jinkela_wire_3130;
    wire new_Jinkela_wire_2118;
    wire new_Jinkela_wire_13638;
    wire new_Jinkela_wire_15525;
    wire new_Jinkela_wire_6773;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_6096;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_11382;
    wire new_Jinkela_wire_11945;
    wire new_Jinkela_wire_7123;
    wire new_Jinkela_wire_3529;
    wire new_Jinkela_wire_7518;
    wire new_Jinkela_wire_18014;
    wire new_Jinkela_wire_17416;
    wire new_Jinkela_wire_8450;
    wire new_Jinkela_wire_3116;
    wire new_Jinkela_wire_5888;
    wire new_Jinkela_wire_8290;
    wire new_Jinkela_wire_7111;
    wire new_Jinkela_wire_18984;
    wire new_Jinkela_wire_10908;
    wire new_Jinkela_wire_12908;
    wire new_Jinkela_wire_6359;
    wire _0324_;
    wire new_Jinkela_wire_13872;
    wire new_Jinkela_wire_4023;
    wire _0203_;
    wire new_Jinkela_wire_13350;
    wire new_Jinkela_wire_21179;
    wire _1703_;
    wire new_Jinkela_wire_2331;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_19677;
    wire new_Jinkela_wire_20310;
    wire new_Jinkela_wire_10193;
    wire new_Jinkela_wire_6723;
    wire new_Jinkela_wire_6825;
    wire new_Jinkela_wire_20817;
    wire new_Jinkela_wire_4620;
    wire new_Jinkela_wire_14521;
    wire new_Jinkela_wire_20586;
    wire _1835_;
    wire new_Jinkela_wire_17038;
    wire new_Jinkela_wire_20756;
    wire new_Jinkela_wire_16566;
    wire new_Jinkela_wire_10528;
    wire new_Jinkela_wire_10085;
    wire new_Jinkela_wire_2394;
    wire new_Jinkela_wire_5340;
    wire new_Jinkela_wire_16647;
    wire new_Jinkela_wire_8225;
    wire new_Jinkela_wire_16825;
    wire new_Jinkela_wire_2391;
    wire new_Jinkela_wire_9720;
    wire new_Jinkela_wire_13469;
    wire new_Jinkela_wire_3999;
    wire new_Jinkela_wire_14243;
    wire new_Jinkela_wire_10674;
    wire new_Jinkela_wire_10267;
    wire new_Jinkela_wire_20615;
    wire new_Jinkela_wire_20613;
    wire new_Jinkela_wire_17050;
    wire new_Jinkela_wire_10350;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_19902;
    wire new_Jinkela_wire_9418;
    wire new_Jinkela_wire_2676;
    wire new_Jinkela_wire_8584;
    wire new_Jinkela_wire_17754;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_18101;
    wire new_Jinkela_wire_15446;
    wire new_Jinkela_wire_14870;
    wire new_Jinkela_wire_10641;
    wire new_Jinkela_wire_6206;
    wire new_Jinkela_wire_16936;
    wire new_Jinkela_wire_19323;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_15470;
    wire new_Jinkela_wire_10693;
    wire new_Jinkela_wire_19768;
    wire new_Jinkela_wire_17325;
    wire new_Jinkela_wire_17166;
    wire new_Jinkela_wire_15355;
    wire new_Jinkela_wire_17949;
    wire new_Jinkela_wire_7823;
    wire new_Jinkela_wire_20641;
    wire new_Jinkela_wire_14195;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_16703;
    wire new_Jinkela_wire_11074;
    wire new_Jinkela_wire_19583;
    wire new_Jinkela_wire_6500;
    wire new_Jinkela_wire_17934;
    wire new_Jinkela_wire_9141;
    wire new_Jinkela_wire_19684;
    wire new_Jinkela_wire_10523;
    wire new_Jinkela_wire_11389;
    wire new_Jinkela_wire_14001;
    wire new_Jinkela_wire_14187;
    wire new_Jinkela_wire_11456;
    wire new_Jinkela_wire_10954;
    wire new_Jinkela_wire_1407;
    wire new_Jinkela_wire_7228;
    wire new_Jinkela_wire_4971;
    wire new_Jinkela_wire_11267;
    wire new_Jinkela_wire_18171;
    wire new_Jinkela_wire_9692;
    wire _1292_;
    wire new_Jinkela_wire_8766;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_16754;
    wire new_Jinkela_wire_8314;
    wire new_Jinkela_wire_18476;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_7308;
    wire new_Jinkela_wire_4011;
    wire new_Jinkela_wire_17032;
    wire new_Jinkela_wire_4645;
    wire new_Jinkela_wire_14805;
    wire new_Jinkela_wire_9838;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_15938;
    wire new_Jinkela_wire_11289;
    wire new_Jinkela_wire_20536;
    wire new_Jinkela_wire_4253;
    wire new_Jinkela_wire_6416;
    wire new_Jinkela_wire_2376;
    wire new_Jinkela_wire_18742;
    wire new_Jinkela_wire_9630;
    wire new_Jinkela_wire_18633;
    wire new_Jinkela_wire_3020;
    wire new_Jinkela_wire_17989;
    wire new_Jinkela_wire_10514;
    wire new_Jinkela_wire_3205;
    wire new_Jinkela_wire_19808;
    wire new_Jinkela_wire_15359;
    wire _1504_;
    wire new_Jinkela_wire_2760;
    wire _0487_;
    wire new_Jinkela_wire_2570;
    wire new_Jinkela_wire_18617;
    wire new_Jinkela_wire_2495;
    wire new_Jinkela_wire_13709;
    wire new_Jinkela_wire_11668;
    wire _0263_;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_17998;
    wire new_Jinkela_wire_20300;
    wire new_Jinkela_wire_9313;
    wire _1066_;
    wire new_Jinkela_wire_11396;
    wire new_Jinkela_wire_13417;
    wire new_Jinkela_wire_5643;
    wire new_Jinkela_wire_20047;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_17102;
    wire new_Jinkela_wire_14507;
    wire new_Jinkela_wire_17100;
    wire new_Jinkela_wire_17356;
    wire new_Jinkela_wire_15476;
    wire new_Jinkela_wire_11156;
    wire new_Jinkela_wire_20371;
    wire new_Jinkela_wire_10852;
    wire new_Jinkela_wire_13155;
    wire new_Jinkela_wire_20013;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_7381;
    wire _0065_;
    wire new_Jinkela_wire_12695;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_17480;
    wire new_Jinkela_wire_15577;
    wire new_Jinkela_wire_2610;
    wire new_Jinkela_wire_13317;
    wire new_Jinkela_wire_19135;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_18166;
    wire new_Jinkela_wire_6542;
    wire new_Jinkela_wire_11937;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_19771;
    wire new_Jinkela_wire_2641;
    wire new_Jinkela_wire_5893;
    wire new_Jinkela_wire_1450;
    wire new_Jinkela_wire_7854;
    wire new_Jinkela_wire_18941;
    wire new_Jinkela_wire_20296;
    wire new_Jinkela_wire_10072;
    wire new_Jinkela_wire_12025;
    wire new_Jinkela_wire_16255;
    wire new_Jinkela_wire_19081;
    wire new_Jinkela_wire_14974;
    wire new_Jinkela_wire_20672;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_2963;
    wire new_Jinkela_wire_8180;
    wire new_Jinkela_wire_11680;
    wire new_Jinkela_wire_4659;
    wire new_Jinkela_wire_2933;
    wire new_Jinkela_wire_9526;
    wire new_Jinkela_wire_5969;
    wire new_Jinkela_wire_11421;
    wire new_Jinkela_wire_20323;
    wire new_Jinkela_wire_6952;
    wire new_Jinkela_wire_5611;
    wire new_Jinkela_wire_19174;
    wire new_Jinkela_wire_3489;
    wire _1100_;
    wire new_Jinkela_wire_4993;
    wire new_Jinkela_wire_20456;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_5510;
    wire new_Jinkela_wire_12914;
    wire new_Jinkela_wire_17119;
    wire new_Jinkela_wire_9428;
    wire new_Jinkela_wire_3759;
    wire _1418_;
    wire new_Jinkela_wire_8322;
    wire _1042_;
    wire _1535_;
    wire _1660_;
    wire new_Jinkela_wire_8640;
    wire new_Jinkela_wire_7664;
    wire new_Jinkela_wire_4342;
    wire new_Jinkela_wire_16521;
    wire new_Jinkela_wire_2646;
    wire _1732_;
    wire new_Jinkela_wire_2039;
    wire _0351_;
    wire new_Jinkela_wire_9684;
    wire new_Jinkela_wire_19129;
    wire new_Jinkela_wire_11134;
    wire new_Jinkela_wire_6119;
    wire new_Jinkela_wire_3689;
    wire new_Jinkela_wire_14527;
    wire new_Jinkela_wire_11020;
    wire new_Jinkela_wire_1962;
    wire _0458_;
    wire new_Jinkela_wire_20516;
    wire new_Jinkela_wire_5988;
    wire new_Jinkela_wire_2465;
    wire new_Jinkela_wire_3390;
    wire new_Jinkela_wire_14659;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_15743;
    wire new_Jinkela_wire_12195;
    wire new_Jinkela_wire_11260;
    wire new_Jinkela_wire_10188;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_13968;
    wire _1523_;
    wire new_Jinkela_wire_19796;
    wire new_Jinkela_wire_9005;
    wire new_Jinkela_wire_4477;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_11898;
    wire new_Jinkela_wire_16917;
    wire new_Jinkela_wire_15338;
    wire new_Jinkela_wire_3963;
    wire new_Jinkela_wire_11272;
    wire new_Jinkela_wire_9977;
    wire new_Jinkela_wire_19260;
    wire new_Jinkela_wire_11905;
    wire _1513_;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_11168;
    wire _0639_;
    wire _0697_;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_14130;
    wire new_Jinkela_wire_12507;
    wire new_Jinkela_wire_18296;
    wire new_Jinkela_wire_13424;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_14612;
    wire new_Jinkela_wire_17587;
    wire new_Jinkela_wire_14909;
    wire new_Jinkela_wire_4567;
    wire new_Jinkela_wire_14210;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_2952;
    wire _0392_;
    wire new_Jinkela_wire_12822;
    wire new_Jinkela_wire_10373;
    wire _0856_;
    wire new_Jinkela_wire_4159;
    wire new_Jinkela_wire_14069;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_5972;
    wire _0590_;
    wire new_Jinkela_wire_5782;
    wire new_Jinkela_wire_18051;
    wire new_Jinkela_wire_12159;
    wire new_Jinkela_wire_3085;
    wire new_Jinkela_wire_17636;
    wire new_Jinkela_wire_2268;
    wire new_Jinkela_wire_14157;
    wire new_Jinkela_wire_20237;
    wire _1108_;
    wire new_Jinkela_wire_3147;
    wire new_Jinkela_wire_4609;
    wire new_Jinkela_wire_11012;
    wire new_Jinkela_wire_12122;
    wire new_Jinkela_wire_17208;
    wire new_Jinkela_wire_15708;
    wire new_Jinkela_wire_17922;
    wire new_Jinkela_wire_5842;
    wire new_Jinkela_wire_19690;
    wire new_Jinkela_wire_8119;
    wire new_Jinkela_wire_11837;
    wire new_Jinkela_wire_14305;
    wire _0067_;
    wire new_Jinkela_wire_10149;
    wire new_Jinkela_wire_16768;
    wire new_Jinkela_wire_18150;
    wire new_Jinkela_wire_12824;
    wire new_Jinkela_wire_15132;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_21111;
    wire new_Jinkela_wire_19452;
    wire new_Jinkela_wire_3258;
    wire new_Jinkela_wire_14273;
    wire new_Jinkela_wire_8723;
    wire new_Jinkela_wire_8726;
    wire new_Jinkela_wire_20822;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_7880;
    wire new_Jinkela_wire_16180;
    wire _0404_;
    wire new_Jinkela_wire_8254;
    wire new_Jinkela_wire_15434;
    wire new_Jinkela_wire_18809;
    wire new_Jinkela_wire_12393;
    wire new_Jinkela_wire_16584;
    wire new_Jinkela_wire_7037;
    wire new_Jinkela_wire_5374;
    wire new_Jinkela_wire_4162;
    wire new_Jinkela_wire_13023;
    wire new_Jinkela_wire_14007;
    wire new_Jinkela_wire_6180;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_1583;
    wire new_Jinkela_wire_20943;
    wire new_Jinkela_wire_8050;
    wire new_Jinkela_wire_16086;
    wire new_Jinkela_wire_2241;
    wire new_Jinkela_wire_10160;
    wire _1605_;
    wire new_Jinkela_wire_14034;
    wire new_Jinkela_wire_20709;
    wire new_Jinkela_wire_15644;
    wire new_Jinkela_wire_15384;
    wire new_Jinkela_wire_18038;
    wire new_Jinkela_wire_4406;
    wire new_Jinkela_wire_11306;
    wire new_Jinkela_wire_3645;
    wire new_Jinkela_wire_2762;
    wire new_Jinkela_wire_14569;
    wire new_Jinkela_wire_5595;
    wire new_Jinkela_wire_14513;
    wire new_Jinkela_wire_7808;
    wire new_Jinkela_wire_183;
    wire _1263_;
    wire new_Jinkela_wire_4191;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_2315;
    wire new_Jinkela_wire_9217;
    wire new_Jinkela_wire_5941;
    wire new_Jinkela_wire_12251;
    wire new_Jinkela_wire_11392;
    wire _1786_;
    wire _1471_;
    wire new_Jinkela_wire_18993;
    wire new_Jinkela_wire_18240;
    wire new_Jinkela_wire_1553;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_3375;
    wire new_Jinkela_wire_14379;
    wire new_Jinkela_wire_14312;
    wire new_Jinkela_wire_7081;
    wire new_Jinkela_wire_16432;
    wire new_Jinkela_wire_2951;
    wire new_Jinkela_wire_2703;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_13506;
    wire new_Jinkela_wire_8060;
    wire new_Jinkela_wire_17067;
    wire new_Jinkela_wire_7965;
    wire new_Jinkela_wire_17943;
    wire _1791_;
    wire _1347_;
    wire new_Jinkela_wire_3800;
    wire new_Jinkela_wire_17126;
    wire new_Jinkela_wire_16495;
    wire new_Jinkela_wire_18480;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_12773;
    wire new_Jinkela_wire_19679;
    wire new_Jinkela_wire_17134;
    wire new_Jinkela_wire_18590;
    wire new_Jinkela_wire_9661;
    wire new_Jinkela_wire_6758;
    wire new_Jinkela_wire_13116;
    wire new_Jinkela_wire_19726;
    wire new_Jinkela_wire_18957;
    wire new_Jinkela_wire_21147;
    wire new_Jinkela_wire_12253;
    wire new_Jinkela_wire_11532;
    wire new_Jinkela_wire_4090;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_15396;
    wire new_Jinkela_wire_241;
    wire _1129_;
    wire new_Jinkela_wire_13590;
    wire new_Jinkela_wire_14992;
    wire new_Jinkela_wire_17026;
    wire new_Jinkela_wire_11006;
    wire new_Jinkela_wire_8020;
    wire _1279_;
    wire new_Jinkela_wire_13222;
    wire new_Jinkela_wire_15151;
    wire new_Jinkela_wire_3749;
    wire new_Jinkela_wire_8126;
    wire _0881_;
    wire new_Jinkela_wire_19947;
    wire new_Jinkela_wire_15117;
    wire new_Jinkela_wire_17383;
    wire new_Jinkela_wire_8309;
    wire _0666_;
    wire new_Jinkela_wire_19366;
    wire new_Jinkela_wire_1503;
    wire new_Jinkela_wire_10436;
    wire new_Jinkela_wire_4105;
    wire new_Jinkela_wire_18153;
    wire new_Jinkela_wire_9760;
    wire new_Jinkela_wire_17912;
    wire new_Jinkela_wire_16176;
    wire new_Jinkela_wire_11838;
    wire new_Jinkela_wire_10097;
    wire new_Jinkela_wire_3203;
    wire new_Jinkela_wire_15473;
    wire new_Jinkela_wire_13594;
    wire new_Jinkela_wire_6240;
    wire new_Jinkela_wire_17517;
    wire _0348_;
    wire _1233_;
    wire new_Jinkela_wire_2262;
    wire new_Jinkela_wire_2073;
    wire new_Jinkela_wire_13024;
    wire _0634_;
    wire new_Jinkela_wire_14054;
    wire new_Jinkela_wire_5480;
    wire new_Jinkela_wire_2695;
    wire new_Jinkela_wire_13687;
    wire new_Jinkela_wire_16736;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_9878;
    wire new_Jinkela_wire_17927;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_2658;
    wire new_Jinkela_wire_7877;
    wire new_Jinkela_wire_9221;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_3979;
    wire new_Jinkela_wire_4743;
    wire new_Jinkela_wire_5489;
    wire new_Jinkela_wire_13422;
    wire new_Jinkela_wire_19650;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_15700;
    wire new_Jinkela_wire_2400;
    wire new_Jinkela_wire_4454;
    wire new_Jinkela_wire_1979;
    wire new_Jinkela_wire_19779;
    wire new_Jinkela_wire_2420;
    wire new_Jinkela_wire_14236;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_18405;
    wire new_Jinkela_wire_5722;
    wire new_Jinkela_wire_13340;
    wire new_Jinkela_wire_3135;
    wire new_Jinkela_wire_18906;
    wire new_Jinkela_wire_3826;
    wire new_Jinkela_wire_4860;
    wire new_Jinkela_wire_20916;
    wire new_Jinkela_wire_19035;
    wire new_Jinkela_wire_2119;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_4781;
    wire new_Jinkela_wire_5493;
    wire new_Jinkela_wire_7670;
    wire new_Jinkela_wire_5323;
    wire new_Jinkela_wire_3579;
    wire _1078_;
    wire new_Jinkela_wire_4027;
    wire new_Jinkela_wire_19575;
    wire new_Jinkela_wire_14554;
    wire new_Jinkela_wire_8749;
    wire new_Jinkela_wire_9548;
    wire new_Jinkela_wire_10850;
    wire new_net_3946;
    wire _0726_;
    wire new_Jinkela_wire_7632;
    wire new_Jinkela_wire_11255;
    wire new_Jinkela_wire_8447;
    wire _1003_;
    wire new_Jinkela_wire_8515;
    wire new_Jinkela_wire_14831;
    wire new_Jinkela_wire_3427;
    wire new_Jinkela_wire_18312;
    wire new_Jinkela_wire_10953;
    wire new_Jinkela_wire_18378;
    wire new_Jinkela_wire_13855;
    wire new_Jinkela_wire_3975;
    wire new_Jinkela_wire_15594;
    wire new_Jinkela_wire_5198;
    wire new_Jinkela_wire_20492;
    wire new_Jinkela_wire_10343;
    wire new_Jinkela_wire_17519;
    wire new_Jinkela_wire_9514;
    wire _1381_;
    wire new_Jinkela_wire_10677;
    wire new_Jinkela_wire_4397;
    wire new_Jinkela_wire_16101;
    wire new_Jinkela_wire_9111;
    wire new_Jinkela_wire_13143;
    wire new_Jinkela_wire_8540;
    wire new_Jinkela_wire_20070;
    wire new_Jinkela_wire_14352;
    wire new_Jinkela_wire_7583;
    wire new_Jinkela_wire_5836;
    wire new_Jinkela_wire_11394;
    wire new_Jinkela_wire_14140;
    wire new_Jinkela_wire_16361;
    wire new_Jinkela_wire_13097;
    wire new_Jinkela_wire_4052;
    wire new_Jinkela_wire_14738;
    wire _0200_;
    wire _0773_;
    wire new_Jinkela_wire_15262;
    wire new_Jinkela_wire_18183;
    wire new_Jinkela_wire_1421;
    wire new_Jinkela_wire_10978;
    wire new_Jinkela_wire_8877;
    wire new_Jinkela_wire_16856;
    wire new_Jinkela_wire_9078;
    wire new_Jinkela_wire_12582;
    wire new_Jinkela_wire_6365;
    wire new_Jinkela_wire_2064;
    wire new_Jinkela_wire_14663;
    wire new_Jinkela_wire_11830;
    wire new_Jinkela_wire_13090;
    wire new_Jinkela_wire_4473;
    wire new_Jinkela_wire_3473;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_12755;
    wire new_Jinkela_wire_15998;
    wire new_Jinkela_wire_8636;
    wire new_Jinkela_wire_13972;
    wire new_Jinkela_wire_19434;
    wire new_Jinkela_wire_4145;
    wire new_Jinkela_wire_17122;
    wire new_Jinkela_wire_7239;
    wire new_Jinkela_wire_18645;
    wire new_Jinkela_wire_2586;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_8734;
    wire new_Jinkela_wire_10938;
    wire new_Jinkela_wire_6445;
    wire new_Jinkela_wire_14397;
    wire new_Jinkela_wire_10974;
    wire new_Jinkela_wire_4505;
    wire new_Jinkela_wire_5739;
    wire new_Jinkela_wire_18059;
    wire new_Jinkela_wire_3544;
    wire new_Jinkela_wire_14785;
    wire new_Jinkela_wire_13187;
    wire new_Jinkela_wire_18836;
    wire new_Jinkela_wire_19077;
    wire new_Jinkela_wire_8159;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_12498;
    wire new_Jinkela_wire_3335;
    wire new_Jinkela_wire_16938;
    wire new_Jinkela_wire_2544;
    wire new_Jinkela_wire_3223;
    wire _0717_;
    wire new_Jinkela_wire_15657;
    wire new_Jinkela_wire_5982;
    wire new_Jinkela_wire_19361;
    wire _1342_;
    wire new_Jinkela_wire_10917;
    wire new_Jinkela_wire_16358;
    wire new_Jinkela_wire_1739;
    wire new_Jinkela_wire_8667;
    wire new_Jinkela_wire_13068;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_21056;
    wire new_Jinkela_wire_16940;
    wire new_Jinkela_wire_4626;
    wire new_Jinkela_wire_19623;
    wire new_Jinkela_wire_9857;
    wire new_Jinkela_wire_9956;
    wire new_Jinkela_wire_17866;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_17160;
    wire new_Jinkela_wire_3055;
    wire new_Jinkela_wire_14773;
    wire new_Jinkela_wire_16298;
    wire new_Jinkela_wire_2076;
    wire new_Jinkela_wire_17857;
    wire new_Jinkela_wire_10083;
    wire new_Jinkela_wire_15404;
    wire new_Jinkela_wire_15968;
    wire new_Jinkela_wire_15850;
    wire new_Jinkela_wire_2510;
    wire new_Jinkela_wire_18070;
    wire new_Jinkela_wire_19109;
    wire _1558_;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_1764;
    wire new_Jinkela_wire_4110;
    wire new_Jinkela_wire_15536;
    wire new_Jinkela_wire_11694;
    wire new_Jinkela_wire_16404;
    wire new_Jinkela_wire_10783;
    wire new_Jinkela_wire_13154;
    wire _0427_;
    wire new_Jinkela_wire_19381;
    wire new_Jinkela_wire_10057;
    wire new_Jinkela_wire_19945;
    wire new_Jinkela_wire_17386;
    wire new_Jinkela_wire_7738;
    wire new_Jinkela_wire_8042;
    wire new_Jinkela_wire_1260;
    wire _0019_;
    wire new_Jinkela_wire_11201;
    wire new_Jinkela_wire_17136;
    wire new_Jinkela_wire_10802;
    wire new_Jinkela_wire_6701;
    wire new_Jinkela_wire_19807;
    wire new_Jinkela_wire_6844;
    wire new_Jinkela_wire_4078;
    wire new_Jinkela_wire_11571;
    wire new_Jinkela_wire_12147;
    wire new_Jinkela_wire_13293;
    wire new_Jinkela_wire_8432;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_10269;
    wire new_Jinkela_wire_16460;
    wire new_Jinkela_wire_18154;
    wire _0631_;
    wire new_Jinkela_wire_8559;
    wire new_Jinkela_wire_19020;
    wire _1615_;
    wire new_Jinkela_wire_7905;
    wire new_Jinkela_wire_10216;
    wire _0475_;
    wire new_Jinkela_wire_3870;
    wire new_Jinkela_wire_14455;
    wire new_Jinkela_wire_15781;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_3257;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_15269;
    wire new_Jinkela_wire_4468;
    wire new_Jinkela_wire_13647;
    wire new_Jinkela_wire_7800;
    wire new_Jinkela_wire_12489;
    wire new_Jinkela_wire_20802;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_20600;
    wire new_Jinkela_wire_13342;
    wire new_Jinkela_wire_14895;
    wire new_Jinkela_wire_20920;
    wire new_Jinkela_wire_5818;
    wire new_Jinkela_wire_15862;
    wire _0688_;
    wire new_Jinkela_wire_8711;
    wire new_Jinkela_wire_13037;
    wire new_Jinkela_wire_10864;
    wire new_Jinkela_wire_3396;
    wire new_Jinkela_wire_16295;
    wire new_Jinkela_wire_5277;
    wire new_Jinkela_wire_3626;
    wire new_Jinkela_wire_11082;
    wire new_Jinkela_wire_15086;
    wire new_Jinkela_wire_18639;
    wire new_Jinkela_wire_7226;
    wire new_Jinkela_wire_14414;
    wire new_Jinkela_wire_11740;
    wire new_Jinkela_wire_16292;
    wire new_Jinkela_wire_14783;
    wire new_Jinkela_wire_18811;
    wire new_Jinkela_wire_6897;
    wire new_Jinkela_wire_5769;
    wire new_Jinkela_wire_14278;
    wire new_Jinkela_wire_8176;
    wire new_Jinkela_wire_4780;
    wire _0833_;
    wire new_Jinkela_wire_18782;
    wire new_Jinkela_wire_4208;
    wire new_Jinkela_wire_6790;
    wire new_Jinkela_wire_9024;
    wire new_Jinkela_wire_14418;
    wire new_Jinkela_wire_17937;
    wire new_Jinkela_wire_21118;
    wire new_Jinkela_wire_20163;
    wire new_Jinkela_wire_18708;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_21306;
    wire new_Jinkela_wire_5538;
    wire new_Jinkela_wire_2847;
    wire new_Jinkela_wire_15307;
    wire new_Jinkela_wire_12658;
    wire new_Jinkela_wire_13128;
    wire new_Jinkela_wire_20340;
    wire new_Jinkela_wire_4003;
    wire _0783_;
    wire new_Jinkela_wire_4069;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_9504;
    wire new_Jinkela_wire_6797;
    wire new_Jinkela_wire_16539;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_12142;
    wire new_Jinkela_wire_12727;
    wire new_Jinkela_wire_2992;
    wire new_Jinkela_wire_19370;
    wire new_Jinkela_wire_18889;
    wire new_Jinkela_wire_15112;
    wire new_Jinkela_wire_3208;
    wire new_Jinkela_wire_8598;
    wire new_Jinkela_wire_2988;
    wire new_Jinkela_wire_21278;
    wire new_Jinkela_wire_18997;
    wire new_Jinkela_wire_13192;
    wire new_Jinkela_wire_20494;
    wire new_Jinkela_wire_6018;
    wire new_Jinkela_wire_4528;
    wire new_Jinkela_wire_13329;
    wire new_Jinkela_wire_10497;
    wire new_Jinkela_wire_5666;
    wire new_Jinkela_wire_5557;
    wire _0985_;
    wire new_Jinkela_wire_17276;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_20980;
    wire new_Jinkela_wire_6628;
    wire new_Jinkela_wire_13078;
    wire new_Jinkela_wire_11195;
    wire new_Jinkela_wire_17363;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_3328;
    wire new_Jinkela_wire_20732;
    wire new_Jinkela_wire_13163;
    wire new_Jinkela_wire_10717;
    wire new_Jinkela_wire_7429;
    wire new_Jinkela_wire_20717;
    wire new_Jinkela_wire_9756;
    wire _1345_;
    wire new_Jinkela_wire_10122;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_16239;
    wire new_Jinkela_wire_9301;
    wire new_Jinkela_wire_15780;
    wire new_Jinkela_wire_17197;
    wire new_Jinkela_wire_5284;
    wire new_Jinkela_wire_4245;
    wire new_Jinkela_wire_6140;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_15959;
    wire new_Jinkela_wire_4644;
    wire new_Jinkela_wire_19619;
    wire new_Jinkela_wire_6939;
    wire new_Jinkela_wire_1688;
    wire new_Jinkela_wire_8956;
    wire _1742_;
    wire new_Jinkela_wire_4822;
    wire new_Jinkela_wire_12478;
    wire new_Jinkela_wire_12750;
    wire _1718_;
    wire new_Jinkela_wire_10491;
    wire new_Jinkela_wire_14947;
    wire new_Jinkela_wire_1857;
    wire _0954_;
    wire new_Jinkela_wire_7801;
    wire new_Jinkela_wire_2593;
    wire _0130_;
    wire new_Jinkela_wire_2475;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_17190;
    wire new_Jinkela_wire_12508;
    wire _0582_;
    wire new_Jinkela_wire_5218;
    wire new_Jinkela_wire_16811;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_19757;
    wire new_Jinkela_wire_9731;
    wire new_Jinkela_wire_4992;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_13184;
    wire new_Jinkela_wire_20585;
    wire new_Jinkela_wire_12396;
    wire new_Jinkela_wire_20054;
    wire new_Jinkela_wire_1754;
    wire new_Jinkela_wire_13439;
    wire new_Jinkela_wire_12048;
    wire new_Jinkela_wire_11145;
    wire new_Jinkela_wire_6069;
    wire new_Jinkela_wire_6923;
    wire new_Jinkela_wire_11639;
    wire new_Jinkela_wire_4271;
    wire new_Jinkela_wire_3287;
    wire new_Jinkela_wire_13628;
    wire new_Jinkela_wire_9535;
    wire _1761_;
    wire _0168_;
    wire _1000_;
    wire new_Jinkela_wire_19365;
    wire new_Jinkela_wire_16090;
    wire new_Jinkela_wire_16945;
    wire new_Jinkela_wire_8480;
    wire new_Jinkela_wire_6061;
    wire new_Jinkela_wire_9325;
    wire new_Jinkela_wire_13918;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_19352;
    wire new_Jinkela_wire_9965;
    wire new_Jinkela_wire_1728;
    wire new_Jinkela_wire_9236;
    wire new_Jinkela_wire_3076;
    wire new_Jinkela_wire_9808;
    wire new_Jinkela_wire_14883;
    wire new_Jinkela_wire_7666;
    wire new_Jinkela_wire_5616;
    wire _0772_;
    wire new_Jinkela_wire_6631;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_20838;
    wire new_Jinkela_wire_2503;
    wire new_Jinkela_wire_1333;
    wire new_Jinkela_wire_7044;
    wire _0637_;
    wire new_Jinkela_wire_18450;
    wire new_Jinkela_wire_11089;
    wire new_Jinkela_wire_10878;
    wire new_Jinkela_wire_3383;
    wire new_Jinkela_wire_19172;
    wire new_Jinkela_wire_7648;
    wire new_Jinkela_wire_14044;
    wire new_Jinkela_wire_6499;
    wire new_Jinkela_wire_7363;
    wire new_Jinkela_wire_13324;
    wire new_Jinkela_wire_21228;
    wire new_Jinkela_wire_12108;
    wire new_Jinkela_wire_20999;
    wire new_Jinkela_wire_11280;
    wire new_Jinkela_wire_11757;
    wire _0989_;
    wire new_Jinkela_wire_14582;
    wire _1149_;
    wire new_Jinkela_wire_16422;
    wire new_Jinkela_wire_3439;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_13562;
    wire new_Jinkela_wire_16857;
    wire new_Jinkela_wire_2552;
    wire new_Jinkela_wire_20825;
    wire new_Jinkela_wire_1327;
    wire _0609_;
    wire new_Jinkela_wire_13274;
    wire new_Jinkela_wire_13585;
    wire new_Jinkela_wire_21290;
    wire new_Jinkela_wire_3869;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_18157;
    wire new_Jinkela_wire_8681;
    wire new_Jinkela_wire_12223;
    wire new_Jinkela_wire_5445;
    wire _0361_;
    wire new_Jinkela_wire_12803;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_12325;
    wire new_Jinkela_wire_7917;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_3858;
    wire new_Jinkela_wire_11930;
    wire new_Jinkela_wire_12918;
    wire new_Jinkela_wire_12706;
    wire new_Jinkela_wire_11527;
    wire new_Jinkela_wire_3070;
    wire _0903_;
    wire _1776_;
    wire new_Jinkela_wire_11736;
    wire new_Jinkela_wire_4316;
    wire new_Jinkela_wire_11200;
    wire _0321_;
    wire new_Jinkela_wire_10991;
    wire new_Jinkela_wire_8613;
    wire new_Jinkela_wire_13699;
    wire _0123_;
    wire new_Jinkela_wire_13836;
    wire new_Jinkela_wire_21271;
    wire new_Jinkela_wire_9894;
    wire new_Jinkela_wire_8543;
    wire new_Jinkela_wire_15799;
    wire new_Jinkela_wire_18938;
    wire new_Jinkela_wire_16105;
    wire new_Jinkela_wire_9263;
    wire new_Jinkela_wire_10040;
    wire new_Jinkela_wire_5399;
    wire new_Jinkela_wire_8550;
    wire new_Jinkela_wire_12047;
    wire new_Jinkela_wire_13328;
    wire new_Jinkela_wire_6088;
    wire new_Jinkela_wire_13237;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_19914;
    wire new_Jinkela_wire_7953;
    wire new_Jinkela_wire_16922;
    wire _0276_;
    wire new_Jinkela_wire_5246;
    wire new_Jinkela_wire_5863;
    wire new_Jinkela_wire_14415;
    wire new_Jinkela_wire_15430;
    wire new_Jinkela_wire_14670;
    wire new_Jinkela_wire_2839;
    wire new_Jinkela_wire_9578;
    wire new_Jinkela_wire_17092;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_15238;
    wire new_Jinkela_wire_15173;
    wire new_Jinkela_wire_15912;
    wire new_Jinkela_wire_3614;
    wire new_Jinkela_wire_4719;
    wire new_Jinkela_wire_11099;
    wire new_Jinkela_wire_19243;
    wire new_Jinkela_wire_9639;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_15219;
    wire new_Jinkela_wire_2350;
    wire _1061_;
    wire new_Jinkela_wire_20445;
    wire new_Jinkela_wire_11080;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_15990;
    wire _1433_;
    wire _0320_;
    wire new_Jinkela_wire_2329;
    wire new_Jinkela_wire_2460;
    wire new_Jinkela_wire_20057;
    wire new_Jinkela_wire_11901;
    wire new_Jinkela_wire_14112;
    wire new_Jinkela_wire_2097;
    wire _0357_;
    wire new_Jinkela_wire_12527;
    wire new_Jinkela_wire_3588;
    wire new_Jinkela_wire_20035;
    wire new_Jinkela_wire_14750;
    wire new_Jinkela_wire_18800;
    wire new_Jinkela_wire_9219;
    wire new_Jinkela_wire_6829;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_9196;
    wire new_Jinkela_wire_20140;
    wire new_Jinkela_wire_12468;
    wire new_Jinkela_wire_3799;
    wire new_Jinkela_wire_7076;
    wire new_Jinkela_wire_19302;
    wire new_Jinkela_wire_3364;
    wire new_Jinkela_wire_13919;
    wire new_Jinkela_wire_16119;
    wire new_Jinkela_wire_1652;
    wire _0840_;
    wire new_Jinkela_wire_2929;
    wire new_Jinkela_wire_13801;
    wire new_Jinkela_wire_10289;
    wire new_Jinkela_wire_20174;
    wire new_Jinkela_wire_21091;
    wire new_Jinkela_wire_18628;
    wire new_Jinkela_wire_18980;
    wire new_Jinkela_wire_13084;
    wire new_Jinkela_wire_3488;
    wire new_Jinkela_wire_19840;
    wire _0001_;
    wire new_Jinkela_wire_20223;
    wire new_Jinkela_wire_4131;
    wire new_Jinkela_wire_13019;
    wire new_Jinkela_wire_16654;
    wire new_Jinkela_wire_10009;
    wire new_Jinkela_wire_18949;
    wire new_Jinkela_wire_8567;
    wire _0673_;
    wire new_Jinkela_wire_10643;
    wire _0496_;
    wire new_Jinkela_wire_3126;
    wire new_Jinkela_wire_4428;
    wire _0336_;
    wire new_Jinkela_wire_2685;
    wire _1712_;
    wire new_Jinkela_wire_9202;
    wire new_Jinkela_wire_17108;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_3317;
    wire new_Jinkela_wire_13170;
    wire new_Jinkela_wire_4508;
    wire new_Jinkela_wire_18422;
    wire _0916_;
    wire new_Jinkela_wire_7067;
    wire new_Jinkela_wire_4395;
    wire new_Jinkela_wire_6581;
    wire new_Jinkela_wire_9715;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_10699;
    wire new_Jinkela_wire_16424;
    wire new_Jinkela_wire_15231;
    wire new_Jinkela_wire_4237;
    wire _0796_;
    wire new_Jinkela_wire_5226;
    wire new_Jinkela_wire_20683;
    wire new_Jinkela_wire_6815;
    wire new_Jinkela_wire_2108;
    wire new_Jinkela_wire_18335;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_1954;
    wire new_Jinkela_wire_9017;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_13689;
    wire new_Jinkela_wire_3060;
    wire new_Jinkela_wire_2415;
    wire new_Jinkela_wire_6837;
    wire _0970_;
    wire new_Jinkela_wire_20885;
    wire new_Jinkela_wire_20149;
    wire new_Jinkela_wire_9135;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_2627;
    wire new_Jinkela_wire_4988;
    wire new_Jinkela_wire_2194;
    wire new_Jinkela_wire_9419;
    wire new_Jinkela_wire_15026;
    wire new_Jinkela_wire_4869;
    wire new_Jinkela_wire_20197;
    wire new_Jinkela_wire_4259;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_9554;
    wire new_Jinkela_wire_20784;
    wire new_Jinkela_wire_1085;
    wire _1631_;
    wire new_Jinkela_wire_15638;
    wire new_Jinkela_wire_10729;
    wire _1265_;
    wire new_Jinkela_wire_12961;
    wire new_Jinkela_wire_19850;
    wire new_Jinkela_wire_19203;
    wire new_Jinkela_wire_14699;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_9092;
    wire new_Jinkela_wire_20334;
    wire new_Jinkela_wire_19426;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_4534;
    wire new_Jinkela_wire_17413;
    wire new_Jinkela_wire_6247;
    wire new_Jinkela_wire_2474;
    wire new_Jinkela_wire_18569;
    wire new_Jinkela_wire_8612;
    wire new_Jinkela_wire_17449;
    wire new_Jinkela_wire_3731;
    wire new_Jinkela_wire_16388;
    wire new_Jinkela_wire_8063;
    wire new_Jinkela_wire_11407;
    wire _1505_;
    wire new_Jinkela_wire_2840;
    wire new_Jinkela_wire_11732;
    wire new_Jinkela_wire_15411;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_17034;
    wire new_Jinkela_wire_8127;
    wire new_Jinkela_wire_14821;
    wire _1198_;
    wire new_Jinkela_wire_7956;
    wire new_Jinkela_wire_10990;
    wire new_Jinkela_wire_18496;
    wire new_Jinkela_wire_14691;
    wire new_Jinkela_wire_8232;
    wire new_Jinkela_wire_20960;
    wire new_Jinkela_wire_13529;
    wire new_Jinkela_wire_7082;
    wire new_Jinkela_wire_9742;
    wire new_Jinkela_wire_10670;
    wire new_Jinkela_wire_14060;
    wire new_Jinkela_wire_975;
    wire _1300_;
    wire new_Jinkela_wire_3207;
    wire new_Jinkela_wire_5050;
    wire new_Jinkela_wire_19812;
    wire new_Jinkela_wire_16517;
    wire new_Jinkela_wire_1003;
    wire _1484_;
    wire new_Jinkela_wire_5704;
    wire new_Jinkela_wire_7166;
    wire new_Jinkela_wire_12798;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_15405;
    wire new_Jinkela_wire_10972;
    wire _0806_;
    wire new_Jinkela_wire_17697;
    wire new_Jinkela_wire_11956;
    wire new_Jinkela_wire_7249;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_4516;
    wire new_Jinkela_wire_4643;
    wire new_Jinkela_wire_5862;
    wire new_Jinkela_wire_4028;
    wire new_Jinkela_wire_16919;
    wire new_Jinkela_wire_16942;
    wire new_Jinkela_wire_18134;
    wire new_Jinkela_wire_20891;
    wire new_Jinkela_wire_12832;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_8818;
    wire new_Jinkela_wire_3849;
    wire new_Jinkela_wire_20073;
    wire new_Jinkela_wire_20776;
    wire new_Jinkela_wire_12363;
    wire new_Jinkela_wire_4984;
    wire new_Jinkela_wire_10696;
    wire new_Jinkela_wire_12751;
    wire new_Jinkela_wire_6436;
    wire new_Jinkela_wire_17154;
    wire new_Jinkela_wire_2286;
    wire new_Jinkela_wire_7026;
    wire new_Jinkela_wire_20235;
    wire new_Jinkela_wire_2877;
    wire new_Jinkela_wire_2157;
    wire new_Jinkela_wire_9178;
    wire new_Jinkela_wire_16589;
    wire new_Jinkela_wire_3164;
    wire new_Jinkela_wire_20893;
    wire new_Jinkela_wire_11030;
    wire _0396_;
    wire new_Jinkela_wire_17566;
    wire new_Jinkela_wire_381;
    wire _0300_;
    wire _1045_;
    wire new_Jinkela_wire_8244;
    wire new_Jinkela_wire_5446;
    wire new_Jinkela_wire_15119;
    wire new_Jinkela_wire_1332;
    wire _0154_;
    wire new_Jinkela_wire_12565;
    wire new_Jinkela_wire_3532;
    wire new_Jinkela_wire_13549;
    wire new_Jinkela_wire_18989;
    wire new_Jinkela_wire_4488;
    wire new_Jinkela_wire_11569;
    wire new_Jinkela_wire_19642;
    wire new_Jinkela_wire_4132;
    wire new_Jinkela_wire_20024;
    wire new_Jinkela_wire_6768;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_12442;
    wire new_Jinkela_wire_5279;
    wire new_Jinkela_wire_13244;
    wire _1429_;
    wire new_Jinkela_wire_4453;
    wire new_Jinkela_wire_14834;
    wire new_Jinkela_wire_13045;
    wire new_Jinkela_wire_18834;
    wire new_Jinkela_wire_5263;
    wire new_Jinkela_wire_12623;
    wire new_Jinkela_wire_11728;
    wire new_Jinkela_wire_17617;
    wire new_Jinkela_wire_21216;
    wire new_Jinkela_wire_14510;
    wire new_Jinkela_wire_7389;
    wire _1337_;
    wire new_Jinkela_wire_13016;
    wire new_Jinkela_wire_18666;
    wire new_Jinkela_wire_4763;
    wire new_Jinkela_wire_3694;
    wire _1204_;
    wire new_Jinkela_wire_21169;
    wire new_Jinkela_wire_2100;
    wire new_Jinkela_wire_21263;
    wire new_Jinkela_wire_2383;
    wire new_Jinkela_wire_10002;
    wire new_Jinkela_wire_13051;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_7095;
    wire new_Jinkela_wire_20870;
    wire new_Jinkela_wire_7866;
    wire _0668_;
    wire _0086_;
    wire new_Jinkela_wire_7122;
    wire new_Jinkela_wire_18709;
    wire new_Jinkela_wire_16983;
    wire new_Jinkela_wire_15819;
    wire new_Jinkela_wire_8035;
    wire new_Jinkela_wire_13552;
    wire new_Jinkela_wire_10203;
    wire new_Jinkela_wire_10143;
    wire new_Jinkela_wire_17782;
    wire new_Jinkela_wire_16951;
    wire new_Jinkela_wire_14859;
    wire new_Jinkela_wire_19617;
    wire new_Jinkela_wire_16147;
    wire new_Jinkela_wire_5282;
    wire new_Jinkela_wire_5240;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_20814;
    wire new_Jinkela_wire_14370;
    wire new_Jinkela_wire_7019;
    wire new_Jinkela_wire_8952;
    wire new_Jinkela_wire_2053;
    wire new_Jinkela_wire_15319;
    wire new_Jinkela_wire_16676;
    wire new_Jinkela_wire_15744;
    wire _1566_;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_14302;
    wire _0316_;
    wire new_Jinkela_wire_21168;
    wire new_Jinkela_wire_4430;
    wire new_Jinkela_wire_1404;
    wire new_Jinkela_wire_19001;
    wire new_Jinkela_wire_16331;
    input N426;
    input N154;
    input N358;
    input N69;
    input N18;
    input N443;
    input N494;
    input N222;
    input N171;
    input N477;
    input N273;
    input N392;
    input N52;
    input N375;
    input N290;
    input N1;
    input N103;
    input N188;
    input N205;
    input N256;
    input N409;
    input N86;
    input N137;
    input N511;
    input N307;
    input N35;
    input N460;
    input N239;
    input N324;
    input N341;
    input N528;
    input N120;
    output N6200;
    output N6280;
    output N6210;
    output N1581;
    output N6270;
    output N6260;
    output N2548;
    output N4946;
    output N5308;
    output N6250;
    output N6220;
    output N5971;
    output N6170;
    output N3552;
    output N6288;
    output N4591;
    output N6240;
    output N6150;
    output N545;
    output N6123;
    output N6180;
    output N6160;
    output N2877;
    output N2223;
    output N3895;
    output N6287;
    output N6190;
    output N5672;
    output N3211;
    output N1901;
    output N6230;
    output N4241;

    bfr new_Jinkela_buffer_10551 (
        .din(new_Jinkela_wire_12750),
        .dout(new_Jinkela_wire_12751)
    );

    bfr new_Jinkela_buffer_10492 (
        .din(new_Jinkela_wire_12669),
        .dout(new_Jinkela_wire_12670)
    );

    bfr new_Jinkela_buffer_10634 (
        .din(new_Jinkela_wire_12835),
        .dout(new_Jinkela_wire_12836)
    );

    bfr new_Jinkela_buffer_10493 (
        .din(new_Jinkela_wire_12670),
        .dout(new_Jinkela_wire_12671)
    );

    bfr new_Jinkela_buffer_10552 (
        .din(new_Jinkela_wire_12751),
        .dout(new_Jinkela_wire_12752)
    );

    bfr new_Jinkela_buffer_10494 (
        .din(new_Jinkela_wire_12671),
        .dout(new_Jinkela_wire_12672)
    );

    bfr new_Jinkela_buffer_10703 (
        .din(new_Jinkela_wire_12908),
        .dout(new_Jinkela_wire_12909)
    );

    bfr new_Jinkela_buffer_10495 (
        .din(new_Jinkela_wire_12672),
        .dout(new_Jinkela_wire_12673)
    );

    bfr new_Jinkela_buffer_10553 (
        .din(new_Jinkela_wire_12752),
        .dout(new_Jinkela_wire_12753)
    );

    bfr new_Jinkela_buffer_10496 (
        .din(new_Jinkela_wire_12673),
        .dout(new_Jinkela_wire_12674)
    );

    bfr new_Jinkela_buffer_10635 (
        .din(new_Jinkela_wire_12836),
        .dout(new_Jinkela_wire_12837)
    );

    bfr new_Jinkela_buffer_10497 (
        .din(new_Jinkela_wire_12674),
        .dout(new_Jinkela_wire_12675)
    );

    bfr new_Jinkela_buffer_10554 (
        .din(new_Jinkela_wire_12753),
        .dout(new_Jinkela_wire_12754)
    );

    bfr new_Jinkela_buffer_10498 (
        .din(new_Jinkela_wire_12675),
        .dout(new_Jinkela_wire_12676)
    );

    spl2 new_Jinkela_splitter_954 (
        .a(_1737_),
        .b(new_Jinkela_wire_13012),
        .c(new_Jinkela_wire_13013)
    );

    bfr new_Jinkela_buffer_10499 (
        .din(new_Jinkela_wire_12676),
        .dout(new_Jinkela_wire_12677)
    );

    bfr new_Jinkela_buffer_10555 (
        .din(new_Jinkela_wire_12754),
        .dout(new_Jinkela_wire_12755)
    );

    bfr new_Jinkela_buffer_10500 (
        .din(new_Jinkela_wire_12677),
        .dout(new_Jinkela_wire_12678)
    );

    bfr new_Jinkela_buffer_10636 (
        .din(new_Jinkela_wire_12837),
        .dout(new_Jinkela_wire_12838)
    );

    bfr new_Jinkela_buffer_10501 (
        .din(new_Jinkela_wire_12678),
        .dout(new_Jinkela_wire_12679)
    );

    bfr new_Jinkela_buffer_10556 (
        .din(new_Jinkela_wire_12755),
        .dout(new_Jinkela_wire_12756)
    );

    bfr new_Jinkela_buffer_10502 (
        .din(new_Jinkela_wire_12679),
        .dout(new_Jinkela_wire_12680)
    );

    bfr new_Jinkela_buffer_10704 (
        .din(new_Jinkela_wire_12909),
        .dout(new_Jinkela_wire_12910)
    );

    bfr new_Jinkela_buffer_10503 (
        .din(new_Jinkela_wire_12680),
        .dout(new_Jinkela_wire_12681)
    );

    bfr new_Jinkela_buffer_10557 (
        .din(new_Jinkela_wire_12756),
        .dout(new_Jinkela_wire_12757)
    );

    bfr new_Jinkela_buffer_10504 (
        .din(new_Jinkela_wire_12681),
        .dout(new_Jinkela_wire_12682)
    );

    bfr new_Jinkela_buffer_10637 (
        .din(new_Jinkela_wire_12838),
        .dout(new_Jinkela_wire_12839)
    );

    bfr new_Jinkela_buffer_10505 (
        .din(new_Jinkela_wire_12682),
        .dout(new_Jinkela_wire_12683)
    );

    bfr new_Jinkela_buffer_10558 (
        .din(new_Jinkela_wire_12757),
        .dout(new_Jinkela_wire_12758)
    );

    bfr new_Jinkela_buffer_10506 (
        .din(new_Jinkela_wire_12683),
        .dout(new_Jinkela_wire_12684)
    );

    bfr new_Jinkela_buffer_10802 (
        .din(_1415_),
        .dout(new_Jinkela_wire_13014)
    );

    bfr new_Jinkela_buffer_10507 (
        .din(new_Jinkela_wire_12684),
        .dout(new_Jinkela_wire_12685)
    );

    bfr new_Jinkela_buffer_10559 (
        .din(new_Jinkela_wire_12758),
        .dout(new_Jinkela_wire_12759)
    );

    bfr new_Jinkela_buffer_10508 (
        .din(new_Jinkela_wire_12685),
        .dout(new_Jinkela_wire_12686)
    );

    bfr new_Jinkela_buffer_10638 (
        .din(new_Jinkela_wire_12839),
        .dout(new_Jinkela_wire_12840)
    );

    bfr new_Jinkela_buffer_10509 (
        .din(new_Jinkela_wire_12686),
        .dout(new_Jinkela_wire_12687)
    );

    bfr new_Jinkela_buffer_10560 (
        .din(new_Jinkela_wire_12759),
        .dout(new_Jinkela_wire_12760)
    );

    bfr new_Jinkela_buffer_10510 (
        .din(new_Jinkela_wire_12687),
        .dout(new_Jinkela_wire_12688)
    );

    bfr new_Jinkela_buffer_10705 (
        .din(new_Jinkela_wire_12910),
        .dout(new_Jinkela_wire_12911)
    );

    bfr new_Jinkela_buffer_10511 (
        .din(new_Jinkela_wire_12688),
        .dout(new_Jinkela_wire_12689)
    );

    bfr new_Jinkela_buffer_10561 (
        .din(new_Jinkela_wire_12760),
        .dout(new_Jinkela_wire_12761)
    );

    bfr new_Jinkela_buffer_10512 (
        .din(new_Jinkela_wire_12689),
        .dout(new_Jinkela_wire_12690)
    );

    bfr new_Jinkela_buffer_17471 (
        .din(new_Jinkela_wire_20825),
        .dout(new_Jinkela_wire_20826)
    );

    spl4L new_Jinkela_splitter_138 (
        .a(new_Jinkela_wire_536),
        .c(new_Jinkela_wire_537),
        .d(new_Jinkela_wire_538),
        .b(new_Jinkela_wire_539),
        .e(new_Jinkela_wire_540)
    );

    spl4L new_Jinkela_splitter_147 (
        .a(new_Jinkela_wire_574),
        .c(new_Jinkela_wire_575),
        .d(new_Jinkela_wire_579),
        .b(new_Jinkela_wire_584),
        .e(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_17379 (
        .din(new_Jinkela_wire_20727),
        .dout(new_Jinkela_wire_20728)
    );

    spl4L new_Jinkela_splitter_139 (
        .a(new_Jinkela_wire_541),
        .c(new_Jinkela_wire_542),
        .d(new_Jinkela_wire_543),
        .b(new_Jinkela_wire_544),
        .e(new_Jinkela_wire_545)
    );

    spl4L new_Jinkela_splitter_141 (
        .a(new_Jinkela_wire_551),
        .c(new_Jinkela_wire_552),
        .d(new_Jinkela_wire_557),
        .b(new_Jinkela_wire_562),
        .e(new_Jinkela_wire_567)
    );

    bfr new_Jinkela_buffer_17552 (
        .din(new_Jinkela_wire_20912),
        .dout(new_Jinkela_wire_20913)
    );

    spl4L new_Jinkela_splitter_143 (
        .a(new_Jinkela_wire_557),
        .c(new_Jinkela_wire_558),
        .d(new_Jinkela_wire_559),
        .b(new_Jinkela_wire_560),
        .e(new_Jinkela_wire_561)
    );

    bfr new_Jinkela_buffer_17380 (
        .din(new_Jinkela_wire_20728),
        .dout(new_Jinkela_wire_20729)
    );

    spl3L new_Jinkela_splitter_137 (
        .a(new_Jinkela_wire_532),
        .d(new_Jinkela_wire_533),
        .b(new_Jinkela_wire_534),
        .c(new_Jinkela_wire_535)
    );

    bfr new_Jinkela_buffer_17472 (
        .din(new_Jinkela_wire_20826),
        .dout(new_Jinkela_wire_20827)
    );

    bfr new_Jinkela_buffer_17381 (
        .din(new_Jinkela_wire_20729),
        .dout(new_Jinkela_wire_20730)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    spl4L new_Jinkela_splitter_140 (
        .a(new_Jinkela_wire_546),
        .c(new_Jinkela_wire_547),
        .d(new_Jinkela_wire_548),
        .b(new_Jinkela_wire_549),
        .e(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_17598 (
        .din(new_Jinkela_wire_20964),
        .dout(new_Jinkela_wire_20965)
    );

    bfr new_Jinkela_buffer_17382 (
        .din(new_Jinkela_wire_20730),
        .dout(new_Jinkela_wire_20731)
    );

    spl3L new_Jinkela_splitter_148 (
        .a(new_Jinkela_wire_575),
        .d(new_Jinkela_wire_576),
        .b(new_Jinkela_wire_577),
        .c(new_Jinkela_wire_578)
    );

    bfr new_Jinkela_buffer_17473 (
        .din(new_Jinkela_wire_20827),
        .dout(new_Jinkela_wire_20828)
    );

    bfr new_Jinkela_buffer_17383 (
        .din(new_Jinkela_wire_20731),
        .dout(new_Jinkela_wire_20732)
    );

    spl4L new_Jinkela_splitter_142 (
        .a(new_Jinkela_wire_552),
        .c(new_Jinkela_wire_553),
        .d(new_Jinkela_wire_554),
        .b(new_Jinkela_wire_555),
        .e(new_Jinkela_wire_556)
    );

    bfr new_Jinkela_buffer_17553 (
        .din(new_Jinkela_wire_20913),
        .dout(new_Jinkela_wire_20914)
    );

    spl4L new_Jinkela_splitter_144 (
        .a(new_Jinkela_wire_562),
        .c(new_Jinkela_wire_563),
        .d(new_Jinkela_wire_564),
        .b(new_Jinkela_wire_565),
        .e(new_Jinkela_wire_566)
    );

    bfr new_Jinkela_buffer_17384 (
        .din(new_Jinkela_wire_20732),
        .dout(new_Jinkela_wire_20733)
    );

    spl4L new_Jinkela_splitter_145 (
        .a(new_Jinkela_wire_567),
        .c(new_Jinkela_wire_568),
        .d(new_Jinkela_wire_569),
        .b(new_Jinkela_wire_570),
        .e(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_17474 (
        .din(new_Jinkela_wire_20828),
        .dout(new_Jinkela_wire_20829)
    );

    spl4L new_Jinkela_splitter_152 (
        .a(new_Jinkela_wire_594),
        .c(new_Jinkela_wire_595),
        .d(new_Jinkela_wire_600),
        .b(new_Jinkela_wire_605),
        .e(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_17385 (
        .din(new_Jinkela_wire_20733),
        .dout(new_Jinkela_wire_20734)
    );

    bfr new_Jinkela_buffer_17625 (
        .din(_0833_),
        .dout(new_Jinkela_wire_20994)
    );

    bfr new_Jinkela_buffer_17386 (
        .din(new_Jinkela_wire_20734),
        .dout(new_Jinkela_wire_20735)
    );

    spl4L new_Jinkela_splitter_149 (
        .a(new_Jinkela_wire_579),
        .c(new_Jinkela_wire_580),
        .d(new_Jinkela_wire_581),
        .b(new_Jinkela_wire_582),
        .e(new_Jinkela_wire_583)
    );

    bfr new_Jinkela_buffer_17475 (
        .din(new_Jinkela_wire_20829),
        .dout(new_Jinkela_wire_20830)
    );

    spl4L new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_600),
        .c(new_Jinkela_wire_601),
        .d(new_Jinkela_wire_602),
        .b(new_Jinkela_wire_603),
        .e(new_Jinkela_wire_604)
    );

    spl4L new_Jinkela_splitter_150 (
        .a(new_Jinkela_wire_584),
        .c(new_Jinkela_wire_585),
        .d(new_Jinkela_wire_586),
        .b(new_Jinkela_wire_587),
        .e(new_Jinkela_wire_588)
    );

    bfr new_Jinkela_buffer_17387 (
        .din(new_Jinkela_wire_20735),
        .dout(new_Jinkela_wire_20736)
    );

    bfr new_Jinkela_buffer_17554 (
        .din(new_Jinkela_wire_20914),
        .dout(new_Jinkela_wire_20915)
    );

    spl4L new_Jinkela_splitter_151 (
        .a(new_Jinkela_wire_589),
        .c(new_Jinkela_wire_590),
        .d(new_Jinkela_wire_591),
        .b(new_Jinkela_wire_592),
        .e(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_17388 (
        .din(new_Jinkela_wire_20736),
        .dout(new_Jinkela_wire_20737)
    );

    spl2 new_Jinkela_splitter_157 (
        .a(N324),
        .b(new_Jinkela_wire_615),
        .c(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_17476 (
        .din(new_Jinkela_wire_20830),
        .dout(new_Jinkela_wire_20831)
    );

    bfr new_Jinkela_buffer_17389 (
        .din(new_Jinkela_wire_20737),
        .dout(new_Jinkela_wire_20738)
    );

    bfr new_Jinkela_buffer_17599 (
        .din(new_Jinkela_wire_20965),
        .dout(new_Jinkela_wire_20966)
    );

    spl4L new_Jinkela_splitter_153 (
        .a(new_Jinkela_wire_595),
        .c(new_Jinkela_wire_596),
        .d(new_Jinkela_wire_597),
        .b(new_Jinkela_wire_598),
        .e(new_Jinkela_wire_599)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_17390 (
        .din(new_Jinkela_wire_20738),
        .dout(new_Jinkela_wire_20739)
    );

    spl4L new_Jinkela_splitter_158 (
        .a(new_Jinkela_wire_617),
        .c(new_Jinkela_wire_618),
        .d(new_Jinkela_wire_622),
        .b(new_Jinkela_wire_627),
        .e(new_Jinkela_wire_632)
    );

    spl4L new_Jinkela_splitter_155 (
        .a(new_Jinkela_wire_605),
        .c(new_Jinkela_wire_606),
        .d(new_Jinkela_wire_607),
        .b(new_Jinkela_wire_608),
        .e(new_Jinkela_wire_609)
    );

    bfr new_Jinkela_buffer_17477 (
        .din(new_Jinkela_wire_20831),
        .dout(new_Jinkela_wire_20832)
    );

    spl4L new_Jinkela_splitter_156 (
        .a(new_Jinkela_wire_610),
        .c(new_Jinkela_wire_611),
        .d(new_Jinkela_wire_612),
        .b(new_Jinkela_wire_613),
        .e(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_17391 (
        .din(new_Jinkela_wire_20739),
        .dout(new_Jinkela_wire_20740)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_17555 (
        .din(new_Jinkela_wire_20915),
        .dout(new_Jinkela_wire_20916)
    );

    spl3L new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_618),
        .d(new_Jinkela_wire_619),
        .b(new_Jinkela_wire_620),
        .c(new_Jinkela_wire_621)
    );

    spl4L new_Jinkela_splitter_177 (
        .a(new_Jinkela_wire_687),
        .c(new_Jinkela_wire_688),
        .d(new_Jinkela_wire_689),
        .b(new_Jinkela_wire_690),
        .e(new_Jinkela_wire_691)
    );

    bfr new_Jinkela_buffer_17392 (
        .din(new_Jinkela_wire_20740),
        .dout(new_Jinkela_wire_20741)
    );

    spl4L new_Jinkela_splitter_160 (
        .a(new_Jinkela_wire_622),
        .c(new_Jinkela_wire_623),
        .d(new_Jinkela_wire_624),
        .b(new_Jinkela_wire_625),
        .e(new_Jinkela_wire_626)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(N341),
        .b(new_Jinkela_wire_637),
        .c(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_17478 (
        .din(new_Jinkela_wire_20832),
        .dout(new_Jinkela_wire_20833)
    );

    bfr new_Jinkela_buffer_17393 (
        .din(new_Jinkela_wire_20741),
        .dout(new_Jinkela_wire_20742)
    );

    spl4L new_Jinkela_splitter_164 (
        .a(new_Jinkela_wire_639),
        .c(new_Jinkela_wire_640),
        .d(new_Jinkela_wire_644),
        .b(new_Jinkela_wire_649),
        .e(new_Jinkela_wire_654)
    );

    spl4L new_Jinkela_splitter_161 (
        .a(new_Jinkela_wire_627),
        .c(new_Jinkela_wire_628),
        .d(new_Jinkela_wire_629),
        .b(new_Jinkela_wire_630),
        .e(new_Jinkela_wire_631)
    );

    bfr new_Jinkela_buffer_17601 (
        .din(_0688_),
        .dout(new_Jinkela_wire_20968)
    );

    spl4L new_Jinkela_splitter_166 (
        .a(new_Jinkela_wire_644),
        .c(new_Jinkela_wire_645),
        .d(new_Jinkela_wire_646),
        .b(new_Jinkela_wire_647),
        .e(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_17394 (
        .din(new_Jinkela_wire_20742),
        .dout(new_Jinkela_wire_20743)
    );

    spl4L new_Jinkela_splitter_162 (
        .a(new_Jinkela_wire_632),
        .c(new_Jinkela_wire_633),
        .d(new_Jinkela_wire_634),
        .b(new_Jinkela_wire_635),
        .e(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_17479 (
        .din(new_Jinkela_wire_20833),
        .dout(new_Jinkela_wire_20834)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_17395 (
        .din(new_Jinkela_wire_20743),
        .dout(new_Jinkela_wire_20744)
    );

    spl3L new_Jinkela_splitter_165 (
        .a(new_Jinkela_wire_640),
        .d(new_Jinkela_wire_641),
        .b(new_Jinkela_wire_642),
        .c(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_17556 (
        .din(new_Jinkela_wire_20916),
        .dout(new_Jinkela_wire_20917)
    );

    bfr new_Jinkela_buffer_17396 (
        .din(new_Jinkela_wire_20744),
        .dout(new_Jinkela_wire_20745)
    );

    spl2 new_Jinkela_splitter_169 (
        .a(N528),
        .b(new_Jinkela_wire_659),
        .c(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_17480 (
        .din(new_Jinkela_wire_20834),
        .dout(new_Jinkela_wire_20835)
    );

    spl4L new_Jinkela_splitter_167 (
        .a(new_Jinkela_wire_649),
        .c(new_Jinkela_wire_650),
        .d(new_Jinkela_wire_651),
        .b(new_Jinkela_wire_652),
        .e(new_Jinkela_wire_653)
    );

    spl4L new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_661),
        .c(new_Jinkela_wire_662),
        .d(new_Jinkela_wire_666),
        .b(new_Jinkela_wire_671),
        .e(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_17397 (
        .din(new_Jinkela_wire_20745),
        .dout(new_Jinkela_wire_20746)
    );

    bfr new_Jinkela_buffer_40 (
        .din(_0481_),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_17600 (
        .din(new_Jinkela_wire_20966),
        .dout(new_Jinkela_wire_20967)
    );

    spl4L new_Jinkela_splitter_168 (
        .a(new_Jinkela_wire_654),
        .c(new_Jinkela_wire_655),
        .d(new_Jinkela_wire_656),
        .b(new_Jinkela_wire_657),
        .e(new_Jinkela_wire_658)
    );

    bfr new_Jinkela_buffer_17398 (
        .din(new_Jinkela_wire_20746),
        .dout(new_Jinkela_wire_20747)
    );

    bfr new_Jinkela_buffer_17481 (
        .din(new_Jinkela_wire_20835),
        .dout(new_Jinkela_wire_20836)
    );

    spl2 new_Jinkela_splitter_180 (
        .a(_1686_),
        .b(new_Jinkela_wire_703),
        .c(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_39 (
        .din(N120),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_17399 (
        .din(new_Jinkela_wire_20747),
        .dout(new_Jinkela_wire_20748)
    );

    spl4L new_Jinkela_splitter_175 (
        .a(new_Jinkela_wire_681),
        .c(new_Jinkela_wire_682),
        .d(new_Jinkela_wire_687),
        .b(new_Jinkela_wire_692),
        .e(new_Jinkela_wire_697)
    );

    bfr new_Jinkela_buffer_7045 (
        .din(new_Jinkela_wire_8806),
        .dout(new_Jinkela_wire_8807)
    );

    bfr new_Jinkela_buffer_10639 (
        .din(new_Jinkela_wire_12840),
        .dout(new_Jinkela_wire_12841)
    );

    bfr new_Jinkela_buffer_7100 (
        .din(new_Jinkela_wire_8879),
        .dout(new_Jinkela_wire_8880)
    );

    bfr new_Jinkela_buffer_10513 (
        .din(new_Jinkela_wire_12690),
        .dout(new_Jinkela_wire_12691)
    );

    bfr new_Jinkela_buffer_7046 (
        .din(new_Jinkela_wire_8807),
        .dout(new_Jinkela_wire_8808)
    );

    bfr new_Jinkela_buffer_10562 (
        .din(new_Jinkela_wire_12761),
        .dout(new_Jinkela_wire_12762)
    );

    bfr new_Jinkela_buffer_7184 (
        .din(new_Jinkela_wire_8967),
        .dout(new_Jinkela_wire_8968)
    );

    bfr new_Jinkela_buffer_10514 (
        .din(new_Jinkela_wire_12691),
        .dout(new_Jinkela_wire_12692)
    );

    bfr new_Jinkela_buffer_7047 (
        .din(new_Jinkela_wire_8808),
        .dout(new_Jinkela_wire_8809)
    );

    bfr new_Jinkela_buffer_10798 (
        .din(new_Jinkela_wire_13007),
        .dout(new_Jinkela_wire_13008)
    );

    bfr new_Jinkela_buffer_7101 (
        .din(new_Jinkela_wire_8880),
        .dout(new_Jinkela_wire_8881)
    );

    bfr new_Jinkela_buffer_10515 (
        .din(new_Jinkela_wire_12692),
        .dout(new_Jinkela_wire_12693)
    );

    bfr new_Jinkela_buffer_7048 (
        .din(new_Jinkela_wire_8809),
        .dout(new_Jinkela_wire_8810)
    );

    bfr new_Jinkela_buffer_10563 (
        .din(new_Jinkela_wire_12762),
        .dout(new_Jinkela_wire_12763)
    );

    bfr new_Jinkela_buffer_10516 (
        .din(new_Jinkela_wire_12693),
        .dout(new_Jinkela_wire_12694)
    );

    bfr new_Jinkela_buffer_7049 (
        .din(new_Jinkela_wire_8810),
        .dout(new_Jinkela_wire_8811)
    );

    bfr new_Jinkela_buffer_10640 (
        .din(new_Jinkela_wire_12841),
        .dout(new_Jinkela_wire_12842)
    );

    bfr new_Jinkela_buffer_7102 (
        .din(new_Jinkela_wire_8881),
        .dout(new_Jinkela_wire_8882)
    );

    bfr new_Jinkela_buffer_10517 (
        .din(new_Jinkela_wire_12694),
        .dout(new_Jinkela_wire_12695)
    );

    bfr new_Jinkela_buffer_7050 (
        .din(new_Jinkela_wire_8811),
        .dout(new_Jinkela_wire_8812)
    );

    bfr new_Jinkela_buffer_10564 (
        .din(new_Jinkela_wire_12763),
        .dout(new_Jinkela_wire_12764)
    );

    bfr new_Jinkela_buffer_7185 (
        .din(new_Jinkela_wire_8968),
        .dout(new_Jinkela_wire_8969)
    );

    bfr new_Jinkela_buffer_10518 (
        .din(new_Jinkela_wire_12695),
        .dout(new_Jinkela_wire_12696)
    );

    bfr new_Jinkela_buffer_7051 (
        .din(new_Jinkela_wire_8812),
        .dout(new_Jinkela_wire_8813)
    );

    bfr new_Jinkela_buffer_10706 (
        .din(new_Jinkela_wire_12911),
        .dout(new_Jinkela_wire_12912)
    );

    bfr new_Jinkela_buffer_7103 (
        .din(new_Jinkela_wire_8882),
        .dout(new_Jinkela_wire_8883)
    );

    bfr new_Jinkela_buffer_10519 (
        .din(new_Jinkela_wire_12696),
        .dout(new_Jinkela_wire_12697)
    );

    bfr new_Jinkela_buffer_7052 (
        .din(new_Jinkela_wire_8813),
        .dout(new_Jinkela_wire_8814)
    );

    bfr new_Jinkela_buffer_10565 (
        .din(new_Jinkela_wire_12764),
        .dout(new_Jinkela_wire_12765)
    );

    bfr new_Jinkela_buffer_7188 (
        .din(new_Jinkela_wire_8971),
        .dout(new_Jinkela_wire_8972)
    );

    bfr new_Jinkela_buffer_10520 (
        .din(new_Jinkela_wire_12697),
        .dout(new_Jinkela_wire_12698)
    );

    bfr new_Jinkela_buffer_7053 (
        .din(new_Jinkela_wire_8814),
        .dout(new_Jinkela_wire_8815)
    );

    bfr new_Jinkela_buffer_10641 (
        .din(new_Jinkela_wire_12842),
        .dout(new_Jinkela_wire_12843)
    );

    bfr new_Jinkela_buffer_7104 (
        .din(new_Jinkela_wire_8883),
        .dout(new_Jinkela_wire_8884)
    );

    bfr new_Jinkela_buffer_10521 (
        .din(new_Jinkela_wire_12698),
        .dout(new_Jinkela_wire_12699)
    );

    bfr new_Jinkela_buffer_7054 (
        .din(new_Jinkela_wire_8815),
        .dout(new_Jinkela_wire_8816)
    );

    bfr new_Jinkela_buffer_10566 (
        .din(new_Jinkela_wire_12765),
        .dout(new_Jinkela_wire_12766)
    );

    bfr new_Jinkela_buffer_10522 (
        .din(new_Jinkela_wire_12699),
        .dout(new_Jinkela_wire_12700)
    );

    bfr new_Jinkela_buffer_7227 (
        .din(_1271_),
        .dout(new_Jinkela_wire_9019)
    );

    bfr new_Jinkela_buffer_7055 (
        .din(new_Jinkela_wire_8816),
        .dout(new_Jinkela_wire_8817)
    );

    bfr new_Jinkela_buffer_10803 (
        .din(_0234_),
        .dout(new_Jinkela_wire_13015)
    );

    bfr new_Jinkela_buffer_7105 (
        .din(new_Jinkela_wire_8884),
        .dout(new_Jinkela_wire_8885)
    );

    bfr new_Jinkela_buffer_10523 (
        .din(new_Jinkela_wire_12700),
        .dout(new_Jinkela_wire_12701)
    );

    bfr new_Jinkela_buffer_7056 (
        .din(new_Jinkela_wire_8817),
        .dout(new_Jinkela_wire_8818)
    );

    bfr new_Jinkela_buffer_10567 (
        .din(new_Jinkela_wire_12766),
        .dout(new_Jinkela_wire_12767)
    );

    bfr new_Jinkela_buffer_7189 (
        .din(new_Jinkela_wire_8972),
        .dout(new_Jinkela_wire_8973)
    );

    bfr new_Jinkela_buffer_10524 (
        .din(new_Jinkela_wire_12701),
        .dout(new_Jinkela_wire_12702)
    );

    bfr new_Jinkela_buffer_7057 (
        .din(new_Jinkela_wire_8818),
        .dout(new_Jinkela_wire_8819)
    );

    bfr new_Jinkela_buffer_10642 (
        .din(new_Jinkela_wire_12843),
        .dout(new_Jinkela_wire_12844)
    );

    bfr new_Jinkela_buffer_7106 (
        .din(new_Jinkela_wire_8885),
        .dout(new_Jinkela_wire_8886)
    );

    bfr new_Jinkela_buffer_10525 (
        .din(new_Jinkela_wire_12702),
        .dout(new_Jinkela_wire_12703)
    );

    bfr new_Jinkela_buffer_7058 (
        .din(new_Jinkela_wire_8819),
        .dout(new_Jinkela_wire_8820)
    );

    bfr new_Jinkela_buffer_10568 (
        .din(new_Jinkela_wire_12767),
        .dout(new_Jinkela_wire_12768)
    );

    bfr new_Jinkela_buffer_7226 (
        .din(new_Jinkela_wire_9013),
        .dout(new_Jinkela_wire_9014)
    );

    bfr new_Jinkela_buffer_10526 (
        .din(new_Jinkela_wire_12703),
        .dout(new_Jinkela_wire_12704)
    );

    spl2 new_Jinkela_splitter_746 (
        .a(_1150_),
        .b(new_Jinkela_wire_9094),
        .c(new_Jinkela_wire_9095)
    );

    bfr new_Jinkela_buffer_7059 (
        .din(new_Jinkela_wire_8820),
        .dout(new_Jinkela_wire_8821)
    );

    bfr new_Jinkela_buffer_10707 (
        .din(new_Jinkela_wire_12912),
        .dout(new_Jinkela_wire_12913)
    );

    bfr new_Jinkela_buffer_7107 (
        .din(new_Jinkela_wire_8886),
        .dout(new_Jinkela_wire_8887)
    );

    bfr new_Jinkela_buffer_10527 (
        .din(new_Jinkela_wire_12704),
        .dout(new_Jinkela_wire_12705)
    );

    bfr new_Jinkela_buffer_7060 (
        .din(new_Jinkela_wire_8821),
        .dout(new_Jinkela_wire_8822)
    );

    bfr new_Jinkela_buffer_10569 (
        .din(new_Jinkela_wire_12768),
        .dout(new_Jinkela_wire_12769)
    );

    bfr new_Jinkela_buffer_7190 (
        .din(new_Jinkela_wire_8973),
        .dout(new_Jinkela_wire_8974)
    );

    bfr new_Jinkela_buffer_10528 (
        .din(new_Jinkela_wire_12705),
        .dout(new_Jinkela_wire_12706)
    );

    bfr new_Jinkela_buffer_7061 (
        .din(new_Jinkela_wire_8822),
        .dout(new_Jinkela_wire_8823)
    );

    bfr new_Jinkela_buffer_10643 (
        .din(new_Jinkela_wire_12844),
        .dout(new_Jinkela_wire_12845)
    );

    bfr new_Jinkela_buffer_7108 (
        .din(new_Jinkela_wire_8887),
        .dout(new_Jinkela_wire_8888)
    );

    bfr new_Jinkela_buffer_10529 (
        .din(new_Jinkela_wire_12706),
        .dout(new_Jinkela_wire_12707)
    );

    bfr new_Jinkela_buffer_7062 (
        .din(new_Jinkela_wire_8823),
        .dout(new_Jinkela_wire_8824)
    );

    bfr new_Jinkela_buffer_10570 (
        .din(new_Jinkela_wire_12769),
        .dout(new_Jinkela_wire_12770)
    );

    bfr new_Jinkela_buffer_7228 (
        .din(_0540_),
        .dout(new_Jinkela_wire_9020)
    );

    bfr new_Jinkela_buffer_10530 (
        .din(new_Jinkela_wire_12707),
        .dout(new_Jinkela_wire_12708)
    );

    spl2 new_Jinkela_splitter_743 (
        .a(new_Jinkela_wire_9014),
        .b(new_Jinkela_wire_9015),
        .c(new_Jinkela_wire_9016)
    );

    bfr new_Jinkela_buffer_7063 (
        .din(new_Jinkela_wire_8824),
        .dout(new_Jinkela_wire_8825)
    );

    bfr new_Jinkela_buffer_10799 (
        .din(new_Jinkela_wire_13008),
        .dout(new_Jinkela_wire_13009)
    );

    bfr new_Jinkela_buffer_7109 (
        .din(new_Jinkela_wire_8888),
        .dout(new_Jinkela_wire_8889)
    );

    spl2 new_Jinkela_splitter_938 (
        .a(new_Jinkela_wire_12708),
        .b(new_Jinkela_wire_12709),
        .c(new_Jinkela_wire_12710)
    );

    bfr new_Jinkela_buffer_7064 (
        .din(new_Jinkela_wire_8825),
        .dout(new_Jinkela_wire_8826)
    );

    bfr new_Jinkela_buffer_10644 (
        .din(new_Jinkela_wire_12845),
        .dout(new_Jinkela_wire_12846)
    );

    bfr new_Jinkela_buffer_7191 (
        .din(new_Jinkela_wire_8974),
        .dout(new_Jinkela_wire_8975)
    );

    bfr new_Jinkela_buffer_10571 (
        .din(new_Jinkela_wire_12770),
        .dout(new_Jinkela_wire_12771)
    );

    bfr new_Jinkela_buffer_7065 (
        .din(new_Jinkela_wire_8826),
        .dout(new_Jinkela_wire_8827)
    );

    bfr new_Jinkela_buffer_10572 (
        .din(new_Jinkela_wire_12771),
        .dout(new_Jinkela_wire_12772)
    );

    bfr new_Jinkela_buffer_7110 (
        .din(new_Jinkela_wire_8889),
        .dout(new_Jinkela_wire_8890)
    );

    bfr new_Jinkela_buffer_10708 (
        .din(new_Jinkela_wire_12913),
        .dout(new_Jinkela_wire_12914)
    );

    bfr new_Jinkela_buffer_3613 (
        .din(new_Jinkela_wire_4794),
        .dout(new_Jinkela_wire_4795)
    );

    bfr new_Jinkela_buffer_14046 (
        .din(new_Jinkela_wire_16733),
        .dout(new_Jinkela_wire_16734)
    );

    bfr new_Jinkela_buffer_13989 (
        .din(new_Jinkela_wire_16672),
        .dout(new_Jinkela_wire_16673)
    );

    bfr new_Jinkela_buffer_3712 (
        .din(new_Jinkela_wire_4923),
        .dout(new_Jinkela_wire_4924)
    );

    bfr new_Jinkela_buffer_3614 (
        .din(new_Jinkela_wire_4795),
        .dout(new_Jinkela_wire_4796)
    );

    bfr new_Jinkela_buffer_13990 (
        .din(new_Jinkela_wire_16673),
        .dout(new_Jinkela_wire_16674)
    );

    bfr new_Jinkela_buffer_3675 (
        .din(new_Jinkela_wire_4868),
        .dout(new_Jinkela_wire_4869)
    );

    spl2 new_Jinkela_splitter_1207 (
        .a(_0187_),
        .b(new_Jinkela_wire_16906),
        .c(new_Jinkela_wire_16907)
    );

    bfr new_Jinkela_buffer_3615 (
        .din(new_Jinkela_wire_4796),
        .dout(new_Jinkela_wire_4797)
    );

    bfr new_Jinkela_buffer_14047 (
        .din(new_Jinkela_wire_16734),
        .dout(new_Jinkela_wire_16735)
    );

    bfr new_Jinkela_buffer_13991 (
        .din(new_Jinkela_wire_16674),
        .dout(new_Jinkela_wire_16675)
    );

    spl2 new_Jinkela_splitter_460 (
        .a(_0500_),
        .b(new_Jinkela_wire_4999),
        .c(new_Jinkela_wire_5000)
    );

    bfr new_Jinkela_buffer_3616 (
        .din(new_Jinkela_wire_4797),
        .dout(new_Jinkela_wire_4798)
    );

    bfr new_Jinkela_buffer_14104 (
        .din(new_Jinkela_wire_16807),
        .dout(new_Jinkela_wire_16808)
    );

    bfr new_Jinkela_buffer_13992 (
        .din(new_Jinkela_wire_16675),
        .dout(new_Jinkela_wire_16676)
    );

    bfr new_Jinkela_buffer_3676 (
        .din(new_Jinkela_wire_4869),
        .dout(new_Jinkela_wire_4870)
    );

    bfr new_Jinkela_buffer_3617 (
        .din(new_Jinkela_wire_4798),
        .dout(new_Jinkela_wire_4799)
    );

    bfr new_Jinkela_buffer_14048 (
        .din(new_Jinkela_wire_16735),
        .dout(new_Jinkela_wire_16736)
    );

    bfr new_Jinkela_buffer_13993 (
        .din(new_Jinkela_wire_16676),
        .dout(new_Jinkela_wire_16677)
    );

    bfr new_Jinkela_buffer_3713 (
        .din(new_Jinkela_wire_4924),
        .dout(new_Jinkela_wire_4925)
    );

    bfr new_Jinkela_buffer_3618 (
        .din(new_Jinkela_wire_4799),
        .dout(new_Jinkela_wire_4800)
    );

    bfr new_Jinkela_buffer_13994 (
        .din(new_Jinkela_wire_16677),
        .dout(new_Jinkela_wire_16678)
    );

    bfr new_Jinkela_buffer_3677 (
        .din(new_Jinkela_wire_4870),
        .dout(new_Jinkela_wire_4871)
    );

    bfr new_Jinkela_buffer_3619 (
        .din(new_Jinkela_wire_4800),
        .dout(new_Jinkela_wire_4801)
    );

    bfr new_Jinkela_buffer_14049 (
        .din(new_Jinkela_wire_16736),
        .dout(new_Jinkela_wire_16737)
    );

    bfr new_Jinkela_buffer_13995 (
        .din(new_Jinkela_wire_16678),
        .dout(new_Jinkela_wire_16679)
    );

    bfr new_Jinkela_buffer_3773 (
        .din(new_Jinkela_wire_4992),
        .dout(new_Jinkela_wire_4993)
    );

    bfr new_Jinkela_buffer_3620 (
        .din(new_Jinkela_wire_4801),
        .dout(new_Jinkela_wire_4802)
    );

    bfr new_Jinkela_buffer_14105 (
        .din(new_Jinkela_wire_16808),
        .dout(new_Jinkela_wire_16809)
    );

    bfr new_Jinkela_buffer_13996 (
        .din(new_Jinkela_wire_16679),
        .dout(new_Jinkela_wire_16680)
    );

    bfr new_Jinkela_buffer_3678 (
        .din(new_Jinkela_wire_4871),
        .dout(new_Jinkela_wire_4872)
    );

    bfr new_Jinkela_buffer_3621 (
        .din(new_Jinkela_wire_4802),
        .dout(new_Jinkela_wire_4803)
    );

    bfr new_Jinkela_buffer_14050 (
        .din(new_Jinkela_wire_16737),
        .dout(new_Jinkela_wire_16738)
    );

    bfr new_Jinkela_buffer_13997 (
        .din(new_Jinkela_wire_16680),
        .dout(new_Jinkela_wire_16681)
    );

    bfr new_Jinkela_buffer_3714 (
        .din(new_Jinkela_wire_4925),
        .dout(new_Jinkela_wire_4926)
    );

    bfr new_Jinkela_buffer_3622 (
        .din(new_Jinkela_wire_4803),
        .dout(new_Jinkela_wire_4804)
    );

    bfr new_Jinkela_buffer_14163 (
        .din(new_Jinkela_wire_16876),
        .dout(new_Jinkela_wire_16877)
    );

    bfr new_Jinkela_buffer_13998 (
        .din(new_Jinkela_wire_16681),
        .dout(new_Jinkela_wire_16682)
    );

    bfr new_Jinkela_buffer_3679 (
        .din(new_Jinkela_wire_4872),
        .dout(new_Jinkela_wire_4873)
    );

    bfr new_Jinkela_buffer_3623 (
        .din(new_Jinkela_wire_4804),
        .dout(new_Jinkela_wire_4805)
    );

    bfr new_Jinkela_buffer_14051 (
        .din(new_Jinkela_wire_16738),
        .dout(new_Jinkela_wire_16739)
    );

    bfr new_Jinkela_buffer_13999 (
        .din(new_Jinkela_wire_16682),
        .dout(new_Jinkela_wire_16683)
    );

    bfr new_Jinkela_buffer_3777 (
        .din(_1017_),
        .dout(new_Jinkela_wire_5001)
    );

    bfr new_Jinkela_buffer_3624 (
        .din(new_Jinkela_wire_4805),
        .dout(new_Jinkela_wire_4806)
    );

    bfr new_Jinkela_buffer_14106 (
        .din(new_Jinkela_wire_16809),
        .dout(new_Jinkela_wire_16810)
    );

    bfr new_Jinkela_buffer_14000 (
        .din(new_Jinkela_wire_16683),
        .dout(new_Jinkela_wire_16684)
    );

    bfr new_Jinkela_buffer_3680 (
        .din(new_Jinkela_wire_4873),
        .dout(new_Jinkela_wire_4874)
    );

    bfr new_Jinkela_buffer_3625 (
        .din(new_Jinkela_wire_4806),
        .dout(new_Jinkela_wire_4807)
    );

    bfr new_Jinkela_buffer_14052 (
        .din(new_Jinkela_wire_16739),
        .dout(new_Jinkela_wire_16740)
    );

    bfr new_Jinkela_buffer_14001 (
        .din(new_Jinkela_wire_16684),
        .dout(new_Jinkela_wire_16685)
    );

    bfr new_Jinkela_buffer_3715 (
        .din(new_Jinkela_wire_4926),
        .dout(new_Jinkela_wire_4927)
    );

    bfr new_Jinkela_buffer_3626 (
        .din(new_Jinkela_wire_4807),
        .dout(new_Jinkela_wire_4808)
    );

    spl2 new_Jinkela_splitter_1208 (
        .a(_1652_),
        .b(new_Jinkela_wire_16909),
        .c(new_Jinkela_wire_16910)
    );

    bfr new_Jinkela_buffer_14002 (
        .din(new_Jinkela_wire_16685),
        .dout(new_Jinkela_wire_16686)
    );

    bfr new_Jinkela_buffer_3681 (
        .din(new_Jinkela_wire_4874),
        .dout(new_Jinkela_wire_4875)
    );

    bfr new_Jinkela_buffer_14190 (
        .din(_0448_),
        .dout(new_Jinkela_wire_16908)
    );

    bfr new_Jinkela_buffer_3627 (
        .din(new_Jinkela_wire_4808),
        .dout(new_Jinkela_wire_4809)
    );

    bfr new_Jinkela_buffer_14053 (
        .din(new_Jinkela_wire_16740),
        .dout(new_Jinkela_wire_16741)
    );

    bfr new_Jinkela_buffer_14003 (
        .din(new_Jinkela_wire_16686),
        .dout(new_Jinkela_wire_16687)
    );

    bfr new_Jinkela_buffer_3774 (
        .din(new_Jinkela_wire_4993),
        .dout(new_Jinkela_wire_4994)
    );

    bfr new_Jinkela_buffer_3628 (
        .din(new_Jinkela_wire_4809),
        .dout(new_Jinkela_wire_4810)
    );

    bfr new_Jinkela_buffer_14107 (
        .din(new_Jinkela_wire_16810),
        .dout(new_Jinkela_wire_16811)
    );

    bfr new_Jinkela_buffer_14004 (
        .din(new_Jinkela_wire_16687),
        .dout(new_Jinkela_wire_16688)
    );

    bfr new_Jinkela_buffer_3682 (
        .din(new_Jinkela_wire_4875),
        .dout(new_Jinkela_wire_4876)
    );

    bfr new_Jinkela_buffer_3629 (
        .din(new_Jinkela_wire_4810),
        .dout(new_Jinkela_wire_4811)
    );

    bfr new_Jinkela_buffer_14054 (
        .din(new_Jinkela_wire_16741),
        .dout(new_Jinkela_wire_16742)
    );

    bfr new_Jinkela_buffer_14005 (
        .din(new_Jinkela_wire_16688),
        .dout(new_Jinkela_wire_16689)
    );

    bfr new_Jinkela_buffer_3716 (
        .din(new_Jinkela_wire_4927),
        .dout(new_Jinkela_wire_4928)
    );

    bfr new_Jinkela_buffer_3630 (
        .din(new_Jinkela_wire_4811),
        .dout(new_Jinkela_wire_4812)
    );

    bfr new_Jinkela_buffer_14164 (
        .din(new_Jinkela_wire_16877),
        .dout(new_Jinkela_wire_16878)
    );

    bfr new_Jinkela_buffer_14006 (
        .din(new_Jinkela_wire_16689),
        .dout(new_Jinkela_wire_16690)
    );

    bfr new_Jinkela_buffer_3683 (
        .din(new_Jinkela_wire_4876),
        .dout(new_Jinkela_wire_4877)
    );

    bfr new_Jinkela_buffer_3631 (
        .din(new_Jinkela_wire_4812),
        .dout(new_Jinkela_wire_4813)
    );

    bfr new_Jinkela_buffer_14055 (
        .din(new_Jinkela_wire_16742),
        .dout(new_Jinkela_wire_16743)
    );

    bfr new_Jinkela_buffer_14007 (
        .din(new_Jinkela_wire_16690),
        .dout(new_Jinkela_wire_16691)
    );

    spl2 new_Jinkela_splitter_462 (
        .a(_1621_),
        .b(new_Jinkela_wire_5043),
        .c(new_Jinkela_wire_5044)
    );

    bfr new_Jinkela_buffer_3632 (
        .din(new_Jinkela_wire_4813),
        .dout(new_Jinkela_wire_4814)
    );

    bfr new_Jinkela_buffer_14108 (
        .din(new_Jinkela_wire_16811),
        .dout(new_Jinkela_wire_16812)
    );

    bfr new_Jinkela_buffer_14008 (
        .din(new_Jinkela_wire_16691),
        .dout(new_Jinkela_wire_16692)
    );

    bfr new_Jinkela_buffer_3684 (
        .din(new_Jinkela_wire_4877),
        .dout(new_Jinkela_wire_4878)
    );

    bfr new_Jinkela_buffer_3633 (
        .din(new_Jinkela_wire_4814),
        .dout(new_Jinkela_wire_4815)
    );

    bfr new_Jinkela_buffer_14056 (
        .din(new_Jinkela_wire_16743),
        .dout(new_Jinkela_wire_16744)
    );

    bfr new_Jinkela_buffer_14009 (
        .din(new_Jinkela_wire_16692),
        .dout(new_Jinkela_wire_16693)
    );

    bfr new_Jinkela_buffer_3717 (
        .din(new_Jinkela_wire_4928),
        .dout(new_Jinkela_wire_4929)
    );

    bfr new_Jinkela_buffer_17557 (
        .din(new_Jinkela_wire_20917),
        .dout(new_Jinkela_wire_20918)
    );

    spl4L new_Jinkela_splitter_173 (
        .a(new_Jinkela_wire_671),
        .c(new_Jinkela_wire_672),
        .d(new_Jinkela_wire_673),
        .b(new_Jinkela_wire_674),
        .e(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_17400 (
        .din(new_Jinkela_wire_20748),
        .dout(new_Jinkela_wire_20749)
    );

    spl4L new_Jinkela_splitter_172 (
        .a(new_Jinkela_wire_666),
        .c(new_Jinkela_wire_667),
        .d(new_Jinkela_wire_668),
        .b(new_Jinkela_wire_669),
        .e(new_Jinkela_wire_670)
    );

    spl3L new_Jinkela_splitter_171 (
        .a(new_Jinkela_wire_662),
        .d(new_Jinkela_wire_663),
        .b(new_Jinkela_wire_664),
        .c(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_17482 (
        .din(new_Jinkela_wire_20836),
        .dout(new_Jinkela_wire_20837)
    );

    bfr new_Jinkela_buffer_17401 (
        .din(new_Jinkela_wire_20749),
        .dout(new_Jinkela_wire_20750)
    );

    spl2 new_Jinkela_splitter_183 (
        .a(_1239_),
        .b(new_Jinkela_wire_714),
        .c(new_Jinkela_wire_715)
    );

    spl4L new_Jinkela_splitter_174 (
        .a(new_Jinkela_wire_676),
        .c(new_Jinkela_wire_677),
        .d(new_Jinkela_wire_678),
        .b(new_Jinkela_wire_679),
        .e(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_17602 (
        .din(new_Jinkela_wire_20968),
        .dout(new_Jinkela_wire_20969)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(_1666_),
        .b(new_Jinkela_wire_708),
        .c(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_17402 (
        .din(new_Jinkela_wire_20750),
        .dout(new_Jinkela_wire_20751)
    );

    bfr new_Jinkela_buffer_41 (
        .din(_0807_),
        .dout(new_Jinkela_wire_705)
    );

    spl4L new_Jinkela_splitter_176 (
        .a(new_Jinkela_wire_682),
        .c(new_Jinkela_wire_683),
        .d(new_Jinkela_wire_684),
        .b(new_Jinkela_wire_685),
        .e(new_Jinkela_wire_686)
    );

    bfr new_Jinkela_buffer_17483 (
        .din(new_Jinkela_wire_20837),
        .dout(new_Jinkela_wire_20838)
    );

    spl4L new_Jinkela_splitter_178 (
        .a(new_Jinkela_wire_692),
        .c(new_Jinkela_wire_693),
        .d(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_695),
        .e(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_17403 (
        .din(new_Jinkela_wire_20751),
        .dout(new_Jinkela_wire_20752)
    );

    bfr new_Jinkela_buffer_17558 (
        .din(new_Jinkela_wire_20918),
        .dout(new_Jinkela_wire_20919)
    );

    bfr new_Jinkela_buffer_17404 (
        .din(new_Jinkela_wire_20752),
        .dout(new_Jinkela_wire_20753)
    );

    spl4L new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_697),
        .c(new_Jinkela_wire_698),
        .d(new_Jinkela_wire_699),
        .b(new_Jinkela_wire_700),
        .e(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_17484 (
        .din(new_Jinkela_wire_20838),
        .dout(new_Jinkela_wire_20839)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(_0152_),
        .b(new_Jinkela_wire_706),
        .c(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_17405 (
        .din(new_Jinkela_wire_20753),
        .dout(new_Jinkela_wire_20754)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    spl2 new_Jinkela_splitter_1535 (
        .a(_0985_),
        .b(new_Jinkela_wire_21094),
        .c(new_Jinkela_wire_21095)
    );

    spl2 new_Jinkela_splitter_184 (
        .a(_1240_),
        .b(new_Jinkela_wire_716),
        .c(new_Jinkela_wire_717)
    );

    bfr new_Jinkela_buffer_17406 (
        .din(new_Jinkela_wire_20754),
        .dout(new_Jinkela_wire_20755)
    );

    bfr new_Jinkela_buffer_17485 (
        .din(new_Jinkela_wire_20839),
        .dout(new_Jinkela_wire_20840)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_17407 (
        .din(new_Jinkela_wire_20755),
        .dout(new_Jinkela_wire_20756)
    );

    spl2 new_Jinkela_splitter_185 (
        .a(_1482_),
        .b(new_Jinkela_wire_718),
        .c(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_17559 (
        .din(new_Jinkela_wire_20919),
        .dout(new_Jinkela_wire_20920)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_17408 (
        .din(new_Jinkela_wire_20756),
        .dout(new_Jinkela_wire_20757)
    );

    bfr new_Jinkela_buffer_46 (
        .din(_1530_),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_17486 (
        .din(new_Jinkela_wire_20840),
        .dout(new_Jinkela_wire_20841)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_17409 (
        .din(new_Jinkela_wire_20757),
        .dout(new_Jinkela_wire_20758)
    );

    bfr new_Jinkela_buffer_47 (
        .din(_0214_),
        .dout(new_Jinkela_wire_723)
    );

    spl2 new_Jinkela_splitter_186 (
        .a(_0976_),
        .b(new_Jinkela_wire_721),
        .c(new_Jinkela_wire_722)
    );

    bfr new_Jinkela_buffer_17603 (
        .din(new_Jinkela_wire_20969),
        .dout(new_Jinkela_wire_20970)
    );

    bfr new_Jinkela_buffer_152 (
        .din(_1176_),
        .dout(new_Jinkela_wire_832)
    );

    bfr new_Jinkela_buffer_17410 (
        .din(new_Jinkela_wire_20758),
        .dout(new_Jinkela_wire_20759)
    );

    spl2 new_Jinkela_splitter_188 (
        .a(_1544_),
        .b(new_Jinkela_wire_830),
        .c(new_Jinkela_wire_831)
    );

    bfr new_Jinkela_buffer_17487 (
        .din(new_Jinkela_wire_20841),
        .dout(new_Jinkela_wire_20842)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_17411 (
        .din(new_Jinkela_wire_20759),
        .dout(new_Jinkela_wire_20760)
    );

    spl2 new_Jinkela_splitter_189 (
        .a(_0979_),
        .b(new_Jinkela_wire_834),
        .c(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_17560 (
        .din(new_Jinkela_wire_20920),
        .dout(new_Jinkela_wire_20921)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_17412 (
        .din(new_Jinkela_wire_20760),
        .dout(new_Jinkela_wire_20761)
    );

    bfr new_Jinkela_buffer_153 (
        .din(_0406_),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_17488 (
        .din(new_Jinkela_wire_20842),
        .dout(new_Jinkela_wire_20843)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_17413 (
        .din(new_Jinkela_wire_20761),
        .dout(new_Jinkela_wire_20762)
    );

    spl2 new_Jinkela_splitter_190 (
        .a(_1389_),
        .b(new_Jinkela_wire_836),
        .c(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_156 (
        .din(_0564_),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_17626 (
        .din(new_Jinkela_wire_20994),
        .dout(new_Jinkela_wire_20995)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_726),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_17414 (
        .din(new_Jinkela_wire_20762),
        .dout(new_Jinkela_wire_20763)
    );

    bfr new_Jinkela_buffer_17489 (
        .din(new_Jinkela_wire_20843),
        .dout(new_Jinkela_wire_20844)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_17415 (
        .din(new_Jinkela_wire_20763),
        .dout(new_Jinkela_wire_20764)
    );

    bfr new_Jinkela_buffer_154 (
        .din(_1086_),
        .dout(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_17561 (
        .din(new_Jinkela_wire_20921),
        .dout(new_Jinkela_wire_20922)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_17416 (
        .din(new_Jinkela_wire_20764),
        .dout(new_Jinkela_wire_20765)
    );

    bfr new_Jinkela_buffer_155 (
        .din(_0763_),
        .dout(new_Jinkela_wire_839)
    );

    bfr new_Jinkela_buffer_17490 (
        .din(new_Jinkela_wire_20844),
        .dout(new_Jinkela_wire_20845)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_729),
        .dout(new_Jinkela_wire_730)
    );

    bfr new_Jinkela_buffer_17417 (
        .din(new_Jinkela_wire_20765),
        .dout(new_Jinkela_wire_20766)
    );

    spl2 new_Jinkela_splitter_191 (
        .a(_1398_),
        .b(new_Jinkela_wire_841),
        .c(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_17604 (
        .din(new_Jinkela_wire_20970),
        .dout(new_Jinkela_wire_20971)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    spl2 new_Jinkela_splitter_1534 (
        .a(_0783_),
        .b(new_Jinkela_wire_21092),
        .c(new_Jinkela_wire_21093)
    );

    bfr new_Jinkela_buffer_17418 (
        .din(new_Jinkela_wire_20766),
        .dout(new_Jinkela_wire_20767)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(_0700_),
        .b(new_Jinkela_wire_843),
        .c(new_Jinkela_wire_844)
    );

    bfr new_Jinkela_buffer_157 (
        .din(_0463_),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_17491 (
        .din(new_Jinkela_wire_20845),
        .dout(new_Jinkela_wire_20846)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_731),
        .dout(new_Jinkela_wire_732)
    );

    bfr new_Jinkela_buffer_17419 (
        .din(new_Jinkela_wire_20767),
        .dout(new_Jinkela_wire_20768)
    );

    bfr new_Jinkela_buffer_17562 (
        .din(new_Jinkela_wire_20922),
        .dout(new_Jinkela_wire_20923)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_17420 (
        .din(new_Jinkela_wire_20768),
        .dout(new_Jinkela_wire_20769)
    );

    bfr new_Jinkela_buffer_7066 (
        .din(new_Jinkela_wire_8827),
        .dout(new_Jinkela_wire_8828)
    );

    bfr new_Jinkela_buffer_3634 (
        .din(new_Jinkela_wire_4815),
        .dout(new_Jinkela_wire_4816)
    );

    bfr new_Jinkela_buffer_3685 (
        .din(new_Jinkela_wire_4878),
        .dout(new_Jinkela_wire_4879)
    );

    bfr new_Jinkela_buffer_7300 (
        .din(_0425_),
        .dout(new_Jinkela_wire_9096)
    );

    bfr new_Jinkela_buffer_7067 (
        .din(new_Jinkela_wire_8828),
        .dout(new_Jinkela_wire_8829)
    );

    bfr new_Jinkela_buffer_3635 (
        .din(new_Jinkela_wire_4816),
        .dout(new_Jinkela_wire_4817)
    );

    bfr new_Jinkela_buffer_7111 (
        .din(new_Jinkela_wire_8890),
        .dout(new_Jinkela_wire_8891)
    );

    spl2 new_Jinkela_splitter_463 (
        .a(_0753_),
        .b(new_Jinkela_wire_5045),
        .c(new_Jinkela_wire_5046)
    );

    bfr new_Jinkela_buffer_7068 (
        .din(new_Jinkela_wire_8829),
        .dout(new_Jinkela_wire_8830)
    );

    bfr new_Jinkela_buffer_3636 (
        .din(new_Jinkela_wire_4817),
        .dout(new_Jinkela_wire_4818)
    );

    bfr new_Jinkela_buffer_7192 (
        .din(new_Jinkela_wire_8975),
        .dout(new_Jinkela_wire_8976)
    );

    bfr new_Jinkela_buffer_3686 (
        .din(new_Jinkela_wire_4879),
        .dout(new_Jinkela_wire_4880)
    );

    bfr new_Jinkela_buffer_7069 (
        .din(new_Jinkela_wire_8830),
        .dout(new_Jinkela_wire_8831)
    );

    bfr new_Jinkela_buffer_3637 (
        .din(new_Jinkela_wire_4818),
        .dout(new_Jinkela_wire_4819)
    );

    bfr new_Jinkela_buffer_7112 (
        .din(new_Jinkela_wire_8891),
        .dout(new_Jinkela_wire_8892)
    );

    bfr new_Jinkela_buffer_3718 (
        .din(new_Jinkela_wire_4929),
        .dout(new_Jinkela_wire_4930)
    );

    bfr new_Jinkela_buffer_7070 (
        .din(new_Jinkela_wire_8831),
        .dout(new_Jinkela_wire_8832)
    );

    bfr new_Jinkela_buffer_3638 (
        .din(new_Jinkela_wire_4819),
        .dout(new_Jinkela_wire_4820)
    );

    bfr new_Jinkela_buffer_7229 (
        .din(new_Jinkela_wire_9020),
        .dout(new_Jinkela_wire_9021)
    );

    bfr new_Jinkela_buffer_3687 (
        .din(new_Jinkela_wire_4880),
        .dout(new_Jinkela_wire_4881)
    );

    bfr new_Jinkela_buffer_7071 (
        .din(new_Jinkela_wire_8832),
        .dout(new_Jinkela_wire_8833)
    );

    bfr new_Jinkela_buffer_3639 (
        .din(new_Jinkela_wire_4820),
        .dout(new_Jinkela_wire_4821)
    );

    bfr new_Jinkela_buffer_7113 (
        .din(new_Jinkela_wire_8892),
        .dout(new_Jinkela_wire_8893)
    );

    bfr new_Jinkela_buffer_3778 (
        .din(new_Jinkela_wire_5001),
        .dout(new_Jinkela_wire_5002)
    );

    bfr new_Jinkela_buffer_7072 (
        .din(new_Jinkela_wire_8833),
        .dout(new_Jinkela_wire_8834)
    );

    bfr new_Jinkela_buffer_3640 (
        .din(new_Jinkela_wire_4821),
        .dout(new_Jinkela_wire_4822)
    );

    bfr new_Jinkela_buffer_7193 (
        .din(new_Jinkela_wire_8976),
        .dout(new_Jinkela_wire_8977)
    );

    bfr new_Jinkela_buffer_3688 (
        .din(new_Jinkela_wire_4881),
        .dout(new_Jinkela_wire_4882)
    );

    bfr new_Jinkela_buffer_7073 (
        .din(new_Jinkela_wire_8834),
        .dout(new_Jinkela_wire_8835)
    );

    bfr new_Jinkela_buffer_3641 (
        .din(new_Jinkela_wire_4822),
        .dout(new_Jinkela_wire_4823)
    );

    bfr new_Jinkela_buffer_7114 (
        .din(new_Jinkela_wire_8893),
        .dout(new_Jinkela_wire_8894)
    );

    bfr new_Jinkela_buffer_3719 (
        .din(new_Jinkela_wire_4930),
        .dout(new_Jinkela_wire_4931)
    );

    spl2 new_Jinkela_splitter_730 (
        .a(new_Jinkela_wire_8835),
        .b(new_Jinkela_wire_8836),
        .c(new_Jinkela_wire_8837)
    );

    spl2 new_Jinkela_splitter_440 (
        .a(new_Jinkela_wire_4823),
        .b(new_Jinkela_wire_4824),
        .c(new_Jinkela_wire_4825)
    );

    bfr new_Jinkela_buffer_7115 (
        .din(new_Jinkela_wire_8894),
        .dout(new_Jinkela_wire_8895)
    );

    bfr new_Jinkela_buffer_3689 (
        .din(new_Jinkela_wire_4882),
        .dout(new_Jinkela_wire_4883)
    );

    bfr new_Jinkela_buffer_7194 (
        .din(new_Jinkela_wire_8977),
        .dout(new_Jinkela_wire_8978)
    );

    bfr new_Jinkela_buffer_3690 (
        .din(new_Jinkela_wire_4883),
        .dout(new_Jinkela_wire_4884)
    );

    bfr new_Jinkela_buffer_7116 (
        .din(new_Jinkela_wire_8895),
        .dout(new_Jinkela_wire_8896)
    );

    bfr new_Jinkela_buffer_3720 (
        .din(new_Jinkela_wire_4931),
        .dout(new_Jinkela_wire_4932)
    );

    bfr new_Jinkela_buffer_3691 (
        .din(new_Jinkela_wire_4884),
        .dout(new_Jinkela_wire_4885)
    );

    bfr new_Jinkela_buffer_7117 (
        .din(new_Jinkela_wire_8896),
        .dout(new_Jinkela_wire_8897)
    );

    bfr new_Jinkela_buffer_3779 (
        .din(new_Jinkela_wire_5002),
        .dout(new_Jinkela_wire_5003)
    );

    bfr new_Jinkela_buffer_7195 (
        .din(new_Jinkela_wire_8978),
        .dout(new_Jinkela_wire_8979)
    );

    bfr new_Jinkela_buffer_3692 (
        .din(new_Jinkela_wire_4885),
        .dout(new_Jinkela_wire_4886)
    );

    bfr new_Jinkela_buffer_7118 (
        .din(new_Jinkela_wire_8897),
        .dout(new_Jinkela_wire_8898)
    );

    bfr new_Jinkela_buffer_3721 (
        .din(new_Jinkela_wire_4932),
        .dout(new_Jinkela_wire_4933)
    );

    bfr new_Jinkela_buffer_7230 (
        .din(new_Jinkela_wire_9021),
        .dout(new_Jinkela_wire_9022)
    );

    bfr new_Jinkela_buffer_3693 (
        .din(new_Jinkela_wire_4886),
        .dout(new_Jinkela_wire_4887)
    );

    bfr new_Jinkela_buffer_7119 (
        .din(new_Jinkela_wire_8898),
        .dout(new_Jinkela_wire_8899)
    );

    bfr new_Jinkela_buffer_3818 (
        .din(_0858_),
        .dout(new_Jinkela_wire_5050)
    );

    bfr new_Jinkela_buffer_7196 (
        .din(new_Jinkela_wire_8979),
        .dout(new_Jinkela_wire_8980)
    );

    bfr new_Jinkela_buffer_3694 (
        .din(new_Jinkela_wire_4887),
        .dout(new_Jinkela_wire_4888)
    );

    bfr new_Jinkela_buffer_7120 (
        .din(new_Jinkela_wire_8899),
        .dout(new_Jinkela_wire_8900)
    );

    bfr new_Jinkela_buffer_3722 (
        .din(new_Jinkela_wire_4933),
        .dout(new_Jinkela_wire_4934)
    );

    spl2 new_Jinkela_splitter_748 (
        .a(_0430_),
        .b(new_Jinkela_wire_9099),
        .c(new_Jinkela_wire_9100)
    );

    bfr new_Jinkela_buffer_3695 (
        .din(new_Jinkela_wire_4888),
        .dout(new_Jinkela_wire_4889)
    );

    spl2 new_Jinkela_splitter_747 (
        .a(_1814_),
        .b(new_Jinkela_wire_9097),
        .c(new_Jinkela_wire_9098)
    );

    bfr new_Jinkela_buffer_7121 (
        .din(new_Jinkela_wire_8900),
        .dout(new_Jinkela_wire_8901)
    );

    bfr new_Jinkela_buffer_3780 (
        .din(new_Jinkela_wire_5003),
        .dout(new_Jinkela_wire_5004)
    );

    bfr new_Jinkela_buffer_7197 (
        .din(new_Jinkela_wire_8980),
        .dout(new_Jinkela_wire_8981)
    );

    bfr new_Jinkela_buffer_3696 (
        .din(new_Jinkela_wire_4889),
        .dout(new_Jinkela_wire_4890)
    );

    bfr new_Jinkela_buffer_7122 (
        .din(new_Jinkela_wire_8901),
        .dout(new_Jinkela_wire_8902)
    );

    bfr new_Jinkela_buffer_3723 (
        .din(new_Jinkela_wire_4934),
        .dout(new_Jinkela_wire_4935)
    );

    bfr new_Jinkela_buffer_7231 (
        .din(new_Jinkela_wire_9022),
        .dout(new_Jinkela_wire_9023)
    );

    bfr new_Jinkela_buffer_3697 (
        .din(new_Jinkela_wire_4890),
        .dout(new_Jinkela_wire_4891)
    );

    bfr new_Jinkela_buffer_7123 (
        .din(new_Jinkela_wire_8902),
        .dout(new_Jinkela_wire_8903)
    );

    bfr new_Jinkela_buffer_3817 (
        .din(new_Jinkela_wire_5046),
        .dout(new_Jinkela_wire_5047)
    );

    bfr new_Jinkela_buffer_3819 (
        .din(_0161_),
        .dout(new_Jinkela_wire_5051)
    );

    bfr new_Jinkela_buffer_7198 (
        .din(new_Jinkela_wire_8981),
        .dout(new_Jinkela_wire_8982)
    );

    bfr new_Jinkela_buffer_3698 (
        .din(new_Jinkela_wire_4891),
        .dout(new_Jinkela_wire_4892)
    );

    bfr new_Jinkela_buffer_7124 (
        .din(new_Jinkela_wire_8903),
        .dout(new_Jinkela_wire_8904)
    );

    bfr new_Jinkela_buffer_3724 (
        .din(new_Jinkela_wire_4935),
        .dout(new_Jinkela_wire_4936)
    );

    spl2 new_Jinkela_splitter_749 (
        .a(_0583_),
        .b(new_Jinkela_wire_9101),
        .c(new_Jinkela_wire_9102)
    );

    bfr new_Jinkela_buffer_3699 (
        .din(new_Jinkela_wire_4892),
        .dout(new_Jinkela_wire_4893)
    );

    bfr new_Jinkela_buffer_7125 (
        .din(new_Jinkela_wire_8904),
        .dout(new_Jinkela_wire_8905)
    );

    bfr new_Jinkela_buffer_3781 (
        .din(new_Jinkela_wire_5004),
        .dout(new_Jinkela_wire_5005)
    );

    bfr new_Jinkela_buffer_7199 (
        .din(new_Jinkela_wire_8982),
        .dout(new_Jinkela_wire_8983)
    );

    bfr new_Jinkela_buffer_3700 (
        .din(new_Jinkela_wire_4893),
        .dout(new_Jinkela_wire_4894)
    );

    bfr new_Jinkela_buffer_7126 (
        .din(new_Jinkela_wire_8905),
        .dout(new_Jinkela_wire_8906)
    );

    bfr new_Jinkela_buffer_3725 (
        .din(new_Jinkela_wire_4936),
        .dout(new_Jinkela_wire_4937)
    );

    bfr new_Jinkela_buffer_7232 (
        .din(new_Jinkela_wire_9023),
        .dout(new_Jinkela_wire_9024)
    );

    spl2 new_Jinkela_splitter_446 (
        .a(new_Jinkela_wire_4894),
        .b(new_Jinkela_wire_4895),
        .c(new_Jinkela_wire_4896)
    );

    bfr new_Jinkela_buffer_10573 (
        .din(new_Jinkela_wire_12772),
        .dout(new_Jinkela_wire_12773)
    );

    bfr new_Jinkela_buffer_10645 (
        .din(new_Jinkela_wire_12846),
        .dout(new_Jinkela_wire_12847)
    );

    bfr new_Jinkela_buffer_10574 (
        .din(new_Jinkela_wire_12773),
        .dout(new_Jinkela_wire_12774)
    );

    spl2 new_Jinkela_splitter_956 (
        .a(_0867_),
        .b(new_Jinkela_wire_13047),
        .c(new_Jinkela_wire_13048)
    );

    bfr new_Jinkela_buffer_10575 (
        .din(new_Jinkela_wire_12774),
        .dout(new_Jinkela_wire_12775)
    );

    bfr new_Jinkela_buffer_10646 (
        .din(new_Jinkela_wire_12847),
        .dout(new_Jinkela_wire_12848)
    );

    bfr new_Jinkela_buffer_10576 (
        .din(new_Jinkela_wire_12775),
        .dout(new_Jinkela_wire_12776)
    );

    bfr new_Jinkela_buffer_10709 (
        .din(new_Jinkela_wire_12914),
        .dout(new_Jinkela_wire_12915)
    );

    bfr new_Jinkela_buffer_10577 (
        .din(new_Jinkela_wire_12776),
        .dout(new_Jinkela_wire_12777)
    );

    bfr new_Jinkela_buffer_10647 (
        .din(new_Jinkela_wire_12848),
        .dout(new_Jinkela_wire_12849)
    );

    bfr new_Jinkela_buffer_10578 (
        .din(new_Jinkela_wire_12777),
        .dout(new_Jinkela_wire_12778)
    );

    bfr new_Jinkela_buffer_10800 (
        .din(new_Jinkela_wire_13009),
        .dout(new_Jinkela_wire_13010)
    );

    bfr new_Jinkela_buffer_10579 (
        .din(new_Jinkela_wire_12778),
        .dout(new_Jinkela_wire_12779)
    );

    bfr new_Jinkela_buffer_10648 (
        .din(new_Jinkela_wire_12849),
        .dout(new_Jinkela_wire_12850)
    );

    bfr new_Jinkela_buffer_10580 (
        .din(new_Jinkela_wire_12779),
        .dout(new_Jinkela_wire_12780)
    );

    bfr new_Jinkela_buffer_10710 (
        .din(new_Jinkela_wire_12915),
        .dout(new_Jinkela_wire_12916)
    );

    bfr new_Jinkela_buffer_10581 (
        .din(new_Jinkela_wire_12780),
        .dout(new_Jinkela_wire_12781)
    );

    bfr new_Jinkela_buffer_10649 (
        .din(new_Jinkela_wire_12850),
        .dout(new_Jinkela_wire_12851)
    );

    bfr new_Jinkela_buffer_10582 (
        .din(new_Jinkela_wire_12781),
        .dout(new_Jinkela_wire_12782)
    );

    spl2 new_Jinkela_splitter_957 (
        .a(_1069_),
        .b(new_Jinkela_wire_13053),
        .c(new_Jinkela_wire_13054)
    );

    bfr new_Jinkela_buffer_10583 (
        .din(new_Jinkela_wire_12782),
        .dout(new_Jinkela_wire_12783)
    );

    bfr new_Jinkela_buffer_10650 (
        .din(new_Jinkela_wire_12851),
        .dout(new_Jinkela_wire_12852)
    );

    bfr new_Jinkela_buffer_10584 (
        .din(new_Jinkela_wire_12783),
        .dout(new_Jinkela_wire_12784)
    );

    bfr new_Jinkela_buffer_10711 (
        .din(new_Jinkela_wire_12916),
        .dout(new_Jinkela_wire_12917)
    );

    bfr new_Jinkela_buffer_10585 (
        .din(new_Jinkela_wire_12784),
        .dout(new_Jinkela_wire_12785)
    );

    bfr new_Jinkela_buffer_10651 (
        .din(new_Jinkela_wire_12852),
        .dout(new_Jinkela_wire_12853)
    );

    bfr new_Jinkela_buffer_10586 (
        .din(new_Jinkela_wire_12785),
        .dout(new_Jinkela_wire_12786)
    );

    bfr new_Jinkela_buffer_10804 (
        .din(new_Jinkela_wire_13015),
        .dout(new_Jinkela_wire_13016)
    );

    bfr new_Jinkela_buffer_10587 (
        .din(new_Jinkela_wire_12786),
        .dout(new_Jinkela_wire_12787)
    );

    bfr new_Jinkela_buffer_10652 (
        .din(new_Jinkela_wire_12853),
        .dout(new_Jinkela_wire_12854)
    );

    bfr new_Jinkela_buffer_10588 (
        .din(new_Jinkela_wire_12787),
        .dout(new_Jinkela_wire_12788)
    );

    bfr new_Jinkela_buffer_10712 (
        .din(new_Jinkela_wire_12917),
        .dout(new_Jinkela_wire_12918)
    );

    bfr new_Jinkela_buffer_10589 (
        .din(new_Jinkela_wire_12788),
        .dout(new_Jinkela_wire_12789)
    );

    bfr new_Jinkela_buffer_10653 (
        .din(new_Jinkela_wire_12854),
        .dout(new_Jinkela_wire_12855)
    );

    bfr new_Jinkela_buffer_10590 (
        .din(new_Jinkela_wire_12789),
        .dout(new_Jinkela_wire_12790)
    );

    bfr new_Jinkela_buffer_10833 (
        .din(new_Jinkela_wire_13048),
        .dout(new_Jinkela_wire_13049)
    );

    bfr new_Jinkela_buffer_10591 (
        .din(new_Jinkela_wire_12790),
        .dout(new_Jinkela_wire_12791)
    );

    bfr new_Jinkela_buffer_10654 (
        .din(new_Jinkela_wire_12855),
        .dout(new_Jinkela_wire_12856)
    );

    bfr new_Jinkela_buffer_10592 (
        .din(new_Jinkela_wire_12791),
        .dout(new_Jinkela_wire_12792)
    );

    bfr new_Jinkela_buffer_10713 (
        .din(new_Jinkela_wire_12918),
        .dout(new_Jinkela_wire_12919)
    );

    bfr new_Jinkela_buffer_10593 (
        .din(new_Jinkela_wire_12792),
        .dout(new_Jinkela_wire_12793)
    );

    bfr new_Jinkela_buffer_10655 (
        .din(new_Jinkela_wire_12856),
        .dout(new_Jinkela_wire_12857)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_17492 (
        .din(new_Jinkela_wire_20846),
        .dout(new_Jinkela_wire_20847)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_17421 (
        .din(new_Jinkela_wire_20769),
        .dout(new_Jinkela_wire_20770)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(_1261_),
        .b(new_Jinkela_wire_846),
        .c(new_Jinkela_wire_847)
    );

    spl2 new_Jinkela_splitter_194 (
        .a(_0863_),
        .b(new_Jinkela_wire_852),
        .c(new_Jinkela_wire_853)
    );

    spl2 new_Jinkela_splitter_1536 (
        .a(_1742_),
        .b(new_Jinkela_wire_21097),
        .c(new_Jinkela_wire_21098)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    bfr new_Jinkela_buffer_17721 (
        .din(_1345_),
        .dout(new_Jinkela_wire_21096)
    );

    bfr new_Jinkela_buffer_17422 (
        .din(new_Jinkela_wire_20770),
        .dout(new_Jinkela_wire_20771)
    );

    bfr new_Jinkela_buffer_17493 (
        .din(new_Jinkela_wire_20847),
        .dout(new_Jinkela_wire_20848)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    bfr new_Jinkela_buffer_17423 (
        .din(new_Jinkela_wire_20771),
        .dout(new_Jinkela_wire_20772)
    );

    spl2 new_Jinkela_splitter_195 (
        .a(_0891_),
        .b(new_Jinkela_wire_854),
        .c(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_17563 (
        .din(new_Jinkela_wire_20923),
        .dout(new_Jinkela_wire_20924)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_17424 (
        .din(new_Jinkela_wire_20772),
        .dout(new_Jinkela_wire_20773)
    );

    bfr new_Jinkela_buffer_17494 (
        .din(new_Jinkela_wire_20848),
        .dout(new_Jinkela_wire_20849)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_737),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_17425 (
        .din(new_Jinkela_wire_20773),
        .dout(new_Jinkela_wire_20774)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_17605 (
        .din(new_Jinkela_wire_20971),
        .dout(new_Jinkela_wire_20972)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_17426 (
        .din(new_Jinkela_wire_20774),
        .dout(new_Jinkela_wire_20775)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_net_3932),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_17495 (
        .din(new_Jinkela_wire_20849),
        .dout(new_Jinkela_wire_20850)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_739),
        .dout(new_Jinkela_wire_740)
    );

    bfr new_Jinkela_buffer_17427 (
        .din(new_Jinkela_wire_20775),
        .dout(new_Jinkela_wire_20776)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_17564 (
        .din(new_Jinkela_wire_20924),
        .dout(new_Jinkela_wire_20925)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_17428 (
        .din(new_Jinkela_wire_20776),
        .dout(new_Jinkela_wire_20777)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    bfr new_Jinkela_buffer_290 (
        .din(_1199_),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_17496 (
        .din(new_Jinkela_wire_20850),
        .dout(new_Jinkela_wire_20851)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_17429 (
        .din(new_Jinkela_wire_20777),
        .dout(new_Jinkela_wire_20778)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_17627 (
        .din(new_Jinkela_wire_20995),
        .dout(new_Jinkela_wire_20996)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_17430 (
        .din(new_Jinkela_wire_20778),
        .dout(new_Jinkela_wire_20779)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_17497 (
        .din(new_Jinkela_wire_20851),
        .dout(new_Jinkela_wire_20852)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_17431 (
        .din(new_Jinkela_wire_20779),
        .dout(new_Jinkela_wire_20780)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    bfr new_Jinkela_buffer_17565 (
        .din(new_Jinkela_wire_20925),
        .dout(new_Jinkela_wire_20926)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_17432 (
        .din(new_Jinkela_wire_20780),
        .dout(new_Jinkela_wire_20781)
    );

    bfr new_Jinkela_buffer_291 (
        .din(_1140_),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_17498 (
        .din(new_Jinkela_wire_20852),
        .dout(new_Jinkela_wire_20853)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_17433 (
        .din(new_Jinkela_wire_20781),
        .dout(new_Jinkela_wire_20782)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_17606 (
        .din(new_Jinkela_wire_20972),
        .dout(new_Jinkela_wire_20973)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_17434 (
        .din(new_Jinkela_wire_20782),
        .dout(new_Jinkela_wire_20783)
    );

    spl2 new_Jinkela_splitter_197 (
        .a(_1166_),
        .b(new_Jinkela_wire_1003),
        .c(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_17499 (
        .din(new_Jinkela_wire_20853),
        .dout(new_Jinkela_wire_20854)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_17435 (
        .din(new_Jinkela_wire_20783),
        .dout(new_Jinkela_wire_20784)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_17566 (
        .din(new_Jinkela_wire_20926),
        .dout(new_Jinkela_wire_20927)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    bfr new_Jinkela_buffer_17436 (
        .din(new_Jinkela_wire_20784),
        .dout(new_Jinkela_wire_20785)
    );

    bfr new_Jinkela_buffer_17500 (
        .din(new_Jinkela_wire_20854),
        .dout(new_Jinkela_wire_20855)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_17437 (
        .din(new_Jinkela_wire_20785),
        .dout(new_Jinkela_wire_20786)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_17438 (
        .din(new_Jinkela_wire_20786),
        .dout(new_Jinkela_wire_20787)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(_0271_),
        .b(new_Jinkela_wire_1009),
        .c(new_Jinkela_wire_1010)
    );

    bfr new_Jinkela_buffer_17501 (
        .din(new_Jinkela_wire_20855),
        .dout(new_Jinkela_wire_20856)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    bfr new_Jinkela_buffer_17439 (
        .din(new_Jinkela_wire_20787),
        .dout(new_Jinkela_wire_20788)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_17567 (
        .din(new_Jinkela_wire_20927),
        .dout(new_Jinkela_wire_20928)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_17440 (
        .din(new_Jinkela_wire_20788),
        .dout(new_Jinkela_wire_20789)
    );

    bfr new_Jinkela_buffer_17502 (
        .din(new_Jinkela_wire_20856),
        .dout(new_Jinkela_wire_20857)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_17441 (
        .din(new_Jinkela_wire_20789),
        .dout(new_Jinkela_wire_20790)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_10594 (
        .din(new_Jinkela_wire_12793),
        .dout(new_Jinkela_wire_12794)
    );

    bfr new_Jinkela_buffer_14195 (
        .din(_1138_),
        .dout(new_Jinkela_wire_16915)
    );

    bfr new_Jinkela_buffer_14191 (
        .din(new_Jinkela_wire_16910),
        .dout(new_Jinkela_wire_16911)
    );

    bfr new_Jinkela_buffer_10805 (
        .din(new_Jinkela_wire_13016),
        .dout(new_Jinkela_wire_13017)
    );

    bfr new_Jinkela_buffer_14057 (
        .din(new_Jinkela_wire_16744),
        .dout(new_Jinkela_wire_16745)
    );

    bfr new_Jinkela_buffer_10595 (
        .din(new_Jinkela_wire_12794),
        .dout(new_Jinkela_wire_12795)
    );

    bfr new_Jinkela_buffer_14109 (
        .din(new_Jinkela_wire_16812),
        .dout(new_Jinkela_wire_16813)
    );

    bfr new_Jinkela_buffer_10656 (
        .din(new_Jinkela_wire_12857),
        .dout(new_Jinkela_wire_12858)
    );

    bfr new_Jinkela_buffer_14058 (
        .din(new_Jinkela_wire_16745),
        .dout(new_Jinkela_wire_16746)
    );

    bfr new_Jinkela_buffer_10596 (
        .din(new_Jinkela_wire_12795),
        .dout(new_Jinkela_wire_12796)
    );

    bfr new_Jinkela_buffer_14165 (
        .din(new_Jinkela_wire_16878),
        .dout(new_Jinkela_wire_16879)
    );

    bfr new_Jinkela_buffer_10714 (
        .din(new_Jinkela_wire_12919),
        .dout(new_Jinkela_wire_12920)
    );

    bfr new_Jinkela_buffer_14059 (
        .din(new_Jinkela_wire_16746),
        .dout(new_Jinkela_wire_16747)
    );

    bfr new_Jinkela_buffer_10597 (
        .din(new_Jinkela_wire_12796),
        .dout(new_Jinkela_wire_12797)
    );

    bfr new_Jinkela_buffer_14110 (
        .din(new_Jinkela_wire_16813),
        .dout(new_Jinkela_wire_16814)
    );

    bfr new_Jinkela_buffer_10657 (
        .din(new_Jinkela_wire_12858),
        .dout(new_Jinkela_wire_12859)
    );

    bfr new_Jinkela_buffer_14060 (
        .din(new_Jinkela_wire_16747),
        .dout(new_Jinkela_wire_16748)
    );

    bfr new_Jinkela_buffer_10598 (
        .din(new_Jinkela_wire_12797),
        .dout(new_Jinkela_wire_12798)
    );

    bfr new_Jinkela_buffer_14061 (
        .din(new_Jinkela_wire_16748),
        .dout(new_Jinkela_wire_16749)
    );

    spl2 new_Jinkela_splitter_958 (
        .a(_1462_),
        .b(new_Jinkela_wire_13055),
        .c(new_Jinkela_wire_13056)
    );

    bfr new_Jinkela_buffer_10599 (
        .din(new_Jinkela_wire_12798),
        .dout(new_Jinkela_wire_12799)
    );

    bfr new_Jinkela_buffer_14111 (
        .din(new_Jinkela_wire_16814),
        .dout(new_Jinkela_wire_16815)
    );

    bfr new_Jinkela_buffer_10658 (
        .din(new_Jinkela_wire_12859),
        .dout(new_Jinkela_wire_12860)
    );

    bfr new_Jinkela_buffer_14062 (
        .din(new_Jinkela_wire_16749),
        .dout(new_Jinkela_wire_16750)
    );

    bfr new_Jinkela_buffer_10600 (
        .din(new_Jinkela_wire_12799),
        .dout(new_Jinkela_wire_12800)
    );

    bfr new_Jinkela_buffer_14166 (
        .din(new_Jinkela_wire_16879),
        .dout(new_Jinkela_wire_16880)
    );

    bfr new_Jinkela_buffer_10715 (
        .din(new_Jinkela_wire_12920),
        .dout(new_Jinkela_wire_12921)
    );

    bfr new_Jinkela_buffer_14063 (
        .din(new_Jinkela_wire_16750),
        .dout(new_Jinkela_wire_16751)
    );

    bfr new_Jinkela_buffer_10601 (
        .din(new_Jinkela_wire_12800),
        .dout(new_Jinkela_wire_12801)
    );

    bfr new_Jinkela_buffer_14112 (
        .din(new_Jinkela_wire_16815),
        .dout(new_Jinkela_wire_16816)
    );

    bfr new_Jinkela_buffer_10659 (
        .din(new_Jinkela_wire_12860),
        .dout(new_Jinkela_wire_12861)
    );

    bfr new_Jinkela_buffer_14064 (
        .din(new_Jinkela_wire_16751),
        .dout(new_Jinkela_wire_16752)
    );

    bfr new_Jinkela_buffer_10602 (
        .din(new_Jinkela_wire_12801),
        .dout(new_Jinkela_wire_12802)
    );

    spl2 new_Jinkela_splitter_1210 (
        .a(_0745_),
        .b(new_Jinkela_wire_16941),
        .c(new_Jinkela_wire_16942)
    );

    bfr new_Jinkela_buffer_10806 (
        .din(new_Jinkela_wire_13017),
        .dout(new_Jinkela_wire_13018)
    );

    bfr new_Jinkela_buffer_14065 (
        .din(new_Jinkela_wire_16752),
        .dout(new_Jinkela_wire_16753)
    );

    bfr new_Jinkela_buffer_10603 (
        .din(new_Jinkela_wire_12802),
        .dout(new_Jinkela_wire_12803)
    );

    bfr new_Jinkela_buffer_14113 (
        .din(new_Jinkela_wire_16816),
        .dout(new_Jinkela_wire_16817)
    );

    bfr new_Jinkela_buffer_10660 (
        .din(new_Jinkela_wire_12861),
        .dout(new_Jinkela_wire_12862)
    );

    bfr new_Jinkela_buffer_14066 (
        .din(new_Jinkela_wire_16753),
        .dout(new_Jinkela_wire_16754)
    );

    bfr new_Jinkela_buffer_10604 (
        .din(new_Jinkela_wire_12803),
        .dout(new_Jinkela_wire_12804)
    );

    bfr new_Jinkela_buffer_14167 (
        .din(new_Jinkela_wire_16880),
        .dout(new_Jinkela_wire_16881)
    );

    bfr new_Jinkela_buffer_10716 (
        .din(new_Jinkela_wire_12921),
        .dout(new_Jinkela_wire_12922)
    );

    bfr new_Jinkela_buffer_14067 (
        .din(new_Jinkela_wire_16754),
        .dout(new_Jinkela_wire_16755)
    );

    bfr new_Jinkela_buffer_10605 (
        .din(new_Jinkela_wire_12804),
        .dout(new_Jinkela_wire_12805)
    );

    bfr new_Jinkela_buffer_14114 (
        .din(new_Jinkela_wire_16817),
        .dout(new_Jinkela_wire_16818)
    );

    bfr new_Jinkela_buffer_10661 (
        .din(new_Jinkela_wire_12862),
        .dout(new_Jinkela_wire_12863)
    );

    bfr new_Jinkela_buffer_14068 (
        .din(new_Jinkela_wire_16755),
        .dout(new_Jinkela_wire_16756)
    );

    bfr new_Jinkela_buffer_10606 (
        .din(new_Jinkela_wire_12805),
        .dout(new_Jinkela_wire_12806)
    );

    spl2 new_Jinkela_splitter_1211 (
        .a(_0327_),
        .b(new_Jinkela_wire_16943),
        .c(new_Jinkela_wire_16944)
    );

    bfr new_Jinkela_buffer_10837 (
        .din(_1601_),
        .dout(new_Jinkela_wire_13057)
    );

    bfr new_Jinkela_buffer_14069 (
        .din(new_Jinkela_wire_16756),
        .dout(new_Jinkela_wire_16757)
    );

    bfr new_Jinkela_buffer_10607 (
        .din(new_Jinkela_wire_12806),
        .dout(new_Jinkela_wire_12807)
    );

    bfr new_Jinkela_buffer_14115 (
        .din(new_Jinkela_wire_16818),
        .dout(new_Jinkela_wire_16819)
    );

    bfr new_Jinkela_buffer_10662 (
        .din(new_Jinkela_wire_12863),
        .dout(new_Jinkela_wire_12864)
    );

    bfr new_Jinkela_buffer_14070 (
        .din(new_Jinkela_wire_16757),
        .dout(new_Jinkela_wire_16758)
    );

    bfr new_Jinkela_buffer_10608 (
        .din(new_Jinkela_wire_12807),
        .dout(new_Jinkela_wire_12808)
    );

    bfr new_Jinkela_buffer_14168 (
        .din(new_Jinkela_wire_16881),
        .dout(new_Jinkela_wire_16882)
    );

    bfr new_Jinkela_buffer_10717 (
        .din(new_Jinkela_wire_12922),
        .dout(new_Jinkela_wire_12923)
    );

    bfr new_Jinkela_buffer_14071 (
        .din(new_Jinkela_wire_16758),
        .dout(new_Jinkela_wire_16759)
    );

    bfr new_Jinkela_buffer_10609 (
        .din(new_Jinkela_wire_12808),
        .dout(new_Jinkela_wire_12809)
    );

    bfr new_Jinkela_buffer_14116 (
        .din(new_Jinkela_wire_16819),
        .dout(new_Jinkela_wire_16820)
    );

    bfr new_Jinkela_buffer_10663 (
        .din(new_Jinkela_wire_12864),
        .dout(new_Jinkela_wire_12865)
    );

    bfr new_Jinkela_buffer_14072 (
        .din(new_Jinkela_wire_16759),
        .dout(new_Jinkela_wire_16760)
    );

    bfr new_Jinkela_buffer_10610 (
        .din(new_Jinkela_wire_12809),
        .dout(new_Jinkela_wire_12810)
    );

    bfr new_Jinkela_buffer_14192 (
        .din(new_Jinkela_wire_16911),
        .dout(new_Jinkela_wire_16912)
    );

    bfr new_Jinkela_buffer_10807 (
        .din(new_Jinkela_wire_13018),
        .dout(new_Jinkela_wire_13019)
    );

    bfr new_Jinkela_buffer_14073 (
        .din(new_Jinkela_wire_16760),
        .dout(new_Jinkela_wire_16761)
    );

    bfr new_Jinkela_buffer_10611 (
        .din(new_Jinkela_wire_12810),
        .dout(new_Jinkela_wire_12811)
    );

    bfr new_Jinkela_buffer_14117 (
        .din(new_Jinkela_wire_16820),
        .dout(new_Jinkela_wire_16821)
    );

    bfr new_Jinkela_buffer_10664 (
        .din(new_Jinkela_wire_12865),
        .dout(new_Jinkela_wire_12866)
    );

    bfr new_Jinkela_buffer_14074 (
        .din(new_Jinkela_wire_16761),
        .dout(new_Jinkela_wire_16762)
    );

    bfr new_Jinkela_buffer_10612 (
        .din(new_Jinkela_wire_12811),
        .dout(new_Jinkela_wire_12812)
    );

    bfr new_Jinkela_buffer_14169 (
        .din(new_Jinkela_wire_16882),
        .dout(new_Jinkela_wire_16883)
    );

    bfr new_Jinkela_buffer_10718 (
        .din(new_Jinkela_wire_12923),
        .dout(new_Jinkela_wire_12924)
    );

    bfr new_Jinkela_buffer_14075 (
        .din(new_Jinkela_wire_16762),
        .dout(new_Jinkela_wire_16763)
    );

    bfr new_Jinkela_buffer_10613 (
        .din(new_Jinkela_wire_12812),
        .dout(new_Jinkela_wire_12813)
    );

    bfr new_Jinkela_buffer_14118 (
        .din(new_Jinkela_wire_16821),
        .dout(new_Jinkela_wire_16822)
    );

    bfr new_Jinkela_buffer_10665 (
        .din(new_Jinkela_wire_12866),
        .dout(new_Jinkela_wire_12867)
    );

    bfr new_Jinkela_buffer_14076 (
        .din(new_Jinkela_wire_16763),
        .dout(new_Jinkela_wire_16764)
    );

    bfr new_Jinkela_buffer_10614 (
        .din(new_Jinkela_wire_12813),
        .dout(new_Jinkela_wire_12814)
    );

    bfr new_Jinkela_buffer_14196 (
        .din(new_Jinkela_wire_16915),
        .dout(new_Jinkela_wire_16916)
    );

    bfr new_Jinkela_buffer_10834 (
        .din(new_Jinkela_wire_13049),
        .dout(new_Jinkela_wire_13050)
    );

    bfr new_Jinkela_buffer_14077 (
        .din(new_Jinkela_wire_16764),
        .dout(new_Jinkela_wire_16765)
    );

    bfr new_Jinkela_buffer_14119 (
        .din(new_Jinkela_wire_16822),
        .dout(new_Jinkela_wire_16823)
    );

    bfr new_Jinkela_buffer_14078 (
        .din(new_Jinkela_wire_16765),
        .dout(new_Jinkela_wire_16766)
    );

    bfr new_Jinkela_buffer_14170 (
        .din(new_Jinkela_wire_16883),
        .dout(new_Jinkela_wire_16884)
    );

    bfr new_Jinkela_buffer_14079 (
        .din(new_Jinkela_wire_16766),
        .dout(new_Jinkela_wire_16767)
    );

    bfr new_Jinkela_buffer_14120 (
        .din(new_Jinkela_wire_16823),
        .dout(new_Jinkela_wire_16824)
    );

    bfr new_Jinkela_buffer_14080 (
        .din(new_Jinkela_wire_16767),
        .dout(new_Jinkela_wire_16768)
    );

    bfr new_Jinkela_buffer_14193 (
        .din(new_Jinkela_wire_16912),
        .dout(new_Jinkela_wire_16913)
    );

    bfr new_Jinkela_buffer_14081 (
        .din(new_Jinkela_wire_16768),
        .dout(new_Jinkela_wire_16769)
    );

    bfr new_Jinkela_buffer_14121 (
        .din(new_Jinkela_wire_16824),
        .dout(new_Jinkela_wire_16825)
    );

    bfr new_Jinkela_buffer_14082 (
        .din(new_Jinkela_wire_16769),
        .dout(new_Jinkela_wire_16770)
    );

    bfr new_Jinkela_buffer_14171 (
        .din(new_Jinkela_wire_16884),
        .dout(new_Jinkela_wire_16885)
    );

    bfr new_Jinkela_buffer_14083 (
        .din(new_Jinkela_wire_16770),
        .dout(new_Jinkela_wire_16771)
    );

    bfr new_Jinkela_buffer_14122 (
        .din(new_Jinkela_wire_16825),
        .dout(new_Jinkela_wire_16826)
    );

    bfr new_Jinkela_buffer_14084 (
        .din(new_Jinkela_wire_16771),
        .dout(new_Jinkela_wire_16772)
    );

    bfr new_Jinkela_buffer_14085 (
        .din(new_Jinkela_wire_16772),
        .dout(new_Jinkela_wire_16773)
    );

    bfr new_Jinkela_buffer_14123 (
        .din(new_Jinkela_wire_16826),
        .dout(new_Jinkela_wire_16827)
    );

    spl2 new_Jinkela_splitter_1193 (
        .a(new_Jinkela_wire_16773),
        .b(new_Jinkela_wire_16774),
        .c(new_Jinkela_wire_16775)
    );

    bfr new_Jinkela_buffer_14124 (
        .din(new_Jinkela_wire_16827),
        .dout(new_Jinkela_wire_16828)
    );

    bfr new_Jinkela_buffer_14172 (
        .din(new_Jinkela_wire_16885),
        .dout(new_Jinkela_wire_16886)
    );

    bfr new_Jinkela_buffer_14194 (
        .din(new_Jinkela_wire_16913),
        .dout(new_Jinkela_wire_16914)
    );

    bfr new_Jinkela_buffer_14125 (
        .din(new_Jinkela_wire_16828),
        .dout(new_Jinkela_wire_16829)
    );

    bfr new_Jinkela_buffer_14173 (
        .din(new_Jinkela_wire_16886),
        .dout(new_Jinkela_wire_16887)
    );

    bfr new_Jinkela_buffer_14126 (
        .din(new_Jinkela_wire_16829),
        .dout(new_Jinkela_wire_16830)
    );

    bfr new_Jinkela_buffer_14197 (
        .din(new_Jinkela_wire_16916),
        .dout(new_Jinkela_wire_16917)
    );

    bfr new_Jinkela_buffer_14127 (
        .din(new_Jinkela_wire_16830),
        .dout(new_Jinkela_wire_16831)
    );

    bfr new_Jinkela_buffer_14174 (
        .din(new_Jinkela_wire_16887),
        .dout(new_Jinkela_wire_16888)
    );

    bfr new_Jinkela_buffer_14128 (
        .din(new_Jinkela_wire_16831),
        .dout(new_Jinkela_wire_16832)
    );

    spl2 new_Jinkela_splitter_1212 (
        .a(_0913_),
        .b(new_Jinkela_wire_16945),
        .c(new_Jinkela_wire_16946)
    );

    bfr new_Jinkela_buffer_14129 (
        .din(new_Jinkela_wire_16832),
        .dout(new_Jinkela_wire_16833)
    );

    bfr new_Jinkela_buffer_14175 (
        .din(new_Jinkela_wire_16888),
        .dout(new_Jinkela_wire_16889)
    );

    bfr new_Jinkela_buffer_14130 (
        .din(new_Jinkela_wire_16833),
        .dout(new_Jinkela_wire_16834)
    );

    bfr new_Jinkela_buffer_14198 (
        .din(new_Jinkela_wire_16917),
        .dout(new_Jinkela_wire_16918)
    );

    bfr new_Jinkela_buffer_14131 (
        .din(new_Jinkela_wire_16834),
        .dout(new_Jinkela_wire_16835)
    );

    bfr new_Jinkela_buffer_14176 (
        .din(new_Jinkela_wire_16889),
        .dout(new_Jinkela_wire_16890)
    );

    bfr new_Jinkela_buffer_14132 (
        .din(new_Jinkela_wire_16835),
        .dout(new_Jinkela_wire_16836)
    );

    spl2 new_Jinkela_splitter_1214 (
        .a(_1075_),
        .b(new_Jinkela_wire_16949),
        .c(new_Jinkela_wire_16950)
    );

    spl2 new_Jinkela_splitter_1213 (
        .a(_1701_),
        .b(new_Jinkela_wire_16947),
        .c(new_Jinkela_wire_16948)
    );

    bfr new_Jinkela_buffer_14133 (
        .din(new_Jinkela_wire_16836),
        .dout(new_Jinkela_wire_16837)
    );

    bfr new_Jinkela_buffer_14177 (
        .din(new_Jinkela_wire_16890),
        .dout(new_Jinkela_wire_16891)
    );

    bfr new_Jinkela_buffer_14134 (
        .din(new_Jinkela_wire_16837),
        .dout(new_Jinkela_wire_16838)
    );

    bfr new_Jinkela_buffer_14199 (
        .din(new_Jinkela_wire_16918),
        .dout(new_Jinkela_wire_16919)
    );

    bfr new_Jinkela_buffer_14135 (
        .din(new_Jinkela_wire_16838),
        .dout(new_Jinkela_wire_16839)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_7127 (
        .din(new_Jinkela_wire_8906),
        .dout(new_Jinkela_wire_8907)
    );

    bfr new_Jinkela_buffer_17608 (
        .din(new_Jinkela_wire_20974),
        .dout(new_Jinkela_wire_20975)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_7200 (
        .din(new_Jinkela_wire_8983),
        .dout(new_Jinkela_wire_8984)
    );

    bfr new_Jinkela_buffer_17442 (
        .din(new_Jinkela_wire_20790),
        .dout(new_Jinkela_wire_20791)
    );

    bfr new_Jinkela_buffer_7128 (
        .din(new_Jinkela_wire_8907),
        .dout(new_Jinkela_wire_8908)
    );

    bfr new_Jinkela_buffer_17503 (
        .din(new_Jinkela_wire_20857),
        .dout(new_Jinkela_wire_20858)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_17443 (
        .din(new_Jinkela_wire_20791),
        .dout(new_Jinkela_wire_20792)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_7129 (
        .din(new_Jinkela_wire_8908),
        .dout(new_Jinkela_wire_8909)
    );

    bfr new_Jinkela_buffer_17568 (
        .din(new_Jinkela_wire_20928),
        .dout(new_Jinkela_wire_20929)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_7201 (
        .din(new_Jinkela_wire_8984),
        .dout(new_Jinkela_wire_8985)
    );

    spl2 new_Jinkela_splitter_1523 (
        .a(new_Jinkela_wire_20792),
        .b(new_Jinkela_wire_20793),
        .c(new_Jinkela_wire_20794)
    );

    bfr new_Jinkela_buffer_7130 (
        .din(new_Jinkela_wire_8909),
        .dout(new_Jinkela_wire_8910)
    );

    spl2 new_Jinkela_splitter_1537 (
        .a(_1718_),
        .b(new_Jinkela_wire_21099),
        .c(new_Jinkela_wire_21100)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_7233 (
        .din(new_Jinkela_wire_9024),
        .dout(new_Jinkela_wire_9025)
    );

    bfr new_Jinkela_buffer_17504 (
        .din(new_Jinkela_wire_20858),
        .dout(new_Jinkela_wire_20859)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_7131 (
        .din(new_Jinkela_wire_8910),
        .dout(new_Jinkela_wire_8911)
    );

    bfr new_Jinkela_buffer_17505 (
        .din(new_Jinkela_wire_20859),
        .dout(new_Jinkela_wire_20860)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_7202 (
        .din(new_Jinkela_wire_8985),
        .dout(new_Jinkela_wire_8986)
    );

    bfr new_Jinkela_buffer_17569 (
        .din(new_Jinkela_wire_20929),
        .dout(new_Jinkela_wire_20930)
    );

    spl2 new_Jinkela_splitter_199 (
        .a(_0018_),
        .b(new_Jinkela_wire_1011),
        .c(new_Jinkela_wire_1012)
    );

    bfr new_Jinkela_buffer_7132 (
        .din(new_Jinkela_wire_8911),
        .dout(new_Jinkela_wire_8912)
    );

    bfr new_Jinkela_buffer_17506 (
        .din(new_Jinkela_wire_20860),
        .dout(new_Jinkela_wire_20861)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    bfr new_Jinkela_buffer_17609 (
        .din(new_Jinkela_wire_20975),
        .dout(new_Jinkela_wire_20976)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_7305 (
        .din(_1691_),
        .dout(new_Jinkela_wire_9107)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_7133 (
        .din(new_Jinkela_wire_8912),
        .dout(new_Jinkela_wire_8913)
    );

    bfr new_Jinkela_buffer_17507 (
        .din(new_Jinkela_wire_20861),
        .dout(new_Jinkela_wire_20862)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_7203 (
        .din(new_Jinkela_wire_8986),
        .dout(new_Jinkela_wire_8987)
    );

    bfr new_Jinkela_buffer_17570 (
        .din(new_Jinkela_wire_20930),
        .dout(new_Jinkela_wire_20931)
    );

    bfr new_Jinkela_buffer_7134 (
        .din(new_Jinkela_wire_8913),
        .dout(new_Jinkela_wire_8914)
    );

    bfr new_Jinkela_buffer_17508 (
        .din(new_Jinkela_wire_20862),
        .dout(new_Jinkela_wire_20863)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    bfr new_Jinkela_buffer_7234 (
        .din(new_Jinkela_wire_9025),
        .dout(new_Jinkela_wire_9026)
    );

    bfr new_Jinkela_buffer_17629 (
        .din(new_Jinkela_wire_20997),
        .dout(new_Jinkela_wire_20998)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_7135 (
        .din(new_Jinkela_wire_8914),
        .dout(new_Jinkela_wire_8915)
    );

    bfr new_Jinkela_buffer_17509 (
        .din(new_Jinkela_wire_20863),
        .dout(new_Jinkela_wire_20864)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_762),
        .dout(new_Jinkela_wire_763)
    );

    bfr new_Jinkela_buffer_7204 (
        .din(new_Jinkela_wire_8987),
        .dout(new_Jinkela_wire_8988)
    );

    bfr new_Jinkela_buffer_17571 (
        .din(new_Jinkela_wire_20931),
        .dout(new_Jinkela_wire_20932)
    );

    bfr new_Jinkela_buffer_7136 (
        .din(new_Jinkela_wire_8915),
        .dout(new_Jinkela_wire_8916)
    );

    bfr new_Jinkela_buffer_17510 (
        .din(new_Jinkela_wire_20864),
        .dout(new_Jinkela_wire_20865)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_763),
        .dout(new_Jinkela_wire_764)
    );

    bfr new_Jinkela_buffer_7301 (
        .din(new_Jinkela_wire_9102),
        .dout(new_Jinkela_wire_9103)
    );

    bfr new_Jinkela_buffer_17610 (
        .din(new_Jinkela_wire_20976),
        .dout(new_Jinkela_wire_20977)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    spl2 new_Jinkela_splitter_751 (
        .a(_0177_),
        .b(new_Jinkela_wire_9173),
        .c(new_Jinkela_wire_9174)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_7137 (
        .din(new_Jinkela_wire_8916),
        .dout(new_Jinkela_wire_8917)
    );

    bfr new_Jinkela_buffer_17511 (
        .din(new_Jinkela_wire_20865),
        .dout(new_Jinkela_wire_20866)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_764),
        .dout(new_Jinkela_wire_765)
    );

    bfr new_Jinkela_buffer_7205 (
        .din(new_Jinkela_wire_8988),
        .dout(new_Jinkela_wire_8989)
    );

    bfr new_Jinkela_buffer_17572 (
        .din(new_Jinkela_wire_20932),
        .dout(new_Jinkela_wire_20933)
    );

    bfr new_Jinkela_buffer_7138 (
        .din(new_Jinkela_wire_8917),
        .dout(new_Jinkela_wire_8918)
    );

    bfr new_Jinkela_buffer_17512 (
        .din(new_Jinkela_wire_20866),
        .dout(new_Jinkela_wire_20867)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_765),
        .dout(new_Jinkela_wire_766)
    );

    bfr new_Jinkela_buffer_7235 (
        .din(new_Jinkela_wire_9026),
        .dout(new_Jinkela_wire_9027)
    );

    bfr new_Jinkela_buffer_17722 (
        .din(new_Jinkela_wire_21100),
        .dout(new_Jinkela_wire_21101)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_7139 (
        .din(new_Jinkela_wire_8918),
        .dout(new_Jinkela_wire_8919)
    );

    bfr new_Jinkela_buffer_17513 (
        .din(new_Jinkela_wire_20867),
        .dout(new_Jinkela_wire_20868)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_7206 (
        .din(new_Jinkela_wire_8989),
        .dout(new_Jinkela_wire_8990)
    );

    bfr new_Jinkela_buffer_17573 (
        .din(new_Jinkela_wire_20933),
        .dout(new_Jinkela_wire_20934)
    );

    bfr new_Jinkela_buffer_7140 (
        .din(new_Jinkela_wire_8919),
        .dout(new_Jinkela_wire_8920)
    );

    bfr new_Jinkela_buffer_17514 (
        .din(new_Jinkela_wire_20868),
        .dout(new_Jinkela_wire_20869)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    bfr new_Jinkela_buffer_17611 (
        .din(new_Jinkela_wire_20977),
        .dout(new_Jinkela_wire_20978)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    spl2 new_Jinkela_splitter_752 (
        .a(_0047_),
        .b(new_Jinkela_wire_9175),
        .c(new_Jinkela_wire_9176)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_871),
        .dout(new_Jinkela_wire_872)
    );

    bfr new_Jinkela_buffer_7141 (
        .din(new_Jinkela_wire_8920),
        .dout(new_Jinkela_wire_8921)
    );

    bfr new_Jinkela_buffer_17515 (
        .din(new_Jinkela_wire_20869),
        .dout(new_Jinkela_wire_20870)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    bfr new_Jinkela_buffer_7207 (
        .din(new_Jinkela_wire_8990),
        .dout(new_Jinkela_wire_8991)
    );

    bfr new_Jinkela_buffer_17574 (
        .din(new_Jinkela_wire_20934),
        .dout(new_Jinkela_wire_20935)
    );

    bfr new_Jinkela_buffer_7142 (
        .din(new_Jinkela_wire_8921),
        .dout(new_Jinkela_wire_8922)
    );

    bfr new_Jinkela_buffer_17516 (
        .din(new_Jinkela_wire_20870),
        .dout(new_Jinkela_wire_20871)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_7236 (
        .din(new_Jinkela_wire_9027),
        .dout(new_Jinkela_wire_9028)
    );

    bfr new_Jinkela_buffer_17630 (
        .din(new_Jinkela_wire_20998),
        .dout(new_Jinkela_wire_20999)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_7143 (
        .din(new_Jinkela_wire_8922),
        .dout(new_Jinkela_wire_8923)
    );

    bfr new_Jinkela_buffer_17517 (
        .din(new_Jinkela_wire_20871),
        .dout(new_Jinkela_wire_20872)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_770),
        .dout(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_7208 (
        .din(new_Jinkela_wire_8991),
        .dout(new_Jinkela_wire_8992)
    );

    bfr new_Jinkela_buffer_17575 (
        .din(new_Jinkela_wire_20935),
        .dout(new_Jinkela_wire_20936)
    );

    bfr new_Jinkela_buffer_315 (
        .din(_0373_),
        .dout(new_Jinkela_wire_1017)
    );

    bfr new_Jinkela_buffer_7144 (
        .din(new_Jinkela_wire_8923),
        .dout(new_Jinkela_wire_8924)
    );

    bfr new_Jinkela_buffer_17518 (
        .din(new_Jinkela_wire_20872),
        .dout(new_Jinkela_wire_20873)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_7302 (
        .din(new_Jinkela_wire_9103),
        .dout(new_Jinkela_wire_9104)
    );

    bfr new_Jinkela_buffer_17612 (
        .din(new_Jinkela_wire_20978),
        .dout(new_Jinkela_wire_20979)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_7145 (
        .din(new_Jinkela_wire_8924),
        .dout(new_Jinkela_wire_8925)
    );

    bfr new_Jinkela_buffer_17519 (
        .din(new_Jinkela_wire_20873),
        .dout(new_Jinkela_wire_20874)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_7209 (
        .din(new_Jinkela_wire_8992),
        .dout(new_Jinkela_wire_8993)
    );

    bfr new_Jinkela_buffer_17576 (
        .din(new_Jinkela_wire_20936),
        .dout(new_Jinkela_wire_20937)
    );

    bfr new_Jinkela_buffer_7146 (
        .din(new_Jinkela_wire_8925),
        .dout(new_Jinkela_wire_8926)
    );

    bfr new_Jinkela_buffer_17520 (
        .din(new_Jinkela_wire_20874),
        .dout(new_Jinkela_wire_20875)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_773),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_7237 (
        .din(new_Jinkela_wire_9028),
        .dout(new_Jinkela_wire_9029)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_17726 (
        .din(_0954_),
        .dout(new_Jinkela_wire_21105)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_7147 (
        .din(new_Jinkela_wire_8926),
        .dout(new_Jinkela_wire_8927)
    );

    bfr new_Jinkela_buffer_17521 (
        .din(new_Jinkela_wire_20875),
        .dout(new_Jinkela_wire_20876)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    bfr new_Jinkela_buffer_7210 (
        .din(new_Jinkela_wire_8993),
        .dout(new_Jinkela_wire_8994)
    );

    bfr new_Jinkela_buffer_17577 (
        .din(new_Jinkela_wire_20937),
        .dout(new_Jinkela_wire_20938)
    );

    bfr new_Jinkela_buffer_10615 (
        .din(new_Jinkela_wire_12814),
        .dout(new_Jinkela_wire_12815)
    );

    bfr new_Jinkela_buffer_10666 (
        .din(new_Jinkela_wire_12867),
        .dout(new_Jinkela_wire_12868)
    );

    bfr new_Jinkela_buffer_10616 (
        .din(new_Jinkela_wire_12815),
        .dout(new_Jinkela_wire_12816)
    );

    bfr new_Jinkela_buffer_10719 (
        .din(new_Jinkela_wire_12924),
        .dout(new_Jinkela_wire_12925)
    );

    bfr new_Jinkela_buffer_10617 (
        .din(new_Jinkela_wire_12816),
        .dout(new_Jinkela_wire_12817)
    );

    bfr new_Jinkela_buffer_10667 (
        .din(new_Jinkela_wire_12868),
        .dout(new_Jinkela_wire_12869)
    );

    bfr new_Jinkela_buffer_10618 (
        .din(new_Jinkela_wire_12817),
        .dout(new_Jinkela_wire_12818)
    );

    bfr new_Jinkela_buffer_10808 (
        .din(new_Jinkela_wire_13019),
        .dout(new_Jinkela_wire_13020)
    );

    bfr new_Jinkela_buffer_10619 (
        .din(new_Jinkela_wire_12818),
        .dout(new_Jinkela_wire_12819)
    );

    bfr new_Jinkela_buffer_10668 (
        .din(new_Jinkela_wire_12869),
        .dout(new_Jinkela_wire_12870)
    );

    bfr new_Jinkela_buffer_10620 (
        .din(new_Jinkela_wire_12819),
        .dout(new_Jinkela_wire_12820)
    );

    bfr new_Jinkela_buffer_10720 (
        .din(new_Jinkela_wire_12925),
        .dout(new_Jinkela_wire_12926)
    );

    bfr new_Jinkela_buffer_10621 (
        .din(new_Jinkela_wire_12820),
        .dout(new_Jinkela_wire_12821)
    );

    bfr new_Jinkela_buffer_10669 (
        .din(new_Jinkela_wire_12870),
        .dout(new_Jinkela_wire_12871)
    );

    bfr new_Jinkela_buffer_10622 (
        .din(new_Jinkela_wire_12821),
        .dout(new_Jinkela_wire_12822)
    );

    spl2 new_Jinkela_splitter_960 (
        .a(_0626_),
        .b(new_Jinkela_wire_13060),
        .c(new_Jinkela_wire_13061)
    );

    bfr new_Jinkela_buffer_10623 (
        .din(new_Jinkela_wire_12822),
        .dout(new_Jinkela_wire_12823)
    );

    bfr new_Jinkela_buffer_10670 (
        .din(new_Jinkela_wire_12871),
        .dout(new_Jinkela_wire_12872)
    );

    bfr new_Jinkela_buffer_10624 (
        .din(new_Jinkela_wire_12823),
        .dout(new_Jinkela_wire_12824)
    );

    bfr new_Jinkela_buffer_10721 (
        .din(new_Jinkela_wire_12926),
        .dout(new_Jinkela_wire_12927)
    );

    bfr new_Jinkela_buffer_10625 (
        .din(new_Jinkela_wire_12824),
        .dout(new_Jinkela_wire_12825)
    );

    bfr new_Jinkela_buffer_10671 (
        .din(new_Jinkela_wire_12872),
        .dout(new_Jinkela_wire_12873)
    );

    bfr new_Jinkela_buffer_10626 (
        .din(new_Jinkela_wire_12825),
        .dout(new_Jinkela_wire_12826)
    );

    bfr new_Jinkela_buffer_10809 (
        .din(new_Jinkela_wire_13020),
        .dout(new_Jinkela_wire_13021)
    );

    bfr new_Jinkela_buffer_10627 (
        .din(new_Jinkela_wire_12826),
        .dout(new_Jinkela_wire_12827)
    );

    bfr new_Jinkela_buffer_10672 (
        .din(new_Jinkela_wire_12873),
        .dout(new_Jinkela_wire_12874)
    );

    bfr new_Jinkela_buffer_10628 (
        .din(new_Jinkela_wire_12827),
        .dout(new_Jinkela_wire_12828)
    );

    bfr new_Jinkela_buffer_10722 (
        .din(new_Jinkela_wire_12927),
        .dout(new_Jinkela_wire_12928)
    );

    spl2 new_Jinkela_splitter_949 (
        .a(new_Jinkela_wire_12828),
        .b(new_Jinkela_wire_12829),
        .c(new_Jinkela_wire_12830)
    );

    bfr new_Jinkela_buffer_10835 (
        .din(new_Jinkela_wire_13050),
        .dout(new_Jinkela_wire_13051)
    );

    bfr new_Jinkela_buffer_10673 (
        .din(new_Jinkela_wire_12874),
        .dout(new_Jinkela_wire_12875)
    );

    bfr new_Jinkela_buffer_10674 (
        .din(new_Jinkela_wire_12875),
        .dout(new_Jinkela_wire_12876)
    );

    bfr new_Jinkela_buffer_10723 (
        .din(new_Jinkela_wire_12928),
        .dout(new_Jinkela_wire_12929)
    );

    bfr new_Jinkela_buffer_10675 (
        .din(new_Jinkela_wire_12876),
        .dout(new_Jinkela_wire_12877)
    );

    bfr new_Jinkela_buffer_10810 (
        .din(new_Jinkela_wire_13021),
        .dout(new_Jinkela_wire_13022)
    );

    bfr new_Jinkela_buffer_10676 (
        .din(new_Jinkela_wire_12877),
        .dout(new_Jinkela_wire_12878)
    );

    bfr new_Jinkela_buffer_10724 (
        .din(new_Jinkela_wire_12929),
        .dout(new_Jinkela_wire_12930)
    );

    bfr new_Jinkela_buffer_10677 (
        .din(new_Jinkela_wire_12878),
        .dout(new_Jinkela_wire_12879)
    );

    spl2 new_Jinkela_splitter_959 (
        .a(_1362_),
        .b(new_Jinkela_wire_13058),
        .c(new_Jinkela_wire_13059)
    );

    bfr new_Jinkela_buffer_10678 (
        .din(new_Jinkela_wire_12879),
        .dout(new_Jinkela_wire_12880)
    );

    bfr new_Jinkela_buffer_10725 (
        .din(new_Jinkela_wire_12930),
        .dout(new_Jinkela_wire_12931)
    );

    bfr new_Jinkela_buffer_10679 (
        .din(new_Jinkela_wire_12880),
        .dout(new_Jinkela_wire_12881)
    );

    bfr new_Jinkela_buffer_7148 (
        .din(new_Jinkela_wire_8927),
        .dout(new_Jinkela_wire_8928)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_775),
        .dout(new_Jinkela_wire_776)
    );

    spl2 new_Jinkela_splitter_465 (
        .a(_0202_),
        .b(new_Jinkela_wire_5052),
        .c(new_Jinkela_wire_5053)
    );

    bfr new_Jinkela_buffer_3726 (
        .din(new_Jinkela_wire_4937),
        .dout(new_Jinkela_wire_4938)
    );

    bfr new_Jinkela_buffer_7306 (
        .din(new_Jinkela_wire_9107),
        .dout(new_Jinkela_wire_9108)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_991),
        .dout(new_Jinkela_wire_992)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_3782 (
        .din(new_Jinkela_wire_5005),
        .dout(new_Jinkela_wire_5006)
    );

    bfr new_Jinkela_buffer_7149 (
        .din(new_Jinkela_wire_8928),
        .dout(new_Jinkela_wire_8929)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_776),
        .dout(new_Jinkela_wire_777)
    );

    bfr new_Jinkela_buffer_3727 (
        .din(new_Jinkela_wire_4938),
        .dout(new_Jinkela_wire_4939)
    );

    bfr new_Jinkela_buffer_7211 (
        .din(new_Jinkela_wire_8994),
        .dout(new_Jinkela_wire_8995)
    );

    spl2 new_Jinkela_splitter_466 (
        .a(_0874_),
        .b(new_Jinkela_wire_5054),
        .c(new_Jinkela_wire_5055)
    );

    bfr new_Jinkela_buffer_7150 (
        .din(new_Jinkela_wire_8929),
        .dout(new_Jinkela_wire_8930)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_777),
        .dout(new_Jinkela_wire_778)
    );

    spl2 new_Jinkela_splitter_464 (
        .a(new_Jinkela_wire_5047),
        .b(new_Jinkela_wire_5048),
        .c(new_Jinkela_wire_5049)
    );

    bfr new_Jinkela_buffer_3728 (
        .din(new_Jinkela_wire_4939),
        .dout(new_Jinkela_wire_4940)
    );

    bfr new_Jinkela_buffer_7238 (
        .din(new_Jinkela_wire_9029),
        .dout(new_Jinkela_wire_9030)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_876),
        .dout(new_Jinkela_wire_877)
    );

    bfr new_Jinkela_buffer_3783 (
        .din(new_Jinkela_wire_5006),
        .dout(new_Jinkela_wire_5007)
    );

    bfr new_Jinkela_buffer_7151 (
        .din(new_Jinkela_wire_8930),
        .dout(new_Jinkela_wire_8931)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_778),
        .dout(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_3729 (
        .din(new_Jinkela_wire_4940),
        .dout(new_Jinkela_wire_4941)
    );

    bfr new_Jinkela_buffer_7212 (
        .din(new_Jinkela_wire_8995),
        .dout(new_Jinkela_wire_8996)
    );

    bfr new_Jinkela_buffer_316 (
        .din(_0984_),
        .dout(new_Jinkela_wire_1018)
    );

    bfr new_Jinkela_buffer_7152 (
        .din(new_Jinkela_wire_8931),
        .dout(new_Jinkela_wire_8932)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_779),
        .dout(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_3730 (
        .din(new_Jinkela_wire_4941),
        .dout(new_Jinkela_wire_4942)
    );

    bfr new_Jinkela_buffer_7303 (
        .din(new_Jinkela_wire_9104),
        .dout(new_Jinkela_wire_9105)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_877),
        .dout(new_Jinkela_wire_878)
    );

    bfr new_Jinkela_buffer_3784 (
        .din(new_Jinkela_wire_5007),
        .dout(new_Jinkela_wire_5008)
    );

    bfr new_Jinkela_buffer_7153 (
        .din(new_Jinkela_wire_8932),
        .dout(new_Jinkela_wire_8933)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_3731 (
        .din(new_Jinkela_wire_4942),
        .dout(new_Jinkela_wire_4943)
    );

    bfr new_Jinkela_buffer_7213 (
        .din(new_Jinkela_wire_8996),
        .dout(new_Jinkela_wire_8997)
    );

    bfr new_Jinkela_buffer_7154 (
        .din(new_Jinkela_wire_8933),
        .dout(new_Jinkela_wire_8934)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_3732 (
        .din(new_Jinkela_wire_4943),
        .dout(new_Jinkela_wire_4944)
    );

    bfr new_Jinkela_buffer_7239 (
        .din(new_Jinkela_wire_9030),
        .dout(new_Jinkela_wire_9031)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_878),
        .dout(new_Jinkela_wire_879)
    );

    bfr new_Jinkela_buffer_3785 (
        .din(new_Jinkela_wire_5008),
        .dout(new_Jinkela_wire_5009)
    );

    bfr new_Jinkela_buffer_7155 (
        .din(new_Jinkela_wire_8934),
        .dout(new_Jinkela_wire_8935)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_3733 (
        .din(new_Jinkela_wire_4944),
        .dout(new_Jinkela_wire_4945)
    );

    bfr new_Jinkela_buffer_7214 (
        .din(new_Jinkela_wire_8997),
        .dout(new_Jinkela_wire_8998)
    );

    bfr new_Jinkela_buffer_7156 (
        .din(new_Jinkela_wire_8935),
        .dout(new_Jinkela_wire_8936)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    spl2 new_Jinkela_splitter_467 (
        .a(_1672_),
        .b(new_Jinkela_wire_5092),
        .c(new_Jinkela_wire_5093)
    );

    bfr new_Jinkela_buffer_3734 (
        .din(new_Jinkela_wire_4945),
        .dout(new_Jinkela_wire_4946)
    );

    bfr new_Jinkela_buffer_7369 (
        .din(_0251_),
        .dout(new_Jinkela_wire_9179)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_879),
        .dout(new_Jinkela_wire_880)
    );

    bfr new_Jinkela_buffer_3786 (
        .din(new_Jinkela_wire_5009),
        .dout(new_Jinkela_wire_5010)
    );

    bfr new_Jinkela_buffer_7157 (
        .din(new_Jinkela_wire_8936),
        .dout(new_Jinkela_wire_8937)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_3735 (
        .din(new_Jinkela_wire_4946),
        .dout(new_Jinkela_wire_4947)
    );

    bfr new_Jinkela_buffer_7215 (
        .din(new_Jinkela_wire_8998),
        .dout(new_Jinkela_wire_8999)
    );

    bfr new_Jinkela_buffer_3820 (
        .din(new_Jinkela_wire_5055),
        .dout(new_Jinkela_wire_5056)
    );

    bfr new_Jinkela_buffer_7158 (
        .din(new_Jinkela_wire_8937),
        .dout(new_Jinkela_wire_8938)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_785),
        .dout(new_Jinkela_wire_786)
    );

    spl2 new_Jinkela_splitter_468 (
        .a(_1094_),
        .b(new_Jinkela_wire_5098),
        .c(new_Jinkela_wire_5099)
    );

    bfr new_Jinkela_buffer_3736 (
        .din(new_Jinkela_wire_4947),
        .dout(new_Jinkela_wire_4948)
    );

    bfr new_Jinkela_buffer_7240 (
        .din(new_Jinkela_wire_9031),
        .dout(new_Jinkela_wire_9032)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_3787 (
        .din(new_Jinkela_wire_5010),
        .dout(new_Jinkela_wire_5011)
    );

    bfr new_Jinkela_buffer_7159 (
        .din(new_Jinkela_wire_8938),
        .dout(new_Jinkela_wire_8939)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_3737 (
        .din(new_Jinkela_wire_4948),
        .dout(new_Jinkela_wire_4949)
    );

    bfr new_Jinkela_buffer_7216 (
        .din(new_Jinkela_wire_8999),
        .dout(new_Jinkela_wire_9000)
    );

    bfr new_Jinkela_buffer_317 (
        .din(_1817_),
        .dout(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_7160 (
        .din(new_Jinkela_wire_8939),
        .dout(new_Jinkela_wire_8940)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_787),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_3738 (
        .din(new_Jinkela_wire_4949),
        .dout(new_Jinkela_wire_4950)
    );

    bfr new_Jinkela_buffer_7304 (
        .din(new_Jinkela_wire_9105),
        .dout(new_Jinkela_wire_9106)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_994),
        .dout(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_3788 (
        .din(new_Jinkela_wire_5011),
        .dout(new_Jinkela_wire_5012)
    );

    bfr new_Jinkela_buffer_7161 (
        .din(new_Jinkela_wire_8940),
        .dout(new_Jinkela_wire_8941)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_3739 (
        .din(new_Jinkela_wire_4950),
        .dout(new_Jinkela_wire_4951)
    );

    bfr new_Jinkela_buffer_7217 (
        .din(new_Jinkela_wire_9000),
        .dout(new_Jinkela_wire_9001)
    );

    bfr new_Jinkela_buffer_3821 (
        .din(new_Jinkela_wire_5056),
        .dout(new_Jinkela_wire_5057)
    );

    bfr new_Jinkela_buffer_7162 (
        .din(new_Jinkela_wire_8941),
        .dout(new_Jinkela_wire_8942)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_3740 (
        .din(new_Jinkela_wire_4951),
        .dout(new_Jinkela_wire_4952)
    );

    bfr new_Jinkela_buffer_7241 (
        .din(new_Jinkela_wire_9032),
        .dout(new_Jinkela_wire_9033)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_1013),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    bfr new_Jinkela_buffer_3789 (
        .din(new_Jinkela_wire_5012),
        .dout(new_Jinkela_wire_5013)
    );

    bfr new_Jinkela_buffer_7163 (
        .din(new_Jinkela_wire_8942),
        .dout(new_Jinkela_wire_8943)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_3741 (
        .din(new_Jinkela_wire_4952),
        .dout(new_Jinkela_wire_4953)
    );

    bfr new_Jinkela_buffer_7218 (
        .din(new_Jinkela_wire_9001),
        .dout(new_Jinkela_wire_9002)
    );

    bfr new_Jinkela_buffer_3856 (
        .din(new_Jinkela_wire_5093),
        .dout(new_Jinkela_wire_5094)
    );

    bfr new_Jinkela_buffer_7164 (
        .din(new_Jinkela_wire_8943),
        .dout(new_Jinkela_wire_8944)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_791),
        .dout(new_Jinkela_wire_792)
    );

    spl2 new_Jinkela_splitter_469 (
        .a(_1392_),
        .b(new_Jinkela_wire_5104),
        .c(new_Jinkela_wire_5105)
    );

    bfr new_Jinkela_buffer_3742 (
        .din(new_Jinkela_wire_4953),
        .dout(new_Jinkela_wire_4954)
    );

    bfr new_Jinkela_buffer_7307 (
        .din(new_Jinkela_wire_9108),
        .dout(new_Jinkela_wire_9109)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    bfr new_Jinkela_buffer_3790 (
        .din(new_Jinkela_wire_5013),
        .dout(new_Jinkela_wire_5014)
    );

    bfr new_Jinkela_buffer_7165 (
        .din(new_Jinkela_wire_8944),
        .dout(new_Jinkela_wire_8945)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    bfr new_Jinkela_buffer_3743 (
        .din(new_Jinkela_wire_4954),
        .dout(new_Jinkela_wire_4955)
    );

    bfr new_Jinkela_buffer_7219 (
        .din(new_Jinkela_wire_9002),
        .dout(new_Jinkela_wire_9003)
    );

    bfr new_Jinkela_buffer_3822 (
        .din(new_Jinkela_wire_5057),
        .dout(new_Jinkela_wire_5058)
    );

    bfr new_Jinkela_buffer_7166 (
        .din(new_Jinkela_wire_8945),
        .dout(new_Jinkela_wire_8946)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_3744 (
        .din(new_Jinkela_wire_4955),
        .dout(new_Jinkela_wire_4956)
    );

    bfr new_Jinkela_buffer_7242 (
        .din(new_Jinkela_wire_9033),
        .dout(new_Jinkela_wire_9034)
    );

    bfr new_Jinkela_buffer_373 (
        .din(_0792_),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    bfr new_Jinkela_buffer_3791 (
        .din(new_Jinkela_wire_5014),
        .dout(new_Jinkela_wire_5015)
    );

    bfr new_Jinkela_buffer_7167 (
        .din(new_Jinkela_wire_8946),
        .dout(new_Jinkela_wire_8947)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    bfr new_Jinkela_buffer_3745 (
        .din(new_Jinkela_wire_4956),
        .dout(new_Jinkela_wire_4957)
    );

    bfr new_Jinkela_buffer_7220 (
        .din(new_Jinkela_wire_9003),
        .dout(new_Jinkela_wire_9004)
    );

    bfr new_Jinkela_buffer_7168 (
        .din(new_Jinkela_wire_8947),
        .dout(new_Jinkela_wire_8948)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    bfr new_Jinkela_buffer_3860 (
        .din(new_Jinkela_wire_5099),
        .dout(new_Jinkela_wire_5100)
    );

    bfr new_Jinkela_buffer_3746 (
        .din(new_Jinkela_wire_4957),
        .dout(new_Jinkela_wire_4958)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    spl2 new_Jinkela_splitter_753 (
        .a(_1307_),
        .b(new_Jinkela_wire_9177),
        .c(new_Jinkela_wire_9178)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_3792 (
        .din(new_Jinkela_wire_5015),
        .dout(new_Jinkela_wire_5016)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_3747 (
        .din(new_Jinkela_wire_4958),
        .dout(new_Jinkela_wire_4959)
    );

    bfr new_Jinkela_buffer_3823 (
        .din(new_Jinkela_wire_5058),
        .dout(new_Jinkela_wire_5059)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_3748 (
        .din(new_Jinkela_wire_4959),
        .dout(new_Jinkela_wire_4960)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    bfr new_Jinkela_buffer_3793 (
        .din(new_Jinkela_wire_5016),
        .dout(new_Jinkela_wire_5017)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_3749 (
        .din(new_Jinkela_wire_4960),
        .dout(new_Jinkela_wire_4961)
    );

    bfr new_Jinkela_buffer_3857 (
        .din(new_Jinkela_wire_5094),
        .dout(new_Jinkela_wire_5095)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    bfr new_Jinkela_buffer_3750 (
        .din(new_Jinkela_wire_4961),
        .dout(new_Jinkela_wire_4962)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_887),
        .dout(new_Jinkela_wire_888)
    );

    bfr new_Jinkela_buffer_3794 (
        .din(new_Jinkela_wire_5017),
        .dout(new_Jinkela_wire_5018)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_3751 (
        .din(new_Jinkela_wire_4962),
        .dout(new_Jinkela_wire_4963)
    );

    bfr new_Jinkela_buffer_3824 (
        .din(new_Jinkela_wire_5059),
        .dout(new_Jinkela_wire_5060)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    bfr new_Jinkela_buffer_3752 (
        .din(new_Jinkela_wire_4963),
        .dout(new_Jinkela_wire_4964)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_888),
        .dout(new_Jinkela_wire_889)
    );

    bfr new_Jinkela_buffer_3795 (
        .din(new_Jinkela_wire_5018),
        .dout(new_Jinkela_wire_5019)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_3753 (
        .din(new_Jinkela_wire_4964),
        .dout(new_Jinkela_wire_4965)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_net_3940),
        .dout(new_Jinkela_wire_1078)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_803),
        .dout(new_Jinkela_wire_804)
    );

    spl2 new_Jinkela_splitter_470 (
        .a(_1719_),
        .b(new_Jinkela_wire_5106),
        .c(new_Jinkela_wire_5107)
    );

    bfr new_Jinkela_buffer_3754 (
        .din(new_Jinkela_wire_4965),
        .dout(new_Jinkela_wire_4966)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_889),
        .dout(new_Jinkela_wire_890)
    );

    bfr new_Jinkela_buffer_3796 (
        .din(new_Jinkela_wire_5019),
        .dout(new_Jinkela_wire_5020)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_804),
        .dout(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_3755 (
        .din(new_Jinkela_wire_4966),
        .dout(new_Jinkela_wire_4967)
    );

    bfr new_Jinkela_buffer_3825 (
        .din(new_Jinkela_wire_5060),
        .dout(new_Jinkela_wire_5061)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_3756 (
        .din(new_Jinkela_wire_4967),
        .dout(new_Jinkela_wire_4968)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_3797 (
        .din(new_Jinkela_wire_5020),
        .dout(new_Jinkela_wire_5021)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_3757 (
        .din(new_Jinkela_wire_4968),
        .dout(new_Jinkela_wire_4969)
    );

    bfr new_Jinkela_buffer_3858 (
        .din(new_Jinkela_wire_5095),
        .dout(new_Jinkela_wire_5096)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_3758 (
        .din(new_Jinkela_wire_4969),
        .dout(new_Jinkela_wire_4970)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_891),
        .dout(new_Jinkela_wire_892)
    );

    bfr new_Jinkela_buffer_3798 (
        .din(new_Jinkela_wire_5021),
        .dout(new_Jinkela_wire_5022)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    bfr new_Jinkela_buffer_3759 (
        .din(new_Jinkela_wire_4970),
        .dout(new_Jinkela_wire_4971)
    );

    bfr new_Jinkela_buffer_3826 (
        .din(new_Jinkela_wire_5061),
        .dout(new_Jinkela_wire_5062)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_3760 (
        .din(new_Jinkela_wire_4971),
        .dout(new_Jinkela_wire_4972)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_3799 (
        .din(new_Jinkela_wire_5022),
        .dout(new_Jinkela_wire_5023)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    bfr new_Jinkela_buffer_3761 (
        .din(new_Jinkela_wire_4972),
        .dout(new_Jinkela_wire_4973)
    );

    bfr new_Jinkela_buffer_3864 (
        .din(_1379_),
        .dout(new_Jinkela_wire_5108)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_3762 (
        .din(new_Jinkela_wire_4973),
        .dout(new_Jinkela_wire_4974)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(new_Jinkela_wire_1000),
        .b(new_Jinkela_wire_1001),
        .c(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_3800 (
        .din(new_Jinkela_wire_5023),
        .dout(new_Jinkela_wire_5024)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_3763 (
        .din(new_Jinkela_wire_4974),
        .dout(new_Jinkela_wire_4975)
    );

    bfr new_Jinkela_buffer_3827 (
        .din(new_Jinkela_wire_5062),
        .dout(new_Jinkela_wire_5063)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_3764 (
        .din(new_Jinkela_wire_4975),
        .dout(new_Jinkela_wire_4976)
    );

    spl2 new_Jinkela_splitter_201 (
        .a(_1747_),
        .b(new_Jinkela_wire_1134),
        .c(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_3801 (
        .din(new_Jinkela_wire_5024),
        .dout(new_Jinkela_wire_5025)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_3765 (
        .din(new_Jinkela_wire_4976),
        .dout(new_Jinkela_wire_4977)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    bfr new_Jinkela_buffer_3859 (
        .din(new_Jinkela_wire_5096),
        .dout(new_Jinkela_wire_5097)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    bfr new_Jinkela_buffer_3766 (
        .din(new_Jinkela_wire_4977),
        .dout(new_Jinkela_wire_4978)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_3802 (
        .din(new_Jinkela_wire_5025),
        .dout(new_Jinkela_wire_5026)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_3767 (
        .din(new_Jinkela_wire_4978),
        .dout(new_Jinkela_wire_4979)
    );

    bfr new_Jinkela_buffer_14178 (
        .din(new_Jinkela_wire_16891),
        .dout(new_Jinkela_wire_16892)
    );

    bfr new_Jinkela_buffer_14136 (
        .din(new_Jinkela_wire_16839),
        .dout(new_Jinkela_wire_16840)
    );

    bfr new_Jinkela_buffer_14137 (
        .din(new_Jinkela_wire_16840),
        .dout(new_Jinkela_wire_16841)
    );

    bfr new_Jinkela_buffer_14179 (
        .din(new_Jinkela_wire_16892),
        .dout(new_Jinkela_wire_16893)
    );

    bfr new_Jinkela_buffer_14138 (
        .din(new_Jinkela_wire_16841),
        .dout(new_Jinkela_wire_16842)
    );

    bfr new_Jinkela_buffer_14200 (
        .din(new_Jinkela_wire_16919),
        .dout(new_Jinkela_wire_16920)
    );

    bfr new_Jinkela_buffer_14139 (
        .din(new_Jinkela_wire_16842),
        .dout(new_Jinkela_wire_16843)
    );

    bfr new_Jinkela_buffer_14180 (
        .din(new_Jinkela_wire_16893),
        .dout(new_Jinkela_wire_16894)
    );

    bfr new_Jinkela_buffer_14140 (
        .din(new_Jinkela_wire_16843),
        .dout(new_Jinkela_wire_16844)
    );

    spl2 new_Jinkela_splitter_1215 (
        .a(_1576_),
        .b(new_Jinkela_wire_16951),
        .c(new_Jinkela_wire_16952)
    );

    bfr new_Jinkela_buffer_14141 (
        .din(new_Jinkela_wire_16844),
        .dout(new_Jinkela_wire_16845)
    );

    bfr new_Jinkela_buffer_14181 (
        .din(new_Jinkela_wire_16894),
        .dout(new_Jinkela_wire_16895)
    );

    bfr new_Jinkela_buffer_14142 (
        .din(new_Jinkela_wire_16845),
        .dout(new_Jinkela_wire_16846)
    );

    bfr new_Jinkela_buffer_14201 (
        .din(new_Jinkela_wire_16920),
        .dout(new_Jinkela_wire_16921)
    );

    bfr new_Jinkela_buffer_14143 (
        .din(new_Jinkela_wire_16846),
        .dout(new_Jinkela_wire_16847)
    );

    bfr new_Jinkela_buffer_14182 (
        .din(new_Jinkela_wire_16895),
        .dout(new_Jinkela_wire_16896)
    );

    bfr new_Jinkela_buffer_14144 (
        .din(new_Jinkela_wire_16847),
        .dout(new_Jinkela_wire_16848)
    );

    spl2 new_Jinkela_splitter_1216 (
        .a(_0107_),
        .b(new_Jinkela_wire_16953),
        .c(new_Jinkela_wire_16954)
    );

    bfr new_Jinkela_buffer_14145 (
        .din(new_Jinkela_wire_16848),
        .dout(new_Jinkela_wire_16849)
    );

    bfr new_Jinkela_buffer_14183 (
        .din(new_Jinkela_wire_16896),
        .dout(new_Jinkela_wire_16897)
    );

    bfr new_Jinkela_buffer_14146 (
        .din(new_Jinkela_wire_16849),
        .dout(new_Jinkela_wire_16850)
    );

    bfr new_Jinkela_buffer_14202 (
        .din(new_Jinkela_wire_16921),
        .dout(new_Jinkela_wire_16922)
    );

    bfr new_Jinkela_buffer_14147 (
        .din(new_Jinkela_wire_16850),
        .dout(new_Jinkela_wire_16851)
    );

    bfr new_Jinkela_buffer_14184 (
        .din(new_Jinkela_wire_16897),
        .dout(new_Jinkela_wire_16898)
    );

    bfr new_Jinkela_buffer_14148 (
        .din(new_Jinkela_wire_16851),
        .dout(new_Jinkela_wire_16852)
    );

    spl2 new_Jinkela_splitter_1217 (
        .a(_1595_),
        .b(new_Jinkela_wire_16955),
        .c(new_Jinkela_wire_16956)
    );

    bfr new_Jinkela_buffer_14149 (
        .din(new_Jinkela_wire_16852),
        .dout(new_Jinkela_wire_16853)
    );

    bfr new_Jinkela_buffer_14185 (
        .din(new_Jinkela_wire_16898),
        .dout(new_Jinkela_wire_16899)
    );

    bfr new_Jinkela_buffer_14150 (
        .din(new_Jinkela_wire_16853),
        .dout(new_Jinkela_wire_16854)
    );

    bfr new_Jinkela_buffer_14203 (
        .din(new_Jinkela_wire_16922),
        .dout(new_Jinkela_wire_16923)
    );

    bfr new_Jinkela_buffer_14151 (
        .din(new_Jinkela_wire_16854),
        .dout(new_Jinkela_wire_16855)
    );

    bfr new_Jinkela_buffer_14186 (
        .din(new_Jinkela_wire_16899),
        .dout(new_Jinkela_wire_16900)
    );

    bfr new_Jinkela_buffer_14152 (
        .din(new_Jinkela_wire_16855),
        .dout(new_Jinkela_wire_16856)
    );

    spl2 new_Jinkela_splitter_1219 (
        .a(_1428_),
        .b(new_Jinkela_wire_16959),
        .c(new_Jinkela_wire_16960)
    );

    spl2 new_Jinkela_splitter_1218 (
        .a(_0534_),
        .b(new_Jinkela_wire_16957),
        .c(new_Jinkela_wire_16958)
    );

    bfr new_Jinkela_buffer_14153 (
        .din(new_Jinkela_wire_16856),
        .dout(new_Jinkela_wire_16857)
    );

    bfr new_Jinkela_buffer_14187 (
        .din(new_Jinkela_wire_16900),
        .dout(new_Jinkela_wire_16901)
    );

    bfr new_Jinkela_buffer_14154 (
        .din(new_Jinkela_wire_16857),
        .dout(new_Jinkela_wire_16858)
    );

    bfr new_Jinkela_buffer_14204 (
        .din(new_Jinkela_wire_16923),
        .dout(new_Jinkela_wire_16924)
    );

    bfr new_Jinkela_buffer_14155 (
        .din(new_Jinkela_wire_16858),
        .dout(new_Jinkela_wire_16859)
    );

    bfr new_Jinkela_buffer_14188 (
        .din(new_Jinkela_wire_16901),
        .dout(new_Jinkela_wire_16902)
    );

    bfr new_Jinkela_buffer_14156 (
        .din(new_Jinkela_wire_16859),
        .dout(new_Jinkela_wire_16860)
    );

    bfr new_Jinkela_buffer_17522 (
        .din(new_Jinkela_wire_20876),
        .dout(new_Jinkela_wire_20877)
    );

    bfr new_Jinkela_buffer_17613 (
        .din(new_Jinkela_wire_20979),
        .dout(new_Jinkela_wire_20980)
    );

    bfr new_Jinkela_buffer_17523 (
        .din(new_Jinkela_wire_20877),
        .dout(new_Jinkela_wire_20878)
    );

    bfr new_Jinkela_buffer_17578 (
        .din(new_Jinkela_wire_20938),
        .dout(new_Jinkela_wire_20939)
    );

    bfr new_Jinkela_buffer_17524 (
        .din(new_Jinkela_wire_20878),
        .dout(new_Jinkela_wire_20879)
    );

    bfr new_Jinkela_buffer_17631 (
        .din(new_Jinkela_wire_20999),
        .dout(new_Jinkela_wire_21000)
    );

    bfr new_Jinkela_buffer_17525 (
        .din(new_Jinkela_wire_20879),
        .dout(new_Jinkela_wire_20880)
    );

    bfr new_Jinkela_buffer_17579 (
        .din(new_Jinkela_wire_20939),
        .dout(new_Jinkela_wire_20940)
    );

    bfr new_Jinkela_buffer_17526 (
        .din(new_Jinkela_wire_20880),
        .dout(new_Jinkela_wire_20881)
    );

    bfr new_Jinkela_buffer_17614 (
        .din(new_Jinkela_wire_20980),
        .dout(new_Jinkela_wire_20981)
    );

    bfr new_Jinkela_buffer_17527 (
        .din(new_Jinkela_wire_20881),
        .dout(new_Jinkela_wire_20882)
    );

    bfr new_Jinkela_buffer_17580 (
        .din(new_Jinkela_wire_20940),
        .dout(new_Jinkela_wire_20941)
    );

    bfr new_Jinkela_buffer_17528 (
        .din(new_Jinkela_wire_20882),
        .dout(new_Jinkela_wire_20883)
    );

    spl2 new_Jinkela_splitter_1538 (
        .a(_0130_),
        .b(new_Jinkela_wire_21106),
        .c(new_Jinkela_wire_21107)
    );

    bfr new_Jinkela_buffer_17529 (
        .din(new_Jinkela_wire_20883),
        .dout(new_Jinkela_wire_20884)
    );

    bfr new_Jinkela_buffer_17581 (
        .din(new_Jinkela_wire_20941),
        .dout(new_Jinkela_wire_20942)
    );

    bfr new_Jinkela_buffer_17530 (
        .din(new_Jinkela_wire_20884),
        .dout(new_Jinkela_wire_20885)
    );

    bfr new_Jinkela_buffer_17615 (
        .din(new_Jinkela_wire_20981),
        .dout(new_Jinkela_wire_20982)
    );

    bfr new_Jinkela_buffer_17531 (
        .din(new_Jinkela_wire_20885),
        .dout(new_Jinkela_wire_20886)
    );

    bfr new_Jinkela_buffer_17582 (
        .din(new_Jinkela_wire_20942),
        .dout(new_Jinkela_wire_20943)
    );

    bfr new_Jinkela_buffer_17532 (
        .din(new_Jinkela_wire_20886),
        .dout(new_Jinkela_wire_20887)
    );

    bfr new_Jinkela_buffer_17632 (
        .din(new_Jinkela_wire_21000),
        .dout(new_Jinkela_wire_21001)
    );

    bfr new_Jinkela_buffer_17533 (
        .din(new_Jinkela_wire_20887),
        .dout(new_Jinkela_wire_20888)
    );

    bfr new_Jinkela_buffer_17583 (
        .din(new_Jinkela_wire_20943),
        .dout(new_Jinkela_wire_20944)
    );

    bfr new_Jinkela_buffer_17534 (
        .din(new_Jinkela_wire_20888),
        .dout(new_Jinkela_wire_20889)
    );

    bfr new_Jinkela_buffer_17616 (
        .din(new_Jinkela_wire_20982),
        .dout(new_Jinkela_wire_20983)
    );

    bfr new_Jinkela_buffer_17535 (
        .din(new_Jinkela_wire_20889),
        .dout(new_Jinkela_wire_20890)
    );

    bfr new_Jinkela_buffer_17584 (
        .din(new_Jinkela_wire_20944),
        .dout(new_Jinkela_wire_20945)
    );

    bfr new_Jinkela_buffer_17536 (
        .din(new_Jinkela_wire_20890),
        .dout(new_Jinkela_wire_20891)
    );

    spl2 new_Jinkela_splitter_1539 (
        .a(_0582_),
        .b(new_Jinkela_wire_21108),
        .c(new_Jinkela_wire_21109)
    );

    bfr new_Jinkela_buffer_17537 (
        .din(new_Jinkela_wire_20891),
        .dout(new_Jinkela_wire_20892)
    );

    bfr new_Jinkela_buffer_17585 (
        .din(new_Jinkela_wire_20945),
        .dout(new_Jinkela_wire_20946)
    );

    bfr new_Jinkela_buffer_17538 (
        .din(new_Jinkela_wire_20892),
        .dout(new_Jinkela_wire_20893)
    );

    bfr new_Jinkela_buffer_17617 (
        .din(new_Jinkela_wire_20983),
        .dout(new_Jinkela_wire_20984)
    );

    bfr new_Jinkela_buffer_17539 (
        .din(new_Jinkela_wire_20893),
        .dout(new_Jinkela_wire_20894)
    );

    bfr new_Jinkela_buffer_17586 (
        .din(new_Jinkela_wire_20946),
        .dout(new_Jinkela_wire_20947)
    );

    bfr new_Jinkela_buffer_17540 (
        .din(new_Jinkela_wire_20894),
        .dout(new_Jinkela_wire_20895)
    );

    bfr new_Jinkela_buffer_17633 (
        .din(new_Jinkela_wire_21001),
        .dout(new_Jinkela_wire_21002)
    );

    bfr new_Jinkela_buffer_17541 (
        .din(new_Jinkela_wire_20895),
        .dout(new_Jinkela_wire_20896)
    );

    bfr new_Jinkela_buffer_17587 (
        .din(new_Jinkela_wire_20947),
        .dout(new_Jinkela_wire_20948)
    );

    bfr new_Jinkela_buffer_17542 (
        .din(new_Jinkela_wire_20896),
        .dout(new_Jinkela_wire_20897)
    );

    bfr new_Jinkela_buffer_17618 (
        .din(new_Jinkela_wire_20984),
        .dout(new_Jinkela_wire_20985)
    );

    bfr new_Jinkela_buffer_7169 (
        .din(new_Jinkela_wire_8948),
        .dout(new_Jinkela_wire_8949)
    );

    bfr new_Jinkela_buffer_7221 (
        .din(new_Jinkela_wire_9004),
        .dout(new_Jinkela_wire_9005)
    );

    bfr new_Jinkela_buffer_7170 (
        .din(new_Jinkela_wire_8949),
        .dout(new_Jinkela_wire_8950)
    );

    bfr new_Jinkela_buffer_7243 (
        .din(new_Jinkela_wire_9034),
        .dout(new_Jinkela_wire_9035)
    );

    bfr new_Jinkela_buffer_7171 (
        .din(new_Jinkela_wire_8950),
        .dout(new_Jinkela_wire_8951)
    );

    bfr new_Jinkela_buffer_7222 (
        .din(new_Jinkela_wire_9005),
        .dout(new_Jinkela_wire_9006)
    );

    bfr new_Jinkela_buffer_7172 (
        .din(new_Jinkela_wire_8951),
        .dout(new_Jinkela_wire_8952)
    );

    bfr new_Jinkela_buffer_7308 (
        .din(new_Jinkela_wire_9109),
        .dout(new_Jinkela_wire_9110)
    );

    bfr new_Jinkela_buffer_7173 (
        .din(new_Jinkela_wire_8952),
        .dout(new_Jinkela_wire_8953)
    );

    bfr new_Jinkela_buffer_7223 (
        .din(new_Jinkela_wire_9006),
        .dout(new_Jinkela_wire_9007)
    );

    bfr new_Jinkela_buffer_7174 (
        .din(new_Jinkela_wire_8953),
        .dout(new_Jinkela_wire_8954)
    );

    bfr new_Jinkela_buffer_7244 (
        .din(new_Jinkela_wire_9035),
        .dout(new_Jinkela_wire_9036)
    );

    bfr new_Jinkela_buffer_7175 (
        .din(new_Jinkela_wire_8954),
        .dout(new_Jinkela_wire_8955)
    );

    bfr new_Jinkela_buffer_7224 (
        .din(new_Jinkela_wire_9007),
        .dout(new_Jinkela_wire_9008)
    );

    bfr new_Jinkela_buffer_7176 (
        .din(new_Jinkela_wire_8955),
        .dout(new_Jinkela_wire_8956)
    );

    spl2 new_Jinkela_splitter_756 (
        .a(_1551_),
        .b(new_Jinkela_wire_9185),
        .c(new_Jinkela_wire_9186)
    );

    bfr new_Jinkela_buffer_7177 (
        .din(new_Jinkela_wire_8956),
        .dout(new_Jinkela_wire_8957)
    );

    bfr new_Jinkela_buffer_7225 (
        .din(new_Jinkela_wire_9008),
        .dout(new_Jinkela_wire_9009)
    );

    bfr new_Jinkela_buffer_7178 (
        .din(new_Jinkela_wire_8957),
        .dout(new_Jinkela_wire_8958)
    );

    bfr new_Jinkela_buffer_7245 (
        .din(new_Jinkela_wire_9036),
        .dout(new_Jinkela_wire_9037)
    );

    bfr new_Jinkela_buffer_7179 (
        .din(new_Jinkela_wire_8958),
        .dout(new_Jinkela_wire_8959)
    );

    spl2 new_Jinkela_splitter_741 (
        .a(new_Jinkela_wire_9009),
        .b(new_Jinkela_wire_9010),
        .c(new_Jinkela_wire_9011)
    );

    bfr new_Jinkela_buffer_7180 (
        .din(new_Jinkela_wire_8959),
        .dout(new_Jinkela_wire_8960)
    );

    bfr new_Jinkela_buffer_7246 (
        .din(new_Jinkela_wire_9037),
        .dout(new_Jinkela_wire_9038)
    );

    spl2 new_Jinkela_splitter_739 (
        .a(new_Jinkela_wire_8960),
        .b(new_Jinkela_wire_8961),
        .c(new_Jinkela_wire_8962)
    );

    spl2 new_Jinkela_splitter_755 (
        .a(_1410_),
        .b(new_Jinkela_wire_9183),
        .c(new_Jinkela_wire_9184)
    );

    bfr new_Jinkela_buffer_7309 (
        .din(new_Jinkela_wire_9110),
        .dout(new_Jinkela_wire_9111)
    );

    bfr new_Jinkela_buffer_7247 (
        .din(new_Jinkela_wire_9038),
        .dout(new_Jinkela_wire_9039)
    );

    bfr new_Jinkela_buffer_7310 (
        .din(new_Jinkela_wire_9111),
        .dout(new_Jinkela_wire_9112)
    );

    bfr new_Jinkela_buffer_7248 (
        .din(new_Jinkela_wire_9039),
        .dout(new_Jinkela_wire_9040)
    );

    bfr new_Jinkela_buffer_7370 (
        .din(new_Jinkela_wire_9179),
        .dout(new_Jinkela_wire_9180)
    );

    bfr new_Jinkela_buffer_7371 (
        .din(_0961_),
        .dout(new_Jinkela_wire_9187)
    );

    bfr new_Jinkela_buffer_7249 (
        .din(new_Jinkela_wire_9040),
        .dout(new_Jinkela_wire_9041)
    );

    bfr new_Jinkela_buffer_7311 (
        .din(new_Jinkela_wire_9112),
        .dout(new_Jinkela_wire_9113)
    );

    bfr new_Jinkela_buffer_7250 (
        .din(new_Jinkela_wire_9041),
        .dout(new_Jinkela_wire_9042)
    );

    bfr new_Jinkela_buffer_7251 (
        .din(new_Jinkela_wire_9042),
        .dout(new_Jinkela_wire_9043)
    );

    bfr new_Jinkela_buffer_7312 (
        .din(new_Jinkela_wire_9113),
        .dout(new_Jinkela_wire_9114)
    );

    bfr new_Jinkela_buffer_7252 (
        .din(new_Jinkela_wire_9043),
        .dout(new_Jinkela_wire_9044)
    );

    spl2 new_Jinkela_splitter_754 (
        .a(new_Jinkela_wire_9180),
        .b(new_Jinkela_wire_9181),
        .c(new_Jinkela_wire_9182)
    );

    bfr new_Jinkela_buffer_7253 (
        .din(new_Jinkela_wire_9044),
        .dout(new_Jinkela_wire_9045)
    );

    bfr new_Jinkela_buffer_7313 (
        .din(new_Jinkela_wire_9114),
        .dout(new_Jinkela_wire_9115)
    );

    bfr new_Jinkela_buffer_7254 (
        .din(new_Jinkela_wire_9045),
        .dout(new_Jinkela_wire_9046)
    );

    bfr new_Jinkela_buffer_10811 (
        .din(new_Jinkela_wire_13022),
        .dout(new_Jinkela_wire_13023)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_10680 (
        .din(new_Jinkela_wire_12881),
        .dout(new_Jinkela_wire_12882)
    );

    spl2 new_Jinkela_splitter_202 (
        .a(_0507_),
        .b(new_Jinkela_wire_1136),
        .c(new_Jinkela_wire_1137)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_10726 (
        .din(new_Jinkela_wire_12931),
        .dout(new_Jinkela_wire_12932)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_10681 (
        .din(new_Jinkela_wire_12882),
        .dout(new_Jinkela_wire_12883)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_10836 (
        .din(new_Jinkela_wire_13051),
        .dout(new_Jinkela_wire_13052)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    bfr new_Jinkela_buffer_10682 (
        .din(new_Jinkela_wire_12883),
        .dout(new_Jinkela_wire_12884)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_10727 (
        .din(new_Jinkela_wire_12932),
        .dout(new_Jinkela_wire_12933)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_10683 (
        .din(new_Jinkela_wire_12884),
        .dout(new_Jinkela_wire_12885)
    );

    bfr new_Jinkela_buffer_10812 (
        .din(new_Jinkela_wire_13023),
        .dout(new_Jinkela_wire_13024)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_821),
        .dout(new_Jinkela_wire_822)
    );

    bfr new_Jinkela_buffer_10684 (
        .din(new_Jinkela_wire_12885),
        .dout(new_Jinkela_wire_12886)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_10728 (
        .din(new_Jinkela_wire_12933),
        .dout(new_Jinkela_wire_12934)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_822),
        .dout(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_10685 (
        .din(new_Jinkela_wire_12886),
        .dout(new_Jinkela_wire_12887)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    bfr new_Jinkela_buffer_10686 (
        .din(new_Jinkela_wire_12887),
        .dout(new_Jinkela_wire_12888)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_1022),
        .dout(new_Jinkela_wire_1023)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_10729 (
        .din(new_Jinkela_wire_12934),
        .dout(new_Jinkela_wire_12935)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    bfr new_Jinkela_buffer_10687 (
        .din(new_Jinkela_wire_12888),
        .dout(new_Jinkela_wire_12889)
    );

    bfr new_Jinkela_buffer_10813 (
        .din(new_Jinkela_wire_13024),
        .dout(new_Jinkela_wire_13025)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_825),
        .dout(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_10688 (
        .din(new_Jinkela_wire_12889),
        .dout(new_Jinkela_wire_12890)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_10730 (
        .din(new_Jinkela_wire_12935),
        .dout(new_Jinkela_wire_12936)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    bfr new_Jinkela_buffer_10689 (
        .din(new_Jinkela_wire_12890),
        .dout(new_Jinkela_wire_12891)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    spl2 new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_827),
        .b(new_Jinkela_wire_828),
        .c(new_Jinkela_wire_829)
    );

    spl2 new_Jinkela_splitter_961 (
        .a(_0958_),
        .b(new_Jinkela_wire_13062),
        .c(new_Jinkela_wire_13063)
    );

    bfr new_Jinkela_buffer_10690 (
        .din(new_Jinkela_wire_12891),
        .dout(new_Jinkela_wire_12892)
    );

    bfr new_Jinkela_buffer_10731 (
        .din(new_Jinkela_wire_12936),
        .dout(new_Jinkela_wire_12937)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_1023),
        .dout(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_10691 (
        .din(new_Jinkela_wire_12892),
        .dout(new_Jinkela_wire_12893)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_10814 (
        .din(new_Jinkela_wire_13025),
        .dout(new_Jinkela_wire_13026)
    );

    bfr new_Jinkela_buffer_10692 (
        .din(new_Jinkela_wire_12893),
        .dout(new_Jinkela_wire_12894)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_10732 (
        .din(new_Jinkela_wire_12937),
        .dout(new_Jinkela_wire_12938)
    );

    bfr new_Jinkela_buffer_10693 (
        .din(new_Jinkela_wire_12894),
        .dout(new_Jinkela_wire_12895)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_10838 (
        .din(_0727_),
        .dout(new_Jinkela_wire_13064)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_1080),
        .dout(new_Jinkela_wire_1081)
    );

    bfr new_Jinkela_buffer_10694 (
        .din(new_Jinkela_wire_12895),
        .dout(new_Jinkela_wire_12896)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_10733 (
        .din(new_Jinkela_wire_12938),
        .dout(new_Jinkela_wire_12939)
    );

    bfr new_Jinkela_buffer_10695 (
        .din(new_Jinkela_wire_12896),
        .dout(new_Jinkela_wire_12897)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_10815 (
        .din(new_Jinkela_wire_13026),
        .dout(new_Jinkela_wire_13027)
    );

    spl2 new_Jinkela_splitter_203 (
        .a(_1636_),
        .b(new_Jinkela_wire_1138),
        .c(new_Jinkela_wire_1139)
    );

    bfr new_Jinkela_buffer_10696 (
        .din(new_Jinkela_wire_12897),
        .dout(new_Jinkela_wire_12898)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_10734 (
        .din(new_Jinkela_wire_12939),
        .dout(new_Jinkela_wire_12940)
    );

    bfr new_Jinkela_buffer_10697 (
        .din(new_Jinkela_wire_12898),
        .dout(new_Jinkela_wire_12899)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(_0136_),
        .b(new_Jinkela_wire_1254),
        .c(new_Jinkela_wire_1255)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_10839 (
        .din(_1813_),
        .dout(new_Jinkela_wire_13067)
    );

    spl2 new_Jinkela_splitter_962 (
        .a(_1335_),
        .b(new_Jinkela_wire_13065),
        .c(new_Jinkela_wire_13066)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_10698 (
        .din(new_Jinkela_wire_12899),
        .dout(new_Jinkela_wire_12900)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_10735 (
        .din(new_Jinkela_wire_12940),
        .dout(new_Jinkela_wire_12941)
    );

    bfr new_Jinkela_buffer_10699 (
        .din(new_Jinkela_wire_12900),
        .dout(new_Jinkela_wire_12901)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_10816 (
        .din(new_Jinkela_wire_13027),
        .dout(new_Jinkela_wire_13028)
    );

    bfr new_Jinkela_buffer_430 (
        .din(_1678_),
        .dout(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_10700 (
        .din(new_Jinkela_wire_12901),
        .dout(new_Jinkela_wire_12902)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_3828 (
        .din(new_Jinkela_wire_5063),
        .dout(new_Jinkela_wire_5064)
    );

    bfr new_Jinkela_buffer_14157 (
        .din(new_Jinkela_wire_16860),
        .dout(new_Jinkela_wire_16861)
    );

    spl2 new_Jinkela_splitter_455 (
        .a(new_Jinkela_wire_4979),
        .b(new_Jinkela_wire_4980),
        .c(new_Jinkela_wire_4981)
    );

    bfr new_Jinkela_buffer_14189 (
        .din(new_Jinkela_wire_16902),
        .dout(new_Jinkela_wire_16903)
    );

    bfr new_Jinkela_buffer_3861 (
        .din(new_Jinkela_wire_5100),
        .dout(new_Jinkela_wire_5101)
    );

    bfr new_Jinkela_buffer_14158 (
        .din(new_Jinkela_wire_16861),
        .dout(new_Jinkela_wire_16862)
    );

    bfr new_Jinkela_buffer_3803 (
        .din(new_Jinkela_wire_5026),
        .dout(new_Jinkela_wire_5027)
    );

    bfr new_Jinkela_buffer_14205 (
        .din(new_Jinkela_wire_16924),
        .dout(new_Jinkela_wire_16925)
    );

    bfr new_Jinkela_buffer_3804 (
        .din(new_Jinkela_wire_5027),
        .dout(new_Jinkela_wire_5028)
    );

    bfr new_Jinkela_buffer_14159 (
        .din(new_Jinkela_wire_16862),
        .dout(new_Jinkela_wire_16863)
    );

    bfr new_Jinkela_buffer_3829 (
        .din(new_Jinkela_wire_5064),
        .dout(new_Jinkela_wire_5065)
    );

    bfr new_Jinkela_buffer_3805 (
        .din(new_Jinkela_wire_5028),
        .dout(new_Jinkela_wire_5029)
    );

    spl2 new_Jinkela_splitter_1220 (
        .a(_0482_),
        .b(new_Jinkela_wire_16961),
        .c(new_Jinkela_wire_16962)
    );

    spl2 new_Jinkela_splitter_1201 (
        .a(new_Jinkela_wire_16863),
        .b(new_Jinkela_wire_16864),
        .c(new_Jinkela_wire_16865)
    );

    spl2 new_Jinkela_splitter_474 (
        .a(_1449_),
        .b(new_Jinkela_wire_5133),
        .c(new_Jinkela_wire_5134)
    );

    spl2 new_Jinkela_splitter_472 (
        .a(_0179_),
        .b(new_Jinkela_wire_5127),
        .c(new_Jinkela_wire_5128)
    );

    bfr new_Jinkela_buffer_3806 (
        .din(new_Jinkela_wire_5029),
        .dout(new_Jinkela_wire_5030)
    );

    spl2 new_Jinkela_splitter_1221 (
        .a(_0185_),
        .b(new_Jinkela_wire_16967),
        .c(new_Jinkela_wire_16968)
    );

    bfr new_Jinkela_buffer_14206 (
        .din(new_Jinkela_wire_16925),
        .dout(new_Jinkela_wire_16926)
    );

    bfr new_Jinkela_buffer_3830 (
        .din(new_Jinkela_wire_5065),
        .dout(new_Jinkela_wire_5066)
    );

    bfr new_Jinkela_buffer_14207 (
        .din(new_Jinkela_wire_16926),
        .dout(new_Jinkela_wire_16927)
    );

    bfr new_Jinkela_buffer_3807 (
        .din(new_Jinkela_wire_5030),
        .dout(new_Jinkela_wire_5031)
    );

    bfr new_Jinkela_buffer_14219 (
        .din(new_Jinkela_wire_16962),
        .dout(new_Jinkela_wire_16963)
    );

    bfr new_Jinkela_buffer_3862 (
        .din(new_Jinkela_wire_5101),
        .dout(new_Jinkela_wire_5102)
    );

    bfr new_Jinkela_buffer_14223 (
        .din(_1677_),
        .dout(new_Jinkela_wire_16969)
    );

    bfr new_Jinkela_buffer_14208 (
        .din(new_Jinkela_wire_16927),
        .dout(new_Jinkela_wire_16928)
    );

    bfr new_Jinkela_buffer_3808 (
        .din(new_Jinkela_wire_5031),
        .dout(new_Jinkela_wire_5032)
    );

    spl2 new_Jinkela_splitter_1222 (
        .a(_1137_),
        .b(new_Jinkela_wire_16971),
        .c(new_Jinkela_wire_16972)
    );

    bfr new_Jinkela_buffer_3831 (
        .din(new_Jinkela_wire_5066),
        .dout(new_Jinkela_wire_5067)
    );

    bfr new_Jinkela_buffer_14209 (
        .din(new_Jinkela_wire_16928),
        .dout(new_Jinkela_wire_16929)
    );

    bfr new_Jinkela_buffer_3809 (
        .din(new_Jinkela_wire_5032),
        .dout(new_Jinkela_wire_5033)
    );

    bfr new_Jinkela_buffer_14220 (
        .din(new_Jinkela_wire_16963),
        .dout(new_Jinkela_wire_16964)
    );

    bfr new_Jinkela_buffer_3880 (
        .din(_1194_),
        .dout(new_Jinkela_wire_5126)
    );

    bfr new_Jinkela_buffer_14210 (
        .din(new_Jinkela_wire_16929),
        .dout(new_Jinkela_wire_16930)
    );

    bfr new_Jinkela_buffer_3810 (
        .din(new_Jinkela_wire_5033),
        .dout(new_Jinkela_wire_5034)
    );

    bfr new_Jinkela_buffer_3832 (
        .din(new_Jinkela_wire_5067),
        .dout(new_Jinkela_wire_5068)
    );

    bfr new_Jinkela_buffer_14224 (
        .din(_0663_),
        .dout(new_Jinkela_wire_16970)
    );

    bfr new_Jinkela_buffer_14211 (
        .din(new_Jinkela_wire_16930),
        .dout(new_Jinkela_wire_16931)
    );

    bfr new_Jinkela_buffer_3811 (
        .din(new_Jinkela_wire_5034),
        .dout(new_Jinkela_wire_5035)
    );

    bfr new_Jinkela_buffer_14221 (
        .din(new_Jinkela_wire_16964),
        .dout(new_Jinkela_wire_16965)
    );

    bfr new_Jinkela_buffer_3863 (
        .din(new_Jinkela_wire_5102),
        .dout(new_Jinkela_wire_5103)
    );

    bfr new_Jinkela_buffer_14212 (
        .din(new_Jinkela_wire_16931),
        .dout(new_Jinkela_wire_16932)
    );

    bfr new_Jinkela_buffer_3812 (
        .din(new_Jinkela_wire_5035),
        .dout(new_Jinkela_wire_5036)
    );

    bfr new_Jinkela_buffer_14225 (
        .din(_1582_),
        .dout(new_Jinkela_wire_16973)
    );

    bfr new_Jinkela_buffer_3833 (
        .din(new_Jinkela_wire_5068),
        .dout(new_Jinkela_wire_5069)
    );

    bfr new_Jinkela_buffer_14213 (
        .din(new_Jinkela_wire_16932),
        .dout(new_Jinkela_wire_16933)
    );

    bfr new_Jinkela_buffer_3813 (
        .din(new_Jinkela_wire_5036),
        .dout(new_Jinkela_wire_5037)
    );

    bfr new_Jinkela_buffer_14222 (
        .din(new_Jinkela_wire_16965),
        .dout(new_Jinkela_wire_16966)
    );

    bfr new_Jinkela_buffer_3865 (
        .din(new_Jinkela_wire_5108),
        .dout(new_Jinkela_wire_5109)
    );

    bfr new_Jinkela_buffer_14214 (
        .din(new_Jinkela_wire_16933),
        .dout(new_Jinkela_wire_16934)
    );

    bfr new_Jinkela_buffer_3814 (
        .din(new_Jinkela_wire_5037),
        .dout(new_Jinkela_wire_5038)
    );

    spl2 new_Jinkela_splitter_1225 (
        .a(_0398_),
        .b(new_Jinkela_wire_17005),
        .c(new_Jinkela_wire_17006)
    );

    bfr new_Jinkela_buffer_3834 (
        .din(new_Jinkela_wire_5069),
        .dout(new_Jinkela_wire_5070)
    );

    bfr new_Jinkela_buffer_14215 (
        .din(new_Jinkela_wire_16934),
        .dout(new_Jinkela_wire_16935)
    );

    bfr new_Jinkela_buffer_3815 (
        .din(new_Jinkela_wire_5038),
        .dout(new_Jinkela_wire_5039)
    );

    spl2 new_Jinkela_splitter_473 (
        .a(_0275_),
        .b(new_Jinkela_wire_5129),
        .c(new_Jinkela_wire_5130)
    );

    bfr new_Jinkela_buffer_3882 (
        .din(new_Jinkela_wire_5131),
        .dout(new_Jinkela_wire_5132)
    );

    spl2 new_Jinkela_splitter_1224 (
        .a(_1522_),
        .b(new_Jinkela_wire_16999),
        .c(new_Jinkela_wire_17000)
    );

    bfr new_Jinkela_buffer_14216 (
        .din(new_Jinkela_wire_16935),
        .dout(new_Jinkela_wire_16936)
    );

    bfr new_Jinkela_buffer_3816 (
        .din(new_Jinkela_wire_5039),
        .dout(new_Jinkela_wire_5040)
    );

    bfr new_Jinkela_buffer_14226 (
        .din(new_Jinkela_wire_16973),
        .dout(new_Jinkela_wire_16974)
    );

    bfr new_Jinkela_buffer_3835 (
        .din(new_Jinkela_wire_5070),
        .dout(new_Jinkela_wire_5071)
    );

    bfr new_Jinkela_buffer_14217 (
        .din(new_Jinkela_wire_16936),
        .dout(new_Jinkela_wire_16937)
    );

    spl2 new_Jinkela_splitter_461 (
        .a(new_Jinkela_wire_5040),
        .b(new_Jinkela_wire_5041),
        .c(new_Jinkela_wire_5042)
    );

    bfr new_Jinkela_buffer_3836 (
        .din(new_Jinkela_wire_5071),
        .dout(new_Jinkela_wire_5072)
    );

    bfr new_Jinkela_buffer_14218 (
        .din(new_Jinkela_wire_16937),
        .dout(new_Jinkela_wire_16938)
    );

    bfr new_Jinkela_buffer_3866 (
        .din(new_Jinkela_wire_5109),
        .dout(new_Jinkela_wire_5110)
    );

    bfr new_Jinkela_buffer_14227 (
        .din(new_Jinkela_wire_16974),
        .dout(new_Jinkela_wire_16975)
    );

    spl2 new_Jinkela_splitter_1209 (
        .a(new_Jinkela_wire_16938),
        .b(new_Jinkela_wire_16939),
        .c(new_Jinkela_wire_16940)
    );

    bfr new_Jinkela_buffer_3837 (
        .din(new_Jinkela_wire_5072),
        .dout(new_Jinkela_wire_5073)
    );

    bfr new_Jinkela_buffer_14228 (
        .din(new_Jinkela_wire_16975),
        .dout(new_Jinkela_wire_16976)
    );

    bfr new_Jinkela_buffer_3867 (
        .din(new_Jinkela_wire_5110),
        .dout(new_Jinkela_wire_5111)
    );

    bfr new_Jinkela_buffer_14249 (
        .din(new_Jinkela_wire_17000),
        .dout(new_Jinkela_wire_17001)
    );

    bfr new_Jinkela_buffer_3838 (
        .din(new_Jinkela_wire_5073),
        .dout(new_Jinkela_wire_5074)
    );

    spl2 new_Jinkela_splitter_1226 (
        .a(_1565_),
        .b(new_Jinkela_wire_17011),
        .c(new_Jinkela_wire_17012)
    );

    bfr new_Jinkela_buffer_3881 (
        .din(_1195_),
        .dout(new_Jinkela_wire_5131)
    );

    bfr new_Jinkela_buffer_14229 (
        .din(new_Jinkela_wire_16976),
        .dout(new_Jinkela_wire_16977)
    );

    bfr new_Jinkela_buffer_3839 (
        .din(new_Jinkela_wire_5074),
        .dout(new_Jinkela_wire_5075)
    );

    bfr new_Jinkela_buffer_14250 (
        .din(new_Jinkela_wire_17001),
        .dout(new_Jinkela_wire_17002)
    );

    bfr new_Jinkela_buffer_3868 (
        .din(new_Jinkela_wire_5111),
        .dout(new_Jinkela_wire_5112)
    );

    bfr new_Jinkela_buffer_14230 (
        .din(new_Jinkela_wire_16977),
        .dout(new_Jinkela_wire_16978)
    );

    bfr new_Jinkela_buffer_3840 (
        .din(new_Jinkela_wire_5075),
        .dout(new_Jinkela_wire_5076)
    );

    bfr new_Jinkela_buffer_14253 (
        .din(new_Jinkela_wire_17006),
        .dout(new_Jinkela_wire_17007)
    );

    bfr new_Jinkela_buffer_3883 (
        .din(_0660_),
        .dout(new_Jinkela_wire_5135)
    );

    spl2 new_Jinkela_splitter_1227 (
        .a(_0040_),
        .b(new_Jinkela_wire_17013),
        .c(new_Jinkela_wire_17014)
    );

    bfr new_Jinkela_buffer_17543 (
        .din(new_Jinkela_wire_20897),
        .dout(new_Jinkela_wire_20898)
    );

    bfr new_Jinkela_buffer_17588 (
        .din(new_Jinkela_wire_20948),
        .dout(new_Jinkela_wire_20949)
    );

    spl2 new_Jinkela_splitter_1526 (
        .a(new_Jinkela_wire_20898),
        .b(new_Jinkela_wire_20899),
        .c(new_Jinkela_wire_20900)
    );

    bfr new_Jinkela_buffer_17589 (
        .din(new_Jinkela_wire_20949),
        .dout(new_Jinkela_wire_20950)
    );

    bfr new_Jinkela_buffer_17723 (
        .din(new_Jinkela_wire_21101),
        .dout(new_Jinkela_wire_21102)
    );

    bfr new_Jinkela_buffer_17619 (
        .din(new_Jinkela_wire_20985),
        .dout(new_Jinkela_wire_20986)
    );

    bfr new_Jinkela_buffer_17590 (
        .din(new_Jinkela_wire_20950),
        .dout(new_Jinkela_wire_20951)
    );

    bfr new_Jinkela_buffer_17634 (
        .din(new_Jinkela_wire_21002),
        .dout(new_Jinkela_wire_21003)
    );

    bfr new_Jinkela_buffer_17591 (
        .din(new_Jinkela_wire_20951),
        .dout(new_Jinkela_wire_20952)
    );

    bfr new_Jinkela_buffer_17620 (
        .din(new_Jinkela_wire_20986),
        .dout(new_Jinkela_wire_20987)
    );

    bfr new_Jinkela_buffer_17592 (
        .din(new_Jinkela_wire_20952),
        .dout(new_Jinkela_wire_20953)
    );

    bfr new_Jinkela_buffer_17593 (
        .din(new_Jinkela_wire_20953),
        .dout(new_Jinkela_wire_20954)
    );

    bfr new_Jinkela_buffer_17621 (
        .din(new_Jinkela_wire_20987),
        .dout(new_Jinkela_wire_20988)
    );

    bfr new_Jinkela_buffer_17594 (
        .din(new_Jinkela_wire_20954),
        .dout(new_Jinkela_wire_20955)
    );

    bfr new_Jinkela_buffer_17635 (
        .din(new_Jinkela_wire_21003),
        .dout(new_Jinkela_wire_21004)
    );

    bfr new_Jinkela_buffer_17595 (
        .din(new_Jinkela_wire_20955),
        .dout(new_Jinkela_wire_20956)
    );

    bfr new_Jinkela_buffer_17622 (
        .din(new_Jinkela_wire_20988),
        .dout(new_Jinkela_wire_20989)
    );

    bfr new_Jinkela_buffer_17596 (
        .din(new_Jinkela_wire_20956),
        .dout(new_Jinkela_wire_20957)
    );

    bfr new_Jinkela_buffer_17724 (
        .din(new_Jinkela_wire_21102),
        .dout(new_Jinkela_wire_21103)
    );

    spl2 new_Jinkela_splitter_1529 (
        .a(new_Jinkela_wire_20957),
        .b(new_Jinkela_wire_20958),
        .c(new_Jinkela_wire_20959)
    );

    bfr new_Jinkela_buffer_17636 (
        .din(new_Jinkela_wire_21004),
        .dout(new_Jinkela_wire_21005)
    );

    bfr new_Jinkela_buffer_17623 (
        .din(new_Jinkela_wire_20989),
        .dout(new_Jinkela_wire_20990)
    );

    bfr new_Jinkela_buffer_17624 (
        .din(new_Jinkela_wire_20990),
        .dout(new_Jinkela_wire_20991)
    );

    spl2 new_Jinkela_splitter_1540 (
        .a(_1761_),
        .b(new_Jinkela_wire_21110),
        .c(new_Jinkela_wire_21111)
    );

    spl2 new_Jinkela_splitter_1532 (
        .a(new_Jinkela_wire_20991),
        .b(new_Jinkela_wire_20992),
        .c(new_Jinkela_wire_20993)
    );

    bfr new_Jinkela_buffer_17725 (
        .din(new_Jinkela_wire_21103),
        .dout(new_Jinkela_wire_21104)
    );

    bfr new_Jinkela_buffer_17637 (
        .din(new_Jinkela_wire_21005),
        .dout(new_Jinkela_wire_21006)
    );

    bfr new_Jinkela_buffer_17638 (
        .din(new_Jinkela_wire_21006),
        .dout(new_Jinkela_wire_21007)
    );

    spl2 new_Jinkela_splitter_1541 (
        .a(_0772_),
        .b(new_Jinkela_wire_21114),
        .c(new_Jinkela_wire_21115)
    );

    bfr new_Jinkela_buffer_17727 (
        .din(_1000_),
        .dout(new_Jinkela_wire_21112)
    );

    bfr new_Jinkela_buffer_17639 (
        .din(new_Jinkela_wire_21007),
        .dout(new_Jinkela_wire_21008)
    );

    bfr new_Jinkela_buffer_17728 (
        .din(_0168_),
        .dout(new_Jinkela_wire_21113)
    );

    bfr new_Jinkela_buffer_17640 (
        .din(new_Jinkela_wire_21008),
        .dout(new_Jinkela_wire_21009)
    );

    bfr new_Jinkela_buffer_17729 (
        .din(_0637_),
        .dout(new_Jinkela_wire_21116)
    );

    bfr new_Jinkela_buffer_17734 (
        .din(_1149_),
        .dout(new_Jinkela_wire_21123)
    );

    bfr new_Jinkela_buffer_17641 (
        .din(new_Jinkela_wire_21009),
        .dout(new_Jinkela_wire_21010)
    );

    bfr new_Jinkela_buffer_17730 (
        .din(new_Jinkela_wire_21118),
        .dout(new_Jinkela_wire_21119)
    );

    bfr new_Jinkela_buffer_17642 (
        .din(new_Jinkela_wire_21010),
        .dout(new_Jinkela_wire_21011)
    );

    spl2 new_Jinkela_splitter_1542 (
        .a(_0989_),
        .b(new_Jinkela_wire_21117),
        .c(new_Jinkela_wire_21118)
    );

    bfr new_Jinkela_buffer_17643 (
        .din(new_Jinkela_wire_21011),
        .dout(new_Jinkela_wire_21012)
    );

    bfr new_Jinkela_buffer_17644 (
        .din(new_Jinkela_wire_21012),
        .dout(new_Jinkela_wire_21013)
    );

    spl2 new_Jinkela_splitter_1543 (
        .a(_0609_),
        .b(new_Jinkela_wire_21124),
        .c(new_Jinkela_wire_21125)
    );

    bfr new_Jinkela_buffer_10736 (
        .din(new_Jinkela_wire_12941),
        .dout(new_Jinkela_wire_12942)
    );

    spl2 new_Jinkela_splitter_950 (
        .a(new_Jinkela_wire_12902),
        .b(new_Jinkela_wire_12903),
        .c(new_Jinkela_wire_12904)
    );

    bfr new_Jinkela_buffer_10737 (
        .din(new_Jinkela_wire_12942),
        .dout(new_Jinkela_wire_12943)
    );

    spl2 new_Jinkela_splitter_965 (
        .a(_0182_),
        .b(new_Jinkela_wire_13147),
        .c(new_Jinkela_wire_13148)
    );

    bfr new_Jinkela_buffer_10817 (
        .din(new_Jinkela_wire_13028),
        .dout(new_Jinkela_wire_13029)
    );

    bfr new_Jinkela_buffer_10738 (
        .din(new_Jinkela_wire_12943),
        .dout(new_Jinkela_wire_12944)
    );

    spl2 new_Jinkela_splitter_964 (
        .a(_1302_),
        .b(new_Jinkela_wire_13141),
        .c(new_Jinkela_wire_13142)
    );

    bfr new_Jinkela_buffer_10739 (
        .din(new_Jinkela_wire_12944),
        .dout(new_Jinkela_wire_12945)
    );

    bfr new_Jinkela_buffer_10818 (
        .din(new_Jinkela_wire_13029),
        .dout(new_Jinkela_wire_13030)
    );

    bfr new_Jinkela_buffer_10740 (
        .din(new_Jinkela_wire_12945),
        .dout(new_Jinkela_wire_12946)
    );

    bfr new_Jinkela_buffer_10840 (
        .din(new_Jinkela_wire_13067),
        .dout(new_Jinkela_wire_13068)
    );

    bfr new_Jinkela_buffer_10741 (
        .din(new_Jinkela_wire_12946),
        .dout(new_Jinkela_wire_12947)
    );

    bfr new_Jinkela_buffer_10819 (
        .din(new_Jinkela_wire_13030),
        .dout(new_Jinkela_wire_13031)
    );

    bfr new_Jinkela_buffer_10742 (
        .din(new_Jinkela_wire_12947),
        .dout(new_Jinkela_wire_12948)
    );

    bfr new_Jinkela_buffer_10743 (
        .din(new_Jinkela_wire_12948),
        .dout(new_Jinkela_wire_12949)
    );

    bfr new_Jinkela_buffer_10820 (
        .din(new_Jinkela_wire_13031),
        .dout(new_Jinkela_wire_13032)
    );

    bfr new_Jinkela_buffer_10744 (
        .din(new_Jinkela_wire_12949),
        .dout(new_Jinkela_wire_12950)
    );

    bfr new_Jinkela_buffer_10841 (
        .din(new_Jinkela_wire_13068),
        .dout(new_Jinkela_wire_13069)
    );

    bfr new_Jinkela_buffer_10745 (
        .din(new_Jinkela_wire_12950),
        .dout(new_Jinkela_wire_12951)
    );

    bfr new_Jinkela_buffer_10821 (
        .din(new_Jinkela_wire_13032),
        .dout(new_Jinkela_wire_13033)
    );

    bfr new_Jinkela_buffer_10746 (
        .din(new_Jinkela_wire_12951),
        .dout(new_Jinkela_wire_12952)
    );

    bfr new_Jinkela_buffer_10911 (
        .din(new_Jinkela_wire_13142),
        .dout(new_Jinkela_wire_13143)
    );

    spl2 new_Jinkela_splitter_966 (
        .a(_0282_),
        .b(new_Jinkela_wire_13149),
        .c(new_Jinkela_wire_13150)
    );

    bfr new_Jinkela_buffer_10747 (
        .din(new_Jinkela_wire_12952),
        .dout(new_Jinkela_wire_12953)
    );

    bfr new_Jinkela_buffer_10822 (
        .din(new_Jinkela_wire_13033),
        .dout(new_Jinkela_wire_13034)
    );

    bfr new_Jinkela_buffer_10748 (
        .din(new_Jinkela_wire_12953),
        .dout(new_Jinkela_wire_12954)
    );

    bfr new_Jinkela_buffer_10842 (
        .din(new_Jinkela_wire_13069),
        .dout(new_Jinkela_wire_13070)
    );

    bfr new_Jinkela_buffer_10749 (
        .din(new_Jinkela_wire_12954),
        .dout(new_Jinkela_wire_12955)
    );

    bfr new_Jinkela_buffer_10823 (
        .din(new_Jinkela_wire_13034),
        .dout(new_Jinkela_wire_13035)
    );

    bfr new_Jinkela_buffer_10750 (
        .din(new_Jinkela_wire_12955),
        .dout(new_Jinkela_wire_12956)
    );

    spl2 new_Jinkela_splitter_967 (
        .a(_1773_),
        .b(new_Jinkela_wire_13151),
        .c(new_Jinkela_wire_13152)
    );

    bfr new_Jinkela_buffer_10751 (
        .din(new_Jinkela_wire_12956),
        .dout(new_Jinkela_wire_12957)
    );

    bfr new_Jinkela_buffer_10824 (
        .din(new_Jinkela_wire_13035),
        .dout(new_Jinkela_wire_13036)
    );

    bfr new_Jinkela_buffer_10752 (
        .din(new_Jinkela_wire_12957),
        .dout(new_Jinkela_wire_12958)
    );

    bfr new_Jinkela_buffer_10843 (
        .din(new_Jinkela_wire_13070),
        .dout(new_Jinkela_wire_13071)
    );

    bfr new_Jinkela_buffer_10753 (
        .din(new_Jinkela_wire_12958),
        .dout(new_Jinkela_wire_12959)
    );

    bfr new_Jinkela_buffer_10825 (
        .din(new_Jinkela_wire_13036),
        .dout(new_Jinkela_wire_13037)
    );

    bfr new_Jinkela_buffer_10754 (
        .din(new_Jinkela_wire_12959),
        .dout(new_Jinkela_wire_12960)
    );

    bfr new_Jinkela_buffer_10912 (
        .din(new_Jinkela_wire_13143),
        .dout(new_Jinkela_wire_13144)
    );

    bfr new_Jinkela_buffer_10755 (
        .din(new_Jinkela_wire_12960),
        .dout(new_Jinkela_wire_12961)
    );

    bfr new_Jinkela_buffer_10826 (
        .din(new_Jinkela_wire_13037),
        .dout(new_Jinkela_wire_13038)
    );

    bfr new_Jinkela_buffer_10756 (
        .din(new_Jinkela_wire_12961),
        .dout(new_Jinkela_wire_12962)
    );

    bfr new_Jinkela_buffer_7481 (
        .din(_0450_),
        .dout(new_Jinkela_wire_9299)
    );

    bfr new_Jinkela_buffer_7255 (
        .din(new_Jinkela_wire_9046),
        .dout(new_Jinkela_wire_9047)
    );

    bfr new_Jinkela_buffer_7314 (
        .din(new_Jinkela_wire_9115),
        .dout(new_Jinkela_wire_9116)
    );

    bfr new_Jinkela_buffer_7256 (
        .din(new_Jinkela_wire_9047),
        .dout(new_Jinkela_wire_9048)
    );

    spl2 new_Jinkela_splitter_759 (
        .a(_1808_),
        .b(new_Jinkela_wire_9347),
        .c(new_Jinkela_wire_9348)
    );

    bfr new_Jinkela_buffer_7257 (
        .din(new_Jinkela_wire_9048),
        .dout(new_Jinkela_wire_9049)
    );

    bfr new_Jinkela_buffer_7315 (
        .din(new_Jinkela_wire_9116),
        .dout(new_Jinkela_wire_9117)
    );

    bfr new_Jinkela_buffer_7258 (
        .din(new_Jinkela_wire_9049),
        .dout(new_Jinkela_wire_9050)
    );

    bfr new_Jinkela_buffer_7372 (
        .din(new_Jinkela_wire_9187),
        .dout(new_Jinkela_wire_9188)
    );

    bfr new_Jinkela_buffer_7259 (
        .din(new_Jinkela_wire_9050),
        .dout(new_Jinkela_wire_9051)
    );

    bfr new_Jinkela_buffer_7316 (
        .din(new_Jinkela_wire_9117),
        .dout(new_Jinkela_wire_9118)
    );

    bfr new_Jinkela_buffer_7260 (
        .din(new_Jinkela_wire_9051),
        .dout(new_Jinkela_wire_9052)
    );

    bfr new_Jinkela_buffer_7527 (
        .din(_0607_),
        .dout(new_Jinkela_wire_9349)
    );

    bfr new_Jinkela_buffer_7261 (
        .din(new_Jinkela_wire_9052),
        .dout(new_Jinkela_wire_9053)
    );

    bfr new_Jinkela_buffer_7317 (
        .din(new_Jinkela_wire_9118),
        .dout(new_Jinkela_wire_9119)
    );

    bfr new_Jinkela_buffer_7262 (
        .din(new_Jinkela_wire_9053),
        .dout(new_Jinkela_wire_9054)
    );

    bfr new_Jinkela_buffer_7373 (
        .din(new_Jinkela_wire_9188),
        .dout(new_Jinkela_wire_9189)
    );

    bfr new_Jinkela_buffer_7263 (
        .din(new_Jinkela_wire_9054),
        .dout(new_Jinkela_wire_9055)
    );

    bfr new_Jinkela_buffer_7318 (
        .din(new_Jinkela_wire_9119),
        .dout(new_Jinkela_wire_9120)
    );

    bfr new_Jinkela_buffer_7264 (
        .din(new_Jinkela_wire_9055),
        .dout(new_Jinkela_wire_9056)
    );

    bfr new_Jinkela_buffer_7482 (
        .din(new_Jinkela_wire_9299),
        .dout(new_Jinkela_wire_9300)
    );

    bfr new_Jinkela_buffer_7265 (
        .din(new_Jinkela_wire_9056),
        .dout(new_Jinkela_wire_9057)
    );

    bfr new_Jinkela_buffer_7319 (
        .din(new_Jinkela_wire_9120),
        .dout(new_Jinkela_wire_9121)
    );

    bfr new_Jinkela_buffer_7266 (
        .din(new_Jinkela_wire_9057),
        .dout(new_Jinkela_wire_9058)
    );

    bfr new_Jinkela_buffer_7374 (
        .din(new_Jinkela_wire_9189),
        .dout(new_Jinkela_wire_9190)
    );

    bfr new_Jinkela_buffer_7267 (
        .din(new_Jinkela_wire_9058),
        .dout(new_Jinkela_wire_9059)
    );

    bfr new_Jinkela_buffer_7320 (
        .din(new_Jinkela_wire_9121),
        .dout(new_Jinkela_wire_9122)
    );

    bfr new_Jinkela_buffer_7268 (
        .din(new_Jinkela_wire_9059),
        .dout(new_Jinkela_wire_9060)
    );

    bfr new_Jinkela_buffer_7528 (
        .din(_0523_),
        .dout(new_Jinkela_wire_9350)
    );

    bfr new_Jinkela_buffer_7269 (
        .din(new_Jinkela_wire_9060),
        .dout(new_Jinkela_wire_9061)
    );

    bfr new_Jinkela_buffer_7321 (
        .din(new_Jinkela_wire_9122),
        .dout(new_Jinkela_wire_9123)
    );

    bfr new_Jinkela_buffer_7270 (
        .din(new_Jinkela_wire_9061),
        .dout(new_Jinkela_wire_9062)
    );

    bfr new_Jinkela_buffer_7375 (
        .din(new_Jinkela_wire_9190),
        .dout(new_Jinkela_wire_9191)
    );

    bfr new_Jinkela_buffer_7271 (
        .din(new_Jinkela_wire_9062),
        .dout(new_Jinkela_wire_9063)
    );

    bfr new_Jinkela_buffer_7322 (
        .din(new_Jinkela_wire_9123),
        .dout(new_Jinkela_wire_9124)
    );

    bfr new_Jinkela_buffer_7272 (
        .din(new_Jinkela_wire_9063),
        .dout(new_Jinkela_wire_9064)
    );

    bfr new_Jinkela_buffer_7483 (
        .din(new_Jinkela_wire_9300),
        .dout(new_Jinkela_wire_9301)
    );

    bfr new_Jinkela_buffer_7273 (
        .din(new_Jinkela_wire_9064),
        .dout(new_Jinkela_wire_9065)
    );

    bfr new_Jinkela_buffer_7323 (
        .din(new_Jinkela_wire_9124),
        .dout(new_Jinkela_wire_9125)
    );

    bfr new_Jinkela_buffer_7274 (
        .din(new_Jinkela_wire_9065),
        .dout(new_Jinkela_wire_9066)
    );

    bfr new_Jinkela_buffer_7376 (
        .din(new_Jinkela_wire_9191),
        .dout(new_Jinkela_wire_9192)
    );

    bfr new_Jinkela_buffer_7275 (
        .din(new_Jinkela_wire_9066),
        .dout(new_Jinkela_wire_9067)
    );

    bfr new_Jinkela_buffer_3841 (
        .din(new_Jinkela_wire_5076),
        .dout(new_Jinkela_wire_5077)
    );

    bfr new_Jinkela_buffer_3869 (
        .din(new_Jinkela_wire_5112),
        .dout(new_Jinkela_wire_5113)
    );

    bfr new_Jinkela_buffer_3842 (
        .din(new_Jinkela_wire_5077),
        .dout(new_Jinkela_wire_5078)
    );

    bfr new_Jinkela_buffer_3843 (
        .din(new_Jinkela_wire_5078),
        .dout(new_Jinkela_wire_5079)
    );

    bfr new_Jinkela_buffer_3870 (
        .din(new_Jinkela_wire_5113),
        .dout(new_Jinkela_wire_5114)
    );

    bfr new_Jinkela_buffer_3844 (
        .din(new_Jinkela_wire_5079),
        .dout(new_Jinkela_wire_5080)
    );

    spl2 new_Jinkela_splitter_476 (
        .a(_0595_),
        .b(new_Jinkela_wire_5142),
        .c(new_Jinkela_wire_5143)
    );

    bfr new_Jinkela_buffer_3884 (
        .din(new_Jinkela_wire_5137),
        .dout(new_Jinkela_wire_5138)
    );

    bfr new_Jinkela_buffer_3845 (
        .din(new_Jinkela_wire_5080),
        .dout(new_Jinkela_wire_5081)
    );

    bfr new_Jinkela_buffer_3871 (
        .din(new_Jinkela_wire_5114),
        .dout(new_Jinkela_wire_5115)
    );

    bfr new_Jinkela_buffer_3846 (
        .din(new_Jinkela_wire_5081),
        .dout(new_Jinkela_wire_5082)
    );

    spl2 new_Jinkela_splitter_475 (
        .a(_0358_),
        .b(new_Jinkela_wire_5136),
        .c(new_Jinkela_wire_5137)
    );

    bfr new_Jinkela_buffer_3847 (
        .din(new_Jinkela_wire_5082),
        .dout(new_Jinkela_wire_5083)
    );

    bfr new_Jinkela_buffer_3872 (
        .din(new_Jinkela_wire_5115),
        .dout(new_Jinkela_wire_5116)
    );

    bfr new_Jinkela_buffer_3848 (
        .din(new_Jinkela_wire_5083),
        .dout(new_Jinkela_wire_5084)
    );

    bfr new_Jinkela_buffer_3849 (
        .din(new_Jinkela_wire_5084),
        .dout(new_Jinkela_wire_5085)
    );

    bfr new_Jinkela_buffer_3873 (
        .din(new_Jinkela_wire_5116),
        .dout(new_Jinkela_wire_5117)
    );

    bfr new_Jinkela_buffer_3850 (
        .din(new_Jinkela_wire_5085),
        .dout(new_Jinkela_wire_5086)
    );

    spl2 new_Jinkela_splitter_477 (
        .a(_0585_),
        .b(new_Jinkela_wire_5144),
        .c(new_Jinkela_wire_5145)
    );

    bfr new_Jinkela_buffer_3851 (
        .din(new_Jinkela_wire_5086),
        .dout(new_Jinkela_wire_5087)
    );

    bfr new_Jinkela_buffer_3874 (
        .din(new_Jinkela_wire_5117),
        .dout(new_Jinkela_wire_5118)
    );

    bfr new_Jinkela_buffer_3852 (
        .din(new_Jinkela_wire_5087),
        .dout(new_Jinkela_wire_5088)
    );

    bfr new_Jinkela_buffer_3853 (
        .din(new_Jinkela_wire_5088),
        .dout(new_Jinkela_wire_5089)
    );

    bfr new_Jinkela_buffer_3875 (
        .din(new_Jinkela_wire_5118),
        .dout(new_Jinkela_wire_5119)
    );

    bfr new_Jinkela_buffer_3854 (
        .din(new_Jinkela_wire_5089),
        .dout(new_Jinkela_wire_5090)
    );

    bfr new_Jinkela_buffer_3885 (
        .din(new_Jinkela_wire_5138),
        .dout(new_Jinkela_wire_5139)
    );

    bfr new_Jinkela_buffer_3855 (
        .din(new_Jinkela_wire_5090),
        .dout(new_Jinkela_wire_5091)
    );

    bfr new_Jinkela_buffer_3876 (
        .din(new_Jinkela_wire_5119),
        .dout(new_Jinkela_wire_5120)
    );

    bfr new_Jinkela_buffer_3888 (
        .din(_0039_),
        .dout(new_Jinkela_wire_5146)
    );

    bfr new_Jinkela_buffer_3877 (
        .din(new_Jinkela_wire_5120),
        .dout(new_Jinkela_wire_5121)
    );

    bfr new_Jinkela_buffer_3886 (
        .din(new_Jinkela_wire_5139),
        .dout(new_Jinkela_wire_5140)
    );

    bfr new_Jinkela_buffer_3878 (
        .din(new_Jinkela_wire_5121),
        .dout(new_Jinkela_wire_5122)
    );

    spl2 new_Jinkela_splitter_479 (
        .a(_0704_),
        .b(new_Jinkela_wire_5149),
        .c(new_Jinkela_wire_5150)
    );

    spl2 new_Jinkela_splitter_478 (
        .a(_1246_),
        .b(new_Jinkela_wire_5147),
        .c(new_Jinkela_wire_5148)
    );

    bfr new_Jinkela_buffer_3879 (
        .din(new_Jinkela_wire_5122),
        .dout(new_Jinkela_wire_5123)
    );

    bfr new_Jinkela_buffer_3887 (
        .din(new_Jinkela_wire_5140),
        .dout(new_Jinkela_wire_5141)
    );

    spl2 new_Jinkela_splitter_471 (
        .a(new_Jinkela_wire_5123),
        .b(new_Jinkela_wire_5124),
        .c(new_Jinkela_wire_5125)
    );

    spl2 new_Jinkela_splitter_480 (
        .a(_1697_),
        .b(new_Jinkela_wire_5151),
        .c(new_Jinkela_wire_5152)
    );

    bfr new_Jinkela_buffer_3893 (
        .din(_1594_),
        .dout(new_Jinkela_wire_5157)
    );

    bfr new_Jinkela_buffer_3889 (
        .din(new_Jinkela_wire_5152),
        .dout(new_Jinkela_wire_5153)
    );

    spl2 new_Jinkela_splitter_481 (
        .a(_0569_),
        .b(new_Jinkela_wire_5158),
        .c(new_Jinkela_wire_5159)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_10844 (
        .din(new_Jinkela_wire_13071),
        .dout(new_Jinkela_wire_13072)
    );

    bfr new_Jinkela_buffer_10757 (
        .din(new_Jinkela_wire_12962),
        .dout(new_Jinkela_wire_12963)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_10827 (
        .din(new_Jinkela_wire_13038),
        .dout(new_Jinkela_wire_13039)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_10758 (
        .din(new_Jinkela_wire_12963),
        .dout(new_Jinkela_wire_12964)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    spl2 new_Jinkela_splitter_970 (
        .a(_1186_),
        .b(new_Jinkela_wire_13195),
        .c(new_Jinkela_wire_13196)
    );

    bfr new_Jinkela_buffer_10759 (
        .din(new_Jinkela_wire_12964),
        .dout(new_Jinkela_wire_12965)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_10828 (
        .din(new_Jinkela_wire_13039),
        .dout(new_Jinkela_wire_13040)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(_0248_),
        .b(new_Jinkela_wire_1256),
        .c(new_Jinkela_wire_1257)
    );

    bfr new_Jinkela_buffer_10760 (
        .din(new_Jinkela_wire_12965),
        .dout(new_Jinkela_wire_12966)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_1030),
        .dout(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    bfr new_Jinkela_buffer_10845 (
        .din(new_Jinkela_wire_13072),
        .dout(new_Jinkela_wire_13073)
    );

    bfr new_Jinkela_buffer_10761 (
        .din(new_Jinkela_wire_12966),
        .dout(new_Jinkela_wire_12967)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_1140),
        .dout(new_Jinkela_wire_1141)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_10829 (
        .din(new_Jinkela_wire_13040),
        .dout(new_Jinkela_wire_13041)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    bfr new_Jinkela_buffer_10762 (
        .din(new_Jinkela_wire_12967),
        .dout(new_Jinkela_wire_12968)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_10913 (
        .din(new_Jinkela_wire_13144),
        .dout(new_Jinkela_wire_13145)
    );

    bfr new_Jinkela_buffer_10763 (
        .din(new_Jinkela_wire_12968),
        .dout(new_Jinkela_wire_12969)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_10830 (
        .din(new_Jinkela_wire_13041),
        .dout(new_Jinkela_wire_13042)
    );

    bfr new_Jinkela_buffer_10764 (
        .din(new_Jinkela_wire_12969),
        .dout(new_Jinkela_wire_12970)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_10846 (
        .din(new_Jinkela_wire_13073),
        .dout(new_Jinkela_wire_13074)
    );

    bfr new_Jinkela_buffer_10765 (
        .din(new_Jinkela_wire_12970),
        .dout(new_Jinkela_wire_12971)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_10831 (
        .din(new_Jinkela_wire_13042),
        .dout(new_Jinkela_wire_13043)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_1084),
        .dout(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_10766 (
        .din(new_Jinkela_wire_12971),
        .dout(new_Jinkela_wire_12972)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_10915 (
        .din(_1018_),
        .dout(new_Jinkela_wire_13153)
    );

    bfr new_Jinkela_buffer_10767 (
        .din(new_Jinkela_wire_12972),
        .dout(new_Jinkela_wire_12973)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_10832 (
        .din(new_Jinkela_wire_13043),
        .dout(new_Jinkela_wire_13044)
    );

    bfr new_Jinkela_buffer_10768 (
        .din(new_Jinkela_wire_12973),
        .dout(new_Jinkela_wire_12974)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_10847 (
        .din(new_Jinkela_wire_13074),
        .dout(new_Jinkela_wire_13075)
    );

    bfr new_Jinkela_buffer_10769 (
        .din(new_Jinkela_wire_12974),
        .dout(new_Jinkela_wire_12975)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_1141),
        .dout(new_Jinkela_wire_1142)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    spl2 new_Jinkela_splitter_955 (
        .a(new_Jinkela_wire_13044),
        .b(new_Jinkela_wire_13045),
        .c(new_Jinkela_wire_13046)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_1085),
        .dout(new_Jinkela_wire_1086)
    );

    bfr new_Jinkela_buffer_10770 (
        .din(new_Jinkela_wire_12975),
        .dout(new_Jinkela_wire_12976)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_10848 (
        .din(new_Jinkela_wire_13075),
        .dout(new_Jinkela_wire_13076)
    );

    bfr new_Jinkela_buffer_10771 (
        .din(new_Jinkela_wire_12976),
        .dout(new_Jinkela_wire_12977)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    bfr new_Jinkela_buffer_10914 (
        .din(new_Jinkela_wire_13145),
        .dout(new_Jinkela_wire_13146)
    );

    bfr new_Jinkela_buffer_10772 (
        .din(new_Jinkela_wire_12977),
        .dout(new_Jinkela_wire_12978)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_10916 (
        .din(_0032_),
        .dout(new_Jinkela_wire_13156)
    );

    spl2 new_Jinkela_splitter_968 (
        .a(_1790_),
        .b(new_Jinkela_wire_13154),
        .c(new_Jinkela_wire_13155)
    );

    bfr new_Jinkela_buffer_10773 (
        .din(new_Jinkela_wire_12978),
        .dout(new_Jinkela_wire_12979)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(_0401_),
        .b(new_Jinkela_wire_1259),
        .c(new_Jinkela_wire_1260)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_10849 (
        .din(new_Jinkela_wire_13076),
        .dout(new_Jinkela_wire_13077)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_1086),
        .dout(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_10774 (
        .din(new_Jinkela_wire_12979),
        .dout(new_Jinkela_wire_12980)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_10775 (
        .din(new_Jinkela_wire_12980),
        .dout(new_Jinkela_wire_12981)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_10850 (
        .din(new_Jinkela_wire_13077),
        .dout(new_Jinkela_wire_13078)
    );

    bfr new_Jinkela_buffer_542 (
        .din(_1510_),
        .dout(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_10776 (
        .din(new_Jinkela_wire_12981),
        .dout(new_Jinkela_wire_12982)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_10917 (
        .din(_0920_),
        .dout(new_Jinkela_wire_13157)
    );

    bfr new_Jinkela_buffer_10777 (
        .din(new_Jinkela_wire_12982),
        .dout(new_Jinkela_wire_12983)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_1142),
        .dout(new_Jinkela_wire_1143)
    );

    bfr new_Jinkela_buffer_14231 (
        .din(new_Jinkela_wire_16978),
        .dout(new_Jinkela_wire_16979)
    );

    bfr new_Jinkela_buffer_14251 (
        .din(new_Jinkela_wire_17002),
        .dout(new_Jinkela_wire_17003)
    );

    bfr new_Jinkela_buffer_14232 (
        .din(new_Jinkela_wire_16979),
        .dout(new_Jinkela_wire_16980)
    );

    bfr new_Jinkela_buffer_14258 (
        .din(new_Jinkela_wire_17017),
        .dout(new_Jinkela_wire_17018)
    );

    bfr new_Jinkela_buffer_14233 (
        .din(new_Jinkela_wire_16980),
        .dout(new_Jinkela_wire_16981)
    );

    bfr new_Jinkela_buffer_14252 (
        .din(new_Jinkela_wire_17003),
        .dout(new_Jinkela_wire_17004)
    );

    bfr new_Jinkela_buffer_14234 (
        .din(new_Jinkela_wire_16981),
        .dout(new_Jinkela_wire_16982)
    );

    bfr new_Jinkela_buffer_14254 (
        .din(new_Jinkela_wire_17007),
        .dout(new_Jinkela_wire_17008)
    );

    bfr new_Jinkela_buffer_14235 (
        .din(new_Jinkela_wire_16982),
        .dout(new_Jinkela_wire_16983)
    );

    bfr new_Jinkela_buffer_14257 (
        .din(_1766_),
        .dout(new_Jinkela_wire_17015)
    );

    bfr new_Jinkela_buffer_14236 (
        .din(new_Jinkela_wire_16983),
        .dout(new_Jinkela_wire_16984)
    );

    bfr new_Jinkela_buffer_14255 (
        .din(new_Jinkela_wire_17008),
        .dout(new_Jinkela_wire_17009)
    );

    bfr new_Jinkela_buffer_14237 (
        .din(new_Jinkela_wire_16984),
        .dout(new_Jinkela_wire_16985)
    );

    spl2 new_Jinkela_splitter_1229 (
        .a(_0090_),
        .b(new_Jinkela_wire_17022),
        .c(new_Jinkela_wire_17023)
    );

    spl2 new_Jinkela_splitter_1228 (
        .a(_0005_),
        .b(new_Jinkela_wire_17016),
        .c(new_Jinkela_wire_17017)
    );

    bfr new_Jinkela_buffer_14238 (
        .din(new_Jinkela_wire_16985),
        .dout(new_Jinkela_wire_16986)
    );

    bfr new_Jinkela_buffer_14256 (
        .din(new_Jinkela_wire_17009),
        .dout(new_Jinkela_wire_17010)
    );

    bfr new_Jinkela_buffer_14239 (
        .din(new_Jinkela_wire_16986),
        .dout(new_Jinkela_wire_16987)
    );

    bfr new_Jinkela_buffer_14240 (
        .din(new_Jinkela_wire_16987),
        .dout(new_Jinkela_wire_16988)
    );

    spl2 new_Jinkela_splitter_1230 (
        .a(_0804_),
        .b(new_Jinkela_wire_17024),
        .c(new_Jinkela_wire_17025)
    );

    bfr new_Jinkela_buffer_14241 (
        .din(new_Jinkela_wire_16988),
        .dout(new_Jinkela_wire_16989)
    );

    bfr new_Jinkela_buffer_14242 (
        .din(new_Jinkela_wire_16989),
        .dout(new_Jinkela_wire_16990)
    );

    bfr new_Jinkela_buffer_14259 (
        .din(new_Jinkela_wire_17018),
        .dout(new_Jinkela_wire_17019)
    );

    bfr new_Jinkela_buffer_14243 (
        .din(new_Jinkela_wire_16990),
        .dout(new_Jinkela_wire_16991)
    );

    spl2 new_Jinkela_splitter_1231 (
        .a(_0384_),
        .b(new_Jinkela_wire_17026),
        .c(new_Jinkela_wire_17027)
    );

    bfr new_Jinkela_buffer_14244 (
        .din(new_Jinkela_wire_16991),
        .dout(new_Jinkela_wire_16992)
    );

    bfr new_Jinkela_buffer_14260 (
        .din(new_Jinkela_wire_17019),
        .dout(new_Jinkela_wire_17020)
    );

    bfr new_Jinkela_buffer_14245 (
        .din(new_Jinkela_wire_16992),
        .dout(new_Jinkela_wire_16993)
    );

    spl2 new_Jinkela_splitter_1232 (
        .a(_0008_),
        .b(new_Jinkela_wire_17028),
        .c(new_Jinkela_wire_17029)
    );

    bfr new_Jinkela_buffer_14246 (
        .din(new_Jinkela_wire_16993),
        .dout(new_Jinkela_wire_16994)
    );

    bfr new_Jinkela_buffer_14261 (
        .din(new_Jinkela_wire_17020),
        .dout(new_Jinkela_wire_17021)
    );

    bfr new_Jinkela_buffer_14247 (
        .din(new_Jinkela_wire_16994),
        .dout(new_Jinkela_wire_16995)
    );

    bfr new_Jinkela_buffer_14263 (
        .din(new_Jinkela_wire_17032),
        .dout(new_Jinkela_wire_17033)
    );

    bfr new_Jinkela_buffer_14262 (
        .din(_1309_),
        .dout(new_Jinkela_wire_17030)
    );

    bfr new_Jinkela_buffer_14248 (
        .din(new_Jinkela_wire_16995),
        .dout(new_Jinkela_wire_16996)
    );

    spl2 new_Jinkela_splitter_1234 (
        .a(_0165_),
        .b(new_Jinkela_wire_17037),
        .c(new_Jinkela_wire_17038)
    );

    spl2 new_Jinkela_splitter_1233 (
        .a(_1160_),
        .b(new_Jinkela_wire_17031),
        .c(new_Jinkela_wire_17032)
    );

    spl2 new_Jinkela_splitter_1223 (
        .a(new_Jinkela_wire_16996),
        .b(new_Jinkela_wire_16997),
        .c(new_Jinkela_wire_16998)
    );

    spl2 new_Jinkela_splitter_1235 (
        .a(_1438_),
        .b(new_Jinkela_wire_17043),
        .c(new_Jinkela_wire_17044)
    );

    bfr new_Jinkela_buffer_14264 (
        .din(new_Jinkela_wire_17033),
        .dout(new_Jinkela_wire_17034)
    );

    bfr new_Jinkela_buffer_14267 (
        .din(new_Jinkela_wire_17038),
        .dout(new_Jinkela_wire_17039)
    );

    spl2 new_Jinkela_splitter_1236 (
        .a(_1027_),
        .b(new_Jinkela_wire_17045),
        .c(new_Jinkela_wire_17046)
    );

    bfr new_Jinkela_buffer_7324 (
        .din(new_Jinkela_wire_9125),
        .dout(new_Jinkela_wire_9126)
    );

    bfr new_Jinkela_buffer_7276 (
        .din(new_Jinkela_wire_9067),
        .dout(new_Jinkela_wire_9068)
    );

    bfr new_Jinkela_buffer_7540 (
        .din(_0221_),
        .dout(new_Jinkela_wire_9364)
    );

    bfr new_Jinkela_buffer_7277 (
        .din(new_Jinkela_wire_9068),
        .dout(new_Jinkela_wire_9069)
    );

    bfr new_Jinkela_buffer_7325 (
        .din(new_Jinkela_wire_9126),
        .dout(new_Jinkela_wire_9127)
    );

    bfr new_Jinkela_buffer_7278 (
        .din(new_Jinkela_wire_9069),
        .dout(new_Jinkela_wire_9070)
    );

    bfr new_Jinkela_buffer_7377 (
        .din(new_Jinkela_wire_9192),
        .dout(new_Jinkela_wire_9193)
    );

    bfr new_Jinkela_buffer_7279 (
        .din(new_Jinkela_wire_9070),
        .dout(new_Jinkela_wire_9071)
    );

    bfr new_Jinkela_buffer_7326 (
        .din(new_Jinkela_wire_9127),
        .dout(new_Jinkela_wire_9128)
    );

    bfr new_Jinkela_buffer_7280 (
        .din(new_Jinkela_wire_9071),
        .dout(new_Jinkela_wire_9072)
    );

    bfr new_Jinkela_buffer_7484 (
        .din(new_Jinkela_wire_9301),
        .dout(new_Jinkela_wire_9302)
    );

    bfr new_Jinkela_buffer_7281 (
        .din(new_Jinkela_wire_9072),
        .dout(new_Jinkela_wire_9073)
    );

    bfr new_Jinkela_buffer_7327 (
        .din(new_Jinkela_wire_9128),
        .dout(new_Jinkela_wire_9129)
    );

    bfr new_Jinkela_buffer_7282 (
        .din(new_Jinkela_wire_9073),
        .dout(new_Jinkela_wire_9074)
    );

    bfr new_Jinkela_buffer_7378 (
        .din(new_Jinkela_wire_9193),
        .dout(new_Jinkela_wire_9194)
    );

    bfr new_Jinkela_buffer_7283 (
        .din(new_Jinkela_wire_9074),
        .dout(new_Jinkela_wire_9075)
    );

    bfr new_Jinkela_buffer_7328 (
        .din(new_Jinkela_wire_9129),
        .dout(new_Jinkela_wire_9130)
    );

    bfr new_Jinkela_buffer_7284 (
        .din(new_Jinkela_wire_9075),
        .dout(new_Jinkela_wire_9076)
    );

    spl2 new_Jinkela_splitter_762 (
        .a(_1005_),
        .b(new_Jinkela_wire_9446),
        .c(new_Jinkela_wire_9447)
    );

    bfr new_Jinkela_buffer_7285 (
        .din(new_Jinkela_wire_9076),
        .dout(new_Jinkela_wire_9077)
    );

    bfr new_Jinkela_buffer_7329 (
        .din(new_Jinkela_wire_9130),
        .dout(new_Jinkela_wire_9131)
    );

    bfr new_Jinkela_buffer_7286 (
        .din(new_Jinkela_wire_9077),
        .dout(new_Jinkela_wire_9078)
    );

    bfr new_Jinkela_buffer_7379 (
        .din(new_Jinkela_wire_9194),
        .dout(new_Jinkela_wire_9195)
    );

    bfr new_Jinkela_buffer_7287 (
        .din(new_Jinkela_wire_9078),
        .dout(new_Jinkela_wire_9079)
    );

    bfr new_Jinkela_buffer_7330 (
        .din(new_Jinkela_wire_9131),
        .dout(new_Jinkela_wire_9132)
    );

    bfr new_Jinkela_buffer_7288 (
        .din(new_Jinkela_wire_9079),
        .dout(new_Jinkela_wire_9080)
    );

    bfr new_Jinkela_buffer_7485 (
        .din(new_Jinkela_wire_9302),
        .dout(new_Jinkela_wire_9303)
    );

    bfr new_Jinkela_buffer_7289 (
        .din(new_Jinkela_wire_9080),
        .dout(new_Jinkela_wire_9081)
    );

    bfr new_Jinkela_buffer_7331 (
        .din(new_Jinkela_wire_9132),
        .dout(new_Jinkela_wire_9133)
    );

    bfr new_Jinkela_buffer_7290 (
        .din(new_Jinkela_wire_9081),
        .dout(new_Jinkela_wire_9082)
    );

    bfr new_Jinkela_buffer_7380 (
        .din(new_Jinkela_wire_9195),
        .dout(new_Jinkela_wire_9196)
    );

    bfr new_Jinkela_buffer_7291 (
        .din(new_Jinkela_wire_9082),
        .dout(new_Jinkela_wire_9083)
    );

    bfr new_Jinkela_buffer_7332 (
        .din(new_Jinkela_wire_9133),
        .dout(new_Jinkela_wire_9134)
    );

    bfr new_Jinkela_buffer_7292 (
        .din(new_Jinkela_wire_9083),
        .dout(new_Jinkela_wire_9084)
    );

    bfr new_Jinkela_buffer_7529 (
        .din(new_Jinkela_wire_9350),
        .dout(new_Jinkela_wire_9351)
    );

    bfr new_Jinkela_buffer_7293 (
        .din(new_Jinkela_wire_9084),
        .dout(new_Jinkela_wire_9085)
    );

    bfr new_Jinkela_buffer_7333 (
        .din(new_Jinkela_wire_9134),
        .dout(new_Jinkela_wire_9135)
    );

    bfr new_Jinkela_buffer_7294 (
        .din(new_Jinkela_wire_9085),
        .dout(new_Jinkela_wire_9086)
    );

    bfr new_Jinkela_buffer_7381 (
        .din(new_Jinkela_wire_9196),
        .dout(new_Jinkela_wire_9197)
    );

    bfr new_Jinkela_buffer_7295 (
        .din(new_Jinkela_wire_9086),
        .dout(new_Jinkela_wire_9087)
    );

    bfr new_Jinkela_buffer_7334 (
        .din(new_Jinkela_wire_9135),
        .dout(new_Jinkela_wire_9136)
    );

    bfr new_Jinkela_buffer_7296 (
        .din(new_Jinkela_wire_9087),
        .dout(new_Jinkela_wire_9088)
    );

    bfr new_Jinkela_buffer_17645 (
        .din(new_Jinkela_wire_21013),
        .dout(new_Jinkela_wire_21014)
    );

    spl2 new_Jinkela_splitter_1544 (
        .a(_0361_),
        .b(new_Jinkela_wire_21146),
        .c(new_Jinkela_wire_21147)
    );

    bfr new_Jinkela_buffer_17735 (
        .din(new_Jinkela_wire_21125),
        .dout(new_Jinkela_wire_21126)
    );

    bfr new_Jinkela_buffer_17646 (
        .din(new_Jinkela_wire_21014),
        .dout(new_Jinkela_wire_21015)
    );

    bfr new_Jinkela_buffer_17731 (
        .din(new_Jinkela_wire_21119),
        .dout(new_Jinkela_wire_21120)
    );

    bfr new_Jinkela_buffer_17647 (
        .din(new_Jinkela_wire_21015),
        .dout(new_Jinkela_wire_21016)
    );

    bfr new_Jinkela_buffer_17648 (
        .din(new_Jinkela_wire_21016),
        .dout(new_Jinkela_wire_21017)
    );

    bfr new_Jinkela_buffer_17732 (
        .din(new_Jinkela_wire_21120),
        .dout(new_Jinkela_wire_21121)
    );

    bfr new_Jinkela_buffer_17649 (
        .din(new_Jinkela_wire_21017),
        .dout(new_Jinkela_wire_21018)
    );

    bfr new_Jinkela_buffer_17756 (
        .din(_0903_),
        .dout(new_Jinkela_wire_21151)
    );

    bfr new_Jinkela_buffer_17650 (
        .din(new_Jinkela_wire_21018),
        .dout(new_Jinkela_wire_21019)
    );

    bfr new_Jinkela_buffer_17733 (
        .din(new_Jinkela_wire_21121),
        .dout(new_Jinkela_wire_21122)
    );

    bfr new_Jinkela_buffer_17651 (
        .din(new_Jinkela_wire_21019),
        .dout(new_Jinkela_wire_21020)
    );

    spl2 new_Jinkela_splitter_1548 (
        .a(_0123_),
        .b(new_Jinkela_wire_21162),
        .c(new_Jinkela_wire_21163)
    );

    bfr new_Jinkela_buffer_17652 (
        .din(new_Jinkela_wire_21020),
        .dout(new_Jinkela_wire_21021)
    );

    bfr new_Jinkela_buffer_17736 (
        .din(new_Jinkela_wire_21126),
        .dout(new_Jinkela_wire_21127)
    );

    bfr new_Jinkela_buffer_17653 (
        .din(new_Jinkela_wire_21021),
        .dout(new_Jinkela_wire_21022)
    );

    bfr new_Jinkela_buffer_17755 (
        .din(new_Jinkela_wire_21147),
        .dout(new_Jinkela_wire_21148)
    );

    bfr new_Jinkela_buffer_17758 (
        .din(_1776_),
        .dout(new_Jinkela_wire_21155)
    );

    bfr new_Jinkela_buffer_17654 (
        .din(new_Jinkela_wire_21022),
        .dout(new_Jinkela_wire_21023)
    );

    bfr new_Jinkela_buffer_17737 (
        .din(new_Jinkela_wire_21127),
        .dout(new_Jinkela_wire_21128)
    );

    bfr new_Jinkela_buffer_17655 (
        .din(new_Jinkela_wire_21023),
        .dout(new_Jinkela_wire_21024)
    );

    bfr new_Jinkela_buffer_17757 (
        .din(new_Jinkela_wire_21151),
        .dout(new_Jinkela_wire_21152)
    );

    bfr new_Jinkela_buffer_17656 (
        .din(new_Jinkela_wire_21024),
        .dout(new_Jinkela_wire_21025)
    );

    bfr new_Jinkela_buffer_17738 (
        .din(new_Jinkela_wire_21128),
        .dout(new_Jinkela_wire_21129)
    );

    bfr new_Jinkela_buffer_17657 (
        .din(new_Jinkela_wire_21025),
        .dout(new_Jinkela_wire_21026)
    );

    spl2 new_Jinkela_splitter_1545 (
        .a(new_Jinkela_wire_21148),
        .b(new_Jinkela_wire_21149),
        .c(new_Jinkela_wire_21150)
    );

    bfr new_Jinkela_buffer_17658 (
        .din(new_Jinkela_wire_21026),
        .dout(new_Jinkela_wire_21027)
    );

    bfr new_Jinkela_buffer_17739 (
        .din(new_Jinkela_wire_21129),
        .dout(new_Jinkela_wire_21130)
    );

    bfr new_Jinkela_buffer_17659 (
        .din(new_Jinkela_wire_21027),
        .dout(new_Jinkela_wire_21028)
    );

    bfr new_Jinkela_buffer_17759 (
        .din(_0321_),
        .dout(new_Jinkela_wire_21156)
    );

    bfr new_Jinkela_buffer_17660 (
        .din(new_Jinkela_wire_21028),
        .dout(new_Jinkela_wire_21029)
    );

    bfr new_Jinkela_buffer_17740 (
        .din(new_Jinkela_wire_21130),
        .dout(new_Jinkela_wire_21131)
    );

    bfr new_Jinkela_buffer_17661 (
        .din(new_Jinkela_wire_21029),
        .dout(new_Jinkela_wire_21030)
    );

    spl2 new_Jinkela_splitter_1546 (
        .a(new_Jinkela_wire_21152),
        .b(new_Jinkela_wire_21153),
        .c(new_Jinkela_wire_21154)
    );

    bfr new_Jinkela_buffer_17662 (
        .din(new_Jinkela_wire_21030),
        .dout(new_Jinkela_wire_21031)
    );

    bfr new_Jinkela_buffer_17741 (
        .din(new_Jinkela_wire_21131),
        .dout(new_Jinkela_wire_21132)
    );

    bfr new_Jinkela_buffer_17663 (
        .din(new_Jinkela_wire_21031),
        .dout(new_Jinkela_wire_21032)
    );

    bfr new_Jinkela_buffer_17664 (
        .din(new_Jinkela_wire_21032),
        .dout(new_Jinkela_wire_21033)
    );

    bfr new_Jinkela_buffer_17742 (
        .din(new_Jinkela_wire_21132),
        .dout(new_Jinkela_wire_21133)
    );

    bfr new_Jinkela_buffer_17665 (
        .din(new_Jinkela_wire_21033),
        .dout(new_Jinkela_wire_21034)
    );

    spl2 new_Jinkela_splitter_1549 (
        .a(_0276_),
        .b(new_Jinkela_wire_21164),
        .c(new_Jinkela_wire_21165)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_1087),
        .dout(new_Jinkela_wire_1088)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_1039),
        .dout(new_Jinkela_wire_1040)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_1040),
        .dout(new_Jinkela_wire_1041)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(_1273_),
        .b(new_Jinkela_wire_1261),
        .c(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_1088),
        .dout(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_1041),
        .dout(new_Jinkela_wire_1042)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_937),
        .dout(new_Jinkela_wire_938)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(_1748_),
        .b(new_Jinkela_wire_1267),
        .c(new_Jinkela_wire_1268)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_1042),
        .dout(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_1143),
        .dout(new_Jinkela_wire_1144)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_1089),
        .dout(new_Jinkela_wire_1090)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_1044),
        .dout(new_Jinkela_wire_1045)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_1090),
        .dout(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_1045),
        .dout(new_Jinkela_wire_1046)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_1046),
        .dout(new_Jinkela_wire_1047)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_1144),
        .dout(new_Jinkela_wire_1145)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_948),
        .dout(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_1091),
        .dout(new_Jinkela_wire_1092)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_1047),
        .dout(new_Jinkela_wire_1048)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_1048),
        .dout(new_Jinkela_wire_1049)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_951),
        .dout(new_Jinkela_wire_952)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_952),
        .dout(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_1049),
        .dout(new_Jinkela_wire_1050)
    );

    bfr new_Jinkela_buffer_10851 (
        .din(new_Jinkela_wire_13078),
        .dout(new_Jinkela_wire_13079)
    );

    bfr new_Jinkela_buffer_10778 (
        .din(new_Jinkela_wire_12983),
        .dout(new_Jinkela_wire_12984)
    );

    bfr new_Jinkela_buffer_10953 (
        .din(_0399_),
        .dout(new_Jinkela_wire_13197)
    );

    bfr new_Jinkela_buffer_10779 (
        .din(new_Jinkela_wire_12984),
        .dout(new_Jinkela_wire_12985)
    );

    bfr new_Jinkela_buffer_10852 (
        .din(new_Jinkela_wire_13079),
        .dout(new_Jinkela_wire_13080)
    );

    bfr new_Jinkela_buffer_10780 (
        .din(new_Jinkela_wire_12985),
        .dout(new_Jinkela_wire_12986)
    );

    bfr new_Jinkela_buffer_10918 (
        .din(new_Jinkela_wire_13157),
        .dout(new_Jinkela_wire_13158)
    );

    bfr new_Jinkela_buffer_10781 (
        .din(new_Jinkela_wire_12986),
        .dout(new_Jinkela_wire_12987)
    );

    bfr new_Jinkela_buffer_10853 (
        .din(new_Jinkela_wire_13080),
        .dout(new_Jinkela_wire_13081)
    );

    bfr new_Jinkela_buffer_10782 (
        .din(new_Jinkela_wire_12987),
        .dout(new_Jinkela_wire_12988)
    );

    spl2 new_Jinkela_splitter_971 (
        .a(_1538_),
        .b(new_Jinkela_wire_13199),
        .c(new_Jinkela_wire_13200)
    );

    bfr new_Jinkela_buffer_10783 (
        .din(new_Jinkela_wire_12988),
        .dout(new_Jinkela_wire_12989)
    );

    bfr new_Jinkela_buffer_10854 (
        .din(new_Jinkela_wire_13081),
        .dout(new_Jinkela_wire_13082)
    );

    bfr new_Jinkela_buffer_10784 (
        .din(new_Jinkela_wire_12989),
        .dout(new_Jinkela_wire_12990)
    );

    bfr new_Jinkela_buffer_10919 (
        .din(new_Jinkela_wire_13158),
        .dout(new_Jinkela_wire_13159)
    );

    bfr new_Jinkela_buffer_10785 (
        .din(new_Jinkela_wire_12990),
        .dout(new_Jinkela_wire_12991)
    );

    bfr new_Jinkela_buffer_10855 (
        .din(new_Jinkela_wire_13082),
        .dout(new_Jinkela_wire_13083)
    );

    bfr new_Jinkela_buffer_10786 (
        .din(new_Jinkela_wire_12991),
        .dout(new_Jinkela_wire_12992)
    );

    bfr new_Jinkela_buffer_10954 (
        .din(_0379_),
        .dout(new_Jinkela_wire_13198)
    );

    bfr new_Jinkela_buffer_10787 (
        .din(new_Jinkela_wire_12992),
        .dout(new_Jinkela_wire_12993)
    );

    bfr new_Jinkela_buffer_10856 (
        .din(new_Jinkela_wire_13083),
        .dout(new_Jinkela_wire_13084)
    );

    bfr new_Jinkela_buffer_10788 (
        .din(new_Jinkela_wire_12993),
        .dout(new_Jinkela_wire_12994)
    );

    bfr new_Jinkela_buffer_10920 (
        .din(new_Jinkela_wire_13159),
        .dout(new_Jinkela_wire_13160)
    );

    bfr new_Jinkela_buffer_10789 (
        .din(new_Jinkela_wire_12994),
        .dout(new_Jinkela_wire_12995)
    );

    bfr new_Jinkela_buffer_10857 (
        .din(new_Jinkela_wire_13084),
        .dout(new_Jinkela_wire_13085)
    );

    bfr new_Jinkela_buffer_10790 (
        .din(new_Jinkela_wire_12995),
        .dout(new_Jinkela_wire_12996)
    );

    spl2 new_Jinkela_splitter_972 (
        .a(_1395_),
        .b(new_Jinkela_wire_13201),
        .c(new_Jinkela_wire_13202)
    );

    spl2 new_Jinkela_splitter_974 (
        .a(_1453_),
        .b(new_Jinkela_wire_13205),
        .c(new_Jinkela_wire_13206)
    );

    bfr new_Jinkela_buffer_10791 (
        .din(new_Jinkela_wire_12996),
        .dout(new_Jinkela_wire_12997)
    );

    bfr new_Jinkela_buffer_10858 (
        .din(new_Jinkela_wire_13085),
        .dout(new_Jinkela_wire_13086)
    );

    bfr new_Jinkela_buffer_10792 (
        .din(new_Jinkela_wire_12997),
        .dout(new_Jinkela_wire_12998)
    );

    bfr new_Jinkela_buffer_10921 (
        .din(new_Jinkela_wire_13160),
        .dout(new_Jinkela_wire_13161)
    );

    bfr new_Jinkela_buffer_10793 (
        .din(new_Jinkela_wire_12998),
        .dout(new_Jinkela_wire_12999)
    );

    bfr new_Jinkela_buffer_10859 (
        .din(new_Jinkela_wire_13086),
        .dout(new_Jinkela_wire_13087)
    );

    bfr new_Jinkela_buffer_10794 (
        .din(new_Jinkela_wire_12999),
        .dout(new_Jinkela_wire_13000)
    );

    bfr new_Jinkela_buffer_10795 (
        .din(new_Jinkela_wire_13000),
        .dout(new_Jinkela_wire_13001)
    );

    bfr new_Jinkela_buffer_10860 (
        .din(new_Jinkela_wire_13087),
        .dout(new_Jinkela_wire_13088)
    );

    bfr new_Jinkela_buffer_10796 (
        .din(new_Jinkela_wire_13001),
        .dout(new_Jinkela_wire_13002)
    );

    bfr new_Jinkela_buffer_10922 (
        .din(new_Jinkela_wire_13161),
        .dout(new_Jinkela_wire_13162)
    );

    spl2 new_Jinkela_splitter_952 (
        .a(new_Jinkela_wire_13002),
        .b(new_Jinkela_wire_13003),
        .c(new_Jinkela_wire_13004)
    );

    spl2 new_Jinkela_splitter_973 (
        .a(_1492_),
        .b(new_Jinkela_wire_13203),
        .c(new_Jinkela_wire_13204)
    );

    bfr new_Jinkela_buffer_10861 (
        .din(new_Jinkela_wire_13088),
        .dout(new_Jinkela_wire_13089)
    );

    bfr new_Jinkela_buffer_3894 (
        .din(_0466_),
        .dout(new_Jinkela_wire_5160)
    );

    bfr new_Jinkela_buffer_3899 (
        .din(_1068_),
        .dout(new_Jinkela_wire_5167)
    );

    bfr new_Jinkela_buffer_3890 (
        .din(new_Jinkela_wire_5153),
        .dout(new_Jinkela_wire_5154)
    );

    bfr new_Jinkela_buffer_3895 (
        .din(new_Jinkela_wire_5162),
        .dout(new_Jinkela_wire_5163)
    );

    bfr new_Jinkela_buffer_3891 (
        .din(new_Jinkela_wire_5154),
        .dout(new_Jinkela_wire_5155)
    );

    spl2 new_Jinkela_splitter_482 (
        .a(_1387_),
        .b(new_Jinkela_wire_5161),
        .c(new_Jinkela_wire_5162)
    );

    bfr new_Jinkela_buffer_3892 (
        .din(new_Jinkela_wire_5155),
        .dout(new_Jinkela_wire_5156)
    );

    bfr new_Jinkela_buffer_3900 (
        .din(_0926_),
        .dout(new_Jinkela_wire_5168)
    );

    spl2 new_Jinkela_splitter_484 (
        .a(_0258_),
        .b(new_Jinkela_wire_5282),
        .c(new_Jinkela_wire_5283)
    );

    bfr new_Jinkela_buffer_3896 (
        .din(new_Jinkela_wire_5163),
        .dout(new_Jinkela_wire_5164)
    );

    spl2 new_Jinkela_splitter_485 (
        .a(_0367_),
        .b(new_Jinkela_wire_5284),
        .c(new_Jinkela_wire_5285)
    );

    bfr new_Jinkela_buffer_3897 (
        .din(new_Jinkela_wire_5164),
        .dout(new_Jinkela_wire_5165)
    );

    bfr new_Jinkela_buffer_3901 (
        .din(new_Jinkela_wire_5168),
        .dout(new_Jinkela_wire_5169)
    );

    bfr new_Jinkela_buffer_3898 (
        .din(new_Jinkela_wire_5165),
        .dout(new_Jinkela_wire_5166)
    );

    bfr new_Jinkela_buffer_3902 (
        .din(new_Jinkela_wire_5169),
        .dout(new_Jinkela_wire_5170)
    );

    spl2 new_Jinkela_splitter_488 (
        .a(_1648_),
        .b(new_Jinkela_wire_5418),
        .c(new_Jinkela_wire_5419)
    );

    bfr new_Jinkela_buffer_4012 (
        .din(_1074_),
        .dout(new_Jinkela_wire_5286)
    );

    bfr new_Jinkela_buffer_3903 (
        .din(new_Jinkela_wire_5170),
        .dout(new_Jinkela_wire_5171)
    );

    bfr new_Jinkela_buffer_4052 (
        .din(_0439_),
        .dout(new_Jinkela_wire_5328)
    );

    bfr new_Jinkela_buffer_3904 (
        .din(new_Jinkela_wire_5171),
        .dout(new_Jinkela_wire_5172)
    );

    bfr new_Jinkela_buffer_4013 (
        .din(new_Jinkela_wire_5286),
        .dout(new_Jinkela_wire_5287)
    );

    bfr new_Jinkela_buffer_3905 (
        .din(new_Jinkela_wire_5172),
        .dout(new_Jinkela_wire_5173)
    );

    bfr new_Jinkela_buffer_4140 (
        .din(_1064_),
        .dout(new_Jinkela_wire_5420)
    );

    bfr new_Jinkela_buffer_3906 (
        .din(new_Jinkela_wire_5173),
        .dout(new_Jinkela_wire_5174)
    );

    bfr new_Jinkela_buffer_4014 (
        .din(new_Jinkela_wire_5287),
        .dout(new_Jinkela_wire_5288)
    );

    bfr new_Jinkela_buffer_3907 (
        .din(new_Jinkela_wire_5174),
        .dout(new_Jinkela_wire_5175)
    );

    bfr new_Jinkela_buffer_4053 (
        .din(new_Jinkela_wire_5328),
        .dout(new_Jinkela_wire_5329)
    );

    bfr new_Jinkela_buffer_3908 (
        .din(new_Jinkela_wire_5175),
        .dout(new_Jinkela_wire_5176)
    );

    bfr new_Jinkela_buffer_4015 (
        .din(new_Jinkela_wire_5288),
        .dout(new_Jinkela_wire_5289)
    );

    bfr new_Jinkela_buffer_3909 (
        .din(new_Jinkela_wire_5176),
        .dout(new_Jinkela_wire_5177)
    );

    spl2 new_Jinkela_splitter_489 (
        .a(_1308_),
        .b(new_Jinkela_wire_5422),
        .c(new_Jinkela_wire_5423)
    );

    bfr new_Jinkela_buffer_3910 (
        .din(new_Jinkela_wire_5177),
        .dout(new_Jinkela_wire_5178)
    );

    bfr new_Jinkela_buffer_4016 (
        .din(new_Jinkela_wire_5289),
        .dout(new_Jinkela_wire_5290)
    );

    bfr new_Jinkela_buffer_3911 (
        .din(new_Jinkela_wire_5178),
        .dout(new_Jinkela_wire_5179)
    );

    bfr new_Jinkela_buffer_4054 (
        .din(new_Jinkela_wire_5329),
        .dout(new_Jinkela_wire_5330)
    );

    bfr new_Jinkela_buffer_3912 (
        .din(new_Jinkela_wire_5179),
        .dout(new_Jinkela_wire_5180)
    );

    bfr new_Jinkela_buffer_4017 (
        .din(new_Jinkela_wire_5290),
        .dout(new_Jinkela_wire_5291)
    );

    bfr new_Jinkela_buffer_3913 (
        .din(new_Jinkela_wire_5180),
        .dout(new_Jinkela_wire_5181)
    );

    bfr new_Jinkela_buffer_4141 (
        .din(_0825_),
        .dout(new_Jinkela_wire_5421)
    );

    bfr new_Jinkela_buffer_3914 (
        .din(new_Jinkela_wire_5181),
        .dout(new_Jinkela_wire_5182)
    );

    bfr new_Jinkela_buffer_4018 (
        .din(new_Jinkela_wire_5291),
        .dout(new_Jinkela_wire_5292)
    );

    bfr new_Jinkela_buffer_3915 (
        .din(new_Jinkela_wire_5182),
        .dout(new_Jinkela_wire_5183)
    );

    bfr new_Jinkela_buffer_7486 (
        .din(new_Jinkela_wire_9303),
        .dout(new_Jinkela_wire_9304)
    );

    bfr new_Jinkela_buffer_14265 (
        .din(new_Jinkela_wire_17034),
        .dout(new_Jinkela_wire_17035)
    );

    bfr new_Jinkela_buffer_17666 (
        .din(new_Jinkela_wire_21034),
        .dout(new_Jinkela_wire_21035)
    );

    bfr new_Jinkela_buffer_7297 (
        .din(new_Jinkela_wire_9088),
        .dout(new_Jinkela_wire_9089)
    );

    bfr new_Jinkela_buffer_17743 (
        .din(new_Jinkela_wire_21133),
        .dout(new_Jinkela_wire_21134)
    );

    bfr new_Jinkela_buffer_7335 (
        .din(new_Jinkela_wire_9136),
        .dout(new_Jinkela_wire_9137)
    );

    bfr new_Jinkela_buffer_14266 (
        .din(new_Jinkela_wire_17035),
        .dout(new_Jinkela_wire_17036)
    );

    bfr new_Jinkela_buffer_17667 (
        .din(new_Jinkela_wire_21035),
        .dout(new_Jinkela_wire_21036)
    );

    bfr new_Jinkela_buffer_7298 (
        .din(new_Jinkela_wire_9089),
        .dout(new_Jinkela_wire_9090)
    );

    bfr new_Jinkela_buffer_14268 (
        .din(new_Jinkela_wire_17039),
        .dout(new_Jinkela_wire_17040)
    );

    bfr new_Jinkela_buffer_17760 (
        .din(new_Jinkela_wire_21156),
        .dout(new_Jinkela_wire_21157)
    );

    bfr new_Jinkela_buffer_7382 (
        .din(new_Jinkela_wire_9197),
        .dout(new_Jinkela_wire_9198)
    );

    bfr new_Jinkela_buffer_17668 (
        .din(new_Jinkela_wire_21036),
        .dout(new_Jinkela_wire_21037)
    );

    spl2 new_Jinkela_splitter_1237 (
        .a(_0133_),
        .b(new_Jinkela_wire_17047),
        .c(new_Jinkela_wire_17048)
    );

    bfr new_Jinkela_buffer_7299 (
        .din(new_Jinkela_wire_9090),
        .dout(new_Jinkela_wire_9091)
    );

    bfr new_Jinkela_buffer_14269 (
        .din(new_Jinkela_wire_17040),
        .dout(new_Jinkela_wire_17041)
    );

    bfr new_Jinkela_buffer_17744 (
        .din(new_Jinkela_wire_21134),
        .dout(new_Jinkela_wire_21135)
    );

    bfr new_Jinkela_buffer_7336 (
        .din(new_Jinkela_wire_9137),
        .dout(new_Jinkela_wire_9138)
    );

    bfr new_Jinkela_buffer_17669 (
        .din(new_Jinkela_wire_21037),
        .dout(new_Jinkela_wire_21038)
    );

    spl2 new_Jinkela_splitter_1238 (
        .a(_1145_),
        .b(new_Jinkela_wire_17049),
        .c(new_Jinkela_wire_17050)
    );

    spl2 new_Jinkela_splitter_745 (
        .a(new_Jinkela_wire_9091),
        .b(new_Jinkela_wire_9092),
        .c(new_Jinkela_wire_9093)
    );

    bfr new_Jinkela_buffer_14270 (
        .din(new_Jinkela_wire_17041),
        .dout(new_Jinkela_wire_17042)
    );

    bfr new_Jinkela_buffer_17765 (
        .din(_0320_),
        .dout(new_Jinkela_wire_21168)
    );

    bfr new_Jinkela_buffer_7337 (
        .din(new_Jinkela_wire_9138),
        .dout(new_Jinkela_wire_9139)
    );

    bfr new_Jinkela_buffer_17670 (
        .din(new_Jinkela_wire_21038),
        .dout(new_Jinkela_wire_21039)
    );

    spl2 new_Jinkela_splitter_1239 (
        .a(_0504_),
        .b(new_Jinkela_wire_17051),
        .c(new_Jinkela_wire_17052)
    );

    bfr new_Jinkela_buffer_17745 (
        .din(new_Jinkela_wire_21135),
        .dout(new_Jinkela_wire_21136)
    );

    bfr new_Jinkela_buffer_7682 (
        .din(_1586_),
        .dout(new_Jinkela_wire_9510)
    );

    spl2 new_Jinkela_splitter_1240 (
        .a(_1563_),
        .b(new_Jinkela_wire_17053),
        .c(new_Jinkela_wire_17054)
    );

    bfr new_Jinkela_buffer_7383 (
        .din(new_Jinkela_wire_9198),
        .dout(new_Jinkela_wire_9199)
    );

    bfr new_Jinkela_buffer_14272 (
        .din(new_Jinkela_wire_17057),
        .dout(new_Jinkela_wire_17058)
    );

    bfr new_Jinkela_buffer_17671 (
        .din(new_Jinkela_wire_21039),
        .dout(new_Jinkela_wire_21040)
    );

    bfr new_Jinkela_buffer_14271 (
        .din(_0197_),
        .dout(new_Jinkela_wire_17055)
    );

    bfr new_Jinkela_buffer_7338 (
        .din(new_Jinkela_wire_9139),
        .dout(new_Jinkela_wire_9140)
    );

    bfr new_Jinkela_buffer_14276 (
        .din(_1391_),
        .dout(new_Jinkela_wire_17062)
    );

    bfr new_Jinkela_buffer_17761 (
        .din(new_Jinkela_wire_21157),
        .dout(new_Jinkela_wire_21158)
    );

    spl2 new_Jinkela_splitter_1241 (
        .a(_1725_),
        .b(new_Jinkela_wire_17056),
        .c(new_Jinkela_wire_17057)
    );

    bfr new_Jinkela_buffer_7487 (
        .din(new_Jinkela_wire_9304),
        .dout(new_Jinkela_wire_9305)
    );

    bfr new_Jinkela_buffer_17672 (
        .din(new_Jinkela_wire_21040),
        .dout(new_Jinkela_wire_21041)
    );

    bfr new_Jinkela_buffer_7339 (
        .din(new_Jinkela_wire_9140),
        .dout(new_Jinkela_wire_9141)
    );

    bfr new_Jinkela_buffer_17746 (
        .din(new_Jinkela_wire_21136),
        .dout(new_Jinkela_wire_21137)
    );

    spl2 new_Jinkela_splitter_1242 (
        .a(_1501_),
        .b(new_Jinkela_wire_17063),
        .c(new_Jinkela_wire_17064)
    );

    bfr new_Jinkela_buffer_7384 (
        .din(new_Jinkela_wire_9199),
        .dout(new_Jinkela_wire_9200)
    );

    spl2 new_Jinkela_splitter_1243 (
        .a(_0020_),
        .b(new_Jinkela_wire_17065),
        .c(new_Jinkela_wire_17066)
    );

    bfr new_Jinkela_buffer_17673 (
        .din(new_Jinkela_wire_21041),
        .dout(new_Jinkela_wire_21042)
    );

    and_bb _1886_ (
        .a(new_Jinkela_wire_9608),
        .b(new_Jinkela_wire_10450),
        .c(_0143_)
    );

    bfr new_Jinkela_buffer_7340 (
        .din(new_Jinkela_wire_9141),
        .dout(new_Jinkela_wire_9142)
    );

    bfr new_Jinkela_buffer_14273 (
        .din(new_Jinkela_wire_17058),
        .dout(new_Jinkela_wire_17059)
    );

    bfr new_Jinkela_buffer_17763 (
        .din(_1061_),
        .dout(new_Jinkela_wire_21166)
    );

    bfr new_Jinkela_buffer_7530 (
        .din(new_Jinkela_wire_9351),
        .dout(new_Jinkela_wire_9352)
    );

    bfr new_Jinkela_buffer_17674 (
        .din(new_Jinkela_wire_21042),
        .dout(new_Jinkela_wire_21043)
    );

    bfr new_Jinkela_buffer_7341 (
        .din(new_Jinkela_wire_9142),
        .dout(new_Jinkela_wire_9143)
    );

    bfr new_Jinkela_buffer_14274 (
        .din(new_Jinkela_wire_17059),
        .dout(new_Jinkela_wire_17060)
    );

    bfr new_Jinkela_buffer_17747 (
        .din(new_Jinkela_wire_21137),
        .dout(new_Jinkela_wire_21138)
    );

    bfr new_Jinkela_buffer_7385 (
        .din(new_Jinkela_wire_9200),
        .dout(new_Jinkela_wire_9201)
    );

    spl2 new_Jinkela_splitter_1244 (
        .a(_1085_),
        .b(new_Jinkela_wire_17067),
        .c(new_Jinkela_wire_17068)
    );

    bfr new_Jinkela_buffer_17675 (
        .din(new_Jinkela_wire_21043),
        .dout(new_Jinkela_wire_21044)
    );

    bfr new_Jinkela_buffer_7342 (
        .din(new_Jinkela_wire_9143),
        .dout(new_Jinkela_wire_9144)
    );

    bfr new_Jinkela_buffer_14275 (
        .din(new_Jinkela_wire_17060),
        .dout(new_Jinkela_wire_17061)
    );

    bfr new_Jinkela_buffer_17762 (
        .din(new_Jinkela_wire_21158),
        .dout(new_Jinkela_wire_21159)
    );

    bfr new_Jinkela_buffer_7488 (
        .din(new_Jinkela_wire_9305),
        .dout(new_Jinkela_wire_9306)
    );

    bfr new_Jinkela_buffer_17676 (
        .din(new_Jinkela_wire_21044),
        .dout(new_Jinkela_wire_21045)
    );

    spl2 new_Jinkela_splitter_1245 (
        .a(_0880_),
        .b(new_Jinkela_wire_17069),
        .c(new_Jinkela_wire_17070)
    );

    bfr new_Jinkela_buffer_7343 (
        .din(new_Jinkela_wire_9144),
        .dout(new_Jinkela_wire_9145)
    );

    bfr new_Jinkela_buffer_17748 (
        .din(new_Jinkela_wire_21138),
        .dout(new_Jinkela_wire_21139)
    );

    spl2 new_Jinkela_splitter_1246 (
        .a(_1699_),
        .b(new_Jinkela_wire_17071),
        .c(new_Jinkela_wire_17072)
    );

    bfr new_Jinkela_buffer_7386 (
        .din(new_Jinkela_wire_9201),
        .dout(new_Jinkela_wire_9202)
    );

    bfr new_Jinkela_buffer_17677 (
        .din(new_Jinkela_wire_21045),
        .dout(new_Jinkela_wire_21046)
    );

    spl2 new_Jinkela_splitter_1247 (
        .a(_0120_),
        .b(new_Jinkela_wire_17073),
        .c(new_Jinkela_wire_17074)
    );

    bfr new_Jinkela_buffer_7344 (
        .din(new_Jinkela_wire_9145),
        .dout(new_Jinkela_wire_9146)
    );

    spl2 new_Jinkela_splitter_1248 (
        .a(_1153_),
        .b(new_Jinkela_wire_17079),
        .c(new_Jinkela_wire_17080)
    );

    bfr new_Jinkela_buffer_17764 (
        .din(_1433_),
        .dout(new_Jinkela_wire_21167)
    );

    bfr new_Jinkela_buffer_7541 (
        .din(new_Jinkela_wire_9364),
        .dout(new_Jinkela_wire_9365)
    );

    bfr new_Jinkela_buffer_14277 (
        .din(new_Jinkela_wire_17074),
        .dout(new_Jinkela_wire_17075)
    );

    bfr new_Jinkela_buffer_17678 (
        .din(new_Jinkela_wire_21046),
        .dout(new_Jinkela_wire_21047)
    );

    spl2 new_Jinkela_splitter_1249 (
        .a(_0156_),
        .b(new_Jinkela_wire_17081),
        .c(new_Jinkela_wire_17082)
    );

    bfr new_Jinkela_buffer_7345 (
        .din(new_Jinkela_wire_9146),
        .dout(new_Jinkela_wire_9147)
    );

    bfr new_Jinkela_buffer_17749 (
        .din(new_Jinkela_wire_21139),
        .dout(new_Jinkela_wire_21140)
    );

    bfr new_Jinkela_buffer_7387 (
        .din(new_Jinkela_wire_9202),
        .dout(new_Jinkela_wire_9203)
    );

    bfr new_Jinkela_buffer_14278 (
        .din(new_Jinkela_wire_17075),
        .dout(new_Jinkela_wire_17076)
    );

    bfr new_Jinkela_buffer_17679 (
        .din(new_Jinkela_wire_21047),
        .dout(new_Jinkela_wire_21048)
    );

    bfr new_Jinkela_buffer_7346 (
        .din(new_Jinkela_wire_9147),
        .dout(new_Jinkela_wire_9148)
    );

    spl2 new_Jinkela_splitter_1547 (
        .a(new_Jinkela_wire_21159),
        .b(new_Jinkela_wire_21160),
        .c(new_Jinkela_wire_21161)
    );

    spl2 new_Jinkela_splitter_1250 (
        .a(_1358_),
        .b(new_Jinkela_wire_17083),
        .c(new_Jinkela_wire_17084)
    );

    bfr new_Jinkela_buffer_7489 (
        .din(new_Jinkela_wire_9306),
        .dout(new_Jinkela_wire_9307)
    );

    bfr new_Jinkela_buffer_14279 (
        .din(new_Jinkela_wire_17076),
        .dout(new_Jinkela_wire_17077)
    );

    bfr new_Jinkela_buffer_17680 (
        .din(new_Jinkela_wire_21048),
        .dout(new_Jinkela_wire_21049)
    );

    bfr new_Jinkela_buffer_7347 (
        .din(new_Jinkela_wire_9148),
        .dout(new_Jinkela_wire_9149)
    );

    bfr new_Jinkela_buffer_17750 (
        .din(new_Jinkela_wire_21140),
        .dout(new_Jinkela_wire_21141)
    );

    spl2 new_Jinkela_splitter_1251 (
        .a(_1581_),
        .b(new_Jinkela_wire_17085),
        .c(new_Jinkela_wire_17086)
    );

    bfr new_Jinkela_buffer_7388 (
        .din(new_Jinkela_wire_9203),
        .dout(new_Jinkela_wire_9204)
    );

    bfr new_Jinkela_buffer_14280 (
        .din(new_Jinkela_wire_17077),
        .dout(new_Jinkela_wire_17078)
    );

    bfr new_Jinkela_buffer_17681 (
        .din(new_Jinkela_wire_21049),
        .dout(new_Jinkela_wire_21050)
    );

    bfr new_Jinkela_buffer_7348 (
        .din(new_Jinkela_wire_9149),
        .dout(new_Jinkela_wire_9150)
    );

    spl2 new_Jinkela_splitter_1551 (
        .a(_0840_),
        .b(new_Jinkela_wire_21175),
        .c(new_Jinkela_wire_21176)
    );

    spl2 new_Jinkela_splitter_1252 (
        .a(_1477_),
        .b(new_Jinkela_wire_17087),
        .c(new_Jinkela_wire_17088)
    );

    bfr new_Jinkela_buffer_7531 (
        .din(new_Jinkela_wire_9352),
        .dout(new_Jinkela_wire_9353)
    );

    bfr new_Jinkela_buffer_17682 (
        .din(new_Jinkela_wire_21050),
        .dout(new_Jinkela_wire_21051)
    );

    bfr new_Jinkela_buffer_14281 (
        .din(_0968_),
        .dout(new_Jinkela_wire_17089)
    );

    bfr new_Jinkela_buffer_7349 (
        .din(new_Jinkela_wire_9150),
        .dout(new_Jinkela_wire_9151)
    );

    spl3L new_Jinkela_splitter_1254 (
        .a(_1587_),
        .d(new_Jinkela_wire_17108),
        .b(new_Jinkela_wire_17109),
        .c(new_Jinkela_wire_17110)
    );

    bfr new_Jinkela_buffer_17751 (
        .din(new_Jinkela_wire_21141),
        .dout(new_Jinkela_wire_21142)
    );

    bfr new_Jinkela_buffer_14282 (
        .din(_1294_),
        .dout(new_Jinkela_wire_17090)
    );

    bfr new_Jinkela_buffer_7389 (
        .din(new_Jinkela_wire_9204),
        .dout(new_Jinkela_wire_9205)
    );

    bfr new_Jinkela_buffer_17683 (
        .din(new_Jinkela_wire_21051),
        .dout(new_Jinkela_wire_21052)
    );

    spl2 new_Jinkela_splitter_1255 (
        .a(_0980_),
        .b(new_Jinkela_wire_17111),
        .c(new_Jinkela_wire_17112)
    );

    bfr new_Jinkela_buffer_7350 (
        .din(new_Jinkela_wire_9151),
        .dout(new_Jinkela_wire_9152)
    );

    bfr new_Jinkela_buffer_14283 (
        .din(new_Jinkela_wire_17090),
        .dout(new_Jinkela_wire_17091)
    );

    bfr new_Jinkela_buffer_17766 (
        .din(_0357_),
        .dout(new_Jinkela_wire_21169)
    );

    bfr new_Jinkela_buffer_7490 (
        .din(new_Jinkela_wire_9307),
        .dout(new_Jinkela_wire_9308)
    );

    bfr new_Jinkela_buffer_14346 (
        .din(new_net_3968),
        .dout(new_Jinkela_wire_17161)
    );

    bfr new_Jinkela_buffer_17684 (
        .din(new_Jinkela_wire_21052),
        .dout(new_Jinkela_wire_21053)
    );

    bfr new_Jinkela_buffer_7351 (
        .din(new_Jinkela_wire_9152),
        .dout(new_Jinkela_wire_9153)
    );

    bfr new_Jinkela_buffer_14284 (
        .din(new_Jinkela_wire_17091),
        .dout(new_Jinkela_wire_17092)
    );

    bfr new_Jinkela_buffer_17752 (
        .din(new_Jinkela_wire_21142),
        .dout(new_Jinkela_wire_21143)
    );

    bfr new_Jinkela_buffer_7390 (
        .din(new_Jinkela_wire_9205),
        .dout(new_Jinkela_wire_9206)
    );

    bfr new_Jinkela_buffer_17685 (
        .din(new_Jinkela_wire_21053),
        .dout(new_Jinkela_wire_21054)
    );

    spl2 new_Jinkela_splitter_1256 (
        .a(_0462_),
        .b(new_Jinkela_wire_17317),
        .c(new_Jinkela_wire_17318)
    );

    bfr new_Jinkela_buffer_7352 (
        .din(new_Jinkela_wire_9153),
        .dout(new_Jinkela_wire_9154)
    );

    bfr new_Jinkela_buffer_14285 (
        .din(new_Jinkela_wire_17092),
        .dout(new_Jinkela_wire_17093)
    );

    spl2 new_Jinkela_splitter_1552 (
        .a(_0001_),
        .b(new_Jinkela_wire_21177),
        .c(new_Jinkela_wire_21178)
    );

    bfr new_Jinkela_buffer_7620 (
        .din(new_Jinkela_wire_9447),
        .dout(new_Jinkela_wire_9448)
    );

    bfr new_Jinkela_buffer_14298 (
        .din(new_Jinkela_wire_17112),
        .dout(new_Jinkela_wire_17113)
    );

    bfr new_Jinkela_buffer_17686 (
        .din(new_Jinkela_wire_21054),
        .dout(new_Jinkela_wire_21055)
    );

    bfr new_Jinkela_buffer_7353 (
        .din(new_Jinkela_wire_9154),
        .dout(new_Jinkela_wire_9155)
    );

    bfr new_Jinkela_buffer_14286 (
        .din(new_Jinkela_wire_17093),
        .dout(new_Jinkela_wire_17094)
    );

    bfr new_Jinkela_buffer_17753 (
        .din(new_Jinkela_wire_21143),
        .dout(new_Jinkela_wire_21144)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_953),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_1050),
        .dout(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_955),
        .dout(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_1145),
        .dout(new_Jinkela_wire_1146)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_1093),
        .dout(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_1051),
        .dout(new_Jinkela_wire_1052)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_957),
        .dout(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_1052),
        .dout(new_Jinkela_wire_1053)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_960),
        .dout(new_Jinkela_wire_961)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_1053),
        .dout(new_Jinkela_wire_1054)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_961),
        .dout(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(_0147_),
        .b(new_Jinkela_wire_1269),
        .c(new_Jinkela_wire_1270)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_1054),
        .dout(new_Jinkela_wire_1055)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_1146),
        .dout(new_Jinkela_wire_1147)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_1095),
        .dout(new_Jinkela_wire_1096)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_1055),
        .dout(new_Jinkela_wire_1056)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_1056),
        .dout(new_Jinkela_wire_1057)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    spl2 new_Jinkela_splitter_211 (
        .a(_0219_),
        .b(new_Jinkela_wire_1275),
        .c(new_Jinkela_wire_1276)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_1057),
        .dout(new_Jinkela_wire_1058)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_969),
        .dout(new_Jinkela_wire_970)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_1058),
        .dout(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_1147),
        .dout(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_972),
        .dout(new_Jinkela_wire_973)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_1097),
        .dout(new_Jinkela_wire_1098)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_1059),
        .dout(new_Jinkela_wire_1060)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_14506 (
        .din(_1700_),
        .dout(new_Jinkela_wire_17323)
    );

    bfr new_Jinkela_buffer_17687 (
        .din(new_Jinkela_wire_21055),
        .dout(new_Jinkela_wire_21056)
    );

    bfr new_Jinkela_buffer_14347 (
        .din(new_Jinkela_wire_17161),
        .dout(new_Jinkela_wire_17162)
    );

    bfr new_Jinkela_buffer_14287 (
        .din(new_Jinkela_wire_17094),
        .dout(new_Jinkela_wire_17095)
    );

    bfr new_Jinkela_buffer_17767 (
        .din(new_Jinkela_wire_21169),
        .dout(new_Jinkela_wire_21170)
    );

    bfr new_Jinkela_buffer_14299 (
        .din(new_Jinkela_wire_17113),
        .dout(new_Jinkela_wire_17114)
    );

    bfr new_Jinkela_buffer_17688 (
        .din(new_Jinkela_wire_21056),
        .dout(new_Jinkela_wire_21057)
    );

    bfr new_Jinkela_buffer_14288 (
        .din(new_Jinkela_wire_17095),
        .dout(new_Jinkela_wire_17096)
    );

    bfr new_Jinkela_buffer_17754 (
        .din(new_Jinkela_wire_21144),
        .dout(new_Jinkela_wire_21145)
    );

    bfr new_Jinkela_buffer_17689 (
        .din(new_Jinkela_wire_21057),
        .dout(new_Jinkela_wire_21058)
    );

    bfr new_Jinkela_buffer_14502 (
        .din(new_Jinkela_wire_17318),
        .dout(new_Jinkela_wire_17319)
    );

    bfr new_Jinkela_buffer_14289 (
        .din(new_Jinkela_wire_17096),
        .dout(new_Jinkela_wire_17097)
    );

    spl2 new_Jinkela_splitter_1553 (
        .a(_0336_),
        .b(new_Jinkela_wire_21181),
        .c(new_Jinkela_wire_21182)
    );

    bfr new_Jinkela_buffer_14300 (
        .din(new_Jinkela_wire_17114),
        .dout(new_Jinkela_wire_17115)
    );

    bfr new_Jinkela_buffer_17690 (
        .din(new_Jinkela_wire_21058),
        .dout(new_Jinkela_wire_21059)
    );

    bfr new_Jinkela_buffer_14290 (
        .din(new_Jinkela_wire_17097),
        .dout(new_Jinkela_wire_17098)
    );

    bfr new_Jinkela_buffer_17768 (
        .din(new_Jinkela_wire_21170),
        .dout(new_Jinkela_wire_21171)
    );

    bfr new_Jinkela_buffer_17691 (
        .din(new_Jinkela_wire_21059),
        .dout(new_Jinkela_wire_21060)
    );

    bfr new_Jinkela_buffer_14348 (
        .din(new_Jinkela_wire_17162),
        .dout(new_Jinkela_wire_17163)
    );

    bfr new_Jinkela_buffer_14291 (
        .din(new_Jinkela_wire_17098),
        .dout(new_Jinkela_wire_17099)
    );

    bfr new_Jinkela_buffer_17770 (
        .din(_0673_),
        .dout(new_Jinkela_wire_21179)
    );

    bfr new_Jinkela_buffer_14301 (
        .din(new_Jinkela_wire_17115),
        .dout(new_Jinkela_wire_17116)
    );

    bfr new_Jinkela_buffer_17692 (
        .din(new_Jinkela_wire_21060),
        .dout(new_Jinkela_wire_21061)
    );

    bfr new_Jinkela_buffer_14292 (
        .din(new_Jinkela_wire_17099),
        .dout(new_Jinkela_wire_17100)
    );

    bfr new_Jinkela_buffer_17769 (
        .din(new_Jinkela_wire_21171),
        .dout(new_Jinkela_wire_21172)
    );

    bfr new_Jinkela_buffer_17693 (
        .din(new_Jinkela_wire_21061),
        .dout(new_Jinkela_wire_21062)
    );

    bfr new_Jinkela_buffer_14293 (
        .din(new_Jinkela_wire_17100),
        .dout(new_Jinkela_wire_17101)
    );

    bfr new_Jinkela_buffer_17771 (
        .din(_0496_),
        .dout(new_Jinkela_wire_21180)
    );

    bfr new_Jinkela_buffer_14302 (
        .din(new_Jinkela_wire_17116),
        .dout(new_Jinkela_wire_17117)
    );

    bfr new_Jinkela_buffer_17694 (
        .din(new_Jinkela_wire_21062),
        .dout(new_Jinkela_wire_21063)
    );

    bfr new_Jinkela_buffer_14294 (
        .din(new_Jinkela_wire_17101),
        .dout(new_Jinkela_wire_17102)
    );

    spl2 new_Jinkela_splitter_1550 (
        .a(new_Jinkela_wire_21172),
        .b(new_Jinkela_wire_21173),
        .c(new_Jinkela_wire_21174)
    );

    bfr new_Jinkela_buffer_17695 (
        .din(new_Jinkela_wire_21063),
        .dout(new_Jinkela_wire_21064)
    );

    bfr new_Jinkela_buffer_14349 (
        .din(new_Jinkela_wire_17163),
        .dout(new_Jinkela_wire_17164)
    );

    bfr new_Jinkela_buffer_14295 (
        .din(new_Jinkela_wire_17102),
        .dout(new_Jinkela_wire_17103)
    );

    bfr new_Jinkela_buffer_17773 (
        .din(new_Jinkela_wire_21185),
        .dout(new_Jinkela_wire_21186)
    );

    bfr new_Jinkela_buffer_14303 (
        .din(new_Jinkela_wire_17117),
        .dout(new_Jinkela_wire_17118)
    );

    bfr new_Jinkela_buffer_17696 (
        .din(new_Jinkela_wire_21064),
        .dout(new_Jinkela_wire_21065)
    );

    bfr new_Jinkela_buffer_14296 (
        .din(new_Jinkela_wire_17103),
        .dout(new_Jinkela_wire_17104)
    );

    bfr new_Jinkela_buffer_17772 (
        .din(_0916_),
        .dout(new_Jinkela_wire_21183)
    );

    spl2 new_Jinkela_splitter_1555 (
        .a(_0970_),
        .b(new_Jinkela_wire_21190),
        .c(new_Jinkela_wire_21191)
    );

    bfr new_Jinkela_buffer_17697 (
        .din(new_Jinkela_wire_21065),
        .dout(new_Jinkela_wire_21066)
    );

    spl2 new_Jinkela_splitter_1258 (
        .a(_0347_),
        .b(new_Jinkela_wire_17357),
        .c(new_Jinkela_wire_17358)
    );

    bfr new_Jinkela_buffer_14297 (
        .din(new_Jinkela_wire_17104),
        .dout(new_Jinkela_wire_17105)
    );

    spl2 new_Jinkela_splitter_1554 (
        .a(_0796_),
        .b(new_Jinkela_wire_21184),
        .c(new_Jinkela_wire_21185)
    );

    bfr new_Jinkela_buffer_14304 (
        .din(new_Jinkela_wire_17118),
        .dout(new_Jinkela_wire_17119)
    );

    bfr new_Jinkela_buffer_17698 (
        .din(new_Jinkela_wire_21066),
        .dout(new_Jinkela_wire_21067)
    );

    spl2 new_Jinkela_splitter_1253 (
        .a(new_Jinkela_wire_17105),
        .b(new_Jinkela_wire_17106),
        .c(new_Jinkela_wire_17107)
    );

    bfr new_Jinkela_buffer_14305 (
        .din(new_Jinkela_wire_17119),
        .dout(new_Jinkela_wire_17120)
    );

    bfr new_Jinkela_buffer_17699 (
        .din(new_Jinkela_wire_21067),
        .dout(new_Jinkela_wire_21068)
    );

    bfr new_Jinkela_buffer_14350 (
        .din(new_Jinkela_wire_17164),
        .dout(new_Jinkela_wire_17165)
    );

    spl2 new_Jinkela_splitter_1556 (
        .a(_1631_),
        .b(new_Jinkela_wire_21192),
        .c(new_Jinkela_wire_21193)
    );

    bfr new_Jinkela_buffer_17700 (
        .din(new_Jinkela_wire_21068),
        .dout(new_Jinkela_wire_21069)
    );

    spl2 new_Jinkela_splitter_1259 (
        .a(_1669_),
        .b(new_Jinkela_wire_17359),
        .c(new_Jinkela_wire_17360)
    );

    bfr new_Jinkela_buffer_14306 (
        .din(new_Jinkela_wire_17120),
        .dout(new_Jinkela_wire_17121)
    );

    bfr new_Jinkela_buffer_14503 (
        .din(new_Jinkela_wire_17319),
        .dout(new_Jinkela_wire_17320)
    );

    bfr new_Jinkela_buffer_17701 (
        .din(new_Jinkela_wire_21069),
        .dout(new_Jinkela_wire_21070)
    );

    bfr new_Jinkela_buffer_14351 (
        .din(new_Jinkela_wire_17165),
        .dout(new_Jinkela_wire_17166)
    );

    bfr new_Jinkela_buffer_14307 (
        .din(new_Jinkela_wire_17121),
        .dout(new_Jinkela_wire_17122)
    );

    bfr new_Jinkela_buffer_17774 (
        .din(new_Jinkela_wire_21186),
        .dout(new_Jinkela_wire_21187)
    );

    bfr new_Jinkela_buffer_17702 (
        .din(new_Jinkela_wire_21070),
        .dout(new_Jinkela_wire_21071)
    );

    bfr new_Jinkela_buffer_14308 (
        .din(new_Jinkela_wire_17122),
        .dout(new_Jinkela_wire_17123)
    );

    bfr new_Jinkela_buffer_17777 (
        .din(_1265_),
        .dout(new_Jinkela_wire_21194)
    );

    bfr new_Jinkela_buffer_14507 (
        .din(new_Jinkela_wire_17323),
        .dout(new_Jinkela_wire_17324)
    );

    bfr new_Jinkela_buffer_17703 (
        .din(new_Jinkela_wire_21071),
        .dout(new_Jinkela_wire_21072)
    );

    bfr new_Jinkela_buffer_14352 (
        .din(new_Jinkela_wire_17166),
        .dout(new_Jinkela_wire_17167)
    );

    bfr new_Jinkela_buffer_14309 (
        .din(new_Jinkela_wire_17123),
        .dout(new_Jinkela_wire_17124)
    );

    bfr new_Jinkela_buffer_17775 (
        .din(new_Jinkela_wire_21187),
        .dout(new_Jinkela_wire_21188)
    );

    bfr new_Jinkela_buffer_17704 (
        .din(new_Jinkela_wire_21072),
        .dout(new_Jinkela_wire_21073)
    );

    bfr new_Jinkela_buffer_14310 (
        .din(new_Jinkela_wire_17124),
        .dout(new_Jinkela_wire_17125)
    );

    bfr new_Jinkela_buffer_17778 (
        .din(_1198_),
        .dout(new_Jinkela_wire_21197)
    );

    spl2 new_Jinkela_splitter_1557 (
        .a(_1505_),
        .b(new_Jinkela_wire_21195),
        .c(new_Jinkela_wire_21196)
    );

    bfr new_Jinkela_buffer_14504 (
        .din(new_Jinkela_wire_17320),
        .dout(new_Jinkela_wire_17321)
    );

    bfr new_Jinkela_buffer_17705 (
        .din(new_Jinkela_wire_21073),
        .dout(new_Jinkela_wire_21074)
    );

    bfr new_Jinkela_buffer_14353 (
        .din(new_Jinkela_wire_17167),
        .dout(new_Jinkela_wire_17168)
    );

    bfr new_Jinkela_buffer_14311 (
        .din(new_Jinkela_wire_17125),
        .dout(new_Jinkela_wire_17126)
    );

    bfr new_Jinkela_buffer_17776 (
        .din(new_Jinkela_wire_21188),
        .dout(new_Jinkela_wire_21189)
    );

    bfr new_Jinkela_buffer_17706 (
        .din(new_Jinkela_wire_21074),
        .dout(new_Jinkela_wire_21075)
    );

    bfr new_Jinkela_buffer_14312 (
        .din(new_Jinkela_wire_17126),
        .dout(new_Jinkela_wire_17127)
    );

    bfr new_Jinkela_buffer_17780 (
        .din(_1484_),
        .dout(new_Jinkela_wire_21199)
    );

    bfr new_Jinkela_buffer_17707 (
        .din(new_Jinkela_wire_21075),
        .dout(new_Jinkela_wire_21076)
    );

    bfr new_Jinkela_buffer_14354 (
        .din(new_Jinkela_wire_17168),
        .dout(new_Jinkela_wire_17169)
    );

    bfr new_Jinkela_buffer_14313 (
        .din(new_Jinkela_wire_17127),
        .dout(new_Jinkela_wire_17128)
    );

    bfr new_Jinkela_buffer_17779 (
        .din(_1300_),
        .dout(new_Jinkela_wire_21198)
    );

    bfr new_Jinkela_buffer_7391 (
        .din(new_Jinkela_wire_9206),
        .dout(new_Jinkela_wire_9207)
    );

    bfr new_Jinkela_buffer_4055 (
        .din(new_Jinkela_wire_5330),
        .dout(new_Jinkela_wire_5331)
    );

    bfr new_Jinkela_buffer_7354 (
        .din(new_Jinkela_wire_9155),
        .dout(new_Jinkela_wire_9156)
    );

    bfr new_Jinkela_buffer_3916 (
        .din(new_Jinkela_wire_5183),
        .dout(new_Jinkela_wire_5184)
    );

    bfr new_Jinkela_buffer_7491 (
        .din(new_Jinkela_wire_9308),
        .dout(new_Jinkela_wire_9309)
    );

    bfr new_Jinkela_buffer_4019 (
        .din(new_Jinkela_wire_5292),
        .dout(new_Jinkela_wire_5293)
    );

    bfr new_Jinkela_buffer_7355 (
        .din(new_Jinkela_wire_9156),
        .dout(new_Jinkela_wire_9157)
    );

    bfr new_Jinkela_buffer_3917 (
        .din(new_Jinkela_wire_5184),
        .dout(new_Jinkela_wire_5185)
    );

    bfr new_Jinkela_buffer_7392 (
        .din(new_Jinkela_wire_9207),
        .dout(new_Jinkela_wire_9208)
    );

    spl2 new_Jinkela_splitter_490 (
        .a(_1469_),
        .b(new_Jinkela_wire_5428),
        .c(new_Jinkela_wire_5429)
    );

    bfr new_Jinkela_buffer_4142 (
        .din(new_Jinkela_wire_5423),
        .dout(new_Jinkela_wire_5424)
    );

    bfr new_Jinkela_buffer_7356 (
        .din(new_Jinkela_wire_9157),
        .dout(new_Jinkela_wire_9158)
    );

    bfr new_Jinkela_buffer_3918 (
        .din(new_Jinkela_wire_5185),
        .dout(new_Jinkela_wire_5186)
    );

    bfr new_Jinkela_buffer_7532 (
        .din(new_Jinkela_wire_9353),
        .dout(new_Jinkela_wire_9354)
    );

    bfr new_Jinkela_buffer_4020 (
        .din(new_Jinkela_wire_5293),
        .dout(new_Jinkela_wire_5294)
    );

    bfr new_Jinkela_buffer_7357 (
        .din(new_Jinkela_wire_9158),
        .dout(new_Jinkela_wire_9159)
    );

    bfr new_Jinkela_buffer_3919 (
        .din(new_Jinkela_wire_5186),
        .dout(new_Jinkela_wire_5187)
    );

    bfr new_Jinkela_buffer_7393 (
        .din(new_Jinkela_wire_9208),
        .dout(new_Jinkela_wire_9209)
    );

    bfr new_Jinkela_buffer_4056 (
        .din(new_Jinkela_wire_5331),
        .dout(new_Jinkela_wire_5332)
    );

    bfr new_Jinkela_buffer_7358 (
        .din(new_Jinkela_wire_9159),
        .dout(new_Jinkela_wire_9160)
    );

    bfr new_Jinkela_buffer_3920 (
        .din(new_Jinkela_wire_5187),
        .dout(new_Jinkela_wire_5188)
    );

    bfr new_Jinkela_buffer_7492 (
        .din(new_Jinkela_wire_9309),
        .dout(new_Jinkela_wire_9310)
    );

    bfr new_Jinkela_buffer_4021 (
        .din(new_Jinkela_wire_5294),
        .dout(new_Jinkela_wire_5295)
    );

    bfr new_Jinkela_buffer_7359 (
        .din(new_Jinkela_wire_9160),
        .dout(new_Jinkela_wire_9161)
    );

    bfr new_Jinkela_buffer_3921 (
        .din(new_Jinkela_wire_5188),
        .dout(new_Jinkela_wire_5189)
    );

    bfr new_Jinkela_buffer_7394 (
        .din(new_Jinkela_wire_9209),
        .dout(new_Jinkela_wire_9210)
    );

    bfr new_Jinkela_buffer_7360 (
        .din(new_Jinkela_wire_9161),
        .dout(new_Jinkela_wire_9162)
    );

    bfr new_Jinkela_buffer_3922 (
        .din(new_Jinkela_wire_5189),
        .dout(new_Jinkela_wire_5190)
    );

    bfr new_Jinkela_buffer_7542 (
        .din(new_Jinkela_wire_9365),
        .dout(new_Jinkela_wire_9366)
    );

    bfr new_Jinkela_buffer_4022 (
        .din(new_Jinkela_wire_5295),
        .dout(new_Jinkela_wire_5296)
    );

    bfr new_Jinkela_buffer_7361 (
        .din(new_Jinkela_wire_9162),
        .dout(new_Jinkela_wire_9163)
    );

    bfr new_Jinkela_buffer_3923 (
        .din(new_Jinkela_wire_5190),
        .dout(new_Jinkela_wire_5191)
    );

    bfr new_Jinkela_buffer_7395 (
        .din(new_Jinkela_wire_9210),
        .dout(new_Jinkela_wire_9211)
    );

    bfr new_Jinkela_buffer_4057 (
        .din(new_Jinkela_wire_5332),
        .dout(new_Jinkela_wire_5333)
    );

    bfr new_Jinkela_buffer_7362 (
        .din(new_Jinkela_wire_9163),
        .dout(new_Jinkela_wire_9164)
    );

    bfr new_Jinkela_buffer_3924 (
        .din(new_Jinkela_wire_5191),
        .dout(new_Jinkela_wire_5192)
    );

    bfr new_Jinkela_buffer_7493 (
        .din(new_Jinkela_wire_9310),
        .dout(new_Jinkela_wire_9311)
    );

    bfr new_Jinkela_buffer_4023 (
        .din(new_Jinkela_wire_5296),
        .dout(new_Jinkela_wire_5297)
    );

    bfr new_Jinkela_buffer_7363 (
        .din(new_Jinkela_wire_9164),
        .dout(new_Jinkela_wire_9165)
    );

    bfr new_Jinkela_buffer_3925 (
        .din(new_Jinkela_wire_5192),
        .dout(new_Jinkela_wire_5193)
    );

    bfr new_Jinkela_buffer_7396 (
        .din(new_Jinkela_wire_9211),
        .dout(new_Jinkela_wire_9212)
    );

    spl2 new_Jinkela_splitter_491 (
        .a(_0738_),
        .b(new_Jinkela_wire_5430),
        .c(new_Jinkela_wire_5431)
    );

    bfr new_Jinkela_buffer_7364 (
        .din(new_Jinkela_wire_9165),
        .dout(new_Jinkela_wire_9166)
    );

    bfr new_Jinkela_buffer_3926 (
        .din(new_Jinkela_wire_5193),
        .dout(new_Jinkela_wire_5194)
    );

    bfr new_Jinkela_buffer_7533 (
        .din(new_Jinkela_wire_9354),
        .dout(new_Jinkela_wire_9355)
    );

    bfr new_Jinkela_buffer_4024 (
        .din(new_Jinkela_wire_5297),
        .dout(new_Jinkela_wire_5298)
    );

    bfr new_Jinkela_buffer_7365 (
        .din(new_Jinkela_wire_9166),
        .dout(new_Jinkela_wire_9167)
    );

    bfr new_Jinkela_buffer_3927 (
        .din(new_Jinkela_wire_5194),
        .dout(new_Jinkela_wire_5195)
    );

    bfr new_Jinkela_buffer_7397 (
        .din(new_Jinkela_wire_9212),
        .dout(new_Jinkela_wire_9213)
    );

    bfr new_Jinkela_buffer_4058 (
        .din(new_Jinkela_wire_5333),
        .dout(new_Jinkela_wire_5334)
    );

    bfr new_Jinkela_buffer_7366 (
        .din(new_Jinkela_wire_9167),
        .dout(new_Jinkela_wire_9168)
    );

    bfr new_Jinkela_buffer_3928 (
        .din(new_Jinkela_wire_5195),
        .dout(new_Jinkela_wire_5196)
    );

    bfr new_Jinkela_buffer_7494 (
        .din(new_Jinkela_wire_9311),
        .dout(new_Jinkela_wire_9312)
    );

    bfr new_Jinkela_buffer_4025 (
        .din(new_Jinkela_wire_5298),
        .dout(new_Jinkela_wire_5299)
    );

    bfr new_Jinkela_buffer_7367 (
        .din(new_Jinkela_wire_9168),
        .dout(new_Jinkela_wire_9169)
    );

    bfr new_Jinkela_buffer_3929 (
        .din(new_Jinkela_wire_5196),
        .dout(new_Jinkela_wire_5197)
    );

    bfr new_Jinkela_buffer_7398 (
        .din(new_Jinkela_wire_9213),
        .dout(new_Jinkela_wire_9214)
    );

    spl2 new_Jinkela_splitter_492 (
        .a(_1083_),
        .b(new_Jinkela_wire_5432),
        .c(new_Jinkela_wire_5433)
    );

    bfr new_Jinkela_buffer_7368 (
        .din(new_Jinkela_wire_9169),
        .dout(new_Jinkela_wire_9170)
    );

    bfr new_Jinkela_buffer_3930 (
        .din(new_Jinkela_wire_5197),
        .dout(new_Jinkela_wire_5198)
    );

    bfr new_Jinkela_buffer_4026 (
        .din(new_Jinkela_wire_5299),
        .dout(new_Jinkela_wire_5300)
    );

    bfr new_Jinkela_buffer_7690 (
        .din(_1739_),
        .dout(new_Jinkela_wire_9520)
    );

    spl2 new_Jinkela_splitter_750 (
        .a(new_Jinkela_wire_9170),
        .b(new_Jinkela_wire_9171),
        .c(new_Jinkela_wire_9172)
    );

    bfr new_Jinkela_buffer_3931 (
        .din(new_Jinkela_wire_5198),
        .dout(new_Jinkela_wire_5199)
    );

    bfr new_Jinkela_buffer_7495 (
        .din(new_Jinkela_wire_9312),
        .dout(new_Jinkela_wire_9313)
    );

    bfr new_Jinkela_buffer_4059 (
        .din(new_Jinkela_wire_5334),
        .dout(new_Jinkela_wire_5335)
    );

    bfr new_Jinkela_buffer_7399 (
        .din(new_Jinkela_wire_9214),
        .dout(new_Jinkela_wire_9215)
    );

    bfr new_Jinkela_buffer_3932 (
        .din(new_Jinkela_wire_5199),
        .dout(new_Jinkela_wire_5200)
    );

    bfr new_Jinkela_buffer_7400 (
        .din(new_Jinkela_wire_9215),
        .dout(new_Jinkela_wire_9216)
    );

    bfr new_Jinkela_buffer_4027 (
        .din(new_Jinkela_wire_5300),
        .dout(new_Jinkela_wire_5301)
    );

    bfr new_Jinkela_buffer_7534 (
        .din(new_Jinkela_wire_9355),
        .dout(new_Jinkela_wire_9356)
    );

    bfr new_Jinkela_buffer_3933 (
        .din(new_Jinkela_wire_5200),
        .dout(new_Jinkela_wire_5201)
    );

    bfr new_Jinkela_buffer_7401 (
        .din(new_Jinkela_wire_9216),
        .dout(new_Jinkela_wire_9217)
    );

    bfr new_Jinkela_buffer_4143 (
        .din(new_Jinkela_wire_5424),
        .dout(new_Jinkela_wire_5425)
    );

    bfr new_Jinkela_buffer_7496 (
        .din(new_Jinkela_wire_9313),
        .dout(new_Jinkela_wire_9314)
    );

    bfr new_Jinkela_buffer_3934 (
        .din(new_Jinkela_wire_5201),
        .dout(new_Jinkela_wire_5202)
    );

    bfr new_Jinkela_buffer_7402 (
        .din(new_Jinkela_wire_9217),
        .dout(new_Jinkela_wire_9218)
    );

    bfr new_Jinkela_buffer_4028 (
        .din(new_Jinkela_wire_5301),
        .dout(new_Jinkela_wire_5302)
    );

    bfr new_Jinkela_buffer_7543 (
        .din(new_Jinkela_wire_9366),
        .dout(new_Jinkela_wire_9367)
    );

    bfr new_Jinkela_buffer_3935 (
        .din(new_Jinkela_wire_5202),
        .dout(new_Jinkela_wire_5203)
    );

    bfr new_Jinkela_buffer_7403 (
        .din(new_Jinkela_wire_9218),
        .dout(new_Jinkela_wire_9219)
    );

    bfr new_Jinkela_buffer_4060 (
        .din(new_Jinkela_wire_5335),
        .dout(new_Jinkela_wire_5336)
    );

    bfr new_Jinkela_buffer_7497 (
        .din(new_Jinkela_wire_9314),
        .dout(new_Jinkela_wire_9315)
    );

    bfr new_Jinkela_buffer_3936 (
        .din(new_Jinkela_wire_5203),
        .dout(new_Jinkela_wire_5204)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_1060),
        .dout(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_976),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_1098),
        .dout(new_Jinkela_wire_1099)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_1061),
        .dout(new_Jinkela_wire_1062)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_1062),
        .dout(new_Jinkela_wire_1063)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_1148),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_980),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_1099),
        .dout(new_Jinkela_wire_1100)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_1270),
        .dout(new_Jinkela_wire_1271)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_1100),
        .dout(new_Jinkela_wire_1101)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_1101),
        .dout(new_Jinkela_wire_1102)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_1068),
        .dout(new_Jinkela_wire_1069)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_1264),
        .dout(new_Jinkela_wire_1265)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_1069),
        .dout(new_Jinkela_wire_1070)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_1070),
        .dout(new_Jinkela_wire_1071)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_1072),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_1073),
        .dout(new_Jinkela_wire_1074)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_net_3938),
        .dout(new_Jinkela_wire_1277)
    );

    spl2 new_Jinkela_splitter_200 (
        .a(new_Jinkela_wire_1074),
        .b(new_Jinkela_wire_1075),
        .c(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_1151),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_1105),
        .dout(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_1265),
        .dout(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    bfr new_Jinkela_buffer_17708 (
        .din(new_Jinkela_wire_21076),
        .dout(new_Jinkela_wire_21077)
    );

    bfr new_Jinkela_buffer_10862 (
        .din(new_Jinkela_wire_13089),
        .dout(new_Jinkela_wire_13090)
    );

    bfr new_Jinkela_buffer_10923 (
        .din(new_Jinkela_wire_13162),
        .dout(new_Jinkela_wire_13163)
    );

    spl2 new_Jinkela_splitter_1558 (
        .a(_0806_),
        .b(new_Jinkela_wire_21200),
        .c(new_Jinkela_wire_21201)
    );

    bfr new_Jinkela_buffer_17709 (
        .din(new_Jinkela_wire_21077),
        .dout(new_Jinkela_wire_21078)
    );

    bfr new_Jinkela_buffer_10863 (
        .din(new_Jinkela_wire_13090),
        .dout(new_Jinkela_wire_13091)
    );

    bfr new_Jinkela_buffer_17781 (
        .din(_0396_),
        .dout(new_Jinkela_wire_21202)
    );

    bfr new_Jinkela_buffer_17710 (
        .din(new_Jinkela_wire_21078),
        .dout(new_Jinkela_wire_21079)
    );

    bfr new_Jinkela_buffer_10864 (
        .din(new_Jinkela_wire_13091),
        .dout(new_Jinkela_wire_13092)
    );

    spl2 new_Jinkela_splitter_1559 (
        .a(_1045_),
        .b(new_Jinkela_wire_21204),
        .c(new_Jinkela_wire_21205)
    );

    bfr new_Jinkela_buffer_10924 (
        .din(new_Jinkela_wire_13163),
        .dout(new_Jinkela_wire_13164)
    );

    bfr new_Jinkela_buffer_17711 (
        .din(new_Jinkela_wire_21079),
        .dout(new_Jinkela_wire_21080)
    );

    bfr new_Jinkela_buffer_10865 (
        .din(new_Jinkela_wire_13092),
        .dout(new_Jinkela_wire_13093)
    );

    spl2 new_Jinkela_splitter_975 (
        .a(_1639_),
        .b(new_Jinkela_wire_13207),
        .c(new_Jinkela_wire_13208)
    );

    bfr new_Jinkela_buffer_17782 (
        .din(_0300_),
        .dout(new_Jinkela_wire_21203)
    );

    bfr new_Jinkela_buffer_17712 (
        .din(new_Jinkela_wire_21080),
        .dout(new_Jinkela_wire_21081)
    );

    bfr new_Jinkela_buffer_10866 (
        .din(new_Jinkela_wire_13093),
        .dout(new_Jinkela_wire_13094)
    );

    spl2 new_Jinkela_splitter_1560 (
        .a(_0154_),
        .b(new_Jinkela_wire_21206),
        .c(new_Jinkela_wire_21207)
    );

    bfr new_Jinkela_buffer_10925 (
        .din(new_Jinkela_wire_13164),
        .dout(new_Jinkela_wire_13165)
    );

    bfr new_Jinkela_buffer_17713 (
        .din(new_Jinkela_wire_21081),
        .dout(new_Jinkela_wire_21082)
    );

    bfr new_Jinkela_buffer_10867 (
        .din(new_Jinkela_wire_13094),
        .dout(new_Jinkela_wire_13095)
    );

    bfr new_Jinkela_buffer_10959 (
        .din(_0155_),
        .dout(new_Jinkela_wire_13213)
    );

    bfr new_Jinkela_buffer_17714 (
        .din(new_Jinkela_wire_21082),
        .dout(new_Jinkela_wire_21083)
    );

    bfr new_Jinkela_buffer_10868 (
        .din(new_Jinkela_wire_13095),
        .dout(new_Jinkela_wire_13096)
    );

    bfr new_Jinkela_buffer_10926 (
        .din(new_Jinkela_wire_13165),
        .dout(new_Jinkela_wire_13166)
    );

    spl2 new_Jinkela_splitter_1561 (
        .a(_1429_),
        .b(new_Jinkela_wire_21208),
        .c(new_Jinkela_wire_21209)
    );

    bfr new_Jinkela_buffer_17715 (
        .din(new_Jinkela_wire_21083),
        .dout(new_Jinkela_wire_21084)
    );

    bfr new_Jinkela_buffer_10869 (
        .din(new_Jinkela_wire_13096),
        .dout(new_Jinkela_wire_13097)
    );

    bfr new_Jinkela_buffer_10955 (
        .din(new_Jinkela_wire_13208),
        .dout(new_Jinkela_wire_13209)
    );

    spl2 new_Jinkela_splitter_976 (
        .a(_1512_),
        .b(new_Jinkela_wire_13214),
        .c(new_Jinkela_wire_13215)
    );

    spl2 new_Jinkela_splitter_1562 (
        .a(_1337_),
        .b(new_Jinkela_wire_21214),
        .c(new_Jinkela_wire_21215)
    );

    bfr new_Jinkela_buffer_17716 (
        .din(new_Jinkela_wire_21084),
        .dout(new_Jinkela_wire_21085)
    );

    bfr new_Jinkela_buffer_10870 (
        .din(new_Jinkela_wire_13097),
        .dout(new_Jinkela_wire_13098)
    );

    bfr new_Jinkela_buffer_17783 (
        .din(new_Jinkela_wire_21209),
        .dout(new_Jinkela_wire_21210)
    );

    bfr new_Jinkela_buffer_10927 (
        .din(new_Jinkela_wire_13166),
        .dout(new_Jinkela_wire_13167)
    );

    spl2 new_Jinkela_splitter_1563 (
        .a(_1204_),
        .b(new_Jinkela_wire_21216),
        .c(new_Jinkela_wire_21217)
    );

    bfr new_Jinkela_buffer_17717 (
        .din(new_Jinkela_wire_21085),
        .dout(new_Jinkela_wire_21086)
    );

    bfr new_Jinkela_buffer_10871 (
        .din(new_Jinkela_wire_13098),
        .dout(new_Jinkela_wire_13099)
    );

    bfr new_Jinkela_buffer_10960 (
        .din(_0091_),
        .dout(new_Jinkela_wire_13216)
    );

    bfr new_Jinkela_buffer_17718 (
        .din(new_Jinkela_wire_21086),
        .dout(new_Jinkela_wire_21087)
    );

    bfr new_Jinkela_buffer_10872 (
        .din(new_Jinkela_wire_13099),
        .dout(new_Jinkela_wire_13100)
    );

    bfr new_Jinkela_buffer_17784 (
        .din(new_Jinkela_wire_21210),
        .dout(new_Jinkela_wire_21211)
    );

    bfr new_Jinkela_buffer_10928 (
        .din(new_Jinkela_wire_13167),
        .dout(new_Jinkela_wire_13168)
    );

    bfr new_Jinkela_buffer_17719 (
        .din(new_Jinkela_wire_21087),
        .dout(new_Jinkela_wire_21088)
    );

    bfr new_Jinkela_buffer_10873 (
        .din(new_Jinkela_wire_13100),
        .dout(new_Jinkela_wire_13101)
    );

    bfr new_Jinkela_buffer_10956 (
        .din(new_Jinkela_wire_13209),
        .dout(new_Jinkela_wire_13210)
    );

    spl2 new_Jinkela_splitter_1564 (
        .a(_0668_),
        .b(new_Jinkela_wire_21218),
        .c(new_Jinkela_wire_21219)
    );

    bfr new_Jinkela_buffer_17720 (
        .din(new_Jinkela_wire_21088),
        .dout(new_Jinkela_wire_21089)
    );

    bfr new_Jinkela_buffer_10874 (
        .din(new_Jinkela_wire_13101),
        .dout(new_Jinkela_wire_13102)
    );

    bfr new_Jinkela_buffer_17785 (
        .din(new_Jinkela_wire_21211),
        .dout(new_Jinkela_wire_21212)
    );

    bfr new_Jinkela_buffer_10929 (
        .din(new_Jinkela_wire_13168),
        .dout(new_Jinkela_wire_13169)
    );

    spl2 new_Jinkela_splitter_1533 (
        .a(new_Jinkela_wire_21089),
        .b(new_Jinkela_wire_21090),
        .c(new_Jinkela_wire_21091)
    );

    bfr new_Jinkela_buffer_10875 (
        .din(new_Jinkela_wire_13102),
        .dout(new_Jinkela_wire_13103)
    );

    bfr new_Jinkela_buffer_17786 (
        .din(new_Jinkela_wire_21212),
        .dout(new_Jinkela_wire_21213)
    );

    bfr new_Jinkela_buffer_11049 (
        .din(_0409_),
        .dout(new_Jinkela_wire_13307)
    );

    bfr new_Jinkela_buffer_17895 (
        .din(_0316_),
        .dout(new_Jinkela_wire_21332)
    );

    bfr new_Jinkela_buffer_10876 (
        .din(new_Jinkela_wire_13103),
        .dout(new_Jinkela_wire_13104)
    );

    bfr new_Jinkela_buffer_17787 (
        .din(_0086_),
        .dout(new_Jinkela_wire_21220)
    );

    bfr new_Jinkela_buffer_10930 (
        .din(new_Jinkela_wire_13169),
        .dout(new_Jinkela_wire_13170)
    );

    spl2 new_Jinkela_splitter_1566 (
        .a(_1566_),
        .b(new_Jinkela_wire_21326),
        .c(new_Jinkela_wire_21327)
    );

    bfr new_Jinkela_buffer_17788 (
        .din(new_Jinkela_wire_21220),
        .dout(new_Jinkela_wire_21221)
    );

    bfr new_Jinkela_buffer_10877 (
        .din(new_Jinkela_wire_13104),
        .dout(new_Jinkela_wire_13105)
    );

    bfr new_Jinkela_buffer_10957 (
        .din(new_Jinkela_wire_13210),
        .dout(new_Jinkela_wire_13211)
    );

    bfr new_Jinkela_buffer_17789 (
        .din(new_Jinkela_wire_21221),
        .dout(new_Jinkela_wire_21222)
    );

    bfr new_Jinkela_buffer_10878 (
        .din(new_Jinkela_wire_13105),
        .dout(new_Jinkela_wire_13106)
    );

    bfr new_Jinkela_buffer_17891 (
        .din(new_Jinkela_wire_21327),
        .dout(new_Jinkela_wire_21328)
    );

    bfr new_Jinkela_buffer_10931 (
        .din(new_Jinkela_wire_13170),
        .dout(new_Jinkela_wire_13171)
    );

    bfr new_Jinkela_buffer_17790 (
        .din(new_Jinkela_wire_21222),
        .dout(new_Jinkela_wire_21223)
    );

    bfr new_Jinkela_buffer_10879 (
        .din(new_Jinkela_wire_13106),
        .dout(new_Jinkela_wire_13107)
    );

    bfr new_Jinkela_buffer_11048 (
        .din(_1400_),
        .dout(new_Jinkela_wire_13306)
    );

    bfr new_Jinkela_buffer_17791 (
        .din(new_Jinkela_wire_21223),
        .dout(new_Jinkela_wire_21224)
    );

    bfr new_Jinkela_buffer_10880 (
        .din(new_Jinkela_wire_13107),
        .dout(new_Jinkela_wire_13108)
    );

    bfr new_Jinkela_buffer_17892 (
        .din(new_Jinkela_wire_21328),
        .dout(new_Jinkela_wire_21329)
    );

    bfr new_Jinkela_buffer_10932 (
        .din(new_Jinkela_wire_13171),
        .dout(new_Jinkela_wire_13172)
    );

    bfr new_Jinkela_buffer_17792 (
        .din(new_Jinkela_wire_21224),
        .dout(new_Jinkela_wire_21225)
    );

    bfr new_Jinkela_buffer_10881 (
        .din(new_Jinkela_wire_13108),
        .dout(new_Jinkela_wire_13109)
    );

    bfr new_Jinkela_buffer_10958 (
        .din(new_Jinkela_wire_13211),
        .dout(new_Jinkela_wire_13212)
    );

    bfr new_Jinkela_buffer_17793 (
        .din(new_Jinkela_wire_21225),
        .dout(new_Jinkela_wire_21226)
    );

    bfr new_Jinkela_buffer_10882 (
        .din(new_Jinkela_wire_13109),
        .dout(new_Jinkela_wire_13110)
    );

    bfr new_Jinkela_buffer_17893 (
        .din(new_Jinkela_wire_21329),
        .dout(new_Jinkela_wire_21330)
    );

    bfr new_Jinkela_buffer_10933 (
        .din(new_Jinkela_wire_13172),
        .dout(new_Jinkela_wire_13173)
    );

    bfr new_Jinkela_buffer_4029 (
        .din(new_Jinkela_wire_5302),
        .dout(new_Jinkela_wire_5303)
    );

    bfr new_Jinkela_buffer_3937 (
        .din(new_Jinkela_wire_5204),
        .dout(new_Jinkela_wire_5205)
    );

    bfr new_Jinkela_buffer_14314 (
        .din(new_Jinkela_wire_17128),
        .dout(new_Jinkela_wire_17129)
    );

    bfr new_Jinkela_buffer_14505 (
        .din(new_Jinkela_wire_17321),
        .dout(new_Jinkela_wire_17322)
    );

    bfr new_Jinkela_buffer_14355 (
        .din(new_Jinkela_wire_17169),
        .dout(new_Jinkela_wire_17170)
    );

    bfr new_Jinkela_buffer_3938 (
        .din(new_Jinkela_wire_5205),
        .dout(new_Jinkela_wire_5206)
    );

    bfr new_Jinkela_buffer_14315 (
        .din(new_Jinkela_wire_17129),
        .dout(new_Jinkela_wire_17130)
    );

    bfr new_Jinkela_buffer_4030 (
        .din(new_Jinkela_wire_5303),
        .dout(new_Jinkela_wire_5304)
    );

    bfr new_Jinkela_buffer_3939 (
        .din(new_Jinkela_wire_5206),
        .dout(new_Jinkela_wire_5207)
    );

    bfr new_Jinkela_buffer_14316 (
        .din(new_Jinkela_wire_17130),
        .dout(new_Jinkela_wire_17131)
    );

    bfr new_Jinkela_buffer_4061 (
        .din(new_Jinkela_wire_5336),
        .dout(new_Jinkela_wire_5337)
    );

    bfr new_Jinkela_buffer_14508 (
        .din(new_Jinkela_wire_17324),
        .dout(new_Jinkela_wire_17325)
    );

    bfr new_Jinkela_buffer_14356 (
        .din(new_Jinkela_wire_17170),
        .dout(new_Jinkela_wire_17171)
    );

    bfr new_Jinkela_buffer_3940 (
        .din(new_Jinkela_wire_5207),
        .dout(new_Jinkela_wire_5208)
    );

    bfr new_Jinkela_buffer_14317 (
        .din(new_Jinkela_wire_17131),
        .dout(new_Jinkela_wire_17132)
    );

    bfr new_Jinkela_buffer_4031 (
        .din(new_Jinkela_wire_5304),
        .dout(new_Jinkela_wire_5305)
    );

    bfr new_Jinkela_buffer_3941 (
        .din(new_Jinkela_wire_5208),
        .dout(new_Jinkela_wire_5209)
    );

    bfr new_Jinkela_buffer_14318 (
        .din(new_Jinkela_wire_17132),
        .dout(new_Jinkela_wire_17133)
    );

    bfr new_Jinkela_buffer_4144 (
        .din(new_Jinkela_wire_5425),
        .dout(new_Jinkela_wire_5426)
    );

    spl2 new_Jinkela_splitter_1260 (
        .a(_0322_),
        .b(new_Jinkela_wire_17361),
        .c(new_Jinkela_wire_17362)
    );

    bfr new_Jinkela_buffer_14357 (
        .din(new_Jinkela_wire_17171),
        .dout(new_Jinkela_wire_17172)
    );

    bfr new_Jinkela_buffer_3942 (
        .din(new_Jinkela_wire_5209),
        .dout(new_Jinkela_wire_5210)
    );

    bfr new_Jinkela_buffer_14319 (
        .din(new_Jinkela_wire_17133),
        .dout(new_Jinkela_wire_17134)
    );

    bfr new_Jinkela_buffer_4032 (
        .din(new_Jinkela_wire_5305),
        .dout(new_Jinkela_wire_5306)
    );

    bfr new_Jinkela_buffer_3943 (
        .din(new_Jinkela_wire_5210),
        .dout(new_Jinkela_wire_5211)
    );

    bfr new_Jinkela_buffer_14320 (
        .din(new_Jinkela_wire_17134),
        .dout(new_Jinkela_wire_17135)
    );

    bfr new_Jinkela_buffer_4062 (
        .din(new_Jinkela_wire_5337),
        .dout(new_Jinkela_wire_5338)
    );

    bfr new_Jinkela_buffer_14509 (
        .din(new_Jinkela_wire_17325),
        .dout(new_Jinkela_wire_17326)
    );

    bfr new_Jinkela_buffer_14358 (
        .din(new_Jinkela_wire_17172),
        .dout(new_Jinkela_wire_17173)
    );

    bfr new_Jinkela_buffer_3944 (
        .din(new_Jinkela_wire_5211),
        .dout(new_Jinkela_wire_5212)
    );

    bfr new_Jinkela_buffer_14321 (
        .din(new_Jinkela_wire_17135),
        .dout(new_Jinkela_wire_17136)
    );

    bfr new_Jinkela_buffer_4033 (
        .din(new_Jinkela_wire_5306),
        .dout(new_Jinkela_wire_5307)
    );

    bfr new_Jinkela_buffer_3945 (
        .din(new_Jinkela_wire_5212),
        .dout(new_Jinkela_wire_5213)
    );

    bfr new_Jinkela_buffer_14322 (
        .din(new_Jinkela_wire_17136),
        .dout(new_Jinkela_wire_17137)
    );

    bfr new_Jinkela_buffer_14594 (
        .din(_0029_),
        .dout(new_Jinkela_wire_17423)
    );

    bfr new_Jinkela_buffer_4146 (
        .din(_0909_),
        .dout(new_Jinkela_wire_5434)
    );

    bfr new_Jinkela_buffer_14359 (
        .din(new_Jinkela_wire_17173),
        .dout(new_Jinkela_wire_17174)
    );

    bfr new_Jinkela_buffer_3946 (
        .din(new_Jinkela_wire_5213),
        .dout(new_Jinkela_wire_5214)
    );

    bfr new_Jinkela_buffer_14323 (
        .din(new_Jinkela_wire_17137),
        .dout(new_Jinkela_wire_17138)
    );

    bfr new_Jinkela_buffer_4034 (
        .din(new_Jinkela_wire_5307),
        .dout(new_Jinkela_wire_5308)
    );

    bfr new_Jinkela_buffer_14538 (
        .din(_0339_),
        .dout(new_Jinkela_wire_17363)
    );

    bfr new_Jinkela_buffer_3947 (
        .din(new_Jinkela_wire_5214),
        .dout(new_Jinkela_wire_5215)
    );

    bfr new_Jinkela_buffer_14324 (
        .din(new_Jinkela_wire_17138),
        .dout(new_Jinkela_wire_17139)
    );

    bfr new_Jinkela_buffer_4063 (
        .din(new_Jinkela_wire_5338),
        .dout(new_Jinkela_wire_5339)
    );

    bfr new_Jinkela_buffer_14510 (
        .din(new_Jinkela_wire_17326),
        .dout(new_Jinkela_wire_17327)
    );

    bfr new_Jinkela_buffer_14360 (
        .din(new_Jinkela_wire_17174),
        .dout(new_Jinkela_wire_17175)
    );

    bfr new_Jinkela_buffer_3948 (
        .din(new_Jinkela_wire_5215),
        .dout(new_Jinkela_wire_5216)
    );

    bfr new_Jinkela_buffer_14325 (
        .din(new_Jinkela_wire_17139),
        .dout(new_Jinkela_wire_17140)
    );

    bfr new_Jinkela_buffer_4035 (
        .din(new_Jinkela_wire_5308),
        .dout(new_Jinkela_wire_5309)
    );

    bfr new_Jinkela_buffer_3949 (
        .din(new_Jinkela_wire_5216),
        .dout(new_Jinkela_wire_5217)
    );

    bfr new_Jinkela_buffer_14326 (
        .din(new_Jinkela_wire_17140),
        .dout(new_Jinkela_wire_17141)
    );

    bfr new_Jinkela_buffer_4145 (
        .din(new_Jinkela_wire_5426),
        .dout(new_Jinkela_wire_5427)
    );

    bfr new_Jinkela_buffer_14361 (
        .din(new_Jinkela_wire_17175),
        .dout(new_Jinkela_wire_17176)
    );

    bfr new_Jinkela_buffer_3950 (
        .din(new_Jinkela_wire_5217),
        .dout(new_Jinkela_wire_5218)
    );

    bfr new_Jinkela_buffer_14327 (
        .din(new_Jinkela_wire_17141),
        .dout(new_Jinkela_wire_17142)
    );

    bfr new_Jinkela_buffer_4036 (
        .din(new_Jinkela_wire_5309),
        .dout(new_Jinkela_wire_5310)
    );

    bfr new_Jinkela_buffer_14546 (
        .din(_1072_),
        .dout(new_Jinkela_wire_17373)
    );

    bfr new_Jinkela_buffer_3951 (
        .din(new_Jinkela_wire_5218),
        .dout(new_Jinkela_wire_5219)
    );

    bfr new_Jinkela_buffer_14328 (
        .din(new_Jinkela_wire_17142),
        .dout(new_Jinkela_wire_17143)
    );

    bfr new_Jinkela_buffer_4064 (
        .din(new_Jinkela_wire_5339),
        .dout(new_Jinkela_wire_5340)
    );

    bfr new_Jinkela_buffer_14511 (
        .din(new_Jinkela_wire_17327),
        .dout(new_Jinkela_wire_17328)
    );

    bfr new_Jinkela_buffer_14362 (
        .din(new_Jinkela_wire_17176),
        .dout(new_Jinkela_wire_17177)
    );

    bfr new_Jinkela_buffer_3952 (
        .din(new_Jinkela_wire_5219),
        .dout(new_Jinkela_wire_5220)
    );

    bfr new_Jinkela_buffer_14329 (
        .din(new_Jinkela_wire_17143),
        .dout(new_Jinkela_wire_17144)
    );

    bfr new_Jinkela_buffer_4037 (
        .din(new_Jinkela_wire_5310),
        .dout(new_Jinkela_wire_5311)
    );

    bfr new_Jinkela_buffer_3953 (
        .din(new_Jinkela_wire_5220),
        .dout(new_Jinkela_wire_5221)
    );

    bfr new_Jinkela_buffer_14330 (
        .din(new_Jinkela_wire_17144),
        .dout(new_Jinkela_wire_17145)
    );

    spl2 new_Jinkela_splitter_494 (
        .a(_0226_),
        .b(new_Jinkela_wire_5437),
        .c(new_Jinkela_wire_5438)
    );

    bfr new_Jinkela_buffer_14539 (
        .din(new_Jinkela_wire_17363),
        .dout(new_Jinkela_wire_17364)
    );

    spl2 new_Jinkela_splitter_493 (
        .a(_1287_),
        .b(new_Jinkela_wire_5435),
        .c(new_Jinkela_wire_5436)
    );

    bfr new_Jinkela_buffer_14363 (
        .din(new_Jinkela_wire_17177),
        .dout(new_Jinkela_wire_17178)
    );

    bfr new_Jinkela_buffer_3954 (
        .din(new_Jinkela_wire_5221),
        .dout(new_Jinkela_wire_5222)
    );

    bfr new_Jinkela_buffer_14331 (
        .din(new_Jinkela_wire_17145),
        .dout(new_Jinkela_wire_17146)
    );

    bfr new_Jinkela_buffer_4038 (
        .din(new_Jinkela_wire_5311),
        .dout(new_Jinkela_wire_5312)
    );

    bfr new_Jinkela_buffer_3955 (
        .din(new_Jinkela_wire_5222),
        .dout(new_Jinkela_wire_5223)
    );

    bfr new_Jinkela_buffer_14332 (
        .din(new_Jinkela_wire_17146),
        .dout(new_Jinkela_wire_17147)
    );

    bfr new_Jinkela_buffer_4065 (
        .din(new_Jinkela_wire_5340),
        .dout(new_Jinkela_wire_5341)
    );

    bfr new_Jinkela_buffer_14512 (
        .din(new_Jinkela_wire_17328),
        .dout(new_Jinkela_wire_17329)
    );

    bfr new_Jinkela_buffer_14364 (
        .din(new_Jinkela_wire_17178),
        .dout(new_Jinkela_wire_17179)
    );

    bfr new_Jinkela_buffer_3956 (
        .din(new_Jinkela_wire_5223),
        .dout(new_Jinkela_wire_5224)
    );

    bfr new_Jinkela_buffer_14333 (
        .din(new_Jinkela_wire_17147),
        .dout(new_Jinkela_wire_17148)
    );

    bfr new_Jinkela_buffer_4039 (
        .din(new_Jinkela_wire_5312),
        .dout(new_Jinkela_wire_5313)
    );

    bfr new_Jinkela_buffer_3957 (
        .din(new_Jinkela_wire_5224),
        .dout(new_Jinkela_wire_5225)
    );

    bfr new_Jinkela_buffer_14334 (
        .din(new_Jinkela_wire_17148),
        .dout(new_Jinkela_wire_17149)
    );

    bfr new_Jinkela_buffer_10883 (
        .din(new_Jinkela_wire_13110),
        .dout(new_Jinkela_wire_13111)
    );

    bfr new_Jinkela_buffer_10961 (
        .din(new_Jinkela_wire_13216),
        .dout(new_Jinkela_wire_13217)
    );

    bfr new_Jinkela_buffer_10884 (
        .din(new_Jinkela_wire_13111),
        .dout(new_Jinkela_wire_13112)
    );

    bfr new_Jinkela_buffer_10934 (
        .din(new_Jinkela_wire_13173),
        .dout(new_Jinkela_wire_13174)
    );

    bfr new_Jinkela_buffer_10885 (
        .din(new_Jinkela_wire_13112),
        .dout(new_Jinkela_wire_13113)
    );

    spl2 new_Jinkela_splitter_978 (
        .a(_0480_),
        .b(new_Jinkela_wire_13308),
        .c(new_Jinkela_wire_13309)
    );

    bfr new_Jinkela_buffer_10886 (
        .din(new_Jinkela_wire_13113),
        .dout(new_Jinkela_wire_13114)
    );

    bfr new_Jinkela_buffer_10935 (
        .din(new_Jinkela_wire_13174),
        .dout(new_Jinkela_wire_13175)
    );

    bfr new_Jinkela_buffer_10887 (
        .din(new_Jinkela_wire_13114),
        .dout(new_Jinkela_wire_13115)
    );

    bfr new_Jinkela_buffer_10962 (
        .din(new_Jinkela_wire_13217),
        .dout(new_Jinkela_wire_13218)
    );

    bfr new_Jinkela_buffer_10888 (
        .din(new_Jinkela_wire_13115),
        .dout(new_Jinkela_wire_13116)
    );

    bfr new_Jinkela_buffer_10936 (
        .din(new_Jinkela_wire_13175),
        .dout(new_Jinkela_wire_13176)
    );

    bfr new_Jinkela_buffer_10889 (
        .din(new_Jinkela_wire_13116),
        .dout(new_Jinkela_wire_13117)
    );

    spl2 new_Jinkela_splitter_979 (
        .a(_0092_),
        .b(new_Jinkela_wire_13310),
        .c(new_Jinkela_wire_13311)
    );

    bfr new_Jinkela_buffer_10890 (
        .din(new_Jinkela_wire_13117),
        .dout(new_Jinkela_wire_13118)
    );

    bfr new_Jinkela_buffer_10937 (
        .din(new_Jinkela_wire_13176),
        .dout(new_Jinkela_wire_13177)
    );

    bfr new_Jinkela_buffer_10891 (
        .din(new_Jinkela_wire_13118),
        .dout(new_Jinkela_wire_13119)
    );

    bfr new_Jinkela_buffer_10963 (
        .din(new_Jinkela_wire_13218),
        .dout(new_Jinkela_wire_13219)
    );

    bfr new_Jinkela_buffer_10892 (
        .din(new_Jinkela_wire_13119),
        .dout(new_Jinkela_wire_13120)
    );

    bfr new_Jinkela_buffer_10938 (
        .din(new_Jinkela_wire_13177),
        .dout(new_Jinkela_wire_13178)
    );

    bfr new_Jinkela_buffer_10893 (
        .din(new_Jinkela_wire_13120),
        .dout(new_Jinkela_wire_13121)
    );

    bfr new_Jinkela_buffer_10894 (
        .din(new_Jinkela_wire_13121),
        .dout(new_Jinkela_wire_13122)
    );

    bfr new_Jinkela_buffer_10939 (
        .din(new_Jinkela_wire_13178),
        .dout(new_Jinkela_wire_13179)
    );

    bfr new_Jinkela_buffer_10895 (
        .din(new_Jinkela_wire_13122),
        .dout(new_Jinkela_wire_13123)
    );

    bfr new_Jinkela_buffer_10964 (
        .din(new_Jinkela_wire_13219),
        .dout(new_Jinkela_wire_13220)
    );

    bfr new_Jinkela_buffer_10896 (
        .din(new_Jinkela_wire_13123),
        .dout(new_Jinkela_wire_13124)
    );

    bfr new_Jinkela_buffer_10940 (
        .din(new_Jinkela_wire_13179),
        .dout(new_Jinkela_wire_13180)
    );

    bfr new_Jinkela_buffer_10897 (
        .din(new_Jinkela_wire_13124),
        .dout(new_Jinkela_wire_13125)
    );

    spl2 new_Jinkela_splitter_980 (
        .a(_0869_),
        .b(new_Jinkela_wire_13312),
        .c(new_Jinkela_wire_13313)
    );

    bfr new_Jinkela_buffer_10898 (
        .din(new_Jinkela_wire_13125),
        .dout(new_Jinkela_wire_13126)
    );

    bfr new_Jinkela_buffer_10941 (
        .din(new_Jinkela_wire_13180),
        .dout(new_Jinkela_wire_13181)
    );

    bfr new_Jinkela_buffer_10899 (
        .din(new_Jinkela_wire_13126),
        .dout(new_Jinkela_wire_13127)
    );

    bfr new_Jinkela_buffer_10965 (
        .din(new_Jinkela_wire_13220),
        .dout(new_Jinkela_wire_13221)
    );

    bfr new_Jinkela_buffer_10900 (
        .din(new_Jinkela_wire_13127),
        .dout(new_Jinkela_wire_13128)
    );

    bfr new_Jinkela_buffer_10942 (
        .din(new_Jinkela_wire_13181),
        .dout(new_Jinkela_wire_13182)
    );

    bfr new_Jinkela_buffer_10901 (
        .din(new_Jinkela_wire_13128),
        .dout(new_Jinkela_wire_13129)
    );

    spl2 new_Jinkela_splitter_982 (
        .a(_1124_),
        .b(new_Jinkela_wire_13316),
        .c(new_Jinkela_wire_13317)
    );

    spl2 new_Jinkela_splitter_981 (
        .a(_1212_),
        .b(new_Jinkela_wire_13314),
        .c(new_Jinkela_wire_13315)
    );

    bfr new_Jinkela_buffer_10902 (
        .din(new_Jinkela_wire_13129),
        .dout(new_Jinkela_wire_13130)
    );

    bfr new_Jinkela_buffer_10943 (
        .din(new_Jinkela_wire_13182),
        .dout(new_Jinkela_wire_13183)
    );

    bfr new_Jinkela_buffer_10903 (
        .din(new_Jinkela_wire_13130),
        .dout(new_Jinkela_wire_13131)
    );

    bfr new_Jinkela_buffer_10966 (
        .din(new_Jinkela_wire_13221),
        .dout(new_Jinkela_wire_13222)
    );

    bfr new_Jinkela_buffer_7404 (
        .din(new_Jinkela_wire_9219),
        .dout(new_Jinkela_wire_9220)
    );

    bfr new_Jinkela_buffer_7535 (
        .din(new_Jinkela_wire_9356),
        .dout(new_Jinkela_wire_9357)
    );

    bfr new_Jinkela_buffer_7405 (
        .din(new_Jinkela_wire_9220),
        .dout(new_Jinkela_wire_9221)
    );

    bfr new_Jinkela_buffer_7498 (
        .din(new_Jinkela_wire_9315),
        .dout(new_Jinkela_wire_9316)
    );

    bfr new_Jinkela_buffer_7406 (
        .din(new_Jinkela_wire_9221),
        .dout(new_Jinkela_wire_9222)
    );

    spl2 new_Jinkela_splitter_764 (
        .a(_1526_),
        .b(new_Jinkela_wire_9521),
        .c(new_Jinkela_wire_9522)
    );

    bfr new_Jinkela_buffer_7407 (
        .din(new_Jinkela_wire_9222),
        .dout(new_Jinkela_wire_9223)
    );

    bfr new_Jinkela_buffer_7499 (
        .din(new_Jinkela_wire_9316),
        .dout(new_Jinkela_wire_9317)
    );

    bfr new_Jinkela_buffer_7408 (
        .din(new_Jinkela_wire_9223),
        .dout(new_Jinkela_wire_9224)
    );

    bfr new_Jinkela_buffer_7536 (
        .din(new_Jinkela_wire_9357),
        .dout(new_Jinkela_wire_9358)
    );

    bfr new_Jinkela_buffer_7409 (
        .din(new_Jinkela_wire_9224),
        .dout(new_Jinkela_wire_9225)
    );

    bfr new_Jinkela_buffer_7500 (
        .din(new_Jinkela_wire_9317),
        .dout(new_Jinkela_wire_9318)
    );

    bfr new_Jinkela_buffer_7410 (
        .din(new_Jinkela_wire_9225),
        .dout(new_Jinkela_wire_9226)
    );

    bfr new_Jinkela_buffer_7544 (
        .din(new_Jinkela_wire_9367),
        .dout(new_Jinkela_wire_9368)
    );

    bfr new_Jinkela_buffer_7411 (
        .din(new_Jinkela_wire_9226),
        .dout(new_Jinkela_wire_9227)
    );

    bfr new_Jinkela_buffer_7501 (
        .din(new_Jinkela_wire_9318),
        .dout(new_Jinkela_wire_9319)
    );

    bfr new_Jinkela_buffer_7412 (
        .din(new_Jinkela_wire_9227),
        .dout(new_Jinkela_wire_9228)
    );

    bfr new_Jinkela_buffer_7537 (
        .din(new_Jinkela_wire_9358),
        .dout(new_Jinkela_wire_9359)
    );

    bfr new_Jinkela_buffer_7413 (
        .din(new_Jinkela_wire_9228),
        .dout(new_Jinkela_wire_9229)
    );

    bfr new_Jinkela_buffer_7502 (
        .din(new_Jinkela_wire_9319),
        .dout(new_Jinkela_wire_9320)
    );

    bfr new_Jinkela_buffer_7414 (
        .din(new_Jinkela_wire_9229),
        .dout(new_Jinkela_wire_9230)
    );

    bfr new_Jinkela_buffer_7621 (
        .din(new_Jinkela_wire_9448),
        .dout(new_Jinkela_wire_9449)
    );

    bfr new_Jinkela_buffer_7415 (
        .din(new_Jinkela_wire_9230),
        .dout(new_Jinkela_wire_9231)
    );

    bfr new_Jinkela_buffer_7503 (
        .din(new_Jinkela_wire_9320),
        .dout(new_Jinkela_wire_9321)
    );

    bfr new_Jinkela_buffer_7416 (
        .din(new_Jinkela_wire_9231),
        .dout(new_Jinkela_wire_9232)
    );

    bfr new_Jinkela_buffer_7538 (
        .din(new_Jinkela_wire_9359),
        .dout(new_Jinkela_wire_9360)
    );

    bfr new_Jinkela_buffer_7417 (
        .din(new_Jinkela_wire_9232),
        .dout(new_Jinkela_wire_9233)
    );

    bfr new_Jinkela_buffer_7504 (
        .din(new_Jinkela_wire_9321),
        .dout(new_Jinkela_wire_9322)
    );

    bfr new_Jinkela_buffer_7418 (
        .din(new_Jinkela_wire_9233),
        .dout(new_Jinkela_wire_9234)
    );

    bfr new_Jinkela_buffer_7545 (
        .din(new_Jinkela_wire_9368),
        .dout(new_Jinkela_wire_9369)
    );

    bfr new_Jinkela_buffer_7419 (
        .din(new_Jinkela_wire_9234),
        .dout(new_Jinkela_wire_9235)
    );

    bfr new_Jinkela_buffer_7505 (
        .din(new_Jinkela_wire_9322),
        .dout(new_Jinkela_wire_9323)
    );

    bfr new_Jinkela_buffer_7420 (
        .din(new_Jinkela_wire_9235),
        .dout(new_Jinkela_wire_9236)
    );

    bfr new_Jinkela_buffer_7539 (
        .din(new_Jinkela_wire_9360),
        .dout(new_Jinkela_wire_9361)
    );

    bfr new_Jinkela_buffer_7421 (
        .din(new_Jinkela_wire_9236),
        .dout(new_Jinkela_wire_9237)
    );

    bfr new_Jinkela_buffer_7506 (
        .din(new_Jinkela_wire_9323),
        .dout(new_Jinkela_wire_9324)
    );

    bfr new_Jinkela_buffer_7422 (
        .din(new_Jinkela_wire_9237),
        .dout(new_Jinkela_wire_9238)
    );

    bfr new_Jinkela_buffer_7683 (
        .din(new_Jinkela_wire_9510),
        .dout(new_Jinkela_wire_9511)
    );

    bfr new_Jinkela_buffer_7423 (
        .din(new_Jinkela_wire_9238),
        .dout(new_Jinkela_wire_9239)
    );

    bfr new_Jinkela_buffer_7507 (
        .din(new_Jinkela_wire_9324),
        .dout(new_Jinkela_wire_9325)
    );

    bfr new_Jinkela_buffer_7424 (
        .din(new_Jinkela_wire_9239),
        .dout(new_Jinkela_wire_9240)
    );

    spl2 new_Jinkela_splitter_760 (
        .a(new_Jinkela_wire_9361),
        .b(new_Jinkela_wire_9362),
        .c(new_Jinkela_wire_9363)
    );

    bfr new_Jinkela_buffer_14365 (
        .din(new_Jinkela_wire_17179),
        .dout(new_Jinkela_wire_17180)
    );

    bfr new_Jinkela_buffer_14335 (
        .din(new_Jinkela_wire_17149),
        .dout(new_Jinkela_wire_17150)
    );

    bfr new_Jinkela_buffer_3958 (
        .din(new_Jinkela_wire_5225),
        .dout(new_Jinkela_wire_5226)
    );

    bfr new_Jinkela_buffer_4040 (
        .din(new_Jinkela_wire_5313),
        .dout(new_Jinkela_wire_5314)
    );

    spl2 new_Jinkela_splitter_1263 (
        .a(_1457_),
        .b(new_Jinkela_wire_17424),
        .c(new_Jinkela_wire_17425)
    );

    bfr new_Jinkela_buffer_14336 (
        .din(new_Jinkela_wire_17150),
        .dout(new_Jinkela_wire_17151)
    );

    bfr new_Jinkela_buffer_3959 (
        .din(new_Jinkela_wire_5226),
        .dout(new_Jinkela_wire_5227)
    );

    bfr new_Jinkela_buffer_14513 (
        .din(new_Jinkela_wire_17329),
        .dout(new_Jinkela_wire_17330)
    );

    bfr new_Jinkela_buffer_4066 (
        .din(new_Jinkela_wire_5341),
        .dout(new_Jinkela_wire_5342)
    );

    bfr new_Jinkela_buffer_14366 (
        .din(new_Jinkela_wire_17180),
        .dout(new_Jinkela_wire_17181)
    );

    bfr new_Jinkela_buffer_14337 (
        .din(new_Jinkela_wire_17151),
        .dout(new_Jinkela_wire_17152)
    );

    bfr new_Jinkela_buffer_3960 (
        .din(new_Jinkela_wire_5227),
        .dout(new_Jinkela_wire_5228)
    );

    bfr new_Jinkela_buffer_4041 (
        .din(new_Jinkela_wire_5314),
        .dout(new_Jinkela_wire_5315)
    );

    bfr new_Jinkela_buffer_14338 (
        .din(new_Jinkela_wire_17152),
        .dout(new_Jinkela_wire_17153)
    );

    bfr new_Jinkela_buffer_3961 (
        .din(new_Jinkela_wire_5228),
        .dout(new_Jinkela_wire_5229)
    );

    bfr new_Jinkela_buffer_14540 (
        .din(new_Jinkela_wire_17364),
        .dout(new_Jinkela_wire_17365)
    );

    spl2 new_Jinkela_splitter_495 (
        .a(_1177_),
        .b(new_Jinkela_wire_5439),
        .c(new_Jinkela_wire_5440)
    );

    bfr new_Jinkela_buffer_14367 (
        .din(new_Jinkela_wire_17181),
        .dout(new_Jinkela_wire_17182)
    );

    bfr new_Jinkela_buffer_14339 (
        .din(new_Jinkela_wire_17153),
        .dout(new_Jinkela_wire_17154)
    );

    bfr new_Jinkela_buffer_3962 (
        .din(new_Jinkela_wire_5229),
        .dout(new_Jinkela_wire_5230)
    );

    bfr new_Jinkela_buffer_4042 (
        .din(new_Jinkela_wire_5315),
        .dout(new_Jinkela_wire_5316)
    );

    bfr new_Jinkela_buffer_14340 (
        .din(new_Jinkela_wire_17154),
        .dout(new_Jinkela_wire_17155)
    );

    bfr new_Jinkela_buffer_3963 (
        .din(new_Jinkela_wire_5230),
        .dout(new_Jinkela_wire_5231)
    );

    bfr new_Jinkela_buffer_14514 (
        .din(new_Jinkela_wire_17330),
        .dout(new_Jinkela_wire_17331)
    );

    bfr new_Jinkela_buffer_4067 (
        .din(new_Jinkela_wire_5342),
        .dout(new_Jinkela_wire_5343)
    );

    bfr new_Jinkela_buffer_14368 (
        .din(new_Jinkela_wire_17182),
        .dout(new_Jinkela_wire_17183)
    );

    bfr new_Jinkela_buffer_14341 (
        .din(new_Jinkela_wire_17155),
        .dout(new_Jinkela_wire_17156)
    );

    bfr new_Jinkela_buffer_3964 (
        .din(new_Jinkela_wire_5231),
        .dout(new_Jinkela_wire_5232)
    );

    bfr new_Jinkela_buffer_4043 (
        .din(new_Jinkela_wire_5316),
        .dout(new_Jinkela_wire_5317)
    );

    bfr new_Jinkela_buffer_14342 (
        .din(new_Jinkela_wire_17156),
        .dout(new_Jinkela_wire_17157)
    );

    bfr new_Jinkela_buffer_3965 (
        .din(new_Jinkela_wire_5232),
        .dout(new_Jinkela_wire_5233)
    );

    bfr new_Jinkela_buffer_14547 (
        .din(new_Jinkela_wire_17373),
        .dout(new_Jinkela_wire_17374)
    );

    spl2 new_Jinkela_splitter_496 (
        .a(_0410_),
        .b(new_Jinkela_wire_5441),
        .c(new_Jinkela_wire_5442)
    );

    bfr new_Jinkela_buffer_14369 (
        .din(new_Jinkela_wire_17183),
        .dout(new_Jinkela_wire_17184)
    );

    bfr new_Jinkela_buffer_14343 (
        .din(new_Jinkela_wire_17157),
        .dout(new_Jinkela_wire_17158)
    );

    bfr new_Jinkela_buffer_3966 (
        .din(new_Jinkela_wire_5233),
        .dout(new_Jinkela_wire_5234)
    );

    bfr new_Jinkela_buffer_4044 (
        .din(new_Jinkela_wire_5317),
        .dout(new_Jinkela_wire_5318)
    );

    bfr new_Jinkela_buffer_14344 (
        .din(new_Jinkela_wire_17158),
        .dout(new_Jinkela_wire_17159)
    );

    bfr new_Jinkela_buffer_3967 (
        .din(new_Jinkela_wire_5234),
        .dout(new_Jinkela_wire_5235)
    );

    bfr new_Jinkela_buffer_14515 (
        .din(new_Jinkela_wire_17331),
        .dout(new_Jinkela_wire_17332)
    );

    bfr new_Jinkela_buffer_4068 (
        .din(new_Jinkela_wire_5343),
        .dout(new_Jinkela_wire_5344)
    );

    bfr new_Jinkela_buffer_14370 (
        .din(new_Jinkela_wire_17184),
        .dout(new_Jinkela_wire_17185)
    );

    bfr new_Jinkela_buffer_14345 (
        .din(new_Jinkela_wire_17159),
        .dout(new_Jinkela_wire_17160)
    );

    bfr new_Jinkela_buffer_3968 (
        .din(new_Jinkela_wire_5235),
        .dout(new_Jinkela_wire_5236)
    );

    bfr new_Jinkela_buffer_4045 (
        .din(new_Jinkela_wire_5318),
        .dout(new_Jinkela_wire_5319)
    );

    bfr new_Jinkela_buffer_14541 (
        .din(new_Jinkela_wire_17365),
        .dout(new_Jinkela_wire_17366)
    );

    bfr new_Jinkela_buffer_3969 (
        .din(new_Jinkela_wire_5236),
        .dout(new_Jinkela_wire_5237)
    );

    bfr new_Jinkela_buffer_14371 (
        .din(new_Jinkela_wire_17185),
        .dout(new_Jinkela_wire_17186)
    );

    spl2 new_Jinkela_splitter_497 (
        .a(_0235_),
        .b(new_Jinkela_wire_5443),
        .c(new_Jinkela_wire_5444)
    );

    bfr new_Jinkela_buffer_14516 (
        .din(new_Jinkela_wire_17332),
        .dout(new_Jinkela_wire_17333)
    );

    bfr new_Jinkela_buffer_3970 (
        .din(new_Jinkela_wire_5237),
        .dout(new_Jinkela_wire_5238)
    );

    bfr new_Jinkela_buffer_14372 (
        .din(new_Jinkela_wire_17186),
        .dout(new_Jinkela_wire_17187)
    );

    bfr new_Jinkela_buffer_4046 (
        .din(new_Jinkela_wire_5319),
        .dout(new_Jinkela_wire_5320)
    );

    bfr new_Jinkela_buffer_14595 (
        .din(_1680_),
        .dout(new_Jinkela_wire_17426)
    );

    bfr new_Jinkela_buffer_3971 (
        .din(new_Jinkela_wire_5238),
        .dout(new_Jinkela_wire_5239)
    );

    bfr new_Jinkela_buffer_14373 (
        .din(new_Jinkela_wire_17187),
        .dout(new_Jinkela_wire_17188)
    );

    bfr new_Jinkela_buffer_4069 (
        .din(new_Jinkela_wire_5344),
        .dout(new_Jinkela_wire_5345)
    );

    bfr new_Jinkela_buffer_14517 (
        .din(new_Jinkela_wire_17333),
        .dout(new_Jinkela_wire_17334)
    );

    bfr new_Jinkela_buffer_3972 (
        .din(new_Jinkela_wire_5239),
        .dout(new_Jinkela_wire_5240)
    );

    bfr new_Jinkela_buffer_14374 (
        .din(new_Jinkela_wire_17188),
        .dout(new_Jinkela_wire_17189)
    );

    bfr new_Jinkela_buffer_4047 (
        .din(new_Jinkela_wire_5320),
        .dout(new_Jinkela_wire_5321)
    );

    bfr new_Jinkela_buffer_14542 (
        .din(new_Jinkela_wire_17366),
        .dout(new_Jinkela_wire_17367)
    );

    bfr new_Jinkela_buffer_3973 (
        .din(new_Jinkela_wire_5240),
        .dout(new_Jinkela_wire_5241)
    );

    bfr new_Jinkela_buffer_14375 (
        .din(new_Jinkela_wire_17189),
        .dout(new_Jinkela_wire_17190)
    );

    spl2 new_Jinkela_splitter_498 (
        .a(_0281_),
        .b(new_Jinkela_wire_5445),
        .c(new_Jinkela_wire_5446)
    );

    bfr new_Jinkela_buffer_14518 (
        .din(new_Jinkela_wire_17334),
        .dout(new_Jinkela_wire_17335)
    );

    bfr new_Jinkela_buffer_3974 (
        .din(new_Jinkela_wire_5241),
        .dout(new_Jinkela_wire_5242)
    );

    bfr new_Jinkela_buffer_14376 (
        .din(new_Jinkela_wire_17190),
        .dout(new_Jinkela_wire_17191)
    );

    bfr new_Jinkela_buffer_4048 (
        .din(new_Jinkela_wire_5321),
        .dout(new_Jinkela_wire_5322)
    );

    bfr new_Jinkela_buffer_14548 (
        .din(new_Jinkela_wire_17374),
        .dout(new_Jinkela_wire_17375)
    );

    bfr new_Jinkela_buffer_3975 (
        .din(new_Jinkela_wire_5242),
        .dout(new_Jinkela_wire_5243)
    );

    bfr new_Jinkela_buffer_14377 (
        .din(new_Jinkela_wire_17191),
        .dout(new_Jinkela_wire_17192)
    );

    bfr new_Jinkela_buffer_4070 (
        .din(new_Jinkela_wire_5345),
        .dout(new_Jinkela_wire_5346)
    );

    bfr new_Jinkela_buffer_14519 (
        .din(new_Jinkela_wire_17335),
        .dout(new_Jinkela_wire_17336)
    );

    bfr new_Jinkela_buffer_3976 (
        .din(new_Jinkela_wire_5243),
        .dout(new_Jinkela_wire_5244)
    );

    bfr new_Jinkela_buffer_14378 (
        .din(new_Jinkela_wire_17192),
        .dout(new_Jinkela_wire_17193)
    );

    bfr new_Jinkela_buffer_4049 (
        .din(new_Jinkela_wire_5322),
        .dout(new_Jinkela_wire_5323)
    );

    bfr new_Jinkela_buffer_14543 (
        .din(new_Jinkela_wire_17367),
        .dout(new_Jinkela_wire_17368)
    );

    bfr new_Jinkela_buffer_3977 (
        .din(new_Jinkela_wire_5244),
        .dout(new_Jinkela_wire_5245)
    );

    bfr new_Jinkela_buffer_14379 (
        .din(new_Jinkela_wire_17193),
        .dout(new_Jinkela_wire_17194)
    );

    spl2 new_Jinkela_splitter_499 (
        .a(_0556_),
        .b(new_Jinkela_wire_5448),
        .c(new_Jinkela_wire_5449)
    );

    bfr new_Jinkela_buffer_4147 (
        .din(_1235_),
        .dout(new_Jinkela_wire_5447)
    );

    bfr new_Jinkela_buffer_14520 (
        .din(new_Jinkela_wire_17336),
        .dout(new_Jinkela_wire_17337)
    );

    bfr new_Jinkela_buffer_3978 (
        .din(new_Jinkela_wire_5245),
        .dout(new_Jinkela_wire_5246)
    );

    bfr new_Jinkela_buffer_14380 (
        .din(new_Jinkela_wire_17194),
        .dout(new_Jinkela_wire_17195)
    );

    bfr new_Jinkela_buffer_10904 (
        .din(new_Jinkela_wire_13131),
        .dout(new_Jinkela_wire_13132)
    );

    bfr new_Jinkela_buffer_10944 (
        .din(new_Jinkela_wire_13183),
        .dout(new_Jinkela_wire_13184)
    );

    bfr new_Jinkela_buffer_10905 (
        .din(new_Jinkela_wire_13132),
        .dout(new_Jinkela_wire_13133)
    );

    bfr new_Jinkela_buffer_10906 (
        .din(new_Jinkela_wire_13133),
        .dout(new_Jinkela_wire_13134)
    );

    bfr new_Jinkela_buffer_10945 (
        .din(new_Jinkela_wire_13184),
        .dout(new_Jinkela_wire_13185)
    );

    bfr new_Jinkela_buffer_10907 (
        .din(new_Jinkela_wire_13134),
        .dout(new_Jinkela_wire_13135)
    );

    bfr new_Jinkela_buffer_10967 (
        .din(new_Jinkela_wire_13222),
        .dout(new_Jinkela_wire_13223)
    );

    bfr new_Jinkela_buffer_10908 (
        .din(new_Jinkela_wire_13135),
        .dout(new_Jinkela_wire_13136)
    );

    bfr new_Jinkela_buffer_10946 (
        .din(new_Jinkela_wire_13185),
        .dout(new_Jinkela_wire_13186)
    );

    bfr new_Jinkela_buffer_10909 (
        .din(new_Jinkela_wire_13136),
        .dout(new_Jinkela_wire_13137)
    );

    bfr new_Jinkela_buffer_11054 (
        .din(_0171_),
        .dout(new_Jinkela_wire_13322)
    );

    bfr new_Jinkela_buffer_10910 (
        .din(new_Jinkela_wire_13137),
        .dout(new_Jinkela_wire_13138)
    );

    bfr new_Jinkela_buffer_10947 (
        .din(new_Jinkela_wire_13186),
        .dout(new_Jinkela_wire_13187)
    );

    spl2 new_Jinkela_splitter_963 (
        .a(new_Jinkela_wire_13138),
        .b(new_Jinkela_wire_13139),
        .c(new_Jinkela_wire_13140)
    );

    bfr new_Jinkela_buffer_10948 (
        .din(new_Jinkela_wire_13187),
        .dout(new_Jinkela_wire_13188)
    );

    bfr new_Jinkela_buffer_10968 (
        .din(new_Jinkela_wire_13223),
        .dout(new_Jinkela_wire_13224)
    );

    bfr new_Jinkela_buffer_11050 (
        .din(new_Jinkela_wire_13317),
        .dout(new_Jinkela_wire_13318)
    );

    spl2 new_Jinkela_splitter_983 (
        .a(_1264_),
        .b(new_Jinkela_wire_13323),
        .c(new_Jinkela_wire_13324)
    );

    bfr new_Jinkela_buffer_10949 (
        .din(new_Jinkela_wire_13188),
        .dout(new_Jinkela_wire_13189)
    );

    bfr new_Jinkela_buffer_10969 (
        .din(new_Jinkela_wire_13224),
        .dout(new_Jinkela_wire_13225)
    );

    bfr new_Jinkela_buffer_10950 (
        .din(new_Jinkela_wire_13189),
        .dout(new_Jinkela_wire_13190)
    );

    bfr new_Jinkela_buffer_11055 (
        .din(_0112_),
        .dout(new_Jinkela_wire_13325)
    );

    bfr new_Jinkela_buffer_10951 (
        .din(new_Jinkela_wire_13190),
        .dout(new_Jinkela_wire_13191)
    );

    bfr new_Jinkela_buffer_10970 (
        .din(new_Jinkela_wire_13225),
        .dout(new_Jinkela_wire_13226)
    );

    bfr new_Jinkela_buffer_10952 (
        .din(new_Jinkela_wire_13191),
        .dout(new_Jinkela_wire_13192)
    );

    bfr new_Jinkela_buffer_11051 (
        .din(new_Jinkela_wire_13318),
        .dout(new_Jinkela_wire_13319)
    );

    spl2 new_Jinkela_splitter_969 (
        .a(new_Jinkela_wire_13192),
        .b(new_Jinkela_wire_13193),
        .c(new_Jinkela_wire_13194)
    );

    spl2 new_Jinkela_splitter_986 (
        .a(_0085_),
        .b(new_Jinkela_wire_13339),
        .c(new_Jinkela_wire_13340)
    );

    bfr new_Jinkela_buffer_10971 (
        .din(new_Jinkela_wire_13226),
        .dout(new_Jinkela_wire_13227)
    );

    bfr new_Jinkela_buffer_10972 (
        .din(new_Jinkela_wire_13227),
        .dout(new_Jinkela_wire_13228)
    );

    bfr new_Jinkela_buffer_11052 (
        .din(new_Jinkela_wire_13319),
        .dout(new_Jinkela_wire_13320)
    );

    bfr new_Jinkela_buffer_10973 (
        .din(new_Jinkela_wire_13228),
        .dout(new_Jinkela_wire_13229)
    );

    spl2 new_Jinkela_splitter_985 (
        .a(_0038_),
        .b(new_Jinkela_wire_13333),
        .c(new_Jinkela_wire_13334)
    );

    bfr new_Jinkela_buffer_10974 (
        .din(new_Jinkela_wire_13229),
        .dout(new_Jinkela_wire_13230)
    );

    bfr new_Jinkela_buffer_11053 (
        .din(new_Jinkela_wire_13320),
        .dout(new_Jinkela_wire_13321)
    );

    bfr new_Jinkela_buffer_10975 (
        .din(new_Jinkela_wire_13230),
        .dout(new_Jinkela_wire_13231)
    );

    bfr new_Jinkela_buffer_11056 (
        .din(new_Jinkela_wire_13325),
        .dout(new_Jinkela_wire_13326)
    );

    bfr new_Jinkela_buffer_10976 (
        .din(new_Jinkela_wire_13231),
        .dout(new_Jinkela_wire_13232)
    );

    bfr new_Jinkela_buffer_11061 (
        .din(new_Jinkela_wire_13334),
        .dout(new_Jinkela_wire_13335)
    );

    bfr new_Jinkela_buffer_10977 (
        .din(new_Jinkela_wire_13232),
        .dout(new_Jinkela_wire_13233)
    );

    bfr new_Jinkela_buffer_11057 (
        .din(new_Jinkela_wire_13326),
        .dout(new_Jinkela_wire_13327)
    );

    bfr new_Jinkela_buffer_10978 (
        .din(new_Jinkela_wire_13233),
        .dout(new_Jinkela_wire_13234)
    );

    bfr new_Jinkela_buffer_7425 (
        .din(new_Jinkela_wire_9240),
        .dout(new_Jinkela_wire_9241)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_1152),
        .dout(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    bfr new_Jinkela_buffer_7508 (
        .din(new_Jinkela_wire_9325),
        .dout(new_Jinkela_wire_9326)
    );

    bfr new_Jinkela_buffer_7426 (
        .din(new_Jinkela_wire_9241),
        .dout(new_Jinkela_wire_9242)
    );

    spl2 new_Jinkela_splitter_213 (
        .a(_1783_),
        .b(new_Jinkela_wire_1283),
        .c(new_Jinkela_wire_1284)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_7622 (
        .din(new_Jinkela_wire_9449),
        .dout(new_Jinkela_wire_9450)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_1277),
        .dout(new_Jinkela_wire_1278)
    );

    bfr new_Jinkela_buffer_7427 (
        .din(new_Jinkela_wire_9242),
        .dout(new_Jinkela_wire_9243)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_1153),
        .dout(new_Jinkela_wire_1154)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_1109),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_7509 (
        .din(new_Jinkela_wire_9326),
        .dout(new_Jinkela_wire_9327)
    );

    bfr new_Jinkela_buffer_7428 (
        .din(new_Jinkela_wire_9243),
        .dout(new_Jinkela_wire_9244)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_1271),
        .dout(new_Jinkela_wire_1272)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_7546 (
        .din(new_Jinkela_wire_9369),
        .dout(new_Jinkela_wire_9370)
    );

    bfr new_Jinkela_buffer_7429 (
        .din(new_Jinkela_wire_9244),
        .dout(new_Jinkela_wire_9245)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_1154),
        .dout(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    bfr new_Jinkela_buffer_7510 (
        .din(new_Jinkela_wire_9327),
        .dout(new_Jinkela_wire_9328)
    );

    bfr new_Jinkela_buffer_7430 (
        .din(new_Jinkela_wire_9245),
        .dout(new_Jinkela_wire_9246)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_7547 (
        .din(new_Jinkela_wire_9370),
        .dout(new_Jinkela_wire_9371)
    );

    spl2 new_Jinkela_splitter_212 (
        .a(_1531_),
        .b(new_Jinkela_wire_1281),
        .c(new_Jinkela_wire_1282)
    );

    bfr new_Jinkela_buffer_7431 (
        .din(new_Jinkela_wire_9246),
        .dout(new_Jinkela_wire_9247)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_1155),
        .dout(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_7511 (
        .din(new_Jinkela_wire_9328),
        .dout(new_Jinkela_wire_9329)
    );

    bfr new_Jinkela_buffer_7432 (
        .din(new_Jinkela_wire_9247),
        .dout(new_Jinkela_wire_9248)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_1272),
        .dout(new_Jinkela_wire_1273)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_7691 (
        .din(_1080_),
        .dout(new_Jinkela_wire_9523)
    );

    bfr new_Jinkela_buffer_7433 (
        .din(new_Jinkela_wire_9248),
        .dout(new_Jinkela_wire_9249)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_1156),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    bfr new_Jinkela_buffer_7512 (
        .din(new_Jinkela_wire_9329),
        .dout(new_Jinkela_wire_9330)
    );

    bfr new_Jinkela_buffer_7434 (
        .din(new_Jinkela_wire_9249),
        .dout(new_Jinkela_wire_9250)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_1116),
        .dout(new_Jinkela_wire_1117)
    );

    bfr new_Jinkela_buffer_7548 (
        .din(new_Jinkela_wire_9371),
        .dout(new_Jinkela_wire_9372)
    );

    bfr new_Jinkela_buffer_556 (
        .din(_0982_),
        .dout(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_7435 (
        .din(new_Jinkela_wire_9250),
        .dout(new_Jinkela_wire_9251)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_7513 (
        .din(new_Jinkela_wire_9330),
        .dout(new_Jinkela_wire_9331)
    );

    bfr new_Jinkela_buffer_7436 (
        .din(new_Jinkela_wire_9251),
        .dout(new_Jinkela_wire_9252)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_1273),
        .dout(new_Jinkela_wire_1274)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    bfr new_Jinkela_buffer_7623 (
        .din(new_Jinkela_wire_9450),
        .dout(new_Jinkela_wire_9451)
    );

    bfr new_Jinkela_buffer_7437 (
        .din(new_Jinkela_wire_9252),
        .dout(new_Jinkela_wire_9253)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    bfr new_Jinkela_buffer_7514 (
        .din(new_Jinkela_wire_9331),
        .dout(new_Jinkela_wire_9332)
    );

    bfr new_Jinkela_buffer_7438 (
        .din(new_Jinkela_wire_9253),
        .dout(new_Jinkela_wire_9254)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_7549 (
        .din(new_Jinkela_wire_9372),
        .dout(new_Jinkela_wire_9373)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_1278),
        .dout(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_7439 (
        .din(new_Jinkela_wire_9254),
        .dout(new_Jinkela_wire_9255)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_1159),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    bfr new_Jinkela_buffer_7515 (
        .din(new_Jinkela_wire_9332),
        .dout(new_Jinkela_wire_9333)
    );

    bfr new_Jinkela_buffer_7440 (
        .din(new_Jinkela_wire_9255),
        .dout(new_Jinkela_wire_9256)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_1122),
        .dout(new_Jinkela_wire_1123)
    );

    bfr new_Jinkela_buffer_7684 (
        .din(new_Jinkela_wire_9511),
        .dout(new_Jinkela_wire_9512)
    );

    bfr new_Jinkela_buffer_7441 (
        .din(new_Jinkela_wire_9256),
        .dout(new_Jinkela_wire_9257)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_1123),
        .dout(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_7516 (
        .din(new_Jinkela_wire_9333),
        .dout(new_Jinkela_wire_9334)
    );

    bfr new_Jinkela_buffer_7442 (
        .din(new_Jinkela_wire_9257),
        .dout(new_Jinkela_wire_9258)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    bfr new_Jinkela_buffer_7550 (
        .din(new_Jinkela_wire_9373),
        .dout(new_Jinkela_wire_9374)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_1279),
        .dout(new_Jinkela_wire_1280)
    );

    bfr new_Jinkela_buffer_7443 (
        .din(new_Jinkela_wire_9258),
        .dout(new_Jinkela_wire_9259)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    bfr new_Jinkela_buffer_7517 (
        .din(new_Jinkela_wire_9334),
        .dout(new_Jinkela_wire_9335)
    );

    bfr new_Jinkela_buffer_7444 (
        .din(new_Jinkela_wire_9259),
        .dout(new_Jinkela_wire_9260)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_1126),
        .dout(new_Jinkela_wire_1127)
    );

    bfr new_Jinkela_buffer_7624 (
        .din(new_Jinkela_wire_9451),
        .dout(new_Jinkela_wire_9452)
    );

    bfr new_Jinkela_buffer_555 (
        .din(_0044_),
        .dout(new_Jinkela_wire_1285)
    );

    bfr new_Jinkela_buffer_7445 (
        .din(new_Jinkela_wire_9260),
        .dout(new_Jinkela_wire_9261)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_1127),
        .dout(new_Jinkela_wire_1128)
    );

    bfr new_Jinkela_buffer_7518 (
        .din(new_Jinkela_wire_9335),
        .dout(new_Jinkela_wire_9336)
    );

    bfr new_Jinkela_buffer_4050 (
        .din(new_Jinkela_wire_5323),
        .dout(new_Jinkela_wire_5324)
    );

    bfr new_Jinkela_buffer_3979 (
        .din(new_Jinkela_wire_5246),
        .dout(new_Jinkela_wire_5247)
    );

    bfr new_Jinkela_buffer_4071 (
        .din(new_Jinkela_wire_5346),
        .dout(new_Jinkela_wire_5347)
    );

    bfr new_Jinkela_buffer_3980 (
        .din(new_Jinkela_wire_5247),
        .dout(new_Jinkela_wire_5248)
    );

    bfr new_Jinkela_buffer_4051 (
        .din(new_Jinkela_wire_5324),
        .dout(new_Jinkela_wire_5325)
    );

    bfr new_Jinkela_buffer_3981 (
        .din(new_Jinkela_wire_5248),
        .dout(new_Jinkela_wire_5249)
    );

    spl2 new_Jinkela_splitter_500 (
        .a(_1044_),
        .b(new_Jinkela_wire_5454),
        .c(new_Jinkela_wire_5455)
    );

    bfr new_Jinkela_buffer_4148 (
        .din(new_Jinkela_wire_5449),
        .dout(new_Jinkela_wire_5450)
    );

    bfr new_Jinkela_buffer_3982 (
        .din(new_Jinkela_wire_5249),
        .dout(new_Jinkela_wire_5250)
    );

    spl2 new_Jinkela_splitter_486 (
        .a(new_Jinkela_wire_5325),
        .b(new_Jinkela_wire_5326),
        .c(new_Jinkela_wire_5327)
    );

    bfr new_Jinkela_buffer_3983 (
        .din(new_Jinkela_wire_5250),
        .dout(new_Jinkela_wire_5251)
    );

    bfr new_Jinkela_buffer_3984 (
        .din(new_Jinkela_wire_5251),
        .dout(new_Jinkela_wire_5252)
    );

    bfr new_Jinkela_buffer_4072 (
        .din(new_Jinkela_wire_5347),
        .dout(new_Jinkela_wire_5348)
    );

    bfr new_Jinkela_buffer_3985 (
        .din(new_Jinkela_wire_5252),
        .dout(new_Jinkela_wire_5253)
    );

    bfr new_Jinkela_buffer_4073 (
        .din(new_Jinkela_wire_5348),
        .dout(new_Jinkela_wire_5349)
    );

    bfr new_Jinkela_buffer_3986 (
        .din(new_Jinkela_wire_5253),
        .dout(new_Jinkela_wire_5254)
    );

    bfr new_Jinkela_buffer_4152 (
        .din(_0680_),
        .dout(new_Jinkela_wire_5456)
    );

    bfr new_Jinkela_buffer_3987 (
        .din(new_Jinkela_wire_5254),
        .dout(new_Jinkela_wire_5255)
    );

    bfr new_Jinkela_buffer_4074 (
        .din(new_Jinkela_wire_5349),
        .dout(new_Jinkela_wire_5350)
    );

    bfr new_Jinkela_buffer_3988 (
        .din(new_Jinkela_wire_5255),
        .dout(new_Jinkela_wire_5256)
    );

    bfr new_Jinkela_buffer_4153 (
        .din(new_Jinkela_wire_5458),
        .dout(new_Jinkela_wire_5459)
    );

    bfr new_Jinkela_buffer_3989 (
        .din(new_Jinkela_wire_5256),
        .dout(new_Jinkela_wire_5257)
    );

    bfr new_Jinkela_buffer_4075 (
        .din(new_Jinkela_wire_5350),
        .dout(new_Jinkela_wire_5351)
    );

    bfr new_Jinkela_buffer_3990 (
        .din(new_Jinkela_wire_5257),
        .dout(new_Jinkela_wire_5258)
    );

    bfr new_Jinkela_buffer_4149 (
        .din(new_Jinkela_wire_5450),
        .dout(new_Jinkela_wire_5451)
    );

    bfr new_Jinkela_buffer_3991 (
        .din(new_Jinkela_wire_5258),
        .dout(new_Jinkela_wire_5259)
    );

    bfr new_Jinkela_buffer_4076 (
        .din(new_Jinkela_wire_5351),
        .dout(new_Jinkela_wire_5352)
    );

    bfr new_Jinkela_buffer_3992 (
        .din(new_Jinkela_wire_5259),
        .dout(new_Jinkela_wire_5260)
    );

    spl2 new_Jinkela_splitter_502 (
        .a(_1768_),
        .b(new_Jinkela_wire_5463),
        .c(new_Jinkela_wire_5464)
    );

    spl2 new_Jinkela_splitter_501 (
        .a(_0012_),
        .b(new_Jinkela_wire_5457),
        .c(new_Jinkela_wire_5458)
    );

    bfr new_Jinkela_buffer_3993 (
        .din(new_Jinkela_wire_5260),
        .dout(new_Jinkela_wire_5261)
    );

    bfr new_Jinkela_buffer_4077 (
        .din(new_Jinkela_wire_5352),
        .dout(new_Jinkela_wire_5353)
    );

    bfr new_Jinkela_buffer_3994 (
        .din(new_Jinkela_wire_5261),
        .dout(new_Jinkela_wire_5262)
    );

    bfr new_Jinkela_buffer_4150 (
        .din(new_Jinkela_wire_5451),
        .dout(new_Jinkela_wire_5452)
    );

    bfr new_Jinkela_buffer_3995 (
        .din(new_Jinkela_wire_5262),
        .dout(new_Jinkela_wire_5263)
    );

    bfr new_Jinkela_buffer_4078 (
        .din(new_Jinkela_wire_5353),
        .dout(new_Jinkela_wire_5354)
    );

    bfr new_Jinkela_buffer_3996 (
        .din(new_Jinkela_wire_5263),
        .dout(new_Jinkela_wire_5264)
    );

    bfr new_Jinkela_buffer_3997 (
        .din(new_Jinkela_wire_5264),
        .dout(new_Jinkela_wire_5265)
    );

    bfr new_Jinkela_buffer_4079 (
        .din(new_Jinkela_wire_5354),
        .dout(new_Jinkela_wire_5355)
    );

    bfr new_Jinkela_buffer_3998 (
        .din(new_Jinkela_wire_5265),
        .dout(new_Jinkela_wire_5266)
    );

    bfr new_Jinkela_buffer_4151 (
        .din(new_Jinkela_wire_5452),
        .dout(new_Jinkela_wire_5453)
    );

    bfr new_Jinkela_buffer_3999 (
        .din(new_Jinkela_wire_5266),
        .dout(new_Jinkela_wire_5267)
    );

    bfr new_Jinkela_buffer_17794 (
        .din(new_Jinkela_wire_21226),
        .dout(new_Jinkela_wire_21227)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_1128),
        .dout(new_Jinkela_wire_1129)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(_0736_),
        .b(new_Jinkela_wire_1334),
        .c(new_Jinkela_wire_1335)
    );

    bfr new_Jinkela_buffer_17795 (
        .din(new_Jinkela_wire_21227),
        .dout(new_Jinkela_wire_21228)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_1163),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_1129),
        .dout(new_Jinkela_wire_1130)
    );

    bfr new_Jinkela_buffer_17894 (
        .din(new_Jinkela_wire_21330),
        .dout(new_Jinkela_wire_21331)
    );

    bfr new_Jinkela_buffer_17796 (
        .din(new_Jinkela_wire_21228),
        .dout(new_Jinkela_wire_21229)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(new_Jinkela_wire_1285),
        .b(new_Jinkela_wire_1286),
        .c(new_Jinkela_wire_1287)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_1130),
        .dout(new_Jinkela_wire_1131)
    );

    bfr new_Jinkela_buffer_17797 (
        .din(new_Jinkela_wire_21229),
        .dout(new_Jinkela_wire_21230)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_1164),
        .dout(new_Jinkela_wire_1165)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_1131),
        .dout(new_Jinkela_wire_1132)
    );

    bfr new_Jinkela_buffer_17798 (
        .din(new_Jinkela_wire_21230),
        .dout(new_Jinkela_wire_21231)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_1288),
        .dout(new_Jinkela_wire_1289)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_1132),
        .dout(new_Jinkela_wire_1133)
    );

    bfr new_Jinkela_buffer_17799 (
        .din(new_Jinkela_wire_21231),
        .dout(new_Jinkela_wire_21232)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_1165),
        .dout(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_600 (
        .din(_1286_),
        .dout(new_Jinkela_wire_1336)
    );

    bfr new_Jinkela_buffer_17800 (
        .din(new_Jinkela_wire_21232),
        .dout(new_Jinkela_wire_21233)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_1166),
        .dout(new_Jinkela_wire_1167)
    );

    spl2 new_Jinkela_splitter_219 (
        .a(_1664_),
        .b(new_Jinkela_wire_1389),
        .c(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_17801 (
        .din(new_Jinkela_wire_21233),
        .dout(new_Jinkela_wire_21234)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_1167),
        .dout(new_Jinkela_wire_1168)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_1289),
        .dout(new_Jinkela_wire_1290)
    );

    bfr new_Jinkela_buffer_17802 (
        .din(new_Jinkela_wire_21234),
        .dout(new_Jinkela_wire_21235)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_1168),
        .dout(new_Jinkela_wire_1169)
    );

    spl2 new_Jinkela_splitter_218 (
        .a(_1775_),
        .b(new_Jinkela_wire_1387),
        .c(new_Jinkela_wire_1388)
    );

    bfr new_Jinkela_buffer_17803 (
        .din(new_Jinkela_wire_21235),
        .dout(new_Jinkela_wire_21236)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_1169),
        .dout(new_Jinkela_wire_1170)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_1290),
        .dout(new_Jinkela_wire_1291)
    );

    bfr new_Jinkela_buffer_17804 (
        .din(new_Jinkela_wire_21236),
        .dout(new_Jinkela_wire_21237)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_1170),
        .dout(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_1336),
        .dout(new_Jinkela_wire_1337)
    );

    bfr new_Jinkela_buffer_17805 (
        .din(new_Jinkela_wire_21237),
        .dout(new_Jinkela_wire_21238)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_1171),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_1291),
        .dout(new_Jinkela_wire_1292)
    );

    bfr new_Jinkela_buffer_17806 (
        .din(new_Jinkela_wire_21238),
        .dout(new_Jinkela_wire_21239)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_1172),
        .dout(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_17807 (
        .din(new_Jinkela_wire_21239),
        .dout(new_Jinkela_wire_21240)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_1173),
        .dout(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_1292),
        .dout(new_Jinkela_wire_1293)
    );

    bfr new_Jinkela_buffer_17808 (
        .din(new_Jinkela_wire_21240),
        .dout(new_Jinkela_wire_21241)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_1174),
        .dout(new_Jinkela_wire_1175)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_1337),
        .dout(new_Jinkela_wire_1338)
    );

    bfr new_Jinkela_buffer_17809 (
        .din(new_Jinkela_wire_21241),
        .dout(new_Jinkela_wire_21242)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_1175),
        .dout(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_1293),
        .dout(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_17810 (
        .din(new_Jinkela_wire_21242),
        .dout(new_Jinkela_wire_21243)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_1176),
        .dout(new_Jinkela_wire_1177)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(_1598_),
        .b(new_Jinkela_wire_1391),
        .c(new_Jinkela_wire_1392)
    );

    bfr new_Jinkela_buffer_17811 (
        .din(new_Jinkela_wire_21243),
        .dout(new_Jinkela_wire_21244)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_1177),
        .dout(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_1294),
        .dout(new_Jinkela_wire_1295)
    );

    bfr new_Jinkela_buffer_17812 (
        .din(new_Jinkela_wire_21244),
        .dout(new_Jinkela_wire_21245)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_1178),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_1338),
        .dout(new_Jinkela_wire_1339)
    );

    bfr new_Jinkela_buffer_17813 (
        .din(new_Jinkela_wire_21245),
        .dout(new_Jinkela_wire_21246)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_1179),
        .dout(new_Jinkela_wire_1180)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_1295),
        .dout(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_17814 (
        .din(new_Jinkela_wire_21246),
        .dout(new_Jinkela_wire_21247)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_net_3972),
        .dout(new_Jinkela_wire_1393)
    );

    bfr new_Jinkela_buffer_16950 (
        .din(new_Jinkela_wire_20202),
        .dout(new_Jinkela_wire_20203)
    );

    spl2 new_Jinkela_splitter_1493 (
        .a(_0263_),
        .b(new_Jinkela_wire_20324),
        .c(new_Jinkela_wire_20325)
    );

    bfr new_Jinkela_buffer_16951 (
        .din(new_Jinkela_wire_20203),
        .dout(new_Jinkela_wire_20204)
    );

    bfr new_Jinkela_buffer_16987 (
        .din(new_Jinkela_wire_20245),
        .dout(new_Jinkela_wire_20246)
    );

    bfr new_Jinkela_buffer_16952 (
        .din(new_Jinkela_wire_20204),
        .dout(new_Jinkela_wire_20205)
    );

    spl2 new_Jinkela_splitter_1490 (
        .a(new_Jinkela_wire_20292),
        .b(new_Jinkela_wire_20293),
        .c(new_Jinkela_wire_20294)
    );

    bfr new_Jinkela_buffer_16953 (
        .din(new_Jinkela_wire_20205),
        .dout(new_Jinkela_wire_20206)
    );

    bfr new_Jinkela_buffer_16988 (
        .din(new_Jinkela_wire_20246),
        .dout(new_Jinkela_wire_20247)
    );

    bfr new_Jinkela_buffer_16954 (
        .din(new_Jinkela_wire_20206),
        .dout(new_Jinkela_wire_20207)
    );

    spl2 new_Jinkela_splitter_1475 (
        .a(new_Jinkela_wire_20207),
        .b(new_Jinkela_wire_20208),
        .c(new_Jinkela_wire_20209)
    );

    bfr new_Jinkela_buffer_17012 (
        .din(new_Jinkela_wire_20296),
        .dout(new_Jinkela_wire_20297)
    );

    bfr new_Jinkela_buffer_16989 (
        .din(new_Jinkela_wire_20247),
        .dout(new_Jinkela_wire_20248)
    );

    bfr new_Jinkela_buffer_16990 (
        .din(new_Jinkela_wire_20248),
        .dout(new_Jinkela_wire_20249)
    );

    bfr new_Jinkela_buffer_17013 (
        .din(new_Jinkela_wire_20297),
        .dout(new_Jinkela_wire_20298)
    );

    bfr new_Jinkela_buffer_16991 (
        .din(new_Jinkela_wire_20249),
        .dout(new_Jinkela_wire_20250)
    );

    spl2 new_Jinkela_splitter_1494 (
        .a(_1066_),
        .b(new_Jinkela_wire_20326),
        .c(new_Jinkela_wire_20327)
    );

    bfr new_Jinkela_buffer_16992 (
        .din(new_Jinkela_wire_20250),
        .dout(new_Jinkela_wire_20251)
    );

    bfr new_Jinkela_buffer_17014 (
        .din(new_Jinkela_wire_20298),
        .dout(new_Jinkela_wire_20299)
    );

    bfr new_Jinkela_buffer_16993 (
        .din(new_Jinkela_wire_20251),
        .dout(new_Jinkela_wire_20252)
    );

    bfr new_Jinkela_buffer_17039 (
        .din(_0065_),
        .dout(new_Jinkela_wire_20332)
    );

    bfr new_Jinkela_buffer_16994 (
        .din(new_Jinkela_wire_20252),
        .dout(new_Jinkela_wire_20253)
    );

    bfr new_Jinkela_buffer_17015 (
        .din(new_Jinkela_wire_20299),
        .dout(new_Jinkela_wire_20300)
    );

    bfr new_Jinkela_buffer_16995 (
        .din(new_Jinkela_wire_20253),
        .dout(new_Jinkela_wire_20254)
    );

    bfr new_Jinkela_buffer_17035 (
        .din(new_Jinkela_wire_20327),
        .dout(new_Jinkela_wire_20328)
    );

    spl2 new_Jinkela_splitter_1495 (
        .a(_1100_),
        .b(new_Jinkela_wire_20333),
        .c(new_Jinkela_wire_20334)
    );

    bfr new_Jinkela_buffer_16996 (
        .din(new_Jinkela_wire_20254),
        .dout(new_Jinkela_wire_20255)
    );

    bfr new_Jinkela_buffer_17016 (
        .din(new_Jinkela_wire_20300),
        .dout(new_Jinkela_wire_20301)
    );

    bfr new_Jinkela_buffer_16997 (
        .din(new_Jinkela_wire_20255),
        .dout(new_Jinkela_wire_20256)
    );

    bfr new_Jinkela_buffer_17044 (
        .din(_1418_),
        .dout(new_Jinkela_wire_20339)
    );

    bfr new_Jinkela_buffer_17040 (
        .din(new_Jinkela_wire_20334),
        .dout(new_Jinkela_wire_20335)
    );

    bfr new_Jinkela_buffer_16998 (
        .din(new_Jinkela_wire_20256),
        .dout(new_Jinkela_wire_20257)
    );

    bfr new_Jinkela_buffer_17017 (
        .din(new_Jinkela_wire_20301),
        .dout(new_Jinkela_wire_20302)
    );

    spl2 new_Jinkela_splitter_1478 (
        .a(new_Jinkela_wire_20257),
        .b(new_Jinkela_wire_20258),
        .c(new_Jinkela_wire_20259)
    );

    bfr new_Jinkela_buffer_17018 (
        .din(new_Jinkela_wire_20302),
        .dout(new_Jinkela_wire_20303)
    );

    bfr new_Jinkela_buffer_17036 (
        .din(new_Jinkela_wire_20328),
        .dout(new_Jinkela_wire_20329)
    );

    bfr new_Jinkela_buffer_17019 (
        .din(new_Jinkela_wire_20303),
        .dout(new_Jinkela_wire_20304)
    );

    bfr new_Jinkela_buffer_17037 (
        .din(new_Jinkela_wire_20329),
        .dout(new_Jinkela_wire_20330)
    );

    bfr new_Jinkela_buffer_17020 (
        .din(new_Jinkela_wire_20304),
        .dout(new_Jinkela_wire_20305)
    );

    spl2 new_Jinkela_splitter_1496 (
        .a(_1042_),
        .b(new_Jinkela_wire_20340),
        .c(new_Jinkela_wire_20341)
    );

    bfr new_Jinkela_buffer_17021 (
        .din(new_Jinkela_wire_20305),
        .dout(new_Jinkela_wire_20306)
    );

    bfr new_Jinkela_buffer_17038 (
        .din(new_Jinkela_wire_20330),
        .dout(new_Jinkela_wire_20331)
    );

    bfr new_Jinkela_buffer_17022 (
        .din(new_Jinkela_wire_20306),
        .dout(new_Jinkela_wire_20307)
    );

    spl2 new_Jinkela_splitter_935 (
        .a(_0803_),
        .b(new_Jinkela_wire_12622),
        .c(new_Jinkela_wire_12623)
    );

    bfr new_Jinkela_buffer_10100 (
        .din(new_Jinkela_wire_12249),
        .dout(new_Jinkela_wire_12250)
    );

    bfr new_Jinkela_buffer_10189 (
        .din(new_Jinkela_wire_12352),
        .dout(new_Jinkela_wire_12353)
    );

    bfr new_Jinkela_buffer_10101 (
        .din(new_Jinkela_wire_12250),
        .dout(new_Jinkela_wire_12251)
    );

    bfr new_Jinkela_buffer_10360 (
        .din(new_Jinkela_wire_12527),
        .dout(new_Jinkela_wire_12528)
    );

    bfr new_Jinkela_buffer_10102 (
        .din(new_Jinkela_wire_12251),
        .dout(new_Jinkela_wire_12252)
    );

    bfr new_Jinkela_buffer_10190 (
        .din(new_Jinkela_wire_12353),
        .dout(new_Jinkela_wire_12354)
    );

    bfr new_Jinkela_buffer_10103 (
        .din(new_Jinkela_wire_12252),
        .dout(new_Jinkela_wire_12253)
    );

    bfr new_Jinkela_buffer_10450 (
        .din(_0013_),
        .dout(new_Jinkela_wire_12624)
    );

    spl2 new_Jinkela_splitter_937 (
        .a(_0163_),
        .b(new_Jinkela_wire_12627),
        .c(new_Jinkela_wire_12628)
    );

    bfr new_Jinkela_buffer_10104 (
        .din(new_Jinkela_wire_12253),
        .dout(new_Jinkela_wire_12254)
    );

    bfr new_Jinkela_buffer_10191 (
        .din(new_Jinkela_wire_12354),
        .dout(new_Jinkela_wire_12355)
    );

    bfr new_Jinkela_buffer_10105 (
        .din(new_Jinkela_wire_12254),
        .dout(new_Jinkela_wire_12255)
    );

    bfr new_Jinkela_buffer_10361 (
        .din(new_Jinkela_wire_12528),
        .dout(new_Jinkela_wire_12529)
    );

    bfr new_Jinkela_buffer_10106 (
        .din(new_Jinkela_wire_12255),
        .dout(new_Jinkela_wire_12256)
    );

    bfr new_Jinkela_buffer_10192 (
        .din(new_Jinkela_wire_12355),
        .dout(new_Jinkela_wire_12356)
    );

    bfr new_Jinkela_buffer_10107 (
        .din(new_Jinkela_wire_12256),
        .dout(new_Jinkela_wire_12257)
    );

    bfr new_Jinkela_buffer_10446 (
        .din(new_Jinkela_wire_12617),
        .dout(new_Jinkela_wire_12618)
    );

    bfr new_Jinkela_buffer_10108 (
        .din(new_Jinkela_wire_12257),
        .dout(new_Jinkela_wire_12258)
    );

    bfr new_Jinkela_buffer_10193 (
        .din(new_Jinkela_wire_12356),
        .dout(new_Jinkela_wire_12357)
    );

    bfr new_Jinkela_buffer_10109 (
        .din(new_Jinkela_wire_12258),
        .dout(new_Jinkela_wire_12259)
    );

    bfr new_Jinkela_buffer_10362 (
        .din(new_Jinkela_wire_12529),
        .dout(new_Jinkela_wire_12530)
    );

    bfr new_Jinkela_buffer_10110 (
        .din(new_Jinkela_wire_12259),
        .dout(new_Jinkela_wire_12260)
    );

    bfr new_Jinkela_buffer_10194 (
        .din(new_Jinkela_wire_12357),
        .dout(new_Jinkela_wire_12358)
    );

    bfr new_Jinkela_buffer_10111 (
        .din(new_Jinkela_wire_12260),
        .dout(new_Jinkela_wire_12261)
    );

    bfr new_Jinkela_buffer_10112 (
        .din(new_Jinkela_wire_12261),
        .dout(new_Jinkela_wire_12262)
    );

    bfr new_Jinkela_buffer_10195 (
        .din(new_Jinkela_wire_12358),
        .dout(new_Jinkela_wire_12359)
    );

    bfr new_Jinkela_buffer_10113 (
        .din(new_Jinkela_wire_12262),
        .dout(new_Jinkela_wire_12263)
    );

    bfr new_Jinkela_buffer_10363 (
        .din(new_Jinkela_wire_12530),
        .dout(new_Jinkela_wire_12531)
    );

    bfr new_Jinkela_buffer_10114 (
        .din(new_Jinkela_wire_12263),
        .dout(new_Jinkela_wire_12264)
    );

    bfr new_Jinkela_buffer_10196 (
        .din(new_Jinkela_wire_12359),
        .dout(new_Jinkela_wire_12360)
    );

    bfr new_Jinkela_buffer_10115 (
        .din(new_Jinkela_wire_12264),
        .dout(new_Jinkela_wire_12265)
    );

    bfr new_Jinkela_buffer_10447 (
        .din(new_Jinkela_wire_12618),
        .dout(new_Jinkela_wire_12619)
    );

    bfr new_Jinkela_buffer_10116 (
        .din(new_Jinkela_wire_12265),
        .dout(new_Jinkela_wire_12266)
    );

    bfr new_Jinkela_buffer_10197 (
        .din(new_Jinkela_wire_12360),
        .dout(new_Jinkela_wire_12361)
    );

    bfr new_Jinkela_buffer_10117 (
        .din(new_Jinkela_wire_12266),
        .dout(new_Jinkela_wire_12267)
    );

    bfr new_Jinkela_buffer_10364 (
        .din(new_Jinkela_wire_12531),
        .dout(new_Jinkela_wire_12532)
    );

    bfr new_Jinkela_buffer_10118 (
        .din(new_Jinkela_wire_12267),
        .dout(new_Jinkela_wire_12268)
    );

    bfr new_Jinkela_buffer_10198 (
        .din(new_Jinkela_wire_12361),
        .dout(new_Jinkela_wire_12362)
    );

    bfr new_Jinkela_buffer_10119 (
        .din(new_Jinkela_wire_12268),
        .dout(new_Jinkela_wire_12269)
    );

    spl2 new_Jinkela_splitter_936 (
        .a(_0017_),
        .b(new_Jinkela_wire_12625),
        .c(new_Jinkela_wire_12626)
    );

    bfr new_Jinkela_buffer_10120 (
        .din(new_Jinkela_wire_12269),
        .dout(new_Jinkela_wire_12270)
    );

    bfr new_Jinkela_buffer_3197 (
        .din(new_Jinkela_wire_4314),
        .dout(new_Jinkela_wire_4315)
    );

    bfr new_Jinkela_buffer_3198 (
        .din(new_Jinkela_wire_4315),
        .dout(new_Jinkela_wire_4316)
    );

    bfr new_Jinkela_buffer_3211 (
        .din(new_Jinkela_wire_4332),
        .dout(new_Jinkela_wire_4333)
    );

    bfr new_Jinkela_buffer_3199 (
        .din(new_Jinkela_wire_4316),
        .dout(new_Jinkela_wire_4317)
    );

    spl2 new_Jinkela_splitter_412 (
        .a(_1285_),
        .b(new_Jinkela_wire_4475),
        .c(new_Jinkela_wire_4476)
    );

    bfr new_Jinkela_buffer_3200 (
        .din(new_Jinkela_wire_4317),
        .dout(new_Jinkela_wire_4318)
    );

    bfr new_Jinkela_buffer_3342 (
        .din(new_Jinkela_wire_4463),
        .dout(new_Jinkela_wire_4464)
    );

    bfr new_Jinkela_buffer_3212 (
        .din(new_Jinkela_wire_4333),
        .dout(new_Jinkela_wire_4334)
    );

    bfr new_Jinkela_buffer_3201 (
        .din(new_Jinkela_wire_4318),
        .dout(new_Jinkela_wire_4319)
    );

    bfr new_Jinkela_buffer_3202 (
        .din(new_Jinkela_wire_4319),
        .dout(new_Jinkela_wire_4320)
    );

    bfr new_Jinkela_buffer_3213 (
        .din(new_Jinkela_wire_4334),
        .dout(new_Jinkela_wire_4335)
    );

    bfr new_Jinkela_buffer_3343 (
        .din(new_Jinkela_wire_4464),
        .dout(new_Jinkela_wire_4465)
    );

    bfr new_Jinkela_buffer_3214 (
        .din(new_Jinkela_wire_4335),
        .dout(new_Jinkela_wire_4336)
    );

    bfr new_Jinkela_buffer_3215 (
        .din(new_Jinkela_wire_4336),
        .dout(new_Jinkela_wire_4337)
    );

    spl2 new_Jinkela_splitter_413 (
        .a(_0576_),
        .b(new_Jinkela_wire_4477),
        .c(new_Jinkela_wire_4478)
    );

    bfr new_Jinkela_buffer_3344 (
        .din(new_Jinkela_wire_4465),
        .dout(new_Jinkela_wire_4466)
    );

    bfr new_Jinkela_buffer_3216 (
        .din(new_Jinkela_wire_4337),
        .dout(new_Jinkela_wire_4338)
    );

    bfr new_Jinkela_buffer_3217 (
        .din(new_Jinkela_wire_4338),
        .dout(new_Jinkela_wire_4339)
    );

    bfr new_Jinkela_buffer_3353 (
        .din(_0647_),
        .dout(new_Jinkela_wire_4483)
    );

    bfr new_Jinkela_buffer_3345 (
        .din(new_Jinkela_wire_4466),
        .dout(new_Jinkela_wire_4467)
    );

    bfr new_Jinkela_buffer_3218 (
        .din(new_Jinkela_wire_4339),
        .dout(new_Jinkela_wire_4340)
    );

    bfr new_Jinkela_buffer_3349 (
        .din(new_Jinkela_wire_4478),
        .dout(new_Jinkela_wire_4479)
    );

    bfr new_Jinkela_buffer_3219 (
        .din(new_Jinkela_wire_4340),
        .dout(new_Jinkela_wire_4341)
    );

    bfr new_Jinkela_buffer_3354 (
        .din(_1324_),
        .dout(new_Jinkela_wire_4484)
    );

    bfr new_Jinkela_buffer_3346 (
        .din(new_Jinkela_wire_4467),
        .dout(new_Jinkela_wire_4468)
    );

    bfr new_Jinkela_buffer_3220 (
        .din(new_Jinkela_wire_4341),
        .dout(new_Jinkela_wire_4342)
    );

    bfr new_Jinkela_buffer_3221 (
        .din(new_Jinkela_wire_4342),
        .dout(new_Jinkela_wire_4343)
    );

    bfr new_Jinkela_buffer_3355 (
        .din(_0128_),
        .dout(new_Jinkela_wire_4485)
    );

    bfr new_Jinkela_buffer_3347 (
        .din(new_Jinkela_wire_4468),
        .dout(new_Jinkela_wire_4469)
    );

    bfr new_Jinkela_buffer_3222 (
        .din(new_Jinkela_wire_4343),
        .dout(new_Jinkela_wire_4344)
    );

    bfr new_Jinkela_buffer_3350 (
        .din(new_Jinkela_wire_4479),
        .dout(new_Jinkela_wire_4480)
    );

    bfr new_Jinkela_buffer_3223 (
        .din(new_Jinkela_wire_4344),
        .dout(new_Jinkela_wire_4345)
    );

    bfr new_Jinkela_buffer_3348 (
        .din(new_Jinkela_wire_4469),
        .dout(new_Jinkela_wire_4470)
    );

    bfr new_Jinkela_buffer_3224 (
        .din(new_Jinkela_wire_4345),
        .dout(new_Jinkela_wire_4346)
    );

    bfr new_Jinkela_buffer_3225 (
        .din(new_Jinkela_wire_4346),
        .dout(new_Jinkela_wire_4347)
    );

    bfr new_Jinkela_buffer_3356 (
        .din(new_net_3936),
        .dout(new_Jinkela_wire_4486)
    );

    spl2 new_Jinkela_splitter_410 (
        .a(new_Jinkela_wire_4470),
        .b(new_Jinkela_wire_4471),
        .c(new_Jinkela_wire_4472)
    );

    bfr new_Jinkela_buffer_3226 (
        .din(new_Jinkela_wire_4347),
        .dout(new_Jinkela_wire_4348)
    );

    bfr new_Jinkela_buffer_3227 (
        .din(new_Jinkela_wire_4348),
        .dout(new_Jinkela_wire_4349)
    );

    bfr new_Jinkela_buffer_3351 (
        .din(new_Jinkela_wire_4480),
        .dout(new_Jinkela_wire_4481)
    );

    bfr new_Jinkela_buffer_3228 (
        .din(new_Jinkela_wire_4349),
        .dout(new_Jinkela_wire_4350)
    );

    bfr new_Jinkela_buffer_6613 (
        .din(new_Jinkela_wire_8332),
        .dout(new_Jinkela_wire_8333)
    );

    bfr new_Jinkela_buffer_6655 (
        .din(new_Jinkela_wire_8378),
        .dout(new_Jinkela_wire_8379)
    );

    bfr new_Jinkela_buffer_6614 (
        .din(new_Jinkela_wire_8333),
        .dout(new_Jinkela_wire_8334)
    );

    bfr new_Jinkela_buffer_6615 (
        .din(new_Jinkela_wire_8334),
        .dout(new_Jinkela_wire_8335)
    );

    bfr new_Jinkela_buffer_6656 (
        .din(new_Jinkela_wire_8379),
        .dout(new_Jinkela_wire_8380)
    );

    bfr new_Jinkela_buffer_6616 (
        .din(new_Jinkela_wire_8335),
        .dout(new_Jinkela_wire_8336)
    );

    bfr new_Jinkela_buffer_6744 (
        .din(new_Jinkela_wire_8469),
        .dout(new_Jinkela_wire_8470)
    );

    bfr new_Jinkela_buffer_6617 (
        .din(new_Jinkela_wire_8336),
        .dout(new_Jinkela_wire_8337)
    );

    bfr new_Jinkela_buffer_6657 (
        .din(new_Jinkela_wire_8380),
        .dout(new_Jinkela_wire_8381)
    );

    bfr new_Jinkela_buffer_6618 (
        .din(new_Jinkela_wire_8337),
        .dout(new_Jinkela_wire_8338)
    );

    bfr new_Jinkela_buffer_6755 (
        .din(new_Jinkela_wire_8486),
        .dout(new_Jinkela_wire_8487)
    );

    bfr new_Jinkela_buffer_6619 (
        .din(new_Jinkela_wire_8338),
        .dout(new_Jinkela_wire_8339)
    );

    bfr new_Jinkela_buffer_6658 (
        .din(new_Jinkela_wire_8381),
        .dout(new_Jinkela_wire_8382)
    );

    bfr new_Jinkela_buffer_6620 (
        .din(new_Jinkela_wire_8339),
        .dout(new_Jinkela_wire_8340)
    );

    bfr new_Jinkela_buffer_6745 (
        .din(new_Jinkela_wire_8470),
        .dout(new_Jinkela_wire_8471)
    );

    bfr new_Jinkela_buffer_6621 (
        .din(new_Jinkela_wire_8340),
        .dout(new_Jinkela_wire_8341)
    );

    bfr new_Jinkela_buffer_6659 (
        .din(new_Jinkela_wire_8382),
        .dout(new_Jinkela_wire_8383)
    );

    bfr new_Jinkela_buffer_6622 (
        .din(new_Jinkela_wire_8341),
        .dout(new_Jinkela_wire_8342)
    );

    spl2 new_Jinkela_splitter_719 (
        .a(_0243_),
        .b(new_Jinkela_wire_8586),
        .c(new_Jinkela_wire_8587)
    );

    bfr new_Jinkela_buffer_6623 (
        .din(new_Jinkela_wire_8342),
        .dout(new_Jinkela_wire_8343)
    );

    bfr new_Jinkela_buffer_6660 (
        .din(new_Jinkela_wire_8383),
        .dout(new_Jinkela_wire_8384)
    );

    bfr new_Jinkela_buffer_6624 (
        .din(new_Jinkela_wire_8343),
        .dout(new_Jinkela_wire_8344)
    );

    bfr new_Jinkela_buffer_6746 (
        .din(new_Jinkela_wire_8471),
        .dout(new_Jinkela_wire_8472)
    );

    bfr new_Jinkela_buffer_6625 (
        .din(new_Jinkela_wire_8344),
        .dout(new_Jinkela_wire_8345)
    );

    bfr new_Jinkela_buffer_6661 (
        .din(new_Jinkela_wire_8384),
        .dout(new_Jinkela_wire_8385)
    );

    bfr new_Jinkela_buffer_6626 (
        .din(new_Jinkela_wire_8345),
        .dout(new_Jinkela_wire_8346)
    );

    bfr new_Jinkela_buffer_6756 (
        .din(new_Jinkela_wire_8487),
        .dout(new_Jinkela_wire_8488)
    );

    bfr new_Jinkela_buffer_6627 (
        .din(new_Jinkela_wire_8346),
        .dout(new_Jinkela_wire_8347)
    );

    bfr new_Jinkela_buffer_6662 (
        .din(new_Jinkela_wire_8385),
        .dout(new_Jinkela_wire_8386)
    );

    bfr new_Jinkela_buffer_6628 (
        .din(new_Jinkela_wire_8347),
        .dout(new_Jinkela_wire_8348)
    );

    bfr new_Jinkela_buffer_6747 (
        .din(new_Jinkela_wire_8472),
        .dout(new_Jinkela_wire_8473)
    );

    bfr new_Jinkela_buffer_6629 (
        .din(new_Jinkela_wire_8348),
        .dout(new_Jinkela_wire_8349)
    );

    bfr new_Jinkela_buffer_6663 (
        .din(new_Jinkela_wire_8386),
        .dout(new_Jinkela_wire_8387)
    );

    bfr new_Jinkela_buffer_6630 (
        .din(new_Jinkela_wire_8349),
        .dout(new_Jinkela_wire_8350)
    );

    spl2 new_Jinkela_splitter_720 (
        .a(_0573_),
        .b(new_Jinkela_wire_8589),
        .c(new_Jinkela_wire_8590)
    );

    bfr new_Jinkela_buffer_6846 (
        .din(_1244_),
        .dout(new_Jinkela_wire_8588)
    );

    bfr new_Jinkela_buffer_6631 (
        .din(new_Jinkela_wire_8350),
        .dout(new_Jinkela_wire_8351)
    );

    bfr new_Jinkela_buffer_6664 (
        .din(new_Jinkela_wire_8387),
        .dout(new_Jinkela_wire_8388)
    );

    bfr new_Jinkela_buffer_6632 (
        .din(new_Jinkela_wire_8351),
        .dout(new_Jinkela_wire_8352)
    );

    bfr new_Jinkela_buffer_6748 (
        .din(new_Jinkela_wire_8473),
        .dout(new_Jinkela_wire_8474)
    );

    bfr new_Jinkela_buffer_6633 (
        .din(new_Jinkela_wire_8352),
        .dout(new_Jinkela_wire_8353)
    );

    bfr new_Jinkela_buffer_6665 (
        .din(new_Jinkela_wire_8388),
        .dout(new_Jinkela_wire_8389)
    );

    bfr new_Jinkela_buffer_10199 (
        .din(new_Jinkela_wire_12362),
        .dout(new_Jinkela_wire_12363)
    );

    bfr new_Jinkela_buffer_6634 (
        .din(new_Jinkela_wire_8353),
        .dout(new_Jinkela_wire_8354)
    );

    bfr new_Jinkela_buffer_13586 (
        .din(new_Jinkela_wire_16241),
        .dout(new_Jinkela_wire_16242)
    );

    bfr new_Jinkela_buffer_3408 (
        .din(_0878_),
        .dout(new_Jinkela_wire_4538)
    );

    bfr new_Jinkela_buffer_6757 (
        .din(new_Jinkela_wire_8488),
        .dout(new_Jinkela_wire_8489)
    );

    bfr new_Jinkela_buffer_3352 (
        .din(new_Jinkela_wire_4481),
        .dout(new_Jinkela_wire_4482)
    );

    bfr new_Jinkela_buffer_10121 (
        .din(new_Jinkela_wire_12270),
        .dout(new_Jinkela_wire_12271)
    );

    bfr new_Jinkela_buffer_3229 (
        .din(new_Jinkela_wire_4350),
        .dout(new_Jinkela_wire_4351)
    );

    bfr new_Jinkela_buffer_13720 (
        .din(new_Jinkela_wire_16381),
        .dout(new_Jinkela_wire_16382)
    );

    bfr new_Jinkela_buffer_10365 (
        .din(new_Jinkela_wire_12532),
        .dout(new_Jinkela_wire_12533)
    );

    bfr new_Jinkela_buffer_6635 (
        .din(new_Jinkela_wire_8354),
        .dout(new_Jinkela_wire_8355)
    );

    bfr new_Jinkela_buffer_13587 (
        .din(new_Jinkela_wire_16242),
        .dout(new_Jinkela_wire_16243)
    );

    bfr new_Jinkela_buffer_10122 (
        .din(new_Jinkela_wire_12271),
        .dout(new_Jinkela_wire_12272)
    );

    bfr new_Jinkela_buffer_6666 (
        .din(new_Jinkela_wire_8389),
        .dout(new_Jinkela_wire_8390)
    );

    bfr new_Jinkela_buffer_13688 (
        .din(new_Jinkela_wire_16345),
        .dout(new_Jinkela_wire_16346)
    );

    bfr new_Jinkela_buffer_3230 (
        .din(new_Jinkela_wire_4351),
        .dout(new_Jinkela_wire_4352)
    );

    bfr new_Jinkela_buffer_10200 (
        .din(new_Jinkela_wire_12363),
        .dout(new_Jinkela_wire_12364)
    );

    bfr new_Jinkela_buffer_6636 (
        .din(new_Jinkela_wire_8355),
        .dout(new_Jinkela_wire_8356)
    );

    bfr new_Jinkela_buffer_13588 (
        .din(new_Jinkela_wire_16243),
        .dout(new_Jinkela_wire_16244)
    );

    bfr new_Jinkela_buffer_3357 (
        .din(new_Jinkela_wire_4486),
        .dout(new_Jinkela_wire_4487)
    );

    bfr new_Jinkela_buffer_10123 (
        .din(new_Jinkela_wire_12272),
        .dout(new_Jinkela_wire_12273)
    );

    bfr new_Jinkela_buffer_6749 (
        .din(new_Jinkela_wire_8474),
        .dout(new_Jinkela_wire_8475)
    );

    bfr new_Jinkela_buffer_13715 (
        .din(new_Jinkela_wire_16374),
        .dout(new_Jinkela_wire_16375)
    );

    bfr new_Jinkela_buffer_3231 (
        .din(new_Jinkela_wire_4352),
        .dout(new_Jinkela_wire_4353)
    );

    bfr new_Jinkela_buffer_10448 (
        .din(new_Jinkela_wire_12619),
        .dout(new_Jinkela_wire_12620)
    );

    bfr new_Jinkela_buffer_6637 (
        .din(new_Jinkela_wire_8356),
        .dout(new_Jinkela_wire_8357)
    );

    bfr new_Jinkela_buffer_13589 (
        .din(new_Jinkela_wire_16244),
        .dout(new_Jinkela_wire_16245)
    );

    spl2 new_Jinkela_splitter_414 (
        .a(_0195_),
        .b(new_Jinkela_wire_4539),
        .c(new_Jinkela_wire_4540)
    );

    bfr new_Jinkela_buffer_6667 (
        .din(new_Jinkela_wire_8390),
        .dout(new_Jinkela_wire_8391)
    );

    spl2 new_Jinkela_splitter_415 (
        .a(_0624_),
        .b(new_Jinkela_wire_4541),
        .c(new_Jinkela_wire_4542)
    );

    bfr new_Jinkela_buffer_10124 (
        .din(new_Jinkela_wire_12273),
        .dout(new_Jinkela_wire_12274)
    );

    bfr new_Jinkela_buffer_3232 (
        .din(new_Jinkela_wire_4353),
        .dout(new_Jinkela_wire_4354)
    );

    bfr new_Jinkela_buffer_13689 (
        .din(new_Jinkela_wire_16346),
        .dout(new_Jinkela_wire_16347)
    );

    bfr new_Jinkela_buffer_10201 (
        .din(new_Jinkela_wire_12364),
        .dout(new_Jinkela_wire_12365)
    );

    bfr new_Jinkela_buffer_6638 (
        .din(new_Jinkela_wire_8357),
        .dout(new_Jinkela_wire_8358)
    );

    bfr new_Jinkela_buffer_13590 (
        .din(new_Jinkela_wire_16245),
        .dout(new_Jinkela_wire_16246)
    );

    bfr new_Jinkela_buffer_3358 (
        .din(new_Jinkela_wire_4487),
        .dout(new_Jinkela_wire_4488)
    );

    bfr new_Jinkela_buffer_10125 (
        .din(new_Jinkela_wire_12274),
        .dout(new_Jinkela_wire_12275)
    );

    bfr new_Jinkela_buffer_6847 (
        .din(_1809_),
        .dout(new_Jinkela_wire_8591)
    );

    bfr new_Jinkela_buffer_3233 (
        .din(new_Jinkela_wire_4354),
        .dout(new_Jinkela_wire_4355)
    );

    bfr new_Jinkela_buffer_13840 (
        .din(_0419_),
        .dout(new_Jinkela_wire_16508)
    );

    bfr new_Jinkela_buffer_10366 (
        .din(new_Jinkela_wire_12533),
        .dout(new_Jinkela_wire_12534)
    );

    spl2 new_Jinkela_splitter_709 (
        .a(new_Jinkela_wire_8358),
        .b(new_Jinkela_wire_8359),
        .c(new_Jinkela_wire_8360)
    );

    bfr new_Jinkela_buffer_13591 (
        .din(new_Jinkela_wire_16246),
        .dout(new_Jinkela_wire_16247)
    );

    bfr new_Jinkela_buffer_3433 (
        .din(_0623_),
        .dout(new_Jinkela_wire_4571)
    );

    bfr new_Jinkela_buffer_10126 (
        .din(new_Jinkela_wire_12275),
        .dout(new_Jinkela_wire_12276)
    );

    bfr new_Jinkela_buffer_6750 (
        .din(new_Jinkela_wire_8475),
        .dout(new_Jinkela_wire_8476)
    );

    bfr new_Jinkela_buffer_13690 (
        .din(new_Jinkela_wire_16347),
        .dout(new_Jinkela_wire_16348)
    );

    bfr new_Jinkela_buffer_3234 (
        .din(new_Jinkela_wire_4355),
        .dout(new_Jinkela_wire_4356)
    );

    bfr new_Jinkela_buffer_10202 (
        .din(new_Jinkela_wire_12365),
        .dout(new_Jinkela_wire_12366)
    );

    bfr new_Jinkela_buffer_6668 (
        .din(new_Jinkela_wire_8391),
        .dout(new_Jinkela_wire_8392)
    );

    bfr new_Jinkela_buffer_13592 (
        .din(new_Jinkela_wire_16247),
        .dout(new_Jinkela_wire_16248)
    );

    bfr new_Jinkela_buffer_3359 (
        .din(new_Jinkela_wire_4488),
        .dout(new_Jinkela_wire_4489)
    );

    bfr new_Jinkela_buffer_10127 (
        .din(new_Jinkela_wire_12276),
        .dout(new_Jinkela_wire_12277)
    );

    bfr new_Jinkela_buffer_6669 (
        .din(new_Jinkela_wire_8392),
        .dout(new_Jinkela_wire_8393)
    );

    bfr new_Jinkela_buffer_13716 (
        .din(new_Jinkela_wire_16375),
        .dout(new_Jinkela_wire_16376)
    );

    bfr new_Jinkela_buffer_3235 (
        .din(new_Jinkela_wire_4356),
        .dout(new_Jinkela_wire_4357)
    );

    spl2 new_Jinkela_splitter_940 (
        .a(_0199_),
        .b(new_Jinkela_wire_12713),
        .c(new_Jinkela_wire_12714)
    );

    bfr new_Jinkela_buffer_6758 (
        .din(new_Jinkela_wire_8489),
        .dout(new_Jinkela_wire_8490)
    );

    bfr new_Jinkela_buffer_13593 (
        .din(new_Jinkela_wire_16248),
        .dout(new_Jinkela_wire_16249)
    );

    bfr new_Jinkela_buffer_10128 (
        .din(new_Jinkela_wire_12277),
        .dout(new_Jinkela_wire_12278)
    );

    bfr new_Jinkela_buffer_6670 (
        .din(new_Jinkela_wire_8393),
        .dout(new_Jinkela_wire_8394)
    );

    bfr new_Jinkela_buffer_13691 (
        .din(new_Jinkela_wire_16348),
        .dout(new_Jinkela_wire_16349)
    );

    bfr new_Jinkela_buffer_3236 (
        .din(new_Jinkela_wire_4357),
        .dout(new_Jinkela_wire_4358)
    );

    bfr new_Jinkela_buffer_10203 (
        .din(new_Jinkela_wire_12366),
        .dout(new_Jinkela_wire_12367)
    );

    bfr new_Jinkela_buffer_6751 (
        .din(new_Jinkela_wire_8476),
        .dout(new_Jinkela_wire_8477)
    );

    bfr new_Jinkela_buffer_13594 (
        .din(new_Jinkela_wire_16249),
        .dout(new_Jinkela_wire_16250)
    );

    bfr new_Jinkela_buffer_3360 (
        .din(new_Jinkela_wire_4489),
        .dout(new_Jinkela_wire_4490)
    );

    bfr new_Jinkela_buffer_10129 (
        .din(new_Jinkela_wire_12278),
        .dout(new_Jinkela_wire_12279)
    );

    bfr new_Jinkela_buffer_6671 (
        .din(new_Jinkela_wire_8394),
        .dout(new_Jinkela_wire_8395)
    );

    bfr new_Jinkela_buffer_13721 (
        .din(new_Jinkela_wire_16382),
        .dout(new_Jinkela_wire_16383)
    );

    bfr new_Jinkela_buffer_3237 (
        .din(new_Jinkela_wire_4358),
        .dout(new_Jinkela_wire_4359)
    );

    bfr new_Jinkela_buffer_10367 (
        .din(new_Jinkela_wire_12534),
        .dout(new_Jinkela_wire_12535)
    );

    spl2 new_Jinkela_splitter_722 (
        .a(_1714_),
        .b(new_Jinkela_wire_8683),
        .c(new_Jinkela_wire_8684)
    );

    bfr new_Jinkela_buffer_13595 (
        .din(new_Jinkela_wire_16250),
        .dout(new_Jinkela_wire_16251)
    );

    bfr new_Jinkela_buffer_3409 (
        .din(_1702_),
        .dout(new_Jinkela_wire_4543)
    );

    bfr new_Jinkela_buffer_10130 (
        .din(new_Jinkela_wire_12279),
        .dout(new_Jinkela_wire_12280)
    );

    bfr new_Jinkela_buffer_6672 (
        .din(new_Jinkela_wire_8395),
        .dout(new_Jinkela_wire_8396)
    );

    bfr new_Jinkela_buffer_13692 (
        .din(new_Jinkela_wire_16349),
        .dout(new_Jinkela_wire_16350)
    );

    bfr new_Jinkela_buffer_3238 (
        .din(new_Jinkela_wire_4359),
        .dout(new_Jinkela_wire_4360)
    );

    bfr new_Jinkela_buffer_10204 (
        .din(new_Jinkela_wire_12367),
        .dout(new_Jinkela_wire_12368)
    );

    spl2 new_Jinkela_splitter_712 (
        .a(new_Jinkela_wire_8477),
        .b(new_Jinkela_wire_8478),
        .c(new_Jinkela_wire_8479)
    );

    bfr new_Jinkela_buffer_13596 (
        .din(new_Jinkela_wire_16251),
        .dout(new_Jinkela_wire_16252)
    );

    bfr new_Jinkela_buffer_3361 (
        .din(new_Jinkela_wire_4490),
        .dout(new_Jinkela_wire_4491)
    );

    bfr new_Jinkela_buffer_10131 (
        .din(new_Jinkela_wire_12280),
        .dout(new_Jinkela_wire_12281)
    );

    bfr new_Jinkela_buffer_6673 (
        .din(new_Jinkela_wire_8396),
        .dout(new_Jinkela_wire_8397)
    );

    bfr new_Jinkela_buffer_13717 (
        .din(new_Jinkela_wire_16376),
        .dout(new_Jinkela_wire_16377)
    );

    bfr new_Jinkela_buffer_3239 (
        .din(new_Jinkela_wire_4360),
        .dout(new_Jinkela_wire_4361)
    );

    bfr new_Jinkela_buffer_13597 (
        .din(new_Jinkela_wire_16252),
        .dout(new_Jinkela_wire_16253)
    );

    spl2 new_Jinkela_splitter_417 (
        .a(_0278_),
        .b(new_Jinkela_wire_4569),
        .c(new_Jinkela_wire_4570)
    );

    bfr new_Jinkela_buffer_6936 (
        .din(_1617_),
        .dout(new_Jinkela_wire_8682)
    );

    bfr new_Jinkela_buffer_10451 (
        .din(_1363_),
        .dout(new_Jinkela_wire_12629)
    );

    bfr new_Jinkela_buffer_6674 (
        .din(new_Jinkela_wire_8397),
        .dout(new_Jinkela_wire_8398)
    );

    bfr new_Jinkela_buffer_3410 (
        .din(new_Jinkela_wire_4543),
        .dout(new_Jinkela_wire_4544)
    );

    bfr new_Jinkela_buffer_10132 (
        .din(new_Jinkela_wire_12281),
        .dout(new_Jinkela_wire_12282)
    );

    bfr new_Jinkela_buffer_3240 (
        .din(new_Jinkela_wire_4361),
        .dout(new_Jinkela_wire_4362)
    );

    bfr new_Jinkela_buffer_13693 (
        .din(new_Jinkela_wire_16350),
        .dout(new_Jinkela_wire_16351)
    );

    bfr new_Jinkela_buffer_10205 (
        .din(new_Jinkela_wire_12368),
        .dout(new_Jinkela_wire_12369)
    );

    bfr new_Jinkela_buffer_6759 (
        .din(new_Jinkela_wire_8490),
        .dout(new_Jinkela_wire_8491)
    );

    bfr new_Jinkela_buffer_13598 (
        .din(new_Jinkela_wire_16253),
        .dout(new_Jinkela_wire_16254)
    );

    bfr new_Jinkela_buffer_3362 (
        .din(new_Jinkela_wire_4491),
        .dout(new_Jinkela_wire_4492)
    );

    bfr new_Jinkela_buffer_10133 (
        .din(new_Jinkela_wire_12282),
        .dout(new_Jinkela_wire_12283)
    );

    bfr new_Jinkela_buffer_6675 (
        .din(new_Jinkela_wire_8398),
        .dout(new_Jinkela_wire_8399)
    );

    bfr new_Jinkela_buffer_3241 (
        .din(new_Jinkela_wire_4362),
        .dout(new_Jinkela_wire_4363)
    );

    bfr new_Jinkela_buffer_13841 (
        .din(_0998_),
        .dout(new_Jinkela_wire_16509)
    );

    bfr new_Jinkela_buffer_10368 (
        .din(new_Jinkela_wire_12535),
        .dout(new_Jinkela_wire_12536)
    );

    bfr new_Jinkela_buffer_6760 (
        .din(new_Jinkela_wire_8491),
        .dout(new_Jinkela_wire_8492)
    );

    bfr new_Jinkela_buffer_13599 (
        .din(new_Jinkela_wire_16254),
        .dout(new_Jinkela_wire_16255)
    );

    bfr new_Jinkela_buffer_6676 (
        .din(new_Jinkela_wire_8399),
        .dout(new_Jinkela_wire_8400)
    );

    bfr new_Jinkela_buffer_3522 (
        .din(_1201_),
        .dout(new_Jinkela_wire_4662)
    );

    bfr new_Jinkela_buffer_10134 (
        .din(new_Jinkela_wire_12283),
        .dout(new_Jinkela_wire_12284)
    );

    bfr new_Jinkela_buffer_3242 (
        .din(new_Jinkela_wire_4363),
        .dout(new_Jinkela_wire_4364)
    );

    bfr new_Jinkela_buffer_13694 (
        .din(new_Jinkela_wire_16351),
        .dout(new_Jinkela_wire_16352)
    );

    bfr new_Jinkela_buffer_10206 (
        .din(new_Jinkela_wire_12369),
        .dout(new_Jinkela_wire_12370)
    );

    bfr new_Jinkela_buffer_6848 (
        .din(new_Jinkela_wire_8591),
        .dout(new_Jinkela_wire_8592)
    );

    bfr new_Jinkela_buffer_13600 (
        .din(new_Jinkela_wire_16255),
        .dout(new_Jinkela_wire_16256)
    );

    bfr new_Jinkela_buffer_3363 (
        .din(new_Jinkela_wire_4492),
        .dout(new_Jinkela_wire_4493)
    );

    bfr new_Jinkela_buffer_10135 (
        .din(new_Jinkela_wire_12284),
        .dout(new_Jinkela_wire_12285)
    );

    bfr new_Jinkela_buffer_6677 (
        .din(new_Jinkela_wire_8400),
        .dout(new_Jinkela_wire_8401)
    );

    spl2 new_Jinkela_splitter_1179 (
        .a(new_Jinkela_wire_16377),
        .b(new_Jinkela_wire_16378),
        .c(new_Jinkela_wire_16379)
    );

    bfr new_Jinkela_buffer_3243 (
        .din(new_Jinkela_wire_4364),
        .dout(new_Jinkela_wire_4365)
    );

    bfr new_Jinkela_buffer_13601 (
        .din(new_Jinkela_wire_16256),
        .dout(new_Jinkela_wire_16257)
    );

    bfr new_Jinkela_buffer_6761 (
        .din(new_Jinkela_wire_8492),
        .dout(new_Jinkela_wire_8493)
    );

    spl2 new_Jinkela_splitter_939 (
        .a(_1623_),
        .b(new_Jinkela_wire_12711),
        .c(new_Jinkela_wire_12712)
    );

    bfr new_Jinkela_buffer_6678 (
        .din(new_Jinkela_wire_8401),
        .dout(new_Jinkela_wire_8402)
    );

    bfr new_Jinkela_buffer_3411 (
        .din(new_Jinkela_wire_4544),
        .dout(new_Jinkela_wire_4545)
    );

    bfr new_Jinkela_buffer_10136 (
        .din(new_Jinkela_wire_12285),
        .dout(new_Jinkela_wire_12286)
    );

    bfr new_Jinkela_buffer_3244 (
        .din(new_Jinkela_wire_4365),
        .dout(new_Jinkela_wire_4366)
    );

    bfr new_Jinkela_buffer_13695 (
        .din(new_Jinkela_wire_16352),
        .dout(new_Jinkela_wire_16353)
    );

    bfr new_Jinkela_buffer_10207 (
        .din(new_Jinkela_wire_12370),
        .dout(new_Jinkela_wire_12371)
    );

    bfr new_Jinkela_buffer_6937 (
        .din(_0802_),
        .dout(new_Jinkela_wire_8685)
    );

    bfr new_Jinkela_buffer_13602 (
        .din(new_Jinkela_wire_16257),
        .dout(new_Jinkela_wire_16258)
    );

    bfr new_Jinkela_buffer_3364 (
        .din(new_Jinkela_wire_4493),
        .dout(new_Jinkela_wire_4494)
    );

    bfr new_Jinkela_buffer_10137 (
        .din(new_Jinkela_wire_12286),
        .dout(new_Jinkela_wire_12287)
    );

    bfr new_Jinkela_buffer_6679 (
        .din(new_Jinkela_wire_8402),
        .dout(new_Jinkela_wire_8403)
    );

    bfr new_Jinkela_buffer_13773 (
        .din(new_Jinkela_wire_16438),
        .dout(new_Jinkela_wire_16439)
    );

    bfr new_Jinkela_buffer_3245 (
        .din(new_Jinkela_wire_4366),
        .dout(new_Jinkela_wire_4367)
    );

    bfr new_Jinkela_buffer_10369 (
        .din(new_Jinkela_wire_12536),
        .dout(new_Jinkela_wire_12537)
    );

    bfr new_Jinkela_buffer_6762 (
        .din(new_Jinkela_wire_8493),
        .dout(new_Jinkela_wire_8494)
    );

    bfr new_Jinkela_buffer_13603 (
        .din(new_Jinkela_wire_16258),
        .dout(new_Jinkela_wire_16259)
    );

    bfr new_Jinkela_buffer_10138 (
        .din(new_Jinkela_wire_12287),
        .dout(new_Jinkela_wire_12288)
    );

    bfr new_Jinkela_buffer_6680 (
        .din(new_Jinkela_wire_8403),
        .dout(new_Jinkela_wire_8404)
    );

    bfr new_Jinkela_buffer_13696 (
        .din(new_Jinkela_wire_16353),
        .dout(new_Jinkela_wire_16354)
    );

    bfr new_Jinkela_buffer_3246 (
        .din(new_Jinkela_wire_4367),
        .dout(new_Jinkela_wire_4368)
    );

    bfr new_Jinkela_buffer_10208 (
        .din(new_Jinkela_wire_12371),
        .dout(new_Jinkela_wire_12372)
    );

    bfr new_Jinkela_buffer_6849 (
        .din(new_Jinkela_wire_8592),
        .dout(new_Jinkela_wire_8593)
    );

    bfr new_Jinkela_buffer_13604 (
        .din(new_Jinkela_wire_16259),
        .dout(new_Jinkela_wire_16260)
    );

    bfr new_Jinkela_buffer_3365 (
        .din(new_Jinkela_wire_4494),
        .dout(new_Jinkela_wire_4495)
    );

    bfr new_Jinkela_buffer_10139 (
        .din(new_Jinkela_wire_12288),
        .dout(new_Jinkela_wire_12289)
    );

    bfr new_Jinkela_buffer_6681 (
        .din(new_Jinkela_wire_8404),
        .dout(new_Jinkela_wire_8405)
    );

    bfr new_Jinkela_buffer_13722 (
        .din(new_Jinkela_wire_16383),
        .dout(new_Jinkela_wire_16384)
    );

    bfr new_Jinkela_buffer_3247 (
        .din(new_Jinkela_wire_4368),
        .dout(new_Jinkela_wire_4369)
    );

    bfr new_Jinkela_buffer_10452 (
        .din(new_Jinkela_wire_12629),
        .dout(new_Jinkela_wire_12630)
    );

    bfr new_Jinkela_buffer_6763 (
        .din(new_Jinkela_wire_8494),
        .dout(new_Jinkela_wire_8495)
    );

    bfr new_Jinkela_buffer_13605 (
        .din(new_Jinkela_wire_16260),
        .dout(new_Jinkela_wire_16261)
    );

    bfr new_Jinkela_buffer_3521 (
        .din(_1397_),
        .dout(new_Jinkela_wire_4661)
    );

    bfr new_Jinkela_buffer_6682 (
        .din(new_Jinkela_wire_8405),
        .dout(new_Jinkela_wire_8406)
    );

    bfr new_Jinkela_buffer_3412 (
        .din(new_Jinkela_wire_4545),
        .dout(new_Jinkela_wire_4546)
    );

    bfr new_Jinkela_buffer_10140 (
        .din(new_Jinkela_wire_12289),
        .dout(new_Jinkela_wire_12290)
    );

    bfr new_Jinkela_buffer_3248 (
        .din(new_Jinkela_wire_4369),
        .dout(new_Jinkela_wire_4370)
    );

    bfr new_Jinkela_buffer_13697 (
        .din(new_Jinkela_wire_16354),
        .dout(new_Jinkela_wire_16355)
    );

    bfr new_Jinkela_buffer_10209 (
        .din(new_Jinkela_wire_12372),
        .dout(new_Jinkela_wire_12373)
    );

    spl2 new_Jinkela_splitter_723 (
        .a(_0055_),
        .b(new_Jinkela_wire_8686),
        .c(new_Jinkela_wire_8687)
    );

    bfr new_Jinkela_buffer_13606 (
        .din(new_Jinkela_wire_16261),
        .dout(new_Jinkela_wire_16262)
    );

    bfr new_Jinkela_buffer_3366 (
        .din(new_Jinkela_wire_4495),
        .dout(new_Jinkela_wire_4496)
    );

    bfr new_Jinkela_buffer_10141 (
        .din(new_Jinkela_wire_12290),
        .dout(new_Jinkela_wire_12291)
    );

    bfr new_Jinkela_buffer_6683 (
        .din(new_Jinkela_wire_8406),
        .dout(new_Jinkela_wire_8407)
    );

    bfr new_Jinkela_buffer_13723 (
        .din(new_Jinkela_wire_16384),
        .dout(new_Jinkela_wire_16385)
    );

    bfr new_Jinkela_buffer_3249 (
        .din(new_Jinkela_wire_4370),
        .dout(new_Jinkela_wire_4371)
    );

    spl2 new_Jinkela_splitter_1497 (
        .a(_1535_),
        .b(new_Jinkela_wire_20346),
        .c(new_Jinkela_wire_20347)
    );

    bfr new_Jinkela_buffer_17045 (
        .din(new_Jinkela_wire_20341),
        .dout(new_Jinkela_wire_20342)
    );

    bfr new_Jinkela_buffer_17023 (
        .din(new_Jinkela_wire_20307),
        .dout(new_Jinkela_wire_20308)
    );

    bfr new_Jinkela_buffer_17041 (
        .din(new_Jinkela_wire_20335),
        .dout(new_Jinkela_wire_20336)
    );

    bfr new_Jinkela_buffer_17024 (
        .din(new_Jinkela_wire_20308),
        .dout(new_Jinkela_wire_20309)
    );

    bfr new_Jinkela_buffer_17025 (
        .din(new_Jinkela_wire_20309),
        .dout(new_Jinkela_wire_20310)
    );

    bfr new_Jinkela_buffer_17042 (
        .din(new_Jinkela_wire_20336),
        .dout(new_Jinkela_wire_20337)
    );

    bfr new_Jinkela_buffer_17026 (
        .din(new_Jinkela_wire_20310),
        .dout(new_Jinkela_wire_20311)
    );

    bfr new_Jinkela_buffer_17049 (
        .din(_1660_),
        .dout(new_Jinkela_wire_20348)
    );

    bfr new_Jinkela_buffer_17027 (
        .din(new_Jinkela_wire_20311),
        .dout(new_Jinkela_wire_20312)
    );

    bfr new_Jinkela_buffer_17043 (
        .din(new_Jinkela_wire_20337),
        .dout(new_Jinkela_wire_20338)
    );

    bfr new_Jinkela_buffer_17028 (
        .din(new_Jinkela_wire_20312),
        .dout(new_Jinkela_wire_20313)
    );

    bfr new_Jinkela_buffer_17050 (
        .din(new_Jinkela_wire_20350),
        .dout(new_Jinkela_wire_20351)
    );

    bfr new_Jinkela_buffer_17029 (
        .din(new_Jinkela_wire_20313),
        .dout(new_Jinkela_wire_20314)
    );

    bfr new_Jinkela_buffer_17046 (
        .din(new_Jinkela_wire_20342),
        .dout(new_Jinkela_wire_20343)
    );

    bfr new_Jinkela_buffer_17030 (
        .din(new_Jinkela_wire_20314),
        .dout(new_Jinkela_wire_20315)
    );

    spl2 new_Jinkela_splitter_1499 (
        .a(_0351_),
        .b(new_Jinkela_wire_20355),
        .c(new_Jinkela_wire_20356)
    );

    spl2 new_Jinkela_splitter_1498 (
        .a(_1732_),
        .b(new_Jinkela_wire_20349),
        .c(new_Jinkela_wire_20350)
    );

    bfr new_Jinkela_buffer_17031 (
        .din(new_Jinkela_wire_20315),
        .dout(new_Jinkela_wire_20316)
    );

    bfr new_Jinkela_buffer_17047 (
        .din(new_Jinkela_wire_20343),
        .dout(new_Jinkela_wire_20344)
    );

    bfr new_Jinkela_buffer_17032 (
        .din(new_Jinkela_wire_20316),
        .dout(new_Jinkela_wire_20317)
    );

    bfr new_Jinkela_buffer_17033 (
        .din(new_Jinkela_wire_20317),
        .dout(new_Jinkela_wire_20318)
    );

    bfr new_Jinkela_buffer_17048 (
        .din(new_Jinkela_wire_20344),
        .dout(new_Jinkela_wire_20345)
    );

    spl2 new_Jinkela_splitter_1491 (
        .a(new_Jinkela_wire_20318),
        .b(new_Jinkela_wire_20319),
        .c(new_Jinkela_wire_20320)
    );

    spl2 new_Jinkela_splitter_1500 (
        .a(_0458_),
        .b(new_Jinkela_wire_20357),
        .c(new_Jinkela_wire_20358)
    );

    bfr new_Jinkela_buffer_17051 (
        .din(new_Jinkela_wire_20351),
        .dout(new_Jinkela_wire_20352)
    );

    bfr new_Jinkela_buffer_17054 (
        .din(_1523_),
        .dout(new_Jinkela_wire_20359)
    );

    bfr new_Jinkela_buffer_17052 (
        .din(new_Jinkela_wire_20352),
        .dout(new_Jinkela_wire_20353)
    );

    spl2 new_Jinkela_splitter_1502 (
        .a(_0639_),
        .b(new_Jinkela_wire_20362),
        .c(new_Jinkela_wire_20363)
    );

    spl2 new_Jinkela_splitter_1501 (
        .a(_1513_),
        .b(new_Jinkela_wire_20360),
        .c(new_Jinkela_wire_20361)
    );

    bfr new_Jinkela_buffer_17053 (
        .din(new_Jinkela_wire_20353),
        .dout(new_Jinkela_wire_20354)
    );

    spl2 new_Jinkela_splitter_1503 (
        .a(_0697_),
        .b(new_Jinkela_wire_20364),
        .c(new_Jinkela_wire_20365)
    );

    bfr new_Jinkela_buffer_17055 (
        .din(_0392_),
        .dout(new_Jinkela_wire_20366)
    );

    spl2 new_Jinkela_splitter_1505 (
        .a(_0590_),
        .b(new_Jinkela_wire_20369),
        .c(new_Jinkela_wire_20370)
    );

    spl2 new_Jinkela_splitter_1504 (
        .a(_0856_),
        .b(new_Jinkela_wire_20367),
        .c(new_Jinkela_wire_20368)
    );

    spl2 new_Jinkela_splitter_1506 (
        .a(_1108_),
        .b(new_Jinkela_wire_20371),
        .c(new_Jinkela_wire_20372)
    );

    spl2 new_Jinkela_splitter_1507 (
        .a(_0067_),
        .b(new_Jinkela_wire_20373),
        .c(new_Jinkela_wire_20374)
    );

    spl2 new_Jinkela_splitter_1508 (
        .a(_0404_),
        .b(new_Jinkela_wire_20375),
        .c(new_Jinkela_wire_20376)
    );

    spl2 new_Jinkela_splitter_1509 (
        .a(_1605_),
        .b(new_Jinkela_wire_20381),
        .c(new_Jinkela_wire_20382)
    );

    bfr new_Jinkela_buffer_17056 (
        .din(new_Jinkela_wire_20376),
        .dout(new_Jinkela_wire_20377)
    );

    spl2 new_Jinkela_splitter_1510 (
        .a(_1263_),
        .b(new_Jinkela_wire_20383),
        .c(new_Jinkela_wire_20384)
    );

    bfr new_Jinkela_buffer_17060 (
        .din(_1786_),
        .dout(new_Jinkela_wire_20385)
    );

    bfr new_Jinkela_buffer_13607 (
        .din(new_Jinkela_wire_16262),
        .dout(new_Jinkela_wire_16263)
    );

    bfr new_Jinkela_buffer_3434 (
        .din(new_Jinkela_wire_4571),
        .dout(new_Jinkela_wire_4572)
    );

    bfr new_Jinkela_buffer_13698 (
        .din(new_Jinkela_wire_16355),
        .dout(new_Jinkela_wire_16356)
    );

    bfr new_Jinkela_buffer_3250 (
        .din(new_Jinkela_wire_4371),
        .dout(new_Jinkela_wire_4372)
    );

    bfr new_Jinkela_buffer_13608 (
        .din(new_Jinkela_wire_16263),
        .dout(new_Jinkela_wire_16264)
    );

    bfr new_Jinkela_buffer_3367 (
        .din(new_Jinkela_wire_4496),
        .dout(new_Jinkela_wire_4497)
    );

    bfr new_Jinkela_buffer_13777 (
        .din(new_Jinkela_wire_16442),
        .dout(new_Jinkela_wire_16443)
    );

    bfr new_Jinkela_buffer_3251 (
        .din(new_Jinkela_wire_4372),
        .dout(new_Jinkela_wire_4373)
    );

    bfr new_Jinkela_buffer_13609 (
        .din(new_Jinkela_wire_16264),
        .dout(new_Jinkela_wire_16265)
    );

    bfr new_Jinkela_buffer_3413 (
        .din(new_Jinkela_wire_4546),
        .dout(new_Jinkela_wire_4547)
    );

    bfr new_Jinkela_buffer_13699 (
        .din(new_Jinkela_wire_16356),
        .dout(new_Jinkela_wire_16357)
    );

    bfr new_Jinkela_buffer_3252 (
        .din(new_Jinkela_wire_4373),
        .dout(new_Jinkela_wire_4374)
    );

    bfr new_Jinkela_buffer_13610 (
        .din(new_Jinkela_wire_16265),
        .dout(new_Jinkela_wire_16266)
    );

    bfr new_Jinkela_buffer_3368 (
        .din(new_Jinkela_wire_4497),
        .dout(new_Jinkela_wire_4498)
    );

    bfr new_Jinkela_buffer_13724 (
        .din(new_Jinkela_wire_16385),
        .dout(new_Jinkela_wire_16386)
    );

    bfr new_Jinkela_buffer_3253 (
        .din(new_Jinkela_wire_4374),
        .dout(new_Jinkela_wire_4375)
    );

    bfr new_Jinkela_buffer_13611 (
        .din(new_Jinkela_wire_16266),
        .dout(new_Jinkela_wire_16267)
    );

    bfr new_Jinkela_buffer_13700 (
        .din(new_Jinkela_wire_16357),
        .dout(new_Jinkela_wire_16358)
    );

    bfr new_Jinkela_buffer_3254 (
        .din(new_Jinkela_wire_4375),
        .dout(new_Jinkela_wire_4376)
    );

    bfr new_Jinkela_buffer_13612 (
        .din(new_Jinkela_wire_16267),
        .dout(new_Jinkela_wire_16268)
    );

    bfr new_Jinkela_buffer_3369 (
        .din(new_Jinkela_wire_4498),
        .dout(new_Jinkela_wire_4499)
    );

    bfr new_Jinkela_buffer_13774 (
        .din(new_Jinkela_wire_16439),
        .dout(new_Jinkela_wire_16440)
    );

    bfr new_Jinkela_buffer_3255 (
        .din(new_Jinkela_wire_4376),
        .dout(new_Jinkela_wire_4377)
    );

    bfr new_Jinkela_buffer_13613 (
        .din(new_Jinkela_wire_16268),
        .dout(new_Jinkela_wire_16269)
    );

    bfr new_Jinkela_buffer_3523 (
        .din(_1318_),
        .dout(new_Jinkela_wire_4663)
    );

    bfr new_Jinkela_buffer_3414 (
        .din(new_Jinkela_wire_4547),
        .dout(new_Jinkela_wire_4548)
    );

    bfr new_Jinkela_buffer_13701 (
        .din(new_Jinkela_wire_16358),
        .dout(new_Jinkela_wire_16359)
    );

    bfr new_Jinkela_buffer_3256 (
        .din(new_Jinkela_wire_4377),
        .dout(new_Jinkela_wire_4378)
    );

    bfr new_Jinkela_buffer_13614 (
        .din(new_Jinkela_wire_16269),
        .dout(new_Jinkela_wire_16270)
    );

    bfr new_Jinkela_buffer_3370 (
        .din(new_Jinkela_wire_4499),
        .dout(new_Jinkela_wire_4500)
    );

    bfr new_Jinkela_buffer_13725 (
        .din(new_Jinkela_wire_16386),
        .dout(new_Jinkela_wire_16387)
    );

    bfr new_Jinkela_buffer_3257 (
        .din(new_Jinkela_wire_4378),
        .dout(new_Jinkela_wire_4379)
    );

    bfr new_Jinkela_buffer_13615 (
        .din(new_Jinkela_wire_16270),
        .dout(new_Jinkela_wire_16271)
    );

    bfr new_Jinkela_buffer_3435 (
        .din(new_Jinkela_wire_4572),
        .dout(new_Jinkela_wire_4573)
    );

    bfr new_Jinkela_buffer_13702 (
        .din(new_Jinkela_wire_16359),
        .dout(new_Jinkela_wire_16360)
    );

    bfr new_Jinkela_buffer_3258 (
        .din(new_Jinkela_wire_4379),
        .dout(new_Jinkela_wire_4380)
    );

    bfr new_Jinkela_buffer_13616 (
        .din(new_Jinkela_wire_16271),
        .dout(new_Jinkela_wire_16272)
    );

    bfr new_Jinkela_buffer_3371 (
        .din(new_Jinkela_wire_4500),
        .dout(new_Jinkela_wire_4501)
    );

    bfr new_Jinkela_buffer_3259 (
        .din(new_Jinkela_wire_4380),
        .dout(new_Jinkela_wire_4381)
    );

    bfr new_Jinkela_buffer_13842 (
        .din(_1799_),
        .dout(new_Jinkela_wire_16510)
    );

    bfr new_Jinkela_buffer_13617 (
        .din(new_Jinkela_wire_16272),
        .dout(new_Jinkela_wire_16273)
    );

    bfr new_Jinkela_buffer_3415 (
        .din(new_Jinkela_wire_4548),
        .dout(new_Jinkela_wire_4549)
    );

    bfr new_Jinkela_buffer_13703 (
        .din(new_Jinkela_wire_16360),
        .dout(new_Jinkela_wire_16361)
    );

    bfr new_Jinkela_buffer_3260 (
        .din(new_Jinkela_wire_4381),
        .dout(new_Jinkela_wire_4382)
    );

    bfr new_Jinkela_buffer_13618 (
        .din(new_Jinkela_wire_16273),
        .dout(new_Jinkela_wire_16274)
    );

    bfr new_Jinkela_buffer_3372 (
        .din(new_Jinkela_wire_4501),
        .dout(new_Jinkela_wire_4502)
    );

    bfr new_Jinkela_buffer_13726 (
        .din(new_Jinkela_wire_16387),
        .dout(new_Jinkela_wire_16388)
    );

    bfr new_Jinkela_buffer_3261 (
        .din(new_Jinkela_wire_4382),
        .dout(new_Jinkela_wire_4383)
    );

    bfr new_Jinkela_buffer_13619 (
        .din(new_Jinkela_wire_16274),
        .dout(new_Jinkela_wire_16275)
    );

    bfr new_Jinkela_buffer_13704 (
        .din(new_Jinkela_wire_16361),
        .dout(new_Jinkela_wire_16362)
    );

    bfr new_Jinkela_buffer_3262 (
        .din(new_Jinkela_wire_4383),
        .dout(new_Jinkela_wire_4384)
    );

    bfr new_Jinkela_buffer_13620 (
        .din(new_Jinkela_wire_16275),
        .dout(new_Jinkela_wire_16276)
    );

    bfr new_Jinkela_buffer_3373 (
        .din(new_Jinkela_wire_4502),
        .dout(new_Jinkela_wire_4503)
    );

    bfr new_Jinkela_buffer_13775 (
        .din(new_Jinkela_wire_16440),
        .dout(new_Jinkela_wire_16441)
    );

    bfr new_Jinkela_buffer_3263 (
        .din(new_Jinkela_wire_4384),
        .dout(new_Jinkela_wire_4385)
    );

    bfr new_Jinkela_buffer_13621 (
        .din(new_Jinkela_wire_16276),
        .dout(new_Jinkela_wire_16277)
    );

    spl2 new_Jinkela_splitter_419 (
        .a(_1508_),
        .b(new_Jinkela_wire_4664),
        .c(new_Jinkela_wire_4665)
    );

    bfr new_Jinkela_buffer_3416 (
        .din(new_Jinkela_wire_4549),
        .dout(new_Jinkela_wire_4550)
    );

    bfr new_Jinkela_buffer_13705 (
        .din(new_Jinkela_wire_16362),
        .dout(new_Jinkela_wire_16363)
    );

    bfr new_Jinkela_buffer_3264 (
        .din(new_Jinkela_wire_4385),
        .dout(new_Jinkela_wire_4386)
    );

    bfr new_Jinkela_buffer_13622 (
        .din(new_Jinkela_wire_16277),
        .dout(new_Jinkela_wire_16278)
    );

    bfr new_Jinkela_buffer_3374 (
        .din(new_Jinkela_wire_4503),
        .dout(new_Jinkela_wire_4504)
    );

    bfr new_Jinkela_buffer_13727 (
        .din(new_Jinkela_wire_16388),
        .dout(new_Jinkela_wire_16389)
    );

    bfr new_Jinkela_buffer_3265 (
        .din(new_Jinkela_wire_4386),
        .dout(new_Jinkela_wire_4387)
    );

    bfr new_Jinkela_buffer_13623 (
        .din(new_Jinkela_wire_16278),
        .dout(new_Jinkela_wire_16279)
    );

    bfr new_Jinkela_buffer_3436 (
        .din(new_Jinkela_wire_4573),
        .dout(new_Jinkela_wire_4574)
    );

    bfr new_Jinkela_buffer_13706 (
        .din(new_Jinkela_wire_16363),
        .dout(new_Jinkela_wire_16364)
    );

    bfr new_Jinkela_buffer_3266 (
        .din(new_Jinkela_wire_4387),
        .dout(new_Jinkela_wire_4388)
    );

    bfr new_Jinkela_buffer_13624 (
        .din(new_Jinkela_wire_16279),
        .dout(new_Jinkela_wire_16280)
    );

    bfr new_Jinkela_buffer_3375 (
        .din(new_Jinkela_wire_4504),
        .dout(new_Jinkela_wire_4505)
    );

    bfr new_Jinkela_buffer_13778 (
        .din(new_Jinkela_wire_16443),
        .dout(new_Jinkela_wire_16444)
    );

    bfr new_Jinkela_buffer_3267 (
        .din(new_Jinkela_wire_4388),
        .dout(new_Jinkela_wire_4389)
    );

    bfr new_Jinkela_buffer_13625 (
        .din(new_Jinkela_wire_16280),
        .dout(new_Jinkela_wire_16281)
    );

    bfr new_Jinkela_buffer_3417 (
        .din(new_Jinkela_wire_4550),
        .dout(new_Jinkela_wire_4551)
    );

    bfr new_Jinkela_buffer_13707 (
        .din(new_Jinkela_wire_16364),
        .dout(new_Jinkela_wire_16365)
    );

    bfr new_Jinkela_buffer_3268 (
        .din(new_Jinkela_wire_4389),
        .dout(new_Jinkela_wire_4390)
    );

    bfr new_Jinkela_buffer_13626 (
        .din(new_Jinkela_wire_16281),
        .dout(new_Jinkela_wire_16282)
    );

    bfr new_Jinkela_buffer_3376 (
        .din(new_Jinkela_wire_4505),
        .dout(new_Jinkela_wire_4506)
    );

    bfr new_Jinkela_buffer_13728 (
        .din(new_Jinkela_wire_16389),
        .dout(new_Jinkela_wire_16390)
    );

    bfr new_Jinkela_buffer_3269 (
        .din(new_Jinkela_wire_4390),
        .dout(new_Jinkela_wire_4391)
    );

    bfr new_Jinkela_buffer_13627 (
        .din(new_Jinkela_wire_16282),
        .dout(new_Jinkela_wire_16283)
    );

    bfr new_Jinkela_buffer_3524 (
        .din(_0056_),
        .dout(new_Jinkela_wire_4666)
    );

    spl2 new_Jinkela_splitter_1178 (
        .a(new_Jinkela_wire_16365),
        .b(new_Jinkela_wire_16366),
        .c(new_Jinkela_wire_16367)
    );

    bfr new_Jinkela_buffer_3270 (
        .din(new_Jinkela_wire_4391),
        .dout(new_Jinkela_wire_4392)
    );

    bfr new_Jinkela_buffer_10370 (
        .din(new_Jinkela_wire_12537),
        .dout(new_Jinkela_wire_12538)
    );

    bfr new_Jinkela_buffer_10142 (
        .din(new_Jinkela_wire_12291),
        .dout(new_Jinkela_wire_12292)
    );

    bfr new_Jinkela_buffer_10210 (
        .din(new_Jinkela_wire_12373),
        .dout(new_Jinkela_wire_12374)
    );

    bfr new_Jinkela_buffer_10143 (
        .din(new_Jinkela_wire_12292),
        .dout(new_Jinkela_wire_12293)
    );

    bfr new_Jinkela_buffer_10144 (
        .din(new_Jinkela_wire_12293),
        .dout(new_Jinkela_wire_12294)
    );

    bfr new_Jinkela_buffer_10211 (
        .din(new_Jinkela_wire_12374),
        .dout(new_Jinkela_wire_12375)
    );

    bfr new_Jinkela_buffer_10145 (
        .din(new_Jinkela_wire_12294),
        .dout(new_Jinkela_wire_12295)
    );

    bfr new_Jinkela_buffer_10371 (
        .din(new_Jinkela_wire_12538),
        .dout(new_Jinkela_wire_12539)
    );

    bfr new_Jinkela_buffer_10146 (
        .din(new_Jinkela_wire_12295),
        .dout(new_Jinkela_wire_12296)
    );

    bfr new_Jinkela_buffer_10212 (
        .din(new_Jinkela_wire_12375),
        .dout(new_Jinkela_wire_12376)
    );

    bfr new_Jinkela_buffer_10147 (
        .din(new_Jinkela_wire_12296),
        .dout(new_Jinkela_wire_12297)
    );

    bfr new_Jinkela_buffer_10453 (
        .din(new_Jinkela_wire_12630),
        .dout(new_Jinkela_wire_12631)
    );

    bfr new_Jinkela_buffer_10148 (
        .din(new_Jinkela_wire_12297),
        .dout(new_Jinkela_wire_12298)
    );

    bfr new_Jinkela_buffer_10213 (
        .din(new_Jinkela_wire_12376),
        .dout(new_Jinkela_wire_12377)
    );

    bfr new_Jinkela_buffer_10149 (
        .din(new_Jinkela_wire_12298),
        .dout(new_Jinkela_wire_12299)
    );

    bfr new_Jinkela_buffer_10372 (
        .din(new_Jinkela_wire_12539),
        .dout(new_Jinkela_wire_12540)
    );

    bfr new_Jinkela_buffer_10150 (
        .din(new_Jinkela_wire_12299),
        .dout(new_Jinkela_wire_12300)
    );

    bfr new_Jinkela_buffer_10214 (
        .din(new_Jinkela_wire_12377),
        .dout(new_Jinkela_wire_12378)
    );

    bfr new_Jinkela_buffer_10151 (
        .din(new_Jinkela_wire_12300),
        .dout(new_Jinkela_wire_12301)
    );

    spl2 new_Jinkela_splitter_941 (
        .a(_1317_),
        .b(new_Jinkela_wire_12715),
        .c(new_Jinkela_wire_12716)
    );

    bfr new_Jinkela_buffer_10152 (
        .din(new_Jinkela_wire_12301),
        .dout(new_Jinkela_wire_12302)
    );

    bfr new_Jinkela_buffer_10215 (
        .din(new_Jinkela_wire_12378),
        .dout(new_Jinkela_wire_12379)
    );

    bfr new_Jinkela_buffer_10153 (
        .din(new_Jinkela_wire_12302),
        .dout(new_Jinkela_wire_12303)
    );

    bfr new_Jinkela_buffer_10373 (
        .din(new_Jinkela_wire_12540),
        .dout(new_Jinkela_wire_12541)
    );

    bfr new_Jinkela_buffer_10154 (
        .din(new_Jinkela_wire_12303),
        .dout(new_Jinkela_wire_12304)
    );

    bfr new_Jinkela_buffer_10216 (
        .din(new_Jinkela_wire_12379),
        .dout(new_Jinkela_wire_12380)
    );

    bfr new_Jinkela_buffer_10155 (
        .din(new_Jinkela_wire_12304),
        .dout(new_Jinkela_wire_12305)
    );

    bfr new_Jinkela_buffer_10454 (
        .din(new_Jinkela_wire_12631),
        .dout(new_Jinkela_wire_12632)
    );

    bfr new_Jinkela_buffer_10156 (
        .din(new_Jinkela_wire_12305),
        .dout(new_Jinkela_wire_12306)
    );

    bfr new_Jinkela_buffer_10217 (
        .din(new_Jinkela_wire_12380),
        .dout(new_Jinkela_wire_12381)
    );

    bfr new_Jinkela_buffer_10157 (
        .din(new_Jinkela_wire_12306),
        .dout(new_Jinkela_wire_12307)
    );

    bfr new_Jinkela_buffer_10374 (
        .din(new_Jinkela_wire_12541),
        .dout(new_Jinkela_wire_12542)
    );

    bfr new_Jinkela_buffer_10158 (
        .din(new_Jinkela_wire_12307),
        .dout(new_Jinkela_wire_12308)
    );

    bfr new_Jinkela_buffer_10218 (
        .din(new_Jinkela_wire_12381),
        .dout(new_Jinkela_wire_12382)
    );

    bfr new_Jinkela_buffer_10159 (
        .din(new_Jinkela_wire_12308),
        .dout(new_Jinkela_wire_12309)
    );

    bfr new_Jinkela_buffer_10535 (
        .din(_1720_),
        .dout(new_Jinkela_wire_12723)
    );

    spl2 new_Jinkela_splitter_942 (
        .a(_0495_),
        .b(new_Jinkela_wire_12717),
        .c(new_Jinkela_wire_12718)
    );

    bfr new_Jinkela_buffer_10160 (
        .din(new_Jinkela_wire_12309),
        .dout(new_Jinkela_wire_12310)
    );

    bfr new_Jinkela_buffer_10219 (
        .din(new_Jinkela_wire_12382),
        .dout(new_Jinkela_wire_12383)
    );

    bfr new_Jinkela_buffer_10161 (
        .din(new_Jinkela_wire_12310),
        .dout(new_Jinkela_wire_12311)
    );

    bfr new_Jinkela_buffer_10375 (
        .din(new_Jinkela_wire_12542),
        .dout(new_Jinkela_wire_12543)
    );

    bfr new_Jinkela_buffer_10162 (
        .din(new_Jinkela_wire_12311),
        .dout(new_Jinkela_wire_12312)
    );

    bfr new_Jinkela_buffer_6764 (
        .din(new_Jinkela_wire_8495),
        .dout(new_Jinkela_wire_8496)
    );

    bfr new_Jinkela_buffer_13628 (
        .din(new_Jinkela_wire_16283),
        .dout(new_Jinkela_wire_16284)
    );

    bfr new_Jinkela_buffer_6684 (
        .din(new_Jinkela_wire_8407),
        .dout(new_Jinkela_wire_8408)
    );

    bfr new_Jinkela_buffer_13729 (
        .din(new_Jinkela_wire_16390),
        .dout(new_Jinkela_wire_16391)
    );

    bfr new_Jinkela_buffer_6850 (
        .din(new_Jinkela_wire_8593),
        .dout(new_Jinkela_wire_8594)
    );

    bfr new_Jinkela_buffer_13629 (
        .din(new_Jinkela_wire_16284),
        .dout(new_Jinkela_wire_16285)
    );

    bfr new_Jinkela_buffer_6685 (
        .din(new_Jinkela_wire_8408),
        .dout(new_Jinkela_wire_8409)
    );

    bfr new_Jinkela_buffer_13843 (
        .din(_1487_),
        .dout(new_Jinkela_wire_16511)
    );

    bfr new_Jinkela_buffer_6765 (
        .din(new_Jinkela_wire_8496),
        .dout(new_Jinkela_wire_8497)
    );

    bfr new_Jinkela_buffer_13630 (
        .din(new_Jinkela_wire_16285),
        .dout(new_Jinkela_wire_16286)
    );

    bfr new_Jinkela_buffer_6686 (
        .din(new_Jinkela_wire_8409),
        .dout(new_Jinkela_wire_8410)
    );

    bfr new_Jinkela_buffer_13779 (
        .din(new_Jinkela_wire_16444),
        .dout(new_Jinkela_wire_16445)
    );

    spl2 new_Jinkela_splitter_725 (
        .a(_0228_),
        .b(new_Jinkela_wire_8691),
        .c(new_Jinkela_wire_8692)
    );

    bfr new_Jinkela_buffer_13631 (
        .din(new_Jinkela_wire_16286),
        .dout(new_Jinkela_wire_16287)
    );

    bfr new_Jinkela_buffer_6687 (
        .din(new_Jinkela_wire_8410),
        .dout(new_Jinkela_wire_8411)
    );

    bfr new_Jinkela_buffer_13730 (
        .din(new_Jinkela_wire_16391),
        .dout(new_Jinkela_wire_16392)
    );

    bfr new_Jinkela_buffer_6766 (
        .din(new_Jinkela_wire_8497),
        .dout(new_Jinkela_wire_8498)
    );

    bfr new_Jinkela_buffer_13632 (
        .din(new_Jinkela_wire_16287),
        .dout(new_Jinkela_wire_16288)
    );

    bfr new_Jinkela_buffer_6688 (
        .din(new_Jinkela_wire_8411),
        .dout(new_Jinkela_wire_8412)
    );

    spl2 new_Jinkela_splitter_1183 (
        .a(_0947_),
        .b(new_Jinkela_wire_16512),
        .c(new_Jinkela_wire_16513)
    );

    bfr new_Jinkela_buffer_6851 (
        .din(new_Jinkela_wire_8594),
        .dout(new_Jinkela_wire_8595)
    );

    bfr new_Jinkela_buffer_13633 (
        .din(new_Jinkela_wire_16288),
        .dout(new_Jinkela_wire_16289)
    );

    bfr new_Jinkela_buffer_6689 (
        .din(new_Jinkela_wire_8412),
        .dout(new_Jinkela_wire_8413)
    );

    bfr new_Jinkela_buffer_13731 (
        .din(new_Jinkela_wire_16392),
        .dout(new_Jinkela_wire_16393)
    );

    bfr new_Jinkela_buffer_6767 (
        .din(new_Jinkela_wire_8498),
        .dout(new_Jinkela_wire_8499)
    );

    bfr new_Jinkela_buffer_13634 (
        .din(new_Jinkela_wire_16289),
        .dout(new_Jinkela_wire_16290)
    );

    bfr new_Jinkela_buffer_6690 (
        .din(new_Jinkela_wire_8413),
        .dout(new_Jinkela_wire_8414)
    );

    bfr new_Jinkela_buffer_13780 (
        .din(new_Jinkela_wire_16445),
        .dout(new_Jinkela_wire_16446)
    );

    bfr new_Jinkela_buffer_6939 (
        .din(_1277_),
        .dout(new_Jinkela_wire_8693)
    );

    bfr new_Jinkela_buffer_13635 (
        .din(new_Jinkela_wire_16290),
        .dout(new_Jinkela_wire_16291)
    );

    bfr new_Jinkela_buffer_6691 (
        .din(new_Jinkela_wire_8414),
        .dout(new_Jinkela_wire_8415)
    );

    bfr new_Jinkela_buffer_13732 (
        .din(new_Jinkela_wire_16393),
        .dout(new_Jinkela_wire_16394)
    );

    bfr new_Jinkela_buffer_6768 (
        .din(new_Jinkela_wire_8499),
        .dout(new_Jinkela_wire_8500)
    );

    bfr new_Jinkela_buffer_13636 (
        .din(new_Jinkela_wire_16291),
        .dout(new_Jinkela_wire_16292)
    );

    bfr new_Jinkela_buffer_6692 (
        .din(new_Jinkela_wire_8415),
        .dout(new_Jinkela_wire_8416)
    );

    spl2 new_Jinkela_splitter_1184 (
        .a(_1402_),
        .b(new_Jinkela_wire_16514),
        .c(new_Jinkela_wire_16515)
    );

    bfr new_Jinkela_buffer_13844 (
        .din(new_Jinkela_wire_16517),
        .dout(new_Jinkela_wire_16518)
    );

    bfr new_Jinkela_buffer_6852 (
        .din(new_Jinkela_wire_8595),
        .dout(new_Jinkela_wire_8596)
    );

    bfr new_Jinkela_buffer_13637 (
        .din(new_Jinkela_wire_16292),
        .dout(new_Jinkela_wire_16293)
    );

    bfr new_Jinkela_buffer_6693 (
        .din(new_Jinkela_wire_8416),
        .dout(new_Jinkela_wire_8417)
    );

    bfr new_Jinkela_buffer_13733 (
        .din(new_Jinkela_wire_16394),
        .dout(new_Jinkela_wire_16395)
    );

    bfr new_Jinkela_buffer_6769 (
        .din(new_Jinkela_wire_8500),
        .dout(new_Jinkela_wire_8501)
    );

    bfr new_Jinkela_buffer_13638 (
        .din(new_Jinkela_wire_16293),
        .dout(new_Jinkela_wire_16294)
    );

    bfr new_Jinkela_buffer_6694 (
        .din(new_Jinkela_wire_8417),
        .dout(new_Jinkela_wire_8418)
    );

    bfr new_Jinkela_buffer_13781 (
        .din(new_Jinkela_wire_16446),
        .dout(new_Jinkela_wire_16447)
    );

    bfr new_Jinkela_buffer_6940 (
        .din(_1282_),
        .dout(new_Jinkela_wire_8694)
    );

    bfr new_Jinkela_buffer_13639 (
        .din(new_Jinkela_wire_16294),
        .dout(new_Jinkela_wire_16295)
    );

    bfr new_Jinkela_buffer_6938 (
        .din(new_Jinkela_wire_8687),
        .dout(new_Jinkela_wire_8688)
    );

    bfr new_Jinkela_buffer_6695 (
        .din(new_Jinkela_wire_8418),
        .dout(new_Jinkela_wire_8419)
    );

    bfr new_Jinkela_buffer_13734 (
        .din(new_Jinkela_wire_16395),
        .dout(new_Jinkela_wire_16396)
    );

    bfr new_Jinkela_buffer_6770 (
        .din(new_Jinkela_wire_8501),
        .dout(new_Jinkela_wire_8502)
    );

    bfr new_Jinkela_buffer_13640 (
        .din(new_Jinkela_wire_16295),
        .dout(new_Jinkela_wire_16296)
    );

    bfr new_Jinkela_buffer_6696 (
        .din(new_Jinkela_wire_8419),
        .dout(new_Jinkela_wire_8420)
    );

    bfr new_Jinkela_buffer_6853 (
        .din(new_Jinkela_wire_8596),
        .dout(new_Jinkela_wire_8597)
    );

    bfr new_Jinkela_buffer_13641 (
        .din(new_Jinkela_wire_16296),
        .dout(new_Jinkela_wire_16297)
    );

    bfr new_Jinkela_buffer_6697 (
        .din(new_Jinkela_wire_8420),
        .dout(new_Jinkela_wire_8421)
    );

    bfr new_Jinkela_buffer_13735 (
        .din(new_Jinkela_wire_16396),
        .dout(new_Jinkela_wire_16397)
    );

    bfr new_Jinkela_buffer_6771 (
        .din(new_Jinkela_wire_8502),
        .dout(new_Jinkela_wire_8503)
    );

    bfr new_Jinkela_buffer_13642 (
        .din(new_Jinkela_wire_16297),
        .dout(new_Jinkela_wire_16298)
    );

    bfr new_Jinkela_buffer_6698 (
        .din(new_Jinkela_wire_8421),
        .dout(new_Jinkela_wire_8422)
    );

    bfr new_Jinkela_buffer_13782 (
        .din(new_Jinkela_wire_16447),
        .dout(new_Jinkela_wire_16448)
    );

    bfr new_Jinkela_buffer_13643 (
        .din(new_Jinkela_wire_16298),
        .dout(new_Jinkela_wire_16299)
    );

    bfr new_Jinkela_buffer_6699 (
        .din(new_Jinkela_wire_8422),
        .dout(new_Jinkela_wire_8423)
    );

    bfr new_Jinkela_buffer_13736 (
        .din(new_Jinkela_wire_16397),
        .dout(new_Jinkela_wire_16398)
    );

    bfr new_Jinkela_buffer_6772 (
        .din(new_Jinkela_wire_8503),
        .dout(new_Jinkela_wire_8504)
    );

    bfr new_Jinkela_buffer_13644 (
        .din(new_Jinkela_wire_16299),
        .dout(new_Jinkela_wire_16300)
    );

    bfr new_Jinkela_buffer_6700 (
        .din(new_Jinkela_wire_8423),
        .dout(new_Jinkela_wire_8424)
    );

    spl2 new_Jinkela_splitter_1185 (
        .a(_1548_),
        .b(new_Jinkela_wire_16516),
        .c(new_Jinkela_wire_16517)
    );

    bfr new_Jinkela_buffer_6854 (
        .din(new_Jinkela_wire_8597),
        .dout(new_Jinkela_wire_8598)
    );

    bfr new_Jinkela_buffer_13645 (
        .din(new_Jinkela_wire_16300),
        .dout(new_Jinkela_wire_16301)
    );

    bfr new_Jinkela_buffer_6701 (
        .din(new_Jinkela_wire_8424),
        .dout(new_Jinkela_wire_8425)
    );

    bfr new_Jinkela_buffer_13737 (
        .din(new_Jinkela_wire_16398),
        .dout(new_Jinkela_wire_16399)
    );

    bfr new_Jinkela_buffer_6773 (
        .din(new_Jinkela_wire_8504),
        .dout(new_Jinkela_wire_8505)
    );

    bfr new_Jinkela_buffer_13646 (
        .din(new_Jinkela_wire_16301),
        .dout(new_Jinkela_wire_16302)
    );

    bfr new_Jinkela_buffer_6702 (
        .din(new_Jinkela_wire_8425),
        .dout(new_Jinkela_wire_8426)
    );

    bfr new_Jinkela_buffer_13783 (
        .din(new_Jinkela_wire_16448),
        .dout(new_Jinkela_wire_16449)
    );

    spl2 new_Jinkela_splitter_727 (
        .a(_1001_),
        .b(new_Jinkela_wire_8760),
        .c(new_Jinkela_wire_8761)
    );

    bfr new_Jinkela_buffer_13647 (
        .din(new_Jinkela_wire_16302),
        .dout(new_Jinkela_wire_16303)
    );

    spl2 new_Jinkela_splitter_724 (
        .a(new_Jinkela_wire_8688),
        .b(new_Jinkela_wire_8689),
        .c(new_Jinkela_wire_8690)
    );

    bfr new_Jinkela_buffer_6703 (
        .din(new_Jinkela_wire_8426),
        .dout(new_Jinkela_wire_8427)
    );

    bfr new_Jinkela_buffer_13738 (
        .din(new_Jinkela_wire_16399),
        .dout(new_Jinkela_wire_16400)
    );

    bfr new_Jinkela_buffer_6774 (
        .din(new_Jinkela_wire_8505),
        .dout(new_Jinkela_wire_8506)
    );

    bfr new_Jinkela_buffer_13648 (
        .din(new_Jinkela_wire_16303),
        .dout(new_Jinkela_wire_16304)
    );

    bfr new_Jinkela_buffer_6704 (
        .din(new_Jinkela_wire_8427),
        .dout(new_Jinkela_wire_8428)
    );

    spl2 new_Jinkela_splitter_1186 (
        .a(_0743_),
        .b(new_Jinkela_wire_16522),
        .c(new_Jinkela_wire_16523)
    );

    bfr new_Jinkela_buffer_10220 (
        .din(new_Jinkela_wire_12383),
        .dout(new_Jinkela_wire_12384)
    );

    bfr new_Jinkela_buffer_17057 (
        .din(new_Jinkela_wire_20377),
        .dout(new_Jinkela_wire_20378)
    );

    bfr new_Jinkela_buffer_3377 (
        .din(new_Jinkela_wire_4506),
        .dout(new_Jinkela_wire_4507)
    );

    bfr new_Jinkela_buffer_10163 (
        .din(new_Jinkela_wire_12312),
        .dout(new_Jinkela_wire_12313)
    );

    spl2 new_Jinkela_splitter_1512 (
        .a(_1791_),
        .b(new_Jinkela_wire_20388),
        .c(new_Jinkela_wire_20389)
    );

    bfr new_Jinkela_buffer_3271 (
        .din(new_Jinkela_wire_4392),
        .dout(new_Jinkela_wire_4393)
    );

    bfr new_Jinkela_buffer_10455 (
        .din(new_Jinkela_wire_12632),
        .dout(new_Jinkela_wire_12633)
    );

    bfr new_Jinkela_buffer_17058 (
        .din(new_Jinkela_wire_20378),
        .dout(new_Jinkela_wire_20379)
    );

    bfr new_Jinkela_buffer_3418 (
        .din(new_Jinkela_wire_4551),
        .dout(new_Jinkela_wire_4552)
    );

    bfr new_Jinkela_buffer_10164 (
        .din(new_Jinkela_wire_12313),
        .dout(new_Jinkela_wire_12314)
    );

    bfr new_Jinkela_buffer_3272 (
        .din(new_Jinkela_wire_4393),
        .dout(new_Jinkela_wire_4394)
    );

    spl2 new_Jinkela_splitter_1511 (
        .a(_1471_),
        .b(new_Jinkela_wire_20386),
        .c(new_Jinkela_wire_20387)
    );

    bfr new_Jinkela_buffer_10221 (
        .din(new_Jinkela_wire_12384),
        .dout(new_Jinkela_wire_12385)
    );

    bfr new_Jinkela_buffer_17059 (
        .din(new_Jinkela_wire_20379),
        .dout(new_Jinkela_wire_20380)
    );

    bfr new_Jinkela_buffer_3378 (
        .din(new_Jinkela_wire_4507),
        .dout(new_Jinkela_wire_4508)
    );

    bfr new_Jinkela_buffer_10165 (
        .din(new_Jinkela_wire_12314),
        .dout(new_Jinkela_wire_12315)
    );

    bfr new_Jinkela_buffer_3273 (
        .din(new_Jinkela_wire_4394),
        .dout(new_Jinkela_wire_4395)
    );

    bfr new_Jinkela_buffer_10376 (
        .din(new_Jinkela_wire_12543),
        .dout(new_Jinkela_wire_12544)
    );

    spl2 new_Jinkela_splitter_1513 (
        .a(_1347_),
        .b(new_Jinkela_wire_20394),
        .c(new_Jinkela_wire_20395)
    );

    bfr new_Jinkela_buffer_3437 (
        .din(new_Jinkela_wire_4574),
        .dout(new_Jinkela_wire_4575)
    );

    bfr new_Jinkela_buffer_10166 (
        .din(new_Jinkela_wire_12315),
        .dout(new_Jinkela_wire_12316)
    );

    bfr new_Jinkela_buffer_17061 (
        .din(new_Jinkela_wire_20389),
        .dout(new_Jinkela_wire_20390)
    );

    bfr new_Jinkela_buffer_3274 (
        .din(new_Jinkela_wire_4395),
        .dout(new_Jinkela_wire_4396)
    );

    spl2 new_Jinkela_splitter_1514 (
        .a(_1129_),
        .b(new_Jinkela_wire_20396),
        .c(new_Jinkela_wire_20397)
    );

    bfr new_Jinkela_buffer_10222 (
        .din(new_Jinkela_wire_12385),
        .dout(new_Jinkela_wire_12386)
    );

    bfr new_Jinkela_buffer_3379 (
        .din(new_Jinkela_wire_4508),
        .dout(new_Jinkela_wire_4509)
    );

    bfr new_Jinkela_buffer_10167 (
        .din(new_Jinkela_wire_12316),
        .dout(new_Jinkela_wire_12317)
    );

    bfr new_Jinkela_buffer_17062 (
        .din(new_Jinkela_wire_20390),
        .dout(new_Jinkela_wire_20391)
    );

    bfr new_Jinkela_buffer_3275 (
        .din(new_Jinkela_wire_4396),
        .dout(new_Jinkela_wire_4397)
    );

    bfr new_Jinkela_buffer_10531 (
        .din(new_Jinkela_wire_12718),
        .dout(new_Jinkela_wire_12719)
    );

    spl2 new_Jinkela_splitter_1515 (
        .a(_1279_),
        .b(new_Jinkela_wire_20398),
        .c(new_Jinkela_wire_20399)
    );

    bfr new_Jinkela_buffer_3419 (
        .din(new_Jinkela_wire_4552),
        .dout(new_Jinkela_wire_4553)
    );

    bfr new_Jinkela_buffer_10168 (
        .din(new_Jinkela_wire_12317),
        .dout(new_Jinkela_wire_12318)
    );

    bfr new_Jinkela_buffer_17063 (
        .din(new_Jinkela_wire_20391),
        .dout(new_Jinkela_wire_20392)
    );

    bfr new_Jinkela_buffer_3276 (
        .din(new_Jinkela_wire_4397),
        .dout(new_Jinkela_wire_4398)
    );

    bfr new_Jinkela_buffer_10223 (
        .din(new_Jinkela_wire_12386),
        .dout(new_Jinkela_wire_12387)
    );

    bfr new_Jinkela_buffer_17209 (
        .din(_0348_),
        .dout(new_Jinkela_wire_20548)
    );

    bfr new_Jinkela_buffer_3380 (
        .din(new_Jinkela_wire_4509),
        .dout(new_Jinkela_wire_4510)
    );

    bfr new_Jinkela_buffer_17065 (
        .din(_0881_),
        .dout(new_Jinkela_wire_20400)
    );

    bfr new_Jinkela_buffer_10169 (
        .din(new_Jinkela_wire_12318),
        .dout(new_Jinkela_wire_12319)
    );

    bfr new_Jinkela_buffer_17064 (
        .din(new_Jinkela_wire_20392),
        .dout(new_Jinkela_wire_20393)
    );

    bfr new_Jinkela_buffer_3277 (
        .din(new_Jinkela_wire_4398),
        .dout(new_Jinkela_wire_4399)
    );

    bfr new_Jinkela_buffer_10377 (
        .din(new_Jinkela_wire_12544),
        .dout(new_Jinkela_wire_12545)
    );

    bfr new_Jinkela_buffer_17177 (
        .din(_0666_),
        .dout(new_Jinkela_wire_20514)
    );

    bfr new_Jinkela_buffer_3525 (
        .din(_0981_),
        .dout(new_Jinkela_wire_4669)
    );

    bfr new_Jinkela_buffer_10170 (
        .din(new_Jinkela_wire_12319),
        .dout(new_Jinkela_wire_12320)
    );

    bfr new_Jinkela_buffer_17066 (
        .din(new_Jinkela_wire_20400),
        .dout(new_Jinkela_wire_20401)
    );

    bfr new_Jinkela_buffer_3278 (
        .din(new_Jinkela_wire_4399),
        .dout(new_Jinkela_wire_4400)
    );

    bfr new_Jinkela_buffer_10224 (
        .din(new_Jinkela_wire_12387),
        .dout(new_Jinkela_wire_12388)
    );

    bfr new_Jinkela_buffer_3381 (
        .din(new_Jinkela_wire_4510),
        .dout(new_Jinkela_wire_4511)
    );

    spl2 new_Jinkela_splitter_1519 (
        .a(_1233_),
        .b(new_Jinkela_wire_20576),
        .c(new_Jinkela_wire_20577)
    );

    bfr new_Jinkela_buffer_10171 (
        .din(new_Jinkela_wire_12320),
        .dout(new_Jinkela_wire_12321)
    );

    bfr new_Jinkela_buffer_17067 (
        .din(new_Jinkela_wire_20401),
        .dout(new_Jinkela_wire_20402)
    );

    bfr new_Jinkela_buffer_3279 (
        .din(new_Jinkela_wire_4400),
        .dout(new_Jinkela_wire_4401)
    );

    bfr new_Jinkela_buffer_10456 (
        .din(new_Jinkela_wire_12633),
        .dout(new_Jinkela_wire_12634)
    );

    bfr new_Jinkela_buffer_17178 (
        .din(new_Jinkela_wire_20514),
        .dout(new_Jinkela_wire_20515)
    );

    bfr new_Jinkela_buffer_3420 (
        .din(new_Jinkela_wire_4553),
        .dout(new_Jinkela_wire_4554)
    );

    bfr new_Jinkela_buffer_10172 (
        .din(new_Jinkela_wire_12321),
        .dout(new_Jinkela_wire_12322)
    );

    bfr new_Jinkela_buffer_17068 (
        .din(new_Jinkela_wire_20402),
        .dout(new_Jinkela_wire_20403)
    );

    bfr new_Jinkela_buffer_3280 (
        .din(new_Jinkela_wire_4401),
        .dout(new_Jinkela_wire_4402)
    );

    bfr new_Jinkela_buffer_10225 (
        .din(new_Jinkela_wire_12388),
        .dout(new_Jinkela_wire_12389)
    );

    bfr new_Jinkela_buffer_3382 (
        .din(new_Jinkela_wire_4511),
        .dout(new_Jinkela_wire_4512)
    );

    bfr new_Jinkela_buffer_17235 (
        .din(_0634_),
        .dout(new_Jinkela_wire_20578)
    );

    bfr new_Jinkela_buffer_10173 (
        .din(new_Jinkela_wire_12322),
        .dout(new_Jinkela_wire_12323)
    );

    bfr new_Jinkela_buffer_17069 (
        .din(new_Jinkela_wire_20403),
        .dout(new_Jinkela_wire_20404)
    );

    bfr new_Jinkela_buffer_3281 (
        .din(new_Jinkela_wire_4402),
        .dout(new_Jinkela_wire_4403)
    );

    bfr new_Jinkela_buffer_10378 (
        .din(new_Jinkela_wire_12545),
        .dout(new_Jinkela_wire_12546)
    );

    bfr new_Jinkela_buffer_17179 (
        .din(new_Jinkela_wire_20515),
        .dout(new_Jinkela_wire_20516)
    );

    bfr new_Jinkela_buffer_3438 (
        .din(new_Jinkela_wire_4575),
        .dout(new_Jinkela_wire_4576)
    );

    bfr new_Jinkela_buffer_10174 (
        .din(new_Jinkela_wire_12323),
        .dout(new_Jinkela_wire_12324)
    );

    bfr new_Jinkela_buffer_17070 (
        .din(new_Jinkela_wire_20404),
        .dout(new_Jinkela_wire_20405)
    );

    bfr new_Jinkela_buffer_3282 (
        .din(new_Jinkela_wire_4403),
        .dout(new_Jinkela_wire_4404)
    );

    bfr new_Jinkela_buffer_10226 (
        .din(new_Jinkela_wire_12389),
        .dout(new_Jinkela_wire_12390)
    );

    bfr new_Jinkela_buffer_17210 (
        .din(new_Jinkela_wire_20548),
        .dout(new_Jinkela_wire_20549)
    );

    bfr new_Jinkela_buffer_3383 (
        .din(new_Jinkela_wire_4512),
        .dout(new_Jinkela_wire_4513)
    );

    bfr new_Jinkela_buffer_10175 (
        .din(new_Jinkela_wire_12324),
        .dout(new_Jinkela_wire_12325)
    );

    bfr new_Jinkela_buffer_17071 (
        .din(new_Jinkela_wire_20405),
        .dout(new_Jinkela_wire_20406)
    );

    bfr new_Jinkela_buffer_3283 (
        .din(new_Jinkela_wire_4404),
        .dout(new_Jinkela_wire_4405)
    );

    bfr new_Jinkela_buffer_17180 (
        .din(new_Jinkela_wire_20516),
        .dout(new_Jinkela_wire_20517)
    );

    bfr new_Jinkela_buffer_10536 (
        .din(_0208_),
        .dout(new_Jinkela_wire_12724)
    );

    bfr new_Jinkela_buffer_3421 (
        .din(new_Jinkela_wire_4554),
        .dout(new_Jinkela_wire_4555)
    );

    bfr new_Jinkela_buffer_10176 (
        .din(new_Jinkela_wire_12325),
        .dout(new_Jinkela_wire_12326)
    );

    bfr new_Jinkela_buffer_17072 (
        .din(new_Jinkela_wire_20406),
        .dout(new_Jinkela_wire_20407)
    );

    bfr new_Jinkela_buffer_3284 (
        .din(new_Jinkela_wire_4405),
        .dout(new_Jinkela_wire_4406)
    );

    bfr new_Jinkela_buffer_10227 (
        .din(new_Jinkela_wire_12390),
        .dout(new_Jinkela_wire_12391)
    );

    bfr new_Jinkela_buffer_17306 (
        .din(new_net_3946),
        .dout(new_Jinkela_wire_20653)
    );

    bfr new_Jinkela_buffer_3384 (
        .din(new_Jinkela_wire_4513),
        .dout(new_Jinkela_wire_4514)
    );

    spl2 new_Jinkela_splitter_924 (
        .a(new_Jinkela_wire_12326),
        .b(new_Jinkela_wire_12327),
        .c(new_Jinkela_wire_12328)
    );

    bfr new_Jinkela_buffer_17073 (
        .din(new_Jinkela_wire_20407),
        .dout(new_Jinkela_wire_20408)
    );

    bfr new_Jinkela_buffer_3285 (
        .din(new_Jinkela_wire_4406),
        .dout(new_Jinkela_wire_4407)
    );

    bfr new_Jinkela_buffer_10228 (
        .din(new_Jinkela_wire_12391),
        .dout(new_Jinkela_wire_12392)
    );

    bfr new_Jinkela_buffer_17181 (
        .din(new_Jinkela_wire_20517),
        .dout(new_Jinkela_wire_20518)
    );

    bfr new_Jinkela_buffer_10379 (
        .din(new_Jinkela_wire_12546),
        .dout(new_Jinkela_wire_12547)
    );

    bfr new_Jinkela_buffer_17074 (
        .din(new_Jinkela_wire_20408),
        .dout(new_Jinkela_wire_20409)
    );

    bfr new_Jinkela_buffer_3286 (
        .din(new_Jinkela_wire_4407),
        .dout(new_Jinkela_wire_4408)
    );

    bfr new_Jinkela_buffer_10457 (
        .din(new_Jinkela_wire_12634),
        .dout(new_Jinkela_wire_12635)
    );

    bfr new_Jinkela_buffer_17211 (
        .din(new_Jinkela_wire_20549),
        .dout(new_Jinkela_wire_20550)
    );

    bfr new_Jinkela_buffer_3385 (
        .din(new_Jinkela_wire_4514),
        .dout(new_Jinkela_wire_4515)
    );

    bfr new_Jinkela_buffer_10229 (
        .din(new_Jinkela_wire_12392),
        .dout(new_Jinkela_wire_12393)
    );

    bfr new_Jinkela_buffer_17075 (
        .din(new_Jinkela_wire_20409),
        .dout(new_Jinkela_wire_20410)
    );

    bfr new_Jinkela_buffer_3287 (
        .din(new_Jinkela_wire_4408),
        .dout(new_Jinkela_wire_4409)
    );

    bfr new_Jinkela_buffer_10380 (
        .din(new_Jinkela_wire_12547),
        .dout(new_Jinkela_wire_12548)
    );

    bfr new_Jinkela_buffer_17182 (
        .din(new_Jinkela_wire_20518),
        .dout(new_Jinkela_wire_20519)
    );

    spl2 new_Jinkela_splitter_420 (
        .a(_1752_),
        .b(new_Jinkela_wire_4667),
        .c(new_Jinkela_wire_4668)
    );

    bfr new_Jinkela_buffer_3422 (
        .din(new_Jinkela_wire_4555),
        .dout(new_Jinkela_wire_4556)
    );

    bfr new_Jinkela_buffer_10230 (
        .din(new_Jinkela_wire_12393),
        .dout(new_Jinkela_wire_12394)
    );

    bfr new_Jinkela_buffer_17076 (
        .din(new_Jinkela_wire_20410),
        .dout(new_Jinkela_wire_20411)
    );

    bfr new_Jinkela_buffer_3288 (
        .din(new_Jinkela_wire_4409),
        .dout(new_Jinkela_wire_4410)
    );

    bfr new_Jinkela_buffer_3386 (
        .din(new_Jinkela_wire_4515),
        .dout(new_Jinkela_wire_4516)
    );

    bfr new_Jinkela_buffer_10537 (
        .din(_0467_),
        .dout(new_Jinkela_wire_12725)
    );

    bfr new_Jinkela_buffer_17281 (
        .din(_1078_),
        .dout(new_Jinkela_wire_20626)
    );

    bfr new_Jinkela_buffer_10231 (
        .din(new_Jinkela_wire_12394),
        .dout(new_Jinkela_wire_12395)
    );

    bfr new_Jinkela_buffer_17077 (
        .din(new_Jinkela_wire_20411),
        .dout(new_Jinkela_wire_20412)
    );

    bfr new_Jinkela_buffer_3289 (
        .din(new_Jinkela_wire_4410),
        .dout(new_Jinkela_wire_4411)
    );

    bfr new_Jinkela_buffer_10381 (
        .din(new_Jinkela_wire_12548),
        .dout(new_Jinkela_wire_12549)
    );

    bfr new_Jinkela_buffer_17183 (
        .din(new_Jinkela_wire_20519),
        .dout(new_Jinkela_wire_20520)
    );

    bfr new_Jinkela_buffer_3439 (
        .din(new_Jinkela_wire_4576),
        .dout(new_Jinkela_wire_4577)
    );

    bfr new_Jinkela_buffer_10232 (
        .din(new_Jinkela_wire_12395),
        .dout(new_Jinkela_wire_12396)
    );

    bfr new_Jinkela_buffer_17078 (
        .din(new_Jinkela_wire_20412),
        .dout(new_Jinkela_wire_20413)
    );

    bfr new_Jinkela_buffer_3290 (
        .din(new_Jinkela_wire_4411),
        .dout(new_Jinkela_wire_4412)
    );

    bfr new_Jinkela_buffer_10458 (
        .din(new_Jinkela_wire_12635),
        .dout(new_Jinkela_wire_12636)
    );

    bfr new_Jinkela_buffer_17212 (
        .din(new_Jinkela_wire_20550),
        .dout(new_Jinkela_wire_20551)
    );

    bfr new_Jinkela_buffer_3387 (
        .din(new_Jinkela_wire_4516),
        .dout(new_Jinkela_wire_4517)
    );

    bfr new_Jinkela_buffer_10233 (
        .din(new_Jinkela_wire_12396),
        .dout(new_Jinkela_wire_12397)
    );

    bfr new_Jinkela_buffer_17079 (
        .din(new_Jinkela_wire_20413),
        .dout(new_Jinkela_wire_20414)
    );

    bfr new_Jinkela_buffer_3291 (
        .din(new_Jinkela_wire_4412),
        .dout(new_Jinkela_wire_4413)
    );

    bfr new_Jinkela_buffer_6855 (
        .din(new_Jinkela_wire_8598),
        .dout(new_Jinkela_wire_8599)
    );

    bfr new_Jinkela_buffer_6705 (
        .din(new_Jinkela_wire_8428),
        .dout(new_Jinkela_wire_8429)
    );

    bfr new_Jinkela_buffer_6775 (
        .din(new_Jinkela_wire_8506),
        .dout(new_Jinkela_wire_8507)
    );

    bfr new_Jinkela_buffer_6706 (
        .din(new_Jinkela_wire_8429),
        .dout(new_Jinkela_wire_8430)
    );

    spl2 new_Jinkela_splitter_728 (
        .a(_1063_),
        .b(new_Jinkela_wire_8762),
        .c(new_Jinkela_wire_8763)
    );

    bfr new_Jinkela_buffer_6707 (
        .din(new_Jinkela_wire_8430),
        .dout(new_Jinkela_wire_8431)
    );

    bfr new_Jinkela_buffer_6776 (
        .din(new_Jinkela_wire_8507),
        .dout(new_Jinkela_wire_8508)
    );

    bfr new_Jinkela_buffer_6708 (
        .din(new_Jinkela_wire_8431),
        .dout(new_Jinkela_wire_8432)
    );

    bfr new_Jinkela_buffer_6856 (
        .din(new_Jinkela_wire_8599),
        .dout(new_Jinkela_wire_8600)
    );

    bfr new_Jinkela_buffer_6709 (
        .din(new_Jinkela_wire_8432),
        .dout(new_Jinkela_wire_8433)
    );

    bfr new_Jinkela_buffer_6777 (
        .din(new_Jinkela_wire_8508),
        .dout(new_Jinkela_wire_8509)
    );

    bfr new_Jinkela_buffer_6710 (
        .din(new_Jinkela_wire_8433),
        .dout(new_Jinkela_wire_8434)
    );

    bfr new_Jinkela_buffer_6941 (
        .din(new_Jinkela_wire_8694),
        .dout(new_Jinkela_wire_8695)
    );

    bfr new_Jinkela_buffer_6711 (
        .din(new_Jinkela_wire_8434),
        .dout(new_Jinkela_wire_8435)
    );

    bfr new_Jinkela_buffer_6778 (
        .din(new_Jinkela_wire_8509),
        .dout(new_Jinkela_wire_8510)
    );

    bfr new_Jinkela_buffer_6712 (
        .din(new_Jinkela_wire_8435),
        .dout(new_Jinkela_wire_8436)
    );

    bfr new_Jinkela_buffer_6857 (
        .din(new_Jinkela_wire_8600),
        .dout(new_Jinkela_wire_8601)
    );

    bfr new_Jinkela_buffer_6713 (
        .din(new_Jinkela_wire_8436),
        .dout(new_Jinkela_wire_8437)
    );

    bfr new_Jinkela_buffer_6779 (
        .din(new_Jinkela_wire_8510),
        .dout(new_Jinkela_wire_8511)
    );

    bfr new_Jinkela_buffer_6714 (
        .din(new_Jinkela_wire_8437),
        .dout(new_Jinkela_wire_8438)
    );

    bfr new_Jinkela_buffer_6715 (
        .din(new_Jinkela_wire_8438),
        .dout(new_Jinkela_wire_8439)
    );

    bfr new_Jinkela_buffer_6780 (
        .din(new_Jinkela_wire_8511),
        .dout(new_Jinkela_wire_8512)
    );

    bfr new_Jinkela_buffer_6716 (
        .din(new_Jinkela_wire_8439),
        .dout(new_Jinkela_wire_8440)
    );

    bfr new_Jinkela_buffer_6858 (
        .din(new_Jinkela_wire_8601),
        .dout(new_Jinkela_wire_8602)
    );

    bfr new_Jinkela_buffer_6717 (
        .din(new_Jinkela_wire_8440),
        .dout(new_Jinkela_wire_8441)
    );

    bfr new_Jinkela_buffer_6781 (
        .din(new_Jinkela_wire_8512),
        .dout(new_Jinkela_wire_8513)
    );

    bfr new_Jinkela_buffer_6718 (
        .din(new_Jinkela_wire_8441),
        .dout(new_Jinkela_wire_8442)
    );

    spl2 new_Jinkela_splitter_729 (
        .a(_0190_),
        .b(new_Jinkela_wire_8764),
        .c(new_Jinkela_wire_8765)
    );

    bfr new_Jinkela_buffer_6719 (
        .din(new_Jinkela_wire_8442),
        .dout(new_Jinkela_wire_8443)
    );

    bfr new_Jinkela_buffer_6782 (
        .din(new_Jinkela_wire_8513),
        .dout(new_Jinkela_wire_8514)
    );

    bfr new_Jinkela_buffer_6720 (
        .din(new_Jinkela_wire_8443),
        .dout(new_Jinkela_wire_8444)
    );

    bfr new_Jinkela_buffer_6859 (
        .din(new_Jinkela_wire_8602),
        .dout(new_Jinkela_wire_8603)
    );

    bfr new_Jinkela_buffer_6721 (
        .din(new_Jinkela_wire_8444),
        .dout(new_Jinkela_wire_8445)
    );

    bfr new_Jinkela_buffer_6783 (
        .din(new_Jinkela_wire_8514),
        .dout(new_Jinkela_wire_8515)
    );

    bfr new_Jinkela_buffer_6722 (
        .din(new_Jinkela_wire_8445),
        .dout(new_Jinkela_wire_8446)
    );

    bfr new_Jinkela_buffer_6942 (
        .din(new_Jinkela_wire_8695),
        .dout(new_Jinkela_wire_8696)
    );

    bfr new_Jinkela_buffer_6723 (
        .din(new_Jinkela_wire_8446),
        .dout(new_Jinkela_wire_8447)
    );

    bfr new_Jinkela_buffer_6784 (
        .din(new_Jinkela_wire_8515),
        .dout(new_Jinkela_wire_8516)
    );

    bfr new_Jinkela_buffer_6724 (
        .din(new_Jinkela_wire_8447),
        .dout(new_Jinkela_wire_8448)
    );

    bfr new_Jinkela_buffer_6860 (
        .din(new_Jinkela_wire_8603),
        .dout(new_Jinkela_wire_8604)
    );

    bfr new_Jinkela_buffer_6725 (
        .din(new_Jinkela_wire_8448),
        .dout(new_Jinkela_wire_8449)
    );

    bfr new_Jinkela_buffer_13649 (
        .din(new_Jinkela_wire_16304),
        .dout(new_Jinkela_wire_16305)
    );

    bfr new_Jinkela_buffer_13739 (
        .din(new_Jinkela_wire_16400),
        .dout(new_Jinkela_wire_16401)
    );

    bfr new_Jinkela_buffer_13650 (
        .din(new_Jinkela_wire_16305),
        .dout(new_Jinkela_wire_16306)
    );

    bfr new_Jinkela_buffer_13784 (
        .din(new_Jinkela_wire_16449),
        .dout(new_Jinkela_wire_16450)
    );

    bfr new_Jinkela_buffer_13651 (
        .din(new_Jinkela_wire_16306),
        .dout(new_Jinkela_wire_16307)
    );

    bfr new_Jinkela_buffer_13740 (
        .din(new_Jinkela_wire_16401),
        .dout(new_Jinkela_wire_16402)
    );

    bfr new_Jinkela_buffer_13652 (
        .din(new_Jinkela_wire_16307),
        .dout(new_Jinkela_wire_16308)
    );

    spl2 new_Jinkela_splitter_1187 (
        .a(_0733_),
        .b(new_Jinkela_wire_16524),
        .c(new_Jinkela_wire_16525)
    );

    bfr new_Jinkela_buffer_13653 (
        .din(new_Jinkela_wire_16308),
        .dout(new_Jinkela_wire_16309)
    );

    bfr new_Jinkela_buffer_13741 (
        .din(new_Jinkela_wire_16402),
        .dout(new_Jinkela_wire_16403)
    );

    bfr new_Jinkela_buffer_13654 (
        .din(new_Jinkela_wire_16309),
        .dout(new_Jinkela_wire_16310)
    );

    bfr new_Jinkela_buffer_13785 (
        .din(new_Jinkela_wire_16450),
        .dout(new_Jinkela_wire_16451)
    );

    bfr new_Jinkela_buffer_13655 (
        .din(new_Jinkela_wire_16310),
        .dout(new_Jinkela_wire_16311)
    );

    bfr new_Jinkela_buffer_13742 (
        .din(new_Jinkela_wire_16403),
        .dout(new_Jinkela_wire_16404)
    );

    bfr new_Jinkela_buffer_13656 (
        .din(new_Jinkela_wire_16311),
        .dout(new_Jinkela_wire_16312)
    );

    bfr new_Jinkela_buffer_13848 (
        .din(new_Jinkela_wire_16525),
        .dout(new_Jinkela_wire_16526)
    );

    bfr new_Jinkela_buffer_13657 (
        .din(new_Jinkela_wire_16312),
        .dout(new_Jinkela_wire_16313)
    );

    bfr new_Jinkela_buffer_13743 (
        .din(new_Jinkela_wire_16404),
        .dout(new_Jinkela_wire_16405)
    );

    bfr new_Jinkela_buffer_13658 (
        .din(new_Jinkela_wire_16313),
        .dout(new_Jinkela_wire_16314)
    );

    bfr new_Jinkela_buffer_13786 (
        .din(new_Jinkela_wire_16451),
        .dout(new_Jinkela_wire_16452)
    );

    bfr new_Jinkela_buffer_13659 (
        .din(new_Jinkela_wire_16314),
        .dout(new_Jinkela_wire_16315)
    );

    bfr new_Jinkela_buffer_13744 (
        .din(new_Jinkela_wire_16405),
        .dout(new_Jinkela_wire_16406)
    );

    bfr new_Jinkela_buffer_13660 (
        .din(new_Jinkela_wire_16315),
        .dout(new_Jinkela_wire_16316)
    );

    bfr new_Jinkela_buffer_13845 (
        .din(new_Jinkela_wire_16518),
        .dout(new_Jinkela_wire_16519)
    );

    bfr new_Jinkela_buffer_13661 (
        .din(new_Jinkela_wire_16316),
        .dout(new_Jinkela_wire_16317)
    );

    bfr new_Jinkela_buffer_13745 (
        .din(new_Jinkela_wire_16406),
        .dout(new_Jinkela_wire_16407)
    );

    bfr new_Jinkela_buffer_13662 (
        .din(new_Jinkela_wire_16317),
        .dout(new_Jinkela_wire_16318)
    );

    bfr new_Jinkela_buffer_13787 (
        .din(new_Jinkela_wire_16452),
        .dout(new_Jinkela_wire_16453)
    );

    bfr new_Jinkela_buffer_13663 (
        .din(new_Jinkela_wire_16318),
        .dout(new_Jinkela_wire_16319)
    );

    bfr new_Jinkela_buffer_13746 (
        .din(new_Jinkela_wire_16407),
        .dout(new_Jinkela_wire_16408)
    );

    bfr new_Jinkela_buffer_13664 (
        .din(new_Jinkela_wire_16319),
        .dout(new_Jinkela_wire_16320)
    );

    spl2 new_Jinkela_splitter_1188 (
        .a(_0035_),
        .b(new_Jinkela_wire_16530),
        .c(new_Jinkela_wire_16531)
    );

    bfr new_Jinkela_buffer_13665 (
        .din(new_Jinkela_wire_16320),
        .dout(new_Jinkela_wire_16321)
    );

    bfr new_Jinkela_buffer_13747 (
        .din(new_Jinkela_wire_16408),
        .dout(new_Jinkela_wire_16409)
    );

    bfr new_Jinkela_buffer_13666 (
        .din(new_Jinkela_wire_16321),
        .dout(new_Jinkela_wire_16322)
    );

    bfr new_Jinkela_buffer_13788 (
        .din(new_Jinkela_wire_16453),
        .dout(new_Jinkela_wire_16454)
    );

    bfr new_Jinkela_buffer_13667 (
        .din(new_Jinkela_wire_16322),
        .dout(new_Jinkela_wire_16323)
    );

    bfr new_Jinkela_buffer_13748 (
        .din(new_Jinkela_wire_16409),
        .dout(new_Jinkela_wire_16410)
    );

    bfr new_Jinkela_buffer_13668 (
        .din(new_Jinkela_wire_16323),
        .dout(new_Jinkela_wire_16324)
    );

    bfr new_Jinkela_buffer_13846 (
        .din(new_Jinkela_wire_16519),
        .dout(new_Jinkela_wire_16520)
    );

    bfr new_Jinkela_buffer_13669 (
        .din(new_Jinkela_wire_16324),
        .dout(new_Jinkela_wire_16325)
    );

    bfr new_Jinkela_buffer_13749 (
        .din(new_Jinkela_wire_16410),
        .dout(new_Jinkela_wire_16411)
    );

    bfr new_Jinkela_buffer_17184 (
        .din(new_Jinkela_wire_20520),
        .dout(new_Jinkela_wire_20521)
    );

    bfr new_Jinkela_buffer_17080 (
        .din(new_Jinkela_wire_20414),
        .dout(new_Jinkela_wire_20415)
    );

    bfr new_Jinkela_buffer_3423 (
        .din(new_Jinkela_wire_4556),
        .dout(new_Jinkela_wire_4557)
    );

    bfr new_Jinkela_buffer_3292 (
        .din(new_Jinkela_wire_4413),
        .dout(new_Jinkela_wire_4414)
    );

    bfr new_Jinkela_buffer_17236 (
        .din(new_Jinkela_wire_20578),
        .dout(new_Jinkela_wire_20579)
    );

    bfr new_Jinkela_buffer_3388 (
        .din(new_Jinkela_wire_4517),
        .dout(new_Jinkela_wire_4518)
    );

    bfr new_Jinkela_buffer_17081 (
        .din(new_Jinkela_wire_20415),
        .dout(new_Jinkela_wire_20416)
    );

    bfr new_Jinkela_buffer_3293 (
        .din(new_Jinkela_wire_4414),
        .dout(new_Jinkela_wire_4415)
    );

    bfr new_Jinkela_buffer_17185 (
        .din(new_Jinkela_wire_20521),
        .dout(new_Jinkela_wire_20522)
    );

    bfr new_Jinkela_buffer_17082 (
        .din(new_Jinkela_wire_20416),
        .dout(new_Jinkela_wire_20417)
    );

    bfr new_Jinkela_buffer_3294 (
        .din(new_Jinkela_wire_4415),
        .dout(new_Jinkela_wire_4416)
    );

    bfr new_Jinkela_buffer_17213 (
        .din(new_Jinkela_wire_20551),
        .dout(new_Jinkela_wire_20552)
    );

    bfr new_Jinkela_buffer_3389 (
        .din(new_Jinkela_wire_4518),
        .dout(new_Jinkela_wire_4519)
    );

    bfr new_Jinkela_buffer_17083 (
        .din(new_Jinkela_wire_20417),
        .dout(new_Jinkela_wire_20418)
    );

    bfr new_Jinkela_buffer_3295 (
        .din(new_Jinkela_wire_4416),
        .dout(new_Jinkela_wire_4417)
    );

    bfr new_Jinkela_buffer_17186 (
        .din(new_Jinkela_wire_20522),
        .dout(new_Jinkela_wire_20523)
    );

    spl2 new_Jinkela_splitter_421 (
        .a(_0274_),
        .b(new_Jinkela_wire_4671),
        .c(new_Jinkela_wire_4672)
    );

    bfr new_Jinkela_buffer_17084 (
        .din(new_Jinkela_wire_20418),
        .dout(new_Jinkela_wire_20419)
    );

    bfr new_Jinkela_buffer_3424 (
        .din(new_Jinkela_wire_4557),
        .dout(new_Jinkela_wire_4558)
    );

    bfr new_Jinkela_buffer_3296 (
        .din(new_Jinkela_wire_4417),
        .dout(new_Jinkela_wire_4418)
    );

    bfr new_Jinkela_buffer_3390 (
        .din(new_Jinkela_wire_4519),
        .dout(new_Jinkela_wire_4520)
    );

    spl2 new_Jinkela_splitter_1522 (
        .a(_0726_),
        .b(new_Jinkela_wire_20677),
        .c(new_Jinkela_wire_20678)
    );

    bfr new_Jinkela_buffer_17085 (
        .din(new_Jinkela_wire_20419),
        .dout(new_Jinkela_wire_20420)
    );

    bfr new_Jinkela_buffer_3297 (
        .din(new_Jinkela_wire_4418),
        .dout(new_Jinkela_wire_4419)
    );

    bfr new_Jinkela_buffer_17187 (
        .din(new_Jinkela_wire_20523),
        .dout(new_Jinkela_wire_20524)
    );

    bfr new_Jinkela_buffer_17086 (
        .din(new_Jinkela_wire_20420),
        .dout(new_Jinkela_wire_20421)
    );

    bfr new_Jinkela_buffer_3440 (
        .din(new_Jinkela_wire_4577),
        .dout(new_Jinkela_wire_4578)
    );

    bfr new_Jinkela_buffer_3298 (
        .din(new_Jinkela_wire_4419),
        .dout(new_Jinkela_wire_4420)
    );

    bfr new_Jinkela_buffer_17214 (
        .din(new_Jinkela_wire_20552),
        .dout(new_Jinkela_wire_20553)
    );

    bfr new_Jinkela_buffer_3391 (
        .din(new_Jinkela_wire_4520),
        .dout(new_Jinkela_wire_4521)
    );

    bfr new_Jinkela_buffer_17087 (
        .din(new_Jinkela_wire_20421),
        .dout(new_Jinkela_wire_20422)
    );

    bfr new_Jinkela_buffer_3299 (
        .din(new_Jinkela_wire_4420),
        .dout(new_Jinkela_wire_4421)
    );

    bfr new_Jinkela_buffer_17188 (
        .din(new_Jinkela_wire_20524),
        .dout(new_Jinkela_wire_20525)
    );

    bfr new_Jinkela_buffer_17088 (
        .din(new_Jinkela_wire_20422),
        .dout(new_Jinkela_wire_20423)
    );

    bfr new_Jinkela_buffer_3425 (
        .din(new_Jinkela_wire_4558),
        .dout(new_Jinkela_wire_4559)
    );

    bfr new_Jinkela_buffer_3300 (
        .din(new_Jinkela_wire_4421),
        .dout(new_Jinkela_wire_4422)
    );

    bfr new_Jinkela_buffer_17237 (
        .din(new_Jinkela_wire_20579),
        .dout(new_Jinkela_wire_20580)
    );

    bfr new_Jinkela_buffer_3392 (
        .din(new_Jinkela_wire_4521),
        .dout(new_Jinkela_wire_4522)
    );

    bfr new_Jinkela_buffer_17089 (
        .din(new_Jinkela_wire_20423),
        .dout(new_Jinkela_wire_20424)
    );

    bfr new_Jinkela_buffer_3301 (
        .din(new_Jinkela_wire_4422),
        .dout(new_Jinkela_wire_4423)
    );

    bfr new_Jinkela_buffer_17189 (
        .din(new_Jinkela_wire_20525),
        .dout(new_Jinkela_wire_20526)
    );

    bfr new_Jinkela_buffer_17090 (
        .din(new_Jinkela_wire_20424),
        .dout(new_Jinkela_wire_20425)
    );

    bfr new_Jinkela_buffer_3302 (
        .din(new_Jinkela_wire_4423),
        .dout(new_Jinkela_wire_4424)
    );

    bfr new_Jinkela_buffer_17215 (
        .din(new_Jinkela_wire_20553),
        .dout(new_Jinkela_wire_20554)
    );

    bfr new_Jinkela_buffer_3393 (
        .din(new_Jinkela_wire_4522),
        .dout(new_Jinkela_wire_4523)
    );

    bfr new_Jinkela_buffer_17091 (
        .din(new_Jinkela_wire_20425),
        .dout(new_Jinkela_wire_20426)
    );

    bfr new_Jinkela_buffer_3303 (
        .din(new_Jinkela_wire_4424),
        .dout(new_Jinkela_wire_4425)
    );

    bfr new_Jinkela_buffer_17190 (
        .din(new_Jinkela_wire_20526),
        .dout(new_Jinkela_wire_20527)
    );

    bfr new_Jinkela_buffer_3526 (
        .din(_0363_),
        .dout(new_Jinkela_wire_4670)
    );

    bfr new_Jinkela_buffer_17092 (
        .din(new_Jinkela_wire_20426),
        .dout(new_Jinkela_wire_20427)
    );

    bfr new_Jinkela_buffer_3426 (
        .din(new_Jinkela_wire_4559),
        .dout(new_Jinkela_wire_4560)
    );

    bfr new_Jinkela_buffer_3304 (
        .din(new_Jinkela_wire_4425),
        .dout(new_Jinkela_wire_4426)
    );

    bfr new_Jinkela_buffer_17282 (
        .din(new_Jinkela_wire_20626),
        .dout(new_Jinkela_wire_20627)
    );

    bfr new_Jinkela_buffer_3394 (
        .din(new_Jinkela_wire_4523),
        .dout(new_Jinkela_wire_4524)
    );

    bfr new_Jinkela_buffer_17093 (
        .din(new_Jinkela_wire_20427),
        .dout(new_Jinkela_wire_20428)
    );

    bfr new_Jinkela_buffer_3305 (
        .din(new_Jinkela_wire_4426),
        .dout(new_Jinkela_wire_4427)
    );

    bfr new_Jinkela_buffer_17191 (
        .din(new_Jinkela_wire_20527),
        .dout(new_Jinkela_wire_20528)
    );

    bfr new_Jinkela_buffer_17094 (
        .din(new_Jinkela_wire_20428),
        .dout(new_Jinkela_wire_20429)
    );

    bfr new_Jinkela_buffer_3441 (
        .din(new_Jinkela_wire_4578),
        .dout(new_Jinkela_wire_4579)
    );

    bfr new_Jinkela_buffer_3306 (
        .din(new_Jinkela_wire_4427),
        .dout(new_Jinkela_wire_4428)
    );

    bfr new_Jinkela_buffer_17216 (
        .din(new_Jinkela_wire_20554),
        .dout(new_Jinkela_wire_20555)
    );

    bfr new_Jinkela_buffer_3395 (
        .din(new_Jinkela_wire_4524),
        .dout(new_Jinkela_wire_4525)
    );

    bfr new_Jinkela_buffer_17095 (
        .din(new_Jinkela_wire_20429),
        .dout(new_Jinkela_wire_20430)
    );

    bfr new_Jinkela_buffer_3307 (
        .din(new_Jinkela_wire_4428),
        .dout(new_Jinkela_wire_4429)
    );

    bfr new_Jinkela_buffer_17192 (
        .din(new_Jinkela_wire_20528),
        .dout(new_Jinkela_wire_20529)
    );

    bfr new_Jinkela_buffer_17096 (
        .din(new_Jinkela_wire_20430),
        .dout(new_Jinkela_wire_20431)
    );

    bfr new_Jinkela_buffer_3427 (
        .din(new_Jinkela_wire_4560),
        .dout(new_Jinkela_wire_4561)
    );

    bfr new_Jinkela_buffer_3308 (
        .din(new_Jinkela_wire_4429),
        .dout(new_Jinkela_wire_4430)
    );

    bfr new_Jinkela_buffer_17238 (
        .din(new_Jinkela_wire_20580),
        .dout(new_Jinkela_wire_20581)
    );

    bfr new_Jinkela_buffer_3396 (
        .din(new_Jinkela_wire_4525),
        .dout(new_Jinkela_wire_4526)
    );

    bfr new_Jinkela_buffer_17097 (
        .din(new_Jinkela_wire_20431),
        .dout(new_Jinkela_wire_20432)
    );

    bfr new_Jinkela_buffer_3309 (
        .din(new_Jinkela_wire_4430),
        .dout(new_Jinkela_wire_4431)
    );

    bfr new_Jinkela_buffer_17193 (
        .din(new_Jinkela_wire_20529),
        .dout(new_Jinkela_wire_20530)
    );

    bfr new_Jinkela_buffer_17098 (
        .din(new_Jinkela_wire_20432),
        .dout(new_Jinkela_wire_20433)
    );

    spl2 new_Jinkela_splitter_422 (
        .a(_0414_),
        .b(new_Jinkela_wire_4673),
        .c(new_Jinkela_wire_4674)
    );

    bfr new_Jinkela_buffer_3310 (
        .din(new_Jinkela_wire_4431),
        .dout(new_Jinkela_wire_4432)
    );

    bfr new_Jinkela_buffer_17217 (
        .din(new_Jinkela_wire_20555),
        .dout(new_Jinkela_wire_20556)
    );

    bfr new_Jinkela_buffer_3397 (
        .din(new_Jinkela_wire_4526),
        .dout(new_Jinkela_wire_4527)
    );

    bfr new_Jinkela_buffer_17099 (
        .din(new_Jinkela_wire_20433),
        .dout(new_Jinkela_wire_20434)
    );

    bfr new_Jinkela_buffer_3311 (
        .din(new_Jinkela_wire_4432),
        .dout(new_Jinkela_wire_4433)
    );

    bfr new_Jinkela_buffer_17194 (
        .din(new_Jinkela_wire_20530),
        .dout(new_Jinkela_wire_20531)
    );

    bfr new_Jinkela_buffer_17100 (
        .din(new_Jinkela_wire_20434),
        .dout(new_Jinkela_wire_20435)
    );

    bfr new_Jinkela_buffer_3428 (
        .din(new_Jinkela_wire_4561),
        .dout(new_Jinkela_wire_4562)
    );

    bfr new_Jinkela_buffer_3312 (
        .din(new_Jinkela_wire_4433),
        .dout(new_Jinkela_wire_4434)
    );

    bfr new_Jinkela_buffer_6785 (
        .din(new_Jinkela_wire_8516),
        .dout(new_Jinkela_wire_8517)
    );

    bfr new_Jinkela_buffer_6726 (
        .din(new_Jinkela_wire_8449),
        .dout(new_Jinkela_wire_8450)
    );

    spl2 new_Jinkela_splitter_731 (
        .a(_1450_),
        .b(new_Jinkela_wire_8839),
        .c(new_Jinkela_wire_8840)
    );

    bfr new_Jinkela_buffer_6727 (
        .din(new_Jinkela_wire_8450),
        .dout(new_Jinkela_wire_8451)
    );

    bfr new_Jinkela_buffer_6786 (
        .din(new_Jinkela_wire_8517),
        .dout(new_Jinkela_wire_8518)
    );

    bfr new_Jinkela_buffer_6728 (
        .din(new_Jinkela_wire_8451),
        .dout(new_Jinkela_wire_8452)
    );

    bfr new_Jinkela_buffer_6861 (
        .din(new_Jinkela_wire_8604),
        .dout(new_Jinkela_wire_8605)
    );

    bfr new_Jinkela_buffer_6729 (
        .din(new_Jinkela_wire_8452),
        .dout(new_Jinkela_wire_8453)
    );

    bfr new_Jinkela_buffer_6787 (
        .din(new_Jinkela_wire_8518),
        .dout(new_Jinkela_wire_8519)
    );

    bfr new_Jinkela_buffer_6730 (
        .din(new_Jinkela_wire_8453),
        .dout(new_Jinkela_wire_8454)
    );

    bfr new_Jinkela_buffer_6943 (
        .din(new_Jinkela_wire_8696),
        .dout(new_Jinkela_wire_8697)
    );

    bfr new_Jinkela_buffer_6731 (
        .din(new_Jinkela_wire_8454),
        .dout(new_Jinkela_wire_8455)
    );

    bfr new_Jinkela_buffer_6788 (
        .din(new_Jinkela_wire_8519),
        .dout(new_Jinkela_wire_8520)
    );

    bfr new_Jinkela_buffer_6732 (
        .din(new_Jinkela_wire_8455),
        .dout(new_Jinkela_wire_8456)
    );

    bfr new_Jinkela_buffer_6862 (
        .din(new_Jinkela_wire_8605),
        .dout(new_Jinkela_wire_8606)
    );

    bfr new_Jinkela_buffer_6733 (
        .din(new_Jinkela_wire_8456),
        .dout(new_Jinkela_wire_8457)
    );

    bfr new_Jinkela_buffer_6789 (
        .din(new_Jinkela_wire_8520),
        .dout(new_Jinkela_wire_8521)
    );

    bfr new_Jinkela_buffer_6734 (
        .din(new_Jinkela_wire_8457),
        .dout(new_Jinkela_wire_8458)
    );

    bfr new_Jinkela_buffer_7004 (
        .din(_0838_),
        .dout(new_Jinkela_wire_8766)
    );

    bfr new_Jinkela_buffer_6735 (
        .din(new_Jinkela_wire_8458),
        .dout(new_Jinkela_wire_8459)
    );

    bfr new_Jinkela_buffer_6790 (
        .din(new_Jinkela_wire_8521),
        .dout(new_Jinkela_wire_8522)
    );

    spl2 new_Jinkela_splitter_711 (
        .a(new_Jinkela_wire_8459),
        .b(new_Jinkela_wire_8460),
        .c(new_Jinkela_wire_8461)
    );

    bfr new_Jinkela_buffer_6791 (
        .din(new_Jinkela_wire_8522),
        .dout(new_Jinkela_wire_8523)
    );

    bfr new_Jinkela_buffer_6863 (
        .din(new_Jinkela_wire_8606),
        .dout(new_Jinkela_wire_8607)
    );

    bfr new_Jinkela_buffer_6944 (
        .din(new_Jinkela_wire_8697),
        .dout(new_Jinkela_wire_8698)
    );

    bfr new_Jinkela_buffer_6792 (
        .din(new_Jinkela_wire_8523),
        .dout(new_Jinkela_wire_8524)
    );

    bfr new_Jinkela_buffer_6864 (
        .din(new_Jinkela_wire_8607),
        .dout(new_Jinkela_wire_8608)
    );

    bfr new_Jinkela_buffer_6793 (
        .din(new_Jinkela_wire_8524),
        .dout(new_Jinkela_wire_8525)
    );

    bfr new_Jinkela_buffer_7074 (
        .din(_0052_),
        .dout(new_Jinkela_wire_8838)
    );

    bfr new_Jinkela_buffer_6794 (
        .din(new_Jinkela_wire_8525),
        .dout(new_Jinkela_wire_8526)
    );

    bfr new_Jinkela_buffer_6865 (
        .din(new_Jinkela_wire_8608),
        .dout(new_Jinkela_wire_8609)
    );

    bfr new_Jinkela_buffer_6795 (
        .din(new_Jinkela_wire_8526),
        .dout(new_Jinkela_wire_8527)
    );

    bfr new_Jinkela_buffer_6945 (
        .din(new_Jinkela_wire_8698),
        .dout(new_Jinkela_wire_8699)
    );

    bfr new_Jinkela_buffer_6796 (
        .din(new_Jinkela_wire_8527),
        .dout(new_Jinkela_wire_8528)
    );

    bfr new_Jinkela_buffer_6866 (
        .din(new_Jinkela_wire_8609),
        .dout(new_Jinkela_wire_8610)
    );

    bfr new_Jinkela_buffer_6797 (
        .din(new_Jinkela_wire_8528),
        .dout(new_Jinkela_wire_8529)
    );

    bfr new_Jinkela_buffer_7005 (
        .din(new_Jinkela_wire_8766),
        .dout(new_Jinkela_wire_8767)
    );

    bfr new_Jinkela_buffer_6798 (
        .din(new_Jinkela_wire_8529),
        .dout(new_Jinkela_wire_8530)
    );

    bfr new_Jinkela_buffer_6867 (
        .din(new_Jinkela_wire_8610),
        .dout(new_Jinkela_wire_8611)
    );

    bfr new_Jinkela_buffer_6799 (
        .din(new_Jinkela_wire_8530),
        .dout(new_Jinkela_wire_8531)
    );

    bfr new_Jinkela_buffer_6946 (
        .din(new_Jinkela_wire_8699),
        .dout(new_Jinkela_wire_8700)
    );

    bfr new_Jinkela_buffer_6800 (
        .din(new_Jinkela_wire_8531),
        .dout(new_Jinkela_wire_8532)
    );

    bfr new_Jinkela_buffer_13670 (
        .din(new_Jinkela_wire_16325),
        .dout(new_Jinkela_wire_16326)
    );

    bfr new_Jinkela_buffer_3398 (
        .din(new_Jinkela_wire_4527),
        .dout(new_Jinkela_wire_4528)
    );

    bfr new_Jinkela_buffer_13789 (
        .din(new_Jinkela_wire_16454),
        .dout(new_Jinkela_wire_16455)
    );

    bfr new_Jinkela_buffer_3313 (
        .din(new_Jinkela_wire_4434),
        .dout(new_Jinkela_wire_4435)
    );

    bfr new_Jinkela_buffer_13671 (
        .din(new_Jinkela_wire_16326),
        .dout(new_Jinkela_wire_16327)
    );

    bfr new_Jinkela_buffer_13750 (
        .din(new_Jinkela_wire_16411),
        .dout(new_Jinkela_wire_16412)
    );

    bfr new_Jinkela_buffer_3442 (
        .din(new_Jinkela_wire_4579),
        .dout(new_Jinkela_wire_4580)
    );

    bfr new_Jinkela_buffer_3314 (
        .din(new_Jinkela_wire_4435),
        .dout(new_Jinkela_wire_4436)
    );

    bfr new_Jinkela_buffer_13672 (
        .din(new_Jinkela_wire_16327),
        .dout(new_Jinkela_wire_16328)
    );

    bfr new_Jinkela_buffer_3399 (
        .din(new_Jinkela_wire_4528),
        .dout(new_Jinkela_wire_4529)
    );

    bfr new_Jinkela_buffer_3315 (
        .din(new_Jinkela_wire_4436),
        .dout(new_Jinkela_wire_4437)
    );

    bfr new_Jinkela_buffer_13852 (
        .din(_1229_),
        .dout(new_Jinkela_wire_16532)
    );

    bfr new_Jinkela_buffer_13673 (
        .din(new_Jinkela_wire_16328),
        .dout(new_Jinkela_wire_16329)
    );

    bfr new_Jinkela_buffer_13751 (
        .din(new_Jinkela_wire_16412),
        .dout(new_Jinkela_wire_16413)
    );

    bfr new_Jinkela_buffer_3429 (
        .din(new_Jinkela_wire_4562),
        .dout(new_Jinkela_wire_4563)
    );

    bfr new_Jinkela_buffer_3316 (
        .din(new_Jinkela_wire_4437),
        .dout(new_Jinkela_wire_4438)
    );

    spl2 new_Jinkela_splitter_1177 (
        .a(new_Jinkela_wire_16329),
        .b(new_Jinkela_wire_16330),
        .c(new_Jinkela_wire_16331)
    );

    bfr new_Jinkela_buffer_3400 (
        .din(new_Jinkela_wire_4529),
        .dout(new_Jinkela_wire_4530)
    );

    bfr new_Jinkela_buffer_13752 (
        .din(new_Jinkela_wire_16413),
        .dout(new_Jinkela_wire_16414)
    );

    bfr new_Jinkela_buffer_3317 (
        .din(new_Jinkela_wire_4438),
        .dout(new_Jinkela_wire_4439)
    );

    bfr new_Jinkela_buffer_13790 (
        .din(new_Jinkela_wire_16455),
        .dout(new_Jinkela_wire_16456)
    );

    bfr new_Jinkela_buffer_13847 (
        .din(new_Jinkela_wire_16520),
        .dout(new_Jinkela_wire_16521)
    );

    bfr new_Jinkela_buffer_3318 (
        .din(new_Jinkela_wire_4439),
        .dout(new_Jinkela_wire_4440)
    );

    bfr new_Jinkela_buffer_13753 (
        .din(new_Jinkela_wire_16414),
        .dout(new_Jinkela_wire_16415)
    );

    bfr new_Jinkela_buffer_3401 (
        .din(new_Jinkela_wire_4530),
        .dout(new_Jinkela_wire_4531)
    );

    bfr new_Jinkela_buffer_13791 (
        .din(new_Jinkela_wire_16456),
        .dout(new_Jinkela_wire_16457)
    );

    bfr new_Jinkela_buffer_3319 (
        .din(new_Jinkela_wire_4440),
        .dout(new_Jinkela_wire_4441)
    );

    bfr new_Jinkela_buffer_13754 (
        .din(new_Jinkela_wire_16415),
        .dout(new_Jinkela_wire_16416)
    );

    bfr new_Jinkela_buffer_3430 (
        .din(new_Jinkela_wire_4563),
        .dout(new_Jinkela_wire_4564)
    );

    bfr new_Jinkela_buffer_3320 (
        .din(new_Jinkela_wire_4441),
        .dout(new_Jinkela_wire_4442)
    );

    bfr new_Jinkela_buffer_13755 (
        .din(new_Jinkela_wire_16416),
        .dout(new_Jinkela_wire_16417)
    );

    bfr new_Jinkela_buffer_3402 (
        .din(new_Jinkela_wire_4531),
        .dout(new_Jinkela_wire_4532)
    );

    bfr new_Jinkela_buffer_13792 (
        .din(new_Jinkela_wire_16457),
        .dout(new_Jinkela_wire_16458)
    );

    bfr new_Jinkela_buffer_3321 (
        .din(new_Jinkela_wire_4442),
        .dout(new_Jinkela_wire_4443)
    );

    bfr new_Jinkela_buffer_13756 (
        .din(new_Jinkela_wire_16417),
        .dout(new_Jinkela_wire_16418)
    );

    bfr new_Jinkela_buffer_13849 (
        .din(new_Jinkela_wire_16526),
        .dout(new_Jinkela_wire_16527)
    );

    bfr new_Jinkela_buffer_3443 (
        .din(new_Jinkela_wire_4580),
        .dout(new_Jinkela_wire_4581)
    );

    bfr new_Jinkela_buffer_3322 (
        .din(new_Jinkela_wire_4443),
        .dout(new_Jinkela_wire_4444)
    );

    bfr new_Jinkela_buffer_13757 (
        .din(new_Jinkela_wire_16418),
        .dout(new_Jinkela_wire_16419)
    );

    bfr new_Jinkela_buffer_3403 (
        .din(new_Jinkela_wire_4532),
        .dout(new_Jinkela_wire_4533)
    );

    bfr new_Jinkela_buffer_13793 (
        .din(new_Jinkela_wire_16458),
        .dout(new_Jinkela_wire_16459)
    );

    bfr new_Jinkela_buffer_3323 (
        .din(new_Jinkela_wire_4444),
        .dout(new_Jinkela_wire_4445)
    );

    bfr new_Jinkela_buffer_13758 (
        .din(new_Jinkela_wire_16419),
        .dout(new_Jinkela_wire_16420)
    );

    bfr new_Jinkela_buffer_13853 (
        .din(_1205_),
        .dout(new_Jinkela_wire_16535)
    );

    bfr new_Jinkela_buffer_3431 (
        .din(new_Jinkela_wire_4564),
        .dout(new_Jinkela_wire_4565)
    );

    bfr new_Jinkela_buffer_3324 (
        .din(new_Jinkela_wire_4445),
        .dout(new_Jinkela_wire_4446)
    );

    spl2 new_Jinkela_splitter_1189 (
        .a(_0706_),
        .b(new_Jinkela_wire_16533),
        .c(new_Jinkela_wire_16534)
    );

    bfr new_Jinkela_buffer_13759 (
        .din(new_Jinkela_wire_16420),
        .dout(new_Jinkela_wire_16421)
    );

    bfr new_Jinkela_buffer_3404 (
        .din(new_Jinkela_wire_4533),
        .dout(new_Jinkela_wire_4534)
    );

    bfr new_Jinkela_buffer_13794 (
        .din(new_Jinkela_wire_16459),
        .dout(new_Jinkela_wire_16460)
    );

    bfr new_Jinkela_buffer_3325 (
        .din(new_Jinkela_wire_4446),
        .dout(new_Jinkela_wire_4447)
    );

    bfr new_Jinkela_buffer_13760 (
        .din(new_Jinkela_wire_16421),
        .dout(new_Jinkela_wire_16422)
    );

    bfr new_Jinkela_buffer_13850 (
        .din(new_Jinkela_wire_16527),
        .dout(new_Jinkela_wire_16528)
    );

    bfr new_Jinkela_buffer_3326 (
        .din(new_Jinkela_wire_4447),
        .dout(new_Jinkela_wire_4448)
    );

    bfr new_Jinkela_buffer_13761 (
        .din(new_Jinkela_wire_16422),
        .dout(new_Jinkela_wire_16423)
    );

    bfr new_Jinkela_buffer_3405 (
        .din(new_Jinkela_wire_4534),
        .dout(new_Jinkela_wire_4535)
    );

    bfr new_Jinkela_buffer_13795 (
        .din(new_Jinkela_wire_16460),
        .dout(new_Jinkela_wire_16461)
    );

    bfr new_Jinkela_buffer_3327 (
        .din(new_Jinkela_wire_4448),
        .dout(new_Jinkela_wire_4449)
    );

    bfr new_Jinkela_buffer_13762 (
        .din(new_Jinkela_wire_16423),
        .dout(new_Jinkela_wire_16424)
    );

    spl2 new_Jinkela_splitter_423 (
        .a(_0518_),
        .b(new_Jinkela_wire_4675),
        .c(new_Jinkela_wire_4676)
    );

    bfr new_Jinkela_buffer_13918 (
        .din(new_net_3926),
        .dout(new_Jinkela_wire_16602)
    );

    bfr new_Jinkela_buffer_3432 (
        .din(new_Jinkela_wire_4565),
        .dout(new_Jinkela_wire_4566)
    );

    bfr new_Jinkela_buffer_3328 (
        .din(new_Jinkela_wire_4449),
        .dout(new_Jinkela_wire_4450)
    );

    bfr new_Jinkela_buffer_13763 (
        .din(new_Jinkela_wire_16424),
        .dout(new_Jinkela_wire_16425)
    );

    bfr new_Jinkela_buffer_3406 (
        .din(new_Jinkela_wire_4535),
        .dout(new_Jinkela_wire_4536)
    );

    bfr new_Jinkela_buffer_13796 (
        .din(new_Jinkela_wire_16461),
        .dout(new_Jinkela_wire_16462)
    );

    bfr new_Jinkela_buffer_3329 (
        .din(new_Jinkela_wire_4450),
        .dout(new_Jinkela_wire_4451)
    );

    bfr new_Jinkela_buffer_13764 (
        .din(new_Jinkela_wire_16425),
        .dout(new_Jinkela_wire_16426)
    );

    bfr new_Jinkela_buffer_13851 (
        .din(new_Jinkela_wire_16528),
        .dout(new_Jinkela_wire_16529)
    );

    bfr new_Jinkela_buffer_3444 (
        .din(new_Jinkela_wire_4581),
        .dout(new_Jinkela_wire_4582)
    );

    bfr new_Jinkela_buffer_3330 (
        .din(new_Jinkela_wire_4451),
        .dout(new_Jinkela_wire_4452)
    );

    bfr new_Jinkela_buffer_13765 (
        .din(new_Jinkela_wire_16426),
        .dout(new_Jinkela_wire_16427)
    );

    bfr new_Jinkela_buffer_3407 (
        .din(new_Jinkela_wire_4536),
        .dout(new_Jinkela_wire_4537)
    );

    bfr new_Jinkela_buffer_13797 (
        .din(new_Jinkela_wire_16462),
        .dout(new_Jinkela_wire_16463)
    );

    bfr new_Jinkela_buffer_3331 (
        .din(new_Jinkela_wire_4452),
        .dout(new_Jinkela_wire_4453)
    );

    bfr new_Jinkela_buffer_13766 (
        .din(new_Jinkela_wire_16427),
        .dout(new_Jinkela_wire_16428)
    );

    spl2 new_Jinkela_splitter_416 (
        .a(new_Jinkela_wire_4566),
        .b(new_Jinkela_wire_4567),
        .c(new_Jinkela_wire_4568)
    );

    bfr new_Jinkela_buffer_3332 (
        .din(new_Jinkela_wire_4453),
        .dout(new_Jinkela_wire_4454)
    );

    bfr new_Jinkela_buffer_13917 (
        .din(_1360_),
        .dout(new_Jinkela_wire_16601)
    );

    bfr new_Jinkela_buffer_13767 (
        .din(new_Jinkela_wire_16428),
        .dout(new_Jinkela_wire_16429)
    );

    bfr new_Jinkela_buffer_13798 (
        .din(new_Jinkela_wire_16463),
        .dout(new_Jinkela_wire_16464)
    );

    bfr new_Jinkela_buffer_3527 (
        .din(_1624_),
        .dout(new_Jinkela_wire_4677)
    );

    bfr new_Jinkela_buffer_3333 (
        .din(new_Jinkela_wire_4454),
        .dout(new_Jinkela_wire_4455)
    );

    bfr new_Jinkela_buffer_17334 (
        .din(_1003_),
        .dout(new_Jinkela_wire_20683)
    );

    bfr new_Jinkela_buffer_17307 (
        .din(new_Jinkela_wire_20653),
        .dout(new_Jinkela_wire_20654)
    );

    bfr new_Jinkela_buffer_17101 (
        .din(new_Jinkela_wire_20435),
        .dout(new_Jinkela_wire_20436)
    );

    bfr new_Jinkela_buffer_17195 (
        .din(new_Jinkela_wire_20531),
        .dout(new_Jinkela_wire_20532)
    );

    bfr new_Jinkela_buffer_17102 (
        .din(new_Jinkela_wire_20436),
        .dout(new_Jinkela_wire_20437)
    );

    bfr new_Jinkela_buffer_17218 (
        .din(new_Jinkela_wire_20556),
        .dout(new_Jinkela_wire_20557)
    );

    bfr new_Jinkela_buffer_17103 (
        .din(new_Jinkela_wire_20437),
        .dout(new_Jinkela_wire_20438)
    );

    bfr new_Jinkela_buffer_17196 (
        .din(new_Jinkela_wire_20532),
        .dout(new_Jinkela_wire_20533)
    );

    bfr new_Jinkela_buffer_17104 (
        .din(new_Jinkela_wire_20438),
        .dout(new_Jinkela_wire_20439)
    );

    bfr new_Jinkela_buffer_17239 (
        .din(new_Jinkela_wire_20581),
        .dout(new_Jinkela_wire_20582)
    );

    bfr new_Jinkela_buffer_17105 (
        .din(new_Jinkela_wire_20439),
        .dout(new_Jinkela_wire_20440)
    );

    bfr new_Jinkela_buffer_17197 (
        .din(new_Jinkela_wire_20533),
        .dout(new_Jinkela_wire_20534)
    );

    bfr new_Jinkela_buffer_17106 (
        .din(new_Jinkela_wire_20440),
        .dout(new_Jinkela_wire_20441)
    );

    bfr new_Jinkela_buffer_17219 (
        .din(new_Jinkela_wire_20557),
        .dout(new_Jinkela_wire_20558)
    );

    bfr new_Jinkela_buffer_17107 (
        .din(new_Jinkela_wire_20441),
        .dout(new_Jinkela_wire_20442)
    );

    bfr new_Jinkela_buffer_17198 (
        .din(new_Jinkela_wire_20534),
        .dout(new_Jinkela_wire_20535)
    );

    bfr new_Jinkela_buffer_17108 (
        .din(new_Jinkela_wire_20442),
        .dout(new_Jinkela_wire_20443)
    );

    bfr new_Jinkela_buffer_17283 (
        .din(new_Jinkela_wire_20627),
        .dout(new_Jinkela_wire_20628)
    );

    bfr new_Jinkela_buffer_17109 (
        .din(new_Jinkela_wire_20443),
        .dout(new_Jinkela_wire_20444)
    );

    bfr new_Jinkela_buffer_17199 (
        .din(new_Jinkela_wire_20535),
        .dout(new_Jinkela_wire_20536)
    );

    bfr new_Jinkela_buffer_17110 (
        .din(new_Jinkela_wire_20444),
        .dout(new_Jinkela_wire_20445)
    );

    bfr new_Jinkela_buffer_17220 (
        .din(new_Jinkela_wire_20558),
        .dout(new_Jinkela_wire_20559)
    );

    bfr new_Jinkela_buffer_17111 (
        .din(new_Jinkela_wire_20445),
        .dout(new_Jinkela_wire_20446)
    );

    bfr new_Jinkela_buffer_17200 (
        .din(new_Jinkela_wire_20536),
        .dout(new_Jinkela_wire_20537)
    );

    bfr new_Jinkela_buffer_17112 (
        .din(new_Jinkela_wire_20446),
        .dout(new_Jinkela_wire_20447)
    );

    bfr new_Jinkela_buffer_17240 (
        .din(new_Jinkela_wire_20582),
        .dout(new_Jinkela_wire_20583)
    );

    bfr new_Jinkela_buffer_17113 (
        .din(new_Jinkela_wire_20447),
        .dout(new_Jinkela_wire_20448)
    );

    bfr new_Jinkela_buffer_17201 (
        .din(new_Jinkela_wire_20537),
        .dout(new_Jinkela_wire_20538)
    );

    bfr new_Jinkela_buffer_17114 (
        .din(new_Jinkela_wire_20448),
        .dout(new_Jinkela_wire_20449)
    );

    bfr new_Jinkela_buffer_17221 (
        .din(new_Jinkela_wire_20559),
        .dout(new_Jinkela_wire_20560)
    );

    bfr new_Jinkela_buffer_17115 (
        .din(new_Jinkela_wire_20449),
        .dout(new_Jinkela_wire_20450)
    );

    bfr new_Jinkela_buffer_17202 (
        .din(new_Jinkela_wire_20538),
        .dout(new_Jinkela_wire_20539)
    );

    bfr new_Jinkela_buffer_17116 (
        .din(new_Jinkela_wire_20450),
        .dout(new_Jinkela_wire_20451)
    );

    bfr new_Jinkela_buffer_17117 (
        .din(new_Jinkela_wire_20451),
        .dout(new_Jinkela_wire_20452)
    );

    bfr new_Jinkela_buffer_17203 (
        .din(new_Jinkela_wire_20539),
        .dout(new_Jinkela_wire_20540)
    );

    bfr new_Jinkela_buffer_17118 (
        .din(new_Jinkela_wire_20452),
        .dout(new_Jinkela_wire_20453)
    );

    bfr new_Jinkela_buffer_17222 (
        .din(new_Jinkela_wire_20560),
        .dout(new_Jinkela_wire_20561)
    );

    bfr new_Jinkela_buffer_17119 (
        .din(new_Jinkela_wire_20453),
        .dout(new_Jinkela_wire_20454)
    );

    bfr new_Jinkela_buffer_17204 (
        .din(new_Jinkela_wire_20540),
        .dout(new_Jinkela_wire_20541)
    );

    bfr new_Jinkela_buffer_17120 (
        .din(new_Jinkela_wire_20454),
        .dout(new_Jinkela_wire_20455)
    );

    bfr new_Jinkela_buffer_17241 (
        .din(new_Jinkela_wire_20583),
        .dout(new_Jinkela_wire_20584)
    );

    bfr new_Jinkela_buffer_17121 (
        .din(new_Jinkela_wire_20455),
        .dout(new_Jinkela_wire_20456)
    );

    bfr new_Jinkela_buffer_10382 (
        .din(new_Jinkela_wire_12549),
        .dout(new_Jinkela_wire_12550)
    );

    bfr new_Jinkela_buffer_10234 (
        .din(new_Jinkela_wire_12397),
        .dout(new_Jinkela_wire_12398)
    );

    bfr new_Jinkela_buffer_10532 (
        .din(new_Jinkela_wire_12719),
        .dout(new_Jinkela_wire_12720)
    );

    bfr new_Jinkela_buffer_10235 (
        .din(new_Jinkela_wire_12398),
        .dout(new_Jinkela_wire_12399)
    );

    bfr new_Jinkela_buffer_10383 (
        .din(new_Jinkela_wire_12550),
        .dout(new_Jinkela_wire_12551)
    );

    bfr new_Jinkela_buffer_10236 (
        .din(new_Jinkela_wire_12399),
        .dout(new_Jinkela_wire_12400)
    );

    bfr new_Jinkela_buffer_10459 (
        .din(new_Jinkela_wire_12636),
        .dout(new_Jinkela_wire_12637)
    );

    bfr new_Jinkela_buffer_10237 (
        .din(new_Jinkela_wire_12400),
        .dout(new_Jinkela_wire_12401)
    );

    bfr new_Jinkela_buffer_10384 (
        .din(new_Jinkela_wire_12551),
        .dout(new_Jinkela_wire_12552)
    );

    bfr new_Jinkela_buffer_10238 (
        .din(new_Jinkela_wire_12401),
        .dout(new_Jinkela_wire_12402)
    );

    spl2 new_Jinkela_splitter_944 (
        .a(_0549_),
        .b(new_Jinkela_wire_12729),
        .c(new_Jinkela_wire_12730)
    );

    bfr new_Jinkela_buffer_10239 (
        .din(new_Jinkela_wire_12402),
        .dout(new_Jinkela_wire_12403)
    );

    bfr new_Jinkela_buffer_10385 (
        .din(new_Jinkela_wire_12552),
        .dout(new_Jinkela_wire_12553)
    );

    bfr new_Jinkela_buffer_10240 (
        .din(new_Jinkela_wire_12403),
        .dout(new_Jinkela_wire_12404)
    );

    bfr new_Jinkela_buffer_10460 (
        .din(new_Jinkela_wire_12637),
        .dout(new_Jinkela_wire_12638)
    );

    bfr new_Jinkela_buffer_10241 (
        .din(new_Jinkela_wire_12404),
        .dout(new_Jinkela_wire_12405)
    );

    bfr new_Jinkela_buffer_10386 (
        .din(new_Jinkela_wire_12553),
        .dout(new_Jinkela_wire_12554)
    );

    bfr new_Jinkela_buffer_10242 (
        .din(new_Jinkela_wire_12405),
        .dout(new_Jinkela_wire_12406)
    );

    bfr new_Jinkela_buffer_10533 (
        .din(new_Jinkela_wire_12720),
        .dout(new_Jinkela_wire_12721)
    );

    bfr new_Jinkela_buffer_10243 (
        .din(new_Jinkela_wire_12406),
        .dout(new_Jinkela_wire_12407)
    );

    bfr new_Jinkela_buffer_10387 (
        .din(new_Jinkela_wire_12554),
        .dout(new_Jinkela_wire_12555)
    );

    bfr new_Jinkela_buffer_10244 (
        .din(new_Jinkela_wire_12407),
        .dout(new_Jinkela_wire_12408)
    );

    bfr new_Jinkela_buffer_10461 (
        .din(new_Jinkela_wire_12638),
        .dout(new_Jinkela_wire_12639)
    );

    bfr new_Jinkela_buffer_10245 (
        .din(new_Jinkela_wire_12408),
        .dout(new_Jinkela_wire_12409)
    );

    bfr new_Jinkela_buffer_10388 (
        .din(new_Jinkela_wire_12555),
        .dout(new_Jinkela_wire_12556)
    );

    bfr new_Jinkela_buffer_10246 (
        .din(new_Jinkela_wire_12409),
        .dout(new_Jinkela_wire_12410)
    );

    spl2 new_Jinkela_splitter_945 (
        .a(_0588_),
        .b(new_Jinkela_wire_12731),
        .c(new_Jinkela_wire_12732)
    );

    bfr new_Jinkela_buffer_10247 (
        .din(new_Jinkela_wire_12410),
        .dout(new_Jinkela_wire_12411)
    );

    bfr new_Jinkela_buffer_10389 (
        .din(new_Jinkela_wire_12556),
        .dout(new_Jinkela_wire_12557)
    );

    bfr new_Jinkela_buffer_10248 (
        .din(new_Jinkela_wire_12411),
        .dout(new_Jinkela_wire_12412)
    );

    bfr new_Jinkela_buffer_10462 (
        .din(new_Jinkela_wire_12639),
        .dout(new_Jinkela_wire_12640)
    );

    bfr new_Jinkela_buffer_10249 (
        .din(new_Jinkela_wire_12412),
        .dout(new_Jinkela_wire_12413)
    );

    bfr new_Jinkela_buffer_10390 (
        .din(new_Jinkela_wire_12557),
        .dout(new_Jinkela_wire_12558)
    );

    bfr new_Jinkela_buffer_10250 (
        .din(new_Jinkela_wire_12413),
        .dout(new_Jinkela_wire_12414)
    );

    bfr new_Jinkela_buffer_10534 (
        .din(new_Jinkela_wire_12721),
        .dout(new_Jinkela_wire_12722)
    );

    bfr new_Jinkela_buffer_10251 (
        .din(new_Jinkela_wire_12414),
        .dout(new_Jinkela_wire_12415)
    );

    bfr new_Jinkela_buffer_10391 (
        .din(new_Jinkela_wire_12558),
        .dout(new_Jinkela_wire_12559)
    );

    bfr new_Jinkela_buffer_10252 (
        .din(new_Jinkela_wire_12415),
        .dout(new_Jinkela_wire_12416)
    );

    bfr new_Jinkela_buffer_10463 (
        .din(new_Jinkela_wire_12640),
        .dout(new_Jinkela_wire_12641)
    );

    bfr new_Jinkela_buffer_10253 (
        .din(new_Jinkela_wire_12416),
        .dout(new_Jinkela_wire_12417)
    );

    bfr new_Jinkela_buffer_10392 (
        .din(new_Jinkela_wire_12559),
        .dout(new_Jinkela_wire_12560)
    );

    bfr new_Jinkela_buffer_10254 (
        .din(new_Jinkela_wire_12417),
        .dout(new_Jinkela_wire_12418)
    );

    bfr new_Jinkela_buffer_3334 (
        .din(new_Jinkela_wire_4455),
        .dout(new_Jinkela_wire_4456)
    );

    bfr new_Jinkela_buffer_3445 (
        .din(new_Jinkela_wire_4582),
        .dout(new_Jinkela_wire_4583)
    );

    spl2 new_Jinkela_splitter_424 (
        .a(_0586_),
        .b(new_Jinkela_wire_4678),
        .c(new_Jinkela_wire_4679)
    );

    bfr new_Jinkela_buffer_3335 (
        .din(new_Jinkela_wire_4456),
        .dout(new_Jinkela_wire_4457)
    );

    spl2 new_Jinkela_splitter_425 (
        .a(_0314_),
        .b(new_Jinkela_wire_4680),
        .c(new_Jinkela_wire_4681)
    );

    bfr new_Jinkela_buffer_3446 (
        .din(new_Jinkela_wire_4583),
        .dout(new_Jinkela_wire_4584)
    );

    bfr new_Jinkela_buffer_3336 (
        .din(new_Jinkela_wire_4457),
        .dout(new_Jinkela_wire_4458)
    );

    bfr new_Jinkela_buffer_3337 (
        .din(new_Jinkela_wire_4458),
        .dout(new_Jinkela_wire_4459)
    );

    bfr new_Jinkela_buffer_3447 (
        .din(new_Jinkela_wire_4584),
        .dout(new_Jinkela_wire_4585)
    );

    bfr new_Jinkela_buffer_3338 (
        .din(new_Jinkela_wire_4459),
        .dout(new_Jinkela_wire_4460)
    );

    bfr new_Jinkela_buffer_3339 (
        .din(new_Jinkela_wire_4460),
        .dout(new_Jinkela_wire_4461)
    );

    spl2 new_Jinkela_splitter_426 (
        .a(_1619_),
        .b(new_Jinkela_wire_4682),
        .c(new_Jinkela_wire_4683)
    );

    bfr new_Jinkela_buffer_3448 (
        .din(new_Jinkela_wire_4585),
        .dout(new_Jinkela_wire_4586)
    );

    spl2 new_Jinkela_splitter_427 (
        .a(_1532_),
        .b(new_Jinkela_wire_4688),
        .c(new_Jinkela_wire_4689)
    );

    bfr new_Jinkela_buffer_3449 (
        .din(new_Jinkela_wire_4586),
        .dout(new_Jinkela_wire_4587)
    );

    bfr new_Jinkela_buffer_3528 (
        .din(new_Jinkela_wire_4683),
        .dout(new_Jinkela_wire_4684)
    );

    spl2 new_Jinkela_splitter_428 (
        .a(_1356_),
        .b(new_Jinkela_wire_4690),
        .c(new_Jinkela_wire_4691)
    );

    bfr new_Jinkela_buffer_3450 (
        .din(new_Jinkela_wire_4587),
        .dout(new_Jinkela_wire_4588)
    );

    bfr new_Jinkela_buffer_3451 (
        .din(new_Jinkela_wire_4588),
        .dout(new_Jinkela_wire_4589)
    );

    bfr new_Jinkela_buffer_3529 (
        .din(new_Jinkela_wire_4684),
        .dout(new_Jinkela_wire_4685)
    );

    bfr new_Jinkela_buffer_3452 (
        .din(new_Jinkela_wire_4589),
        .dout(new_Jinkela_wire_4590)
    );

    spl2 new_Jinkela_splitter_429 (
        .a(_0272_),
        .b(new_Jinkela_wire_4696),
        .c(new_Jinkela_wire_4697)
    );

    bfr new_Jinkela_buffer_3453 (
        .din(new_Jinkela_wire_4590),
        .dout(new_Jinkela_wire_4591)
    );

    bfr new_Jinkela_buffer_3530 (
        .din(new_Jinkela_wire_4685),
        .dout(new_Jinkela_wire_4686)
    );

    bfr new_Jinkela_buffer_3454 (
        .din(new_Jinkela_wire_4591),
        .dout(new_Jinkela_wire_4592)
    );

    bfr new_Jinkela_buffer_3532 (
        .din(new_Jinkela_wire_4691),
        .dout(new_Jinkela_wire_4692)
    );

    spl2 new_Jinkela_splitter_430 (
        .a(_0025_),
        .b(new_Jinkela_wire_4702),
        .c(new_Jinkela_wire_4703)
    );

    bfr new_Jinkela_buffer_3455 (
        .din(new_Jinkela_wire_4592),
        .dout(new_Jinkela_wire_4593)
    );

    bfr new_Jinkela_buffer_3531 (
        .din(new_Jinkela_wire_4686),
        .dout(new_Jinkela_wire_4687)
    );

    bfr new_Jinkela_buffer_3456 (
        .din(new_Jinkela_wire_4593),
        .dout(new_Jinkela_wire_4594)
    );

    bfr new_Jinkela_buffer_3457 (
        .din(new_Jinkela_wire_4594),
        .dout(new_Jinkela_wire_4595)
    );

    bfr new_Jinkela_buffer_3533 (
        .din(new_Jinkela_wire_4692),
        .dout(new_Jinkela_wire_4693)
    );

    bfr new_Jinkela_buffer_3458 (
        .din(new_Jinkela_wire_4595),
        .dout(new_Jinkela_wire_4596)
    );

    bfr new_Jinkela_buffer_3536 (
        .din(new_Jinkela_wire_4697),
        .dout(new_Jinkela_wire_4698)
    );

    bfr new_Jinkela_buffer_3544 (
        .din(_0865_),
        .dout(new_Jinkela_wire_4708)
    );

    bfr new_Jinkela_buffer_3459 (
        .din(new_Jinkela_wire_4596),
        .dout(new_Jinkela_wire_4597)
    );

    bfr new_Jinkela_buffer_3534 (
        .din(new_Jinkela_wire_4693),
        .dout(new_Jinkela_wire_4694)
    );

    bfr new_Jinkela_buffer_3460 (
        .din(new_Jinkela_wire_4597),
        .dout(new_Jinkela_wire_4598)
    );

    bfr new_Jinkela_buffer_3540 (
        .din(new_Jinkela_wire_4703),
        .dout(new_Jinkela_wire_4704)
    );

    bfr new_Jinkela_buffer_3461 (
        .din(new_Jinkela_wire_4598),
        .dout(new_Jinkela_wire_4599)
    );

    bfr new_Jinkela_buffer_3535 (
        .din(new_Jinkela_wire_4694),
        .dout(new_Jinkela_wire_4695)
    );

    bfr new_Jinkela_buffer_3462 (
        .din(new_Jinkela_wire_4599),
        .dout(new_Jinkela_wire_4600)
    );

    bfr new_Jinkela_buffer_17205 (
        .din(new_Jinkela_wire_20541),
        .dout(new_Jinkela_wire_20542)
    );

    bfr new_Jinkela_buffer_10538 (
        .din(new_Jinkela_wire_12725),
        .dout(new_Jinkela_wire_12726)
    );

    bfr new_Jinkela_buffer_17122 (
        .din(new_Jinkela_wire_20456),
        .dout(new_Jinkela_wire_20457)
    );

    bfr new_Jinkela_buffer_10255 (
        .din(new_Jinkela_wire_12418),
        .dout(new_Jinkela_wire_12419)
    );

    bfr new_Jinkela_buffer_17223 (
        .din(new_Jinkela_wire_20561),
        .dout(new_Jinkela_wire_20562)
    );

    bfr new_Jinkela_buffer_10393 (
        .din(new_Jinkela_wire_12560),
        .dout(new_Jinkela_wire_12561)
    );

    bfr new_Jinkela_buffer_17123 (
        .din(new_Jinkela_wire_20457),
        .dout(new_Jinkela_wire_20458)
    );

    bfr new_Jinkela_buffer_10256 (
        .din(new_Jinkela_wire_12419),
        .dout(new_Jinkela_wire_12420)
    );

    bfr new_Jinkela_buffer_17206 (
        .din(new_Jinkela_wire_20542),
        .dout(new_Jinkela_wire_20543)
    );

    bfr new_Jinkela_buffer_10464 (
        .din(new_Jinkela_wire_12641),
        .dout(new_Jinkela_wire_12642)
    );

    bfr new_Jinkela_buffer_17124 (
        .din(new_Jinkela_wire_20458),
        .dout(new_Jinkela_wire_20459)
    );

    bfr new_Jinkela_buffer_10257 (
        .din(new_Jinkela_wire_12420),
        .dout(new_Jinkela_wire_12421)
    );

    bfr new_Jinkela_buffer_17284 (
        .din(new_Jinkela_wire_20628),
        .dout(new_Jinkela_wire_20629)
    );

    bfr new_Jinkela_buffer_10394 (
        .din(new_Jinkela_wire_12561),
        .dout(new_Jinkela_wire_12562)
    );

    bfr new_Jinkela_buffer_17125 (
        .din(new_Jinkela_wire_20459),
        .dout(new_Jinkela_wire_20460)
    );

    bfr new_Jinkela_buffer_10258 (
        .din(new_Jinkela_wire_12421),
        .dout(new_Jinkela_wire_12422)
    );

    bfr new_Jinkela_buffer_17207 (
        .din(new_Jinkela_wire_20543),
        .dout(new_Jinkela_wire_20544)
    );

    bfr new_Jinkela_buffer_17126 (
        .din(new_Jinkela_wire_20460),
        .dout(new_Jinkela_wire_20461)
    );

    bfr new_Jinkela_buffer_10259 (
        .din(new_Jinkela_wire_12422),
        .dout(new_Jinkela_wire_12423)
    );

    bfr new_Jinkela_buffer_17224 (
        .din(new_Jinkela_wire_20562),
        .dout(new_Jinkela_wire_20563)
    );

    bfr new_Jinkela_buffer_10395 (
        .din(new_Jinkela_wire_12562),
        .dout(new_Jinkela_wire_12563)
    );

    bfr new_Jinkela_buffer_17127 (
        .din(new_Jinkela_wire_20461),
        .dout(new_Jinkela_wire_20462)
    );

    bfr new_Jinkela_buffer_10260 (
        .din(new_Jinkela_wire_12423),
        .dout(new_Jinkela_wire_12424)
    );

    bfr new_Jinkela_buffer_17208 (
        .din(new_Jinkela_wire_20544),
        .dout(new_Jinkela_wire_20545)
    );

    bfr new_Jinkela_buffer_10465 (
        .din(new_Jinkela_wire_12642),
        .dout(new_Jinkela_wire_12643)
    );

    bfr new_Jinkela_buffer_17128 (
        .din(new_Jinkela_wire_20462),
        .dout(new_Jinkela_wire_20463)
    );

    bfr new_Jinkela_buffer_10261 (
        .din(new_Jinkela_wire_12424),
        .dout(new_Jinkela_wire_12425)
    );

    bfr new_Jinkela_buffer_17242 (
        .din(new_Jinkela_wire_20584),
        .dout(new_Jinkela_wire_20585)
    );

    bfr new_Jinkela_buffer_10396 (
        .din(new_Jinkela_wire_12563),
        .dout(new_Jinkela_wire_12564)
    );

    bfr new_Jinkela_buffer_17129 (
        .din(new_Jinkela_wire_20463),
        .dout(new_Jinkela_wire_20464)
    );

    bfr new_Jinkela_buffer_10262 (
        .din(new_Jinkela_wire_12425),
        .dout(new_Jinkela_wire_12426)
    );

    spl2 new_Jinkela_splitter_1517 (
        .a(new_Jinkela_wire_20545),
        .b(new_Jinkela_wire_20546),
        .c(new_Jinkela_wire_20547)
    );

    spl2 new_Jinkela_splitter_943 (
        .a(new_Jinkela_wire_12726),
        .b(new_Jinkela_wire_12727),
        .c(new_Jinkela_wire_12728)
    );

    bfr new_Jinkela_buffer_17130 (
        .din(new_Jinkela_wire_20464),
        .dout(new_Jinkela_wire_20465)
    );

    bfr new_Jinkela_buffer_10263 (
        .din(new_Jinkela_wire_12426),
        .dout(new_Jinkela_wire_12427)
    );

    bfr new_Jinkela_buffer_10397 (
        .din(new_Jinkela_wire_12564),
        .dout(new_Jinkela_wire_12565)
    );

    bfr new_Jinkela_buffer_17308 (
        .din(new_Jinkela_wire_20654),
        .dout(new_Jinkela_wire_20655)
    );

    bfr new_Jinkela_buffer_17131 (
        .din(new_Jinkela_wire_20465),
        .dout(new_Jinkela_wire_20466)
    );

    bfr new_Jinkela_buffer_10264 (
        .din(new_Jinkela_wire_12427),
        .dout(new_Jinkela_wire_12428)
    );

    bfr new_Jinkela_buffer_17225 (
        .din(new_Jinkela_wire_20563),
        .dout(new_Jinkela_wire_20564)
    );

    bfr new_Jinkela_buffer_10466 (
        .din(new_Jinkela_wire_12643),
        .dout(new_Jinkela_wire_12644)
    );

    bfr new_Jinkela_buffer_17132 (
        .din(new_Jinkela_wire_20466),
        .dout(new_Jinkela_wire_20467)
    );

    bfr new_Jinkela_buffer_10265 (
        .din(new_Jinkela_wire_12428),
        .dout(new_Jinkela_wire_12429)
    );

    bfr new_Jinkela_buffer_17226 (
        .din(new_Jinkela_wire_20564),
        .dout(new_Jinkela_wire_20565)
    );

    bfr new_Jinkela_buffer_10398 (
        .din(new_Jinkela_wire_12565),
        .dout(new_Jinkela_wire_12566)
    );

    bfr new_Jinkela_buffer_17133 (
        .din(new_Jinkela_wire_20467),
        .dout(new_Jinkela_wire_20468)
    );

    bfr new_Jinkela_buffer_10266 (
        .din(new_Jinkela_wire_12429),
        .dout(new_Jinkela_wire_12430)
    );

    bfr new_Jinkela_buffer_17243 (
        .din(new_Jinkela_wire_20585),
        .dout(new_Jinkela_wire_20586)
    );

    spl2 new_Jinkela_splitter_947 (
        .a(_1440_),
        .b(new_Jinkela_wire_12735),
        .c(new_Jinkela_wire_12736)
    );

    bfr new_Jinkela_buffer_17134 (
        .din(new_Jinkela_wire_20468),
        .dout(new_Jinkela_wire_20469)
    );

    bfr new_Jinkela_buffer_10267 (
        .din(new_Jinkela_wire_12430),
        .dout(new_Jinkela_wire_12431)
    );

    bfr new_Jinkela_buffer_17227 (
        .din(new_Jinkela_wire_20565),
        .dout(new_Jinkela_wire_20566)
    );

    bfr new_Jinkela_buffer_10399 (
        .din(new_Jinkela_wire_12566),
        .dout(new_Jinkela_wire_12567)
    );

    bfr new_Jinkela_buffer_17135 (
        .din(new_Jinkela_wire_20469),
        .dout(new_Jinkela_wire_20470)
    );

    bfr new_Jinkela_buffer_10268 (
        .din(new_Jinkela_wire_12431),
        .dout(new_Jinkela_wire_12432)
    );

    bfr new_Jinkela_buffer_17285 (
        .din(new_Jinkela_wire_20629),
        .dout(new_Jinkela_wire_20630)
    );

    bfr new_Jinkela_buffer_10467 (
        .din(new_Jinkela_wire_12644),
        .dout(new_Jinkela_wire_12645)
    );

    bfr new_Jinkela_buffer_17136 (
        .din(new_Jinkela_wire_20470),
        .dout(new_Jinkela_wire_20471)
    );

    bfr new_Jinkela_buffer_10269 (
        .din(new_Jinkela_wire_12432),
        .dout(new_Jinkela_wire_12433)
    );

    bfr new_Jinkela_buffer_17228 (
        .din(new_Jinkela_wire_20566),
        .dout(new_Jinkela_wire_20567)
    );

    bfr new_Jinkela_buffer_10400 (
        .din(new_Jinkela_wire_12567),
        .dout(new_Jinkela_wire_12568)
    );

    bfr new_Jinkela_buffer_17137 (
        .din(new_Jinkela_wire_20471),
        .dout(new_Jinkela_wire_20472)
    );

    bfr new_Jinkela_buffer_10270 (
        .din(new_Jinkela_wire_12433),
        .dout(new_Jinkela_wire_12434)
    );

    bfr new_Jinkela_buffer_17244 (
        .din(new_Jinkela_wire_20586),
        .dout(new_Jinkela_wire_20587)
    );

    spl2 new_Jinkela_splitter_946 (
        .a(_0965_),
        .b(new_Jinkela_wire_12733),
        .c(new_Jinkela_wire_12734)
    );

    bfr new_Jinkela_buffer_17138 (
        .din(new_Jinkela_wire_20472),
        .dout(new_Jinkela_wire_20473)
    );

    bfr new_Jinkela_buffer_10271 (
        .din(new_Jinkela_wire_12434),
        .dout(new_Jinkela_wire_12435)
    );

    bfr new_Jinkela_buffer_17229 (
        .din(new_Jinkela_wire_20567),
        .dout(new_Jinkela_wire_20568)
    );

    bfr new_Jinkela_buffer_10401 (
        .din(new_Jinkela_wire_12568),
        .dout(new_Jinkela_wire_12569)
    );

    bfr new_Jinkela_buffer_17139 (
        .din(new_Jinkela_wire_20473),
        .dout(new_Jinkela_wire_20474)
    );

    bfr new_Jinkela_buffer_10272 (
        .din(new_Jinkela_wire_12435),
        .dout(new_Jinkela_wire_12436)
    );

    bfr new_Jinkela_buffer_10468 (
        .din(new_Jinkela_wire_12645),
        .dout(new_Jinkela_wire_12646)
    );

    bfr new_Jinkela_buffer_17330 (
        .din(new_Jinkela_wire_20678),
        .dout(new_Jinkela_wire_20679)
    );

    bfr new_Jinkela_buffer_17140 (
        .din(new_Jinkela_wire_20474),
        .dout(new_Jinkela_wire_20475)
    );

    bfr new_Jinkela_buffer_10273 (
        .din(new_Jinkela_wire_12436),
        .dout(new_Jinkela_wire_12437)
    );

    bfr new_Jinkela_buffer_17230 (
        .din(new_Jinkela_wire_20568),
        .dout(new_Jinkela_wire_20569)
    );

    bfr new_Jinkela_buffer_10402 (
        .din(new_Jinkela_wire_12569),
        .dout(new_Jinkela_wire_12570)
    );

    bfr new_Jinkela_buffer_17141 (
        .din(new_Jinkela_wire_20475),
        .dout(new_Jinkela_wire_20476)
    );

    bfr new_Jinkela_buffer_10274 (
        .din(new_Jinkela_wire_12437),
        .dout(new_Jinkela_wire_12438)
    );

    bfr new_Jinkela_buffer_17245 (
        .din(new_Jinkela_wire_20587),
        .dout(new_Jinkela_wire_20588)
    );

    bfr new_Jinkela_buffer_10540 (
        .din(_0683_),
        .dout(new_Jinkela_wire_12738)
    );

    bfr new_Jinkela_buffer_10539 (
        .din(_1161_),
        .dout(new_Jinkela_wire_12737)
    );

    bfr new_Jinkela_buffer_17142 (
        .din(new_Jinkela_wire_20476),
        .dout(new_Jinkela_wire_20477)
    );

    bfr new_Jinkela_buffer_10275 (
        .din(new_Jinkela_wire_12438),
        .dout(new_Jinkela_wire_12439)
    );

    spl4L new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_24),
        .c(new_Jinkela_wire_25),
        .d(new_Jinkela_wire_29),
        .b(new_Jinkela_wire_34),
        .e(new_Jinkela_wire_39)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(N426),
        .b(new_Jinkela_wire_0),
        .c(new_Jinkela_wire_2)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(N154),
        .b(new_Jinkela_wire_22),
        .c(new_Jinkela_wire_24)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_6868 (
        .din(new_Jinkela_wire_8611),
        .dout(new_Jinkela_wire_8612)
    );

    bfr new_Jinkela_buffer_10403 (
        .din(new_Jinkela_wire_12570),
        .dout(new_Jinkela_wire_12571)
    );

    bfr new_Jinkela_buffer_17231 (
        .din(new_Jinkela_wire_20569),
        .dout(new_Jinkela_wire_20570)
    );

    bfr new_Jinkela_buffer_6801 (
        .din(new_Jinkela_wire_8532),
        .dout(new_Jinkela_wire_8533)
    );

    bfr new_Jinkela_buffer_10276 (
        .din(new_Jinkela_wire_12439),
        .dout(new_Jinkela_wire_12440)
    );

    bfr new_Jinkela_buffer_17143 (
        .din(new_Jinkela_wire_20477),
        .dout(new_Jinkela_wire_20478)
    );

    spl2 new_Jinkela_splitter_732 (
        .a(_1812_),
        .b(new_Jinkela_wire_8841),
        .c(new_Jinkela_wire_8842)
    );

    bfr new_Jinkela_buffer_10469 (
        .din(new_Jinkela_wire_12646),
        .dout(new_Jinkela_wire_12647)
    );

    bfr new_Jinkela_buffer_17286 (
        .din(new_Jinkela_wire_20630),
        .dout(new_Jinkela_wire_20631)
    );

    spl2 new_Jinkela_splitter_734 (
        .a(_1102_),
        .b(new_Jinkela_wire_8849),
        .c(new_Jinkela_wire_8850)
    );

    bfr new_Jinkela_buffer_6802 (
        .din(new_Jinkela_wire_8533),
        .dout(new_Jinkela_wire_8534)
    );

    bfr new_Jinkela_buffer_10277 (
        .din(new_Jinkela_wire_12440),
        .dout(new_Jinkela_wire_12441)
    );

    bfr new_Jinkela_buffer_17144 (
        .din(new_Jinkela_wire_20478),
        .dout(new_Jinkela_wire_20479)
    );

    bfr new_Jinkela_buffer_6869 (
        .din(new_Jinkela_wire_8612),
        .dout(new_Jinkela_wire_8613)
    );

    bfr new_Jinkela_buffer_10404 (
        .din(new_Jinkela_wire_12571),
        .dout(new_Jinkela_wire_12572)
    );

    bfr new_Jinkela_buffer_17232 (
        .din(new_Jinkela_wire_20570),
        .dout(new_Jinkela_wire_20571)
    );

    bfr new_Jinkela_buffer_6803 (
        .din(new_Jinkela_wire_8534),
        .dout(new_Jinkela_wire_8535)
    );

    bfr new_Jinkela_buffer_10278 (
        .din(new_Jinkela_wire_12441),
        .dout(new_Jinkela_wire_12442)
    );

    bfr new_Jinkela_buffer_17145 (
        .din(new_Jinkela_wire_20479),
        .dout(new_Jinkela_wire_20480)
    );

    bfr new_Jinkela_buffer_6947 (
        .din(new_Jinkela_wire_8700),
        .dout(new_Jinkela_wire_8701)
    );

    bfr new_Jinkela_buffer_17246 (
        .din(new_Jinkela_wire_20588),
        .dout(new_Jinkela_wire_20589)
    );

    spl2 new_Jinkela_splitter_948 (
        .a(_1755_),
        .b(new_Jinkela_wire_12739),
        .c(new_Jinkela_wire_12740)
    );

    bfr new_Jinkela_buffer_6804 (
        .din(new_Jinkela_wire_8535),
        .dout(new_Jinkela_wire_8536)
    );

    bfr new_Jinkela_buffer_10279 (
        .din(new_Jinkela_wire_12442),
        .dout(new_Jinkela_wire_12443)
    );

    bfr new_Jinkela_buffer_17146 (
        .din(new_Jinkela_wire_20480),
        .dout(new_Jinkela_wire_20481)
    );

    bfr new_Jinkela_buffer_6870 (
        .din(new_Jinkela_wire_8613),
        .dout(new_Jinkela_wire_8614)
    );

    bfr new_Jinkela_buffer_10405 (
        .din(new_Jinkela_wire_12572),
        .dout(new_Jinkela_wire_12573)
    );

    bfr new_Jinkela_buffer_17233 (
        .din(new_Jinkela_wire_20571),
        .dout(new_Jinkela_wire_20572)
    );

    bfr new_Jinkela_buffer_6805 (
        .din(new_Jinkela_wire_8536),
        .dout(new_Jinkela_wire_8537)
    );

    bfr new_Jinkela_buffer_10280 (
        .din(new_Jinkela_wire_12443),
        .dout(new_Jinkela_wire_12444)
    );

    bfr new_Jinkela_buffer_17147 (
        .din(new_Jinkela_wire_20481),
        .dout(new_Jinkela_wire_20482)
    );

    bfr new_Jinkela_buffer_7006 (
        .din(new_Jinkela_wire_8767),
        .dout(new_Jinkela_wire_8768)
    );

    bfr new_Jinkela_buffer_10470 (
        .din(new_Jinkela_wire_12647),
        .dout(new_Jinkela_wire_12648)
    );

    bfr new_Jinkela_buffer_17309 (
        .din(new_Jinkela_wire_20655),
        .dout(new_Jinkela_wire_20656)
    );

    bfr new_Jinkela_buffer_6806 (
        .din(new_Jinkela_wire_8537),
        .dout(new_Jinkela_wire_8538)
    );

    bfr new_Jinkela_buffer_10281 (
        .din(new_Jinkela_wire_12444),
        .dout(new_Jinkela_wire_12445)
    );

    bfr new_Jinkela_buffer_17148 (
        .din(new_Jinkela_wire_20482),
        .dout(new_Jinkela_wire_20483)
    );

    bfr new_Jinkela_buffer_6871 (
        .din(new_Jinkela_wire_8614),
        .dout(new_Jinkela_wire_8615)
    );

    bfr new_Jinkela_buffer_10406 (
        .din(new_Jinkela_wire_12573),
        .dout(new_Jinkela_wire_12574)
    );

    bfr new_Jinkela_buffer_17234 (
        .din(new_Jinkela_wire_20572),
        .dout(new_Jinkela_wire_20573)
    );

    bfr new_Jinkela_buffer_6807 (
        .din(new_Jinkela_wire_8538),
        .dout(new_Jinkela_wire_8539)
    );

    bfr new_Jinkela_buffer_10282 (
        .din(new_Jinkela_wire_12445),
        .dout(new_Jinkela_wire_12446)
    );

    bfr new_Jinkela_buffer_17149 (
        .din(new_Jinkela_wire_20483),
        .dout(new_Jinkela_wire_20484)
    );

    bfr new_Jinkela_buffer_6948 (
        .din(new_Jinkela_wire_8701),
        .dout(new_Jinkela_wire_8702)
    );

    bfr new_Jinkela_buffer_10541 (
        .din(_0703_),
        .dout(new_Jinkela_wire_12741)
    );

    bfr new_Jinkela_buffer_17247 (
        .din(new_Jinkela_wire_20589),
        .dout(new_Jinkela_wire_20590)
    );

    bfr new_Jinkela_buffer_6808 (
        .din(new_Jinkela_wire_8539),
        .dout(new_Jinkela_wire_8540)
    );

    bfr new_Jinkela_buffer_10283 (
        .din(new_Jinkela_wire_12446),
        .dout(new_Jinkela_wire_12447)
    );

    bfr new_Jinkela_buffer_17150 (
        .din(new_Jinkela_wire_20484),
        .dout(new_Jinkela_wire_20485)
    );

    bfr new_Jinkela_buffer_6872 (
        .din(new_Jinkela_wire_8615),
        .dout(new_Jinkela_wire_8616)
    );

    bfr new_Jinkela_buffer_10407 (
        .din(new_Jinkela_wire_12574),
        .dout(new_Jinkela_wire_12575)
    );

    spl2 new_Jinkela_splitter_1518 (
        .a(new_Jinkela_wire_20573),
        .b(new_Jinkela_wire_20574),
        .c(new_Jinkela_wire_20575)
    );

    bfr new_Jinkela_buffer_6809 (
        .din(new_Jinkela_wire_8540),
        .dout(new_Jinkela_wire_8541)
    );

    bfr new_Jinkela_buffer_10284 (
        .din(new_Jinkela_wire_12447),
        .dout(new_Jinkela_wire_12448)
    );

    bfr new_Jinkela_buffer_17151 (
        .din(new_Jinkela_wire_20485),
        .dout(new_Jinkela_wire_20486)
    );

    bfr new_Jinkela_buffer_10471 (
        .din(new_Jinkela_wire_12648),
        .dout(new_Jinkela_wire_12649)
    );

    bfr new_Jinkela_buffer_17248 (
        .din(new_Jinkela_wire_20590),
        .dout(new_Jinkela_wire_20591)
    );

    bfr new_Jinkela_buffer_6810 (
        .din(new_Jinkela_wire_8541),
        .dout(new_Jinkela_wire_8542)
    );

    bfr new_Jinkela_buffer_10285 (
        .din(new_Jinkela_wire_12448),
        .dout(new_Jinkela_wire_12449)
    );

    bfr new_Jinkela_buffer_17152 (
        .din(new_Jinkela_wire_20486),
        .dout(new_Jinkela_wire_20487)
    );

    bfr new_Jinkela_buffer_6873 (
        .din(new_Jinkela_wire_8616),
        .dout(new_Jinkela_wire_8617)
    );

    bfr new_Jinkela_buffer_10408 (
        .din(new_Jinkela_wire_12575),
        .dout(new_Jinkela_wire_12576)
    );

    bfr new_Jinkela_buffer_17287 (
        .din(new_Jinkela_wire_20631),
        .dout(new_Jinkela_wire_20632)
    );

    bfr new_Jinkela_buffer_6811 (
        .din(new_Jinkela_wire_8542),
        .dout(new_Jinkela_wire_8543)
    );

    bfr new_Jinkela_buffer_10286 (
        .din(new_Jinkela_wire_12449),
        .dout(new_Jinkela_wire_12450)
    );

    bfr new_Jinkela_buffer_17153 (
        .din(new_Jinkela_wire_20487),
        .dout(new_Jinkela_wire_20488)
    );

    bfr new_Jinkela_buffer_6949 (
        .din(new_Jinkela_wire_8702),
        .dout(new_Jinkela_wire_8703)
    );

    spl2 new_Jinkela_splitter_951 (
        .a(_0166_),
        .b(new_Jinkela_wire_12905),
        .c(new_Jinkela_wire_12906)
    );

    bfr new_Jinkela_buffer_17444 (
        .din(_1381_),
        .dout(new_Jinkela_wire_20795)
    );

    bfr new_Jinkela_buffer_6812 (
        .din(new_Jinkela_wire_8543),
        .dout(new_Jinkela_wire_8544)
    );

    bfr new_Jinkela_buffer_10287 (
        .din(new_Jinkela_wire_12450),
        .dout(new_Jinkela_wire_12451)
    );

    bfr new_Jinkela_buffer_17154 (
        .din(new_Jinkela_wire_20488),
        .dout(new_Jinkela_wire_20489)
    );

    bfr new_Jinkela_buffer_6874 (
        .din(new_Jinkela_wire_8617),
        .dout(new_Jinkela_wire_8618)
    );

    bfr new_Jinkela_buffer_10409 (
        .din(new_Jinkela_wire_12576),
        .dout(new_Jinkela_wire_12577)
    );

    bfr new_Jinkela_buffer_17249 (
        .din(new_Jinkela_wire_20591),
        .dout(new_Jinkela_wire_20592)
    );

    bfr new_Jinkela_buffer_6813 (
        .din(new_Jinkela_wire_8544),
        .dout(new_Jinkela_wire_8545)
    );

    bfr new_Jinkela_buffer_10288 (
        .din(new_Jinkela_wire_12451),
        .dout(new_Jinkela_wire_12452)
    );

    bfr new_Jinkela_buffer_17155 (
        .din(new_Jinkela_wire_20489),
        .dout(new_Jinkela_wire_20490)
    );

    bfr new_Jinkela_buffer_7007 (
        .din(new_Jinkela_wire_8768),
        .dout(new_Jinkela_wire_8769)
    );

    bfr new_Jinkela_buffer_10472 (
        .din(new_Jinkela_wire_12649),
        .dout(new_Jinkela_wire_12650)
    );

    bfr new_Jinkela_buffer_17288 (
        .din(new_Jinkela_wire_20632),
        .dout(new_Jinkela_wire_20633)
    );

    bfr new_Jinkela_buffer_6814 (
        .din(new_Jinkela_wire_8545),
        .dout(new_Jinkela_wire_8546)
    );

    bfr new_Jinkela_buffer_10289 (
        .din(new_Jinkela_wire_12452),
        .dout(new_Jinkela_wire_12453)
    );

    bfr new_Jinkela_buffer_17156 (
        .din(new_Jinkela_wire_20490),
        .dout(new_Jinkela_wire_20491)
    );

    bfr new_Jinkela_buffer_6875 (
        .din(new_Jinkela_wire_8618),
        .dout(new_Jinkela_wire_8619)
    );

    bfr new_Jinkela_buffer_10410 (
        .din(new_Jinkela_wire_12577),
        .dout(new_Jinkela_wire_12578)
    );

    bfr new_Jinkela_buffer_17250 (
        .din(new_Jinkela_wire_20592),
        .dout(new_Jinkela_wire_20593)
    );

    bfr new_Jinkela_buffer_6815 (
        .din(new_Jinkela_wire_8546),
        .dout(new_Jinkela_wire_8547)
    );

    bfr new_Jinkela_buffer_10290 (
        .din(new_Jinkela_wire_12453),
        .dout(new_Jinkela_wire_12454)
    );

    bfr new_Jinkela_buffer_17157 (
        .din(new_Jinkela_wire_20491),
        .dout(new_Jinkela_wire_20492)
    );

    bfr new_Jinkela_buffer_6950 (
        .din(new_Jinkela_wire_8703),
        .dout(new_Jinkela_wire_8704)
    );

    bfr new_Jinkela_buffer_10629 (
        .din(_1459_),
        .dout(new_Jinkela_wire_12831)
    );

    bfr new_Jinkela_buffer_17310 (
        .din(new_Jinkela_wire_20656),
        .dout(new_Jinkela_wire_20657)
    );

    bfr new_Jinkela_buffer_6816 (
        .din(new_Jinkela_wire_8547),
        .dout(new_Jinkela_wire_8548)
    );

    bfr new_Jinkela_buffer_10291 (
        .din(new_Jinkela_wire_12454),
        .dout(new_Jinkela_wire_12455)
    );

    bfr new_Jinkela_buffer_17158 (
        .din(new_Jinkela_wire_20492),
        .dout(new_Jinkela_wire_20493)
    );

    bfr new_Jinkela_buffer_6876 (
        .din(new_Jinkela_wire_8619),
        .dout(new_Jinkela_wire_8620)
    );

    bfr new_Jinkela_buffer_10411 (
        .din(new_Jinkela_wire_12578),
        .dout(new_Jinkela_wire_12579)
    );

    bfr new_Jinkela_buffer_17251 (
        .din(new_Jinkela_wire_20593),
        .dout(new_Jinkela_wire_20594)
    );

    bfr new_Jinkela_buffer_6817 (
        .din(new_Jinkela_wire_8548),
        .dout(new_Jinkela_wire_8549)
    );

    bfr new_Jinkela_buffer_10292 (
        .din(new_Jinkela_wire_12455),
        .dout(new_Jinkela_wire_12456)
    );

    bfr new_Jinkela_buffer_17159 (
        .din(new_Jinkela_wire_20493),
        .dout(new_Jinkela_wire_20494)
    );

    bfr new_Jinkela_buffer_10473 (
        .din(new_Jinkela_wire_12650),
        .dout(new_Jinkela_wire_12651)
    );

    bfr new_Jinkela_buffer_17289 (
        .din(new_Jinkela_wire_20633),
        .dout(new_Jinkela_wire_20634)
    );

    spl2 new_Jinkela_splitter_733 (
        .a(_1172_),
        .b(new_Jinkela_wire_8843),
        .c(new_Jinkela_wire_8844)
    );

    bfr new_Jinkela_buffer_6818 (
        .din(new_Jinkela_wire_8549),
        .dout(new_Jinkela_wire_8550)
    );

    bfr new_Jinkela_buffer_10293 (
        .din(new_Jinkela_wire_12456),
        .dout(new_Jinkela_wire_12457)
    );

    bfr new_Jinkela_buffer_17160 (
        .din(new_Jinkela_wire_20494),
        .dout(new_Jinkela_wire_20495)
    );

    bfr new_Jinkela_buffer_6877 (
        .din(new_Jinkela_wire_8620),
        .dout(new_Jinkela_wire_8621)
    );

    bfr new_Jinkela_buffer_10412 (
        .din(new_Jinkela_wire_12579),
        .dout(new_Jinkela_wire_12580)
    );

    bfr new_Jinkela_buffer_17252 (
        .din(new_Jinkela_wire_20594),
        .dout(new_Jinkela_wire_20595)
    );

    bfr new_Jinkela_buffer_6819 (
        .din(new_Jinkela_wire_8550),
        .dout(new_Jinkela_wire_8551)
    );

    bfr new_Jinkela_buffer_10294 (
        .din(new_Jinkela_wire_12457),
        .dout(new_Jinkela_wire_12458)
    );

    bfr new_Jinkela_buffer_17161 (
        .din(new_Jinkela_wire_20495),
        .dout(new_Jinkela_wire_20496)
    );

    bfr new_Jinkela_buffer_6951 (
        .din(new_Jinkela_wire_8704),
        .dout(new_Jinkela_wire_8705)
    );

    bfr new_Jinkela_buffer_10542 (
        .din(new_Jinkela_wire_12741),
        .dout(new_Jinkela_wire_12742)
    );

    spl2 new_Jinkela_splitter_1525 (
        .a(_0200_),
        .b(new_Jinkela_wire_20805),
        .c(new_Jinkela_wire_20806)
    );

    bfr new_Jinkela_buffer_6820 (
        .din(new_Jinkela_wire_8551),
        .dout(new_Jinkela_wire_8552)
    );

    bfr new_Jinkela_buffer_10295 (
        .din(new_Jinkela_wire_12458),
        .dout(new_Jinkela_wire_12459)
    );

    bfr new_Jinkela_buffer_17162 (
        .din(new_Jinkela_wire_20496),
        .dout(new_Jinkela_wire_20497)
    );

    bfr new_Jinkela_buffer_6878 (
        .din(new_Jinkela_wire_8621),
        .dout(new_Jinkela_wire_8622)
    );

    bfr new_Jinkela_buffer_10413 (
        .din(new_Jinkela_wire_12580),
        .dout(new_Jinkela_wire_12581)
    );

    bfr new_Jinkela_buffer_17253 (
        .din(new_Jinkela_wire_20595),
        .dout(new_Jinkela_wire_20596)
    );

    bfr new_Jinkela_buffer_6821 (
        .din(new_Jinkela_wire_8552),
        .dout(new_Jinkela_wire_8553)
    );

    bfr new_Jinkela_buffer_10296 (
        .din(new_Jinkela_wire_12459),
        .dout(new_Jinkela_wire_12460)
    );

    bfr new_Jinkela_buffer_17163 (
        .din(new_Jinkela_wire_20497),
        .dout(new_Jinkela_wire_20498)
    );

    bfr new_Jinkela_buffer_13768 (
        .din(new_Jinkela_wire_16429),
        .dout(new_Jinkela_wire_16430)
    );

    bfr new_Jinkela_buffer_13854 (
        .din(new_Jinkela_wire_16535),
        .dout(new_Jinkela_wire_16536)
    );

    bfr new_Jinkela_buffer_13769 (
        .din(new_Jinkela_wire_16430),
        .dout(new_Jinkela_wire_16431)
    );

    bfr new_Jinkela_buffer_13799 (
        .din(new_Jinkela_wire_16464),
        .dout(new_Jinkela_wire_16465)
    );

    bfr new_Jinkela_buffer_13770 (
        .din(new_Jinkela_wire_16431),
        .dout(new_Jinkela_wire_16432)
    );

    spl2 new_Jinkela_splitter_1191 (
        .a(_0253_),
        .b(new_Jinkela_wire_16694),
        .c(new_Jinkela_wire_16695)
    );

    bfr new_Jinkela_buffer_13771 (
        .din(new_Jinkela_wire_16432),
        .dout(new_Jinkela_wire_16433)
    );

    bfr new_Jinkela_buffer_13800 (
        .din(new_Jinkela_wire_16465),
        .dout(new_Jinkela_wire_16466)
    );

    spl2 new_Jinkela_splitter_1180 (
        .a(new_Jinkela_wire_16433),
        .b(new_Jinkela_wire_16434),
        .c(new_Jinkela_wire_16435)
    );

    bfr new_Jinkela_buffer_13801 (
        .din(new_Jinkela_wire_16466),
        .dout(new_Jinkela_wire_16467)
    );

    bfr new_Jinkela_buffer_13855 (
        .din(new_Jinkela_wire_16536),
        .dout(new_Jinkela_wire_16537)
    );

    spl2 new_Jinkela_splitter_1192 (
        .a(_1750_),
        .b(new_Jinkela_wire_16700),
        .c(new_Jinkela_wire_16701)
    );

    bfr new_Jinkela_buffer_13919 (
        .din(new_Jinkela_wire_16602),
        .dout(new_Jinkela_wire_16603)
    );

    bfr new_Jinkela_buffer_13802 (
        .din(new_Jinkela_wire_16467),
        .dout(new_Jinkela_wire_16468)
    );

    bfr new_Jinkela_buffer_13856 (
        .din(new_Jinkela_wire_16537),
        .dout(new_Jinkela_wire_16538)
    );

    bfr new_Jinkela_buffer_13803 (
        .din(new_Jinkela_wire_16468),
        .dout(new_Jinkela_wire_16469)
    );

    bfr new_Jinkela_buffer_14010 (
        .din(new_Jinkela_wire_16695),
        .dout(new_Jinkela_wire_16696)
    );

    bfr new_Jinkela_buffer_13804 (
        .din(new_Jinkela_wire_16469),
        .dout(new_Jinkela_wire_16470)
    );

    bfr new_Jinkela_buffer_13857 (
        .din(new_Jinkela_wire_16538),
        .dout(new_Jinkela_wire_16539)
    );

    bfr new_Jinkela_buffer_13805 (
        .din(new_Jinkela_wire_16470),
        .dout(new_Jinkela_wire_16471)
    );

    bfr new_Jinkela_buffer_13920 (
        .din(new_Jinkela_wire_16603),
        .dout(new_Jinkela_wire_16604)
    );

    bfr new_Jinkela_buffer_13806 (
        .din(new_Jinkela_wire_16471),
        .dout(new_Jinkela_wire_16472)
    );

    bfr new_Jinkela_buffer_13858 (
        .din(new_Jinkela_wire_16539),
        .dout(new_Jinkela_wire_16540)
    );

    bfr new_Jinkela_buffer_13807 (
        .din(new_Jinkela_wire_16472),
        .dout(new_Jinkela_wire_16473)
    );

    bfr new_Jinkela_buffer_13808 (
        .din(new_Jinkela_wire_16473),
        .dout(new_Jinkela_wire_16474)
    );

    bfr new_Jinkela_buffer_13859 (
        .din(new_Jinkela_wire_16540),
        .dout(new_Jinkela_wire_16541)
    );

    bfr new_Jinkela_buffer_13809 (
        .din(new_Jinkela_wire_16474),
        .dout(new_Jinkela_wire_16475)
    );

    bfr new_Jinkela_buffer_13921 (
        .din(new_Jinkela_wire_16604),
        .dout(new_Jinkela_wire_16605)
    );

    bfr new_Jinkela_buffer_13810 (
        .din(new_Jinkela_wire_16475),
        .dout(new_Jinkela_wire_16476)
    );

    bfr new_Jinkela_buffer_13860 (
        .din(new_Jinkela_wire_16541),
        .dout(new_Jinkela_wire_16542)
    );

    bfr new_Jinkela_buffer_13811 (
        .din(new_Jinkela_wire_16476),
        .dout(new_Jinkela_wire_16477)
    );

    bfr new_Jinkela_buffer_14014 (
        .din(_0095_),
        .dout(new_Jinkela_wire_16702)
    );

    bfr new_Jinkela_buffer_13812 (
        .din(new_Jinkela_wire_16477),
        .dout(new_Jinkela_wire_16478)
    );

    bfr new_Jinkela_buffer_13861 (
        .din(new_Jinkela_wire_16542),
        .dout(new_Jinkela_wire_16543)
    );

    bfr new_Jinkela_buffer_13813 (
        .din(new_Jinkela_wire_16478),
        .dout(new_Jinkela_wire_16479)
    );

    bfr new_Jinkela_buffer_14086 (
        .din(_1736_),
        .dout(new_Jinkela_wire_16776)
    );

    bfr new_Jinkela_buffer_13922 (
        .din(new_Jinkela_wire_16605),
        .dout(new_Jinkela_wire_16606)
    );

    bfr new_Jinkela_buffer_13814 (
        .din(new_Jinkela_wire_16479),
        .dout(new_Jinkela_wire_16480)
    );

    bfr new_Jinkela_buffer_13862 (
        .din(new_Jinkela_wire_16543),
        .dout(new_Jinkela_wire_16544)
    );

    bfr new_Jinkela_buffer_13815 (
        .din(new_Jinkela_wire_16480),
        .dout(new_Jinkela_wire_16481)
    );

    bfr new_Jinkela_buffer_13816 (
        .din(new_Jinkela_wire_16481),
        .dout(new_Jinkela_wire_16482)
    );

    bfr new_Jinkela_buffer_13863 (
        .din(new_Jinkela_wire_16544),
        .dout(new_Jinkela_wire_16545)
    );

    spl4L new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_2),
        .c(new_Jinkela_wire_3),
        .d(new_Jinkela_wire_7),
        .b(new_Jinkela_wire_12),
        .e(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_7008 (
        .din(new_Jinkela_wire_8769),
        .dout(new_Jinkela_wire_8770)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_0),
        .dout(new_Jinkela_wire_1)
    );

    bfr new_Jinkela_buffer_6822 (
        .din(new_Jinkela_wire_8553),
        .dout(new_Jinkela_wire_8554)
    );

    bfr new_Jinkela_buffer_6879 (
        .din(new_Jinkela_wire_8622),
        .dout(new_Jinkela_wire_8623)
    );

    spl4L new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_7),
        .c(new_Jinkela_wire_8),
        .d(new_Jinkela_wire_9),
        .b(new_Jinkela_wire_10),
        .e(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_6823 (
        .din(new_Jinkela_wire_8554),
        .dout(new_Jinkela_wire_8555)
    );

    spl3L new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_3),
        .d(new_Jinkela_wire_4),
        .b(new_Jinkela_wire_5),
        .c(new_Jinkela_wire_6)
    );

    bfr new_Jinkela_buffer_6952 (
        .din(new_Jinkela_wire_8705),
        .dout(new_Jinkela_wire_8706)
    );

    spl4L new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_12),
        .c(new_Jinkela_wire_13),
        .d(new_Jinkela_wire_14),
        .b(new_Jinkela_wire_15),
        .e(new_Jinkela_wire_16)
    );

    bfr new_Jinkela_buffer_6824 (
        .din(new_Jinkela_wire_8555),
        .dout(new_Jinkela_wire_8556)
    );

    spl4L new_Jinkela_splitter_9 (
        .a(new_Jinkela_wire_29),
        .c(new_Jinkela_wire_30),
        .d(new_Jinkela_wire_31),
        .b(new_Jinkela_wire_32),
        .e(new_Jinkela_wire_33)
    );

    bfr new_Jinkela_buffer_6880 (
        .din(new_Jinkela_wire_8623),
        .dout(new_Jinkela_wire_8624)
    );

    spl4L new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_17),
        .c(new_Jinkela_wire_18),
        .d(new_Jinkela_wire_19),
        .b(new_Jinkela_wire_20),
        .e(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_6825 (
        .din(new_Jinkela_wire_8556),
        .dout(new_Jinkela_wire_8557)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_44),
        .dout(new_Jinkela_wire_45)
    );

    bfr new_Jinkela_buffer_7075 (
        .din(new_Jinkela_wire_8844),
        .dout(new_Jinkela_wire_8845)
    );

    spl3L new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_25),
        .d(new_Jinkela_wire_26),
        .b(new_Jinkela_wire_27),
        .c(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_6826 (
        .din(new_Jinkela_wire_8557),
        .dout(new_Jinkela_wire_8558)
    );

    bfr new_Jinkela_buffer_6881 (
        .din(new_Jinkela_wire_8624),
        .dout(new_Jinkela_wire_8625)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(N358),
        .b(new_Jinkela_wire_44),
        .c(new_Jinkela_wire_46)
    );

    bfr new_Jinkela_buffer_6827 (
        .din(new_Jinkela_wire_8558),
        .dout(new_Jinkela_wire_8559)
    );

    spl4L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_34),
        .c(new_Jinkela_wire_35),
        .d(new_Jinkela_wire_36),
        .b(new_Jinkela_wire_37),
        .e(new_Jinkela_wire_38)
    );

    spl4L new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_46),
        .c(new_Jinkela_wire_47),
        .d(new_Jinkela_wire_51),
        .b(new_Jinkela_wire_56),
        .e(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_6953 (
        .din(new_Jinkela_wire_8706),
        .dout(new_Jinkela_wire_8707)
    );

    spl4L new_Jinkela_splitter_15 (
        .a(new_Jinkela_wire_51),
        .c(new_Jinkela_wire_52),
        .d(new_Jinkela_wire_53),
        .b(new_Jinkela_wire_54),
        .e(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_6828 (
        .din(new_Jinkela_wire_8559),
        .dout(new_Jinkela_wire_8560)
    );

    spl4L new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_39),
        .c(new_Jinkela_wire_40),
        .d(new_Jinkela_wire_41),
        .b(new_Jinkela_wire_42),
        .e(new_Jinkela_wire_43)
    );

    bfr new_Jinkela_buffer_6882 (
        .din(new_Jinkela_wire_8625),
        .dout(new_Jinkela_wire_8626)
    );

    spl4L new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_66),
        .c(new_Jinkela_wire_67),
        .d(new_Jinkela_wire_68),
        .b(new_Jinkela_wire_69),
        .e(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_6829 (
        .din(new_Jinkela_wire_8560),
        .dout(new_Jinkela_wire_8561)
    );

    spl3L new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_47),
        .d(new_Jinkela_wire_48),
        .b(new_Jinkela_wire_49),
        .c(new_Jinkela_wire_50)
    );

    bfr new_Jinkela_buffer_7009 (
        .din(new_Jinkela_wire_8770),
        .dout(new_Jinkela_wire_8771)
    );

    bfr new_Jinkela_buffer_6830 (
        .din(new_Jinkela_wire_8561),
        .dout(new_Jinkela_wire_8562)
    );

    spl4L new_Jinkela_splitter_18 (
        .a(N69),
        .c(new_Jinkela_wire_66),
        .d(new_Jinkela_wire_71),
        .b(new_Jinkela_wire_76),
        .e(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_6883 (
        .din(new_Jinkela_wire_8626),
        .dout(new_Jinkela_wire_8627)
    );

    spl4L new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_56),
        .c(new_Jinkela_wire_57),
        .d(new_Jinkela_wire_58),
        .b(new_Jinkela_wire_59),
        .e(new_Jinkela_wire_60)
    );

    spl4L new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_71),
        .c(new_Jinkela_wire_72),
        .d(new_Jinkela_wire_73),
        .b(new_Jinkela_wire_74),
        .e(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_6831 (
        .din(new_Jinkela_wire_8562),
        .dout(new_Jinkela_wire_8563)
    );

    spl4L new_Jinkela_splitter_23 (
        .a(new_Jinkela_wire_86),
        .c(new_Jinkela_wire_87),
        .d(new_Jinkela_wire_92),
        .b(new_Jinkela_wire_97),
        .e(new_Jinkela_wire_102)
    );

    bfr new_Jinkela_buffer_6954 (
        .din(new_Jinkela_wire_8707),
        .dout(new_Jinkela_wire_8708)
    );

    spl4L new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_61),
        .c(new_Jinkela_wire_62),
        .d(new_Jinkela_wire_63),
        .b(new_Jinkela_wire_64),
        .e(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_6832 (
        .din(new_Jinkela_wire_8563),
        .dout(new_Jinkela_wire_8564)
    );

    bfr new_Jinkela_buffer_3 (
        .din(N18),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_6884 (
        .din(new_Jinkela_wire_8627),
        .dout(new_Jinkela_wire_8628)
    );

    spl4L new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_81),
        .c(new_Jinkela_wire_82),
        .d(new_Jinkela_wire_83),
        .b(new_Jinkela_wire_84),
        .e(new_Jinkela_wire_85)
    );

    spl4L new_Jinkela_splitter_21 (
        .a(new_Jinkela_wire_76),
        .c(new_Jinkela_wire_77),
        .d(new_Jinkela_wire_78),
        .b(new_Jinkela_wire_79),
        .e(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_6833 (
        .din(new_Jinkela_wire_8564),
        .dout(new_Jinkela_wire_8565)
    );

    spl2 new_Jinkela_splitter_735 (
        .a(_1057_),
        .b(new_Jinkela_wire_8851),
        .c(new_Jinkela_wire_8852)
    );

    spl4L new_Jinkela_splitter_24 (
        .a(new_Jinkela_wire_87),
        .c(new_Jinkela_wire_88),
        .d(new_Jinkela_wire_89),
        .b(new_Jinkela_wire_90),
        .e(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_6834 (
        .din(new_Jinkela_wire_8565),
        .dout(new_Jinkela_wire_8566)
    );

    bfr new_Jinkela_buffer_6885 (
        .din(new_Jinkela_wire_8628),
        .dout(new_Jinkela_wire_8629)
    );

    spl2 new_Jinkela_splitter_28 (
        .a(N443),
        .b(new_Jinkela_wire_107),
        .c(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_6835 (
        .din(new_Jinkela_wire_8566),
        .dout(new_Jinkela_wire_8567)
    );

    spl4L new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_97),
        .c(new_Jinkela_wire_98),
        .d(new_Jinkela_wire_99),
        .b(new_Jinkela_wire_100),
        .e(new_Jinkela_wire_101)
    );

    bfr new_Jinkela_buffer_6955 (
        .din(new_Jinkela_wire_8708),
        .dout(new_Jinkela_wire_8709)
    );

    spl4L new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_92),
        .c(new_Jinkela_wire_93),
        .d(new_Jinkela_wire_94),
        .b(new_Jinkela_wire_95),
        .e(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_6836 (
        .din(new_Jinkela_wire_8567),
        .dout(new_Jinkela_wire_8568)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_107),
        .dout(new_Jinkela_wire_108)
    );

    spl4L new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_109),
        .c(new_Jinkela_wire_110),
        .d(new_Jinkela_wire_114),
        .b(new_Jinkela_wire_119),
        .e(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_6886 (
        .din(new_Jinkela_wire_8629),
        .dout(new_Jinkela_wire_8630)
    );

    bfr new_Jinkela_buffer_6837 (
        .din(new_Jinkela_wire_8568),
        .dout(new_Jinkela_wire_8569)
    );

    spl4L new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_102),
        .c(new_Jinkela_wire_103),
        .d(new_Jinkela_wire_104),
        .b(new_Jinkela_wire_105),
        .e(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_7010 (
        .din(new_Jinkela_wire_8771),
        .dout(new_Jinkela_wire_8772)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_6838 (
        .din(new_Jinkela_wire_8569),
        .dout(new_Jinkela_wire_8570)
    );

    spl3L new_Jinkela_splitter_30 (
        .a(new_Jinkela_wire_110),
        .d(new_Jinkela_wire_111),
        .b(new_Jinkela_wire_112),
        .c(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_6887 (
        .din(new_Jinkela_wire_8630),
        .dout(new_Jinkela_wire_8631)
    );

    spl4L new_Jinkela_splitter_31 (
        .a(new_Jinkela_wire_114),
        .c(new_Jinkela_wire_115),
        .d(new_Jinkela_wire_116),
        .b(new_Jinkela_wire_117),
        .e(new_Jinkela_wire_118)
    );

    spl2 new_Jinkela_splitter_34 (
        .a(N494),
        .b(new_Jinkela_wire_129),
        .c(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_6839 (
        .din(new_Jinkela_wire_8570),
        .dout(new_Jinkela_wire_8571)
    );

    bfr new_Jinkela_buffer_6956 (
        .din(new_Jinkela_wire_8709),
        .dout(new_Jinkela_wire_8710)
    );

    spl4L new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_131),
        .c(new_Jinkela_wire_132),
        .d(new_Jinkela_wire_136),
        .b(new_Jinkela_wire_141),
        .e(new_Jinkela_wire_146)
    );

    spl4L new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_119),
        .c(new_Jinkela_wire_120),
        .d(new_Jinkela_wire_121),
        .b(new_Jinkela_wire_122),
        .e(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_6840 (
        .din(new_Jinkela_wire_8571),
        .dout(new_Jinkela_wire_8572)
    );

    bfr new_Jinkela_buffer_10 (
        .din(N171),
        .dout(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_6888 (
        .din(new_Jinkela_wire_8631),
        .dout(new_Jinkela_wire_8632)
    );

    spl4L new_Jinkela_splitter_33 (
        .a(new_Jinkela_wire_124),
        .c(new_Jinkela_wire_125),
        .d(new_Jinkela_wire_126),
        .b(new_Jinkela_wire_127),
        .e(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_6841 (
        .din(new_Jinkela_wire_8572),
        .dout(new_Jinkela_wire_8573)
    );

    spl4L new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_154),
        .c(new_Jinkela_wire_155),
        .d(new_Jinkela_wire_160),
        .b(new_Jinkela_wire_165),
        .e(new_Jinkela_wire_170)
    );

    spl2 new_Jinkela_splitter_736 (
        .a(_0142_),
        .b(new_Jinkela_wire_8853),
        .c(new_Jinkela_wire_8854)
    );

    spl2 new_Jinkela_splitter_40 (
        .a(N222),
        .b(new_Jinkela_wire_151),
        .c(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_6842 (
        .din(new_Jinkela_wire_8573),
        .dout(new_Jinkela_wire_8574)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_10474 (
        .din(new_Jinkela_wire_12651),
        .dout(new_Jinkela_wire_12652)
    );

    bfr new_Jinkela_buffer_17290 (
        .din(new_Jinkela_wire_20634),
        .dout(new_Jinkela_wire_20635)
    );

    bfr new_Jinkela_buffer_10297 (
        .din(new_Jinkela_wire_12460),
        .dout(new_Jinkela_wire_12461)
    );

    bfr new_Jinkela_buffer_17164 (
        .din(new_Jinkela_wire_20498),
        .dout(new_Jinkela_wire_20499)
    );

    bfr new_Jinkela_buffer_10414 (
        .din(new_Jinkela_wire_12581),
        .dout(new_Jinkela_wire_12582)
    );

    bfr new_Jinkela_buffer_17254 (
        .din(new_Jinkela_wire_20596),
        .dout(new_Jinkela_wire_20597)
    );

    bfr new_Jinkela_buffer_10298 (
        .din(new_Jinkela_wire_12461),
        .dout(new_Jinkela_wire_12462)
    );

    bfr new_Jinkela_buffer_17165 (
        .din(new_Jinkela_wire_20499),
        .dout(new_Jinkela_wire_20500)
    );

    bfr new_Jinkela_buffer_17331 (
        .din(new_Jinkela_wire_20679),
        .dout(new_Jinkela_wire_20680)
    );

    bfr new_Jinkela_buffer_17311 (
        .din(new_Jinkela_wire_20657),
        .dout(new_Jinkela_wire_20658)
    );

    bfr new_Jinkela_buffer_10299 (
        .din(new_Jinkela_wire_12462),
        .dout(new_Jinkela_wire_12463)
    );

    bfr new_Jinkela_buffer_17166 (
        .din(new_Jinkela_wire_20500),
        .dout(new_Jinkela_wire_20501)
    );

    bfr new_Jinkela_buffer_10415 (
        .din(new_Jinkela_wire_12582),
        .dout(new_Jinkela_wire_12583)
    );

    bfr new_Jinkela_buffer_17255 (
        .din(new_Jinkela_wire_20597),
        .dout(new_Jinkela_wire_20598)
    );

    bfr new_Jinkela_buffer_10300 (
        .din(new_Jinkela_wire_12463),
        .dout(new_Jinkela_wire_12464)
    );

    bfr new_Jinkela_buffer_17167 (
        .din(new_Jinkela_wire_20501),
        .dout(new_Jinkela_wire_20502)
    );

    bfr new_Jinkela_buffer_10475 (
        .din(new_Jinkela_wire_12652),
        .dout(new_Jinkela_wire_12653)
    );

    bfr new_Jinkela_buffer_17291 (
        .din(new_Jinkela_wire_20635),
        .dout(new_Jinkela_wire_20636)
    );

    bfr new_Jinkela_buffer_10301 (
        .din(new_Jinkela_wire_12464),
        .dout(new_Jinkela_wire_12465)
    );

    bfr new_Jinkela_buffer_17168 (
        .din(new_Jinkela_wire_20502),
        .dout(new_Jinkela_wire_20503)
    );

    bfr new_Jinkela_buffer_10416 (
        .din(new_Jinkela_wire_12583),
        .dout(new_Jinkela_wire_12584)
    );

    bfr new_Jinkela_buffer_17256 (
        .din(new_Jinkela_wire_20598),
        .dout(new_Jinkela_wire_20599)
    );

    bfr new_Jinkela_buffer_10302 (
        .din(new_Jinkela_wire_12465),
        .dout(new_Jinkela_wire_12466)
    );

    bfr new_Jinkela_buffer_17169 (
        .din(new_Jinkela_wire_20503),
        .dout(new_Jinkela_wire_20504)
    );

    bfr new_Jinkela_buffer_10543 (
        .din(new_Jinkela_wire_12742),
        .dout(new_Jinkela_wire_12743)
    );

    bfr new_Jinkela_buffer_10303 (
        .din(new_Jinkela_wire_12466),
        .dout(new_Jinkela_wire_12467)
    );

    bfr new_Jinkela_buffer_17170 (
        .din(new_Jinkela_wire_20504),
        .dout(new_Jinkela_wire_20505)
    );

    bfr new_Jinkela_buffer_10417 (
        .din(new_Jinkela_wire_12584),
        .dout(new_Jinkela_wire_12585)
    );

    bfr new_Jinkela_buffer_17257 (
        .din(new_Jinkela_wire_20599),
        .dout(new_Jinkela_wire_20600)
    );

    bfr new_Jinkela_buffer_10304 (
        .din(new_Jinkela_wire_12467),
        .dout(new_Jinkela_wire_12468)
    );

    bfr new_Jinkela_buffer_17171 (
        .din(new_Jinkela_wire_20505),
        .dout(new_Jinkela_wire_20506)
    );

    bfr new_Jinkela_buffer_10476 (
        .din(new_Jinkela_wire_12653),
        .dout(new_Jinkela_wire_12654)
    );

    bfr new_Jinkela_buffer_17292 (
        .din(new_Jinkela_wire_20636),
        .dout(new_Jinkela_wire_20637)
    );

    bfr new_Jinkela_buffer_10305 (
        .din(new_Jinkela_wire_12468),
        .dout(new_Jinkela_wire_12469)
    );

    bfr new_Jinkela_buffer_17172 (
        .din(new_Jinkela_wire_20506),
        .dout(new_Jinkela_wire_20507)
    );

    bfr new_Jinkela_buffer_10418 (
        .din(new_Jinkela_wire_12585),
        .dout(new_Jinkela_wire_12586)
    );

    bfr new_Jinkela_buffer_17258 (
        .din(new_Jinkela_wire_20600),
        .dout(new_Jinkela_wire_20601)
    );

    bfr new_Jinkela_buffer_10306 (
        .din(new_Jinkela_wire_12469),
        .dout(new_Jinkela_wire_12470)
    );

    bfr new_Jinkela_buffer_17173 (
        .din(new_Jinkela_wire_20507),
        .dout(new_Jinkela_wire_20508)
    );

    bfr new_Jinkela_buffer_10630 (
        .din(new_Jinkela_wire_12831),
        .dout(new_Jinkela_wire_12832)
    );

    bfr new_Jinkela_buffer_17335 (
        .din(new_Jinkela_wire_20683),
        .dout(new_Jinkela_wire_20684)
    );

    bfr new_Jinkela_buffer_17312 (
        .din(new_Jinkela_wire_20658),
        .dout(new_Jinkela_wire_20659)
    );

    bfr new_Jinkela_buffer_10307 (
        .din(new_Jinkela_wire_12470),
        .dout(new_Jinkela_wire_12471)
    );

    bfr new_Jinkela_buffer_17174 (
        .din(new_Jinkela_wire_20508),
        .dout(new_Jinkela_wire_20509)
    );

    bfr new_Jinkela_buffer_10419 (
        .din(new_Jinkela_wire_12586),
        .dout(new_Jinkela_wire_12587)
    );

    bfr new_Jinkela_buffer_17259 (
        .din(new_Jinkela_wire_20601),
        .dout(new_Jinkela_wire_20602)
    );

    bfr new_Jinkela_buffer_10308 (
        .din(new_Jinkela_wire_12471),
        .dout(new_Jinkela_wire_12472)
    );

    bfr new_Jinkela_buffer_17175 (
        .din(new_Jinkela_wire_20509),
        .dout(new_Jinkela_wire_20510)
    );

    bfr new_Jinkela_buffer_10477 (
        .din(new_Jinkela_wire_12654),
        .dout(new_Jinkela_wire_12655)
    );

    bfr new_Jinkela_buffer_17293 (
        .din(new_Jinkela_wire_20637),
        .dout(new_Jinkela_wire_20638)
    );

    bfr new_Jinkela_buffer_10309 (
        .din(new_Jinkela_wire_12472),
        .dout(new_Jinkela_wire_12473)
    );

    bfr new_Jinkela_buffer_17176 (
        .din(new_Jinkela_wire_20510),
        .dout(new_Jinkela_wire_20511)
    );

    bfr new_Jinkela_buffer_10420 (
        .din(new_Jinkela_wire_12587),
        .dout(new_Jinkela_wire_12588)
    );

    bfr new_Jinkela_buffer_17260 (
        .din(new_Jinkela_wire_20602),
        .dout(new_Jinkela_wire_20603)
    );

    bfr new_Jinkela_buffer_10310 (
        .din(new_Jinkela_wire_12473),
        .dout(new_Jinkela_wire_12474)
    );

    spl2 new_Jinkela_splitter_1516 (
        .a(new_Jinkela_wire_20511),
        .b(new_Jinkela_wire_20512),
        .c(new_Jinkela_wire_20513)
    );

    bfr new_Jinkela_buffer_10544 (
        .din(new_Jinkela_wire_12743),
        .dout(new_Jinkela_wire_12744)
    );

    bfr new_Jinkela_buffer_17261 (
        .din(new_Jinkela_wire_20603),
        .dout(new_Jinkela_wire_20604)
    );

    bfr new_Jinkela_buffer_10311 (
        .din(new_Jinkela_wire_12474),
        .dout(new_Jinkela_wire_12475)
    );

    bfr new_Jinkela_buffer_10421 (
        .din(new_Jinkela_wire_12588),
        .dout(new_Jinkela_wire_12589)
    );

    bfr new_Jinkela_buffer_17294 (
        .din(new_Jinkela_wire_20638),
        .dout(new_Jinkela_wire_20639)
    );

    bfr new_Jinkela_buffer_10312 (
        .din(new_Jinkela_wire_12475),
        .dout(new_Jinkela_wire_12476)
    );

    bfr new_Jinkela_buffer_17262 (
        .din(new_Jinkela_wire_20604),
        .dout(new_Jinkela_wire_20605)
    );

    bfr new_Jinkela_buffer_10478 (
        .din(new_Jinkela_wire_12655),
        .dout(new_Jinkela_wire_12656)
    );

    bfr new_Jinkela_buffer_17332 (
        .din(new_Jinkela_wire_20680),
        .dout(new_Jinkela_wire_20681)
    );

    bfr new_Jinkela_buffer_17313 (
        .din(new_Jinkela_wire_20659),
        .dout(new_Jinkela_wire_20660)
    );

    bfr new_Jinkela_buffer_10313 (
        .din(new_Jinkela_wire_12476),
        .dout(new_Jinkela_wire_12477)
    );

    bfr new_Jinkela_buffer_17263 (
        .din(new_Jinkela_wire_20605),
        .dout(new_Jinkela_wire_20606)
    );

    bfr new_Jinkela_buffer_10422 (
        .din(new_Jinkela_wire_12589),
        .dout(new_Jinkela_wire_12590)
    );

    bfr new_Jinkela_buffer_17295 (
        .din(new_Jinkela_wire_20639),
        .dout(new_Jinkela_wire_20640)
    );

    bfr new_Jinkela_buffer_10314 (
        .din(new_Jinkela_wire_12477),
        .dout(new_Jinkela_wire_12478)
    );

    bfr new_Jinkela_buffer_17264 (
        .din(new_Jinkela_wire_20606),
        .dout(new_Jinkela_wire_20607)
    );

    bfr new_Jinkela_buffer_10797 (
        .din(new_Jinkela_wire_13006),
        .dout(new_Jinkela_wire_13007)
    );

    bfr new_Jinkela_buffer_10315 (
        .din(new_Jinkela_wire_12478),
        .dout(new_Jinkela_wire_12479)
    );

    bfr new_Jinkela_buffer_17265 (
        .din(new_Jinkela_wire_20607),
        .dout(new_Jinkela_wire_20608)
    );

    bfr new_Jinkela_buffer_10423 (
        .din(new_Jinkela_wire_12590),
        .dout(new_Jinkela_wire_12591)
    );

    bfr new_Jinkela_buffer_17296 (
        .din(new_Jinkela_wire_20640),
        .dout(new_Jinkela_wire_20641)
    );

    bfr new_Jinkela_buffer_10316 (
        .din(new_Jinkela_wire_12479),
        .dout(new_Jinkela_wire_12480)
    );

    bfr new_Jinkela_buffer_17266 (
        .din(new_Jinkela_wire_20608),
        .dout(new_Jinkela_wire_20609)
    );

    bfr new_Jinkela_buffer_10479 (
        .din(new_Jinkela_wire_12656),
        .dout(new_Jinkela_wire_12657)
    );

    bfr new_Jinkela_buffer_17314 (
        .din(new_Jinkela_wire_20660),
        .dout(new_Jinkela_wire_20661)
    );

    bfr new_Jinkela_buffer_10317 (
        .din(new_Jinkela_wire_12480),
        .dout(new_Jinkela_wire_12481)
    );

    bfr new_Jinkela_buffer_17267 (
        .din(new_Jinkela_wire_20609),
        .dout(new_Jinkela_wire_20610)
    );

    bfr new_Jinkela_buffer_13817 (
        .din(new_Jinkela_wire_16482),
        .dout(new_Jinkela_wire_16483)
    );

    bfr new_Jinkela_buffer_14011 (
        .din(new_Jinkela_wire_16696),
        .dout(new_Jinkela_wire_16697)
    );

    bfr new_Jinkela_buffer_13923 (
        .din(new_Jinkela_wire_16606),
        .dout(new_Jinkela_wire_16607)
    );

    bfr new_Jinkela_buffer_13818 (
        .din(new_Jinkela_wire_16483),
        .dout(new_Jinkela_wire_16484)
    );

    bfr new_Jinkela_buffer_13864 (
        .din(new_Jinkela_wire_16545),
        .dout(new_Jinkela_wire_16546)
    );

    bfr new_Jinkela_buffer_13819 (
        .din(new_Jinkela_wire_16484),
        .dout(new_Jinkela_wire_16485)
    );

    bfr new_Jinkela_buffer_13820 (
        .din(new_Jinkela_wire_16485),
        .dout(new_Jinkela_wire_16486)
    );

    bfr new_Jinkela_buffer_13865 (
        .din(new_Jinkela_wire_16546),
        .dout(new_Jinkela_wire_16547)
    );

    bfr new_Jinkela_buffer_13821 (
        .din(new_Jinkela_wire_16486),
        .dout(new_Jinkela_wire_16487)
    );

    bfr new_Jinkela_buffer_13924 (
        .din(new_Jinkela_wire_16607),
        .dout(new_Jinkela_wire_16608)
    );

    bfr new_Jinkela_buffer_13822 (
        .din(new_Jinkela_wire_16487),
        .dout(new_Jinkela_wire_16488)
    );

    bfr new_Jinkela_buffer_13866 (
        .din(new_Jinkela_wire_16547),
        .dout(new_Jinkela_wire_16548)
    );

    bfr new_Jinkela_buffer_13823 (
        .din(new_Jinkela_wire_16488),
        .dout(new_Jinkela_wire_16489)
    );

    spl2 new_Jinkela_splitter_1194 (
        .a(_1641_),
        .b(new_Jinkela_wire_16777),
        .c(new_Jinkela_wire_16778)
    );

    bfr new_Jinkela_buffer_13824 (
        .din(new_Jinkela_wire_16489),
        .dout(new_Jinkela_wire_16490)
    );

    bfr new_Jinkela_buffer_13867 (
        .din(new_Jinkela_wire_16548),
        .dout(new_Jinkela_wire_16549)
    );

    bfr new_Jinkela_buffer_13825 (
        .din(new_Jinkela_wire_16490),
        .dout(new_Jinkela_wire_16491)
    );

    bfr new_Jinkela_buffer_14012 (
        .din(new_Jinkela_wire_16697),
        .dout(new_Jinkela_wire_16698)
    );

    bfr new_Jinkela_buffer_13925 (
        .din(new_Jinkela_wire_16608),
        .dout(new_Jinkela_wire_16609)
    );

    bfr new_Jinkela_buffer_13826 (
        .din(new_Jinkela_wire_16491),
        .dout(new_Jinkela_wire_16492)
    );

    bfr new_Jinkela_buffer_13868 (
        .din(new_Jinkela_wire_16549),
        .dout(new_Jinkela_wire_16550)
    );

    bfr new_Jinkela_buffer_13827 (
        .din(new_Jinkela_wire_16492),
        .dout(new_Jinkela_wire_16493)
    );

    bfr new_Jinkela_buffer_13828 (
        .din(new_Jinkela_wire_16493),
        .dout(new_Jinkela_wire_16494)
    );

    bfr new_Jinkela_buffer_13869 (
        .din(new_Jinkela_wire_16550),
        .dout(new_Jinkela_wire_16551)
    );

    bfr new_Jinkela_buffer_13829 (
        .din(new_Jinkela_wire_16494),
        .dout(new_Jinkela_wire_16495)
    );

    bfr new_Jinkela_buffer_14015 (
        .din(new_Jinkela_wire_16702),
        .dout(new_Jinkela_wire_16703)
    );

    bfr new_Jinkela_buffer_13926 (
        .din(new_Jinkela_wire_16609),
        .dout(new_Jinkela_wire_16610)
    );

    bfr new_Jinkela_buffer_13830 (
        .din(new_Jinkela_wire_16495),
        .dout(new_Jinkela_wire_16496)
    );

    bfr new_Jinkela_buffer_13870 (
        .din(new_Jinkela_wire_16551),
        .dout(new_Jinkela_wire_16552)
    );

    bfr new_Jinkela_buffer_13831 (
        .din(new_Jinkela_wire_16496),
        .dout(new_Jinkela_wire_16497)
    );

    bfr new_Jinkela_buffer_13832 (
        .din(new_Jinkela_wire_16497),
        .dout(new_Jinkela_wire_16498)
    );

    bfr new_Jinkela_buffer_13871 (
        .din(new_Jinkela_wire_16552),
        .dout(new_Jinkela_wire_16553)
    );

    bfr new_Jinkela_buffer_13833 (
        .din(new_Jinkela_wire_16498),
        .dout(new_Jinkela_wire_16499)
    );

    bfr new_Jinkela_buffer_14013 (
        .din(new_Jinkela_wire_16698),
        .dout(new_Jinkela_wire_16699)
    );

    bfr new_Jinkela_buffer_13927 (
        .din(new_Jinkela_wire_16610),
        .dout(new_Jinkela_wire_16611)
    );

    bfr new_Jinkela_buffer_13834 (
        .din(new_Jinkela_wire_16499),
        .dout(new_Jinkela_wire_16500)
    );

    bfr new_Jinkela_buffer_13872 (
        .din(new_Jinkela_wire_16553),
        .dout(new_Jinkela_wire_16554)
    );

    bfr new_Jinkela_buffer_13835 (
        .din(new_Jinkela_wire_16500),
        .dout(new_Jinkela_wire_16501)
    );

    bfr new_Jinkela_buffer_13836 (
        .din(new_Jinkela_wire_16501),
        .dout(new_Jinkela_wire_16502)
    );

    bfr new_Jinkela_buffer_13873 (
        .din(new_Jinkela_wire_16554),
        .dout(new_Jinkela_wire_16555)
    );

    bfr new_Jinkela_buffer_13837 (
        .din(new_Jinkela_wire_16502),
        .dout(new_Jinkela_wire_16503)
    );

    spl2 new_Jinkela_splitter_1195 (
        .a(_1728_),
        .b(new_Jinkela_wire_16779),
        .c(new_Jinkela_wire_16780)
    );

    bfr new_Jinkela_buffer_13928 (
        .din(new_Jinkela_wire_16611),
        .dout(new_Jinkela_wire_16612)
    );

    bfr new_Jinkela_buffer_6889 (
        .din(new_Jinkela_wire_8632),
        .dout(new_Jinkela_wire_8633)
    );

    bfr new_Jinkela_buffer_6843 (
        .din(new_Jinkela_wire_8574),
        .dout(new_Jinkela_wire_8575)
    );

    bfr new_Jinkela_buffer_6957 (
        .din(new_Jinkela_wire_8710),
        .dout(new_Jinkela_wire_8711)
    );

    bfr new_Jinkela_buffer_6844 (
        .din(new_Jinkela_wire_8575),
        .dout(new_Jinkela_wire_8576)
    );

    bfr new_Jinkela_buffer_6890 (
        .din(new_Jinkela_wire_8633),
        .dout(new_Jinkela_wire_8634)
    );

    bfr new_Jinkela_buffer_6845 (
        .din(new_Jinkela_wire_8576),
        .dout(new_Jinkela_wire_8577)
    );

    bfr new_Jinkela_buffer_7011 (
        .din(new_Jinkela_wire_8772),
        .dout(new_Jinkela_wire_8773)
    );

    spl2 new_Jinkela_splitter_715 (
        .a(new_Jinkela_wire_8577),
        .b(new_Jinkela_wire_8578),
        .c(new_Jinkela_wire_8579)
    );

    bfr new_Jinkela_buffer_6958 (
        .din(new_Jinkela_wire_8711),
        .dout(new_Jinkela_wire_8712)
    );

    bfr new_Jinkela_buffer_6891 (
        .din(new_Jinkela_wire_8634),
        .dout(new_Jinkela_wire_8635)
    );

    bfr new_Jinkela_buffer_6892 (
        .din(new_Jinkela_wire_8635),
        .dout(new_Jinkela_wire_8636)
    );

    bfr new_Jinkela_buffer_7076 (
        .din(new_Jinkela_wire_8845),
        .dout(new_Jinkela_wire_8846)
    );

    bfr new_Jinkela_buffer_6893 (
        .din(new_Jinkela_wire_8636),
        .dout(new_Jinkela_wire_8637)
    );

    bfr new_Jinkela_buffer_6959 (
        .din(new_Jinkela_wire_8712),
        .dout(new_Jinkela_wire_8713)
    );

    bfr new_Jinkela_buffer_6894 (
        .din(new_Jinkela_wire_8637),
        .dout(new_Jinkela_wire_8638)
    );

    bfr new_Jinkela_buffer_7012 (
        .din(new_Jinkela_wire_8773),
        .dout(new_Jinkela_wire_8774)
    );

    bfr new_Jinkela_buffer_6895 (
        .din(new_Jinkela_wire_8638),
        .dout(new_Jinkela_wire_8639)
    );

    bfr new_Jinkela_buffer_6960 (
        .din(new_Jinkela_wire_8713),
        .dout(new_Jinkela_wire_8714)
    );

    bfr new_Jinkela_buffer_6896 (
        .din(new_Jinkela_wire_8639),
        .dout(new_Jinkela_wire_8640)
    );

    bfr new_Jinkela_buffer_7093 (
        .din(_1684_),
        .dout(new_Jinkela_wire_8873)
    );

    bfr new_Jinkela_buffer_6897 (
        .din(new_Jinkela_wire_8640),
        .dout(new_Jinkela_wire_8641)
    );

    bfr new_Jinkela_buffer_6961 (
        .din(new_Jinkela_wire_8714),
        .dout(new_Jinkela_wire_8715)
    );

    bfr new_Jinkela_buffer_6898 (
        .din(new_Jinkela_wire_8641),
        .dout(new_Jinkela_wire_8642)
    );

    bfr new_Jinkela_buffer_7013 (
        .din(new_Jinkela_wire_8774),
        .dout(new_Jinkela_wire_8775)
    );

    bfr new_Jinkela_buffer_6899 (
        .din(new_Jinkela_wire_8642),
        .dout(new_Jinkela_wire_8643)
    );

    bfr new_Jinkela_buffer_6962 (
        .din(new_Jinkela_wire_8715),
        .dout(new_Jinkela_wire_8716)
    );

    bfr new_Jinkela_buffer_6900 (
        .din(new_Jinkela_wire_8643),
        .dout(new_Jinkela_wire_8644)
    );

    bfr new_Jinkela_buffer_7077 (
        .din(new_Jinkela_wire_8846),
        .dout(new_Jinkela_wire_8847)
    );

    bfr new_Jinkela_buffer_6901 (
        .din(new_Jinkela_wire_8644),
        .dout(new_Jinkela_wire_8645)
    );

    bfr new_Jinkela_buffer_6963 (
        .din(new_Jinkela_wire_8716),
        .dout(new_Jinkela_wire_8717)
    );

    bfr new_Jinkela_buffer_6902 (
        .din(new_Jinkela_wire_8645),
        .dout(new_Jinkela_wire_8646)
    );

    bfr new_Jinkela_buffer_7014 (
        .din(new_Jinkela_wire_8775),
        .dout(new_Jinkela_wire_8776)
    );

    bfr new_Jinkela_buffer_6903 (
        .din(new_Jinkela_wire_8646),
        .dout(new_Jinkela_wire_8647)
    );

    bfr new_Jinkela_buffer_6964 (
        .din(new_Jinkela_wire_8717),
        .dout(new_Jinkela_wire_8718)
    );

    bfr new_Jinkela_buffer_6904 (
        .din(new_Jinkela_wire_8647),
        .dout(new_Jinkela_wire_8648)
    );

    bfr new_Jinkela_buffer_6905 (
        .din(new_Jinkela_wire_8648),
        .dout(new_Jinkela_wire_8649)
    );

    bfr new_Jinkela_buffer_6965 (
        .din(new_Jinkela_wire_8718),
        .dout(new_Jinkela_wire_8719)
    );

    bfr new_Jinkela_buffer_6906 (
        .din(new_Jinkela_wire_8649),
        .dout(new_Jinkela_wire_8650)
    );

    bfr new_Jinkela_buffer_7015 (
        .din(new_Jinkela_wire_8776),
        .dout(new_Jinkela_wire_8777)
    );

    bfr new_Jinkela_buffer_6907 (
        .din(new_Jinkela_wire_8650),
        .dout(new_Jinkela_wire_8651)
    );

    bfr new_Jinkela_buffer_6966 (
        .din(new_Jinkela_wire_8719),
        .dout(new_Jinkela_wire_8720)
    );

    bfr new_Jinkela_buffer_3537 (
        .din(new_Jinkela_wire_4698),
        .dout(new_Jinkela_wire_4699)
    );

    bfr new_Jinkela_buffer_10424 (
        .din(new_Jinkela_wire_12591),
        .dout(new_Jinkela_wire_12592)
    );

    bfr new_Jinkela_buffer_3463 (
        .din(new_Jinkela_wire_4600),
        .dout(new_Jinkela_wire_4601)
    );

    bfr new_Jinkela_buffer_10318 (
        .din(new_Jinkela_wire_12481),
        .dout(new_Jinkela_wire_12482)
    );

    bfr new_Jinkela_buffer_10545 (
        .din(new_Jinkela_wire_12744),
        .dout(new_Jinkela_wire_12745)
    );

    spl2 new_Jinkela_splitter_431 (
        .a(_0543_),
        .b(new_Jinkela_wire_4709),
        .c(new_Jinkela_wire_4710)
    );

    bfr new_Jinkela_buffer_3464 (
        .din(new_Jinkela_wire_4601),
        .dout(new_Jinkela_wire_4602)
    );

    bfr new_Jinkela_buffer_10319 (
        .din(new_Jinkela_wire_12482),
        .dout(new_Jinkela_wire_12483)
    );

    bfr new_Jinkela_buffer_3538 (
        .din(new_Jinkela_wire_4699),
        .dout(new_Jinkela_wire_4700)
    );

    bfr new_Jinkela_buffer_10425 (
        .din(new_Jinkela_wire_12592),
        .dout(new_Jinkela_wire_12593)
    );

    bfr new_Jinkela_buffer_3465 (
        .din(new_Jinkela_wire_4602),
        .dout(new_Jinkela_wire_4603)
    );

    bfr new_Jinkela_buffer_10320 (
        .din(new_Jinkela_wire_12483),
        .dout(new_Jinkela_wire_12484)
    );

    spl2 new_Jinkela_splitter_432 (
        .a(_0485_),
        .b(new_Jinkela_wire_4711),
        .c(new_Jinkela_wire_4712)
    );

    bfr new_Jinkela_buffer_10480 (
        .din(new_Jinkela_wire_12657),
        .dout(new_Jinkela_wire_12658)
    );

    bfr new_Jinkela_buffer_3466 (
        .din(new_Jinkela_wire_4603),
        .dout(new_Jinkela_wire_4604)
    );

    bfr new_Jinkela_buffer_10321 (
        .din(new_Jinkela_wire_12484),
        .dout(new_Jinkela_wire_12485)
    );

    bfr new_Jinkela_buffer_3539 (
        .din(new_Jinkela_wire_4700),
        .dout(new_Jinkela_wire_4701)
    );

    bfr new_Jinkela_buffer_10426 (
        .din(new_Jinkela_wire_12593),
        .dout(new_Jinkela_wire_12594)
    );

    bfr new_Jinkela_buffer_3467 (
        .din(new_Jinkela_wire_4604),
        .dout(new_Jinkela_wire_4605)
    );

    bfr new_Jinkela_buffer_10322 (
        .din(new_Jinkela_wire_12485),
        .dout(new_Jinkela_wire_12486)
    );

    bfr new_Jinkela_buffer_3541 (
        .din(new_Jinkela_wire_4704),
        .dout(new_Jinkela_wire_4705)
    );

    bfr new_Jinkela_buffer_10631 (
        .din(new_Jinkela_wire_12832),
        .dout(new_Jinkela_wire_12833)
    );

    bfr new_Jinkela_buffer_3468 (
        .din(new_Jinkela_wire_4605),
        .dout(new_Jinkela_wire_4606)
    );

    bfr new_Jinkela_buffer_10323 (
        .din(new_Jinkela_wire_12486),
        .dout(new_Jinkela_wire_12487)
    );

    bfr new_Jinkela_buffer_10427 (
        .din(new_Jinkela_wire_12594),
        .dout(new_Jinkela_wire_12595)
    );

    bfr new_Jinkela_buffer_3469 (
        .din(new_Jinkela_wire_4606),
        .dout(new_Jinkela_wire_4607)
    );

    bfr new_Jinkela_buffer_10324 (
        .din(new_Jinkela_wire_12487),
        .dout(new_Jinkela_wire_12488)
    );

    bfr new_Jinkela_buffer_3542 (
        .din(new_Jinkela_wire_4705),
        .dout(new_Jinkela_wire_4706)
    );

    bfr new_Jinkela_buffer_10481 (
        .din(new_Jinkela_wire_12658),
        .dout(new_Jinkela_wire_12659)
    );

    bfr new_Jinkela_buffer_3470 (
        .din(new_Jinkela_wire_4607),
        .dout(new_Jinkela_wire_4608)
    );

    bfr new_Jinkela_buffer_10325 (
        .din(new_Jinkela_wire_12488),
        .dout(new_Jinkela_wire_12489)
    );

    bfr new_Jinkela_buffer_10428 (
        .din(new_Jinkela_wire_12595),
        .dout(new_Jinkela_wire_12596)
    );

    spl2 new_Jinkela_splitter_433 (
        .a(_1643_),
        .b(new_Jinkela_wire_4713),
        .c(new_Jinkela_wire_4714)
    );

    bfr new_Jinkela_buffer_3471 (
        .din(new_Jinkela_wire_4608),
        .dout(new_Jinkela_wire_4609)
    );

    bfr new_Jinkela_buffer_10326 (
        .din(new_Jinkela_wire_12489),
        .dout(new_Jinkela_wire_12490)
    );

    bfr new_Jinkela_buffer_3543 (
        .din(new_Jinkela_wire_4706),
        .dout(new_Jinkela_wire_4707)
    );

    bfr new_Jinkela_buffer_10546 (
        .din(new_Jinkela_wire_12745),
        .dout(new_Jinkela_wire_12746)
    );

    bfr new_Jinkela_buffer_3472 (
        .din(new_Jinkela_wire_4609),
        .dout(new_Jinkela_wire_4610)
    );

    bfr new_Jinkela_buffer_10327 (
        .din(new_Jinkela_wire_12490),
        .dout(new_Jinkela_wire_12491)
    );

    bfr new_Jinkela_buffer_10429 (
        .din(new_Jinkela_wire_12596),
        .dout(new_Jinkela_wire_12597)
    );

    spl2 new_Jinkela_splitter_434 (
        .a(_0873_),
        .b(new_Jinkela_wire_4715),
        .c(new_Jinkela_wire_4716)
    );

    bfr new_Jinkela_buffer_3473 (
        .din(new_Jinkela_wire_4610),
        .dout(new_Jinkela_wire_4611)
    );

    bfr new_Jinkela_buffer_10328 (
        .din(new_Jinkela_wire_12491),
        .dout(new_Jinkela_wire_12492)
    );

    bfr new_Jinkela_buffer_10482 (
        .din(new_Jinkela_wire_12659),
        .dout(new_Jinkela_wire_12660)
    );

    spl2 new_Jinkela_splitter_435 (
        .a(_1609_),
        .b(new_Jinkela_wire_4717),
        .c(new_Jinkela_wire_4718)
    );

    bfr new_Jinkela_buffer_3474 (
        .din(new_Jinkela_wire_4611),
        .dout(new_Jinkela_wire_4612)
    );

    bfr new_Jinkela_buffer_10329 (
        .din(new_Jinkela_wire_12492),
        .dout(new_Jinkela_wire_12493)
    );

    bfr new_Jinkela_buffer_10430 (
        .din(new_Jinkela_wire_12597),
        .dout(new_Jinkela_wire_12598)
    );

    bfr new_Jinkela_buffer_3545 (
        .din(_0902_),
        .dout(new_Jinkela_wire_4719)
    );

    bfr new_Jinkela_buffer_3475 (
        .din(new_Jinkela_wire_4612),
        .dout(new_Jinkela_wire_4613)
    );

    bfr new_Jinkela_buffer_10330 (
        .din(new_Jinkela_wire_12493),
        .dout(new_Jinkela_wire_12494)
    );

    spl2 new_Jinkela_splitter_437 (
        .a(_0083_),
        .b(new_Jinkela_wire_4722),
        .c(new_Jinkela_wire_4723)
    );

    bfr new_Jinkela_buffer_10701 (
        .din(_1562_),
        .dout(new_Jinkela_wire_12907)
    );

    spl2 new_Jinkela_splitter_436 (
        .a(_1081_),
        .b(new_Jinkela_wire_4720),
        .c(new_Jinkela_wire_4721)
    );

    spl2 new_Jinkela_splitter_953 (
        .a(_0071_),
        .b(new_Jinkela_wire_13005),
        .c(new_Jinkela_wire_13006)
    );

    bfr new_Jinkela_buffer_3476 (
        .din(new_Jinkela_wire_4613),
        .dout(new_Jinkela_wire_4614)
    );

    bfr new_Jinkela_buffer_10331 (
        .din(new_Jinkela_wire_12494),
        .dout(new_Jinkela_wire_12495)
    );

    bfr new_Jinkela_buffer_10431 (
        .din(new_Jinkela_wire_12598),
        .dout(new_Jinkela_wire_12599)
    );

    bfr new_Jinkela_buffer_3477 (
        .din(new_Jinkela_wire_4614),
        .dout(new_Jinkela_wire_4615)
    );

    bfr new_Jinkela_buffer_10332 (
        .din(new_Jinkela_wire_12495),
        .dout(new_Jinkela_wire_12496)
    );

    bfr new_Jinkela_buffer_10483 (
        .din(new_Jinkela_wire_12660),
        .dout(new_Jinkela_wire_12661)
    );

    spl2 new_Jinkela_splitter_438 (
        .a(_0159_),
        .b(new_Jinkela_wire_4724),
        .c(new_Jinkela_wire_4725)
    );

    bfr new_Jinkela_buffer_3478 (
        .din(new_Jinkela_wire_4615),
        .dout(new_Jinkela_wire_4616)
    );

    bfr new_Jinkela_buffer_10333 (
        .din(new_Jinkela_wire_12496),
        .dout(new_Jinkela_wire_12497)
    );

    bfr new_Jinkela_buffer_3569 (
        .din(new_Jinkela_wire_4750),
        .dout(new_Jinkela_wire_4751)
    );

    bfr new_Jinkela_buffer_10432 (
        .din(new_Jinkela_wire_12599),
        .dout(new_Jinkela_wire_12600)
    );

    spl2 new_Jinkela_splitter_439 (
        .a(_1305_),
        .b(new_Jinkela_wire_4726),
        .c(new_Jinkela_wire_4727)
    );

    bfr new_Jinkela_buffer_3479 (
        .din(new_Jinkela_wire_4616),
        .dout(new_Jinkela_wire_4617)
    );

    bfr new_Jinkela_buffer_10334 (
        .din(new_Jinkela_wire_12497),
        .dout(new_Jinkela_wire_12498)
    );

    bfr new_Jinkela_buffer_10547 (
        .din(new_Jinkela_wire_12746),
        .dout(new_Jinkela_wire_12747)
    );

    bfr new_Jinkela_buffer_3480 (
        .din(new_Jinkela_wire_4617),
        .dout(new_Jinkela_wire_4618)
    );

    bfr new_Jinkela_buffer_10335 (
        .din(new_Jinkela_wire_12498),
        .dout(new_Jinkela_wire_12499)
    );

    bfr new_Jinkela_buffer_10433 (
        .din(new_Jinkela_wire_12600),
        .dout(new_Jinkela_wire_12601)
    );

    bfr new_Jinkela_buffer_3481 (
        .din(new_Jinkela_wire_4618),
        .dout(new_Jinkela_wire_4619)
    );

    bfr new_Jinkela_buffer_10336 (
        .din(new_Jinkela_wire_12499),
        .dout(new_Jinkela_wire_12500)
    );

    bfr new_Jinkela_buffer_3701 (
        .din(_1756_),
        .dout(new_Jinkela_wire_4913)
    );

    bfr new_Jinkela_buffer_10484 (
        .din(new_Jinkela_wire_12661),
        .dout(new_Jinkela_wire_12662)
    );

    bfr new_Jinkela_buffer_3570 (
        .din(new_Jinkela_wire_4751),
        .dout(new_Jinkela_wire_4752)
    );

    bfr new_Jinkela_buffer_3482 (
        .din(new_Jinkela_wire_4619),
        .dout(new_Jinkela_wire_4620)
    );

    bfr new_Jinkela_buffer_10337 (
        .din(new_Jinkela_wire_12500),
        .dout(new_Jinkela_wire_12501)
    );

    bfr new_Jinkela_buffer_10434 (
        .din(new_Jinkela_wire_12601),
        .dout(new_Jinkela_wire_12602)
    );

    bfr new_Jinkela_buffer_3653 (
        .din(new_Jinkela_wire_4846),
        .dout(new_Jinkela_wire_4847)
    );

    bfr new_Jinkela_buffer_3483 (
        .din(new_Jinkela_wire_4620),
        .dout(new_Jinkela_wire_4621)
    );

    bfr new_Jinkela_buffer_10338 (
        .din(new_Jinkela_wire_12501),
        .dout(new_Jinkela_wire_12502)
    );

    bfr new_Jinkela_buffer_13838 (
        .din(new_Jinkela_wire_16503),
        .dout(new_Jinkela_wire_16504)
    );

    bfr new_Jinkela_buffer_13874 (
        .din(new_Jinkela_wire_16555),
        .dout(new_Jinkela_wire_16556)
    );

    bfr new_Jinkela_buffer_13839 (
        .din(new_Jinkela_wire_16504),
        .dout(new_Jinkela_wire_16505)
    );

    spl2 new_Jinkela_splitter_1182 (
        .a(new_Jinkela_wire_16505),
        .b(new_Jinkela_wire_16506),
        .c(new_Jinkela_wire_16507)
    );

    bfr new_Jinkela_buffer_14016 (
        .din(new_Jinkela_wire_16703),
        .dout(new_Jinkela_wire_16704)
    );

    bfr new_Jinkela_buffer_13929 (
        .din(new_Jinkela_wire_16612),
        .dout(new_Jinkela_wire_16613)
    );

    bfr new_Jinkela_buffer_13875 (
        .din(new_Jinkela_wire_16556),
        .dout(new_Jinkela_wire_16557)
    );

    bfr new_Jinkela_buffer_13876 (
        .din(new_Jinkela_wire_16557),
        .dout(new_Jinkela_wire_16558)
    );

    bfr new_Jinkela_buffer_13877 (
        .din(new_Jinkela_wire_16558),
        .dout(new_Jinkela_wire_16559)
    );

    bfr new_Jinkela_buffer_13930 (
        .din(new_Jinkela_wire_16613),
        .dout(new_Jinkela_wire_16614)
    );

    bfr new_Jinkela_buffer_13878 (
        .din(new_Jinkela_wire_16559),
        .dout(new_Jinkela_wire_16560)
    );

    bfr new_Jinkela_buffer_13879 (
        .din(new_Jinkela_wire_16560),
        .dout(new_Jinkela_wire_16561)
    );

    bfr new_Jinkela_buffer_14017 (
        .din(new_Jinkela_wire_16704),
        .dout(new_Jinkela_wire_16705)
    );

    bfr new_Jinkela_buffer_13931 (
        .din(new_Jinkela_wire_16614),
        .dout(new_Jinkela_wire_16615)
    );

    bfr new_Jinkela_buffer_13880 (
        .din(new_Jinkela_wire_16561),
        .dout(new_Jinkela_wire_16562)
    );

    bfr new_Jinkela_buffer_13881 (
        .din(new_Jinkela_wire_16562),
        .dout(new_Jinkela_wire_16563)
    );

    bfr new_Jinkela_buffer_13932 (
        .din(new_Jinkela_wire_16615),
        .dout(new_Jinkela_wire_16616)
    );

    bfr new_Jinkela_buffer_13882 (
        .din(new_Jinkela_wire_16563),
        .dout(new_Jinkela_wire_16564)
    );

    spl2 new_Jinkela_splitter_1196 (
        .a(_0081_),
        .b(new_Jinkela_wire_16781),
        .c(new_Jinkela_wire_16782)
    );

    bfr new_Jinkela_buffer_13883 (
        .din(new_Jinkela_wire_16564),
        .dout(new_Jinkela_wire_16565)
    );

    bfr new_Jinkela_buffer_14018 (
        .din(new_Jinkela_wire_16705),
        .dout(new_Jinkela_wire_16706)
    );

    bfr new_Jinkela_buffer_13933 (
        .din(new_Jinkela_wire_16616),
        .dout(new_Jinkela_wire_16617)
    );

    bfr new_Jinkela_buffer_13884 (
        .din(new_Jinkela_wire_16565),
        .dout(new_Jinkela_wire_16566)
    );

    bfr new_Jinkela_buffer_13885 (
        .din(new_Jinkela_wire_16566),
        .dout(new_Jinkela_wire_16567)
    );

    bfr new_Jinkela_buffer_14087 (
        .din(new_Jinkela_wire_16784),
        .dout(new_Jinkela_wire_16785)
    );

    bfr new_Jinkela_buffer_13934 (
        .din(new_Jinkela_wire_16617),
        .dout(new_Jinkela_wire_16618)
    );

    bfr new_Jinkela_buffer_13886 (
        .din(new_Jinkela_wire_16567),
        .dout(new_Jinkela_wire_16568)
    );

    spl2 new_Jinkela_splitter_1197 (
        .a(_1765_),
        .b(new_Jinkela_wire_16783),
        .c(new_Jinkela_wire_16784)
    );

    bfr new_Jinkela_buffer_13887 (
        .din(new_Jinkela_wire_16568),
        .dout(new_Jinkela_wire_16569)
    );

    bfr new_Jinkela_buffer_14019 (
        .din(new_Jinkela_wire_16706),
        .dout(new_Jinkela_wire_16707)
    );

    bfr new_Jinkela_buffer_13935 (
        .din(new_Jinkela_wire_16618),
        .dout(new_Jinkela_wire_16619)
    );

    bfr new_Jinkela_buffer_13888 (
        .din(new_Jinkela_wire_16569),
        .dout(new_Jinkela_wire_16570)
    );

    bfr new_Jinkela_buffer_13889 (
        .din(new_Jinkela_wire_16570),
        .dout(new_Jinkela_wire_16571)
    );

    bfr new_Jinkela_buffer_13936 (
        .din(new_Jinkela_wire_16619),
        .dout(new_Jinkela_wire_16620)
    );

    bfr new_Jinkela_buffer_13890 (
        .din(new_Jinkela_wire_16571),
        .dout(new_Jinkela_wire_16572)
    );

    bfr new_Jinkela_buffer_14091 (
        .din(_1806_),
        .dout(new_Jinkela_wire_16789)
    );

    bfr new_Jinkela_buffer_13891 (
        .din(new_Jinkela_wire_16572),
        .dout(new_Jinkela_wire_16573)
    );

    bfr new_Jinkela_buffer_14020 (
        .din(new_Jinkela_wire_16707),
        .dout(new_Jinkela_wire_16708)
    );

    bfr new_Jinkela_buffer_13937 (
        .din(new_Jinkela_wire_16620),
        .dout(new_Jinkela_wire_16621)
    );

    bfr new_Jinkela_buffer_13892 (
        .din(new_Jinkela_wire_16573),
        .dout(new_Jinkela_wire_16574)
    );

    bfr new_Jinkela_buffer_13893 (
        .din(new_Jinkela_wire_16574),
        .dout(new_Jinkela_wire_16575)
    );

    spl4L new_Jinkela_splitter_38 (
        .a(new_Jinkela_wire_141),
        .c(new_Jinkela_wire_142),
        .d(new_Jinkela_wire_143),
        .b(new_Jinkela_wire_144),
        .e(new_Jinkela_wire_145)
    );

    spl4L new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_136),
        .c(new_Jinkela_wire_137),
        .d(new_Jinkela_wire_138),
        .b(new_Jinkela_wire_139),
        .e(new_Jinkela_wire_140)
    );

    spl3L new_Jinkela_splitter_36 (
        .a(new_Jinkela_wire_132),
        .d(new_Jinkela_wire_133),
        .b(new_Jinkela_wire_134),
        .c(new_Jinkela_wire_135)
    );

    spl4L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_160),
        .c(new_Jinkela_wire_161),
        .d(new_Jinkela_wire_162),
        .b(new_Jinkela_wire_163),
        .e(new_Jinkela_wire_164)
    );

    spl4L new_Jinkela_splitter_39 (
        .a(new_Jinkela_wire_146),
        .c(new_Jinkela_wire_147),
        .d(new_Jinkela_wire_148),
        .b(new_Jinkela_wire_149),
        .e(new_Jinkela_wire_150)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_177),
        .c(new_Jinkela_wire_178),
        .d(new_Jinkela_wire_183),
        .b(new_Jinkela_wire_188),
        .e(new_Jinkela_wire_193)
    );

    spl4L new_Jinkela_splitter_48 (
        .a(new_Jinkela_wire_183),
        .c(new_Jinkela_wire_184),
        .d(new_Jinkela_wire_185),
        .b(new_Jinkela_wire_186),
        .e(new_Jinkela_wire_187)
    );

    spl4L new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_155),
        .c(new_Jinkela_wire_156),
        .d(new_Jinkela_wire_157),
        .b(new_Jinkela_wire_158),
        .e(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    spl4L new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_165),
        .c(new_Jinkela_wire_166),
        .d(new_Jinkela_wire_167),
        .b(new_Jinkela_wire_168),
        .e(new_Jinkela_wire_169)
    );

    spl4L new_Jinkela_splitter_45 (
        .a(new_Jinkela_wire_170),
        .c(new_Jinkela_wire_171),
        .d(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_173),
        .e(new_Jinkela_wire_174)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(N477),
        .b(new_Jinkela_wire_198),
        .c(new_Jinkela_wire_200)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    spl4L new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_178),
        .c(new_Jinkela_wire_179),
        .d(new_Jinkela_wire_180),
        .b(new_Jinkela_wire_181),
        .e(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    spl4L new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_200),
        .c(new_Jinkela_wire_201),
        .d(new_Jinkela_wire_205),
        .b(new_Jinkela_wire_210),
        .e(new_Jinkela_wire_215)
    );

    spl4L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_188),
        .c(new_Jinkela_wire_189),
        .d(new_Jinkela_wire_190),
        .b(new_Jinkela_wire_191),
        .e(new_Jinkela_wire_192)
    );

    spl4L new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_193),
        .c(new_Jinkela_wire_194),
        .d(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_196),
        .e(new_Jinkela_wire_197)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    spl3L new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_201),
        .d(new_Jinkela_wire_202),
        .b(new_Jinkela_wire_203),
        .c(new_Jinkela_wire_204)
    );

    spl4L new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_270),
        .c(new_Jinkela_wire_271),
        .d(new_Jinkela_wire_272),
        .b(new_Jinkela_wire_273),
        .e(new_Jinkela_wire_274)
    );

    spl4L new_Jinkela_splitter_54 (
        .a(new_Jinkela_wire_205),
        .c(new_Jinkela_wire_206),
        .d(new_Jinkela_wire_207),
        .b(new_Jinkela_wire_208),
        .e(new_Jinkela_wire_209)
    );

    spl2 new_Jinkela_splitter_57 (
        .a(N273),
        .b(new_Jinkela_wire_220),
        .c(new_Jinkela_wire_222)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_222),
        .c(new_Jinkela_wire_223),
        .d(new_Jinkela_wire_227),
        .b(new_Jinkela_wire_232),
        .e(new_Jinkela_wire_237)
    );

    spl4L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_210),
        .c(new_Jinkela_wire_211),
        .d(new_Jinkela_wire_212),
        .b(new_Jinkela_wire_213),
        .e(new_Jinkela_wire_214)
    );

    spl4L new_Jinkela_splitter_60 (
        .a(new_Jinkela_wire_227),
        .c(new_Jinkela_wire_228),
        .d(new_Jinkela_wire_229),
        .b(new_Jinkela_wire_230),
        .e(new_Jinkela_wire_231)
    );

    spl4L new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_215),
        .c(new_Jinkela_wire_216),
        .d(new_Jinkela_wire_217),
        .b(new_Jinkela_wire_218),
        .e(new_Jinkela_wire_219)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_242),
        .dout(new_Jinkela_wire_243)
    );

    spl3L new_Jinkela_splitter_59 (
        .a(new_Jinkela_wire_223),
        .d(new_Jinkela_wire_224),
        .b(new_Jinkela_wire_225),
        .c(new_Jinkela_wire_226)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(N392),
        .b(new_Jinkela_wire_242),
        .c(new_Jinkela_wire_244)
    );

    spl4L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_232),
        .c(new_Jinkela_wire_233),
        .d(new_Jinkela_wire_234),
        .b(new_Jinkela_wire_235),
        .e(new_Jinkela_wire_236)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_244),
        .c(new_Jinkela_wire_245),
        .d(new_Jinkela_wire_249),
        .b(new_Jinkela_wire_254),
        .e(new_Jinkela_wire_259)
    );

    spl4L new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_249),
        .c(new_Jinkela_wire_250),
        .d(new_Jinkela_wire_251),
        .b(new_Jinkela_wire_252),
        .e(new_Jinkela_wire_253)
    );

    spl2 new_Jinkela_splitter_80 (
        .a(N290),
        .b(new_Jinkela_wire_307),
        .c(new_Jinkela_wire_311)
    );

    spl4L new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_237),
        .c(new_Jinkela_wire_238),
        .d(new_Jinkela_wire_239),
        .b(new_Jinkela_wire_240),
        .e(new_Jinkela_wire_241)
    );

    spl4L new_Jinkela_splitter_69 (
        .a(new_Jinkela_wire_264),
        .c(new_Jinkela_wire_265),
        .d(new_Jinkela_wire_270),
        .b(new_Jinkela_wire_275),
        .e(new_Jinkela_wire_280)
    );

    spl3L new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_245),
        .d(new_Jinkela_wire_246),
        .b(new_Jinkela_wire_247),
        .c(new_Jinkela_wire_248)
    );

    bfr new_Jinkela_buffer_14 (
        .din(N52),
        .dout(new_Jinkela_wire_264)
    );

    spl4L new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_254),
        .c(new_Jinkela_wire_255),
        .d(new_Jinkela_wire_256),
        .b(new_Jinkela_wire_257),
        .e(new_Jinkela_wire_258)
    );

    spl4L new_Jinkela_splitter_75 (
        .a(new_Jinkela_wire_287),
        .c(new_Jinkela_wire_288),
        .d(new_Jinkela_wire_292),
        .b(new_Jinkela_wire_297),
        .e(new_Jinkela_wire_302)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(N375),
        .b(new_Jinkela_wire_285),
        .c(new_Jinkela_wire_287)
    );

    spl4L new_Jinkela_splitter_68 (
        .a(new_Jinkela_wire_259),
        .c(new_Jinkela_wire_260),
        .d(new_Jinkela_wire_261),
        .b(new_Jinkela_wire_262),
        .e(new_Jinkela_wire_263)
    );

    spl2 new_Jinkela_splitter_441 (
        .a(_0215_),
        .b(new_Jinkela_wire_4826),
        .c(new_Jinkela_wire_4827)
    );

    bfr new_Jinkela_buffer_3484 (
        .din(new_Jinkela_wire_4621),
        .dout(new_Jinkela_wire_4622)
    );

    bfr new_Jinkela_buffer_3642 (
        .din(_0871_),
        .dout(new_Jinkela_wire_4828)
    );

    bfr new_Jinkela_buffer_3485 (
        .din(new_Jinkela_wire_4622),
        .dout(new_Jinkela_wire_4623)
    );

    bfr new_Jinkela_buffer_3547 (
        .din(new_Jinkela_wire_4728),
        .dout(new_Jinkela_wire_4729)
    );

    bfr new_Jinkela_buffer_3486 (
        .din(new_Jinkela_wire_4623),
        .dout(new_Jinkela_wire_4624)
    );

    bfr new_Jinkela_buffer_3487 (
        .din(new_Jinkela_wire_4624),
        .dout(new_Jinkela_wire_4625)
    );

    bfr new_Jinkela_buffer_3548 (
        .din(new_Jinkela_wire_4729),
        .dout(new_Jinkela_wire_4730)
    );

    bfr new_Jinkela_buffer_3488 (
        .din(new_Jinkela_wire_4625),
        .dout(new_Jinkela_wire_4626)
    );

    spl2 new_Jinkela_splitter_443 (
        .a(_1382_),
        .b(new_Jinkela_wire_4831),
        .c(new_Jinkela_wire_4832)
    );

    spl2 new_Jinkela_splitter_442 (
        .a(_1159_),
        .b(new_Jinkela_wire_4829),
        .c(new_Jinkela_wire_4830)
    );

    bfr new_Jinkela_buffer_3489 (
        .din(new_Jinkela_wire_4626),
        .dout(new_Jinkela_wire_4627)
    );

    bfr new_Jinkela_buffer_3549 (
        .din(new_Jinkela_wire_4730),
        .dout(new_Jinkela_wire_4731)
    );

    bfr new_Jinkela_buffer_3490 (
        .din(new_Jinkela_wire_4627),
        .dout(new_Jinkela_wire_4628)
    );

    bfr new_Jinkela_buffer_3491 (
        .din(new_Jinkela_wire_4628),
        .dout(new_Jinkela_wire_4629)
    );

    bfr new_Jinkela_buffer_3550 (
        .din(new_Jinkela_wire_4731),
        .dout(new_Jinkela_wire_4732)
    );

    bfr new_Jinkela_buffer_3492 (
        .din(new_Jinkela_wire_4629),
        .dout(new_Jinkela_wire_4630)
    );

    bfr new_Jinkela_buffer_3643 (
        .din(_1741_),
        .dout(new_Jinkela_wire_4833)
    );

    bfr new_Jinkela_buffer_3493 (
        .din(new_Jinkela_wire_4630),
        .dout(new_Jinkela_wire_4631)
    );

    bfr new_Jinkela_buffer_3551 (
        .din(new_Jinkela_wire_4732),
        .dout(new_Jinkela_wire_4733)
    );

    bfr new_Jinkela_buffer_3494 (
        .din(new_Jinkela_wire_4631),
        .dout(new_Jinkela_wire_4632)
    );

    spl2 new_Jinkela_splitter_445 (
        .a(_1120_),
        .b(new_Jinkela_wire_4836),
        .c(new_Jinkela_wire_4837)
    );

    spl2 new_Jinkela_splitter_444 (
        .a(_1734_),
        .b(new_Jinkela_wire_4834),
        .c(new_Jinkela_wire_4835)
    );

    bfr new_Jinkela_buffer_3495 (
        .din(new_Jinkela_wire_4632),
        .dout(new_Jinkela_wire_4633)
    );

    bfr new_Jinkela_buffer_3552 (
        .din(new_Jinkela_wire_4733),
        .dout(new_Jinkela_wire_4734)
    );

    bfr new_Jinkela_buffer_3496 (
        .din(new_Jinkela_wire_4633),
        .dout(new_Jinkela_wire_4634)
    );

    bfr new_Jinkela_buffer_3497 (
        .din(new_Jinkela_wire_4634),
        .dout(new_Jinkela_wire_4635)
    );

    bfr new_Jinkela_buffer_3553 (
        .din(new_Jinkela_wire_4734),
        .dout(new_Jinkela_wire_4735)
    );

    bfr new_Jinkela_buffer_3498 (
        .din(new_Jinkela_wire_4635),
        .dout(new_Jinkela_wire_4636)
    );

    bfr new_Jinkela_buffer_3644 (
        .din(_0075_),
        .dout(new_Jinkela_wire_4838)
    );

    bfr new_Jinkela_buffer_3499 (
        .din(new_Jinkela_wire_4636),
        .dout(new_Jinkela_wire_4637)
    );

    bfr new_Jinkela_buffer_3554 (
        .din(new_Jinkela_wire_4735),
        .dout(new_Jinkela_wire_4736)
    );

    bfr new_Jinkela_buffer_3500 (
        .din(new_Jinkela_wire_4637),
        .dout(new_Jinkela_wire_4638)
    );

    spl2 new_Jinkela_splitter_447 (
        .a(_0907_),
        .b(new_Jinkela_wire_4897),
        .c(new_Jinkela_wire_4898)
    );

    bfr new_Jinkela_buffer_3645 (
        .din(_0100_),
        .dout(new_Jinkela_wire_4839)
    );

    bfr new_Jinkela_buffer_3501 (
        .din(new_Jinkela_wire_4638),
        .dout(new_Jinkela_wire_4639)
    );

    bfr new_Jinkela_buffer_3555 (
        .din(new_Jinkela_wire_4736),
        .dout(new_Jinkela_wire_4737)
    );

    bfr new_Jinkela_buffer_3502 (
        .din(new_Jinkela_wire_4639),
        .dout(new_Jinkela_wire_4640)
    );

    spl2 new_Jinkela_splitter_448 (
        .a(_0638_),
        .b(new_Jinkela_wire_4899),
        .c(new_Jinkela_wire_4900)
    );

    bfr new_Jinkela_buffer_3503 (
        .din(new_Jinkela_wire_4640),
        .dout(new_Jinkela_wire_4641)
    );

    bfr new_Jinkela_buffer_3556 (
        .din(new_Jinkela_wire_4737),
        .dout(new_Jinkela_wire_4738)
    );

    bfr new_Jinkela_buffer_3546 (
        .din(_0331_),
        .dout(new_Jinkela_wire_4728)
    );

    bfr new_Jinkela_buffer_3504 (
        .din(new_Jinkela_wire_4641),
        .dout(new_Jinkela_wire_4642)
    );

    bfr new_Jinkela_buffer_10632 (
        .din(new_Jinkela_wire_12833),
        .dout(new_Jinkela_wire_12834)
    );

    bfr new_Jinkela_buffer_10339 (
        .din(new_Jinkela_wire_12502),
        .dout(new_Jinkela_wire_12503)
    );

    bfr new_Jinkela_buffer_10435 (
        .din(new_Jinkela_wire_12602),
        .dout(new_Jinkela_wire_12603)
    );

    bfr new_Jinkela_buffer_10340 (
        .din(new_Jinkela_wire_12503),
        .dout(new_Jinkela_wire_12504)
    );

    bfr new_Jinkela_buffer_10485 (
        .din(new_Jinkela_wire_12662),
        .dout(new_Jinkela_wire_12663)
    );

    bfr new_Jinkela_buffer_10341 (
        .din(new_Jinkela_wire_12504),
        .dout(new_Jinkela_wire_12505)
    );

    bfr new_Jinkela_buffer_10436 (
        .din(new_Jinkela_wire_12603),
        .dout(new_Jinkela_wire_12604)
    );

    bfr new_Jinkela_buffer_10342 (
        .din(new_Jinkela_wire_12505),
        .dout(new_Jinkela_wire_12506)
    );

    bfr new_Jinkela_buffer_10548 (
        .din(new_Jinkela_wire_12747),
        .dout(new_Jinkela_wire_12748)
    );

    bfr new_Jinkela_buffer_10343 (
        .din(new_Jinkela_wire_12506),
        .dout(new_Jinkela_wire_12507)
    );

    bfr new_Jinkela_buffer_10437 (
        .din(new_Jinkela_wire_12604),
        .dout(new_Jinkela_wire_12605)
    );

    bfr new_Jinkela_buffer_10344 (
        .din(new_Jinkela_wire_12507),
        .dout(new_Jinkela_wire_12508)
    );

    bfr new_Jinkela_buffer_10486 (
        .din(new_Jinkela_wire_12663),
        .dout(new_Jinkela_wire_12664)
    );

    bfr new_Jinkela_buffer_10345 (
        .din(new_Jinkela_wire_12508),
        .dout(new_Jinkela_wire_12509)
    );

    bfr new_Jinkela_buffer_10438 (
        .din(new_Jinkela_wire_12605),
        .dout(new_Jinkela_wire_12606)
    );

    bfr new_Jinkela_buffer_10346 (
        .din(new_Jinkela_wire_12509),
        .dout(new_Jinkela_wire_12510)
    );

    bfr new_Jinkela_buffer_10702 (
        .din(new_Jinkela_wire_12907),
        .dout(new_Jinkela_wire_12908)
    );

    bfr new_Jinkela_buffer_10347 (
        .din(new_Jinkela_wire_12510),
        .dout(new_Jinkela_wire_12511)
    );

    bfr new_Jinkela_buffer_10439 (
        .din(new_Jinkela_wire_12606),
        .dout(new_Jinkela_wire_12607)
    );

    bfr new_Jinkela_buffer_10348 (
        .din(new_Jinkela_wire_12511),
        .dout(new_Jinkela_wire_12512)
    );

    bfr new_Jinkela_buffer_10487 (
        .din(new_Jinkela_wire_12664),
        .dout(new_Jinkela_wire_12665)
    );

    bfr new_Jinkela_buffer_10349 (
        .din(new_Jinkela_wire_12512),
        .dout(new_Jinkela_wire_12513)
    );

    bfr new_Jinkela_buffer_10440 (
        .din(new_Jinkela_wire_12607),
        .dout(new_Jinkela_wire_12608)
    );

    bfr new_Jinkela_buffer_10350 (
        .din(new_Jinkela_wire_12513),
        .dout(new_Jinkela_wire_12514)
    );

    bfr new_Jinkela_buffer_10549 (
        .din(new_Jinkela_wire_12748),
        .dout(new_Jinkela_wire_12749)
    );

    bfr new_Jinkela_buffer_10351 (
        .din(new_Jinkela_wire_12514),
        .dout(new_Jinkela_wire_12515)
    );

    bfr new_Jinkela_buffer_10441 (
        .din(new_Jinkela_wire_12608),
        .dout(new_Jinkela_wire_12609)
    );

    bfr new_Jinkela_buffer_10352 (
        .din(new_Jinkela_wire_12515),
        .dout(new_Jinkela_wire_12516)
    );

    bfr new_Jinkela_buffer_10488 (
        .din(new_Jinkela_wire_12665),
        .dout(new_Jinkela_wire_12666)
    );

    bfr new_Jinkela_buffer_10353 (
        .din(new_Jinkela_wire_12516),
        .dout(new_Jinkela_wire_12517)
    );

    bfr new_Jinkela_buffer_10442 (
        .din(new_Jinkela_wire_12609),
        .dout(new_Jinkela_wire_12610)
    );

    bfr new_Jinkela_buffer_10354 (
        .din(new_Jinkela_wire_12517),
        .dout(new_Jinkela_wire_12518)
    );

    bfr new_Jinkela_buffer_10633 (
        .din(new_Jinkela_wire_12834),
        .dout(new_Jinkela_wire_12835)
    );

    bfr new_Jinkela_buffer_10355 (
        .din(new_Jinkela_wire_12518),
        .dout(new_Jinkela_wire_12519)
    );

    bfr new_Jinkela_buffer_10443 (
        .din(new_Jinkela_wire_12610),
        .dout(new_Jinkela_wire_12611)
    );

    bfr new_Jinkela_buffer_10489 (
        .din(new_Jinkela_wire_12666),
        .dout(new_Jinkela_wire_12667)
    );

    bfr new_Jinkela_buffer_10444 (
        .din(new_Jinkela_wire_12611),
        .dout(new_Jinkela_wire_12612)
    );

    bfr new_Jinkela_buffer_10550 (
        .din(new_Jinkela_wire_12749),
        .dout(new_Jinkela_wire_12750)
    );

    spl2 new_Jinkela_splitter_933 (
        .a(new_Jinkela_wire_12612),
        .b(new_Jinkela_wire_12613),
        .c(new_Jinkela_wire_12614)
    );

    bfr new_Jinkela_buffer_10801 (
        .din(_1427_),
        .dout(new_Jinkela_wire_13011)
    );

    bfr new_Jinkela_buffer_10490 (
        .din(new_Jinkela_wire_12667),
        .dout(new_Jinkela_wire_12668)
    );

    bfr new_Jinkela_buffer_10491 (
        .din(new_Jinkela_wire_12668),
        .dout(new_Jinkela_wire_12669)
    );

    bfr new_Jinkela_buffer_6908 (
        .din(new_Jinkela_wire_8651),
        .dout(new_Jinkela_wire_8652)
    );

    bfr new_Jinkela_buffer_7078 (
        .din(new_Jinkela_wire_8847),
        .dout(new_Jinkela_wire_8848)
    );

    bfr new_Jinkela_buffer_6909 (
        .din(new_Jinkela_wire_8652),
        .dout(new_Jinkela_wire_8653)
    );

    bfr new_Jinkela_buffer_6967 (
        .din(new_Jinkela_wire_8720),
        .dout(new_Jinkela_wire_8721)
    );

    bfr new_Jinkela_buffer_6910 (
        .din(new_Jinkela_wire_8653),
        .dout(new_Jinkela_wire_8654)
    );

    bfr new_Jinkela_buffer_7016 (
        .din(new_Jinkela_wire_8777),
        .dout(new_Jinkela_wire_8778)
    );

    bfr new_Jinkela_buffer_6911 (
        .din(new_Jinkela_wire_8654),
        .dout(new_Jinkela_wire_8655)
    );

    bfr new_Jinkela_buffer_6968 (
        .din(new_Jinkela_wire_8721),
        .dout(new_Jinkela_wire_8722)
    );

    bfr new_Jinkela_buffer_6912 (
        .din(new_Jinkela_wire_8655),
        .dout(new_Jinkela_wire_8656)
    );

    bfr new_Jinkela_buffer_7087 (
        .din(_0158_),
        .dout(new_Jinkela_wire_8865)
    );

    bfr new_Jinkela_buffer_6913 (
        .din(new_Jinkela_wire_8656),
        .dout(new_Jinkela_wire_8657)
    );

    bfr new_Jinkela_buffer_6969 (
        .din(new_Jinkela_wire_8722),
        .dout(new_Jinkela_wire_8723)
    );

    bfr new_Jinkela_buffer_6914 (
        .din(new_Jinkela_wire_8657),
        .dout(new_Jinkela_wire_8658)
    );

    bfr new_Jinkela_buffer_7017 (
        .din(new_Jinkela_wire_8778),
        .dout(new_Jinkela_wire_8779)
    );

    bfr new_Jinkela_buffer_6915 (
        .din(new_Jinkela_wire_8658),
        .dout(new_Jinkela_wire_8659)
    );

    bfr new_Jinkela_buffer_6970 (
        .din(new_Jinkela_wire_8723),
        .dout(new_Jinkela_wire_8724)
    );

    bfr new_Jinkela_buffer_6916 (
        .din(new_Jinkela_wire_8659),
        .dout(new_Jinkela_wire_8660)
    );

    bfr new_Jinkela_buffer_7088 (
        .din(_1481_),
        .dout(new_Jinkela_wire_8866)
    );

    bfr new_Jinkela_buffer_6917 (
        .din(new_Jinkela_wire_8660),
        .dout(new_Jinkela_wire_8661)
    );

    bfr new_Jinkela_buffer_6971 (
        .din(new_Jinkela_wire_8724),
        .dout(new_Jinkela_wire_8725)
    );

    bfr new_Jinkela_buffer_6918 (
        .din(new_Jinkela_wire_8661),
        .dout(new_Jinkela_wire_8662)
    );

    bfr new_Jinkela_buffer_7018 (
        .din(new_Jinkela_wire_8779),
        .dout(new_Jinkela_wire_8780)
    );

    bfr new_Jinkela_buffer_6919 (
        .din(new_Jinkela_wire_8662),
        .dout(new_Jinkela_wire_8663)
    );

    bfr new_Jinkela_buffer_6972 (
        .din(new_Jinkela_wire_8725),
        .dout(new_Jinkela_wire_8726)
    );

    bfr new_Jinkela_buffer_6920 (
        .din(new_Jinkela_wire_8663),
        .dout(new_Jinkela_wire_8664)
    );

    bfr new_Jinkela_buffer_7080 (
        .din(new_Jinkela_wire_8855),
        .dout(new_Jinkela_wire_8856)
    );

    bfr new_Jinkela_buffer_6921 (
        .din(new_Jinkela_wire_8664),
        .dout(new_Jinkela_wire_8665)
    );

    bfr new_Jinkela_buffer_6973 (
        .din(new_Jinkela_wire_8726),
        .dout(new_Jinkela_wire_8727)
    );

    bfr new_Jinkela_buffer_6922 (
        .din(new_Jinkela_wire_8665),
        .dout(new_Jinkela_wire_8666)
    );

    bfr new_Jinkela_buffer_7019 (
        .din(new_Jinkela_wire_8780),
        .dout(new_Jinkela_wire_8781)
    );

    bfr new_Jinkela_buffer_6923 (
        .din(new_Jinkela_wire_8666),
        .dout(new_Jinkela_wire_8667)
    );

    bfr new_Jinkela_buffer_6974 (
        .din(new_Jinkela_wire_8727),
        .dout(new_Jinkela_wire_8728)
    );

    bfr new_Jinkela_buffer_6924 (
        .din(new_Jinkela_wire_8667),
        .dout(new_Jinkela_wire_8668)
    );

    spl2 new_Jinkela_splitter_738 (
        .a(_1529_),
        .b(new_Jinkela_wire_8867),
        .c(new_Jinkela_wire_8868)
    );

    bfr new_Jinkela_buffer_6925 (
        .din(new_Jinkela_wire_8668),
        .dout(new_Jinkela_wire_8669)
    );

    bfr new_Jinkela_buffer_6975 (
        .din(new_Jinkela_wire_8728),
        .dout(new_Jinkela_wire_8729)
    );

    bfr new_Jinkela_buffer_6926 (
        .din(new_Jinkela_wire_8669),
        .dout(new_Jinkela_wire_8670)
    );

    bfr new_Jinkela_buffer_7020 (
        .din(new_Jinkela_wire_8781),
        .dout(new_Jinkela_wire_8782)
    );

    bfr new_Jinkela_buffer_6927 (
        .din(new_Jinkela_wire_8670),
        .dout(new_Jinkela_wire_8671)
    );

    bfr new_Jinkela_buffer_6976 (
        .din(new_Jinkela_wire_8729),
        .dout(new_Jinkela_wire_8730)
    );

    bfr new_Jinkela_buffer_6928 (
        .din(new_Jinkela_wire_8671),
        .dout(new_Jinkela_wire_8672)
    );

    bfr new_Jinkela_buffer_7081 (
        .din(new_Jinkela_wire_8856),
        .dout(new_Jinkela_wire_8857)
    );

    bfr new_Jinkela_buffer_7079 (
        .din(_1632_),
        .dout(new_Jinkela_wire_8855)
    );

    bfr new_Jinkela_buffer_3646 (
        .din(new_Jinkela_wire_4839),
        .dout(new_Jinkela_wire_4840)
    );

    bfr new_Jinkela_buffer_17297 (
        .din(new_Jinkela_wire_20641),
        .dout(new_Jinkela_wire_20642)
    );

    bfr new_Jinkela_buffer_3505 (
        .din(new_Jinkela_wire_4642),
        .dout(new_Jinkela_wire_4643)
    );

    bfr new_Jinkela_buffer_17268 (
        .din(new_Jinkela_wire_20610),
        .dout(new_Jinkela_wire_20611)
    );

    bfr new_Jinkela_buffer_3557 (
        .din(new_Jinkela_wire_4738),
        .dout(new_Jinkela_wire_4739)
    );

    bfr new_Jinkela_buffer_17456 (
        .din(_0773_),
        .dout(new_Jinkela_wire_20811)
    );

    bfr new_Jinkela_buffer_3506 (
        .din(new_Jinkela_wire_4643),
        .dout(new_Jinkela_wire_4644)
    );

    bfr new_Jinkela_buffer_17269 (
        .din(new_Jinkela_wire_20611),
        .dout(new_Jinkela_wire_20612)
    );

    bfr new_Jinkela_buffer_17298 (
        .din(new_Jinkela_wire_20642),
        .dout(new_Jinkela_wire_20643)
    );

    bfr new_Jinkela_buffer_3507 (
        .din(new_Jinkela_wire_4644),
        .dout(new_Jinkela_wire_4645)
    );

    bfr new_Jinkela_buffer_17270 (
        .din(new_Jinkela_wire_20612),
        .dout(new_Jinkela_wire_20613)
    );

    bfr new_Jinkela_buffer_3558 (
        .din(new_Jinkela_wire_4739),
        .dout(new_Jinkela_wire_4740)
    );

    bfr new_Jinkela_buffer_17333 (
        .din(new_Jinkela_wire_20681),
        .dout(new_Jinkela_wire_20682)
    );

    bfr new_Jinkela_buffer_17315 (
        .din(new_Jinkela_wire_20661),
        .dout(new_Jinkela_wire_20662)
    );

    bfr new_Jinkela_buffer_3508 (
        .din(new_Jinkela_wire_4645),
        .dout(new_Jinkela_wire_4646)
    );

    bfr new_Jinkela_buffer_17271 (
        .din(new_Jinkela_wire_20613),
        .dout(new_Jinkela_wire_20614)
    );

    bfr new_Jinkela_buffer_3647 (
        .din(new_Jinkela_wire_4840),
        .dout(new_Jinkela_wire_4841)
    );

    bfr new_Jinkela_buffer_17299 (
        .din(new_Jinkela_wire_20643),
        .dout(new_Jinkela_wire_20644)
    );

    bfr new_Jinkela_buffer_3509 (
        .din(new_Jinkela_wire_4646),
        .dout(new_Jinkela_wire_4647)
    );

    bfr new_Jinkela_buffer_17272 (
        .din(new_Jinkela_wire_20614),
        .dout(new_Jinkela_wire_20615)
    );

    bfr new_Jinkela_buffer_3559 (
        .din(new_Jinkela_wire_4740),
        .dout(new_Jinkela_wire_4741)
    );

    bfr new_Jinkela_buffer_3510 (
        .din(new_Jinkela_wire_4647),
        .dout(new_Jinkela_wire_4648)
    );

    bfr new_Jinkela_buffer_17273 (
        .din(new_Jinkela_wire_20615),
        .dout(new_Jinkela_wire_20616)
    );

    bfr new_Jinkela_buffer_17300 (
        .din(new_Jinkela_wire_20644),
        .dout(new_Jinkela_wire_20645)
    );

    spl2 new_Jinkela_splitter_449 (
        .a(_1460_),
        .b(new_Jinkela_wire_4901),
        .c(new_Jinkela_wire_4902)
    );

    bfr new_Jinkela_buffer_3511 (
        .din(new_Jinkela_wire_4648),
        .dout(new_Jinkela_wire_4649)
    );

    bfr new_Jinkela_buffer_17274 (
        .din(new_Jinkela_wire_20616),
        .dout(new_Jinkela_wire_20617)
    );

    bfr new_Jinkela_buffer_3560 (
        .din(new_Jinkela_wire_4741),
        .dout(new_Jinkela_wire_4742)
    );

    bfr new_Jinkela_buffer_17336 (
        .din(new_Jinkela_wire_20684),
        .dout(new_Jinkela_wire_20685)
    );

    bfr new_Jinkela_buffer_17316 (
        .din(new_Jinkela_wire_20662),
        .dout(new_Jinkela_wire_20663)
    );

    bfr new_Jinkela_buffer_3512 (
        .din(new_Jinkela_wire_4649),
        .dout(new_Jinkela_wire_4650)
    );

    bfr new_Jinkela_buffer_17275 (
        .din(new_Jinkela_wire_20617),
        .dout(new_Jinkela_wire_20618)
    );

    bfr new_Jinkela_buffer_3648 (
        .din(new_Jinkela_wire_4841),
        .dout(new_Jinkela_wire_4842)
    );

    bfr new_Jinkela_buffer_17301 (
        .din(new_Jinkela_wire_20645),
        .dout(new_Jinkela_wire_20646)
    );

    bfr new_Jinkela_buffer_3513 (
        .din(new_Jinkela_wire_4650),
        .dout(new_Jinkela_wire_4651)
    );

    bfr new_Jinkela_buffer_17276 (
        .din(new_Jinkela_wire_20618),
        .dout(new_Jinkela_wire_20619)
    );

    bfr new_Jinkela_buffer_3561 (
        .din(new_Jinkela_wire_4742),
        .dout(new_Jinkela_wire_4743)
    );

    bfr new_Jinkela_buffer_3514 (
        .din(new_Jinkela_wire_4651),
        .dout(new_Jinkela_wire_4652)
    );

    bfr new_Jinkela_buffer_17277 (
        .din(new_Jinkela_wire_20619),
        .dout(new_Jinkela_wire_20620)
    );

    bfr new_Jinkela_buffer_17302 (
        .din(new_Jinkela_wire_20646),
        .dout(new_Jinkela_wire_20647)
    );

    spl2 new_Jinkela_splitter_450 (
        .a(_1744_),
        .b(new_Jinkela_wire_4903),
        .c(new_Jinkela_wire_4904)
    );

    bfr new_Jinkela_buffer_3515 (
        .din(new_Jinkela_wire_4652),
        .dout(new_Jinkela_wire_4653)
    );

    bfr new_Jinkela_buffer_17278 (
        .din(new_Jinkela_wire_20620),
        .dout(new_Jinkela_wire_20621)
    );

    bfr new_Jinkela_buffer_3562 (
        .din(new_Jinkela_wire_4743),
        .dout(new_Jinkela_wire_4744)
    );

    bfr new_Jinkela_buffer_17445 (
        .din(new_Jinkela_wire_20795),
        .dout(new_Jinkela_wire_20796)
    );

    bfr new_Jinkela_buffer_17317 (
        .din(new_Jinkela_wire_20663),
        .dout(new_Jinkela_wire_20664)
    );

    bfr new_Jinkela_buffer_3516 (
        .din(new_Jinkela_wire_4653),
        .dout(new_Jinkela_wire_4654)
    );

    bfr new_Jinkela_buffer_17279 (
        .din(new_Jinkela_wire_20621),
        .dout(new_Jinkela_wire_20622)
    );

    bfr new_Jinkela_buffer_3649 (
        .din(new_Jinkela_wire_4842),
        .dout(new_Jinkela_wire_4843)
    );

    bfr new_Jinkela_buffer_17303 (
        .din(new_Jinkela_wire_20647),
        .dout(new_Jinkela_wire_20648)
    );

    bfr new_Jinkela_buffer_3517 (
        .din(new_Jinkela_wire_4654),
        .dout(new_Jinkela_wire_4655)
    );

    bfr new_Jinkela_buffer_17280 (
        .din(new_Jinkela_wire_20622),
        .dout(new_Jinkela_wire_20623)
    );

    bfr new_Jinkela_buffer_3563 (
        .din(new_Jinkela_wire_4744),
        .dout(new_Jinkela_wire_4745)
    );

    bfr new_Jinkela_buffer_3518 (
        .din(new_Jinkela_wire_4655),
        .dout(new_Jinkela_wire_4656)
    );

    spl2 new_Jinkela_splitter_1520 (
        .a(new_Jinkela_wire_20623),
        .b(new_Jinkela_wire_20624),
        .c(new_Jinkela_wire_20625)
    );

    bfr new_Jinkela_buffer_17337 (
        .din(new_Jinkela_wire_20685),
        .dout(new_Jinkela_wire_20686)
    );

    spl2 new_Jinkela_splitter_451 (
        .a(_1599_),
        .b(new_Jinkela_wire_4905),
        .c(new_Jinkela_wire_4906)
    );

    bfr new_Jinkela_buffer_17318 (
        .din(new_Jinkela_wire_20664),
        .dout(new_Jinkela_wire_20665)
    );

    bfr new_Jinkela_buffer_3519 (
        .din(new_Jinkela_wire_4656),
        .dout(new_Jinkela_wire_4657)
    );

    bfr new_Jinkela_buffer_17304 (
        .din(new_Jinkela_wire_20648),
        .dout(new_Jinkela_wire_20649)
    );

    bfr new_Jinkela_buffer_3564 (
        .din(new_Jinkela_wire_4745),
        .dout(new_Jinkela_wire_4746)
    );

    bfr new_Jinkela_buffer_17305 (
        .din(new_Jinkela_wire_20649),
        .dout(new_Jinkela_wire_20650)
    );

    bfr new_Jinkela_buffer_3520 (
        .din(new_Jinkela_wire_4657),
        .dout(new_Jinkela_wire_4658)
    );

    bfr new_Jinkela_buffer_3650 (
        .din(new_Jinkela_wire_4843),
        .dout(new_Jinkela_wire_4844)
    );

    spl2 new_Jinkela_splitter_1521 (
        .a(new_Jinkela_wire_20650),
        .b(new_Jinkela_wire_20651),
        .c(new_Jinkela_wire_20652)
    );

    spl2 new_Jinkela_splitter_418 (
        .a(new_Jinkela_wire_4658),
        .b(new_Jinkela_wire_4659),
        .c(new_Jinkela_wire_4660)
    );

    spl2 new_Jinkela_splitter_454 (
        .a(_0492_),
        .b(new_Jinkela_wire_4911),
        .c(new_Jinkela_wire_4912)
    );

    spl2 new_Jinkela_splitter_452 (
        .a(_0532_),
        .b(new_Jinkela_wire_4907),
        .c(new_Jinkela_wire_4908)
    );

    bfr new_Jinkela_buffer_17319 (
        .din(new_Jinkela_wire_20665),
        .dout(new_Jinkela_wire_20666)
    );

    bfr new_Jinkela_buffer_3565 (
        .din(new_Jinkela_wire_4746),
        .dout(new_Jinkela_wire_4747)
    );

    bfr new_Jinkela_buffer_17338 (
        .din(new_Jinkela_wire_20686),
        .dout(new_Jinkela_wire_20687)
    );

    bfr new_Jinkela_buffer_17320 (
        .din(new_Jinkela_wire_20666),
        .dout(new_Jinkela_wire_20667)
    );

    bfr new_Jinkela_buffer_3566 (
        .din(new_Jinkela_wire_4747),
        .dout(new_Jinkela_wire_4748)
    );

    bfr new_Jinkela_buffer_3651 (
        .din(new_Jinkela_wire_4844),
        .dout(new_Jinkela_wire_4845)
    );

    bfr new_Jinkela_buffer_17446 (
        .din(new_Jinkela_wire_20796),
        .dout(new_Jinkela_wire_20797)
    );

    bfr new_Jinkela_buffer_17321 (
        .din(new_Jinkela_wire_20667),
        .dout(new_Jinkela_wire_20668)
    );

    bfr new_Jinkela_buffer_3567 (
        .din(new_Jinkela_wire_4748),
        .dout(new_Jinkela_wire_4749)
    );

    bfr new_Jinkela_buffer_17339 (
        .din(new_Jinkela_wire_20687),
        .dout(new_Jinkela_wire_20688)
    );

    spl2 new_Jinkela_splitter_453 (
        .a(_0041_),
        .b(new_Jinkela_wire_4909),
        .c(new_Jinkela_wire_4910)
    );

    bfr new_Jinkela_buffer_17322 (
        .din(new_Jinkela_wire_20668),
        .dout(new_Jinkela_wire_20669)
    );

    bfr new_Jinkela_buffer_3568 (
        .din(new_Jinkela_wire_4749),
        .dout(new_Jinkela_wire_4750)
    );

    bfr new_Jinkela_buffer_3652 (
        .din(new_Jinkela_wire_4845),
        .dout(new_Jinkela_wire_4846)
    );

    bfr new_Jinkela_buffer_17452 (
        .din(new_Jinkela_wire_20806),
        .dout(new_Jinkela_wire_20807)
    );

    bfr new_Jinkela_buffer_17323 (
        .din(new_Jinkela_wire_20669),
        .dout(new_Jinkela_wire_20670)
    );

    bfr new_Jinkela_buffer_13938 (
        .din(new_Jinkela_wire_16621),
        .dout(new_Jinkela_wire_16622)
    );

    bfr new_Jinkela_buffer_13894 (
        .din(new_Jinkela_wire_16575),
        .dout(new_Jinkela_wire_16576)
    );

    spl2 new_Jinkela_splitter_1198 (
        .a(_0801_),
        .b(new_Jinkela_wire_16790),
        .c(new_Jinkela_wire_16791)
    );

    bfr new_Jinkela_buffer_13895 (
        .din(new_Jinkela_wire_16576),
        .dout(new_Jinkela_wire_16577)
    );

    bfr new_Jinkela_buffer_14021 (
        .din(new_Jinkela_wire_16708),
        .dout(new_Jinkela_wire_16709)
    );

    bfr new_Jinkela_buffer_13939 (
        .din(new_Jinkela_wire_16622),
        .dout(new_Jinkela_wire_16623)
    );

    bfr new_Jinkela_buffer_13896 (
        .din(new_Jinkela_wire_16577),
        .dout(new_Jinkela_wire_16578)
    );

    bfr new_Jinkela_buffer_13897 (
        .din(new_Jinkela_wire_16578),
        .dout(new_Jinkela_wire_16579)
    );

    spl2 new_Jinkela_splitter_1199 (
        .a(_0986_),
        .b(new_Jinkela_wire_16796),
        .c(new_Jinkela_wire_16797)
    );

    bfr new_Jinkela_buffer_13940 (
        .din(new_Jinkela_wire_16623),
        .dout(new_Jinkela_wire_16624)
    );

    bfr new_Jinkela_buffer_13898 (
        .din(new_Jinkela_wire_16579),
        .dout(new_Jinkela_wire_16580)
    );

    bfr new_Jinkela_buffer_14092 (
        .din(new_Jinkela_wire_16791),
        .dout(new_Jinkela_wire_16792)
    );

    bfr new_Jinkela_buffer_13899 (
        .din(new_Jinkela_wire_16580),
        .dout(new_Jinkela_wire_16581)
    );

    bfr new_Jinkela_buffer_14022 (
        .din(new_Jinkela_wire_16709),
        .dout(new_Jinkela_wire_16710)
    );

    bfr new_Jinkela_buffer_13941 (
        .din(new_Jinkela_wire_16624),
        .dout(new_Jinkela_wire_16625)
    );

    bfr new_Jinkela_buffer_13900 (
        .din(new_Jinkela_wire_16581),
        .dout(new_Jinkela_wire_16582)
    );

    bfr new_Jinkela_buffer_13901 (
        .din(new_Jinkela_wire_16582),
        .dout(new_Jinkela_wire_16583)
    );

    bfr new_Jinkela_buffer_14088 (
        .din(new_Jinkela_wire_16785),
        .dout(new_Jinkela_wire_16786)
    );

    bfr new_Jinkela_buffer_13942 (
        .din(new_Jinkela_wire_16625),
        .dout(new_Jinkela_wire_16626)
    );

    bfr new_Jinkela_buffer_13902 (
        .din(new_Jinkela_wire_16583),
        .dout(new_Jinkela_wire_16584)
    );

    bfr new_Jinkela_buffer_13903 (
        .din(new_Jinkela_wire_16584),
        .dout(new_Jinkela_wire_16585)
    );

    bfr new_Jinkela_buffer_14023 (
        .din(new_Jinkela_wire_16710),
        .dout(new_Jinkela_wire_16711)
    );

    bfr new_Jinkela_buffer_13943 (
        .din(new_Jinkela_wire_16626),
        .dout(new_Jinkela_wire_16627)
    );

    bfr new_Jinkela_buffer_13904 (
        .din(new_Jinkela_wire_16585),
        .dout(new_Jinkela_wire_16586)
    );

    bfr new_Jinkela_buffer_13905 (
        .din(new_Jinkela_wire_16586),
        .dout(new_Jinkela_wire_16587)
    );

    bfr new_Jinkela_buffer_13944 (
        .din(new_Jinkela_wire_16627),
        .dout(new_Jinkela_wire_16628)
    );

    bfr new_Jinkela_buffer_13906 (
        .din(new_Jinkela_wire_16587),
        .dout(new_Jinkela_wire_16588)
    );

    bfr new_Jinkela_buffer_13907 (
        .din(new_Jinkela_wire_16588),
        .dout(new_Jinkela_wire_16589)
    );

    bfr new_Jinkela_buffer_14024 (
        .din(new_Jinkela_wire_16711),
        .dout(new_Jinkela_wire_16712)
    );

    bfr new_Jinkela_buffer_13945 (
        .din(new_Jinkela_wire_16628),
        .dout(new_Jinkela_wire_16629)
    );

    bfr new_Jinkela_buffer_13908 (
        .din(new_Jinkela_wire_16589),
        .dout(new_Jinkela_wire_16590)
    );

    bfr new_Jinkela_buffer_13909 (
        .din(new_Jinkela_wire_16590),
        .dout(new_Jinkela_wire_16591)
    );

    bfr new_Jinkela_buffer_14089 (
        .din(new_Jinkela_wire_16786),
        .dout(new_Jinkela_wire_16787)
    );

    bfr new_Jinkela_buffer_13946 (
        .din(new_Jinkela_wire_16629),
        .dout(new_Jinkela_wire_16630)
    );

    bfr new_Jinkela_buffer_13910 (
        .din(new_Jinkela_wire_16591),
        .dout(new_Jinkela_wire_16592)
    );

    bfr new_Jinkela_buffer_13911 (
        .din(new_Jinkela_wire_16592),
        .dout(new_Jinkela_wire_16593)
    );

    bfr new_Jinkela_buffer_14025 (
        .din(new_Jinkela_wire_16712),
        .dout(new_Jinkela_wire_16713)
    );

    bfr new_Jinkela_buffer_13947 (
        .din(new_Jinkela_wire_16630),
        .dout(new_Jinkela_wire_16631)
    );

    bfr new_Jinkela_buffer_13912 (
        .din(new_Jinkela_wire_16593),
        .dout(new_Jinkela_wire_16594)
    );

    bfr new_Jinkela_buffer_13913 (
        .din(new_Jinkela_wire_16594),
        .dout(new_Jinkela_wire_16595)
    );

    bfr new_Jinkela_buffer_13948 (
        .din(new_Jinkela_wire_16631),
        .dout(new_Jinkela_wire_16632)
    );

    bfr new_Jinkela_buffer_13914 (
        .din(new_Jinkela_wire_16595),
        .dout(new_Jinkela_wire_16596)
    );

    bfr new_Jinkela_buffer_6929 (
        .din(new_Jinkela_wire_8672),
        .dout(new_Jinkela_wire_8673)
    );

    bfr new_Jinkela_buffer_6977 (
        .din(new_Jinkela_wire_8730),
        .dout(new_Jinkela_wire_8731)
    );

    bfr new_Jinkela_buffer_6930 (
        .din(new_Jinkela_wire_8673),
        .dout(new_Jinkela_wire_8674)
    );

    bfr new_Jinkela_buffer_7021 (
        .din(new_Jinkela_wire_8782),
        .dout(new_Jinkela_wire_8783)
    );

    bfr new_Jinkela_buffer_6931 (
        .din(new_Jinkela_wire_8674),
        .dout(new_Jinkela_wire_8675)
    );

    bfr new_Jinkela_buffer_6978 (
        .din(new_Jinkela_wire_8731),
        .dout(new_Jinkela_wire_8732)
    );

    bfr new_Jinkela_buffer_6932 (
        .din(new_Jinkela_wire_8675),
        .dout(new_Jinkela_wire_8676)
    );

    bfr new_Jinkela_buffer_7082 (
        .din(new_Jinkela_wire_8857),
        .dout(new_Jinkela_wire_8858)
    );

    bfr new_Jinkela_buffer_6933 (
        .din(new_Jinkela_wire_8676),
        .dout(new_Jinkela_wire_8677)
    );

    bfr new_Jinkela_buffer_6979 (
        .din(new_Jinkela_wire_8732),
        .dout(new_Jinkela_wire_8733)
    );

    bfr new_Jinkela_buffer_6934 (
        .din(new_Jinkela_wire_8677),
        .dout(new_Jinkela_wire_8678)
    );

    bfr new_Jinkela_buffer_7022 (
        .din(new_Jinkela_wire_8783),
        .dout(new_Jinkela_wire_8784)
    );

    bfr new_Jinkela_buffer_6935 (
        .din(new_Jinkela_wire_8678),
        .dout(new_Jinkela_wire_8679)
    );

    bfr new_Jinkela_buffer_6980 (
        .din(new_Jinkela_wire_8733),
        .dout(new_Jinkela_wire_8734)
    );

    spl2 new_Jinkela_splitter_721 (
        .a(new_Jinkela_wire_8679),
        .b(new_Jinkela_wire_8680),
        .c(new_Jinkela_wire_8681)
    );

    bfr new_Jinkela_buffer_6981 (
        .din(new_Jinkela_wire_8734),
        .dout(new_Jinkela_wire_8735)
    );

    bfr new_Jinkela_buffer_7089 (
        .din(new_Jinkela_wire_8868),
        .dout(new_Jinkela_wire_8869)
    );

    bfr new_Jinkela_buffer_7023 (
        .din(new_Jinkela_wire_8784),
        .dout(new_Jinkela_wire_8785)
    );

    bfr new_Jinkela_buffer_6982 (
        .din(new_Jinkela_wire_8735),
        .dout(new_Jinkela_wire_8736)
    );

    bfr new_Jinkela_buffer_7083 (
        .din(new_Jinkela_wire_8858),
        .dout(new_Jinkela_wire_8859)
    );

    bfr new_Jinkela_buffer_6983 (
        .din(new_Jinkela_wire_8736),
        .dout(new_Jinkela_wire_8737)
    );

    bfr new_Jinkela_buffer_7024 (
        .din(new_Jinkela_wire_8785),
        .dout(new_Jinkela_wire_8786)
    );

    bfr new_Jinkela_buffer_6984 (
        .din(new_Jinkela_wire_8737),
        .dout(new_Jinkela_wire_8738)
    );

    bfr new_Jinkela_buffer_7181 (
        .din(_1537_),
        .dout(new_Jinkela_wire_8963)
    );

    bfr new_Jinkela_buffer_6985 (
        .din(new_Jinkela_wire_8738),
        .dout(new_Jinkela_wire_8739)
    );

    bfr new_Jinkela_buffer_7025 (
        .din(new_Jinkela_wire_8786),
        .dout(new_Jinkela_wire_8787)
    );

    bfr new_Jinkela_buffer_6986 (
        .din(new_Jinkela_wire_8739),
        .dout(new_Jinkela_wire_8740)
    );

    bfr new_Jinkela_buffer_7084 (
        .din(new_Jinkela_wire_8859),
        .dout(new_Jinkela_wire_8860)
    );

    bfr new_Jinkela_buffer_6987 (
        .din(new_Jinkela_wire_8740),
        .dout(new_Jinkela_wire_8741)
    );

    bfr new_Jinkela_buffer_7026 (
        .din(new_Jinkela_wire_8787),
        .dout(new_Jinkela_wire_8788)
    );

    bfr new_Jinkela_buffer_6988 (
        .din(new_Jinkela_wire_8741),
        .dout(new_Jinkela_wire_8742)
    );

    spl2 new_Jinkela_splitter_740 (
        .a(_0312_),
        .b(new_Jinkela_wire_8964),
        .c(new_Jinkela_wire_8965)
    );

    bfr new_Jinkela_buffer_6989 (
        .din(new_Jinkela_wire_8742),
        .dout(new_Jinkela_wire_8743)
    );

    bfr new_Jinkela_buffer_7027 (
        .din(new_Jinkela_wire_8788),
        .dout(new_Jinkela_wire_8789)
    );

    bfr new_Jinkela_buffer_6990 (
        .din(new_Jinkela_wire_8743),
        .dout(new_Jinkela_wire_8744)
    );

    bfr new_Jinkela_buffer_7085 (
        .din(new_Jinkela_wire_8860),
        .dout(new_Jinkela_wire_8861)
    );

    bfr new_Jinkela_buffer_6991 (
        .din(new_Jinkela_wire_8744),
        .dout(new_Jinkela_wire_8745)
    );

    bfr new_Jinkela_buffer_7028 (
        .din(new_Jinkela_wire_8789),
        .dout(new_Jinkela_wire_8790)
    );

    bfr new_Jinkela_buffer_6992 (
        .din(new_Jinkela_wire_8745),
        .dout(new_Jinkela_wire_8746)
    );

    bfr new_Jinkela_buffer_7090 (
        .din(new_Jinkela_wire_8869),
        .dout(new_Jinkela_wire_8870)
    );

    bfr new_Jinkela_buffer_6993 (
        .din(new_Jinkela_wire_8746),
        .dout(new_Jinkela_wire_8747)
    );

    bfr new_Jinkela_buffer_7029 (
        .din(new_Jinkela_wire_8790),
        .dout(new_Jinkela_wire_8791)
    );

    spl4L new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_265),
        .c(new_Jinkela_wire_266),
        .d(new_Jinkela_wire_267),
        .b(new_Jinkela_wire_268),
        .e(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    spl4L new_Jinkela_splitter_72 (
        .a(new_Jinkela_wire_275),
        .c(new_Jinkela_wire_276),
        .d(new_Jinkela_wire_277),
        .b(new_Jinkela_wire_278),
        .e(new_Jinkela_wire_279)
    );

    spl3L new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_288),
        .d(new_Jinkela_wire_289),
        .b(new_Jinkela_wire_290),
        .c(new_Jinkela_wire_291)
    );

    spl4L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_280),
        .c(new_Jinkela_wire_281),
        .d(new_Jinkela_wire_282),
        .b(new_Jinkela_wire_283),
        .e(new_Jinkela_wire_284)
    );

    spl4L new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_311),
        .c(new_Jinkela_wire_312),
        .d(new_Jinkela_wire_314),
        .b(new_Jinkela_wire_319),
        .e(new_Jinkela_wire_324)
    );

    spl3L new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_307),
        .d(new_Jinkela_wire_308),
        .b(new_Jinkela_wire_309),
        .c(new_Jinkela_wire_310)
    );

    spl4L new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_292),
        .c(new_Jinkela_wire_293),
        .d(new_Jinkela_wire_294),
        .b(new_Jinkela_wire_295),
        .e(new_Jinkela_wire_296)
    );

    spl4L new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_357),
        .c(new_Jinkela_wire_358),
        .d(new_Jinkela_wire_359),
        .b(new_Jinkela_wire_360),
        .e(new_Jinkela_wire_361)
    );

    spl4L new_Jinkela_splitter_78 (
        .a(new_Jinkela_wire_297),
        .c(new_Jinkela_wire_298),
        .d(new_Jinkela_wire_299),
        .b(new_Jinkela_wire_300),
        .e(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    spl4L new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_319),
        .c(new_Jinkela_wire_320),
        .d(new_Jinkela_wire_321),
        .b(new_Jinkela_wire_322),
        .e(new_Jinkela_wire_323)
    );

    spl4L new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_302),
        .c(new_Jinkela_wire_303),
        .d(new_Jinkela_wire_304),
        .b(new_Jinkela_wire_305),
        .e(new_Jinkela_wire_306)
    );

    spl4L new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_331),
        .c(new_Jinkela_wire_332),
        .d(new_Jinkela_wire_336),
        .b(new_Jinkela_wire_341),
        .e(new_Jinkela_wire_346)
    );

    spl4L new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_336),
        .c(new_Jinkela_wire_337),
        .d(new_Jinkela_wire_338),
        .b(new_Jinkela_wire_339),
        .e(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_329),
        .dout(new_Jinkela_wire_330)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(N1),
        .b(new_Jinkela_wire_329),
        .c(new_Jinkela_wire_331)
    );

    spl4L new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_314),
        .c(new_Jinkela_wire_315),
        .d(new_Jinkela_wire_316),
        .b(new_Jinkela_wire_317),
        .e(new_Jinkela_wire_318)
    );

    spl4L new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_324),
        .c(new_Jinkela_wire_325),
        .d(new_Jinkela_wire_326),
        .b(new_Jinkela_wire_327),
        .e(new_Jinkela_wire_328)
    );

    spl4L new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_351),
        .c(new_Jinkela_wire_352),
        .d(new_Jinkela_wire_357),
        .b(new_Jinkela_wire_362),
        .e(new_Jinkela_wire_367)
    );

    spl3L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_332),
        .d(new_Jinkela_wire_333),
        .b(new_Jinkela_wire_334),
        .c(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_18 (
        .din(N103),
        .dout(new_Jinkela_wire_351)
    );

    spl4L new_Jinkela_splitter_90 (
        .a(new_Jinkela_wire_341),
        .c(new_Jinkela_wire_342),
        .d(new_Jinkela_wire_343),
        .b(new_Jinkela_wire_344),
        .e(new_Jinkela_wire_345)
    );

    spl4L new_Jinkela_splitter_91 (
        .a(new_Jinkela_wire_346),
        .c(new_Jinkela_wire_347),
        .d(new_Jinkela_wire_348),
        .b(new_Jinkela_wire_349),
        .e(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_19 (
        .din(N188),
        .dout(new_Jinkela_wire_372)
    );

    spl4L new_Jinkela_splitter_100 (
        .a(new_Jinkela_wire_383),
        .c(new_Jinkela_wire_384),
        .d(new_Jinkela_wire_385),
        .b(new_Jinkela_wire_386),
        .e(new_Jinkela_wire_387)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(N409),
        .b(new_Jinkela_wire_443),
        .c(new_Jinkela_wire_445)
    );

    spl4L new_Jinkela_splitter_93 (
        .a(new_Jinkela_wire_352),
        .c(new_Jinkela_wire_353),
        .d(new_Jinkela_wire_354),
        .b(new_Jinkela_wire_355),
        .e(new_Jinkela_wire_356)
    );

    spl4L new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_372),
        .c(new_Jinkela_wire_373),
        .d(new_Jinkela_wire_378),
        .b(new_Jinkela_wire_383),
        .e(new_Jinkela_wire_388)
    );

    spl4L new_Jinkela_splitter_95 (
        .a(new_Jinkela_wire_362),
        .c(new_Jinkela_wire_363),
        .d(new_Jinkela_wire_364),
        .b(new_Jinkela_wire_365),
        .e(new_Jinkela_wire_366)
    );

    spl4L new_Jinkela_splitter_96 (
        .a(new_Jinkela_wire_367),
        .c(new_Jinkela_wire_368),
        .d(new_Jinkela_wire_369),
        .b(new_Jinkela_wire_370),
        .e(new_Jinkela_wire_371)
    );

    bfr new_Jinkela_buffer_20 (
        .din(N205),
        .dout(new_Jinkela_wire_393)
    );

    spl4L new_Jinkela_splitter_105 (
        .a(new_Jinkela_wire_404),
        .c(new_Jinkela_wire_405),
        .d(new_Jinkela_wire_406),
        .b(new_Jinkela_wire_407),
        .e(new_Jinkela_wire_408)
    );

    spl4L new_Jinkela_splitter_98 (
        .a(new_Jinkela_wire_373),
        .c(new_Jinkela_wire_374),
        .d(new_Jinkela_wire_375),
        .b(new_Jinkela_wire_376),
        .e(new_Jinkela_wire_377)
    );

    spl4L new_Jinkela_splitter_99 (
        .a(new_Jinkela_wire_378),
        .c(new_Jinkela_wire_379),
        .d(new_Jinkela_wire_380),
        .b(new_Jinkela_wire_381),
        .e(new_Jinkela_wire_382)
    );

    spl4L new_Jinkela_splitter_102 (
        .a(new_Jinkela_wire_393),
        .c(new_Jinkela_wire_394),
        .d(new_Jinkela_wire_399),
        .b(new_Jinkela_wire_404),
        .e(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    spl4L new_Jinkela_splitter_101 (
        .a(new_Jinkela_wire_388),
        .c(new_Jinkela_wire_389),
        .d(new_Jinkela_wire_390),
        .b(new_Jinkela_wire_391),
        .e(new_Jinkela_wire_392)
    );

    spl4L new_Jinkela_splitter_108 (
        .a(new_Jinkela_wire_417),
        .c(new_Jinkela_wire_418),
        .d(new_Jinkela_wire_423),
        .b(new_Jinkela_wire_428),
        .e(new_Jinkela_wire_433)
    );

    spl4L new_Jinkela_splitter_103 (
        .a(new_Jinkela_wire_394),
        .c(new_Jinkela_wire_395),
        .d(new_Jinkela_wire_396),
        .b(new_Jinkela_wire_397),
        .e(new_Jinkela_wire_398)
    );

    spl4L new_Jinkela_splitter_104 (
        .a(new_Jinkela_wire_399),
        .c(new_Jinkela_wire_400),
        .d(new_Jinkela_wire_401),
        .b(new_Jinkela_wire_402),
        .e(new_Jinkela_wire_403)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(N256),
        .b(new_Jinkela_wire_414),
        .c(new_Jinkela_wire_417)
    );

    bfr new_Jinkela_buffer_17544 (
        .din(_0717_),
        .dout(new_Jinkela_wire_20901)
    );

    bfr new_Jinkela_buffer_17340 (
        .din(new_Jinkela_wire_20688),
        .dout(new_Jinkela_wire_20689)
    );

    bfr new_Jinkela_buffer_17324 (
        .din(new_Jinkela_wire_20670),
        .dout(new_Jinkela_wire_20671)
    );

    bfr new_Jinkela_buffer_17447 (
        .din(new_Jinkela_wire_20797),
        .dout(new_Jinkela_wire_20798)
    );

    bfr new_Jinkela_buffer_17325 (
        .din(new_Jinkela_wire_20671),
        .dout(new_Jinkela_wire_20672)
    );

    bfr new_Jinkela_buffer_17341 (
        .din(new_Jinkela_wire_20689),
        .dout(new_Jinkela_wire_20690)
    );

    bfr new_Jinkela_buffer_17326 (
        .din(new_Jinkela_wire_20672),
        .dout(new_Jinkela_wire_20673)
    );

    bfr new_Jinkela_buffer_17327 (
        .din(new_Jinkela_wire_20673),
        .dout(new_Jinkela_wire_20674)
    );

    bfr new_Jinkela_buffer_17545 (
        .din(_1342_),
        .dout(new_Jinkela_wire_20902)
    );

    bfr new_Jinkela_buffer_17342 (
        .din(new_Jinkela_wire_20690),
        .dout(new_Jinkela_wire_20691)
    );

    bfr new_Jinkela_buffer_17328 (
        .din(new_Jinkela_wire_20674),
        .dout(new_Jinkela_wire_20675)
    );

    bfr new_Jinkela_buffer_17448 (
        .din(new_Jinkela_wire_20798),
        .dout(new_Jinkela_wire_20799)
    );

    bfr new_Jinkela_buffer_17329 (
        .din(new_Jinkela_wire_20675),
        .dout(new_Jinkela_wire_20676)
    );

    bfr new_Jinkela_buffer_17343 (
        .din(new_Jinkela_wire_20691),
        .dout(new_Jinkela_wire_20692)
    );

    bfr new_Jinkela_buffer_17453 (
        .din(new_Jinkela_wire_20807),
        .dout(new_Jinkela_wire_20808)
    );

    bfr new_Jinkela_buffer_17344 (
        .din(new_Jinkela_wire_20692),
        .dout(new_Jinkela_wire_20693)
    );

    bfr new_Jinkela_buffer_17449 (
        .din(new_Jinkela_wire_20799),
        .dout(new_Jinkela_wire_20800)
    );

    bfr new_Jinkela_buffer_17345 (
        .din(new_Jinkela_wire_20693),
        .dout(new_Jinkela_wire_20694)
    );

    bfr new_Jinkela_buffer_17457 (
        .din(new_Jinkela_wire_20811),
        .dout(new_Jinkela_wire_20812)
    );

    bfr new_Jinkela_buffer_17346 (
        .din(new_Jinkela_wire_20694),
        .dout(new_Jinkela_wire_20695)
    );

    bfr new_Jinkela_buffer_17450 (
        .din(new_Jinkela_wire_20800),
        .dout(new_Jinkela_wire_20801)
    );

    bfr new_Jinkela_buffer_17347 (
        .din(new_Jinkela_wire_20695),
        .dout(new_Jinkela_wire_20696)
    );

    bfr new_Jinkela_buffer_17454 (
        .din(new_Jinkela_wire_20808),
        .dout(new_Jinkela_wire_20809)
    );

    bfr new_Jinkela_buffer_17348 (
        .din(new_Jinkela_wire_20696),
        .dout(new_Jinkela_wire_20697)
    );

    bfr new_Jinkela_buffer_17451 (
        .din(new_Jinkela_wire_20801),
        .dout(new_Jinkela_wire_20802)
    );

    bfr new_Jinkela_buffer_17349 (
        .din(new_Jinkela_wire_20697),
        .dout(new_Jinkela_wire_20698)
    );

    spl2 new_Jinkela_splitter_1527 (
        .a(_1558_),
        .b(new_Jinkela_wire_20903),
        .c(new_Jinkela_wire_20904)
    );

    bfr new_Jinkela_buffer_17350 (
        .din(new_Jinkela_wire_20698),
        .dout(new_Jinkela_wire_20699)
    );

    spl2 new_Jinkela_splitter_1524 (
        .a(new_Jinkela_wire_20802),
        .b(new_Jinkela_wire_20803),
        .c(new_Jinkela_wire_20804)
    );

    bfr new_Jinkela_buffer_17351 (
        .din(new_Jinkela_wire_20699),
        .dout(new_Jinkela_wire_20700)
    );

    bfr new_Jinkela_buffer_17458 (
        .din(new_Jinkela_wire_20812),
        .dout(new_Jinkela_wire_20813)
    );

    bfr new_Jinkela_buffer_17352 (
        .din(new_Jinkela_wire_20700),
        .dout(new_Jinkela_wire_20701)
    );

    bfr new_Jinkela_buffer_17455 (
        .din(new_Jinkela_wire_20809),
        .dout(new_Jinkela_wire_20810)
    );

    bfr new_Jinkela_buffer_17353 (
        .din(new_Jinkela_wire_20701),
        .dout(new_Jinkela_wire_20702)
    );

    spl2 new_Jinkela_splitter_1528 (
        .a(_0427_),
        .b(new_Jinkela_wire_20905),
        .c(new_Jinkela_wire_20906)
    );

    bfr new_Jinkela_buffer_17354 (
        .din(new_Jinkela_wire_20702),
        .dout(new_Jinkela_wire_20703)
    );

    bfr new_Jinkela_buffer_17459 (
        .din(new_Jinkela_wire_20813),
        .dout(new_Jinkela_wire_20814)
    );

    bfr new_Jinkela_buffer_17355 (
        .din(new_Jinkela_wire_20703),
        .dout(new_Jinkela_wire_20704)
    );

    bfr new_Jinkela_buffer_17546 (
        .din(_0019_),
        .dout(new_Jinkela_wire_20907)
    );

    bfr new_Jinkela_buffer_17356 (
        .din(new_Jinkela_wire_20704),
        .dout(new_Jinkela_wire_20705)
    );

    bfr new_Jinkela_buffer_17460 (
        .din(new_Jinkela_wire_20814),
        .dout(new_Jinkela_wire_20815)
    );

    bfr new_Jinkela_buffer_17357 (
        .din(new_Jinkela_wire_20705),
        .dout(new_Jinkela_wire_20706)
    );

    spl2 new_Jinkela_splitter_1200 (
        .a(_1021_),
        .b(new_Jinkela_wire_16798),
        .c(new_Jinkela_wire_16799)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_443),
        .dout(new_Jinkela_wire_444)
    );

    bfr new_Jinkela_buffer_13915 (
        .din(new_Jinkela_wire_16596),
        .dout(new_Jinkela_wire_16597)
    );

    spl4L new_Jinkela_splitter_106 (
        .a(new_Jinkela_wire_409),
        .c(new_Jinkela_wire_410),
        .d(new_Jinkela_wire_411),
        .b(new_Jinkela_wire_412),
        .e(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_14026 (
        .din(new_Jinkela_wire_16713),
        .dout(new_Jinkela_wire_16714)
    );

    bfr new_Jinkela_buffer_13949 (
        .din(new_Jinkela_wire_16632),
        .dout(new_Jinkela_wire_16633)
    );

    spl4L new_Jinkela_splitter_114 (
        .a(new_Jinkela_wire_445),
        .c(new_Jinkela_wire_446),
        .d(new_Jinkela_wire_450),
        .b(new_Jinkela_wire_455),
        .e(new_Jinkela_wire_460)
    );

    bfr new_Jinkela_buffer_13916 (
        .din(new_Jinkela_wire_16597),
        .dout(new_Jinkela_wire_16598)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    spl4L new_Jinkela_splitter_121 (
        .a(new_Jinkela_wire_471),
        .c(new_Jinkela_wire_472),
        .d(new_Jinkela_wire_473),
        .b(new_Jinkela_wire_474),
        .e(new_Jinkela_wire_475)
    );

    spl4L new_Jinkela_splitter_110 (
        .a(new_Jinkela_wire_423),
        .c(new_Jinkela_wire_424),
        .d(new_Jinkela_wire_425),
        .b(new_Jinkela_wire_426),
        .e(new_Jinkela_wire_427)
    );

    spl2 new_Jinkela_splitter_1190 (
        .a(new_Jinkela_wire_16598),
        .b(new_Jinkela_wire_16599),
        .c(new_Jinkela_wire_16600)
    );

    spl4L new_Jinkela_splitter_109 (
        .a(new_Jinkela_wire_418),
        .c(new_Jinkela_wire_419),
        .d(new_Jinkela_wire_420),
        .b(new_Jinkela_wire_421),
        .e(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_14090 (
        .din(new_Jinkela_wire_16787),
        .dout(new_Jinkela_wire_16788)
    );

    bfr new_Jinkela_buffer_13950 (
        .din(new_Jinkela_wire_16633),
        .dout(new_Jinkela_wire_16634)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_437),
        .dout(new_Jinkela_wire_438)
    );

    bfr new_Jinkela_buffer_14027 (
        .din(new_Jinkela_wire_16714),
        .dout(new_Jinkela_wire_16715)
    );

    bfr new_Jinkela_buffer_13951 (
        .din(new_Jinkela_wire_16634),
        .dout(new_Jinkela_wire_16635)
    );

    spl4L new_Jinkela_splitter_111 (
        .a(new_Jinkela_wire_428),
        .c(new_Jinkela_wire_429),
        .d(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_431),
        .e(new_Jinkela_wire_432)
    );

    spl4L new_Jinkela_splitter_112 (
        .a(new_Jinkela_wire_433),
        .c(new_Jinkela_wire_434),
        .d(new_Jinkela_wire_435),
        .b(new_Jinkela_wire_436),
        .e(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_13952 (
        .din(new_Jinkela_wire_16635),
        .dout(new_Jinkela_wire_16636)
    );

    spl4L new_Jinkela_splitter_119 (
        .a(new_Jinkela_wire_465),
        .c(new_Jinkela_wire_466),
        .d(new_Jinkela_wire_471),
        .b(new_Jinkela_wire_476),
        .e(new_Jinkela_wire_481)
    );

    spl3L new_Jinkela_splitter_115 (
        .a(new_Jinkela_wire_446),
        .d(new_Jinkela_wire_447),
        .b(new_Jinkela_wire_448),
        .c(new_Jinkela_wire_449)
    );

    bfr new_Jinkela_buffer_14028 (
        .din(new_Jinkela_wire_16715),
        .dout(new_Jinkela_wire_16716)
    );

    bfr new_Jinkela_buffer_13953 (
        .din(new_Jinkela_wire_16636),
        .dout(new_Jinkela_wire_16637)
    );

    spl4L new_Jinkela_splitter_116 (
        .a(new_Jinkela_wire_450),
        .c(new_Jinkela_wire_451),
        .d(new_Jinkela_wire_452),
        .b(new_Jinkela_wire_453),
        .e(new_Jinkela_wire_454)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_438),
        .dout(new_Jinkela_wire_439)
    );

    bfr new_Jinkela_buffer_14093 (
        .din(new_Jinkela_wire_16792),
        .dout(new_Jinkela_wire_16793)
    );

    bfr new_Jinkela_buffer_13954 (
        .din(new_Jinkela_wire_16637),
        .dout(new_Jinkela_wire_16638)
    );

    bfr new_Jinkela_buffer_29 (
        .din(N86),
        .dout(new_Jinkela_wire_465)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    bfr new_Jinkela_buffer_14029 (
        .din(new_Jinkela_wire_16716),
        .dout(new_Jinkela_wire_16717)
    );

    bfr new_Jinkela_buffer_13955 (
        .din(new_Jinkela_wire_16638),
        .dout(new_Jinkela_wire_16639)
    );

    spl4L new_Jinkela_splitter_117 (
        .a(new_Jinkela_wire_455),
        .c(new_Jinkela_wire_456),
        .d(new_Jinkela_wire_457),
        .b(new_Jinkela_wire_458),
        .e(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    spl2 new_Jinkela_splitter_1203 (
        .a(_0832_),
        .b(new_Jinkela_wire_16868),
        .c(new_Jinkela_wire_16869)
    );

    bfr new_Jinkela_buffer_13956 (
        .din(new_Jinkela_wire_16639),
        .dout(new_Jinkela_wire_16640)
    );

    bfr new_Jinkela_buffer_14096 (
        .din(_1571_),
        .dout(new_Jinkela_wire_16800)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_441),
        .dout(new_Jinkela_wire_442)
    );

    bfr new_Jinkela_buffer_14030 (
        .din(new_Jinkela_wire_16717),
        .dout(new_Jinkela_wire_16718)
    );

    bfr new_Jinkela_buffer_13957 (
        .din(new_Jinkela_wire_16640),
        .dout(new_Jinkela_wire_16641)
    );

    spl4L new_Jinkela_splitter_118 (
        .a(new_Jinkela_wire_460),
        .c(new_Jinkela_wire_461),
        .d(new_Jinkela_wire_462),
        .b(new_Jinkela_wire_463),
        .e(new_Jinkela_wire_464)
    );

    bfr new_Jinkela_buffer_14094 (
        .din(new_Jinkela_wire_16793),
        .dout(new_Jinkela_wire_16794)
    );

    bfr new_Jinkela_buffer_13958 (
        .din(new_Jinkela_wire_16641),
        .dout(new_Jinkela_wire_16642)
    );

    bfr new_Jinkela_buffer_30 (
        .din(N137),
        .dout(new_Jinkela_wire_486)
    );

    spl4L new_Jinkela_splitter_127 (
        .a(new_Jinkela_wire_497),
        .c(new_Jinkela_wire_498),
        .d(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_500),
        .e(new_Jinkela_wire_501)
    );

    bfr new_Jinkela_buffer_14031 (
        .din(new_Jinkela_wire_16718),
        .dout(new_Jinkela_wire_16719)
    );

    bfr new_Jinkela_buffer_13959 (
        .din(new_Jinkela_wire_16642),
        .dout(new_Jinkela_wire_16643)
    );

    spl4L new_Jinkela_splitter_120 (
        .a(new_Jinkela_wire_466),
        .c(new_Jinkela_wire_467),
        .d(new_Jinkela_wire_468),
        .b(new_Jinkela_wire_469),
        .e(new_Jinkela_wire_470)
    );

    spl4L new_Jinkela_splitter_124 (
        .a(new_Jinkela_wire_486),
        .c(new_Jinkela_wire_487),
        .d(new_Jinkela_wire_492),
        .b(new_Jinkela_wire_497),
        .e(new_Jinkela_wire_502)
    );

    bfr new_Jinkela_buffer_13960 (
        .din(new_Jinkela_wire_16643),
        .dout(new_Jinkela_wire_16644)
    );

    spl4L new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_476),
        .c(new_Jinkela_wire_477),
        .d(new_Jinkela_wire_478),
        .b(new_Jinkela_wire_479),
        .e(new_Jinkela_wire_480)
    );

    spl4L new_Jinkela_splitter_123 (
        .a(new_Jinkela_wire_481),
        .c(new_Jinkela_wire_482),
        .d(new_Jinkela_wire_483),
        .b(new_Jinkela_wire_484),
        .e(new_Jinkela_wire_485)
    );

    spl2 new_Jinkela_splitter_1202 (
        .a(_0034_),
        .b(new_Jinkela_wire_16866),
        .c(new_Jinkela_wire_16867)
    );

    bfr new_Jinkela_buffer_14032 (
        .din(new_Jinkela_wire_16719),
        .dout(new_Jinkela_wire_16720)
    );

    spl2 new_Jinkela_splitter_129 (
        .a(N511),
        .b(new_Jinkela_wire_507),
        .c(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_13961 (
        .din(new_Jinkela_wire_16644),
        .dout(new_Jinkela_wire_16645)
    );

    bfr new_Jinkela_buffer_33 (
        .din(N35),
        .dout(new_Jinkela_wire_551)
    );

    spl4L new_Jinkela_splitter_125 (
        .a(new_Jinkela_wire_487),
        .c(new_Jinkela_wire_488),
        .d(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_490),
        .e(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_14095 (
        .din(new_Jinkela_wire_16794),
        .dout(new_Jinkela_wire_16795)
    );

    spl4L new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_492),
        .c(new_Jinkela_wire_493),
        .d(new_Jinkela_wire_494),
        .b(new_Jinkela_wire_495),
        .e(new_Jinkela_wire_496)
    );

    bfr new_Jinkela_buffer_13962 (
        .din(new_Jinkela_wire_16645),
        .dout(new_Jinkela_wire_16646)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    spl4L new_Jinkela_splitter_130 (
        .a(new_Jinkela_wire_509),
        .c(new_Jinkela_wire_510),
        .d(new_Jinkela_wire_514),
        .b(new_Jinkela_wire_519),
        .e(new_Jinkela_wire_524)
    );

    bfr new_Jinkela_buffer_14033 (
        .din(new_Jinkela_wire_16720),
        .dout(new_Jinkela_wire_16721)
    );

    bfr new_Jinkela_buffer_13963 (
        .din(new_Jinkela_wire_16646),
        .dout(new_Jinkela_wire_16647)
    );

    spl4L new_Jinkela_splitter_128 (
        .a(new_Jinkela_wire_502),
        .c(new_Jinkela_wire_503),
        .d(new_Jinkela_wire_504),
        .b(new_Jinkela_wire_505),
        .e(new_Jinkela_wire_506)
    );

    bfr new_Jinkela_buffer_14097 (
        .din(new_Jinkela_wire_16800),
        .dout(new_Jinkela_wire_16801)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    bfr new_Jinkela_buffer_13964 (
        .din(new_Jinkela_wire_16647),
        .dout(new_Jinkela_wire_16648)
    );

    spl3L new_Jinkela_splitter_131 (
        .a(new_Jinkela_wire_510),
        .d(new_Jinkela_wire_511),
        .b(new_Jinkela_wire_512),
        .c(new_Jinkela_wire_513)
    );

    bfr new_Jinkela_buffer_35 (
        .din(N239),
        .dout(new_Jinkela_wire_594)
    );

    bfr new_Jinkela_buffer_14034 (
        .din(new_Jinkela_wire_16721),
        .dout(new_Jinkela_wire_16722)
    );

    spl4L new_Jinkela_splitter_132 (
        .a(new_Jinkela_wire_514),
        .c(new_Jinkela_wire_515),
        .d(new_Jinkela_wire_516),
        .b(new_Jinkela_wire_517),
        .e(new_Jinkela_wire_518)
    );

    bfr new_Jinkela_buffer_13965 (
        .din(new_Jinkela_wire_16648),
        .dout(new_Jinkela_wire_16649)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(N307),
        .b(new_Jinkela_wire_529),
        .c(new_Jinkela_wire_531)
    );

    spl2 new_Jinkela_splitter_1204 (
        .a(_0775_),
        .b(new_Jinkela_wire_16870),
        .c(new_Jinkela_wire_16871)
    );

    spl4L new_Jinkela_splitter_136 (
        .a(new_Jinkela_wire_531),
        .c(new_Jinkela_wire_532),
        .d(new_Jinkela_wire_536),
        .b(new_Jinkela_wire_541),
        .e(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_13966 (
        .din(new_Jinkela_wire_16649),
        .dout(new_Jinkela_wire_16650)
    );

    spl4L new_Jinkela_splitter_133 (
        .a(new_Jinkela_wire_519),
        .c(new_Jinkela_wire_520),
        .d(new_Jinkela_wire_521),
        .b(new_Jinkela_wire_522),
        .e(new_Jinkela_wire_523)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(N460),
        .b(new_Jinkela_wire_572),
        .c(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_14035 (
        .din(new_Jinkela_wire_16722),
        .dout(new_Jinkela_wire_16723)
    );

    bfr new_Jinkela_buffer_13967 (
        .din(new_Jinkela_wire_16650),
        .dout(new_Jinkela_wire_16651)
    );

    spl4L new_Jinkela_splitter_134 (
        .a(new_Jinkela_wire_524),
        .c(new_Jinkela_wire_525),
        .d(new_Jinkela_wire_526),
        .b(new_Jinkela_wire_527),
        .e(new_Jinkela_wire_528)
    );

    bfr new_Jinkela_buffer_3571 (
        .din(new_Jinkela_wire_4752),
        .dout(new_Jinkela_wire_4753)
    );

    bfr new_Jinkela_buffer_3768 (
        .din(_0562_),
        .dout(new_Jinkela_wire_4982)
    );

    bfr new_Jinkela_buffer_3572 (
        .din(new_Jinkela_wire_4753),
        .dout(new_Jinkela_wire_4754)
    );

    bfr new_Jinkela_buffer_3654 (
        .din(new_Jinkela_wire_4847),
        .dout(new_Jinkela_wire_4848)
    );

    bfr new_Jinkela_buffer_3573 (
        .din(new_Jinkela_wire_4754),
        .dout(new_Jinkela_wire_4755)
    );

    bfr new_Jinkela_buffer_3702 (
        .din(_0778_),
        .dout(new_Jinkela_wire_4914)
    );

    bfr new_Jinkela_buffer_3574 (
        .din(new_Jinkela_wire_4755),
        .dout(new_Jinkela_wire_4756)
    );

    bfr new_Jinkela_buffer_3655 (
        .din(new_Jinkela_wire_4848),
        .dout(new_Jinkela_wire_4849)
    );

    bfr new_Jinkela_buffer_3575 (
        .din(new_Jinkela_wire_4756),
        .dout(new_Jinkela_wire_4757)
    );

    spl2 new_Jinkela_splitter_457 (
        .a(_1603_),
        .b(new_Jinkela_wire_4986),
        .c(new_Jinkela_wire_4987)
    );

    bfr new_Jinkela_buffer_3576 (
        .din(new_Jinkela_wire_4757),
        .dout(new_Jinkela_wire_4758)
    );

    bfr new_Jinkela_buffer_3656 (
        .din(new_Jinkela_wire_4849),
        .dout(new_Jinkela_wire_4850)
    );

    bfr new_Jinkela_buffer_3577 (
        .din(new_Jinkela_wire_4758),
        .dout(new_Jinkela_wire_4759)
    );

    bfr new_Jinkela_buffer_3703 (
        .din(new_Jinkela_wire_4914),
        .dout(new_Jinkela_wire_4915)
    );

    bfr new_Jinkela_buffer_3578 (
        .din(new_Jinkela_wire_4759),
        .dout(new_Jinkela_wire_4760)
    );

    bfr new_Jinkela_buffer_3657 (
        .din(new_Jinkela_wire_4850),
        .dout(new_Jinkela_wire_4851)
    );

    bfr new_Jinkela_buffer_3579 (
        .din(new_Jinkela_wire_4760),
        .dout(new_Jinkela_wire_4761)
    );

    bfr new_Jinkela_buffer_3770 (
        .din(_1179_),
        .dout(new_Jinkela_wire_4988)
    );

    bfr new_Jinkela_buffer_3580 (
        .din(new_Jinkela_wire_4761),
        .dout(new_Jinkela_wire_4762)
    );

    bfr new_Jinkela_buffer_3658 (
        .din(new_Jinkela_wire_4851),
        .dout(new_Jinkela_wire_4852)
    );

    bfr new_Jinkela_buffer_3581 (
        .din(new_Jinkela_wire_4762),
        .dout(new_Jinkela_wire_4763)
    );

    bfr new_Jinkela_buffer_3704 (
        .din(new_Jinkela_wire_4915),
        .dout(new_Jinkela_wire_4916)
    );

    bfr new_Jinkela_buffer_3582 (
        .din(new_Jinkela_wire_4763),
        .dout(new_Jinkela_wire_4764)
    );

    bfr new_Jinkela_buffer_3659 (
        .din(new_Jinkela_wire_4852),
        .dout(new_Jinkela_wire_4853)
    );

    bfr new_Jinkela_buffer_3583 (
        .din(new_Jinkela_wire_4764),
        .dout(new_Jinkela_wire_4765)
    );

    bfr new_Jinkela_buffer_3769 (
        .din(new_Jinkela_wire_4982),
        .dout(new_Jinkela_wire_4983)
    );

    spl2 new_Jinkela_splitter_458 (
        .a(_0470_),
        .b(new_Jinkela_wire_4989),
        .c(new_Jinkela_wire_4990)
    );

    bfr new_Jinkela_buffer_3584 (
        .din(new_Jinkela_wire_4765),
        .dout(new_Jinkela_wire_4766)
    );

    bfr new_Jinkela_buffer_3660 (
        .din(new_Jinkela_wire_4853),
        .dout(new_Jinkela_wire_4854)
    );

    bfr new_Jinkela_buffer_3585 (
        .din(new_Jinkela_wire_4766),
        .dout(new_Jinkela_wire_4767)
    );

    bfr new_Jinkela_buffer_3705 (
        .din(new_Jinkela_wire_4916),
        .dout(new_Jinkela_wire_4917)
    );

    bfr new_Jinkela_buffer_3586 (
        .din(new_Jinkela_wire_4767),
        .dout(new_Jinkela_wire_4768)
    );

    bfr new_Jinkela_buffer_3661 (
        .din(new_Jinkela_wire_4854),
        .dout(new_Jinkela_wire_4855)
    );

    bfr new_Jinkela_buffer_3587 (
        .din(new_Jinkela_wire_4768),
        .dout(new_Jinkela_wire_4769)
    );

    bfr new_Jinkela_buffer_3588 (
        .din(new_Jinkela_wire_4769),
        .dout(new_Jinkela_wire_4770)
    );

    bfr new_Jinkela_buffer_3662 (
        .din(new_Jinkela_wire_4855),
        .dout(new_Jinkela_wire_4856)
    );

    bfr new_Jinkela_buffer_3589 (
        .din(new_Jinkela_wire_4770),
        .dout(new_Jinkela_wire_4771)
    );

    bfr new_Jinkela_buffer_3706 (
        .din(new_Jinkela_wire_4917),
        .dout(new_Jinkela_wire_4918)
    );

    bfr new_Jinkela_buffer_3590 (
        .din(new_Jinkela_wire_4771),
        .dout(new_Jinkela_wire_4772)
    );

    bfr new_Jinkela_buffer_3663 (
        .din(new_Jinkela_wire_4856),
        .dout(new_Jinkela_wire_4857)
    );

    bfr new_Jinkela_buffer_3591 (
        .din(new_Jinkela_wire_4772),
        .dout(new_Jinkela_wire_4773)
    );

    spl2 new_Jinkela_splitter_456 (
        .a(new_Jinkela_wire_4983),
        .b(new_Jinkela_wire_4984),
        .c(new_Jinkela_wire_4985)
    );

    bfr new_Jinkela_buffer_6994 (
        .din(new_Jinkela_wire_8747),
        .dout(new_Jinkela_wire_8748)
    );

    spl2 new_Jinkela_splitter_1530 (
        .a(_1615_),
        .b(new_Jinkela_wire_20960),
        .c(new_Jinkela_wire_20961)
    );

    bfr new_Jinkela_buffer_7086 (
        .din(new_Jinkela_wire_8861),
        .dout(new_Jinkela_wire_8862)
    );

    bfr new_Jinkela_buffer_17358 (
        .din(new_Jinkela_wire_20706),
        .dout(new_Jinkela_wire_20707)
    );

    bfr new_Jinkela_buffer_6995 (
        .din(new_Jinkela_wire_8748),
        .dout(new_Jinkela_wire_8749)
    );

    bfr new_Jinkela_buffer_17461 (
        .din(new_Jinkela_wire_20815),
        .dout(new_Jinkela_wire_20816)
    );

    bfr new_Jinkela_buffer_7030 (
        .din(new_Jinkela_wire_8791),
        .dout(new_Jinkela_wire_8792)
    );

    bfr new_Jinkela_buffer_17359 (
        .din(new_Jinkela_wire_20707),
        .dout(new_Jinkela_wire_20708)
    );

    bfr new_Jinkela_buffer_6996 (
        .din(new_Jinkela_wire_8749),
        .dout(new_Jinkela_wire_8750)
    );

    bfr new_Jinkela_buffer_17547 (
        .din(_0631_),
        .dout(new_Jinkela_wire_20908)
    );

    bfr new_Jinkela_buffer_7094 (
        .din(new_Jinkela_wire_8873),
        .dout(new_Jinkela_wire_8874)
    );

    bfr new_Jinkela_buffer_17360 (
        .din(new_Jinkela_wire_20708),
        .dout(new_Jinkela_wire_20709)
    );

    bfr new_Jinkela_buffer_6997 (
        .din(new_Jinkela_wire_8750),
        .dout(new_Jinkela_wire_8751)
    );

    bfr new_Jinkela_buffer_17462 (
        .din(new_Jinkela_wire_20816),
        .dout(new_Jinkela_wire_20817)
    );

    bfr new_Jinkela_buffer_7031 (
        .din(new_Jinkela_wire_8792),
        .dout(new_Jinkela_wire_8793)
    );

    bfr new_Jinkela_buffer_17361 (
        .din(new_Jinkela_wire_20709),
        .dout(new_Jinkela_wire_20710)
    );

    bfr new_Jinkela_buffer_6998 (
        .din(new_Jinkela_wire_8751),
        .dout(new_Jinkela_wire_8752)
    );

    spl2 new_Jinkela_splitter_1531 (
        .a(_0475_),
        .b(new_Jinkela_wire_20962),
        .c(new_Jinkela_wire_20963)
    );

    spl2 new_Jinkela_splitter_737 (
        .a(new_Jinkela_wire_8862),
        .b(new_Jinkela_wire_8863),
        .c(new_Jinkela_wire_8864)
    );

    bfr new_Jinkela_buffer_17362 (
        .din(new_Jinkela_wire_20710),
        .dout(new_Jinkela_wire_20711)
    );

    bfr new_Jinkela_buffer_6999 (
        .din(new_Jinkela_wire_8752),
        .dout(new_Jinkela_wire_8753)
    );

    bfr new_Jinkela_buffer_17463 (
        .din(new_Jinkela_wire_20817),
        .dout(new_Jinkela_wire_20818)
    );

    bfr new_Jinkela_buffer_7032 (
        .din(new_Jinkela_wire_8793),
        .dout(new_Jinkela_wire_8794)
    );

    bfr new_Jinkela_buffer_17363 (
        .din(new_Jinkela_wire_20711),
        .dout(new_Jinkela_wire_20712)
    );

    bfr new_Jinkela_buffer_7000 (
        .din(new_Jinkela_wire_8753),
        .dout(new_Jinkela_wire_8754)
    );

    bfr new_Jinkela_buffer_17548 (
        .din(new_Jinkela_wire_20908),
        .dout(new_Jinkela_wire_20909)
    );

    bfr new_Jinkela_buffer_7186 (
        .din(_0955_),
        .dout(new_Jinkela_wire_8970)
    );

    bfr new_Jinkela_buffer_17364 (
        .din(new_Jinkela_wire_20712),
        .dout(new_Jinkela_wire_20713)
    );

    bfr new_Jinkela_buffer_7182 (
        .din(new_Jinkela_wire_8965),
        .dout(new_Jinkela_wire_8966)
    );

    bfr new_Jinkela_buffer_7001 (
        .din(new_Jinkela_wire_8754),
        .dout(new_Jinkela_wire_8755)
    );

    bfr new_Jinkela_buffer_17464 (
        .din(new_Jinkela_wire_20818),
        .dout(new_Jinkela_wire_20819)
    );

    bfr new_Jinkela_buffer_7033 (
        .din(new_Jinkela_wire_8794),
        .dout(new_Jinkela_wire_8795)
    );

    bfr new_Jinkela_buffer_17365 (
        .din(new_Jinkela_wire_20713),
        .dout(new_Jinkela_wire_20714)
    );

    bfr new_Jinkela_buffer_7002 (
        .din(new_Jinkela_wire_8755),
        .dout(new_Jinkela_wire_8756)
    );

    bfr new_Jinkela_buffer_17607 (
        .din(new_Jinkela_wire_20973),
        .dout(new_Jinkela_wire_20974)
    );

    bfr new_Jinkela_buffer_7091 (
        .din(new_Jinkela_wire_8870),
        .dout(new_Jinkela_wire_8871)
    );

    bfr new_Jinkela_buffer_17366 (
        .din(new_Jinkela_wire_20714),
        .dout(new_Jinkela_wire_20715)
    );

    bfr new_Jinkela_buffer_7003 (
        .din(new_Jinkela_wire_8756),
        .dout(new_Jinkela_wire_8757)
    );

    bfr new_Jinkela_buffer_17465 (
        .din(new_Jinkela_wire_20819),
        .dout(new_Jinkela_wire_20820)
    );

    bfr new_Jinkela_buffer_7034 (
        .din(new_Jinkela_wire_8795),
        .dout(new_Jinkela_wire_8796)
    );

    bfr new_Jinkela_buffer_17367 (
        .din(new_Jinkela_wire_20715),
        .dout(new_Jinkela_wire_20716)
    );

    spl2 new_Jinkela_splitter_726 (
        .a(new_Jinkela_wire_8757),
        .b(new_Jinkela_wire_8758),
        .c(new_Jinkela_wire_8759)
    );

    bfr new_Jinkela_buffer_17549 (
        .din(new_Jinkela_wire_20909),
        .dout(new_Jinkela_wire_20910)
    );

    bfr new_Jinkela_buffer_7035 (
        .din(new_Jinkela_wire_8796),
        .dout(new_Jinkela_wire_8797)
    );

    bfr new_Jinkela_buffer_17368 (
        .din(new_Jinkela_wire_20716),
        .dout(new_Jinkela_wire_20717)
    );

    bfr new_Jinkela_buffer_7092 (
        .din(new_Jinkela_wire_8871),
        .dout(new_Jinkela_wire_8872)
    );

    bfr new_Jinkela_buffer_17466 (
        .din(new_Jinkela_wire_20820),
        .dout(new_Jinkela_wire_20821)
    );

    bfr new_Jinkela_buffer_7095 (
        .din(new_Jinkela_wire_8874),
        .dout(new_Jinkela_wire_8875)
    );

    bfr new_Jinkela_buffer_17369 (
        .din(new_Jinkela_wire_20717),
        .dout(new_Jinkela_wire_20718)
    );

    bfr new_Jinkela_buffer_7036 (
        .din(new_Jinkela_wire_8797),
        .dout(new_Jinkela_wire_8798)
    );

    bfr new_Jinkela_buffer_17370 (
        .din(new_Jinkela_wire_20718),
        .dout(new_Jinkela_wire_20719)
    );

    bfr new_Jinkela_buffer_7037 (
        .din(new_Jinkela_wire_8798),
        .dout(new_Jinkela_wire_8799)
    );

    bfr new_Jinkela_buffer_17467 (
        .din(new_Jinkela_wire_20821),
        .dout(new_Jinkela_wire_20822)
    );

    bfr new_Jinkela_buffer_7096 (
        .din(new_Jinkela_wire_8875),
        .dout(new_Jinkela_wire_8876)
    );

    bfr new_Jinkela_buffer_17371 (
        .din(new_Jinkela_wire_20719),
        .dout(new_Jinkela_wire_20720)
    );

    bfr new_Jinkela_buffer_7038 (
        .din(new_Jinkela_wire_8799),
        .dout(new_Jinkela_wire_8800)
    );

    bfr new_Jinkela_buffer_17550 (
        .din(new_Jinkela_wire_20910),
        .dout(new_Jinkela_wire_20911)
    );

    bfr new_Jinkela_buffer_17372 (
        .din(new_Jinkela_wire_20720),
        .dout(new_Jinkela_wire_20721)
    );

    spl2 new_Jinkela_splitter_742 (
        .a(_1383_),
        .b(new_Jinkela_wire_9012),
        .c(new_Jinkela_wire_9013)
    );

    bfr new_Jinkela_buffer_7039 (
        .din(new_Jinkela_wire_8800),
        .dout(new_Jinkela_wire_8801)
    );

    bfr new_Jinkela_buffer_17468 (
        .din(new_Jinkela_wire_20822),
        .dout(new_Jinkela_wire_20823)
    );

    bfr new_Jinkela_buffer_7097 (
        .din(new_Jinkela_wire_8876),
        .dout(new_Jinkela_wire_8877)
    );

    bfr new_Jinkela_buffer_17373 (
        .din(new_Jinkela_wire_20721),
        .dout(new_Jinkela_wire_20722)
    );

    bfr new_Jinkela_buffer_7040 (
        .din(new_Jinkela_wire_8801),
        .dout(new_Jinkela_wire_8802)
    );

    bfr new_Jinkela_buffer_17597 (
        .din(new_Jinkela_wire_20963),
        .dout(new_Jinkela_wire_20964)
    );

    bfr new_Jinkela_buffer_17374 (
        .din(new_Jinkela_wire_20722),
        .dout(new_Jinkela_wire_20723)
    );

    spl2 new_Jinkela_splitter_744 (
        .a(_1090_),
        .b(new_Jinkela_wire_9017),
        .c(new_Jinkela_wire_9018)
    );

    bfr new_Jinkela_buffer_7041 (
        .din(new_Jinkela_wire_8802),
        .dout(new_Jinkela_wire_8803)
    );

    bfr new_Jinkela_buffer_17469 (
        .din(new_Jinkela_wire_20823),
        .dout(new_Jinkela_wire_20824)
    );

    bfr new_Jinkela_buffer_7098 (
        .din(new_Jinkela_wire_8877),
        .dout(new_Jinkela_wire_8878)
    );

    bfr new_Jinkela_buffer_17375 (
        .din(new_Jinkela_wire_20723),
        .dout(new_Jinkela_wire_20724)
    );

    bfr new_Jinkela_buffer_7042 (
        .din(new_Jinkela_wire_8803),
        .dout(new_Jinkela_wire_8804)
    );

    bfr new_Jinkela_buffer_17551 (
        .din(new_Jinkela_wire_20911),
        .dout(new_Jinkela_wire_20912)
    );

    bfr new_Jinkela_buffer_7183 (
        .din(new_Jinkela_wire_8966),
        .dout(new_Jinkela_wire_8967)
    );

    bfr new_Jinkela_buffer_17376 (
        .din(new_Jinkela_wire_20724),
        .dout(new_Jinkela_wire_20725)
    );

    bfr new_Jinkela_buffer_7043 (
        .din(new_Jinkela_wire_8804),
        .dout(new_Jinkela_wire_8805)
    );

    bfr new_Jinkela_buffer_17470 (
        .din(new_Jinkela_wire_20824),
        .dout(new_Jinkela_wire_20825)
    );

    bfr new_Jinkela_buffer_7099 (
        .din(new_Jinkela_wire_8878),
        .dout(new_Jinkela_wire_8879)
    );

    bfr new_Jinkela_buffer_17377 (
        .din(new_Jinkela_wire_20725),
        .dout(new_Jinkela_wire_20726)
    );

    bfr new_Jinkela_buffer_7044 (
        .din(new_Jinkela_wire_8805),
        .dout(new_Jinkela_wire_8806)
    );

    bfr new_Jinkela_buffer_17628 (
        .din(new_Jinkela_wire_20996),
        .dout(new_Jinkela_wire_20997)
    );

    bfr new_Jinkela_buffer_7187 (
        .din(new_Jinkela_wire_8970),
        .dout(new_Jinkela_wire_8971)
    );

    bfr new_Jinkela_buffer_17378 (
        .din(new_Jinkela_wire_20726),
        .dout(new_Jinkela_wire_20727)
    );

    bfr new_Jinkela_buffer_3592 (
        .din(new_Jinkela_wire_4773),
        .dout(new_Jinkela_wire_4774)
    );

    bfr new_Jinkela_buffer_14098 (
        .din(new_Jinkela_wire_16801),
        .dout(new_Jinkela_wire_16802)
    );

    bfr new_Jinkela_buffer_13968 (
        .din(new_Jinkela_wire_16651),
        .dout(new_Jinkela_wire_16652)
    );

    bfr new_Jinkela_buffer_3664 (
        .din(new_Jinkela_wire_4857),
        .dout(new_Jinkela_wire_4858)
    );

    bfr new_Jinkela_buffer_3593 (
        .din(new_Jinkela_wire_4774),
        .dout(new_Jinkela_wire_4775)
    );

    bfr new_Jinkela_buffer_14036 (
        .din(new_Jinkela_wire_16723),
        .dout(new_Jinkela_wire_16724)
    );

    bfr new_Jinkela_buffer_13969 (
        .din(new_Jinkela_wire_16652),
        .dout(new_Jinkela_wire_16653)
    );

    bfr new_Jinkela_buffer_3707 (
        .din(new_Jinkela_wire_4918),
        .dout(new_Jinkela_wire_4919)
    );

    bfr new_Jinkela_buffer_3594 (
        .din(new_Jinkela_wire_4775),
        .dout(new_Jinkela_wire_4776)
    );

    spl2 new_Jinkela_splitter_1205 (
        .a(_0759_),
        .b(new_Jinkela_wire_16874),
        .c(new_Jinkela_wire_16875)
    );

    bfr new_Jinkela_buffer_13970 (
        .din(new_Jinkela_wire_16653),
        .dout(new_Jinkela_wire_16654)
    );

    bfr new_Jinkela_buffer_3665 (
        .din(new_Jinkela_wire_4858),
        .dout(new_Jinkela_wire_4859)
    );

    bfr new_Jinkela_buffer_3595 (
        .din(new_Jinkela_wire_4776),
        .dout(new_Jinkela_wire_4777)
    );

    bfr new_Jinkela_buffer_14037 (
        .din(new_Jinkela_wire_16724),
        .dout(new_Jinkela_wire_16725)
    );

    bfr new_Jinkela_buffer_13971 (
        .din(new_Jinkela_wire_16654),
        .dout(new_Jinkela_wire_16655)
    );

    bfr new_Jinkela_buffer_3596 (
        .din(new_Jinkela_wire_4777),
        .dout(new_Jinkela_wire_4778)
    );

    bfr new_Jinkela_buffer_14099 (
        .din(new_Jinkela_wire_16802),
        .dout(new_Jinkela_wire_16803)
    );

    bfr new_Jinkela_buffer_13972 (
        .din(new_Jinkela_wire_16655),
        .dout(new_Jinkela_wire_16656)
    );

    bfr new_Jinkela_buffer_3666 (
        .din(new_Jinkela_wire_4859),
        .dout(new_Jinkela_wire_4860)
    );

    bfr new_Jinkela_buffer_3597 (
        .din(new_Jinkela_wire_4778),
        .dout(new_Jinkela_wire_4779)
    );

    bfr new_Jinkela_buffer_14038 (
        .din(new_Jinkela_wire_16725),
        .dout(new_Jinkela_wire_16726)
    );

    bfr new_Jinkela_buffer_13973 (
        .din(new_Jinkela_wire_16656),
        .dout(new_Jinkela_wire_16657)
    );

    bfr new_Jinkela_buffer_3708 (
        .din(new_Jinkela_wire_4919),
        .dout(new_Jinkela_wire_4920)
    );

    bfr new_Jinkela_buffer_3598 (
        .din(new_Jinkela_wire_4779),
        .dout(new_Jinkela_wire_4780)
    );

    bfr new_Jinkela_buffer_13974 (
        .din(new_Jinkela_wire_16657),
        .dout(new_Jinkela_wire_16658)
    );

    bfr new_Jinkela_buffer_3667 (
        .din(new_Jinkela_wire_4860),
        .dout(new_Jinkela_wire_4861)
    );

    bfr new_Jinkela_buffer_14160 (
        .din(_0650_),
        .dout(new_Jinkela_wire_16872)
    );

    bfr new_Jinkela_buffer_3599 (
        .din(new_Jinkela_wire_4780),
        .dout(new_Jinkela_wire_4781)
    );

    bfr new_Jinkela_buffer_14039 (
        .din(new_Jinkela_wire_16726),
        .dout(new_Jinkela_wire_16727)
    );

    bfr new_Jinkela_buffer_13975 (
        .din(new_Jinkela_wire_16658),
        .dout(new_Jinkela_wire_16659)
    );

    spl2 new_Jinkela_splitter_459 (
        .a(_0002_),
        .b(new_Jinkela_wire_4995),
        .c(new_Jinkela_wire_4996)
    );

    bfr new_Jinkela_buffer_3771 (
        .din(new_Jinkela_wire_4990),
        .dout(new_Jinkela_wire_4991)
    );

    bfr new_Jinkela_buffer_3600 (
        .din(new_Jinkela_wire_4781),
        .dout(new_Jinkela_wire_4782)
    );

    bfr new_Jinkela_buffer_14100 (
        .din(new_Jinkela_wire_16803),
        .dout(new_Jinkela_wire_16804)
    );

    bfr new_Jinkela_buffer_13976 (
        .din(new_Jinkela_wire_16659),
        .dout(new_Jinkela_wire_16660)
    );

    bfr new_Jinkela_buffer_3668 (
        .din(new_Jinkela_wire_4861),
        .dout(new_Jinkela_wire_4862)
    );

    bfr new_Jinkela_buffer_3601 (
        .din(new_Jinkela_wire_4782),
        .dout(new_Jinkela_wire_4783)
    );

    bfr new_Jinkela_buffer_14040 (
        .din(new_Jinkela_wire_16727),
        .dout(new_Jinkela_wire_16728)
    );

    bfr new_Jinkela_buffer_13977 (
        .din(new_Jinkela_wire_16660),
        .dout(new_Jinkela_wire_16661)
    );

    bfr new_Jinkela_buffer_3709 (
        .din(new_Jinkela_wire_4920),
        .dout(new_Jinkela_wire_4921)
    );

    bfr new_Jinkela_buffer_3602 (
        .din(new_Jinkela_wire_4783),
        .dout(new_Jinkela_wire_4784)
    );

    bfr new_Jinkela_buffer_13978 (
        .din(new_Jinkela_wire_16661),
        .dout(new_Jinkela_wire_16662)
    );

    bfr new_Jinkela_buffer_3669 (
        .din(new_Jinkela_wire_4862),
        .dout(new_Jinkela_wire_4863)
    );

    bfr new_Jinkela_buffer_14161 (
        .din(_0247_),
        .dout(new_Jinkela_wire_16873)
    );

    bfr new_Jinkela_buffer_3603 (
        .din(new_Jinkela_wire_4784),
        .dout(new_Jinkela_wire_4785)
    );

    bfr new_Jinkela_buffer_14041 (
        .din(new_Jinkela_wire_16728),
        .dout(new_Jinkela_wire_16729)
    );

    bfr new_Jinkela_buffer_13979 (
        .din(new_Jinkela_wire_16662),
        .dout(new_Jinkela_wire_16663)
    );

    bfr new_Jinkela_buffer_3775 (
        .din(_1673_),
        .dout(new_Jinkela_wire_4997)
    );

    bfr new_Jinkela_buffer_3604 (
        .din(new_Jinkela_wire_4785),
        .dout(new_Jinkela_wire_4786)
    );

    bfr new_Jinkela_buffer_14101 (
        .din(new_Jinkela_wire_16804),
        .dout(new_Jinkela_wire_16805)
    );

    bfr new_Jinkela_buffer_13980 (
        .din(new_Jinkela_wire_16663),
        .dout(new_Jinkela_wire_16664)
    );

    bfr new_Jinkela_buffer_3670 (
        .din(new_Jinkela_wire_4863),
        .dout(new_Jinkela_wire_4864)
    );

    bfr new_Jinkela_buffer_3605 (
        .din(new_Jinkela_wire_4786),
        .dout(new_Jinkela_wire_4787)
    );

    bfr new_Jinkela_buffer_14042 (
        .din(new_Jinkela_wire_16729),
        .dout(new_Jinkela_wire_16730)
    );

    bfr new_Jinkela_buffer_13981 (
        .din(new_Jinkela_wire_16664),
        .dout(new_Jinkela_wire_16665)
    );

    bfr new_Jinkela_buffer_3710 (
        .din(new_Jinkela_wire_4921),
        .dout(new_Jinkela_wire_4922)
    );

    bfr new_Jinkela_buffer_3606 (
        .din(new_Jinkela_wire_4787),
        .dout(new_Jinkela_wire_4788)
    );

    spl2 new_Jinkela_splitter_1206 (
        .a(_0377_),
        .b(new_Jinkela_wire_16904),
        .c(new_Jinkela_wire_16905)
    );

    bfr new_Jinkela_buffer_13982 (
        .din(new_Jinkela_wire_16665),
        .dout(new_Jinkela_wire_16666)
    );

    bfr new_Jinkela_buffer_3671 (
        .din(new_Jinkela_wire_4864),
        .dout(new_Jinkela_wire_4865)
    );

    bfr new_Jinkela_buffer_14162 (
        .din(new_Jinkela_wire_16875),
        .dout(new_Jinkela_wire_16876)
    );

    bfr new_Jinkela_buffer_3607 (
        .din(new_Jinkela_wire_4788),
        .dout(new_Jinkela_wire_4789)
    );

    bfr new_Jinkela_buffer_14043 (
        .din(new_Jinkela_wire_16730),
        .dout(new_Jinkela_wire_16731)
    );

    bfr new_Jinkela_buffer_13983 (
        .din(new_Jinkela_wire_16666),
        .dout(new_Jinkela_wire_16667)
    );

    bfr new_Jinkela_buffer_3776 (
        .din(_0789_),
        .dout(new_Jinkela_wire_4998)
    );

    bfr new_Jinkela_buffer_3608 (
        .din(new_Jinkela_wire_4789),
        .dout(new_Jinkela_wire_4790)
    );

    bfr new_Jinkela_buffer_14102 (
        .din(new_Jinkela_wire_16805),
        .dout(new_Jinkela_wire_16806)
    );

    bfr new_Jinkela_buffer_13984 (
        .din(new_Jinkela_wire_16667),
        .dout(new_Jinkela_wire_16668)
    );

    bfr new_Jinkela_buffer_3672 (
        .din(new_Jinkela_wire_4865),
        .dout(new_Jinkela_wire_4866)
    );

    bfr new_Jinkela_buffer_3609 (
        .din(new_Jinkela_wire_4790),
        .dout(new_Jinkela_wire_4791)
    );

    bfr new_Jinkela_buffer_14044 (
        .din(new_Jinkela_wire_16731),
        .dout(new_Jinkela_wire_16732)
    );

    bfr new_Jinkela_buffer_13985 (
        .din(new_Jinkela_wire_16668),
        .dout(new_Jinkela_wire_16669)
    );

    bfr new_Jinkela_buffer_3711 (
        .din(new_Jinkela_wire_4922),
        .dout(new_Jinkela_wire_4923)
    );

    bfr new_Jinkela_buffer_3610 (
        .din(new_Jinkela_wire_4791),
        .dout(new_Jinkela_wire_4792)
    );

    bfr new_Jinkela_buffer_13986 (
        .din(new_Jinkela_wire_16669),
        .dout(new_Jinkela_wire_16670)
    );

    bfr new_Jinkela_buffer_3673 (
        .din(new_Jinkela_wire_4866),
        .dout(new_Jinkela_wire_4867)
    );

    bfr new_Jinkela_buffer_3611 (
        .din(new_Jinkela_wire_4792),
        .dout(new_Jinkela_wire_4793)
    );

    bfr new_Jinkela_buffer_14045 (
        .din(new_Jinkela_wire_16732),
        .dout(new_Jinkela_wire_16733)
    );

    bfr new_Jinkela_buffer_13987 (
        .din(new_Jinkela_wire_16670),
        .dout(new_Jinkela_wire_16671)
    );

    bfr new_Jinkela_buffer_3772 (
        .din(new_Jinkela_wire_4991),
        .dout(new_Jinkela_wire_4992)
    );

    bfr new_Jinkela_buffer_3612 (
        .din(new_Jinkela_wire_4793),
        .dout(new_Jinkela_wire_4794)
    );

    bfr new_Jinkela_buffer_14103 (
        .din(new_Jinkela_wire_16806),
        .dout(new_Jinkela_wire_16807)
    );

    bfr new_Jinkela_buffer_13988 (
        .din(new_Jinkela_wire_16671),
        .dout(new_Jinkela_wire_16672)
    );

    bfr new_Jinkela_buffer_3674 (
        .din(new_Jinkela_wire_4867),
        .dout(new_Jinkela_wire_4868)
    );

    bfr new_Jinkela_buffer_9608 (
        .din(new_Jinkela_wire_11701),
        .dout(new_Jinkela_wire_11702)
    );

    bfr new_Jinkela_buffer_9924 (
        .din(new_Jinkela_wire_12047),
        .dout(new_Jinkela_wire_12048)
    );

    bfr new_Jinkela_buffer_9609 (
        .din(new_Jinkela_wire_11702),
        .dout(new_Jinkela_wire_11703)
    );

    bfr new_Jinkela_buffer_9668 (
        .din(new_Jinkela_wire_11767),
        .dout(new_Jinkela_wire_11768)
    );

    bfr new_Jinkela_buffer_9610 (
        .din(new_Jinkela_wire_11703),
        .dout(new_Jinkela_wire_11704)
    );

    bfr new_Jinkela_buffer_9745 (
        .din(new_Jinkela_wire_11854),
        .dout(new_Jinkela_wire_11855)
    );

    bfr new_Jinkela_buffer_9611 (
        .din(new_Jinkela_wire_11704),
        .dout(new_Jinkela_wire_11705)
    );

    bfr new_Jinkela_buffer_9669 (
        .din(new_Jinkela_wire_11768),
        .dout(new_Jinkela_wire_11769)
    );

    bfr new_Jinkela_buffer_9612 (
        .din(new_Jinkela_wire_11705),
        .dout(new_Jinkela_wire_11706)
    );

    bfr new_Jinkela_buffer_9848 (
        .din(new_Jinkela_wire_11967),
        .dout(new_Jinkela_wire_11968)
    );

    bfr new_Jinkela_buffer_9613 (
        .din(new_Jinkela_wire_11706),
        .dout(new_Jinkela_wire_11707)
    );

    bfr new_Jinkela_buffer_9670 (
        .din(new_Jinkela_wire_11769),
        .dout(new_Jinkela_wire_11770)
    );

    bfr new_Jinkela_buffer_9614 (
        .din(new_Jinkela_wire_11707),
        .dout(new_Jinkela_wire_11708)
    );

    bfr new_Jinkela_buffer_9746 (
        .din(new_Jinkela_wire_11855),
        .dout(new_Jinkela_wire_11856)
    );

    bfr new_Jinkela_buffer_9615 (
        .din(new_Jinkela_wire_11708),
        .dout(new_Jinkela_wire_11709)
    );

    bfr new_Jinkela_buffer_9671 (
        .din(new_Jinkela_wire_11770),
        .dout(new_Jinkela_wire_11771)
    );

    bfr new_Jinkela_buffer_9616 (
        .din(new_Jinkela_wire_11709),
        .dout(new_Jinkela_wire_11710)
    );

    spl2 new_Jinkela_splitter_913 (
        .a(_0923_),
        .b(new_Jinkela_wire_12056),
        .c(new_Jinkela_wire_12057)
    );

    bfr new_Jinkela_buffer_9617 (
        .din(new_Jinkela_wire_11710),
        .dout(new_Jinkela_wire_11711)
    );

    bfr new_Jinkela_buffer_9672 (
        .din(new_Jinkela_wire_11771),
        .dout(new_Jinkela_wire_11772)
    );

    bfr new_Jinkela_buffer_9618 (
        .din(new_Jinkela_wire_11711),
        .dout(new_Jinkela_wire_11712)
    );

    bfr new_Jinkela_buffer_9747 (
        .din(new_Jinkela_wire_11856),
        .dout(new_Jinkela_wire_11857)
    );

    bfr new_Jinkela_buffer_9619 (
        .din(new_Jinkela_wire_11712),
        .dout(new_Jinkela_wire_11713)
    );

    bfr new_Jinkela_buffer_9673 (
        .din(new_Jinkela_wire_11772),
        .dout(new_Jinkela_wire_11773)
    );

    bfr new_Jinkela_buffer_9620 (
        .din(new_Jinkela_wire_11713),
        .dout(new_Jinkela_wire_11714)
    );

    bfr new_Jinkela_buffer_9849 (
        .din(new_Jinkela_wire_11968),
        .dout(new_Jinkela_wire_11969)
    );

    bfr new_Jinkela_buffer_9621 (
        .din(new_Jinkela_wire_11714),
        .dout(new_Jinkela_wire_11715)
    );

    bfr new_Jinkela_buffer_9674 (
        .din(new_Jinkela_wire_11773),
        .dout(new_Jinkela_wire_11774)
    );

    bfr new_Jinkela_buffer_9622 (
        .din(new_Jinkela_wire_11715),
        .dout(new_Jinkela_wire_11716)
    );

    bfr new_Jinkela_buffer_9748 (
        .din(new_Jinkela_wire_11857),
        .dout(new_Jinkela_wire_11858)
    );

    bfr new_Jinkela_buffer_9623 (
        .din(new_Jinkela_wire_11716),
        .dout(new_Jinkela_wire_11717)
    );

    bfr new_Jinkela_buffer_9675 (
        .din(new_Jinkela_wire_11774),
        .dout(new_Jinkela_wire_11775)
    );

    bfr new_Jinkela_buffer_9624 (
        .din(new_Jinkela_wire_11717),
        .dout(new_Jinkela_wire_11718)
    );

    bfr new_Jinkela_buffer_9925 (
        .din(new_Jinkela_wire_12048),
        .dout(new_Jinkela_wire_12049)
    );

    bfr new_Jinkela_buffer_9625 (
        .din(new_Jinkela_wire_11718),
        .dout(new_Jinkela_wire_11719)
    );

    bfr new_Jinkela_buffer_9676 (
        .din(new_Jinkela_wire_11775),
        .dout(new_Jinkela_wire_11776)
    );

    spl2 new_Jinkela_splitter_896 (
        .a(new_Jinkela_wire_11719),
        .b(new_Jinkela_wire_11720),
        .c(new_Jinkela_wire_11721)
    );

    bfr new_Jinkela_buffer_9677 (
        .din(new_Jinkela_wire_11776),
        .dout(new_Jinkela_wire_11777)
    );

    bfr new_Jinkela_buffer_9749 (
        .din(new_Jinkela_wire_11858),
        .dout(new_Jinkela_wire_11859)
    );

    bfr new_Jinkela_buffer_9850 (
        .din(new_Jinkela_wire_11969),
        .dout(new_Jinkela_wire_11970)
    );

    bfr new_Jinkela_buffer_9678 (
        .din(new_Jinkela_wire_11777),
        .dout(new_Jinkela_wire_11778)
    );

    bfr new_Jinkela_buffer_9750 (
        .din(new_Jinkela_wire_11859),
        .dout(new_Jinkela_wire_11860)
    );

    bfr new_Jinkela_buffer_6213 (
        .din(new_Jinkela_wire_7886),
        .dout(new_Jinkela_wire_7887)
    );

    bfr new_Jinkela_buffer_6154 (
        .din(new_Jinkela_wire_7811),
        .dout(new_Jinkela_wire_7812)
    );

    bfr new_Jinkela_buffer_6304 (
        .din(new_Jinkela_wire_7983),
        .dout(new_Jinkela_wire_7984)
    );

    bfr new_Jinkela_buffer_6155 (
        .din(new_Jinkela_wire_7812),
        .dout(new_Jinkela_wire_7813)
    );

    bfr new_Jinkela_buffer_6214 (
        .din(new_Jinkela_wire_7887),
        .dout(new_Jinkela_wire_7888)
    );

    bfr new_Jinkela_buffer_6156 (
        .din(new_Jinkela_wire_7813),
        .dout(new_Jinkela_wire_7814)
    );

    spl2 new_Jinkela_splitter_691 (
        .a(_1258_),
        .b(new_Jinkela_wire_8025),
        .c(new_Jinkela_wire_8026)
    );

    bfr new_Jinkela_buffer_6337 (
        .din(new_Jinkela_wire_8020),
        .dout(new_Jinkela_wire_8021)
    );

    bfr new_Jinkela_buffer_6157 (
        .din(new_Jinkela_wire_7814),
        .dout(new_Jinkela_wire_7815)
    );

    bfr new_Jinkela_buffer_6215 (
        .din(new_Jinkela_wire_7888),
        .dout(new_Jinkela_wire_7889)
    );

    bfr new_Jinkela_buffer_6158 (
        .din(new_Jinkela_wire_7815),
        .dout(new_Jinkela_wire_7816)
    );

    bfr new_Jinkela_buffer_6305 (
        .din(new_Jinkela_wire_7984),
        .dout(new_Jinkela_wire_7985)
    );

    bfr new_Jinkela_buffer_6159 (
        .din(new_Jinkela_wire_7816),
        .dout(new_Jinkela_wire_7817)
    );

    bfr new_Jinkela_buffer_6216 (
        .din(new_Jinkela_wire_7889),
        .dout(new_Jinkela_wire_7890)
    );

    bfr new_Jinkela_buffer_6160 (
        .din(new_Jinkela_wire_7817),
        .dout(new_Jinkela_wire_7818)
    );

    bfr new_Jinkela_buffer_6161 (
        .din(new_Jinkela_wire_7818),
        .dout(new_Jinkela_wire_7819)
    );

    bfr new_Jinkela_buffer_6217 (
        .din(new_Jinkela_wire_7890),
        .dout(new_Jinkela_wire_7891)
    );

    bfr new_Jinkela_buffer_6162 (
        .din(new_Jinkela_wire_7819),
        .dout(new_Jinkela_wire_7820)
    );

    bfr new_Jinkela_buffer_6306 (
        .din(new_Jinkela_wire_7985),
        .dout(new_Jinkela_wire_7986)
    );

    bfr new_Jinkela_buffer_6163 (
        .din(new_Jinkela_wire_7820),
        .dout(new_Jinkela_wire_7821)
    );

    bfr new_Jinkela_buffer_6218 (
        .din(new_Jinkela_wire_7891),
        .dout(new_Jinkela_wire_7892)
    );

    bfr new_Jinkela_buffer_6164 (
        .din(new_Jinkela_wire_7821),
        .dout(new_Jinkela_wire_7822)
    );

    spl2 new_Jinkela_splitter_692 (
        .a(_0616_),
        .b(new_Jinkela_wire_8027),
        .c(new_Jinkela_wire_8028)
    );

    bfr new_Jinkela_buffer_6165 (
        .din(new_Jinkela_wire_7822),
        .dout(new_Jinkela_wire_7823)
    );

    bfr new_Jinkela_buffer_6219 (
        .din(new_Jinkela_wire_7892),
        .dout(new_Jinkela_wire_7893)
    );

    bfr new_Jinkela_buffer_6166 (
        .din(new_Jinkela_wire_7823),
        .dout(new_Jinkela_wire_7824)
    );

    bfr new_Jinkela_buffer_6307 (
        .din(new_Jinkela_wire_7986),
        .dout(new_Jinkela_wire_7987)
    );

    bfr new_Jinkela_buffer_6167 (
        .din(new_Jinkela_wire_7824),
        .dout(new_Jinkela_wire_7825)
    );

    bfr new_Jinkela_buffer_6220 (
        .din(new_Jinkela_wire_7893),
        .dout(new_Jinkela_wire_7894)
    );

    bfr new_Jinkela_buffer_6168 (
        .din(new_Jinkela_wire_7825),
        .dout(new_Jinkela_wire_7826)
    );

    bfr new_Jinkela_buffer_6341 (
        .din(_0097_),
        .dout(new_Jinkela_wire_8029)
    );

    bfr new_Jinkela_buffer_6169 (
        .din(new_Jinkela_wire_7826),
        .dout(new_Jinkela_wire_7827)
    );

    bfr new_Jinkela_buffer_6221 (
        .din(new_Jinkela_wire_7894),
        .dout(new_Jinkela_wire_7895)
    );

    bfr new_Jinkela_buffer_6170 (
        .din(new_Jinkela_wire_7827),
        .dout(new_Jinkela_wire_7828)
    );

    bfr new_Jinkela_buffer_6308 (
        .din(new_Jinkela_wire_7987),
        .dout(new_Jinkela_wire_7988)
    );

    bfr new_Jinkela_buffer_6171 (
        .din(new_Jinkela_wire_7828),
        .dout(new_Jinkela_wire_7829)
    );

    bfr new_Jinkela_buffer_6222 (
        .din(new_Jinkela_wire_7895),
        .dout(new_Jinkela_wire_7896)
    );

    bfr new_Jinkela_buffer_6172 (
        .din(new_Jinkela_wire_7829),
        .dout(new_Jinkela_wire_7830)
    );

    bfr new_Jinkela_buffer_6338 (
        .din(new_Jinkela_wire_8021),
        .dout(new_Jinkela_wire_8022)
    );

    spl2 new_Jinkela_splitter_678 (
        .a(new_Jinkela_wire_7830),
        .b(new_Jinkela_wire_7831),
        .c(new_Jinkela_wire_7832)
    );

    bfr new_Jinkela_buffer_6309 (
        .din(new_Jinkela_wire_7988),
        .dout(new_Jinkela_wire_7989)
    );

    bfr new_Jinkela_buffer_6223 (
        .din(new_Jinkela_wire_7896),
        .dout(new_Jinkela_wire_7897)
    );

    bfr new_Jinkela_buffer_13116 (
        .din(new_Jinkela_wire_15649),
        .dout(new_Jinkela_wire_15650)
    );

    spl2 new_Jinkela_splitter_1148 (
        .a(_0997_),
        .b(new_Jinkela_wire_15837),
        .c(new_Jinkela_wire_15838)
    );

    bfr new_Jinkela_buffer_13117 (
        .din(new_Jinkela_wire_15650),
        .dout(new_Jinkela_wire_15651)
    );

    bfr new_Jinkela_buffer_13189 (
        .din(new_Jinkela_wire_15784),
        .dout(new_Jinkela_wire_15785)
    );

    bfr new_Jinkela_buffer_13118 (
        .din(new_Jinkela_wire_15651),
        .dout(new_Jinkela_wire_15652)
    );

    bfr new_Jinkela_buffer_13293 (
        .din(_0042_),
        .dout(new_Jinkela_wire_15893)
    );

    bfr new_Jinkela_buffer_13239 (
        .din(new_Jinkela_wire_15838),
        .dout(new_Jinkela_wire_15839)
    );

    bfr new_Jinkela_buffer_13119 (
        .din(new_Jinkela_wire_15652),
        .dout(new_Jinkela_wire_15653)
    );

    bfr new_Jinkela_buffer_13190 (
        .din(new_Jinkela_wire_15785),
        .dout(new_Jinkela_wire_15786)
    );

    bfr new_Jinkela_buffer_13120 (
        .din(new_Jinkela_wire_15653),
        .dout(new_Jinkela_wire_15654)
    );

    bfr new_Jinkela_buffer_13121 (
        .din(new_Jinkela_wire_15654),
        .dout(new_Jinkela_wire_15655)
    );

    bfr new_Jinkela_buffer_13191 (
        .din(new_Jinkela_wire_15786),
        .dout(new_Jinkela_wire_15787)
    );

    bfr new_Jinkela_buffer_13122 (
        .din(new_Jinkela_wire_15655),
        .dout(new_Jinkela_wire_15656)
    );

    bfr new_Jinkela_buffer_13294 (
        .din(_1458_),
        .dout(new_Jinkela_wire_15894)
    );

    bfr new_Jinkela_buffer_13123 (
        .din(new_Jinkela_wire_15656),
        .dout(new_Jinkela_wire_15657)
    );

    bfr new_Jinkela_buffer_13192 (
        .din(new_Jinkela_wire_15787),
        .dout(new_Jinkela_wire_15788)
    );

    bfr new_Jinkela_buffer_13124 (
        .din(new_Jinkela_wire_15657),
        .dout(new_Jinkela_wire_15658)
    );

    bfr new_Jinkela_buffer_13310 (
        .din(_0625_),
        .dout(new_Jinkela_wire_15912)
    );

    bfr new_Jinkela_buffer_13125 (
        .din(new_Jinkela_wire_15658),
        .dout(new_Jinkela_wire_15659)
    );

    bfr new_Jinkela_buffer_13193 (
        .din(new_Jinkela_wire_15788),
        .dout(new_Jinkela_wire_15789)
    );

    spl2 new_Jinkela_splitter_1116 (
        .a(new_Jinkela_wire_15659),
        .b(new_Jinkela_wire_15660),
        .c(new_Jinkela_wire_15661)
    );

    bfr new_Jinkela_buffer_13194 (
        .din(new_Jinkela_wire_15789),
        .dout(new_Jinkela_wire_15790)
    );

    bfr new_Jinkela_buffer_13240 (
        .din(new_Jinkela_wire_15839),
        .dout(new_Jinkela_wire_15840)
    );

    spl2 new_Jinkela_splitter_1151 (
        .a(_0735_),
        .b(new_Jinkela_wire_15994),
        .c(new_Jinkela_wire_15995)
    );

    bfr new_Jinkela_buffer_13195 (
        .din(new_Jinkela_wire_15790),
        .dout(new_Jinkela_wire_15791)
    );

    bfr new_Jinkela_buffer_13241 (
        .din(new_Jinkela_wire_15840),
        .dout(new_Jinkela_wire_15841)
    );

    bfr new_Jinkela_buffer_13196 (
        .din(new_Jinkela_wire_15791),
        .dout(new_Jinkela_wire_15792)
    );

    bfr new_Jinkela_buffer_13295 (
        .din(new_Jinkela_wire_15894),
        .dout(new_Jinkela_wire_15895)
    );

    bfr new_Jinkela_buffer_13197 (
        .din(new_Jinkela_wire_15792),
        .dout(new_Jinkela_wire_15793)
    );

    bfr new_Jinkela_buffer_13242 (
        .din(new_Jinkela_wire_15841),
        .dout(new_Jinkela_wire_15842)
    );

    bfr new_Jinkela_buffer_13198 (
        .din(new_Jinkela_wire_15793),
        .dout(new_Jinkela_wire_15794)
    );

    spl2 new_Jinkela_splitter_1152 (
        .a(_0279_),
        .b(new_Jinkela_wire_15996),
        .c(new_Jinkela_wire_15997)
    );

    bfr new_Jinkela_buffer_13199 (
        .din(new_Jinkela_wire_15794),
        .dout(new_Jinkela_wire_15795)
    );

    bfr new_Jinkela_buffer_13243 (
        .din(new_Jinkela_wire_15842),
        .dout(new_Jinkela_wire_15843)
    );

    bfr new_Jinkela_buffer_13200 (
        .din(new_Jinkela_wire_15795),
        .dout(new_Jinkela_wire_15796)
    );

    bfr new_Jinkela_buffer_13296 (
        .din(new_Jinkela_wire_15895),
        .dout(new_Jinkela_wire_15896)
    );

    bfr new_Jinkela_buffer_13201 (
        .din(new_Jinkela_wire_15796),
        .dout(new_Jinkela_wire_15797)
    );

    bfr new_Jinkela_buffer_13244 (
        .din(new_Jinkela_wire_15843),
        .dout(new_Jinkela_wire_15844)
    );

    bfr new_Jinkela_buffer_13202 (
        .din(new_Jinkela_wire_15797),
        .dout(new_Jinkela_wire_15798)
    );

    bfr new_Jinkela_buffer_13311 (
        .din(new_Jinkela_wire_15912),
        .dout(new_Jinkela_wire_15913)
    );

    bfr new_Jinkela_buffer_13203 (
        .din(new_Jinkela_wire_15798),
        .dout(new_Jinkela_wire_15799)
    );

    bfr new_Jinkela_buffer_13245 (
        .din(new_Jinkela_wire_15844),
        .dout(new_Jinkela_wire_15845)
    );

    and_ii _3054_ (
        .a(new_Jinkela_wire_13720),
        .b(new_Jinkela_wire_828),
        .c(_0309_)
    );

    or_bb _3053_ (
        .a(new_Jinkela_wire_19109),
        .b(new_Jinkela_wire_8019),
        .c(_0308_)
    );

    and_bb _3052_ (
        .a(new_Jinkela_wire_14197),
        .b(new_Jinkela_wire_4827),
        .c(_0306_)
    );

    bfr new_Jinkela_buffer_2805 (
        .din(new_Jinkela_wire_3854),
        .dout(new_Jinkela_wire_3855)
    );

    bfr new_Jinkela_buffer_2752 (
        .din(new_Jinkela_wire_3795),
        .dout(new_Jinkela_wire_3796)
    );

    bfr new_Jinkela_buffer_2844 (
        .din(new_Jinkela_wire_3905),
        .dout(new_Jinkela_wire_3906)
    );

    bfr new_Jinkela_buffer_2753 (
        .din(new_Jinkela_wire_3796),
        .dout(new_Jinkela_wire_3797)
    );

    bfr new_Jinkela_buffer_2806 (
        .din(new_Jinkela_wire_3855),
        .dout(new_Jinkela_wire_3856)
    );

    bfr new_Jinkela_buffer_2754 (
        .din(new_Jinkela_wire_3797),
        .dout(new_Jinkela_wire_3798)
    );

    bfr new_Jinkela_buffer_2895 (
        .din(new_Jinkela_wire_3966),
        .dout(new_Jinkela_wire_3967)
    );

    bfr new_Jinkela_buffer_2755 (
        .din(new_Jinkela_wire_3798),
        .dout(new_Jinkela_wire_3799)
    );

    bfr new_Jinkela_buffer_2807 (
        .din(new_Jinkela_wire_3856),
        .dout(new_Jinkela_wire_3857)
    );

    bfr new_Jinkela_buffer_2756 (
        .din(new_Jinkela_wire_3799),
        .dout(new_Jinkela_wire_3800)
    );

    bfr new_Jinkela_buffer_2845 (
        .din(new_Jinkela_wire_3906),
        .dout(new_Jinkela_wire_3907)
    );

    bfr new_Jinkela_buffer_2757 (
        .din(new_Jinkela_wire_3800),
        .dout(new_Jinkela_wire_3801)
    );

    bfr new_Jinkela_buffer_2808 (
        .din(new_Jinkela_wire_3857),
        .dout(new_Jinkela_wire_3858)
    );

    bfr new_Jinkela_buffer_2758 (
        .din(new_Jinkela_wire_3801),
        .dout(new_Jinkela_wire_3802)
    );

    bfr new_Jinkela_buffer_2759 (
        .din(new_Jinkela_wire_3802),
        .dout(new_Jinkela_wire_3803)
    );

    bfr new_Jinkela_buffer_2809 (
        .din(new_Jinkela_wire_3858),
        .dout(new_Jinkela_wire_3859)
    );

    bfr new_Jinkela_buffer_2760 (
        .din(new_Jinkela_wire_3803),
        .dout(new_Jinkela_wire_3804)
    );

    bfr new_Jinkela_buffer_2846 (
        .din(new_Jinkela_wire_3907),
        .dout(new_Jinkela_wire_3908)
    );

    bfr new_Jinkela_buffer_2761 (
        .din(new_Jinkela_wire_3804),
        .dout(new_Jinkela_wire_3805)
    );

    bfr new_Jinkela_buffer_2810 (
        .din(new_Jinkela_wire_3859),
        .dout(new_Jinkela_wire_3860)
    );

    bfr new_Jinkela_buffer_2762 (
        .din(new_Jinkela_wire_3805),
        .dout(new_Jinkela_wire_3806)
    );

    bfr new_Jinkela_buffer_2896 (
        .din(new_Jinkela_wire_3967),
        .dout(new_Jinkela_wire_3968)
    );

    bfr new_Jinkela_buffer_2763 (
        .din(new_Jinkela_wire_3806),
        .dout(new_Jinkela_wire_3807)
    );

    bfr new_Jinkela_buffer_2811 (
        .din(new_Jinkela_wire_3860),
        .dout(new_Jinkela_wire_3861)
    );

    bfr new_Jinkela_buffer_2764 (
        .din(new_Jinkela_wire_3807),
        .dout(new_Jinkela_wire_3808)
    );

    bfr new_Jinkela_buffer_2847 (
        .din(new_Jinkela_wire_3908),
        .dout(new_Jinkela_wire_3909)
    );

    bfr new_Jinkela_buffer_2765 (
        .din(new_Jinkela_wire_3808),
        .dout(new_Jinkela_wire_3809)
    );

    bfr new_Jinkela_buffer_2812 (
        .din(new_Jinkela_wire_3861),
        .dout(new_Jinkela_wire_3862)
    );

    bfr new_Jinkela_buffer_2766 (
        .din(new_Jinkela_wire_3809),
        .dout(new_Jinkela_wire_3810)
    );

    spl2 new_Jinkela_splitter_388 (
        .a(_1396_),
        .b(new_Jinkela_wire_4080),
        .c(new_Jinkela_wire_4081)
    );

    bfr new_Jinkela_buffer_2767 (
        .din(new_Jinkela_wire_3810),
        .dout(new_Jinkela_wire_3811)
    );

    bfr new_Jinkela_buffer_2813 (
        .din(new_Jinkela_wire_3862),
        .dout(new_Jinkela_wire_3863)
    );

    spl2 new_Jinkela_splitter_371 (
        .a(new_Jinkela_wire_3811),
        .b(new_Jinkela_wire_3812),
        .c(new_Jinkela_wire_3813)
    );

    bfr new_Jinkela_buffer_2814 (
        .din(new_Jinkela_wire_3863),
        .dout(new_Jinkela_wire_3864)
    );

    bfr new_Jinkela_buffer_2848 (
        .din(new_Jinkela_wire_3909),
        .dout(new_Jinkela_wire_3910)
    );

    bfr new_Jinkela_buffer_2897 (
        .din(new_Jinkela_wire_3968),
        .dout(new_Jinkela_wire_3969)
    );

    bfr new_Jinkela_buffer_2815 (
        .din(new_Jinkela_wire_3864),
        .dout(new_Jinkela_wire_3865)
    );

    bfr new_Jinkela_buffer_2849 (
        .din(new_Jinkela_wire_3910),
        .dout(new_Jinkela_wire_3911)
    );

    bfr new_Jinkela_buffer_2816 (
        .din(new_Jinkela_wire_3865),
        .dout(new_Jinkela_wire_3866)
    );

    bfr new_Jinkela_buffer_2998 (
        .din(new_Jinkela_wire_4075),
        .dout(new_Jinkela_wire_4076)
    );

    bfr new_Jinkela_buffer_3002 (
        .din(_1173_),
        .dout(new_Jinkela_wire_4082)
    );

    bfr new_Jinkela_buffer_2817 (
        .din(new_Jinkela_wire_3866),
        .dout(new_Jinkela_wire_3867)
    );

    and_bb _3592_ (
        .a(new_Jinkela_wire_6522),
        .b(new_Jinkela_wire_17635),
        .c(_0892_)
    );

    or_bb _3593_ (
        .a(new_Jinkela_wire_15682),
        .b(new_Jinkela_wire_854),
        .c(_0894_)
    );

    and_ii _3594_ (
        .a(new_Jinkela_wire_6992),
        .b(new_Jinkela_wire_9693),
        .c(_0895_)
    );

    and_bb _3595_ (
        .a(new_Jinkela_wire_6993),
        .b(new_Jinkela_wire_9694),
        .c(_0896_)
    );

    or_bb _3596_ (
        .a(new_Jinkela_wire_6367),
        .b(new_Jinkela_wire_10073),
        .c(_0897_)
    );

    and_ii _3597_ (
        .a(new_Jinkela_wire_11432),
        .b(new_Jinkela_wire_5689),
        .c(_0898_)
    );

    and_bb _3598_ (
        .a(new_Jinkela_wire_11433),
        .b(new_Jinkela_wire_5690),
        .c(_0899_)
    );

    or_bb _3599_ (
        .a(new_Jinkela_wire_14078),
        .b(new_Jinkela_wire_19911),
        .c(_0900_)
    );

    and_ii _3600_ (
        .a(new_Jinkela_wire_3964),
        .b(new_Jinkela_wire_7968),
        .c(_0901_)
    );

    and_bb _3601_ (
        .a(new_Jinkela_wire_3965),
        .b(new_Jinkela_wire_7969),
        .c(_0902_)
    );

    or_bb _3602_ (
        .a(new_Jinkela_wire_4719),
        .b(new_Jinkela_wire_4245),
        .c(_0903_)
    );

    and_ii _3603_ (
        .a(new_Jinkela_wire_21153),
        .b(new_Jinkela_wire_3120),
        .c(_0905_)
    );

    and_bb _3604_ (
        .a(new_Jinkela_wire_21154),
        .b(new_Jinkela_wire_3121),
        .c(_0906_)
    );

    or_bb _3605_ (
        .a(new_Jinkela_wire_18222),
        .b(new_Jinkela_wire_19290),
        .c(_0907_)
    );

    and_ii _3606_ (
        .a(new_Jinkela_wire_4897),
        .b(new_Jinkela_wire_11338),
        .c(_0908_)
    );

    and_bb _3607_ (
        .a(new_Jinkela_wire_4898),
        .b(new_Jinkela_wire_11339),
        .c(_0909_)
    );

    or_bb _3608_ (
        .a(new_Jinkela_wire_5434),
        .b(new_Jinkela_wire_6370),
        .c(_0910_)
    );

    and_ii _3609_ (
        .a(new_Jinkela_wire_15674),
        .b(new_Jinkela_wire_1771),
        .c(_0911_)
    );

    and_bb _3610_ (
        .a(new_Jinkela_wire_15675),
        .b(new_Jinkela_wire_1772),
        .c(_0912_)
    );

    or_bb _3611_ (
        .a(new_Jinkela_wire_7972),
        .b(new_Jinkela_wire_19128),
        .c(_0913_)
    );

    and_ii _3612_ (
        .a(new_Jinkela_wire_16945),
        .b(new_Jinkela_wire_20512),
        .c(_0914_)
    );

    and_bb _3613_ (
        .a(new_Jinkela_wire_16946),
        .b(new_Jinkela_wire_20513),
        .c(_0916_)
    );

    or_bb _3614_ (
        .a(new_Jinkela_wire_21183),
        .b(new_Jinkela_wire_19558),
        .c(_0917_)
    );

    and_ii _3615_ (
        .a(new_Jinkela_wire_4473),
        .b(new_Jinkela_wire_17069),
        .c(_0918_)
    );

    and_bb _3616_ (
        .a(new_Jinkela_wire_4474),
        .b(new_Jinkela_wire_17070),
        .c(_0919_)
    );

    and_ii _3617_ (
        .a(new_Jinkela_wire_7719),
        .b(new_Jinkela_wire_10399),
        .c(_0920_)
    );

    and_bb _3618_ (
        .a(new_Jinkela_wire_13193),
        .b(new_Jinkela_wire_3437),
        .c(_0921_)
    );

    and_ii _3619_ (
        .a(new_Jinkela_wire_13194),
        .b(new_Jinkela_wire_3438),
        .c(_0922_)
    );

    or_bb _3620_ (
        .a(new_Jinkela_wire_15671),
        .b(new_Jinkela_wire_3711),
        .c(new_net_3924)
    );

    or_bb _3621_ (
        .a(new_Jinkela_wire_3712),
        .b(new_Jinkela_wire_10440),
        .c(_0923_)
    );

    and_ii _3622_ (
        .a(new_Jinkela_wire_19559),
        .b(new_Jinkela_wire_19133),
        .c(_0924_)
    );

    and_bb _3623_ (
        .a(new_Jinkela_wire_400),
        .b(new_Jinkela_wire_680),
        .c(_0926_)
    );

    and_ii _3624_ (
        .a(new_Jinkela_wire_6371),
        .b(new_Jinkela_wire_19295),
        .c(_0927_)
    );

    and_bb _3625_ (
        .a(new_Jinkela_wire_158),
        .b(new_Jinkela_wire_518),
        .c(_0928_)
    );

    and_ii _3626_ (
        .a(new_Jinkela_wire_4246),
        .b(new_Jinkela_wire_19916),
        .c(_0929_)
    );

    and_bb _3627_ (
        .a(new_Jinkela_wire_601),
        .b(new_Jinkela_wire_133),
        .c(_0930_)
    );

    and_bb _3628_ (
        .a(new_Jinkela_wire_425),
        .b(new_Jinkela_wire_202),
        .c(_0931_)
    );

    and_ii _3629_ (
        .a(new_Jinkela_wire_10074),
        .b(new_Jinkela_wire_859),
        .c(_0932_)
    );

    and_ii _3630_ (
        .a(new_Jinkela_wire_12067),
        .b(new_Jinkela_wire_11134),
        .c(_0933_)
    );

    and_bb _3631_ (
        .a(new_Jinkela_wire_12068),
        .b(new_Jinkela_wire_11135),
        .c(_0934_)
    );

    or_bb _3632_ (
        .a(new_Jinkela_wire_14212),
        .b(new_Jinkela_wire_18944),
        .c(_0935_)
    );

    and_ii _3633_ (
        .a(new_Jinkela_wire_17532),
        .b(new_Jinkela_wire_3812),
        .c(_0937_)
    );

    bfr new_Jinkela_buffer_9679 (
        .din(new_Jinkela_wire_11778),
        .dout(new_Jinkela_wire_11779)
    );

    bfr new_Jinkela_buffer_9680 (
        .din(new_Jinkela_wire_11779),
        .dout(new_Jinkela_wire_11780)
    );

    bfr new_Jinkela_buffer_9751 (
        .din(new_Jinkela_wire_11860),
        .dout(new_Jinkela_wire_11861)
    );

    bfr new_Jinkela_buffer_9681 (
        .din(new_Jinkela_wire_11780),
        .dout(new_Jinkela_wire_11781)
    );

    bfr new_Jinkela_buffer_9851 (
        .din(new_Jinkela_wire_11970),
        .dout(new_Jinkela_wire_11971)
    );

    bfr new_Jinkela_buffer_9682 (
        .din(new_Jinkela_wire_11781),
        .dout(new_Jinkela_wire_11782)
    );

    bfr new_Jinkela_buffer_9752 (
        .din(new_Jinkela_wire_11861),
        .dout(new_Jinkela_wire_11862)
    );

    bfr new_Jinkela_buffer_9683 (
        .din(new_Jinkela_wire_11782),
        .dout(new_Jinkela_wire_11783)
    );

    bfr new_Jinkela_buffer_9926 (
        .din(new_Jinkela_wire_12049),
        .dout(new_Jinkela_wire_12050)
    );

    bfr new_Jinkela_buffer_9684 (
        .din(new_Jinkela_wire_11783),
        .dout(new_Jinkela_wire_11784)
    );

    bfr new_Jinkela_buffer_9753 (
        .din(new_Jinkela_wire_11862),
        .dout(new_Jinkela_wire_11863)
    );

    bfr new_Jinkela_buffer_9685 (
        .din(new_Jinkela_wire_11784),
        .dout(new_Jinkela_wire_11785)
    );

    bfr new_Jinkela_buffer_9852 (
        .din(new_Jinkela_wire_11971),
        .dout(new_Jinkela_wire_11972)
    );

    bfr new_Jinkela_buffer_9686 (
        .din(new_Jinkela_wire_11785),
        .dout(new_Jinkela_wire_11786)
    );

    bfr new_Jinkela_buffer_9754 (
        .din(new_Jinkela_wire_11863),
        .dout(new_Jinkela_wire_11864)
    );

    bfr new_Jinkela_buffer_9687 (
        .din(new_Jinkela_wire_11786),
        .dout(new_Jinkela_wire_11787)
    );

    spl2 new_Jinkela_splitter_914 (
        .a(_0664_),
        .b(new_Jinkela_wire_12058),
        .c(new_Jinkela_wire_12059)
    );

    bfr new_Jinkela_buffer_9688 (
        .din(new_Jinkela_wire_11787),
        .dout(new_Jinkela_wire_11788)
    );

    bfr new_Jinkela_buffer_9755 (
        .din(new_Jinkela_wire_11864),
        .dout(new_Jinkela_wire_11865)
    );

    bfr new_Jinkela_buffer_9689 (
        .din(new_Jinkela_wire_11788),
        .dout(new_Jinkela_wire_11789)
    );

    bfr new_Jinkela_buffer_9853 (
        .din(new_Jinkela_wire_11972),
        .dout(new_Jinkela_wire_11973)
    );

    bfr new_Jinkela_buffer_9690 (
        .din(new_Jinkela_wire_11789),
        .dout(new_Jinkela_wire_11790)
    );

    bfr new_Jinkela_buffer_9756 (
        .din(new_Jinkela_wire_11865),
        .dout(new_Jinkela_wire_11866)
    );

    bfr new_Jinkela_buffer_9691 (
        .din(new_Jinkela_wire_11790),
        .dout(new_Jinkela_wire_11791)
    );

    spl2 new_Jinkela_splitter_915 (
        .a(_0599_),
        .b(new_Jinkela_wire_12060),
        .c(new_Jinkela_wire_12061)
    );

    bfr new_Jinkela_buffer_9692 (
        .din(new_Jinkela_wire_11791),
        .dout(new_Jinkela_wire_11792)
    );

    bfr new_Jinkela_buffer_9757 (
        .din(new_Jinkela_wire_11866),
        .dout(new_Jinkela_wire_11867)
    );

    bfr new_Jinkela_buffer_9693 (
        .din(new_Jinkela_wire_11792),
        .dout(new_Jinkela_wire_11793)
    );

    bfr new_Jinkela_buffer_9854 (
        .din(new_Jinkela_wire_11973),
        .dout(new_Jinkela_wire_11974)
    );

    bfr new_Jinkela_buffer_9694 (
        .din(new_Jinkela_wire_11793),
        .dout(new_Jinkela_wire_11794)
    );

    bfr new_Jinkela_buffer_9758 (
        .din(new_Jinkela_wire_11867),
        .dout(new_Jinkela_wire_11868)
    );

    bfr new_Jinkela_buffer_9695 (
        .din(new_Jinkela_wire_11794),
        .dout(new_Jinkela_wire_11795)
    );

    bfr new_Jinkela_buffer_9928 (
        .din(_0244_),
        .dout(new_Jinkela_wire_12062)
    );

    bfr new_Jinkela_buffer_9696 (
        .din(new_Jinkela_wire_11795),
        .dout(new_Jinkela_wire_11796)
    );

    bfr new_Jinkela_buffer_9759 (
        .din(new_Jinkela_wire_11868),
        .dout(new_Jinkela_wire_11869)
    );

    bfr new_Jinkela_buffer_9697 (
        .din(new_Jinkela_wire_11796),
        .dout(new_Jinkela_wire_11797)
    );

    bfr new_Jinkela_buffer_9855 (
        .din(new_Jinkela_wire_11974),
        .dout(new_Jinkela_wire_11975)
    );

    bfr new_Jinkela_buffer_9698 (
        .din(new_Jinkela_wire_11797),
        .dout(new_Jinkela_wire_11798)
    );

    bfr new_Jinkela_buffer_9760 (
        .din(new_Jinkela_wire_11869),
        .dout(new_Jinkela_wire_11870)
    );

    bfr new_Jinkela_buffer_9699 (
        .din(new_Jinkela_wire_11798),
        .dout(new_Jinkela_wire_11799)
    );

    spl2 new_Jinkela_splitter_917 (
        .a(_0222_),
        .b(new_Jinkela_wire_12065),
        .c(new_Jinkela_wire_12066)
    );

    spl2 new_Jinkela_splitter_916 (
        .a(_0677_),
        .b(new_Jinkela_wire_12063),
        .c(new_Jinkela_wire_12064)
    );

    bfr new_Jinkela_buffer_16579 (
        .din(new_Jinkela_wire_19777),
        .dout(new_Jinkela_wire_19778)
    );

    bfr new_Jinkela_buffer_16600 (
        .din(new_Jinkela_wire_19808),
        .dout(new_Jinkela_wire_19809)
    );

    bfr new_Jinkela_buffer_16580 (
        .din(new_Jinkela_wire_19778),
        .dout(new_Jinkela_wire_19779)
    );

    bfr new_Jinkela_buffer_16706 (
        .din(new_Jinkela_wire_19922),
        .dout(new_Jinkela_wire_19923)
    );

    bfr new_Jinkela_buffer_16581 (
        .din(new_Jinkela_wire_19779),
        .dout(new_Jinkela_wire_19780)
    );

    bfr new_Jinkela_buffer_16601 (
        .din(new_Jinkela_wire_19809),
        .dout(new_Jinkela_wire_19810)
    );

    spl2 new_Jinkela_splitter_1448 (
        .a(new_Jinkela_wire_19780),
        .b(new_Jinkela_wire_19781),
        .c(new_Jinkela_wire_19782)
    );

    bfr new_Jinkela_buffer_16602 (
        .din(new_Jinkela_wire_19810),
        .dout(new_Jinkela_wire_19811)
    );

    bfr new_Jinkela_buffer_16709 (
        .din(_0241_),
        .dout(new_Jinkela_wire_19934)
    );

    bfr new_Jinkela_buffer_16707 (
        .din(new_Jinkela_wire_19923),
        .dout(new_Jinkela_wire_19924)
    );

    bfr new_Jinkela_buffer_16603 (
        .din(new_Jinkela_wire_19811),
        .dout(new_Jinkela_wire_19812)
    );

    spl2 new_Jinkela_splitter_1463 (
        .a(_0651_),
        .b(new_Jinkela_wire_19962),
        .c(new_Jinkela_wire_19963)
    );

    spl2 new_Jinkela_splitter_1458 (
        .a(new_Jinkela_wire_19927),
        .b(new_Jinkela_wire_19928),
        .c(new_Jinkela_wire_19929)
    );

    bfr new_Jinkela_buffer_16604 (
        .din(new_Jinkela_wire_19812),
        .dout(new_Jinkela_wire_19813)
    );

    spl2 new_Jinkela_splitter_1462 (
        .a(_1787_),
        .b(new_Jinkela_wire_19960),
        .c(new_Jinkela_wire_19961)
    );

    bfr new_Jinkela_buffer_16605 (
        .din(new_Jinkela_wire_19813),
        .dout(new_Jinkela_wire_19814)
    );

    bfr new_Jinkela_buffer_16710 (
        .din(new_Jinkela_wire_19934),
        .dout(new_Jinkela_wire_19935)
    );

    bfr new_Jinkela_buffer_16606 (
        .din(new_Jinkela_wire_19814),
        .dout(new_Jinkela_wire_19815)
    );

    bfr new_Jinkela_buffer_16607 (
        .din(new_Jinkela_wire_19815),
        .dout(new_Jinkela_wire_19816)
    );

    bfr new_Jinkela_buffer_16608 (
        .din(new_Jinkela_wire_19816),
        .dout(new_Jinkela_wire_19817)
    );

    bfr new_Jinkela_buffer_16711 (
        .din(new_Jinkela_wire_19935),
        .dout(new_Jinkela_wire_19936)
    );

    bfr new_Jinkela_buffer_16609 (
        .din(new_Jinkela_wire_19817),
        .dout(new_Jinkela_wire_19818)
    );

    spl2 new_Jinkela_splitter_1464 (
        .a(_0371_),
        .b(new_Jinkela_wire_19964),
        .c(new_Jinkela_wire_19965)
    );

    bfr new_Jinkela_buffer_16610 (
        .din(new_Jinkela_wire_19818),
        .dout(new_Jinkela_wire_19819)
    );

    bfr new_Jinkela_buffer_16712 (
        .din(new_Jinkela_wire_19936),
        .dout(new_Jinkela_wire_19937)
    );

    bfr new_Jinkela_buffer_16611 (
        .din(new_Jinkela_wire_19819),
        .dout(new_Jinkela_wire_19820)
    );

    spl2 new_Jinkela_splitter_1465 (
        .a(_1029_),
        .b(new_Jinkela_wire_19970),
        .c(new_Jinkela_wire_19971)
    );

    bfr new_Jinkela_buffer_16612 (
        .din(new_Jinkela_wire_19820),
        .dout(new_Jinkela_wire_19821)
    );

    bfr new_Jinkela_buffer_16713 (
        .din(new_Jinkela_wire_19937),
        .dout(new_Jinkela_wire_19938)
    );

    bfr new_Jinkela_buffer_16613 (
        .din(new_Jinkela_wire_19821),
        .dout(new_Jinkela_wire_19822)
    );

    bfr new_Jinkela_buffer_16733 (
        .din(new_Jinkela_wire_19965),
        .dout(new_Jinkela_wire_19966)
    );

    spl2 new_Jinkela_splitter_1466 (
        .a(_0315_),
        .b(new_Jinkela_wire_19972),
        .c(new_Jinkela_wire_19973)
    );

    bfr new_Jinkela_buffer_16614 (
        .din(new_Jinkela_wire_19822),
        .dout(new_Jinkela_wire_19823)
    );

    bfr new_Jinkela_buffer_16714 (
        .din(new_Jinkela_wire_19938),
        .dout(new_Jinkela_wire_19939)
    );

    bfr new_Jinkela_buffer_16615 (
        .din(new_Jinkela_wire_19823),
        .dout(new_Jinkela_wire_19824)
    );

    bfr new_Jinkela_buffer_16737 (
        .din(_1092_),
        .dout(new_Jinkela_wire_19974)
    );

    bfr new_Jinkela_buffer_16616 (
        .din(new_Jinkela_wire_19824),
        .dout(new_Jinkela_wire_19825)
    );

    bfr new_Jinkela_buffer_16715 (
        .din(new_Jinkela_wire_19939),
        .dout(new_Jinkela_wire_19940)
    );

    bfr new_Jinkela_buffer_16617 (
        .din(new_Jinkela_wire_19825),
        .dout(new_Jinkela_wire_19826)
    );

    bfr new_Jinkela_buffer_16734 (
        .din(new_Jinkela_wire_19966),
        .dout(new_Jinkela_wire_19967)
    );

    bfr new_Jinkela_buffer_16716 (
        .din(new_Jinkela_wire_19940),
        .dout(new_Jinkela_wire_19941)
    );

    bfr new_Jinkela_buffer_16618 (
        .din(new_Jinkela_wire_19826),
        .dout(new_Jinkela_wire_19827)
    );

    bfr new_Jinkela_buffer_2850 (
        .din(new_Jinkela_wire_3911),
        .dout(new_Jinkela_wire_3912)
    );

    bfr new_Jinkela_buffer_6224 (
        .din(new_Jinkela_wire_7897),
        .dout(new_Jinkela_wire_7898)
    );

    bfr new_Jinkela_buffer_2818 (
        .din(new_Jinkela_wire_3867),
        .dout(new_Jinkela_wire_3868)
    );

    bfr new_Jinkela_buffer_6485 (
        .din(_1012_),
        .dout(new_Jinkela_wire_8185)
    );

    bfr new_Jinkela_buffer_6354 (
        .din(new_Jinkela_wire_8041),
        .dout(new_Jinkela_wire_8042)
    );

    bfr new_Jinkela_buffer_2898 (
        .din(new_Jinkela_wire_3969),
        .dout(new_Jinkela_wire_3970)
    );

    bfr new_Jinkela_buffer_6225 (
        .din(new_Jinkela_wire_7898),
        .dout(new_Jinkela_wire_7899)
    );

    bfr new_Jinkela_buffer_2819 (
        .din(new_Jinkela_wire_3868),
        .dout(new_Jinkela_wire_3869)
    );

    bfr new_Jinkela_buffer_6310 (
        .din(new_Jinkela_wire_7989),
        .dout(new_Jinkela_wire_7990)
    );

    bfr new_Jinkela_buffer_2851 (
        .din(new_Jinkela_wire_3912),
        .dout(new_Jinkela_wire_3913)
    );

    bfr new_Jinkela_buffer_6226 (
        .din(new_Jinkela_wire_7899),
        .dout(new_Jinkela_wire_7900)
    );

    bfr new_Jinkela_buffer_2820 (
        .din(new_Jinkela_wire_3869),
        .dout(new_Jinkela_wire_3870)
    );

    bfr new_Jinkela_buffer_6339 (
        .din(new_Jinkela_wire_8022),
        .dout(new_Jinkela_wire_8023)
    );

    bfr new_Jinkela_buffer_3003 (
        .din(_1280_),
        .dout(new_Jinkela_wire_4085)
    );

    bfr new_Jinkela_buffer_6227 (
        .din(new_Jinkela_wire_7900),
        .dout(new_Jinkela_wire_7901)
    );

    bfr new_Jinkela_buffer_2821 (
        .din(new_Jinkela_wire_3870),
        .dout(new_Jinkela_wire_3871)
    );

    bfr new_Jinkela_buffer_6311 (
        .din(new_Jinkela_wire_7990),
        .dout(new_Jinkela_wire_7991)
    );

    bfr new_Jinkela_buffer_2852 (
        .din(new_Jinkela_wire_3913),
        .dout(new_Jinkela_wire_3914)
    );

    bfr new_Jinkela_buffer_6228 (
        .din(new_Jinkela_wire_7901),
        .dout(new_Jinkela_wire_7902)
    );

    bfr new_Jinkela_buffer_2822 (
        .din(new_Jinkela_wire_3871),
        .dout(new_Jinkela_wire_3872)
    );

    spl2 new_Jinkela_splitter_698 (
        .a(_0630_),
        .b(new_Jinkela_wire_8183),
        .c(new_Jinkela_wire_8184)
    );

    bfr new_Jinkela_buffer_6486 (
        .din(_1409_),
        .dout(new_Jinkela_wire_8186)
    );

    bfr new_Jinkela_buffer_2899 (
        .din(new_Jinkela_wire_3970),
        .dout(new_Jinkela_wire_3971)
    );

    bfr new_Jinkela_buffer_6229 (
        .din(new_Jinkela_wire_7902),
        .dout(new_Jinkela_wire_7903)
    );

    bfr new_Jinkela_buffer_2823 (
        .din(new_Jinkela_wire_3872),
        .dout(new_Jinkela_wire_3873)
    );

    bfr new_Jinkela_buffer_6312 (
        .din(new_Jinkela_wire_7991),
        .dout(new_Jinkela_wire_7992)
    );

    bfr new_Jinkela_buffer_2853 (
        .din(new_Jinkela_wire_3914),
        .dout(new_Jinkela_wire_3915)
    );

    bfr new_Jinkela_buffer_6230 (
        .din(new_Jinkela_wire_7903),
        .dout(new_Jinkela_wire_7904)
    );

    bfr new_Jinkela_buffer_2824 (
        .din(new_Jinkela_wire_3873),
        .dout(new_Jinkela_wire_3874)
    );

    bfr new_Jinkela_buffer_6340 (
        .din(new_Jinkela_wire_8023),
        .dout(new_Jinkela_wire_8024)
    );

    bfr new_Jinkela_buffer_2999 (
        .din(new_Jinkela_wire_4076),
        .dout(new_Jinkela_wire_4077)
    );

    bfr new_Jinkela_buffer_6231 (
        .din(new_Jinkela_wire_7904),
        .dout(new_Jinkela_wire_7905)
    );

    bfr new_Jinkela_buffer_2825 (
        .din(new_Jinkela_wire_3874),
        .dout(new_Jinkela_wire_3875)
    );

    bfr new_Jinkela_buffer_6313 (
        .din(new_Jinkela_wire_7992),
        .dout(new_Jinkela_wire_7993)
    );

    bfr new_Jinkela_buffer_2854 (
        .din(new_Jinkela_wire_3915),
        .dout(new_Jinkela_wire_3916)
    );

    bfr new_Jinkela_buffer_6232 (
        .din(new_Jinkela_wire_7905),
        .dout(new_Jinkela_wire_7906)
    );

    bfr new_Jinkela_buffer_2826 (
        .din(new_Jinkela_wire_3875),
        .dout(new_Jinkela_wire_3876)
    );

    bfr new_Jinkela_buffer_6413 (
        .din(new_Jinkela_wire_8104),
        .dout(new_Jinkela_wire_8105)
    );

    bfr new_Jinkela_buffer_2900 (
        .din(new_Jinkela_wire_3971),
        .dout(new_Jinkela_wire_3972)
    );

    bfr new_Jinkela_buffer_6233 (
        .din(new_Jinkela_wire_7906),
        .dout(new_Jinkela_wire_7907)
    );

    spl2 new_Jinkela_splitter_374 (
        .a(new_Jinkela_wire_3876),
        .b(new_Jinkela_wire_3877),
        .c(new_Jinkela_wire_3878)
    );

    bfr new_Jinkela_buffer_6314 (
        .din(new_Jinkela_wire_7993),
        .dout(new_Jinkela_wire_7994)
    );

    bfr new_Jinkela_buffer_6234 (
        .din(new_Jinkela_wire_7907),
        .dout(new_Jinkela_wire_7908)
    );

    spl2 new_Jinkela_splitter_389 (
        .a(_1694_),
        .b(new_Jinkela_wire_4083),
        .c(new_Jinkela_wire_4084)
    );

    bfr new_Jinkela_buffer_2855 (
        .din(new_Jinkela_wire_3916),
        .dout(new_Jinkela_wire_3917)
    );

    bfr new_Jinkela_buffer_6355 (
        .din(new_Jinkela_wire_8042),
        .dout(new_Jinkela_wire_8043)
    );

    bfr new_Jinkela_buffer_2856 (
        .din(new_Jinkela_wire_3917),
        .dout(new_Jinkela_wire_3918)
    );

    bfr new_Jinkela_buffer_6235 (
        .din(new_Jinkela_wire_7908),
        .dout(new_Jinkela_wire_7909)
    );

    bfr new_Jinkela_buffer_2901 (
        .din(new_Jinkela_wire_3972),
        .dout(new_Jinkela_wire_3973)
    );

    bfr new_Jinkela_buffer_6315 (
        .din(new_Jinkela_wire_7994),
        .dout(new_Jinkela_wire_7995)
    );

    bfr new_Jinkela_buffer_2857 (
        .din(new_Jinkela_wire_3918),
        .dout(new_Jinkela_wire_3919)
    );

    bfr new_Jinkela_buffer_6236 (
        .din(new_Jinkela_wire_7909),
        .dout(new_Jinkela_wire_7910)
    );

    bfr new_Jinkela_buffer_3000 (
        .din(new_Jinkela_wire_4077),
        .dout(new_Jinkela_wire_4078)
    );

    bfr new_Jinkela_buffer_2858 (
        .din(new_Jinkela_wire_3919),
        .dout(new_Jinkela_wire_3920)
    );

    bfr new_Jinkela_buffer_6237 (
        .din(new_Jinkela_wire_7910),
        .dout(new_Jinkela_wire_7911)
    );

    bfr new_Jinkela_buffer_2902 (
        .din(new_Jinkela_wire_3973),
        .dout(new_Jinkela_wire_3974)
    );

    bfr new_Jinkela_buffer_6316 (
        .din(new_Jinkela_wire_7995),
        .dout(new_Jinkela_wire_7996)
    );

    bfr new_Jinkela_buffer_2859 (
        .din(new_Jinkela_wire_3920),
        .dout(new_Jinkela_wire_3921)
    );

    bfr new_Jinkela_buffer_6238 (
        .din(new_Jinkela_wire_7911),
        .dout(new_Jinkela_wire_7912)
    );

    spl2 new_Jinkela_splitter_393 (
        .a(_1422_),
        .b(new_Jinkela_wire_4164),
        .c(new_Jinkela_wire_4165)
    );

    bfr new_Jinkela_buffer_6356 (
        .din(new_Jinkela_wire_8043),
        .dout(new_Jinkela_wire_8044)
    );

    bfr new_Jinkela_buffer_2860 (
        .din(new_Jinkela_wire_3921),
        .dout(new_Jinkela_wire_3922)
    );

    bfr new_Jinkela_buffer_6239 (
        .din(new_Jinkela_wire_7912),
        .dout(new_Jinkela_wire_7913)
    );

    bfr new_Jinkela_buffer_2903 (
        .din(new_Jinkela_wire_3974),
        .dout(new_Jinkela_wire_3975)
    );

    bfr new_Jinkela_buffer_6317 (
        .din(new_Jinkela_wire_7996),
        .dout(new_Jinkela_wire_7997)
    );

    bfr new_Jinkela_buffer_2861 (
        .din(new_Jinkela_wire_3922),
        .dout(new_Jinkela_wire_3923)
    );

    bfr new_Jinkela_buffer_6240 (
        .din(new_Jinkela_wire_7913),
        .dout(new_Jinkela_wire_7914)
    );

    bfr new_Jinkela_buffer_3001 (
        .din(new_Jinkela_wire_4078),
        .dout(new_Jinkela_wire_4079)
    );

    bfr new_Jinkela_buffer_6414 (
        .din(new_Jinkela_wire_8105),
        .dout(new_Jinkela_wire_8106)
    );

    bfr new_Jinkela_buffer_2862 (
        .din(new_Jinkela_wire_3923),
        .dout(new_Jinkela_wire_3924)
    );

    bfr new_Jinkela_buffer_6241 (
        .din(new_Jinkela_wire_7914),
        .dout(new_Jinkela_wire_7915)
    );

    bfr new_Jinkela_buffer_2904 (
        .din(new_Jinkela_wire_3975),
        .dout(new_Jinkela_wire_3976)
    );

    bfr new_Jinkela_buffer_6318 (
        .din(new_Jinkela_wire_7997),
        .dout(new_Jinkela_wire_7998)
    );

    bfr new_Jinkela_buffer_2863 (
        .din(new_Jinkela_wire_3924),
        .dout(new_Jinkela_wire_3925)
    );

    bfr new_Jinkela_buffer_6242 (
        .din(new_Jinkela_wire_7915),
        .dout(new_Jinkela_wire_7916)
    );

    spl2 new_Jinkela_splitter_391 (
        .a(_0206_),
        .b(new_Jinkela_wire_4159),
        .c(new_Jinkela_wire_4160)
    );

    bfr new_Jinkela_buffer_6357 (
        .din(new_Jinkela_wire_8044),
        .dout(new_Jinkela_wire_8045)
    );

    bfr new_Jinkela_buffer_2864 (
        .din(new_Jinkela_wire_3925),
        .dout(new_Jinkela_wire_3926)
    );

    bfr new_Jinkela_buffer_6243 (
        .din(new_Jinkela_wire_7916),
        .dout(new_Jinkela_wire_7917)
    );

    bfr new_Jinkela_buffer_2905 (
        .din(new_Jinkela_wire_3976),
        .dout(new_Jinkela_wire_3977)
    );

    bfr new_Jinkela_buffer_6319 (
        .din(new_Jinkela_wire_7998),
        .dout(new_Jinkela_wire_7999)
    );

    bfr new_Jinkela_buffer_2865 (
        .din(new_Jinkela_wire_3926),
        .dout(new_Jinkela_wire_3927)
    );

    bfr new_Jinkela_buffer_6244 (
        .din(new_Jinkela_wire_7917),
        .dout(new_Jinkela_wire_7918)
    );

    bfr new_Jinkela_buffer_3004 (
        .din(new_Jinkela_wire_4085),
        .dout(new_Jinkela_wire_4086)
    );

    bfr new_Jinkela_buffer_9700 (
        .din(new_Jinkela_wire_11799),
        .dout(new_Jinkela_wire_11800)
    );

    bfr new_Jinkela_buffer_9761 (
        .din(new_Jinkela_wire_11870),
        .dout(new_Jinkela_wire_11871)
    );

    bfr new_Jinkela_buffer_9701 (
        .din(new_Jinkela_wire_11800),
        .dout(new_Jinkela_wire_11801)
    );

    bfr new_Jinkela_buffer_9856 (
        .din(new_Jinkela_wire_11975),
        .dout(new_Jinkela_wire_11976)
    );

    bfr new_Jinkela_buffer_9702 (
        .din(new_Jinkela_wire_11801),
        .dout(new_Jinkela_wire_11802)
    );

    bfr new_Jinkela_buffer_9762 (
        .din(new_Jinkela_wire_11871),
        .dout(new_Jinkela_wire_11872)
    );

    bfr new_Jinkela_buffer_9703 (
        .din(new_Jinkela_wire_11802),
        .dout(new_Jinkela_wire_11803)
    );

    bfr new_Jinkela_buffer_9704 (
        .din(new_Jinkela_wire_11803),
        .dout(new_Jinkela_wire_11804)
    );

    bfr new_Jinkela_buffer_9763 (
        .din(new_Jinkela_wire_11872),
        .dout(new_Jinkela_wire_11873)
    );

    bfr new_Jinkela_buffer_9705 (
        .din(new_Jinkela_wire_11804),
        .dout(new_Jinkela_wire_11805)
    );

    bfr new_Jinkela_buffer_9857 (
        .din(new_Jinkela_wire_11976),
        .dout(new_Jinkela_wire_11977)
    );

    bfr new_Jinkela_buffer_9706 (
        .din(new_Jinkela_wire_11805),
        .dout(new_Jinkela_wire_11806)
    );

    bfr new_Jinkela_buffer_9764 (
        .din(new_Jinkela_wire_11873),
        .dout(new_Jinkela_wire_11874)
    );

    bfr new_Jinkela_buffer_9707 (
        .din(new_Jinkela_wire_11806),
        .dout(new_Jinkela_wire_11807)
    );

    spl2 new_Jinkela_splitter_918 (
        .a(_0932_),
        .b(new_Jinkela_wire_12067),
        .c(new_Jinkela_wire_12068)
    );

    bfr new_Jinkela_buffer_9708 (
        .din(new_Jinkela_wire_11807),
        .dout(new_Jinkela_wire_11808)
    );

    bfr new_Jinkela_buffer_9765 (
        .din(new_Jinkela_wire_11874),
        .dout(new_Jinkela_wire_11875)
    );

    bfr new_Jinkela_buffer_9709 (
        .din(new_Jinkela_wire_11808),
        .dout(new_Jinkela_wire_11809)
    );

    bfr new_Jinkela_buffer_9858 (
        .din(new_Jinkela_wire_11977),
        .dout(new_Jinkela_wire_11978)
    );

    bfr new_Jinkela_buffer_9710 (
        .din(new_Jinkela_wire_11809),
        .dout(new_Jinkela_wire_11810)
    );

    bfr new_Jinkela_buffer_9766 (
        .din(new_Jinkela_wire_11875),
        .dout(new_Jinkela_wire_11876)
    );

    bfr new_Jinkela_buffer_9711 (
        .din(new_Jinkela_wire_11810),
        .dout(new_Jinkela_wire_11811)
    );

    spl2 new_Jinkela_splitter_921 (
        .a(_1606_),
        .b(new_Jinkela_wire_12105),
        .c(new_Jinkela_wire_12106)
    );

    bfr new_Jinkela_buffer_9929 (
        .din(_1580_),
        .dout(new_Jinkela_wire_12069)
    );

    bfr new_Jinkela_buffer_9712 (
        .din(new_Jinkela_wire_11811),
        .dout(new_Jinkela_wire_11812)
    );

    bfr new_Jinkela_buffer_9767 (
        .din(new_Jinkela_wire_11876),
        .dout(new_Jinkela_wire_11877)
    );

    bfr new_Jinkela_buffer_9713 (
        .din(new_Jinkela_wire_11812),
        .dout(new_Jinkela_wire_11813)
    );

    bfr new_Jinkela_buffer_9859 (
        .din(new_Jinkela_wire_11978),
        .dout(new_Jinkela_wire_11979)
    );

    bfr new_Jinkela_buffer_9714 (
        .din(new_Jinkela_wire_11813),
        .dout(new_Jinkela_wire_11814)
    );

    bfr new_Jinkela_buffer_9768 (
        .din(new_Jinkela_wire_11877),
        .dout(new_Jinkela_wire_11878)
    );

    bfr new_Jinkela_buffer_9715 (
        .din(new_Jinkela_wire_11814),
        .dout(new_Jinkela_wire_11815)
    );

    spl2 new_Jinkela_splitter_920 (
        .a(_0037_),
        .b(new_Jinkela_wire_12103),
        .c(new_Jinkela_wire_12104)
    );

    bfr new_Jinkela_buffer_9716 (
        .din(new_Jinkela_wire_11815),
        .dout(new_Jinkela_wire_11816)
    );

    bfr new_Jinkela_buffer_9769 (
        .din(new_Jinkela_wire_11878),
        .dout(new_Jinkela_wire_11879)
    );

    bfr new_Jinkela_buffer_9717 (
        .din(new_Jinkela_wire_11816),
        .dout(new_Jinkela_wire_11817)
    );

    bfr new_Jinkela_buffer_9860 (
        .din(new_Jinkela_wire_11979),
        .dout(new_Jinkela_wire_11980)
    );

    bfr new_Jinkela_buffer_9718 (
        .din(new_Jinkela_wire_11817),
        .dout(new_Jinkela_wire_11818)
    );

    bfr new_Jinkela_buffer_9770 (
        .din(new_Jinkela_wire_11879),
        .dout(new_Jinkela_wire_11880)
    );

    bfr new_Jinkela_buffer_9719 (
        .din(new_Jinkela_wire_11818),
        .dout(new_Jinkela_wire_11819)
    );

    bfr new_Jinkela_buffer_9930 (
        .din(new_Jinkela_wire_12069),
        .dout(new_Jinkela_wire_12070)
    );

    bfr new_Jinkela_buffer_9720 (
        .din(new_Jinkela_wire_11819),
        .dout(new_Jinkela_wire_11820)
    );

    bfr new_Jinkela_buffer_9771 (
        .din(new_Jinkela_wire_11880),
        .dout(new_Jinkela_wire_11881)
    );

    and_bb _3634_ (
        .a(new_Jinkela_wire_17533),
        .b(new_Jinkela_wire_3813),
        .c(_0938_)
    );

    or_bb _3635_ (
        .a(new_Jinkela_wire_18298),
        .b(new_Jinkela_wire_3483),
        .c(_0939_)
    );

    and_ii _3636_ (
        .a(new_Jinkela_wire_11044),
        .b(new_Jinkela_wire_2954),
        .c(_0940_)
    );

    and_bb _3637_ (
        .a(new_Jinkela_wire_11045),
        .b(new_Jinkela_wire_2955),
        .c(_0941_)
    );

    or_bb _3638_ (
        .a(new_Jinkela_wire_17991),
        .b(new_Jinkela_wire_6960),
        .c(_0942_)
    );

    and_ii _3639_ (
        .a(new_Jinkela_wire_3718),
        .b(new_Jinkela_wire_2589),
        .c(_0943_)
    );

    and_bb _3640_ (
        .a(new_Jinkela_wire_3719),
        .b(new_Jinkela_wire_2590),
        .c(_0944_)
    );

    or_bb _3641_ (
        .a(new_Jinkela_wire_5537),
        .b(new_Jinkela_wire_3182),
        .c(_0945_)
    );

    and_ii _3642_ (
        .a(new_Jinkela_wire_2322),
        .b(new_Jinkela_wire_5725),
        .c(_0946_)
    );

    and_bb _3643_ (
        .a(new_Jinkela_wire_2323),
        .b(new_Jinkela_wire_5726),
        .c(_0948_)
    );

    or_bb _3644_ (
        .a(new_Jinkela_wire_3721),
        .b(new_Jinkela_wire_18309),
        .c(_0949_)
    );

    and_ii _3645_ (
        .a(new_Jinkela_wire_14032),
        .b(new_Jinkela_wire_5280),
        .c(_0950_)
    );

    and_bb _3646_ (
        .a(new_Jinkela_wire_14033),
        .b(new_Jinkela_wire_5281),
        .c(_0951_)
    );

    or_bb _3647_ (
        .a(new_Jinkela_wire_2119),
        .b(new_Jinkela_wire_3245),
        .c(_0952_)
    );

    and_ii _3648_ (
        .a(new_Jinkela_wire_12329),
        .b(new_Jinkela_wire_19048),
        .c(_0953_)
    );

    and_bb _3649_ (
        .a(new_Jinkela_wire_12330),
        .b(new_Jinkela_wire_19049),
        .c(_0954_)
    );

    and_ii _3650_ (
        .a(new_Jinkela_wire_21105),
        .b(new_Jinkela_wire_19685),
        .c(_0955_)
    );

    and_bb _3651_ (
        .a(new_Jinkela_wire_9010),
        .b(new_Jinkela_wire_12056),
        .c(_0956_)
    );

    and_ii _3652_ (
        .a(new_Jinkela_wire_9011),
        .b(new_Jinkela_wire_12057),
        .c(_0957_)
    );

    or_bb _3653_ (
        .a(new_Jinkela_wire_7750),
        .b(new_Jinkela_wire_18805),
        .c(new_net_3948)
    );

    and_ii _3654_ (
        .a(new_Jinkela_wire_18806),
        .b(new_Jinkela_wire_19730),
        .c(_0959_)
    );

    and_ii _3655_ (
        .a(new_Jinkela_wire_3246),
        .b(new_Jinkela_wire_18314),
        .c(_0960_)
    );

    and_bb _3656_ (
        .a(new_Jinkela_wire_157),
        .b(new_Jinkela_wire_669),
        .c(_0961_)
    );

    and_ii _3657_ (
        .a(new_Jinkela_wire_3183),
        .b(new_Jinkela_wire_6965),
        .c(_0962_)
    );

    and_bb _3658_ (
        .a(new_Jinkela_wire_609),
        .b(new_Jinkela_wire_525),
        .c(_0963_)
    );

    and_bb _3659_ (
        .a(new_Jinkela_wire_420),
        .b(new_Jinkela_wire_137),
        .c(_0964_)
    );

    and_ii _3660_ (
        .a(new_Jinkela_wire_3484),
        .b(new_Jinkela_wire_18949),
        .c(_0965_)
    );

    and_ii _3661_ (
        .a(new_Jinkela_wire_12733),
        .b(new_Jinkela_wire_8578),
        .c(_0966_)
    );

    and_bb _3662_ (
        .a(new_Jinkela_wire_12734),
        .b(new_Jinkela_wire_8579),
        .c(_0967_)
    );

    or_bb _3663_ (
        .a(new_Jinkela_wire_14689),
        .b(new_Jinkela_wire_6848),
        .c(_0969_)
    );

    and_ii _3664_ (
        .a(new_Jinkela_wire_5685),
        .b(new_Jinkela_wire_7689),
        .c(_0970_)
    );

    and_bb _3665_ (
        .a(new_Jinkela_wire_5686),
        .b(new_Jinkela_wire_7690),
        .c(_0971_)
    );

    or_bb _3666_ (
        .a(new_Jinkela_wire_18572),
        .b(new_Jinkela_wire_21190),
        .c(_0972_)
    );

    and_ii _3667_ (
        .a(new_Jinkela_wire_1631),
        .b(new_Jinkela_wire_20263),
        .c(_0973_)
    );

    and_bb _3668_ (
        .a(new_Jinkela_wire_1632),
        .b(new_Jinkela_wire_20264),
        .c(_0974_)
    );

    or_bb _3669_ (
        .a(new_Jinkela_wire_19158),
        .b(new_Jinkela_wire_17536),
        .c(_0975_)
    );

    and_ii _3670_ (
        .a(new_Jinkela_wire_17673),
        .b(new_Jinkela_wire_9297),
        .c(_0976_)
    );

    and_bb _3671_ (
        .a(new_Jinkela_wire_17674),
        .b(new_Jinkela_wire_9298),
        .c(_0977_)
    );

    or_bb _3672_ (
        .a(new_Jinkela_wire_11399),
        .b(new_Jinkela_wire_721),
        .c(_0978_)
    );

    and_ii _3673_ (
        .a(new_Jinkela_wire_19124),
        .b(new_Jinkela_wire_10684),
        .c(_0980_)
    );

    and_bb _3674_ (
        .a(new_Jinkela_wire_19125),
        .b(new_Jinkela_wire_10685),
        .c(_0981_)
    );

    and_ii _3675_ (
        .a(new_Jinkela_wire_4669),
        .b(new_Jinkela_wire_17111),
        .c(_0982_)
    );

    bfr new_Jinkela_buffer_6245 (
        .din(new_Jinkela_wire_7918),
        .dout(new_Jinkela_wire_7919)
    );

    bfr new_Jinkela_buffer_13204 (
        .din(new_Jinkela_wire_15799),
        .dout(new_Jinkela_wire_15800)
    );

    bfr new_Jinkela_buffer_16619 (
        .din(new_Jinkela_wire_19827),
        .dout(new_Jinkela_wire_19828)
    );

    bfr new_Jinkela_buffer_6320 (
        .din(new_Jinkela_wire_7999),
        .dout(new_Jinkela_wire_8000)
    );

    bfr new_Jinkela_buffer_13297 (
        .din(new_Jinkela_wire_15896),
        .dout(new_Jinkela_wire_15897)
    );

    spl2 new_Jinkela_splitter_1468 (
        .a(_1651_),
        .b(new_Jinkela_wire_20039),
        .c(new_Jinkela_wire_20040)
    );

    bfr new_Jinkela_buffer_6246 (
        .din(new_Jinkela_wire_7919),
        .dout(new_Jinkela_wire_7920)
    );

    bfr new_Jinkela_buffer_13205 (
        .din(new_Jinkela_wire_15800),
        .dout(new_Jinkela_wire_15801)
    );

    bfr new_Jinkela_buffer_16620 (
        .din(new_Jinkela_wire_19828),
        .dout(new_Jinkela_wire_19829)
    );

    spl2 new_Jinkela_splitter_694 (
        .a(_0391_),
        .b(new_Jinkela_wire_8095),
        .c(new_Jinkela_wire_8096)
    );

    bfr new_Jinkela_buffer_13246 (
        .din(new_Jinkela_wire_15845),
        .dout(new_Jinkela_wire_15846)
    );

    bfr new_Jinkela_buffer_16717 (
        .din(new_Jinkela_wire_19941),
        .dout(new_Jinkela_wire_19942)
    );

    bfr new_Jinkela_buffer_6247 (
        .din(new_Jinkela_wire_7920),
        .dout(new_Jinkela_wire_7921)
    );

    bfr new_Jinkela_buffer_13206 (
        .din(new_Jinkela_wire_15801),
        .dout(new_Jinkela_wire_15802)
    );

    bfr new_Jinkela_buffer_16621 (
        .din(new_Jinkela_wire_19829),
        .dout(new_Jinkela_wire_19830)
    );

    bfr new_Jinkela_buffer_6321 (
        .din(new_Jinkela_wire_8000),
        .dout(new_Jinkela_wire_8001)
    );

    bfr new_Jinkela_buffer_16735 (
        .din(new_Jinkela_wire_19967),
        .dout(new_Jinkela_wire_19968)
    );

    bfr new_Jinkela_buffer_6248 (
        .din(new_Jinkela_wire_7921),
        .dout(new_Jinkela_wire_7922)
    );

    bfr new_Jinkela_buffer_13207 (
        .din(new_Jinkela_wire_15802),
        .dout(new_Jinkela_wire_15803)
    );

    bfr new_Jinkela_buffer_16622 (
        .din(new_Jinkela_wire_19830),
        .dout(new_Jinkela_wire_19831)
    );

    bfr new_Jinkela_buffer_6409 (
        .din(_0837_),
        .dout(new_Jinkela_wire_8101)
    );

    bfr new_Jinkela_buffer_13247 (
        .din(new_Jinkela_wire_15846),
        .dout(new_Jinkela_wire_15847)
    );

    bfr new_Jinkela_buffer_16718 (
        .din(new_Jinkela_wire_19942),
        .dout(new_Jinkela_wire_19943)
    );

    bfr new_Jinkela_buffer_6342 (
        .din(new_Jinkela_wire_8029),
        .dout(new_Jinkela_wire_8030)
    );

    bfr new_Jinkela_buffer_6249 (
        .din(new_Jinkela_wire_7922),
        .dout(new_Jinkela_wire_7923)
    );

    bfr new_Jinkela_buffer_13208 (
        .din(new_Jinkela_wire_15803),
        .dout(new_Jinkela_wire_15804)
    );

    bfr new_Jinkela_buffer_16623 (
        .din(new_Jinkela_wire_19831),
        .dout(new_Jinkela_wire_19832)
    );

    bfr new_Jinkela_buffer_6322 (
        .din(new_Jinkela_wire_8001),
        .dout(new_Jinkela_wire_8002)
    );

    bfr new_Jinkela_buffer_13298 (
        .din(new_Jinkela_wire_15897),
        .dout(new_Jinkela_wire_15898)
    );

    bfr new_Jinkela_buffer_16738 (
        .din(_0779_),
        .dout(new_Jinkela_wire_19975)
    );

    bfr new_Jinkela_buffer_6250 (
        .din(new_Jinkela_wire_7923),
        .dout(new_Jinkela_wire_7924)
    );

    bfr new_Jinkela_buffer_13209 (
        .din(new_Jinkela_wire_15804),
        .dout(new_Jinkela_wire_15805)
    );

    bfr new_Jinkela_buffer_16624 (
        .din(new_Jinkela_wire_19832),
        .dout(new_Jinkela_wire_19833)
    );

    bfr new_Jinkela_buffer_13248 (
        .din(new_Jinkela_wire_15847),
        .dout(new_Jinkela_wire_15848)
    );

    bfr new_Jinkela_buffer_16719 (
        .din(new_Jinkela_wire_19943),
        .dout(new_Jinkela_wire_19944)
    );

    bfr new_Jinkela_buffer_6251 (
        .din(new_Jinkela_wire_7924),
        .dout(new_Jinkela_wire_7925)
    );

    bfr new_Jinkela_buffer_13210 (
        .din(new_Jinkela_wire_15805),
        .dout(new_Jinkela_wire_15806)
    );

    bfr new_Jinkela_buffer_16625 (
        .din(new_Jinkela_wire_19833),
        .dout(new_Jinkela_wire_19834)
    );

    bfr new_Jinkela_buffer_6323 (
        .din(new_Jinkela_wire_8002),
        .dout(new_Jinkela_wire_8003)
    );

    bfr new_Jinkela_buffer_13312 (
        .din(new_Jinkela_wire_15913),
        .dout(new_Jinkela_wire_15914)
    );

    bfr new_Jinkela_buffer_16736 (
        .din(new_Jinkela_wire_19968),
        .dout(new_Jinkela_wire_19969)
    );

    bfr new_Jinkela_buffer_6252 (
        .din(new_Jinkela_wire_7925),
        .dout(new_Jinkela_wire_7926)
    );

    bfr new_Jinkela_buffer_13211 (
        .din(new_Jinkela_wire_15806),
        .dout(new_Jinkela_wire_15807)
    );

    bfr new_Jinkela_buffer_16626 (
        .din(new_Jinkela_wire_19834),
        .dout(new_Jinkela_wire_19835)
    );

    bfr new_Jinkela_buffer_13249 (
        .din(new_Jinkela_wire_15848),
        .dout(new_Jinkela_wire_15849)
    );

    bfr new_Jinkela_buffer_16720 (
        .din(new_Jinkela_wire_19944),
        .dout(new_Jinkela_wire_19945)
    );

    bfr new_Jinkela_buffer_6343 (
        .din(new_Jinkela_wire_8030),
        .dout(new_Jinkela_wire_8031)
    );

    bfr new_Jinkela_buffer_6253 (
        .din(new_Jinkela_wire_7926),
        .dout(new_Jinkela_wire_7927)
    );

    bfr new_Jinkela_buffer_13212 (
        .din(new_Jinkela_wire_15807),
        .dout(new_Jinkela_wire_15808)
    );

    bfr new_Jinkela_buffer_16627 (
        .din(new_Jinkela_wire_19835),
        .dout(new_Jinkela_wire_19836)
    );

    bfr new_Jinkela_buffer_6324 (
        .din(new_Jinkela_wire_8003),
        .dout(new_Jinkela_wire_8004)
    );

    bfr new_Jinkela_buffer_13299 (
        .din(new_Jinkela_wire_15898),
        .dout(new_Jinkela_wire_15899)
    );

    spl2 new_Jinkela_splitter_1469 (
        .a(_1298_),
        .b(new_Jinkela_wire_20041),
        .c(new_Jinkela_wire_20042)
    );

    bfr new_Jinkela_buffer_6254 (
        .din(new_Jinkela_wire_7927),
        .dout(new_Jinkela_wire_7928)
    );

    bfr new_Jinkela_buffer_13213 (
        .din(new_Jinkela_wire_15808),
        .dout(new_Jinkela_wire_15809)
    );

    bfr new_Jinkela_buffer_16628 (
        .din(new_Jinkela_wire_19836),
        .dout(new_Jinkela_wire_19837)
    );

    bfr new_Jinkela_buffer_13250 (
        .din(new_Jinkela_wire_15849),
        .dout(new_Jinkela_wire_15850)
    );

    bfr new_Jinkela_buffer_16721 (
        .din(new_Jinkela_wire_19945),
        .dout(new_Jinkela_wire_19946)
    );

    bfr new_Jinkela_buffer_6405 (
        .din(new_Jinkela_wire_8096),
        .dout(new_Jinkela_wire_8097)
    );

    bfr new_Jinkela_buffer_6255 (
        .din(new_Jinkela_wire_7928),
        .dout(new_Jinkela_wire_7929)
    );

    bfr new_Jinkela_buffer_13214 (
        .din(new_Jinkela_wire_15809),
        .dout(new_Jinkela_wire_15810)
    );

    bfr new_Jinkela_buffer_16629 (
        .din(new_Jinkela_wire_19837),
        .dout(new_Jinkela_wire_19838)
    );

    bfr new_Jinkela_buffer_6325 (
        .din(new_Jinkela_wire_8004),
        .dout(new_Jinkela_wire_8005)
    );

    bfr new_Jinkela_buffer_16739 (
        .din(new_Jinkela_wire_19975),
        .dout(new_Jinkela_wire_19976)
    );

    spl2 new_Jinkela_splitter_1153 (
        .a(_1249_),
        .b(new_Jinkela_wire_16002),
        .c(new_Jinkela_wire_16003)
    );

    bfr new_Jinkela_buffer_6256 (
        .din(new_Jinkela_wire_7929),
        .dout(new_Jinkela_wire_7930)
    );

    bfr new_Jinkela_buffer_13215 (
        .din(new_Jinkela_wire_15810),
        .dout(new_Jinkela_wire_15811)
    );

    bfr new_Jinkela_buffer_16630 (
        .din(new_Jinkela_wire_19838),
        .dout(new_Jinkela_wire_19839)
    );

    bfr new_Jinkela_buffer_6483 (
        .din(_0822_),
        .dout(new_Jinkela_wire_8177)
    );

    bfr new_Jinkela_buffer_13251 (
        .din(new_Jinkela_wire_15850),
        .dout(new_Jinkela_wire_15851)
    );

    bfr new_Jinkela_buffer_16722 (
        .din(new_Jinkela_wire_19946),
        .dout(new_Jinkela_wire_19947)
    );

    bfr new_Jinkela_buffer_6344 (
        .din(new_Jinkela_wire_8031),
        .dout(new_Jinkela_wire_8032)
    );

    bfr new_Jinkela_buffer_6257 (
        .din(new_Jinkela_wire_7930),
        .dout(new_Jinkela_wire_7931)
    );

    bfr new_Jinkela_buffer_13216 (
        .din(new_Jinkela_wire_15811),
        .dout(new_Jinkela_wire_15812)
    );

    bfr new_Jinkela_buffer_16631 (
        .din(new_Jinkela_wire_19839),
        .dout(new_Jinkela_wire_19840)
    );

    bfr new_Jinkela_buffer_6326 (
        .din(new_Jinkela_wire_8005),
        .dout(new_Jinkela_wire_8006)
    );

    bfr new_Jinkela_buffer_13300 (
        .din(new_Jinkela_wire_15899),
        .dout(new_Jinkela_wire_15900)
    );

    bfr new_Jinkela_buffer_6258 (
        .din(new_Jinkela_wire_7931),
        .dout(new_Jinkela_wire_7932)
    );

    bfr new_Jinkela_buffer_13217 (
        .din(new_Jinkela_wire_15812),
        .dout(new_Jinkela_wire_15813)
    );

    bfr new_Jinkela_buffer_16632 (
        .din(new_Jinkela_wire_19840),
        .dout(new_Jinkela_wire_19841)
    );

    bfr new_Jinkela_buffer_13252 (
        .din(new_Jinkela_wire_15851),
        .dout(new_Jinkela_wire_15852)
    );

    bfr new_Jinkela_buffer_16723 (
        .din(new_Jinkela_wire_19947),
        .dout(new_Jinkela_wire_19948)
    );

    bfr new_Jinkela_buffer_6259 (
        .din(new_Jinkela_wire_7932),
        .dout(new_Jinkela_wire_7933)
    );

    bfr new_Jinkela_buffer_13218 (
        .din(new_Jinkela_wire_15813),
        .dout(new_Jinkela_wire_15814)
    );

    bfr new_Jinkela_buffer_16633 (
        .din(new_Jinkela_wire_19841),
        .dout(new_Jinkela_wire_19842)
    );

    bfr new_Jinkela_buffer_6327 (
        .din(new_Jinkela_wire_8006),
        .dout(new_Jinkela_wire_8007)
    );

    bfr new_Jinkela_buffer_13313 (
        .din(new_Jinkela_wire_15914),
        .dout(new_Jinkela_wire_15915)
    );

    bfr new_Jinkela_buffer_16740 (
        .din(new_Jinkela_wire_19976),
        .dout(new_Jinkela_wire_19977)
    );

    bfr new_Jinkela_buffer_6260 (
        .din(new_Jinkela_wire_7933),
        .dout(new_Jinkela_wire_7934)
    );

    bfr new_Jinkela_buffer_13219 (
        .din(new_Jinkela_wire_15814),
        .dout(new_Jinkela_wire_15815)
    );

    bfr new_Jinkela_buffer_16634 (
        .din(new_Jinkela_wire_19842),
        .dout(new_Jinkela_wire_19843)
    );

    spl2 new_Jinkela_splitter_696 (
        .a(_0440_),
        .b(new_Jinkela_wire_8178),
        .c(new_Jinkela_wire_8179)
    );

    bfr new_Jinkela_buffer_13253 (
        .din(new_Jinkela_wire_15852),
        .dout(new_Jinkela_wire_15853)
    );

    bfr new_Jinkela_buffer_16724 (
        .din(new_Jinkela_wire_19948),
        .dout(new_Jinkela_wire_19949)
    );

    bfr new_Jinkela_buffer_6345 (
        .din(new_Jinkela_wire_8032),
        .dout(new_Jinkela_wire_8033)
    );

    bfr new_Jinkela_buffer_6261 (
        .din(new_Jinkela_wire_7934),
        .dout(new_Jinkela_wire_7935)
    );

    bfr new_Jinkela_buffer_13220 (
        .din(new_Jinkela_wire_15815),
        .dout(new_Jinkela_wire_15816)
    );

    bfr new_Jinkela_buffer_16635 (
        .din(new_Jinkela_wire_19843),
        .dout(new_Jinkela_wire_19844)
    );

    bfr new_Jinkela_buffer_6328 (
        .din(new_Jinkela_wire_8007),
        .dout(new_Jinkela_wire_8008)
    );

    bfr new_Jinkela_buffer_13301 (
        .din(new_Jinkela_wire_15900),
        .dout(new_Jinkela_wire_15901)
    );

    bfr new_Jinkela_buffer_16801 (
        .din(_1241_),
        .dout(new_Jinkela_wire_20046)
    );

    bfr new_Jinkela_buffer_6262 (
        .din(new_Jinkela_wire_7935),
        .dout(new_Jinkela_wire_7936)
    );

    bfr new_Jinkela_buffer_13221 (
        .din(new_Jinkela_wire_15816),
        .dout(new_Jinkela_wire_15817)
    );

    bfr new_Jinkela_buffer_16636 (
        .din(new_Jinkela_wire_19844),
        .dout(new_Jinkela_wire_19845)
    );

    bfr new_Jinkela_buffer_13254 (
        .din(new_Jinkela_wire_15853),
        .dout(new_Jinkela_wire_15854)
    );

    bfr new_Jinkela_buffer_16725 (
        .din(new_Jinkela_wire_19949),
        .dout(new_Jinkela_wire_19950)
    );

    bfr new_Jinkela_buffer_6406 (
        .din(new_Jinkela_wire_8097),
        .dout(new_Jinkela_wire_8098)
    );

    bfr new_Jinkela_buffer_6263 (
        .din(new_Jinkela_wire_7936),
        .dout(new_Jinkela_wire_7937)
    );

    bfr new_Jinkela_buffer_13222 (
        .din(new_Jinkela_wire_15817),
        .dout(new_Jinkela_wire_15818)
    );

    bfr new_Jinkela_buffer_16637 (
        .din(new_Jinkela_wire_19845),
        .dout(new_Jinkela_wire_19846)
    );

    bfr new_Jinkela_buffer_6329 (
        .din(new_Jinkela_wire_8008),
        .dout(new_Jinkela_wire_8009)
    );

    bfr new_Jinkela_buffer_13390 (
        .din(new_Jinkela_wire_15997),
        .dout(new_Jinkela_wire_15998)
    );

    bfr new_Jinkela_buffer_16741 (
        .din(new_Jinkela_wire_19977),
        .dout(new_Jinkela_wire_19978)
    );

    spl2 new_Jinkela_splitter_1154 (
        .a(_1349_),
        .b(new_Jinkela_wire_16008),
        .c(new_Jinkela_wire_16009)
    );

    bfr new_Jinkela_buffer_6264 (
        .din(new_Jinkela_wire_7937),
        .dout(new_Jinkela_wire_7938)
    );

    bfr new_Jinkela_buffer_13223 (
        .din(new_Jinkela_wire_15818),
        .dout(new_Jinkela_wire_15819)
    );

    bfr new_Jinkela_buffer_16638 (
        .din(new_Jinkela_wire_19846),
        .dout(new_Jinkela_wire_19847)
    );

    bfr new_Jinkela_buffer_13255 (
        .din(new_Jinkela_wire_15854),
        .dout(new_Jinkela_wire_15855)
    );

    bfr new_Jinkela_buffer_16726 (
        .din(new_Jinkela_wire_19950),
        .dout(new_Jinkela_wire_19951)
    );

    bfr new_Jinkela_buffer_6265 (
        .din(new_Jinkela_wire_7938),
        .dout(new_Jinkela_wire_7939)
    );

    bfr new_Jinkela_buffer_13224 (
        .din(new_Jinkela_wire_15819),
        .dout(new_Jinkela_wire_15820)
    );

    bfr new_Jinkela_buffer_16639 (
        .din(new_Jinkela_wire_19847),
        .dout(new_Jinkela_wire_19848)
    );

    bfr new_Jinkela_buffer_6330 (
        .din(new_Jinkela_wire_8009),
        .dout(new_Jinkela_wire_8010)
    );

    bfr new_Jinkela_buffer_13302 (
        .din(new_Jinkela_wire_15901),
        .dout(new_Jinkela_wire_15902)
    );

    bfr new_Jinkela_buffer_16800 (
        .din(new_Jinkela_wire_20042),
        .dout(new_Jinkela_wire_20043)
    );

    bfr new_Jinkela_buffer_16802 (
        .din(_1733_),
        .dout(new_Jinkela_wire_20047)
    );

    bfr new_Jinkela_buffer_9721 (
        .din(new_Jinkela_wire_11820),
        .dout(new_Jinkela_wire_11821)
    );

    bfr new_Jinkela_buffer_9861 (
        .din(new_Jinkela_wire_11980),
        .dout(new_Jinkela_wire_11981)
    );

    bfr new_Jinkela_buffer_9722 (
        .din(new_Jinkela_wire_11821),
        .dout(new_Jinkela_wire_11822)
    );

    bfr new_Jinkela_buffer_9772 (
        .din(new_Jinkela_wire_11881),
        .dout(new_Jinkela_wire_11882)
    );

    spl2 new_Jinkela_splitter_899 (
        .a(new_Jinkela_wire_11822),
        .b(new_Jinkela_wire_11823),
        .c(new_Jinkela_wire_11824)
    );

    bfr new_Jinkela_buffer_9773 (
        .din(new_Jinkela_wire_11882),
        .dout(new_Jinkela_wire_11883)
    );

    bfr new_Jinkela_buffer_9862 (
        .din(new_Jinkela_wire_11981),
        .dout(new_Jinkela_wire_11982)
    );

    bfr new_Jinkela_buffer_9774 (
        .din(new_Jinkela_wire_11883),
        .dout(new_Jinkela_wire_11884)
    );

    bfr new_Jinkela_buffer_9931 (
        .din(new_Jinkela_wire_12070),
        .dout(new_Jinkela_wire_12071)
    );

    bfr new_Jinkela_buffer_9775 (
        .din(new_Jinkela_wire_11884),
        .dout(new_Jinkela_wire_11885)
    );

    bfr new_Jinkela_buffer_9863 (
        .din(new_Jinkela_wire_11982),
        .dout(new_Jinkela_wire_11983)
    );

    bfr new_Jinkela_buffer_9776 (
        .din(new_Jinkela_wire_11885),
        .dout(new_Jinkela_wire_11886)
    );

    bfr new_Jinkela_buffer_9965 (
        .din(new_net_3920),
        .dout(new_Jinkela_wire_12111)
    );

    bfr new_Jinkela_buffer_9777 (
        .din(new_Jinkela_wire_11886),
        .dout(new_Jinkela_wire_11887)
    );

    bfr new_Jinkela_buffer_9864 (
        .din(new_Jinkela_wire_11983),
        .dout(new_Jinkela_wire_11984)
    );

    bfr new_Jinkela_buffer_9778 (
        .din(new_Jinkela_wire_11887),
        .dout(new_Jinkela_wire_11888)
    );

    bfr new_Jinkela_buffer_9932 (
        .din(new_Jinkela_wire_12071),
        .dout(new_Jinkela_wire_12072)
    );

    bfr new_Jinkela_buffer_9779 (
        .din(new_Jinkela_wire_11888),
        .dout(new_Jinkela_wire_11889)
    );

    bfr new_Jinkela_buffer_9865 (
        .din(new_Jinkela_wire_11984),
        .dout(new_Jinkela_wire_11985)
    );

    bfr new_Jinkela_buffer_9780 (
        .din(new_Jinkela_wire_11889),
        .dout(new_Jinkela_wire_11890)
    );

    bfr new_Jinkela_buffer_9961 (
        .din(new_Jinkela_wire_12106),
        .dout(new_Jinkela_wire_12107)
    );

    bfr new_Jinkela_buffer_10025 (
        .din(_1575_),
        .dout(new_Jinkela_wire_12171)
    );

    bfr new_Jinkela_buffer_9781 (
        .din(new_Jinkela_wire_11890),
        .dout(new_Jinkela_wire_11891)
    );

    bfr new_Jinkela_buffer_9866 (
        .din(new_Jinkela_wire_11985),
        .dout(new_Jinkela_wire_11986)
    );

    bfr new_Jinkela_buffer_9782 (
        .din(new_Jinkela_wire_11891),
        .dout(new_Jinkela_wire_11892)
    );

    bfr new_Jinkela_buffer_9933 (
        .din(new_Jinkela_wire_12072),
        .dout(new_Jinkela_wire_12073)
    );

    bfr new_Jinkela_buffer_9783 (
        .din(new_Jinkela_wire_11892),
        .dout(new_Jinkela_wire_11893)
    );

    bfr new_Jinkela_buffer_9867 (
        .din(new_Jinkela_wire_11986),
        .dout(new_Jinkela_wire_11987)
    );

    bfr new_Jinkela_buffer_9784 (
        .din(new_Jinkela_wire_11893),
        .dout(new_Jinkela_wire_11894)
    );

    spl2 new_Jinkela_splitter_923 (
        .a(_0659_),
        .b(new_Jinkela_wire_12221),
        .c(new_Jinkela_wire_12222)
    );

    bfr new_Jinkela_buffer_9966 (
        .din(new_Jinkela_wire_12111),
        .dout(new_Jinkela_wire_12112)
    );

    bfr new_Jinkela_buffer_9785 (
        .din(new_Jinkela_wire_11894),
        .dout(new_Jinkela_wire_11895)
    );

    bfr new_Jinkela_buffer_9868 (
        .din(new_Jinkela_wire_11987),
        .dout(new_Jinkela_wire_11988)
    );

    bfr new_Jinkela_buffer_9786 (
        .din(new_Jinkela_wire_11895),
        .dout(new_Jinkela_wire_11896)
    );

    bfr new_Jinkela_buffer_9934 (
        .din(new_Jinkela_wire_12073),
        .dout(new_Jinkela_wire_12074)
    );

    bfr new_Jinkela_buffer_9787 (
        .din(new_Jinkela_wire_11896),
        .dout(new_Jinkela_wire_11897)
    );

    bfr new_Jinkela_buffer_9869 (
        .din(new_Jinkela_wire_11988),
        .dout(new_Jinkela_wire_11989)
    );

    bfr new_Jinkela_buffer_9788 (
        .din(new_Jinkela_wire_11897),
        .dout(new_Jinkela_wire_11898)
    );

    bfr new_Jinkela_buffer_9962 (
        .din(new_Jinkela_wire_12107),
        .dout(new_Jinkela_wire_12108)
    );

    bfr new_Jinkela_buffer_9789 (
        .din(new_Jinkela_wire_11898),
        .dout(new_Jinkela_wire_11899)
    );

    bfr new_Jinkela_buffer_9870 (
        .din(new_Jinkela_wire_11989),
        .dout(new_Jinkela_wire_11990)
    );

    bfr new_Jinkela_buffer_9790 (
        .din(new_Jinkela_wire_11899),
        .dout(new_Jinkela_wire_11900)
    );

    bfr new_Jinkela_buffer_9935 (
        .din(new_Jinkela_wire_12074),
        .dout(new_Jinkela_wire_12075)
    );

    bfr new_Jinkela_buffer_2866 (
        .din(new_Jinkela_wire_3927),
        .dout(new_Jinkela_wire_3928)
    );

    bfr new_Jinkela_buffer_13225 (
        .din(new_Jinkela_wire_15820),
        .dout(new_Jinkela_wire_15821)
    );

    bfr new_Jinkela_buffer_2906 (
        .din(new_Jinkela_wire_3977),
        .dout(new_Jinkela_wire_3978)
    );

    bfr new_Jinkela_buffer_13256 (
        .din(new_Jinkela_wire_15855),
        .dout(new_Jinkela_wire_15856)
    );

    bfr new_Jinkela_buffer_2867 (
        .din(new_Jinkela_wire_3928),
        .dout(new_Jinkela_wire_3929)
    );

    bfr new_Jinkela_buffer_13226 (
        .din(new_Jinkela_wire_15821),
        .dout(new_Jinkela_wire_15822)
    );

    bfr new_Jinkela_buffer_13314 (
        .din(new_Jinkela_wire_15915),
        .dout(new_Jinkela_wire_15916)
    );

    bfr new_Jinkela_buffer_2868 (
        .din(new_Jinkela_wire_3929),
        .dout(new_Jinkela_wire_3930)
    );

    bfr new_Jinkela_buffer_13227 (
        .din(new_Jinkela_wire_15822),
        .dout(new_Jinkela_wire_15823)
    );

    bfr new_Jinkela_buffer_2907 (
        .din(new_Jinkela_wire_3978),
        .dout(new_Jinkela_wire_3979)
    );

    bfr new_Jinkela_buffer_13257 (
        .din(new_Jinkela_wire_15856),
        .dout(new_Jinkela_wire_15857)
    );

    bfr new_Jinkela_buffer_2869 (
        .din(new_Jinkela_wire_3930),
        .dout(new_Jinkela_wire_3931)
    );

    bfr new_Jinkela_buffer_13228 (
        .din(new_Jinkela_wire_15823),
        .dout(new_Jinkela_wire_15824)
    );

    bfr new_Jinkela_buffer_3005 (
        .din(new_Jinkela_wire_4086),
        .dout(new_Jinkela_wire_4087)
    );

    bfr new_Jinkela_buffer_13303 (
        .din(new_Jinkela_wire_15902),
        .dout(new_Jinkela_wire_15903)
    );

    bfr new_Jinkela_buffer_2870 (
        .din(new_Jinkela_wire_3931),
        .dout(new_Jinkela_wire_3932)
    );

    bfr new_Jinkela_buffer_13229 (
        .din(new_Jinkela_wire_15824),
        .dout(new_Jinkela_wire_15825)
    );

    bfr new_Jinkela_buffer_2908 (
        .din(new_Jinkela_wire_3979),
        .dout(new_Jinkela_wire_3980)
    );

    bfr new_Jinkela_buffer_13258 (
        .din(new_Jinkela_wire_15857),
        .dout(new_Jinkela_wire_15858)
    );

    bfr new_Jinkela_buffer_2871 (
        .din(new_Jinkela_wire_3932),
        .dout(new_Jinkela_wire_3933)
    );

    bfr new_Jinkela_buffer_13230 (
        .din(new_Jinkela_wire_15825),
        .dout(new_Jinkela_wire_15826)
    );

    bfr new_Jinkela_buffer_13394 (
        .din(new_Jinkela_wire_16003),
        .dout(new_Jinkela_wire_16004)
    );

    bfr new_Jinkela_buffer_3076 (
        .din(_0707_),
        .dout(new_Jinkela_wire_4166)
    );

    bfr new_Jinkela_buffer_2872 (
        .din(new_Jinkela_wire_3933),
        .dout(new_Jinkela_wire_3934)
    );

    bfr new_Jinkela_buffer_13231 (
        .din(new_Jinkela_wire_15826),
        .dout(new_Jinkela_wire_15827)
    );

    bfr new_Jinkela_buffer_2909 (
        .din(new_Jinkela_wire_3980),
        .dout(new_Jinkela_wire_3981)
    );

    bfr new_Jinkela_buffer_13259 (
        .din(new_Jinkela_wire_15858),
        .dout(new_Jinkela_wire_15859)
    );

    bfr new_Jinkela_buffer_2873 (
        .din(new_Jinkela_wire_3934),
        .dout(new_Jinkela_wire_3935)
    );

    bfr new_Jinkela_buffer_13232 (
        .din(new_Jinkela_wire_15827),
        .dout(new_Jinkela_wire_15828)
    );

    bfr new_Jinkela_buffer_3006 (
        .din(new_Jinkela_wire_4087),
        .dout(new_Jinkela_wire_4088)
    );

    bfr new_Jinkela_buffer_13304 (
        .din(new_Jinkela_wire_15903),
        .dout(new_Jinkela_wire_15904)
    );

    bfr new_Jinkela_buffer_2874 (
        .din(new_Jinkela_wire_3935),
        .dout(new_Jinkela_wire_3936)
    );

    bfr new_Jinkela_buffer_13233 (
        .din(new_Jinkela_wire_15828),
        .dout(new_Jinkela_wire_15829)
    );

    bfr new_Jinkela_buffer_2910 (
        .din(new_Jinkela_wire_3981),
        .dout(new_Jinkela_wire_3982)
    );

    bfr new_Jinkela_buffer_13260 (
        .din(new_Jinkela_wire_15859),
        .dout(new_Jinkela_wire_15860)
    );

    bfr new_Jinkela_buffer_2875 (
        .din(new_Jinkela_wire_3936),
        .dout(new_Jinkela_wire_3937)
    );

    bfr new_Jinkela_buffer_13234 (
        .din(new_Jinkela_wire_15829),
        .dout(new_Jinkela_wire_15830)
    );

    bfr new_Jinkela_buffer_3075 (
        .din(new_Jinkela_wire_4160),
        .dout(new_Jinkela_wire_4161)
    );

    bfr new_Jinkela_buffer_13315 (
        .din(new_Jinkela_wire_15916),
        .dout(new_Jinkela_wire_15917)
    );

    spl2 new_Jinkela_splitter_395 (
        .a(_1071_),
        .b(new_Jinkela_wire_4238),
        .c(new_Jinkela_wire_4239)
    );

    bfr new_Jinkela_buffer_2876 (
        .din(new_Jinkela_wire_3937),
        .dout(new_Jinkela_wire_3938)
    );

    bfr new_Jinkela_buffer_13235 (
        .din(new_Jinkela_wire_15830),
        .dout(new_Jinkela_wire_15831)
    );

    bfr new_Jinkela_buffer_2911 (
        .din(new_Jinkela_wire_3982),
        .dout(new_Jinkela_wire_3983)
    );

    bfr new_Jinkela_buffer_13261 (
        .din(new_Jinkela_wire_15860),
        .dout(new_Jinkela_wire_15861)
    );

    bfr new_Jinkela_buffer_2877 (
        .din(new_Jinkela_wire_3938),
        .dout(new_Jinkela_wire_3939)
    );

    bfr new_Jinkela_buffer_13236 (
        .din(new_Jinkela_wire_15831),
        .dout(new_Jinkela_wire_15832)
    );

    bfr new_Jinkela_buffer_3007 (
        .din(new_Jinkela_wire_4088),
        .dout(new_Jinkela_wire_4089)
    );

    bfr new_Jinkela_buffer_13305 (
        .din(new_Jinkela_wire_15904),
        .dout(new_Jinkela_wire_15905)
    );

    bfr new_Jinkela_buffer_2878 (
        .din(new_Jinkela_wire_3939),
        .dout(new_Jinkela_wire_3940)
    );

    spl2 new_Jinkela_splitter_1147 (
        .a(new_Jinkela_wire_15832),
        .b(new_Jinkela_wire_15833),
        .c(new_Jinkela_wire_15834)
    );

    bfr new_Jinkela_buffer_2912 (
        .din(new_Jinkela_wire_3983),
        .dout(new_Jinkela_wire_3984)
    );

    bfr new_Jinkela_buffer_13391 (
        .din(new_Jinkela_wire_15998),
        .dout(new_Jinkela_wire_15999)
    );

    bfr new_Jinkela_buffer_2879 (
        .din(new_Jinkela_wire_3940),
        .dout(new_Jinkela_wire_3941)
    );

    bfr new_Jinkela_buffer_13262 (
        .din(new_Jinkela_wire_15861),
        .dout(new_Jinkela_wire_15862)
    );

    bfr new_Jinkela_buffer_13263 (
        .din(new_Jinkela_wire_15862),
        .dout(new_Jinkela_wire_15863)
    );

    spl2 new_Jinkela_splitter_392 (
        .a(new_Jinkela_wire_4161),
        .b(new_Jinkela_wire_4162),
        .c(new_Jinkela_wire_4163)
    );

    bfr new_Jinkela_buffer_2880 (
        .din(new_Jinkela_wire_3941),
        .dout(new_Jinkela_wire_3942)
    );

    bfr new_Jinkela_buffer_13306 (
        .din(new_Jinkela_wire_15905),
        .dout(new_Jinkela_wire_15906)
    );

    bfr new_Jinkela_buffer_2913 (
        .din(new_Jinkela_wire_3984),
        .dout(new_Jinkela_wire_3985)
    );

    bfr new_Jinkela_buffer_13264 (
        .din(new_Jinkela_wire_15863),
        .dout(new_Jinkela_wire_15864)
    );

    bfr new_Jinkela_buffer_2881 (
        .din(new_Jinkela_wire_3942),
        .dout(new_Jinkela_wire_3943)
    );

    bfr new_Jinkela_buffer_13316 (
        .din(new_Jinkela_wire_15917),
        .dout(new_Jinkela_wire_15918)
    );

    bfr new_Jinkela_buffer_3008 (
        .din(new_Jinkela_wire_4089),
        .dout(new_Jinkela_wire_4090)
    );

    bfr new_Jinkela_buffer_13265 (
        .din(new_Jinkela_wire_15864),
        .dout(new_Jinkela_wire_15865)
    );

    bfr new_Jinkela_buffer_2882 (
        .din(new_Jinkela_wire_3943),
        .dout(new_Jinkela_wire_3944)
    );

    bfr new_Jinkela_buffer_13307 (
        .din(new_Jinkela_wire_15906),
        .dout(new_Jinkela_wire_15907)
    );

    bfr new_Jinkela_buffer_2914 (
        .din(new_Jinkela_wire_3985),
        .dout(new_Jinkela_wire_3986)
    );

    bfr new_Jinkela_buffer_13266 (
        .din(new_Jinkela_wire_15865),
        .dout(new_Jinkela_wire_15866)
    );

    bfr new_Jinkela_buffer_2883 (
        .din(new_Jinkela_wire_3944),
        .dout(new_Jinkela_wire_3945)
    );

    spl2 new_Jinkela_splitter_1155 (
        .a(_1310_),
        .b(new_Jinkela_wire_16010),
        .c(new_Jinkela_wire_16011)
    );

    bfr new_Jinkela_buffer_13267 (
        .din(new_Jinkela_wire_15866),
        .dout(new_Jinkela_wire_15867)
    );

    bfr new_Jinkela_buffer_3146 (
        .din(_1676_),
        .dout(new_Jinkela_wire_4240)
    );

    bfr new_Jinkela_buffer_2884 (
        .din(new_Jinkela_wire_3945),
        .dout(new_Jinkela_wire_3946)
    );

    bfr new_Jinkela_buffer_13308 (
        .din(new_Jinkela_wire_15907),
        .dout(new_Jinkela_wire_15908)
    );

    bfr new_Jinkela_buffer_2915 (
        .din(new_Jinkela_wire_3986),
        .dout(new_Jinkela_wire_3987)
    );

    bfr new_Jinkela_buffer_13268 (
        .din(new_Jinkela_wire_15867),
        .dout(new_Jinkela_wire_15868)
    );

    bfr new_Jinkela_buffer_2885 (
        .din(new_Jinkela_wire_3946),
        .dout(new_Jinkela_wire_3947)
    );

    bfr new_Jinkela_buffer_13317 (
        .din(new_Jinkela_wire_15918),
        .dout(new_Jinkela_wire_15919)
    );

    bfr new_Jinkela_buffer_3009 (
        .din(new_Jinkela_wire_4090),
        .dout(new_Jinkela_wire_4091)
    );

    bfr new_Jinkela_buffer_13269 (
        .din(new_Jinkela_wire_15868),
        .dout(new_Jinkela_wire_15869)
    );

    bfr new_Jinkela_buffer_2886 (
        .din(new_Jinkela_wire_3947),
        .dout(new_Jinkela_wire_3948)
    );

    bfr new_Jinkela_buffer_13309 (
        .din(new_Jinkela_wire_15908),
        .dout(new_Jinkela_wire_15909)
    );

    bfr new_Jinkela_buffer_2916 (
        .din(new_Jinkela_wire_3987),
        .dout(new_Jinkela_wire_3988)
    );

    bfr new_Jinkela_buffer_13270 (
        .din(new_Jinkela_wire_15869),
        .dout(new_Jinkela_wire_15870)
    );

    bfr new_Jinkela_buffer_6266 (
        .din(new_Jinkela_wire_7939),
        .dout(new_Jinkela_wire_7940)
    );

    bfr new_Jinkela_buffer_6410 (
        .din(new_Jinkela_wire_8101),
        .dout(new_Jinkela_wire_8102)
    );

    bfr new_Jinkela_buffer_6267 (
        .din(new_Jinkela_wire_7940),
        .dout(new_Jinkela_wire_7941)
    );

    bfr new_Jinkela_buffer_6331 (
        .din(new_Jinkela_wire_8010),
        .dout(new_Jinkela_wire_8011)
    );

    bfr new_Jinkela_buffer_6268 (
        .din(new_Jinkela_wire_7941),
        .dout(new_Jinkela_wire_7942)
    );

    bfr new_Jinkela_buffer_6347 (
        .din(new_Jinkela_wire_8034),
        .dout(new_Jinkela_wire_8035)
    );

    bfr new_Jinkela_buffer_6269 (
        .din(new_Jinkela_wire_7942),
        .dout(new_Jinkela_wire_7943)
    );

    bfr new_Jinkela_buffer_6332 (
        .din(new_Jinkela_wire_8011),
        .dout(new_Jinkela_wire_8012)
    );

    bfr new_Jinkela_buffer_6270 (
        .din(new_Jinkela_wire_7943),
        .dout(new_Jinkela_wire_7944)
    );

    bfr new_Jinkela_buffer_6407 (
        .din(new_Jinkela_wire_8098),
        .dout(new_Jinkela_wire_8099)
    );

    bfr new_Jinkela_buffer_6271 (
        .din(new_Jinkela_wire_7944),
        .dout(new_Jinkela_wire_7945)
    );

    bfr new_Jinkela_buffer_6333 (
        .din(new_Jinkela_wire_8012),
        .dout(new_Jinkela_wire_8013)
    );

    bfr new_Jinkela_buffer_6272 (
        .din(new_Jinkela_wire_7945),
        .dout(new_Jinkela_wire_7946)
    );

    bfr new_Jinkela_buffer_6348 (
        .din(new_Jinkela_wire_8035),
        .dout(new_Jinkela_wire_8036)
    );

    bfr new_Jinkela_buffer_6273 (
        .din(new_Jinkela_wire_7946),
        .dout(new_Jinkela_wire_7947)
    );

    bfr new_Jinkela_buffer_6334 (
        .din(new_Jinkela_wire_8013),
        .dout(new_Jinkela_wire_8014)
    );

    bfr new_Jinkela_buffer_6274 (
        .din(new_Jinkela_wire_7947),
        .dout(new_Jinkela_wire_7948)
    );

    bfr new_Jinkela_buffer_6484 (
        .din(_1351_),
        .dout(new_Jinkela_wire_8180)
    );

    bfr new_Jinkela_buffer_6275 (
        .din(new_Jinkela_wire_7948),
        .dout(new_Jinkela_wire_7949)
    );

    bfr new_Jinkela_buffer_6335 (
        .din(new_Jinkela_wire_8014),
        .dout(new_Jinkela_wire_8015)
    );

    bfr new_Jinkela_buffer_6276 (
        .din(new_Jinkela_wire_7949),
        .dout(new_Jinkela_wire_7950)
    );

    bfr new_Jinkela_buffer_6349 (
        .din(new_Jinkela_wire_8036),
        .dout(new_Jinkela_wire_8037)
    );

    bfr new_Jinkela_buffer_6277 (
        .din(new_Jinkela_wire_7950),
        .dout(new_Jinkela_wire_7951)
    );

    spl2 new_Jinkela_splitter_689 (
        .a(new_Jinkela_wire_8015),
        .b(new_Jinkela_wire_8016),
        .c(new_Jinkela_wire_8017)
    );

    bfr new_Jinkela_buffer_6278 (
        .din(new_Jinkela_wire_7951),
        .dout(new_Jinkela_wire_7952)
    );

    bfr new_Jinkela_buffer_6350 (
        .din(new_Jinkela_wire_8037),
        .dout(new_Jinkela_wire_8038)
    );

    bfr new_Jinkela_buffer_6279 (
        .din(new_Jinkela_wire_7952),
        .dout(new_Jinkela_wire_7953)
    );

    bfr new_Jinkela_buffer_6408 (
        .din(new_Jinkela_wire_8099),
        .dout(new_Jinkela_wire_8100)
    );

    bfr new_Jinkela_buffer_6280 (
        .din(new_Jinkela_wire_7953),
        .dout(new_Jinkela_wire_7954)
    );

    bfr new_Jinkela_buffer_6411 (
        .din(new_Jinkela_wire_8102),
        .dout(new_Jinkela_wire_8103)
    );

    bfr new_Jinkela_buffer_6281 (
        .din(new_Jinkela_wire_7954),
        .dout(new_Jinkela_wire_7955)
    );

    bfr new_Jinkela_buffer_6351 (
        .din(new_Jinkela_wire_8038),
        .dout(new_Jinkela_wire_8039)
    );

    bfr new_Jinkela_buffer_6282 (
        .din(new_Jinkela_wire_7955),
        .dout(new_Jinkela_wire_7956)
    );

    spl2 new_Jinkela_splitter_697 (
        .a(_1013_),
        .b(new_Jinkela_wire_8181),
        .c(new_Jinkela_wire_8182)
    );

    bfr new_Jinkela_buffer_6283 (
        .din(new_Jinkela_wire_7956),
        .dout(new_Jinkela_wire_7957)
    );

    bfr new_Jinkela_buffer_6352 (
        .din(new_Jinkela_wire_8039),
        .dout(new_Jinkela_wire_8040)
    );

    bfr new_Jinkela_buffer_6284 (
        .din(new_Jinkela_wire_7957),
        .dout(new_Jinkela_wire_7958)
    );

    bfr new_Jinkela_buffer_6412 (
        .din(new_Jinkela_wire_8103),
        .dout(new_Jinkela_wire_8104)
    );

    bfr new_Jinkela_buffer_6285 (
        .din(new_Jinkela_wire_7958),
        .dout(new_Jinkela_wire_7959)
    );

    bfr new_Jinkela_buffer_6353 (
        .din(new_Jinkela_wire_8040),
        .dout(new_Jinkela_wire_8041)
    );

    bfr new_Jinkela_buffer_6286 (
        .din(new_Jinkela_wire_7959),
        .dout(new_Jinkela_wire_7960)
    );

    bfr new_Jinkela_buffer_6346 (
        .din(new_Jinkela_wire_8033),
        .dout(new_Jinkela_wire_8034)
    );

    and_bi _3676_ (
        .a(new_Jinkela_wire_1332),
        .b(new_Jinkela_wire_10560),
        .c(_0983_)
    );

    bfr new_Jinkela_buffer_16640 (
        .din(new_Jinkela_wire_19848),
        .dout(new_Jinkela_wire_19849)
    );

    and_bi _3677_ (
        .a(new_Jinkela_wire_10561),
        .b(new_Jinkela_wire_1333),
        .c(_0984_)
    );

    bfr new_Jinkela_buffer_16727 (
        .din(new_Jinkela_wire_19951),
        .dout(new_Jinkela_wire_19952)
    );

    or_bb _3678_ (
        .a(new_Jinkela_wire_1018),
        .b(new_Jinkela_wire_10682),
        .c(new_net_3972)
    );

    bfr new_Jinkela_buffer_16641 (
        .din(new_Jinkela_wire_19849),
        .dout(new_Jinkela_wire_19850)
    );

    and_ii _3679_ (
        .a(new_Jinkela_wire_10683),
        .b(new_Jinkela_wire_17160),
        .c(_0985_)
    );

    bfr new_Jinkela_buffer_16742 (
        .din(new_Jinkela_wire_19978),
        .dout(new_Jinkela_wire_19979)
    );

    and_ii _3680_ (
        .a(new_Jinkela_wire_722),
        .b(new_Jinkela_wire_17541),
        .c(_0986_)
    );

    bfr new_Jinkela_buffer_16642 (
        .din(new_Jinkela_wire_19850),
        .dout(new_Jinkela_wire_19851)
    );

    and_bb _3681_ (
        .a(new_Jinkela_wire_603),
        .b(new_Jinkela_wire_672),
        .c(_0987_)
    );

    bfr new_Jinkela_buffer_16728 (
        .din(new_Jinkela_wire_19952),
        .dout(new_Jinkela_wire_19953)
    );

    and_bb _3682_ (
        .a(new_Jinkela_wire_416),
        .b(new_Jinkela_wire_521),
        .c(_0988_)
    );

    bfr new_Jinkela_buffer_16643 (
        .din(new_Jinkela_wire_19851),
        .dout(new_Jinkela_wire_19852)
    );

    and_ii _3683_ (
        .a(new_Jinkela_wire_21191),
        .b(new_Jinkela_wire_6853),
        .c(_0990_)
    );

    bfr new_Jinkela_buffer_16803 (
        .din(_0526_),
        .dout(new_Jinkela_wire_20048)
    );

    and_ii _3684_ (
        .a(new_Jinkela_wire_10097),
        .b(new_Jinkela_wire_11720),
        .c(_0991_)
    );

    bfr new_Jinkela_buffer_16644 (
        .din(new_Jinkela_wire_19852),
        .dout(new_Jinkela_wire_19853)
    );

    and_bb _3685_ (
        .a(new_Jinkela_wire_10098),
        .b(new_Jinkela_wire_11721),
        .c(_0992_)
    );

    bfr new_Jinkela_buffer_16729 (
        .din(new_Jinkela_wire_19953),
        .dout(new_Jinkela_wire_19954)
    );

    or_bb _3686_ (
        .a(new_Jinkela_wire_2261),
        .b(new_Jinkela_wire_15676),
        .c(_0993_)
    );

    bfr new_Jinkela_buffer_16645 (
        .din(new_Jinkela_wire_19853),
        .dout(new_Jinkela_wire_19854)
    );

    and_ii _3687_ (
        .a(new_Jinkela_wire_10751),
        .b(new_Jinkela_wire_14536),
        .c(_0994_)
    );

    bfr new_Jinkela_buffer_16743 (
        .din(new_Jinkela_wire_19979),
        .dout(new_Jinkela_wire_19980)
    );

    and_bb _3688_ (
        .a(new_Jinkela_wire_10752),
        .b(new_Jinkela_wire_14537),
        .c(_0995_)
    );

    bfr new_Jinkela_buffer_16646 (
        .din(new_Jinkela_wire_19854),
        .dout(new_Jinkela_wire_19855)
    );

    or_bb _3689_ (
        .a(new_Jinkela_wire_14265),
        .b(new_Jinkela_wire_2257),
        .c(_0996_)
    );

    bfr new_Jinkela_buffer_16730 (
        .din(new_Jinkela_wire_19954),
        .dout(new_Jinkela_wire_19955)
    );

    and_ii _3690_ (
        .a(new_Jinkela_wire_14004),
        .b(new_Jinkela_wire_16796),
        .c(_0997_)
    );

    bfr new_Jinkela_buffer_16647 (
        .din(new_Jinkela_wire_19855),
        .dout(new_Jinkela_wire_19856)
    );

    and_bb _3691_ (
        .a(new_Jinkela_wire_14005),
        .b(new_Jinkela_wire_16797),
        .c(_0998_)
    );

    spl2 new_Jinkela_splitter_1470 (
        .a(new_Jinkela_wire_20043),
        .b(new_Jinkela_wire_20044),
        .c(new_Jinkela_wire_20045)
    );

    and_ii _3692_ (
        .a(new_Jinkela_wire_16509),
        .b(new_Jinkela_wire_15837),
        .c(_0999_)
    );

    bfr new_Jinkela_buffer_16648 (
        .din(new_Jinkela_wire_19856),
        .dout(new_Jinkela_wire_19857)
    );

    and_bi _3693_ (
        .a(new_Jinkela_wire_15833),
        .b(new_Jinkela_wire_21094),
        .c(_1001_)
    );

    bfr new_Jinkela_buffer_16731 (
        .din(new_Jinkela_wire_19955),
        .dout(new_Jinkela_wire_19956)
    );

    and_bi _3694_ (
        .a(new_Jinkela_wire_21095),
        .b(new_Jinkela_wire_15834),
        .c(_1002_)
    );

    bfr new_Jinkela_buffer_16649 (
        .din(new_Jinkela_wire_19857),
        .dout(new_Jinkela_wire_19858)
    );

    or_bb _3695_ (
        .a(new_Jinkela_wire_11400),
        .b(new_Jinkela_wire_8760),
        .c(new_net_3938)
    );

    bfr new_Jinkela_buffer_16744 (
        .din(new_Jinkela_wire_19980),
        .dout(new_Jinkela_wire_19981)
    );

    and_bb _3696_ (
        .a(new_Jinkela_wire_421),
        .b(new_Jinkela_wire_663),
        .c(_1003_)
    );

    bfr new_Jinkela_buffer_16650 (
        .din(new_Jinkela_wire_19858),
        .dout(new_Jinkela_wire_19859)
    );

    and_ii _3697_ (
        .a(new_Jinkela_wire_2258),
        .b(new_Jinkela_wire_15681),
        .c(_1004_)
    );

    bfr new_Jinkela_buffer_16732 (
        .din(new_Jinkela_wire_19956),
        .dout(new_Jinkela_wire_19957)
    );

    or_bb _3698_ (
        .a(new_Jinkela_wire_13997),
        .b(new_Jinkela_wire_20793),
        .c(_1005_)
    );

    bfr new_Jinkela_buffer_16651 (
        .din(new_Jinkela_wire_19859),
        .dout(new_Jinkela_wire_19860)
    );

    and_ii _3699_ (
        .a(new_Jinkela_wire_8761),
        .b(new_Jinkela_wire_15892),
        .c(_1006_)
    );

    and_bb _3700_ (
        .a(new_Jinkela_wire_13998),
        .b(new_Jinkela_wire_20794),
        .c(_1007_)
    );

    bfr new_Jinkela_buffer_16652 (
        .din(new_Jinkela_wire_19860),
        .dout(new_Jinkela_wire_19861)
    );

    and_bi _3701_ (
        .a(new_Jinkela_wire_9446),
        .b(new_Jinkela_wire_20219),
        .c(_1008_)
    );

    spl2 new_Jinkela_splitter_1461 (
        .a(new_Jinkela_wire_19957),
        .b(new_Jinkela_wire_19958),
        .c(new_Jinkela_wire_19959)
    );

    and_bi _3702_ (
        .a(new_Jinkela_wire_8359),
        .b(new_Jinkela_wire_13584),
        .c(_1009_)
    );

    bfr new_Jinkela_buffer_16653 (
        .din(new_Jinkela_wire_19861),
        .dout(new_Jinkela_wire_19862)
    );

    and_bi _3703_ (
        .a(new_Jinkela_wire_9509),
        .b(new_Jinkela_wire_2124),
        .c(N6287)
    );

    bfr new_Jinkela_buffer_16885 (
        .din(_0145_),
        .dout(new_Jinkela_wire_20134)
    );

    spl2 new_Jinkela_splitter_1471 (
        .a(_1353_),
        .b(new_Jinkela_wire_20049),
        .c(new_Jinkela_wire_20050)
    );

    and_bi _3704_ (
        .a(new_Jinkela_wire_13585),
        .b(new_Jinkela_wire_8360),
        .c(_1011_)
    );

    bfr new_Jinkela_buffer_16654 (
        .din(new_Jinkela_wire_19862),
        .dout(new_Jinkela_wire_19863)
    );

    or_bb _3705_ (
        .a(new_Jinkela_wire_6376),
        .b(new_Jinkela_wire_2125),
        .c(N6288)
    );

    bfr new_Jinkela_buffer_16745 (
        .din(new_Jinkela_wire_19981),
        .dout(new_Jinkela_wire_19982)
    );

    and_bb _3706_ (
        .a(new_Jinkela_wire_9743),
        .b(new_Jinkela_wire_20286),
        .c(_1012_)
    );

    bfr new_Jinkela_buffer_16655 (
        .din(new_Jinkela_wire_19863),
        .dout(new_Jinkela_wire_19864)
    );

    and_bi _3707_ (
        .a(new_Jinkela_wire_4159),
        .b(new_Jinkela_wire_8185),
        .c(new_net_3940)
    );

    bfr new_Jinkela_buffer_16746 (
        .din(new_Jinkela_wire_19982),
        .dout(new_Jinkela_wire_19983)
    );

    bfr new_Jinkela_buffer_16656 (
        .din(new_Jinkela_wire_19864),
        .dout(new_Jinkela_wire_19865)
    );

    bfr new_Jinkela_buffer_16804 (
        .din(_0441_),
        .dout(new_Jinkela_wire_20051)
    );

    bfr new_Jinkela_buffer_16657 (
        .din(new_Jinkela_wire_19865),
        .dout(new_Jinkela_wire_19866)
    );

    bfr new_Jinkela_buffer_16747 (
        .din(new_Jinkela_wire_19983),
        .dout(new_Jinkela_wire_19984)
    );

    bfr new_Jinkela_buffer_16658 (
        .din(new_Jinkela_wire_19866),
        .dout(new_Jinkela_wire_19867)
    );

    bfr new_Jinkela_buffer_16884 (
        .din(_1256_),
        .dout(new_Jinkela_wire_20133)
    );

    bfr new_Jinkela_buffer_16659 (
        .din(new_Jinkela_wire_19867),
        .dout(new_Jinkela_wire_19868)
    );

    bfr new_Jinkela_buffer_16748 (
        .din(new_Jinkela_wire_19984),
        .dout(new_Jinkela_wire_19985)
    );

    bfr new_Jinkela_buffer_16660 (
        .din(new_Jinkela_wire_19868),
        .dout(new_Jinkela_wire_19869)
    );

    bfr new_Jinkela_buffer_16805 (
        .din(new_Jinkela_wire_20051),
        .dout(new_Jinkela_wire_20052)
    );

    bfr new_Jinkela_buffer_2887 (
        .din(new_Jinkela_wire_3948),
        .dout(new_Jinkela_wire_3949)
    );

    bfr new_Jinkela_buffer_13392 (
        .din(new_Jinkela_wire_15999),
        .dout(new_Jinkela_wire_16000)
    );

    spl2 new_Jinkela_splitter_397 (
        .a(_1579_),
        .b(new_Jinkela_wire_4243),
        .c(new_Jinkela_wire_4244)
    );

    bfr new_Jinkela_buffer_13271 (
        .din(new_Jinkela_wire_15870),
        .dout(new_Jinkela_wire_15871)
    );

    bfr new_Jinkela_buffer_3077 (
        .din(new_Jinkela_wire_4166),
        .dout(new_Jinkela_wire_4167)
    );

    spl2 new_Jinkela_splitter_380 (
        .a(new_Jinkela_wire_3949),
        .b(new_Jinkela_wire_3950),
        .c(new_Jinkela_wire_3951)
    );

    spl2 new_Jinkela_splitter_1149 (
        .a(new_Jinkela_wire_15909),
        .b(new_Jinkela_wire_15910),
        .c(new_Jinkela_wire_15911)
    );

    bfr new_Jinkela_buffer_3010 (
        .din(new_Jinkela_wire_4091),
        .dout(new_Jinkela_wire_4092)
    );

    bfr new_Jinkela_buffer_13272 (
        .din(new_Jinkela_wire_15871),
        .dout(new_Jinkela_wire_15872)
    );

    bfr new_Jinkela_buffer_2917 (
        .din(new_Jinkela_wire_3988),
        .dout(new_Jinkela_wire_3989)
    );

    bfr new_Jinkela_buffer_13492 (
        .din(new_Jinkela_wire_16129),
        .dout(new_Jinkela_wire_16130)
    );

    bfr new_Jinkela_buffer_13419 (
        .din(new_Jinkela_wire_16032),
        .dout(new_Jinkela_wire_16033)
    );

    bfr new_Jinkela_buffer_2918 (
        .din(new_Jinkela_wire_3989),
        .dout(new_Jinkela_wire_3990)
    );

    bfr new_Jinkela_buffer_13273 (
        .din(new_Jinkela_wire_15872),
        .dout(new_Jinkela_wire_15873)
    );

    bfr new_Jinkela_buffer_13318 (
        .din(new_Jinkela_wire_15919),
        .dout(new_Jinkela_wire_15920)
    );

    bfr new_Jinkela_buffer_2919 (
        .din(new_Jinkela_wire_3990),
        .dout(new_Jinkela_wire_3991)
    );

    bfr new_Jinkela_buffer_13274 (
        .din(new_Jinkela_wire_15873),
        .dout(new_Jinkela_wire_15874)
    );

    bfr new_Jinkela_buffer_3011 (
        .din(new_Jinkela_wire_4092),
        .dout(new_Jinkela_wire_4093)
    );

    bfr new_Jinkela_buffer_13319 (
        .din(new_Jinkela_wire_15920),
        .dout(new_Jinkela_wire_15921)
    );

    bfr new_Jinkela_buffer_2920 (
        .din(new_Jinkela_wire_3991),
        .dout(new_Jinkela_wire_3992)
    );

    bfr new_Jinkela_buffer_13275 (
        .din(new_Jinkela_wire_15874),
        .dout(new_Jinkela_wire_15875)
    );

    bfr new_Jinkela_buffer_3078 (
        .din(new_Jinkela_wire_4167),
        .dout(new_Jinkela_wire_4168)
    );

    bfr new_Jinkela_buffer_13393 (
        .din(new_Jinkela_wire_16000),
        .dout(new_Jinkela_wire_16001)
    );

    bfr new_Jinkela_buffer_2921 (
        .din(new_Jinkela_wire_3992),
        .dout(new_Jinkela_wire_3993)
    );

    bfr new_Jinkela_buffer_13276 (
        .din(new_Jinkela_wire_15875),
        .dout(new_Jinkela_wire_15876)
    );

    bfr new_Jinkela_buffer_3012 (
        .din(new_Jinkela_wire_4093),
        .dout(new_Jinkela_wire_4094)
    );

    bfr new_Jinkela_buffer_13320 (
        .din(new_Jinkela_wire_15921),
        .dout(new_Jinkela_wire_15922)
    );

    bfr new_Jinkela_buffer_2922 (
        .din(new_Jinkela_wire_3993),
        .dout(new_Jinkela_wire_3994)
    );

    bfr new_Jinkela_buffer_13277 (
        .din(new_Jinkela_wire_15876),
        .dout(new_Jinkela_wire_15877)
    );

    bfr new_Jinkela_buffer_13395 (
        .din(new_Jinkela_wire_16004),
        .dout(new_Jinkela_wire_16005)
    );

    spl2 new_Jinkela_splitter_396 (
        .a(_0000_),
        .b(new_Jinkela_wire_4241),
        .c(new_Jinkela_wire_4242)
    );

    bfr new_Jinkela_buffer_2923 (
        .din(new_Jinkela_wire_3994),
        .dout(new_Jinkela_wire_3995)
    );

    bfr new_Jinkela_buffer_13278 (
        .din(new_Jinkela_wire_15877),
        .dout(new_Jinkela_wire_15878)
    );

    bfr new_Jinkela_buffer_3013 (
        .din(new_Jinkela_wire_4094),
        .dout(new_Jinkela_wire_4095)
    );

    bfr new_Jinkela_buffer_13321 (
        .din(new_Jinkela_wire_15922),
        .dout(new_Jinkela_wire_15923)
    );

    bfr new_Jinkela_buffer_2924 (
        .din(new_Jinkela_wire_3995),
        .dout(new_Jinkela_wire_3996)
    );

    bfr new_Jinkela_buffer_13279 (
        .din(new_Jinkela_wire_15878),
        .dout(new_Jinkela_wire_15879)
    );

    bfr new_Jinkela_buffer_3079 (
        .din(new_Jinkela_wire_4168),
        .dout(new_Jinkela_wire_4169)
    );

    spl2 new_Jinkela_splitter_1170 (
        .a(_1025_),
        .b(new_Jinkela_wire_16192),
        .c(new_Jinkela_wire_16193)
    );

    bfr new_Jinkela_buffer_2925 (
        .din(new_Jinkela_wire_3996),
        .dout(new_Jinkela_wire_3997)
    );

    bfr new_Jinkela_buffer_13280 (
        .din(new_Jinkela_wire_15879),
        .dout(new_Jinkela_wire_15880)
    );

    bfr new_Jinkela_buffer_3014 (
        .din(new_Jinkela_wire_4095),
        .dout(new_Jinkela_wire_4096)
    );

    bfr new_Jinkela_buffer_13322 (
        .din(new_Jinkela_wire_15923),
        .dout(new_Jinkela_wire_15924)
    );

    bfr new_Jinkela_buffer_2926 (
        .din(new_Jinkela_wire_3997),
        .dout(new_Jinkela_wire_3998)
    );

    bfr new_Jinkela_buffer_13281 (
        .din(new_Jinkela_wire_15880),
        .dout(new_Jinkela_wire_15881)
    );

    bfr new_Jinkela_buffer_13396 (
        .din(new_Jinkela_wire_16005),
        .dout(new_Jinkela_wire_16006)
    );

    bfr new_Jinkela_buffer_2927 (
        .din(new_Jinkela_wire_3998),
        .dout(new_Jinkela_wire_3999)
    );

    bfr new_Jinkela_buffer_13282 (
        .din(new_Jinkela_wire_15881),
        .dout(new_Jinkela_wire_15882)
    );

    bfr new_Jinkela_buffer_3015 (
        .din(new_Jinkela_wire_4096),
        .dout(new_Jinkela_wire_4097)
    );

    bfr new_Jinkela_buffer_13323 (
        .din(new_Jinkela_wire_15924),
        .dout(new_Jinkela_wire_15925)
    );

    bfr new_Jinkela_buffer_2928 (
        .din(new_Jinkela_wire_3999),
        .dout(new_Jinkela_wire_4000)
    );

    bfr new_Jinkela_buffer_13283 (
        .din(new_Jinkela_wire_15882),
        .dout(new_Jinkela_wire_15883)
    );

    bfr new_Jinkela_buffer_3080 (
        .din(new_Jinkela_wire_4169),
        .dout(new_Jinkela_wire_4170)
    );

    bfr new_Jinkela_buffer_2929 (
        .din(new_Jinkela_wire_4000),
        .dout(new_Jinkela_wire_4001)
    );

    bfr new_Jinkela_buffer_13284 (
        .din(new_Jinkela_wire_15883),
        .dout(new_Jinkela_wire_15884)
    );

    bfr new_Jinkela_buffer_3016 (
        .din(new_Jinkela_wire_4097),
        .dout(new_Jinkela_wire_4098)
    );

    bfr new_Jinkela_buffer_13324 (
        .din(new_Jinkela_wire_15925),
        .dout(new_Jinkela_wire_15926)
    );

    bfr new_Jinkela_buffer_2930 (
        .din(new_Jinkela_wire_4001),
        .dout(new_Jinkela_wire_4002)
    );

    bfr new_Jinkela_buffer_13285 (
        .din(new_Jinkela_wire_15884),
        .dout(new_Jinkela_wire_15885)
    );

    bfr new_Jinkela_buffer_13397 (
        .din(new_Jinkela_wire_16006),
        .dout(new_Jinkela_wire_16007)
    );

    spl2 new_Jinkela_splitter_398 (
        .a(_0901_),
        .b(new_Jinkela_wire_4245),
        .c(new_Jinkela_wire_4246)
    );

    bfr new_Jinkela_buffer_2931 (
        .din(new_Jinkela_wire_4002),
        .dout(new_Jinkela_wire_4003)
    );

    bfr new_Jinkela_buffer_13286 (
        .din(new_Jinkela_wire_15885),
        .dout(new_Jinkela_wire_15886)
    );

    bfr new_Jinkela_buffer_3017 (
        .din(new_Jinkela_wire_4098),
        .dout(new_Jinkela_wire_4099)
    );

    bfr new_Jinkela_buffer_13325 (
        .din(new_Jinkela_wire_15926),
        .dout(new_Jinkela_wire_15927)
    );

    bfr new_Jinkela_buffer_2932 (
        .din(new_Jinkela_wire_4003),
        .dout(new_Jinkela_wire_4004)
    );

    bfr new_Jinkela_buffer_13287 (
        .din(new_Jinkela_wire_15886),
        .dout(new_Jinkela_wire_15887)
    );

    bfr new_Jinkela_buffer_3081 (
        .din(new_Jinkela_wire_4170),
        .dout(new_Jinkela_wire_4171)
    );

    bfr new_Jinkela_buffer_13420 (
        .din(new_Jinkela_wire_16033),
        .dout(new_Jinkela_wire_16034)
    );

    bfr new_Jinkela_buffer_2933 (
        .din(new_Jinkela_wire_4004),
        .dout(new_Jinkela_wire_4005)
    );

    bfr new_Jinkela_buffer_13288 (
        .din(new_Jinkela_wire_15887),
        .dout(new_Jinkela_wire_15888)
    );

    bfr new_Jinkela_buffer_3018 (
        .din(new_Jinkela_wire_4099),
        .dout(new_Jinkela_wire_4100)
    );

    bfr new_Jinkela_buffer_13326 (
        .din(new_Jinkela_wire_15927),
        .dout(new_Jinkela_wire_15928)
    );

    bfr new_Jinkela_buffer_2934 (
        .din(new_Jinkela_wire_4005),
        .dout(new_Jinkela_wire_4006)
    );

    bfr new_Jinkela_buffer_13289 (
        .din(new_Jinkela_wire_15888),
        .dout(new_Jinkela_wire_15889)
    );

    bfr new_Jinkela_buffer_3148 (
        .din(_0815_),
        .dout(new_Jinkela_wire_4248)
    );

    bfr new_Jinkela_buffer_3147 (
        .din(_1746_),
        .dout(new_Jinkela_wire_4247)
    );

    bfr new_Jinkela_buffer_13495 (
        .din(new_Jinkela_wire_16132),
        .dout(new_Jinkela_wire_16133)
    );

    bfr new_Jinkela_buffer_2935 (
        .din(new_Jinkela_wire_4006),
        .dout(new_Jinkela_wire_4007)
    );

    bfr new_Jinkela_buffer_13290 (
        .din(new_Jinkela_wire_15889),
        .dout(new_Jinkela_wire_15890)
    );

    bfr new_Jinkela_buffer_3019 (
        .din(new_Jinkela_wire_4100),
        .dout(new_Jinkela_wire_4101)
    );

    bfr new_Jinkela_buffer_13327 (
        .din(new_Jinkela_wire_15928),
        .dout(new_Jinkela_wire_15929)
    );

    bfr new_Jinkela_buffer_2936 (
        .din(new_Jinkela_wire_4007),
        .dout(new_Jinkela_wire_4008)
    );

    bfr new_Jinkela_buffer_13291 (
        .din(new_Jinkela_wire_15890),
        .dout(new_Jinkela_wire_15891)
    );

    bfr new_Jinkela_buffer_6287 (
        .din(new_Jinkela_wire_7960),
        .dout(new_Jinkela_wire_7961)
    );

    bfr new_Jinkela_buffer_9791 (
        .din(new_Jinkela_wire_11900),
        .dout(new_Jinkela_wire_11901)
    );

    bfr new_Jinkela_buffer_16661 (
        .din(new_Jinkela_wire_19869),
        .dout(new_Jinkela_wire_19870)
    );

    bfr new_Jinkela_buffer_6358 (
        .din(new_Jinkela_wire_8045),
        .dout(new_Jinkela_wire_8046)
    );

    bfr new_Jinkela_buffer_9871 (
        .din(new_Jinkela_wire_11990),
        .dout(new_Jinkela_wire_11991)
    );

    bfr new_Jinkela_buffer_16749 (
        .din(new_Jinkela_wire_19985),
        .dout(new_Jinkela_wire_19986)
    );

    bfr new_Jinkela_buffer_6288 (
        .din(new_Jinkela_wire_7961),
        .dout(new_Jinkela_wire_7962)
    );

    bfr new_Jinkela_buffer_9792 (
        .din(new_Jinkela_wire_11901),
        .dout(new_Jinkela_wire_11902)
    );

    bfr new_Jinkela_buffer_16662 (
        .din(new_Jinkela_wire_19870),
        .dout(new_Jinkela_wire_19871)
    );

    bfr new_Jinkela_buffer_6415 (
        .din(new_Jinkela_wire_8106),
        .dout(new_Jinkela_wire_8107)
    );

    bfr new_Jinkela_buffer_16886 (
        .din(_0376_),
        .dout(new_Jinkela_wire_20135)
    );

    bfr new_Jinkela_buffer_6289 (
        .din(new_Jinkela_wire_7962),
        .dout(new_Jinkela_wire_7963)
    );

    bfr new_Jinkela_buffer_9793 (
        .din(new_Jinkela_wire_11902),
        .dout(new_Jinkela_wire_11903)
    );

    bfr new_Jinkela_buffer_16663 (
        .din(new_Jinkela_wire_19871),
        .dout(new_Jinkela_wire_19872)
    );

    bfr new_Jinkela_buffer_6359 (
        .din(new_Jinkela_wire_8046),
        .dout(new_Jinkela_wire_8047)
    );

    bfr new_Jinkela_buffer_9872 (
        .din(new_Jinkela_wire_11991),
        .dout(new_Jinkela_wire_11992)
    );

    bfr new_Jinkela_buffer_16750 (
        .din(new_Jinkela_wire_19986),
        .dout(new_Jinkela_wire_19987)
    );

    bfr new_Jinkela_buffer_6290 (
        .din(new_Jinkela_wire_7963),
        .dout(new_Jinkela_wire_7964)
    );

    bfr new_Jinkela_buffer_9794 (
        .din(new_Jinkela_wire_11903),
        .dout(new_Jinkela_wire_11904)
    );

    bfr new_Jinkela_buffer_16664 (
        .din(new_Jinkela_wire_19872),
        .dout(new_Jinkela_wire_19873)
    );

    bfr new_Jinkela_buffer_9936 (
        .din(new_Jinkela_wire_12075),
        .dout(new_Jinkela_wire_12076)
    );

    bfr new_Jinkela_buffer_16806 (
        .din(new_Jinkela_wire_20052),
        .dout(new_Jinkela_wire_20053)
    );

    bfr new_Jinkela_buffer_6487 (
        .din(new_net_3964),
        .dout(new_Jinkela_wire_8187)
    );

    bfr new_Jinkela_buffer_6291 (
        .din(new_Jinkela_wire_7964),
        .dout(new_Jinkela_wire_7965)
    );

    bfr new_Jinkela_buffer_9795 (
        .din(new_Jinkela_wire_11904),
        .dout(new_Jinkela_wire_11905)
    );

    bfr new_Jinkela_buffer_16665 (
        .din(new_Jinkela_wire_19873),
        .dout(new_Jinkela_wire_19874)
    );

    bfr new_Jinkela_buffer_6360 (
        .din(new_Jinkela_wire_8047),
        .dout(new_Jinkela_wire_8048)
    );

    bfr new_Jinkela_buffer_9873 (
        .din(new_Jinkela_wire_11992),
        .dout(new_Jinkela_wire_11993)
    );

    bfr new_Jinkela_buffer_16751 (
        .din(new_Jinkela_wire_19987),
        .dout(new_Jinkela_wire_19988)
    );

    bfr new_Jinkela_buffer_6292 (
        .din(new_Jinkela_wire_7965),
        .dout(new_Jinkela_wire_7966)
    );

    bfr new_Jinkela_buffer_9796 (
        .din(new_Jinkela_wire_11905),
        .dout(new_Jinkela_wire_11906)
    );

    bfr new_Jinkela_buffer_16666 (
        .din(new_Jinkela_wire_19874),
        .dout(new_Jinkela_wire_19875)
    );

    bfr new_Jinkela_buffer_6416 (
        .din(new_Jinkela_wire_8107),
        .dout(new_Jinkela_wire_8108)
    );

    bfr new_Jinkela_buffer_9963 (
        .din(new_Jinkela_wire_12108),
        .dout(new_Jinkela_wire_12109)
    );

    spl2 new_Jinkela_splitter_1473 (
        .a(_0642_),
        .b(new_Jinkela_wire_20136),
        .c(new_Jinkela_wire_20137)
    );

    bfr new_Jinkela_buffer_6293 (
        .din(new_Jinkela_wire_7966),
        .dout(new_Jinkela_wire_7967)
    );

    bfr new_Jinkela_buffer_9797 (
        .din(new_Jinkela_wire_11906),
        .dout(new_Jinkela_wire_11907)
    );

    bfr new_Jinkela_buffer_16667 (
        .din(new_Jinkela_wire_19875),
        .dout(new_Jinkela_wire_19876)
    );

    bfr new_Jinkela_buffer_6361 (
        .din(new_Jinkela_wire_8048),
        .dout(new_Jinkela_wire_8049)
    );

    bfr new_Jinkela_buffer_9874 (
        .din(new_Jinkela_wire_11993),
        .dout(new_Jinkela_wire_11994)
    );

    bfr new_Jinkela_buffer_16752 (
        .din(new_Jinkela_wire_19988),
        .dout(new_Jinkela_wire_19989)
    );

    spl2 new_Jinkela_splitter_686 (
        .a(new_Jinkela_wire_7967),
        .b(new_Jinkela_wire_7968),
        .c(new_Jinkela_wire_7969)
    );

    bfr new_Jinkela_buffer_9798 (
        .din(new_Jinkela_wire_11907),
        .dout(new_Jinkela_wire_11908)
    );

    bfr new_Jinkela_buffer_16668 (
        .din(new_Jinkela_wire_19876),
        .dout(new_Jinkela_wire_19877)
    );

    bfr new_Jinkela_buffer_6362 (
        .din(new_Jinkela_wire_8049),
        .dout(new_Jinkela_wire_8050)
    );

    bfr new_Jinkela_buffer_9937 (
        .din(new_Jinkela_wire_12076),
        .dout(new_Jinkela_wire_12077)
    );

    bfr new_Jinkela_buffer_16807 (
        .din(new_Jinkela_wire_20053),
        .dout(new_Jinkela_wire_20054)
    );

    bfr new_Jinkela_buffer_9799 (
        .din(new_Jinkela_wire_11908),
        .dout(new_Jinkela_wire_11909)
    );

    bfr new_Jinkela_buffer_16669 (
        .din(new_Jinkela_wire_19877),
        .dout(new_Jinkela_wire_19878)
    );

    bfr new_Jinkela_buffer_6507 (
        .din(_1597_),
        .dout(new_Jinkela_wire_8207)
    );

    bfr new_Jinkela_buffer_6417 (
        .din(new_Jinkela_wire_8108),
        .dout(new_Jinkela_wire_8109)
    );

    bfr new_Jinkela_buffer_9875 (
        .din(new_Jinkela_wire_11994),
        .dout(new_Jinkela_wire_11995)
    );

    bfr new_Jinkela_buffer_16753 (
        .din(new_Jinkela_wire_19989),
        .dout(new_Jinkela_wire_19990)
    );

    bfr new_Jinkela_buffer_6363 (
        .din(new_Jinkela_wire_8050),
        .dout(new_Jinkela_wire_8051)
    );

    bfr new_Jinkela_buffer_9800 (
        .din(new_Jinkela_wire_11909),
        .dout(new_Jinkela_wire_11910)
    );

    bfr new_Jinkela_buffer_16670 (
        .din(new_Jinkela_wire_19878),
        .dout(new_Jinkela_wire_19879)
    );

    spl2 new_Jinkela_splitter_1474 (
        .a(_1097_),
        .b(new_Jinkela_wire_20142),
        .c(new_Jinkela_wire_20143)
    );

    bfr new_Jinkela_buffer_6488 (
        .din(new_Jinkela_wire_8187),
        .dout(new_Jinkela_wire_8188)
    );

    bfr new_Jinkela_buffer_9967 (
        .din(new_Jinkela_wire_12112),
        .dout(new_Jinkela_wire_12113)
    );

    bfr new_Jinkela_buffer_16887 (
        .din(new_Jinkela_wire_20137),
        .dout(new_Jinkela_wire_20138)
    );

    bfr new_Jinkela_buffer_6364 (
        .din(new_Jinkela_wire_8051),
        .dout(new_Jinkela_wire_8052)
    );

    bfr new_Jinkela_buffer_9801 (
        .din(new_Jinkela_wire_11910),
        .dout(new_Jinkela_wire_11911)
    );

    bfr new_Jinkela_buffer_16671 (
        .din(new_Jinkela_wire_19879),
        .dout(new_Jinkela_wire_19880)
    );

    bfr new_Jinkela_buffer_6418 (
        .din(new_Jinkela_wire_8109),
        .dout(new_Jinkela_wire_8110)
    );

    bfr new_Jinkela_buffer_9876 (
        .din(new_Jinkela_wire_11995),
        .dout(new_Jinkela_wire_11996)
    );

    bfr new_Jinkela_buffer_16754 (
        .din(new_Jinkela_wire_19990),
        .dout(new_Jinkela_wire_19991)
    );

    bfr new_Jinkela_buffer_6365 (
        .din(new_Jinkela_wire_8052),
        .dout(new_Jinkela_wire_8053)
    );

    bfr new_Jinkela_buffer_9802 (
        .din(new_Jinkela_wire_11911),
        .dout(new_Jinkela_wire_11912)
    );

    bfr new_Jinkela_buffer_16672 (
        .din(new_Jinkela_wire_19880),
        .dout(new_Jinkela_wire_19881)
    );

    bfr new_Jinkela_buffer_9938 (
        .din(new_Jinkela_wire_12077),
        .dout(new_Jinkela_wire_12078)
    );

    bfr new_Jinkela_buffer_16808 (
        .din(new_Jinkela_wire_20054),
        .dout(new_Jinkela_wire_20055)
    );

    bfr new_Jinkela_buffer_6508 (
        .din(_1774_),
        .dout(new_Jinkela_wire_8208)
    );

    bfr new_Jinkela_buffer_6366 (
        .din(new_Jinkela_wire_8053),
        .dout(new_Jinkela_wire_8054)
    );

    bfr new_Jinkela_buffer_9803 (
        .din(new_Jinkela_wire_11912),
        .dout(new_Jinkela_wire_11913)
    );

    bfr new_Jinkela_buffer_16673 (
        .din(new_Jinkela_wire_19881),
        .dout(new_Jinkela_wire_19882)
    );

    bfr new_Jinkela_buffer_6419 (
        .din(new_Jinkela_wire_8110),
        .dout(new_Jinkela_wire_8111)
    );

    bfr new_Jinkela_buffer_9877 (
        .din(new_Jinkela_wire_11996),
        .dout(new_Jinkela_wire_11997)
    );

    bfr new_Jinkela_buffer_16755 (
        .din(new_Jinkela_wire_19991),
        .dout(new_Jinkela_wire_19992)
    );

    bfr new_Jinkela_buffer_6367 (
        .din(new_Jinkela_wire_8054),
        .dout(new_Jinkela_wire_8055)
    );

    bfr new_Jinkela_buffer_9804 (
        .din(new_Jinkela_wire_11913),
        .dout(new_Jinkela_wire_11914)
    );

    bfr new_Jinkela_buffer_16674 (
        .din(new_Jinkela_wire_19882),
        .dout(new_Jinkela_wire_19883)
    );

    bfr new_Jinkela_buffer_9964 (
        .din(new_Jinkela_wire_12109),
        .dout(new_Jinkela_wire_12110)
    );

    bfr new_Jinkela_buffer_6489 (
        .din(new_Jinkela_wire_8188),
        .dout(new_Jinkela_wire_8189)
    );

    bfr new_Jinkela_buffer_6368 (
        .din(new_Jinkela_wire_8055),
        .dout(new_Jinkela_wire_8056)
    );

    bfr new_Jinkela_buffer_9805 (
        .din(new_Jinkela_wire_11914),
        .dout(new_Jinkela_wire_11915)
    );

    bfr new_Jinkela_buffer_16675 (
        .din(new_Jinkela_wire_19883),
        .dout(new_Jinkela_wire_19884)
    );

    bfr new_Jinkela_buffer_6420 (
        .din(new_Jinkela_wire_8111),
        .dout(new_Jinkela_wire_8112)
    );

    bfr new_Jinkela_buffer_9878 (
        .din(new_Jinkela_wire_11997),
        .dout(new_Jinkela_wire_11998)
    );

    bfr new_Jinkela_buffer_16756 (
        .din(new_Jinkela_wire_19992),
        .dout(new_Jinkela_wire_19993)
    );

    bfr new_Jinkela_buffer_6369 (
        .din(new_Jinkela_wire_8056),
        .dout(new_Jinkela_wire_8057)
    );

    bfr new_Jinkela_buffer_9806 (
        .din(new_Jinkela_wire_11915),
        .dout(new_Jinkela_wire_11916)
    );

    bfr new_Jinkela_buffer_16676 (
        .din(new_Jinkela_wire_19884),
        .dout(new_Jinkela_wire_19885)
    );

    bfr new_Jinkela_buffer_9939 (
        .din(new_Jinkela_wire_12078),
        .dout(new_Jinkela_wire_12079)
    );

    bfr new_Jinkela_buffer_16809 (
        .din(new_Jinkela_wire_20055),
        .dout(new_Jinkela_wire_20056)
    );

    bfr new_Jinkela_buffer_6509 (
        .din(_1461_),
        .dout(new_Jinkela_wire_8209)
    );

    bfr new_Jinkela_buffer_6370 (
        .din(new_Jinkela_wire_8057),
        .dout(new_Jinkela_wire_8058)
    );

    bfr new_Jinkela_buffer_9807 (
        .din(new_Jinkela_wire_11916),
        .dout(new_Jinkela_wire_11917)
    );

    bfr new_Jinkela_buffer_16677 (
        .din(new_Jinkela_wire_19885),
        .dout(new_Jinkela_wire_19886)
    );

    bfr new_Jinkela_buffer_6421 (
        .din(new_Jinkela_wire_8112),
        .dout(new_Jinkela_wire_8113)
    );

    bfr new_Jinkela_buffer_9879 (
        .din(new_Jinkela_wire_11998),
        .dout(new_Jinkela_wire_11999)
    );

    bfr new_Jinkela_buffer_16757 (
        .din(new_Jinkela_wire_19993),
        .dout(new_Jinkela_wire_19994)
    );

    bfr new_Jinkela_buffer_6371 (
        .din(new_Jinkela_wire_8058),
        .dout(new_Jinkela_wire_8059)
    );

    bfr new_Jinkela_buffer_9808 (
        .din(new_Jinkela_wire_11917),
        .dout(new_Jinkela_wire_11918)
    );

    bfr new_Jinkela_buffer_16678 (
        .din(new_Jinkela_wire_19886),
        .dout(new_Jinkela_wire_19887)
    );

    spl2 new_Jinkela_splitter_700 (
        .a(_1165_),
        .b(new_Jinkela_wire_8276),
        .c(new_Jinkela_wire_8277)
    );

    bfr new_Jinkela_buffer_6490 (
        .din(new_Jinkela_wire_8189),
        .dout(new_Jinkela_wire_8190)
    );

    spl2 new_Jinkela_splitter_925 (
        .a(_0952_),
        .b(new_Jinkela_wire_12329),
        .c(new_Jinkela_wire_12330)
    );

    bfr new_Jinkela_buffer_16891 (
        .din(_0225_),
        .dout(new_Jinkela_wire_20144)
    );

    bfr new_Jinkela_buffer_6372 (
        .din(new_Jinkela_wire_8059),
        .dout(new_Jinkela_wire_8060)
    );

    bfr new_Jinkela_buffer_9809 (
        .din(new_Jinkela_wire_11918),
        .dout(new_Jinkela_wire_11919)
    );

    bfr new_Jinkela_buffer_16679 (
        .din(new_Jinkela_wire_19887),
        .dout(new_Jinkela_wire_19888)
    );

    bfr new_Jinkela_buffer_6422 (
        .din(new_Jinkela_wire_8113),
        .dout(new_Jinkela_wire_8114)
    );

    bfr new_Jinkela_buffer_9880 (
        .din(new_Jinkela_wire_11999),
        .dout(new_Jinkela_wire_12000)
    );

    bfr new_Jinkela_buffer_16758 (
        .din(new_Jinkela_wire_19994),
        .dout(new_Jinkela_wire_19995)
    );

    bfr new_Jinkela_buffer_6373 (
        .din(new_Jinkela_wire_8060),
        .dout(new_Jinkela_wire_8061)
    );

    bfr new_Jinkela_buffer_9810 (
        .din(new_Jinkela_wire_11919),
        .dout(new_Jinkela_wire_11920)
    );

    bfr new_Jinkela_buffer_16680 (
        .din(new_Jinkela_wire_19888),
        .dout(new_Jinkela_wire_19889)
    );

    bfr new_Jinkela_buffer_9940 (
        .din(new_Jinkela_wire_12079),
        .dout(new_Jinkela_wire_12080)
    );

    bfr new_Jinkela_buffer_16810 (
        .din(new_Jinkela_wire_20056),
        .dout(new_Jinkela_wire_20057)
    );

    bfr new_Jinkela_buffer_6374 (
        .din(new_Jinkela_wire_8061),
        .dout(new_Jinkela_wire_8062)
    );

    bfr new_Jinkela_buffer_9811 (
        .din(new_Jinkela_wire_11920),
        .dout(new_Jinkela_wire_11921)
    );

    bfr new_Jinkela_buffer_16681 (
        .din(new_Jinkela_wire_19889),
        .dout(new_Jinkela_wire_19890)
    );

    bfr new_Jinkela_buffer_6423 (
        .din(new_Jinkela_wire_8114),
        .dout(new_Jinkela_wire_8115)
    );

    bfr new_Jinkela_buffer_9881 (
        .din(new_Jinkela_wire_12000),
        .dout(new_Jinkela_wire_12001)
    );

    bfr new_Jinkela_buffer_16759 (
        .din(new_Jinkela_wire_19995),
        .dout(new_Jinkela_wire_19996)
    );

    spl2 new_Jinkela_splitter_1157 (
        .a(_1616_),
        .b(new_Jinkela_wire_16102),
        .c(new_Jinkela_wire_16103)
    );

    bfr new_Jinkela_buffer_13292 (
        .din(new_Jinkela_wire_15891),
        .dout(new_Jinkela_wire_15892)
    );

    bfr new_Jinkela_buffer_13328 (
        .din(new_Jinkela_wire_15929),
        .dout(new_Jinkela_wire_15930)
    );

    spl2 new_Jinkela_splitter_1158 (
        .a(_0685_),
        .b(new_Jinkela_wire_16104),
        .c(new_Jinkela_wire_16105)
    );

    bfr new_Jinkela_buffer_13329 (
        .din(new_Jinkela_wire_15930),
        .dout(new_Jinkela_wire_15931)
    );

    bfr new_Jinkela_buffer_13399 (
        .din(new_Jinkela_wire_16012),
        .dout(new_Jinkela_wire_16013)
    );

    bfr new_Jinkela_buffer_13330 (
        .din(new_Jinkela_wire_15931),
        .dout(new_Jinkela_wire_15932)
    );

    bfr new_Jinkela_buffer_13331 (
        .din(new_Jinkela_wire_15932),
        .dout(new_Jinkela_wire_15933)
    );

    bfr new_Jinkela_buffer_13400 (
        .din(new_Jinkela_wire_16013),
        .dout(new_Jinkela_wire_16014)
    );

    bfr new_Jinkela_buffer_13332 (
        .din(new_Jinkela_wire_15933),
        .dout(new_Jinkela_wire_15934)
    );

    spl2 new_Jinkela_splitter_1159 (
        .a(_1556_),
        .b(new_Jinkela_wire_16106),
        .c(new_Jinkela_wire_16107)
    );

    bfr new_Jinkela_buffer_13333 (
        .din(new_Jinkela_wire_15934),
        .dout(new_Jinkela_wire_15935)
    );

    bfr new_Jinkela_buffer_13401 (
        .din(new_Jinkela_wire_16014),
        .dout(new_Jinkela_wire_16015)
    );

    bfr new_Jinkela_buffer_13334 (
        .din(new_Jinkela_wire_15935),
        .dout(new_Jinkela_wire_15936)
    );

    spl2 new_Jinkela_splitter_1161 (
        .a(_1127_),
        .b(new_Jinkela_wire_16111),
        .c(new_Jinkela_wire_16112)
    );

    bfr new_Jinkela_buffer_13335 (
        .din(new_Jinkela_wire_15936),
        .dout(new_Jinkela_wire_15937)
    );

    bfr new_Jinkela_buffer_13402 (
        .din(new_Jinkela_wire_16015),
        .dout(new_Jinkela_wire_16016)
    );

    bfr new_Jinkela_buffer_13336 (
        .din(new_Jinkela_wire_15937),
        .dout(new_Jinkela_wire_15938)
    );

    bfr new_Jinkela_buffer_13486 (
        .din(new_Jinkela_wire_16107),
        .dout(new_Jinkela_wire_16108)
    );

    bfr new_Jinkela_buffer_13487 (
        .din(_0201_),
        .dout(new_Jinkela_wire_16113)
    );

    bfr new_Jinkela_buffer_13337 (
        .din(new_Jinkela_wire_15938),
        .dout(new_Jinkela_wire_15939)
    );

    bfr new_Jinkela_buffer_13403 (
        .din(new_Jinkela_wire_16016),
        .dout(new_Jinkela_wire_16017)
    );

    bfr new_Jinkela_buffer_13338 (
        .din(new_Jinkela_wire_15939),
        .dout(new_Jinkela_wire_15940)
    );

    spl2 new_Jinkela_splitter_1162 (
        .a(_0261_),
        .b(new_Jinkela_wire_16114),
        .c(new_Jinkela_wire_16115)
    );

    bfr new_Jinkela_buffer_13339 (
        .din(new_Jinkela_wire_15940),
        .dout(new_Jinkela_wire_15941)
    );

    bfr new_Jinkela_buffer_13404 (
        .din(new_Jinkela_wire_16017),
        .dout(new_Jinkela_wire_16018)
    );

    bfr new_Jinkela_buffer_13340 (
        .din(new_Jinkela_wire_15941),
        .dout(new_Jinkela_wire_15942)
    );

    spl2 new_Jinkela_splitter_1163 (
        .a(_0372_),
        .b(new_Jinkela_wire_16116),
        .c(new_Jinkela_wire_16117)
    );

    spl2 new_Jinkela_splitter_1160 (
        .a(new_Jinkela_wire_16108),
        .b(new_Jinkela_wire_16109),
        .c(new_Jinkela_wire_16110)
    );

    bfr new_Jinkela_buffer_13341 (
        .din(new_Jinkela_wire_15942),
        .dout(new_Jinkela_wire_15943)
    );

    bfr new_Jinkela_buffer_13405 (
        .din(new_Jinkela_wire_16018),
        .dout(new_Jinkela_wire_16019)
    );

    bfr new_Jinkela_buffer_13342 (
        .din(new_Jinkela_wire_15943),
        .dout(new_Jinkela_wire_15944)
    );

    bfr new_Jinkela_buffer_13343 (
        .din(new_Jinkela_wire_15944),
        .dout(new_Jinkela_wire_15945)
    );

    bfr new_Jinkela_buffer_13406 (
        .din(new_Jinkela_wire_16019),
        .dout(new_Jinkela_wire_16020)
    );

    bfr new_Jinkela_buffer_13344 (
        .din(new_Jinkela_wire_15945),
        .dout(new_Jinkela_wire_15946)
    );

    bfr new_Jinkela_buffer_13488 (
        .din(_1188_),
        .dout(new_Jinkela_wire_16120)
    );

    bfr new_Jinkela_buffer_13345 (
        .din(new_Jinkela_wire_15946),
        .dout(new_Jinkela_wire_15947)
    );

    bfr new_Jinkela_buffer_13407 (
        .din(new_Jinkela_wire_16020),
        .dout(new_Jinkela_wire_16021)
    );

    bfr new_Jinkela_buffer_13346 (
        .din(new_Jinkela_wire_15947),
        .dout(new_Jinkela_wire_15948)
    );

    spl2 new_Jinkela_splitter_1164 (
        .a(_1355_),
        .b(new_Jinkela_wire_16118),
        .c(new_Jinkela_wire_16119)
    );

    bfr new_Jinkela_buffer_13347 (
        .din(new_Jinkela_wire_15948),
        .dout(new_Jinkela_wire_15949)
    );

    bfr new_Jinkela_buffer_13408 (
        .din(new_Jinkela_wire_16021),
        .dout(new_Jinkela_wire_16022)
    );

    bfr new_Jinkela_buffer_13398 (
        .din(_0333_),
        .dout(new_Jinkela_wire_16012)
    );

    bfr new_Jinkela_buffer_9812 (
        .din(new_Jinkela_wire_11921),
        .dout(new_Jinkela_wire_11922)
    );

    bfr new_Jinkela_buffer_3082 (
        .din(new_Jinkela_wire_4171),
        .dout(new_Jinkela_wire_4172)
    );

    bfr new_Jinkela_buffer_16682 (
        .din(new_Jinkela_wire_19890),
        .dout(new_Jinkela_wire_19891)
    );

    bfr new_Jinkela_buffer_10026 (
        .din(new_Jinkela_wire_12171),
        .dout(new_Jinkela_wire_12172)
    );

    bfr new_Jinkela_buffer_2937 (
        .din(new_Jinkela_wire_4008),
        .dout(new_Jinkela_wire_4009)
    );

    bfr new_Jinkela_buffer_9968 (
        .din(new_Jinkela_wire_12113),
        .dout(new_Jinkela_wire_12114)
    );

    bfr new_Jinkela_buffer_16959 (
        .din(_0594_),
        .dout(new_Jinkela_wire_20216)
    );

    bfr new_Jinkela_buffer_9813 (
        .din(new_Jinkela_wire_11922),
        .dout(new_Jinkela_wire_11923)
    );

    bfr new_Jinkela_buffer_3020 (
        .din(new_Jinkela_wire_4101),
        .dout(new_Jinkela_wire_4102)
    );

    bfr new_Jinkela_buffer_16683 (
        .din(new_Jinkela_wire_19891),
        .dout(new_Jinkela_wire_19892)
    );

    bfr new_Jinkela_buffer_9882 (
        .din(new_Jinkela_wire_12001),
        .dout(new_Jinkela_wire_12002)
    );

    bfr new_Jinkela_buffer_2938 (
        .din(new_Jinkela_wire_4009),
        .dout(new_Jinkela_wire_4010)
    );

    bfr new_Jinkela_buffer_16760 (
        .din(new_Jinkela_wire_19996),
        .dout(new_Jinkela_wire_19997)
    );

    bfr new_Jinkela_buffer_16684 (
        .din(new_Jinkela_wire_19892),
        .dout(new_Jinkela_wire_19893)
    );

    bfr new_Jinkela_buffer_9814 (
        .din(new_Jinkela_wire_11923),
        .dout(new_Jinkela_wire_11924)
    );

    spl2 new_Jinkela_splitter_399 (
        .a(_0503_),
        .b(new_Jinkela_wire_4249),
        .c(new_Jinkela_wire_4250)
    );

    bfr new_Jinkela_buffer_9941 (
        .din(new_Jinkela_wire_12080),
        .dout(new_Jinkela_wire_12081)
    );

    bfr new_Jinkela_buffer_2939 (
        .din(new_Jinkela_wire_4010),
        .dout(new_Jinkela_wire_4011)
    );

    bfr new_Jinkela_buffer_16811 (
        .din(new_Jinkela_wire_20057),
        .dout(new_Jinkela_wire_20058)
    );

    bfr new_Jinkela_buffer_9815 (
        .din(new_Jinkela_wire_11924),
        .dout(new_Jinkela_wire_11925)
    );

    bfr new_Jinkela_buffer_3021 (
        .din(new_Jinkela_wire_4102),
        .dout(new_Jinkela_wire_4103)
    );

    bfr new_Jinkela_buffer_16685 (
        .din(new_Jinkela_wire_19893),
        .dout(new_Jinkela_wire_19894)
    );

    bfr new_Jinkela_buffer_9883 (
        .din(new_Jinkela_wire_12002),
        .dout(new_Jinkela_wire_12003)
    );

    bfr new_Jinkela_buffer_2940 (
        .din(new_Jinkela_wire_4011),
        .dout(new_Jinkela_wire_4012)
    );

    bfr new_Jinkela_buffer_16761 (
        .din(new_Jinkela_wire_19997),
        .dout(new_Jinkela_wire_19998)
    );

    bfr new_Jinkela_buffer_9816 (
        .din(new_Jinkela_wire_11925),
        .dout(new_Jinkela_wire_11926)
    );

    bfr new_Jinkela_buffer_3083 (
        .din(new_Jinkela_wire_4172),
        .dout(new_Jinkela_wire_4173)
    );

    bfr new_Jinkela_buffer_16686 (
        .din(new_Jinkela_wire_19894),
        .dout(new_Jinkela_wire_19895)
    );

    bfr new_Jinkela_buffer_16888 (
        .din(new_Jinkela_wire_20138),
        .dout(new_Jinkela_wire_20139)
    );

    bfr new_Jinkela_buffer_2941 (
        .din(new_Jinkela_wire_4012),
        .dout(new_Jinkela_wire_4013)
    );

    bfr new_Jinkela_buffer_9817 (
        .din(new_Jinkela_wire_11926),
        .dout(new_Jinkela_wire_11927)
    );

    bfr new_Jinkela_buffer_3022 (
        .din(new_Jinkela_wire_4103),
        .dout(new_Jinkela_wire_4104)
    );

    bfr new_Jinkela_buffer_16687 (
        .din(new_Jinkela_wire_19895),
        .dout(new_Jinkela_wire_19896)
    );

    bfr new_Jinkela_buffer_9884 (
        .din(new_Jinkela_wire_12003),
        .dout(new_Jinkela_wire_12004)
    );

    bfr new_Jinkela_buffer_2942 (
        .din(new_Jinkela_wire_4013),
        .dout(new_Jinkela_wire_4014)
    );

    bfr new_Jinkela_buffer_16762 (
        .din(new_Jinkela_wire_19998),
        .dout(new_Jinkela_wire_19999)
    );

    bfr new_Jinkela_buffer_9818 (
        .din(new_Jinkela_wire_11927),
        .dout(new_Jinkela_wire_11928)
    );

    spl2 new_Jinkela_splitter_400 (
        .a(_1767_),
        .b(new_Jinkela_wire_4251),
        .c(new_Jinkela_wire_4252)
    );

    bfr new_Jinkela_buffer_16688 (
        .din(new_Jinkela_wire_19896),
        .dout(new_Jinkela_wire_19897)
    );

    bfr new_Jinkela_buffer_3150 (
        .din(new_Jinkela_wire_4253),
        .dout(new_Jinkela_wire_4254)
    );

    bfr new_Jinkela_buffer_9942 (
        .din(new_Jinkela_wire_12081),
        .dout(new_Jinkela_wire_12082)
    );

    bfr new_Jinkela_buffer_2943 (
        .din(new_Jinkela_wire_4014),
        .dout(new_Jinkela_wire_4015)
    );

    bfr new_Jinkela_buffer_16812 (
        .din(new_Jinkela_wire_20058),
        .dout(new_Jinkela_wire_20059)
    );

    bfr new_Jinkela_buffer_9819 (
        .din(new_Jinkela_wire_11928),
        .dout(new_Jinkela_wire_11929)
    );

    bfr new_Jinkela_buffer_3023 (
        .din(new_Jinkela_wire_4104),
        .dout(new_Jinkela_wire_4105)
    );

    bfr new_Jinkela_buffer_16689 (
        .din(new_Jinkela_wire_19897),
        .dout(new_Jinkela_wire_19898)
    );

    bfr new_Jinkela_buffer_9885 (
        .din(new_Jinkela_wire_12004),
        .dout(new_Jinkela_wire_12005)
    );

    bfr new_Jinkela_buffer_2944 (
        .din(new_Jinkela_wire_4015),
        .dout(new_Jinkela_wire_4016)
    );

    bfr new_Jinkela_buffer_16763 (
        .din(new_Jinkela_wire_19999),
        .dout(new_Jinkela_wire_20000)
    );

    bfr new_Jinkela_buffer_9820 (
        .din(new_Jinkela_wire_11929),
        .dout(new_Jinkela_wire_11930)
    );

    bfr new_Jinkela_buffer_3084 (
        .din(new_Jinkela_wire_4173),
        .dout(new_Jinkela_wire_4174)
    );

    bfr new_Jinkela_buffer_16690 (
        .din(new_Jinkela_wire_19898),
        .dout(new_Jinkela_wire_19899)
    );

    bfr new_Jinkela_buffer_10073 (
        .din(_0769_),
        .dout(new_Jinkela_wire_12223)
    );

    bfr new_Jinkela_buffer_2945 (
        .din(new_Jinkela_wire_4016),
        .dout(new_Jinkela_wire_4017)
    );

    bfr new_Jinkela_buffer_9969 (
        .din(new_Jinkela_wire_12114),
        .dout(new_Jinkela_wire_12115)
    );

    spl2 new_Jinkela_splitter_1476 (
        .a(_0861_),
        .b(new_Jinkela_wire_20210),
        .c(new_Jinkela_wire_20211)
    );

    bfr new_Jinkela_buffer_9821 (
        .din(new_Jinkela_wire_11930),
        .dout(new_Jinkela_wire_11931)
    );

    bfr new_Jinkela_buffer_3024 (
        .din(new_Jinkela_wire_4105),
        .dout(new_Jinkela_wire_4106)
    );

    bfr new_Jinkela_buffer_16691 (
        .din(new_Jinkela_wire_19899),
        .dout(new_Jinkela_wire_19900)
    );

    bfr new_Jinkela_buffer_9886 (
        .din(new_Jinkela_wire_12005),
        .dout(new_Jinkela_wire_12006)
    );

    bfr new_Jinkela_buffer_2946 (
        .din(new_Jinkela_wire_4017),
        .dout(new_Jinkela_wire_4018)
    );

    bfr new_Jinkela_buffer_16764 (
        .din(new_Jinkela_wire_20000),
        .dout(new_Jinkela_wire_20001)
    );

    bfr new_Jinkela_buffer_16692 (
        .din(new_Jinkela_wire_19900),
        .dout(new_Jinkela_wire_19901)
    );

    bfr new_Jinkela_buffer_9822 (
        .din(new_Jinkela_wire_11931),
        .dout(new_Jinkela_wire_11932)
    );

    bfr new_Jinkela_buffer_9943 (
        .din(new_Jinkela_wire_12082),
        .dout(new_Jinkela_wire_12083)
    );

    bfr new_Jinkela_buffer_2947 (
        .din(new_Jinkela_wire_4018),
        .dout(new_Jinkela_wire_4019)
    );

    bfr new_Jinkela_buffer_16813 (
        .din(new_Jinkela_wire_20059),
        .dout(new_Jinkela_wire_20060)
    );

    bfr new_Jinkela_buffer_9823 (
        .din(new_Jinkela_wire_11932),
        .dout(new_Jinkela_wire_11933)
    );

    bfr new_Jinkela_buffer_3025 (
        .din(new_Jinkela_wire_4106),
        .dout(new_Jinkela_wire_4107)
    );

    bfr new_Jinkela_buffer_16693 (
        .din(new_Jinkela_wire_19901),
        .dout(new_Jinkela_wire_19902)
    );

    bfr new_Jinkela_buffer_9887 (
        .din(new_Jinkela_wire_12006),
        .dout(new_Jinkela_wire_12007)
    );

    bfr new_Jinkela_buffer_2948 (
        .din(new_Jinkela_wire_4019),
        .dout(new_Jinkela_wire_4020)
    );

    bfr new_Jinkela_buffer_16765 (
        .din(new_Jinkela_wire_20001),
        .dout(new_Jinkela_wire_20002)
    );

    bfr new_Jinkela_buffer_9824 (
        .din(new_Jinkela_wire_11933),
        .dout(new_Jinkela_wire_11934)
    );

    bfr new_Jinkela_buffer_3085 (
        .din(new_Jinkela_wire_4174),
        .dout(new_Jinkela_wire_4175)
    );

    bfr new_Jinkela_buffer_16694 (
        .din(new_Jinkela_wire_19902),
        .dout(new_Jinkela_wire_19903)
    );

    bfr new_Jinkela_buffer_16889 (
        .din(new_Jinkela_wire_20139),
        .dout(new_Jinkela_wire_20140)
    );

    bfr new_Jinkela_buffer_2949 (
        .din(new_Jinkela_wire_4020),
        .dout(new_Jinkela_wire_4021)
    );

    bfr new_Jinkela_buffer_9825 (
        .din(new_Jinkela_wire_11934),
        .dout(new_Jinkela_wire_11935)
    );

    bfr new_Jinkela_buffer_3026 (
        .din(new_Jinkela_wire_4107),
        .dout(new_Jinkela_wire_4108)
    );

    bfr new_Jinkela_buffer_16695 (
        .din(new_Jinkela_wire_19903),
        .dout(new_Jinkela_wire_19904)
    );

    bfr new_Jinkela_buffer_9888 (
        .din(new_Jinkela_wire_12007),
        .dout(new_Jinkela_wire_12008)
    );

    bfr new_Jinkela_buffer_2950 (
        .din(new_Jinkela_wire_4021),
        .dout(new_Jinkela_wire_4022)
    );

    bfr new_Jinkela_buffer_16766 (
        .din(new_Jinkela_wire_20002),
        .dout(new_Jinkela_wire_20003)
    );

    bfr new_Jinkela_buffer_16696 (
        .din(new_Jinkela_wire_19904),
        .dout(new_Jinkela_wire_19905)
    );

    bfr new_Jinkela_buffer_9826 (
        .din(new_Jinkela_wire_11935),
        .dout(new_Jinkela_wire_11936)
    );

    bfr new_Jinkela_buffer_3149 (
        .din(new_net_3948),
        .dout(new_Jinkela_wire_4253)
    );

    bfr new_Jinkela_buffer_9944 (
        .din(new_Jinkela_wire_12083),
        .dout(new_Jinkela_wire_12084)
    );

    bfr new_Jinkela_buffer_2951 (
        .din(new_Jinkela_wire_4022),
        .dout(new_Jinkela_wire_4023)
    );

    bfr new_Jinkela_buffer_16814 (
        .din(new_Jinkela_wire_20060),
        .dout(new_Jinkela_wire_20061)
    );

    bfr new_Jinkela_buffer_9827 (
        .din(new_Jinkela_wire_11936),
        .dout(new_Jinkela_wire_11937)
    );

    bfr new_Jinkela_buffer_3027 (
        .din(new_Jinkela_wire_4108),
        .dout(new_Jinkela_wire_4109)
    );

    spl2 new_Jinkela_splitter_1453 (
        .a(new_Jinkela_wire_19905),
        .b(new_Jinkela_wire_19906),
        .c(new_Jinkela_wire_19907)
    );

    bfr new_Jinkela_buffer_9889 (
        .din(new_Jinkela_wire_12008),
        .dout(new_Jinkela_wire_12009)
    );

    bfr new_Jinkela_buffer_2952 (
        .din(new_Jinkela_wire_4023),
        .dout(new_Jinkela_wire_4024)
    );

    bfr new_Jinkela_buffer_16892 (
        .din(new_Jinkela_wire_20144),
        .dout(new_Jinkela_wire_20145)
    );

    bfr new_Jinkela_buffer_9828 (
        .din(new_Jinkela_wire_11937),
        .dout(new_Jinkela_wire_11938)
    );

    bfr new_Jinkela_buffer_3086 (
        .din(new_Jinkela_wire_4175),
        .dout(new_Jinkela_wire_4176)
    );

    bfr new_Jinkela_buffer_16767 (
        .din(new_Jinkela_wire_20003),
        .dout(new_Jinkela_wire_20004)
    );

    bfr new_Jinkela_buffer_10027 (
        .din(new_Jinkela_wire_12172),
        .dout(new_Jinkela_wire_12173)
    );

    bfr new_Jinkela_buffer_2953 (
        .din(new_Jinkela_wire_4024),
        .dout(new_Jinkela_wire_4025)
    );

    bfr new_Jinkela_buffer_16768 (
        .din(new_Jinkela_wire_20004),
        .dout(new_Jinkela_wire_20005)
    );

    bfr new_Jinkela_buffer_9970 (
        .din(new_Jinkela_wire_12115),
        .dout(new_Jinkela_wire_12116)
    );

    bfr new_Jinkela_buffer_9829 (
        .din(new_Jinkela_wire_11938),
        .dout(new_Jinkela_wire_11939)
    );

    bfr new_Jinkela_buffer_3028 (
        .din(new_Jinkela_wire_4109),
        .dout(new_Jinkela_wire_4110)
    );

    bfr new_Jinkela_buffer_16815 (
        .din(new_Jinkela_wire_20061),
        .dout(new_Jinkela_wire_20062)
    );

    bfr new_Jinkela_buffer_9890 (
        .din(new_Jinkela_wire_12009),
        .dout(new_Jinkela_wire_12010)
    );

    bfr new_Jinkela_buffer_2954 (
        .din(new_Jinkela_wire_4025),
        .dout(new_Jinkela_wire_4026)
    );

    bfr new_Jinkela_buffer_16769 (
        .din(new_Jinkela_wire_20005),
        .dout(new_Jinkela_wire_20006)
    );

    bfr new_Jinkela_buffer_9830 (
        .din(new_Jinkela_wire_11939),
        .dout(new_Jinkela_wire_11940)
    );

    spl2 new_Jinkela_splitter_402 (
        .a(_0428_),
        .b(new_Jinkela_wire_4283),
        .c(new_Jinkela_wire_4284)
    );

    bfr new_Jinkela_buffer_16890 (
        .din(new_Jinkela_wire_20140),
        .dout(new_Jinkela_wire_20141)
    );

    bfr new_Jinkela_buffer_3161 (
        .din(_0709_),
        .dout(new_Jinkela_wire_4265)
    );

    bfr new_Jinkela_buffer_9945 (
        .din(new_Jinkela_wire_12084),
        .dout(new_Jinkela_wire_12085)
    );

    bfr new_Jinkela_buffer_2955 (
        .din(new_Jinkela_wire_4026),
        .dout(new_Jinkela_wire_4027)
    );

    bfr new_Jinkela_buffer_16770 (
        .din(new_Jinkela_wire_20006),
        .dout(new_Jinkela_wire_20007)
    );

    bfr new_Jinkela_buffer_9831 (
        .din(new_Jinkela_wire_11940),
        .dout(new_Jinkela_wire_11941)
    );

    bfr new_Jinkela_buffer_3029 (
        .din(new_Jinkela_wire_4110),
        .dout(new_Jinkela_wire_4111)
    );

    bfr new_Jinkela_buffer_16816 (
        .din(new_Jinkela_wire_20062),
        .dout(new_Jinkela_wire_20063)
    );

    bfr new_Jinkela_buffer_9891 (
        .din(new_Jinkela_wire_12010),
        .dout(new_Jinkela_wire_12011)
    );

    bfr new_Jinkela_buffer_2956 (
        .din(new_Jinkela_wire_4027),
        .dout(new_Jinkela_wire_4028)
    );

    bfr new_Jinkela_buffer_16771 (
        .din(new_Jinkela_wire_20007),
        .dout(new_Jinkela_wire_20008)
    );

    bfr new_Jinkela_buffer_9832 (
        .din(new_Jinkela_wire_11941),
        .dout(new_Jinkela_wire_11942)
    );

    bfr new_Jinkela_buffer_3087 (
        .din(new_Jinkela_wire_4176),
        .dout(new_Jinkela_wire_4177)
    );

    bfr new_Jinkela_buffer_16955 (
        .din(new_Jinkela_wire_20211),
        .dout(new_Jinkela_wire_20212)
    );

    bfr new_Jinkela_buffer_16772 (
        .din(new_Jinkela_wire_20008),
        .dout(new_Jinkela_wire_20009)
    );

    bfr new_Jinkela_buffer_2957 (
        .din(new_Jinkela_wire_4028),
        .dout(new_Jinkela_wire_4029)
    );

    and_bb _3055_ (
        .a(new_Jinkela_wire_13721),
        .b(new_Jinkela_wire_829),
        .c(_0310_)
    );

    or_ii _1884_ (
        .a(new_Jinkela_wire_10680),
        .b(new_Jinkela_wire_14204),
        .c(_0121_)
    );

    bfr new_Jinkela_buffer_6375 (
        .din(new_Jinkela_wire_8062),
        .dout(new_Jinkela_wire_8063)
    );

    bfr new_Jinkela_buffer_3030 (
        .din(new_Jinkela_wire_4111),
        .dout(new_Jinkela_wire_4112)
    );

    bfr new_Jinkela_buffer_9833 (
        .din(new_Jinkela_wire_11942),
        .dout(new_Jinkela_wire_11943)
    );

    bfr new_Jinkela_buffer_9892 (
        .din(new_Jinkela_wire_12011),
        .dout(new_Jinkela_wire_12012)
    );

    bfr new_Jinkela_buffer_2958 (
        .din(new_Jinkela_wire_4029),
        .dout(new_Jinkela_wire_4030)
    );

    bfr new_Jinkela_buffer_6491 (
        .din(new_Jinkela_wire_8190),
        .dout(new_Jinkela_wire_8191)
    );

    bfr new_Jinkela_buffer_9834 (
        .din(new_Jinkela_wire_11943),
        .dout(new_Jinkela_wire_11944)
    );

    bfr new_Jinkela_buffer_6376 (
        .din(new_Jinkela_wire_8063),
        .dout(new_Jinkela_wire_8064)
    );

    bfr new_Jinkela_buffer_6424 (
        .din(new_Jinkela_wire_8115),
        .dout(new_Jinkela_wire_8116)
    );

    bfr new_Jinkela_buffer_2959 (
        .din(new_Jinkela_wire_4030),
        .dout(new_Jinkela_wire_4031)
    );

    bfr new_Jinkela_buffer_9946 (
        .din(new_Jinkela_wire_12085),
        .dout(new_Jinkela_wire_12086)
    );

    bfr new_Jinkela_buffer_6377 (
        .din(new_Jinkela_wire_8064),
        .dout(new_Jinkela_wire_8065)
    );

    bfr new_Jinkela_buffer_3031 (
        .din(new_Jinkela_wire_4112),
        .dout(new_Jinkela_wire_4113)
    );

    bfr new_Jinkela_buffer_9835 (
        .din(new_Jinkela_wire_11944),
        .dout(new_Jinkela_wire_11945)
    );

    bfr new_Jinkela_buffer_9893 (
        .din(new_Jinkela_wire_12012),
        .dout(new_Jinkela_wire_12013)
    );

    bfr new_Jinkela_buffer_2960 (
        .din(new_Jinkela_wire_4031),
        .dout(new_Jinkela_wire_4032)
    );

    spl2 new_Jinkela_splitter_701 (
        .a(_1329_),
        .b(new_Jinkela_wire_8278),
        .c(new_Jinkela_wire_8279)
    );

    bfr new_Jinkela_buffer_6378 (
        .din(new_Jinkela_wire_8065),
        .dout(new_Jinkela_wire_8066)
    );

    bfr new_Jinkela_buffer_3088 (
        .din(new_Jinkela_wire_4177),
        .dout(new_Jinkela_wire_4178)
    );

    bfr new_Jinkela_buffer_9836 (
        .din(new_Jinkela_wire_11945),
        .dout(new_Jinkela_wire_11946)
    );

    bfr new_Jinkela_buffer_6425 (
        .din(new_Jinkela_wire_8116),
        .dout(new_Jinkela_wire_8117)
    );

    bfr new_Jinkela_buffer_2961 (
        .din(new_Jinkela_wire_4032),
        .dout(new_Jinkela_wire_4033)
    );

    bfr new_Jinkela_buffer_9971 (
        .din(new_Jinkela_wire_12116),
        .dout(new_Jinkela_wire_12117)
    );

    bfr new_Jinkela_buffer_6379 (
        .din(new_Jinkela_wire_8066),
        .dout(new_Jinkela_wire_8067)
    );

    bfr new_Jinkela_buffer_3032 (
        .din(new_Jinkela_wire_4113),
        .dout(new_Jinkela_wire_4114)
    );

    bfr new_Jinkela_buffer_9837 (
        .din(new_Jinkela_wire_11946),
        .dout(new_Jinkela_wire_11947)
    );

    bfr new_Jinkela_buffer_6510 (
        .din(new_Jinkela_wire_8209),
        .dout(new_Jinkela_wire_8210)
    );

    bfr new_Jinkela_buffer_2962 (
        .din(new_Jinkela_wire_4033),
        .dout(new_Jinkela_wire_4034)
    );

    bfr new_Jinkela_buffer_9894 (
        .din(new_Jinkela_wire_12013),
        .dout(new_Jinkela_wire_12014)
    );

    bfr new_Jinkela_buffer_6492 (
        .din(new_Jinkela_wire_8191),
        .dout(new_Jinkela_wire_8192)
    );

    bfr new_Jinkela_buffer_9838 (
        .din(new_Jinkela_wire_11947),
        .dout(new_Jinkela_wire_11948)
    );

    bfr new_Jinkela_buffer_6380 (
        .din(new_Jinkela_wire_8067),
        .dout(new_Jinkela_wire_8068)
    );

    bfr new_Jinkela_buffer_3151 (
        .din(new_Jinkela_wire_4254),
        .dout(new_Jinkela_wire_4255)
    );

    bfr new_Jinkela_buffer_6426 (
        .din(new_Jinkela_wire_8117),
        .dout(new_Jinkela_wire_8118)
    );

    bfr new_Jinkela_buffer_2963 (
        .din(new_Jinkela_wire_4034),
        .dout(new_Jinkela_wire_4035)
    );

    bfr new_Jinkela_buffer_9947 (
        .din(new_Jinkela_wire_12086),
        .dout(new_Jinkela_wire_12087)
    );

    bfr new_Jinkela_buffer_6381 (
        .din(new_Jinkela_wire_8068),
        .dout(new_Jinkela_wire_8069)
    );

    bfr new_Jinkela_buffer_3033 (
        .din(new_Jinkela_wire_4114),
        .dout(new_Jinkela_wire_4115)
    );

    bfr new_Jinkela_buffer_9839 (
        .din(new_Jinkela_wire_11948),
        .dout(new_Jinkela_wire_11949)
    );

    bfr new_Jinkela_buffer_9895 (
        .din(new_Jinkela_wire_12014),
        .dout(new_Jinkela_wire_12015)
    );

    bfr new_Jinkela_buffer_2964 (
        .din(new_Jinkela_wire_4035),
        .dout(new_Jinkela_wire_4036)
    );

    bfr new_Jinkela_buffer_6382 (
        .din(new_Jinkela_wire_8069),
        .dout(new_Jinkela_wire_8070)
    );

    bfr new_Jinkela_buffer_3089 (
        .din(new_Jinkela_wire_4178),
        .dout(new_Jinkela_wire_4179)
    );

    bfr new_Jinkela_buffer_9840 (
        .din(new_Jinkela_wire_11949),
        .dout(new_Jinkela_wire_11950)
    );

    bfr new_Jinkela_buffer_6427 (
        .din(new_Jinkela_wire_8118),
        .dout(new_Jinkela_wire_8119)
    );

    bfr new_Jinkela_buffer_2965 (
        .din(new_Jinkela_wire_4036),
        .dout(new_Jinkela_wire_4037)
    );

    spl2 new_Jinkela_splitter_926 (
        .a(_1626_),
        .b(new_Jinkela_wire_12331),
        .c(new_Jinkela_wire_12332)
    );

    bfr new_Jinkela_buffer_6383 (
        .din(new_Jinkela_wire_8070),
        .dout(new_Jinkela_wire_8071)
    );

    bfr new_Jinkela_buffer_3034 (
        .din(new_Jinkela_wire_4115),
        .dout(new_Jinkela_wire_4116)
    );

    bfr new_Jinkela_buffer_9841 (
        .din(new_Jinkela_wire_11950),
        .dout(new_Jinkela_wire_11951)
    );

    bfr new_Jinkela_buffer_9896 (
        .din(new_Jinkela_wire_12015),
        .dout(new_Jinkela_wire_12016)
    );

    bfr new_Jinkela_buffer_2966 (
        .din(new_Jinkela_wire_4037),
        .dout(new_Jinkela_wire_4038)
    );

    bfr new_Jinkela_buffer_6493 (
        .din(new_Jinkela_wire_8192),
        .dout(new_Jinkela_wire_8193)
    );

    spl2 new_Jinkela_splitter_904 (
        .a(new_Jinkela_wire_11951),
        .b(new_Jinkela_wire_11952),
        .c(new_Jinkela_wire_11953)
    );

    bfr new_Jinkela_buffer_6384 (
        .din(new_Jinkela_wire_8071),
        .dout(new_Jinkela_wire_8072)
    );

    spl2 new_Jinkela_splitter_403 (
        .a(_1231_),
        .b(new_Jinkela_wire_4285),
        .c(new_Jinkela_wire_4286)
    );

    bfr new_Jinkela_buffer_6428 (
        .din(new_Jinkela_wire_8119),
        .dout(new_Jinkela_wire_8120)
    );

    bfr new_Jinkela_buffer_2967 (
        .din(new_Jinkela_wire_4038),
        .dout(new_Jinkela_wire_4039)
    );

    bfr new_Jinkela_buffer_9897 (
        .din(new_Jinkela_wire_12016),
        .dout(new_Jinkela_wire_12017)
    );

    bfr new_Jinkela_buffer_6385 (
        .din(new_Jinkela_wire_8072),
        .dout(new_Jinkela_wire_8073)
    );

    bfr new_Jinkela_buffer_3035 (
        .din(new_Jinkela_wire_4116),
        .dout(new_Jinkela_wire_4117)
    );

    bfr new_Jinkela_buffer_9948 (
        .din(new_Jinkela_wire_12087),
        .dout(new_Jinkela_wire_12088)
    );

    bfr new_Jinkela_buffer_10028 (
        .din(new_Jinkela_wire_12173),
        .dout(new_Jinkela_wire_12174)
    );

    bfr new_Jinkela_buffer_2968 (
        .din(new_Jinkela_wire_4039),
        .dout(new_Jinkela_wire_4040)
    );

    bfr new_Jinkela_buffer_9972 (
        .din(new_Jinkela_wire_12117),
        .dout(new_Jinkela_wire_12118)
    );

    bfr new_Jinkela_buffer_6386 (
        .din(new_Jinkela_wire_8073),
        .dout(new_Jinkela_wire_8074)
    );

    bfr new_Jinkela_buffer_3090 (
        .din(new_Jinkela_wire_4179),
        .dout(new_Jinkela_wire_4180)
    );

    bfr new_Jinkela_buffer_9898 (
        .din(new_Jinkela_wire_12017),
        .dout(new_Jinkela_wire_12018)
    );

    bfr new_Jinkela_buffer_6429 (
        .din(new_Jinkela_wire_8120),
        .dout(new_Jinkela_wire_8121)
    );

    bfr new_Jinkela_buffer_2969 (
        .din(new_Jinkela_wire_4040),
        .dout(new_Jinkela_wire_4041)
    );

    bfr new_Jinkela_buffer_9949 (
        .din(new_Jinkela_wire_12088),
        .dout(new_Jinkela_wire_12089)
    );

    bfr new_Jinkela_buffer_6387 (
        .din(new_Jinkela_wire_8074),
        .dout(new_Jinkela_wire_8075)
    );

    bfr new_Jinkela_buffer_3036 (
        .din(new_Jinkela_wire_4117),
        .dout(new_Jinkela_wire_4118)
    );

    bfr new_Jinkela_buffer_9899 (
        .din(new_Jinkela_wire_12018),
        .dout(new_Jinkela_wire_12019)
    );

    bfr new_Jinkela_buffer_6511 (
        .din(new_Jinkela_wire_8210),
        .dout(new_Jinkela_wire_8211)
    );

    bfr new_Jinkela_buffer_2970 (
        .din(new_Jinkela_wire_4041),
        .dout(new_Jinkela_wire_4042)
    );

    bfr new_Jinkela_buffer_6494 (
        .din(new_Jinkela_wire_8193),
        .dout(new_Jinkela_wire_8194)
    );

    bfr new_Jinkela_buffer_6388 (
        .din(new_Jinkela_wire_8075),
        .dout(new_Jinkela_wire_8076)
    );

    bfr new_Jinkela_buffer_3162 (
        .din(new_Jinkela_wire_4265),
        .dout(new_Jinkela_wire_4266)
    );

    bfr new_Jinkela_buffer_9900 (
        .din(new_Jinkela_wire_12019),
        .dout(new_Jinkela_wire_12020)
    );

    bfr new_Jinkela_buffer_3152 (
        .din(new_Jinkela_wire_4255),
        .dout(new_Jinkela_wire_4256)
    );

    bfr new_Jinkela_buffer_6430 (
        .din(new_Jinkela_wire_8121),
        .dout(new_Jinkela_wire_8122)
    );

    bfr new_Jinkela_buffer_2971 (
        .din(new_Jinkela_wire_4042),
        .dout(new_Jinkela_wire_4043)
    );

    bfr new_Jinkela_buffer_9950 (
        .din(new_Jinkela_wire_12089),
        .dout(new_Jinkela_wire_12090)
    );

    bfr new_Jinkela_buffer_6389 (
        .din(new_Jinkela_wire_8076),
        .dout(new_Jinkela_wire_8077)
    );

    bfr new_Jinkela_buffer_3037 (
        .din(new_Jinkela_wire_4118),
        .dout(new_Jinkela_wire_4119)
    );

    bfr new_Jinkela_buffer_9901 (
        .din(new_Jinkela_wire_12020),
        .dout(new_Jinkela_wire_12021)
    );

    bfr new_Jinkela_buffer_10074 (
        .din(new_Jinkela_wire_12223),
        .dout(new_Jinkela_wire_12224)
    );

    bfr new_Jinkela_buffer_2972 (
        .din(new_Jinkela_wire_4043),
        .dout(new_Jinkela_wire_4044)
    );

    bfr new_Jinkela_buffer_9973 (
        .din(new_Jinkela_wire_12118),
        .dout(new_Jinkela_wire_12119)
    );

    bfr new_Jinkela_buffer_6390 (
        .din(new_Jinkela_wire_8077),
        .dout(new_Jinkela_wire_8078)
    );

    bfr new_Jinkela_buffer_3091 (
        .din(new_Jinkela_wire_4180),
        .dout(new_Jinkela_wire_4181)
    );

    bfr new_Jinkela_buffer_9902 (
        .din(new_Jinkela_wire_12021),
        .dout(new_Jinkela_wire_12022)
    );

    bfr new_Jinkela_buffer_6431 (
        .din(new_Jinkela_wire_8122),
        .dout(new_Jinkela_wire_8123)
    );

    bfr new_Jinkela_buffer_2973 (
        .din(new_Jinkela_wire_4044),
        .dout(new_Jinkela_wire_4045)
    );

    bfr new_Jinkela_buffer_9951 (
        .din(new_Jinkela_wire_12090),
        .dout(new_Jinkela_wire_12091)
    );

    bfr new_Jinkela_buffer_6391 (
        .din(new_Jinkela_wire_8078),
        .dout(new_Jinkela_wire_8079)
    );

    bfr new_Jinkela_buffer_3038 (
        .din(new_Jinkela_wire_4119),
        .dout(new_Jinkela_wire_4120)
    );

    bfr new_Jinkela_buffer_9903 (
        .din(new_Jinkela_wire_12022),
        .dout(new_Jinkela_wire_12023)
    );

    spl2 new_Jinkela_splitter_703 (
        .a(_1088_),
        .b(new_Jinkela_wire_8282),
        .c(new_Jinkela_wire_8283)
    );

    bfr new_Jinkela_buffer_2974 (
        .din(new_Jinkela_wire_4045),
        .dout(new_Jinkela_wire_4046)
    );

    bfr new_Jinkela_buffer_6495 (
        .din(new_Jinkela_wire_8194),
        .dout(new_Jinkela_wire_8195)
    );

    bfr new_Jinkela_buffer_9904 (
        .din(new_Jinkela_wire_12023),
        .dout(new_Jinkela_wire_12024)
    );

    bfr new_Jinkela_buffer_6392 (
        .din(new_Jinkela_wire_8079),
        .dout(new_Jinkela_wire_8080)
    );

    bfr new_Jinkela_buffer_6432 (
        .din(new_Jinkela_wire_8123),
        .dout(new_Jinkela_wire_8124)
    );

    bfr new_Jinkela_buffer_2975 (
        .din(new_Jinkela_wire_4046),
        .dout(new_Jinkela_wire_4047)
    );

    bfr new_Jinkela_buffer_9952 (
        .din(new_Jinkela_wire_12091),
        .dout(new_Jinkela_wire_12092)
    );

    bfr new_Jinkela_buffer_6393 (
        .din(new_Jinkela_wire_8080),
        .dout(new_Jinkela_wire_8081)
    );

    bfr new_Jinkela_buffer_3039 (
        .din(new_Jinkela_wire_4120),
        .dout(new_Jinkela_wire_4121)
    );

    bfr new_Jinkela_buffer_9905 (
        .din(new_Jinkela_wire_12024),
        .dout(new_Jinkela_wire_12025)
    );

    bfr new_Jinkela_buffer_10029 (
        .din(new_Jinkela_wire_12174),
        .dout(new_Jinkela_wire_12175)
    );

    bfr new_Jinkela_buffer_2976 (
        .din(new_Jinkela_wire_4047),
        .dout(new_Jinkela_wire_4048)
    );

    spl2 new_Jinkela_splitter_702 (
        .a(_0050_),
        .b(new_Jinkela_wire_8280),
        .c(new_Jinkela_wire_8281)
    );

    bfr new_Jinkela_buffer_9974 (
        .din(new_Jinkela_wire_12119),
        .dout(new_Jinkela_wire_12120)
    );

    bfr new_Jinkela_buffer_6394 (
        .din(new_Jinkela_wire_8081),
        .dout(new_Jinkela_wire_8082)
    );

    bfr new_Jinkela_buffer_3092 (
        .din(new_Jinkela_wire_4181),
        .dout(new_Jinkela_wire_4182)
    );

    bfr new_Jinkela_buffer_9906 (
        .din(new_Jinkela_wire_12025),
        .dout(new_Jinkela_wire_12026)
    );

    bfr new_Jinkela_buffer_6433 (
        .din(new_Jinkela_wire_8124),
        .dout(new_Jinkela_wire_8125)
    );

    bfr new_Jinkela_buffer_2977 (
        .din(new_Jinkela_wire_4048),
        .dout(new_Jinkela_wire_4049)
    );

    bfr new_Jinkela_buffer_9953 (
        .din(new_Jinkela_wire_12092),
        .dout(new_Jinkela_wire_12093)
    );

    bfr new_Jinkela_buffer_6395 (
        .din(new_Jinkela_wire_8082),
        .dout(new_Jinkela_wire_8083)
    );

    bfr new_Jinkela_buffer_3040 (
        .din(new_Jinkela_wire_4121),
        .dout(new_Jinkela_wire_4122)
    );

    bfr new_Jinkela_buffer_9907 (
        .din(new_Jinkela_wire_12026),
        .dout(new_Jinkela_wire_12027)
    );

    bfr new_Jinkela_buffer_6512 (
        .din(new_Jinkela_wire_8211),
        .dout(new_Jinkela_wire_8212)
    );

    bfr new_Jinkela_buffer_2978 (
        .din(new_Jinkela_wire_4049),
        .dout(new_Jinkela_wire_4050)
    );

    bfr new_Jinkela_buffer_6496 (
        .din(new_Jinkela_wire_8195),
        .dout(new_Jinkela_wire_8196)
    );

    bfr new_Jinkela_buffer_13348 (
        .din(new_Jinkela_wire_15949),
        .dout(new_Jinkela_wire_15950)
    );

    spl2 new_Jinkela_splitter_1166 (
        .a(_0720_),
        .b(new_Jinkela_wire_16123),
        .c(new_Jinkela_wire_16124)
    );

    bfr new_Jinkela_buffer_13349 (
        .din(new_Jinkela_wire_15950),
        .dout(new_Jinkela_wire_15951)
    );

    bfr new_Jinkela_buffer_13409 (
        .din(new_Jinkela_wire_16022),
        .dout(new_Jinkela_wire_16023)
    );

    bfr new_Jinkela_buffer_13350 (
        .din(new_Jinkela_wire_15951),
        .dout(new_Jinkela_wire_15952)
    );

    spl2 new_Jinkela_splitter_1165 (
        .a(_0207_),
        .b(new_Jinkela_wire_16121),
        .c(new_Jinkela_wire_16122)
    );

    bfr new_Jinkela_buffer_13351 (
        .din(new_Jinkela_wire_15952),
        .dout(new_Jinkela_wire_15953)
    );

    bfr new_Jinkela_buffer_13410 (
        .din(new_Jinkela_wire_16023),
        .dout(new_Jinkela_wire_16024)
    );

    bfr new_Jinkela_buffer_13352 (
        .din(new_Jinkela_wire_15953),
        .dout(new_Jinkela_wire_15954)
    );

    bfr new_Jinkela_buffer_13353 (
        .din(new_Jinkela_wire_15954),
        .dout(new_Jinkela_wire_15955)
    );

    bfr new_Jinkela_buffer_13411 (
        .din(new_Jinkela_wire_16024),
        .dout(new_Jinkela_wire_16025)
    );

    bfr new_Jinkela_buffer_13354 (
        .din(new_Jinkela_wire_15955),
        .dout(new_Jinkela_wire_15956)
    );

    spl2 new_Jinkela_splitter_1167 (
        .a(_1600_),
        .b(new_Jinkela_wire_16125),
        .c(new_Jinkela_wire_16126)
    );

    bfr new_Jinkela_buffer_13355 (
        .din(new_Jinkela_wire_15956),
        .dout(new_Jinkela_wire_15957)
    );

    bfr new_Jinkela_buffer_13412 (
        .din(new_Jinkela_wire_16025),
        .dout(new_Jinkela_wire_16026)
    );

    bfr new_Jinkela_buffer_13356 (
        .din(new_Jinkela_wire_15957),
        .dout(new_Jinkela_wire_15958)
    );

    bfr new_Jinkela_buffer_13493 (
        .din(_1369_),
        .dout(new_Jinkela_wire_16131)
    );

    bfr new_Jinkela_buffer_13357 (
        .din(new_Jinkela_wire_15958),
        .dout(new_Jinkela_wire_15959)
    );

    bfr new_Jinkela_buffer_13413 (
        .din(new_Jinkela_wire_16026),
        .dout(new_Jinkela_wire_16027)
    );

    bfr new_Jinkela_buffer_13358 (
        .din(new_Jinkela_wire_15959),
        .dout(new_Jinkela_wire_15960)
    );

    bfr new_Jinkela_buffer_13489 (
        .din(new_Jinkela_wire_16126),
        .dout(new_Jinkela_wire_16127)
    );

    spl2 new_Jinkela_splitter_1169 (
        .a(_0818_),
        .b(new_Jinkela_wire_16190),
        .c(new_Jinkela_wire_16191)
    );

    bfr new_Jinkela_buffer_13359 (
        .din(new_Jinkela_wire_15960),
        .dout(new_Jinkela_wire_15961)
    );

    bfr new_Jinkela_buffer_13414 (
        .din(new_Jinkela_wire_16027),
        .dout(new_Jinkela_wire_16028)
    );

    bfr new_Jinkela_buffer_13360 (
        .din(new_Jinkela_wire_15961),
        .dout(new_Jinkela_wire_15962)
    );

    bfr new_Jinkela_buffer_13361 (
        .din(new_Jinkela_wire_15962),
        .dout(new_Jinkela_wire_15963)
    );

    bfr new_Jinkela_buffer_13415 (
        .din(new_Jinkela_wire_16028),
        .dout(new_Jinkela_wire_16029)
    );

    bfr new_Jinkela_buffer_13362 (
        .din(new_Jinkela_wire_15963),
        .dout(new_Jinkela_wire_15964)
    );

    bfr new_Jinkela_buffer_13490 (
        .din(new_Jinkela_wire_16127),
        .dout(new_Jinkela_wire_16128)
    );

    bfr new_Jinkela_buffer_13363 (
        .din(new_Jinkela_wire_15964),
        .dout(new_Jinkela_wire_15965)
    );

    bfr new_Jinkela_buffer_13416 (
        .din(new_Jinkela_wire_16029),
        .dout(new_Jinkela_wire_16030)
    );

    bfr new_Jinkela_buffer_13364 (
        .din(new_Jinkela_wire_15965),
        .dout(new_Jinkela_wire_15966)
    );

    bfr new_Jinkela_buffer_13494 (
        .din(new_Jinkela_wire_16131),
        .dout(new_Jinkela_wire_16132)
    );

    bfr new_Jinkela_buffer_13365 (
        .din(new_Jinkela_wire_15966),
        .dout(new_Jinkela_wire_15967)
    );

    bfr new_Jinkela_buffer_13417 (
        .din(new_Jinkela_wire_16030),
        .dout(new_Jinkela_wire_16031)
    );

    bfr new_Jinkela_buffer_13366 (
        .din(new_Jinkela_wire_15967),
        .dout(new_Jinkela_wire_15968)
    );

    bfr new_Jinkela_buffer_13491 (
        .din(new_Jinkela_wire_16128),
        .dout(new_Jinkela_wire_16129)
    );

    bfr new_Jinkela_buffer_13367 (
        .din(new_Jinkela_wire_15968),
        .dout(new_Jinkela_wire_15969)
    );

    bfr new_Jinkela_buffer_13418 (
        .din(new_Jinkela_wire_16031),
        .dout(new_Jinkela_wire_16032)
    );

    bfr new_Jinkela_buffer_13368 (
        .din(new_Jinkela_wire_15969),
        .dout(new_Jinkela_wire_15970)
    );

    spl2 new_Jinkela_splitter_1171 (
        .a(_0860_),
        .b(new_Jinkela_wire_16194),
        .c(new_Jinkela_wire_16195)
    );

    bfr new_Jinkela_buffer_6396 (
        .din(new_Jinkela_wire_8083),
        .dout(new_Jinkela_wire_8084)
    );

    bfr new_Jinkela_buffer_6434 (
        .din(new_Jinkela_wire_8125),
        .dout(new_Jinkela_wire_8126)
    );

    bfr new_Jinkela_buffer_6397 (
        .din(new_Jinkela_wire_8084),
        .dout(new_Jinkela_wire_8085)
    );

    bfr new_Jinkela_buffer_6398 (
        .din(new_Jinkela_wire_8085),
        .dout(new_Jinkela_wire_8086)
    );

    bfr new_Jinkela_buffer_6435 (
        .din(new_Jinkela_wire_8126),
        .dout(new_Jinkela_wire_8127)
    );

    bfr new_Jinkela_buffer_6399 (
        .din(new_Jinkela_wire_8086),
        .dout(new_Jinkela_wire_8087)
    );

    bfr new_Jinkela_buffer_6497 (
        .din(new_Jinkela_wire_8196),
        .dout(new_Jinkela_wire_8197)
    );

    bfr new_Jinkela_buffer_6400 (
        .din(new_Jinkela_wire_8087),
        .dout(new_Jinkela_wire_8088)
    );

    bfr new_Jinkela_buffer_6436 (
        .din(new_Jinkela_wire_8127),
        .dout(new_Jinkela_wire_8128)
    );

    bfr new_Jinkela_buffer_6401 (
        .din(new_Jinkela_wire_8088),
        .dout(new_Jinkela_wire_8089)
    );

    bfr new_Jinkela_buffer_6402 (
        .din(new_Jinkela_wire_8089),
        .dout(new_Jinkela_wire_8090)
    );

    bfr new_Jinkela_buffer_6437 (
        .din(new_Jinkela_wire_8128),
        .dout(new_Jinkela_wire_8129)
    );

    bfr new_Jinkela_buffer_6403 (
        .din(new_Jinkela_wire_8090),
        .dout(new_Jinkela_wire_8091)
    );

    bfr new_Jinkela_buffer_6513 (
        .din(new_Jinkela_wire_8212),
        .dout(new_Jinkela_wire_8213)
    );

    bfr new_Jinkela_buffer_6498 (
        .din(new_Jinkela_wire_8197),
        .dout(new_Jinkela_wire_8198)
    );

    bfr new_Jinkela_buffer_6404 (
        .din(new_Jinkela_wire_8091),
        .dout(new_Jinkela_wire_8092)
    );

    bfr new_Jinkela_buffer_6438 (
        .din(new_Jinkela_wire_8129),
        .dout(new_Jinkela_wire_8130)
    );

    spl2 new_Jinkela_splitter_693 (
        .a(new_Jinkela_wire_8092),
        .b(new_Jinkela_wire_8093),
        .c(new_Jinkela_wire_8094)
    );

    bfr new_Jinkela_buffer_6439 (
        .din(new_Jinkela_wire_8130),
        .dout(new_Jinkela_wire_8131)
    );

    bfr new_Jinkela_buffer_6499 (
        .din(new_Jinkela_wire_8198),
        .dout(new_Jinkela_wire_8199)
    );

    bfr new_Jinkela_buffer_6440 (
        .din(new_Jinkela_wire_8131),
        .dout(new_Jinkela_wire_8132)
    );

    spl2 new_Jinkela_splitter_704 (
        .a(_0242_),
        .b(new_Jinkela_wire_8288),
        .c(new_Jinkela_wire_8289)
    );

    bfr new_Jinkela_buffer_6441 (
        .din(new_Jinkela_wire_8132),
        .dout(new_Jinkela_wire_8133)
    );

    bfr new_Jinkela_buffer_6514 (
        .din(new_Jinkela_wire_8213),
        .dout(new_Jinkela_wire_8214)
    );

    bfr new_Jinkela_buffer_6500 (
        .din(new_Jinkela_wire_8199),
        .dout(new_Jinkela_wire_8200)
    );

    bfr new_Jinkela_buffer_6442 (
        .din(new_Jinkela_wire_8133),
        .dout(new_Jinkela_wire_8134)
    );

    bfr new_Jinkela_buffer_6443 (
        .din(new_Jinkela_wire_8134),
        .dout(new_Jinkela_wire_8135)
    );

    bfr new_Jinkela_buffer_6574 (
        .din(new_Jinkela_wire_8283),
        .dout(new_Jinkela_wire_8284)
    );

    bfr new_Jinkela_buffer_6501 (
        .din(new_Jinkela_wire_8200),
        .dout(new_Jinkela_wire_8201)
    );

    bfr new_Jinkela_buffer_6444 (
        .din(new_Jinkela_wire_8135),
        .dout(new_Jinkela_wire_8136)
    );

    spl2 new_Jinkela_splitter_705 (
        .a(_1010_),
        .b(new_Jinkela_wire_8290),
        .c(new_Jinkela_wire_8291)
    );

    bfr new_Jinkela_buffer_6445 (
        .din(new_Jinkela_wire_8136),
        .dout(new_Jinkela_wire_8137)
    );

    bfr new_Jinkela_buffer_6515 (
        .din(new_Jinkela_wire_8214),
        .dout(new_Jinkela_wire_8215)
    );

    bfr new_Jinkela_buffer_6502 (
        .din(new_Jinkela_wire_8201),
        .dout(new_Jinkela_wire_8202)
    );

    bfr new_Jinkela_buffer_6446 (
        .din(new_Jinkela_wire_8137),
        .dout(new_Jinkela_wire_8138)
    );

    bfr new_Jinkela_buffer_6447 (
        .din(new_Jinkela_wire_8138),
        .dout(new_Jinkela_wire_8139)
    );

    spl2 new_Jinkela_splitter_706 (
        .a(_1541_),
        .b(new_Jinkela_wire_8292),
        .c(new_Jinkela_wire_8293)
    );

    bfr new_Jinkela_buffer_6503 (
        .din(new_Jinkela_wire_8202),
        .dout(new_Jinkela_wire_8203)
    );

    bfr new_Jinkela_buffer_6448 (
        .din(new_Jinkela_wire_8139),
        .dout(new_Jinkela_wire_8140)
    );

    bfr new_Jinkela_buffer_6449 (
        .din(new_Jinkela_wire_8140),
        .dout(new_Jinkela_wire_8141)
    );

    bfr new_Jinkela_buffer_6516 (
        .din(new_Jinkela_wire_8215),
        .dout(new_Jinkela_wire_8216)
    );

    bfr new_Jinkela_buffer_6504 (
        .din(new_Jinkela_wire_8203),
        .dout(new_Jinkela_wire_8204)
    );

    bfr new_Jinkela_buffer_13369 (
        .din(new_Jinkela_wire_15970),
        .dout(new_Jinkela_wire_15971)
    );

    bfr new_Jinkela_buffer_3153 (
        .din(new_Jinkela_wire_4256),
        .dout(new_Jinkela_wire_4257)
    );

    bfr new_Jinkela_buffer_13421 (
        .din(new_Jinkela_wire_16034),
        .dout(new_Jinkela_wire_16035)
    );

    bfr new_Jinkela_buffer_2979 (
        .din(new_Jinkela_wire_4050),
        .dout(new_Jinkela_wire_4051)
    );

    bfr new_Jinkela_buffer_13370 (
        .din(new_Jinkela_wire_15971),
        .dout(new_Jinkela_wire_15972)
    );

    bfr new_Jinkela_buffer_3041 (
        .din(new_Jinkela_wire_4122),
        .dout(new_Jinkela_wire_4123)
    );

    bfr new_Jinkela_buffer_2980 (
        .din(new_Jinkela_wire_4051),
        .dout(new_Jinkela_wire_4052)
    );

    bfr new_Jinkela_buffer_13371 (
        .din(new_Jinkela_wire_15972),
        .dout(new_Jinkela_wire_15973)
    );

    bfr new_Jinkela_buffer_3093 (
        .din(new_Jinkela_wire_4182),
        .dout(new_Jinkela_wire_4183)
    );

    bfr new_Jinkela_buffer_13422 (
        .din(new_Jinkela_wire_16035),
        .dout(new_Jinkela_wire_16036)
    );

    bfr new_Jinkela_buffer_2981 (
        .din(new_Jinkela_wire_4052),
        .dout(new_Jinkela_wire_4053)
    );

    bfr new_Jinkela_buffer_13372 (
        .din(new_Jinkela_wire_15973),
        .dout(new_Jinkela_wire_15974)
    );

    bfr new_Jinkela_buffer_3042 (
        .din(new_Jinkela_wire_4123),
        .dout(new_Jinkela_wire_4124)
    );

    bfr new_Jinkela_buffer_13496 (
        .din(new_Jinkela_wire_16133),
        .dout(new_Jinkela_wire_16134)
    );

    bfr new_Jinkela_buffer_2982 (
        .din(new_Jinkela_wire_4053),
        .dout(new_Jinkela_wire_4054)
    );

    bfr new_Jinkela_buffer_13373 (
        .din(new_Jinkela_wire_15974),
        .dout(new_Jinkela_wire_15975)
    );

    bfr new_Jinkela_buffer_3177 (
        .din(new_Jinkela_wire_4286),
        .dout(new_Jinkela_wire_4287)
    );

    bfr new_Jinkela_buffer_13423 (
        .din(new_Jinkela_wire_16036),
        .dout(new_Jinkela_wire_16037)
    );

    bfr new_Jinkela_buffer_2983 (
        .din(new_Jinkela_wire_4054),
        .dout(new_Jinkela_wire_4055)
    );

    bfr new_Jinkela_buffer_13374 (
        .din(new_Jinkela_wire_15975),
        .dout(new_Jinkela_wire_15976)
    );

    bfr new_Jinkela_buffer_3043 (
        .din(new_Jinkela_wire_4124),
        .dout(new_Jinkela_wire_4125)
    );

    bfr new_Jinkela_buffer_2984 (
        .din(new_Jinkela_wire_4055),
        .dout(new_Jinkela_wire_4056)
    );

    bfr new_Jinkela_buffer_13554 (
        .din(_1232_),
        .dout(new_Jinkela_wire_16200)
    );

    bfr new_Jinkela_buffer_13375 (
        .din(new_Jinkela_wire_15976),
        .dout(new_Jinkela_wire_15977)
    );

    bfr new_Jinkela_buffer_3094 (
        .din(new_Jinkela_wire_4183),
        .dout(new_Jinkela_wire_4184)
    );

    bfr new_Jinkela_buffer_13424 (
        .din(new_Jinkela_wire_16037),
        .dout(new_Jinkela_wire_16038)
    );

    bfr new_Jinkela_buffer_2985 (
        .din(new_Jinkela_wire_4056),
        .dout(new_Jinkela_wire_4057)
    );

    bfr new_Jinkela_buffer_13376 (
        .din(new_Jinkela_wire_15977),
        .dout(new_Jinkela_wire_15978)
    );

    bfr new_Jinkela_buffer_3044 (
        .din(new_Jinkela_wire_4125),
        .dout(new_Jinkela_wire_4126)
    );

    bfr new_Jinkela_buffer_13497 (
        .din(new_Jinkela_wire_16134),
        .dout(new_Jinkela_wire_16135)
    );

    bfr new_Jinkela_buffer_2986 (
        .din(new_Jinkela_wire_4057),
        .dout(new_Jinkela_wire_4058)
    );

    bfr new_Jinkela_buffer_13377 (
        .din(new_Jinkela_wire_15978),
        .dout(new_Jinkela_wire_15979)
    );

    bfr new_Jinkela_buffer_3163 (
        .din(new_Jinkela_wire_4266),
        .dout(new_Jinkela_wire_4267)
    );

    bfr new_Jinkela_buffer_3154 (
        .din(new_Jinkela_wire_4257),
        .dout(new_Jinkela_wire_4258)
    );

    bfr new_Jinkela_buffer_13425 (
        .din(new_Jinkela_wire_16038),
        .dout(new_Jinkela_wire_16039)
    );

    bfr new_Jinkela_buffer_2987 (
        .din(new_Jinkela_wire_4058),
        .dout(new_Jinkela_wire_4059)
    );

    bfr new_Jinkela_buffer_13378 (
        .din(new_Jinkela_wire_15979),
        .dout(new_Jinkela_wire_15980)
    );

    bfr new_Jinkela_buffer_3045 (
        .din(new_Jinkela_wire_4126),
        .dout(new_Jinkela_wire_4127)
    );

    bfr new_Jinkela_buffer_13550 (
        .din(new_Jinkela_wire_16195),
        .dout(new_Jinkela_wire_16196)
    );

    bfr new_Jinkela_buffer_2988 (
        .din(new_Jinkela_wire_4059),
        .dout(new_Jinkela_wire_4060)
    );

    spl2 new_Jinkela_splitter_1172 (
        .a(_0817_),
        .b(new_Jinkela_wire_16201),
        .c(new_Jinkela_wire_16202)
    );

    bfr new_Jinkela_buffer_13379 (
        .din(new_Jinkela_wire_15980),
        .dout(new_Jinkela_wire_15981)
    );

    bfr new_Jinkela_buffer_3095 (
        .din(new_Jinkela_wire_4184),
        .dout(new_Jinkela_wire_4185)
    );

    bfr new_Jinkela_buffer_13426 (
        .din(new_Jinkela_wire_16039),
        .dout(new_Jinkela_wire_16040)
    );

    bfr new_Jinkela_buffer_2989 (
        .din(new_Jinkela_wire_4060),
        .dout(new_Jinkela_wire_4061)
    );

    bfr new_Jinkela_buffer_13380 (
        .din(new_Jinkela_wire_15981),
        .dout(new_Jinkela_wire_15982)
    );

    bfr new_Jinkela_buffer_3046 (
        .din(new_Jinkela_wire_4127),
        .dout(new_Jinkela_wire_4128)
    );

    bfr new_Jinkela_buffer_13498 (
        .din(new_Jinkela_wire_16135),
        .dout(new_Jinkela_wire_16136)
    );

    bfr new_Jinkela_buffer_2990 (
        .din(new_Jinkela_wire_4061),
        .dout(new_Jinkela_wire_4062)
    );

    bfr new_Jinkela_buffer_13381 (
        .din(new_Jinkela_wire_15982),
        .dout(new_Jinkela_wire_15983)
    );

    bfr new_Jinkela_buffer_13427 (
        .din(new_Jinkela_wire_16040),
        .dout(new_Jinkela_wire_16041)
    );

    bfr new_Jinkela_buffer_2991 (
        .din(new_Jinkela_wire_4062),
        .dout(new_Jinkela_wire_4063)
    );

    bfr new_Jinkela_buffer_13382 (
        .din(new_Jinkela_wire_15983),
        .dout(new_Jinkela_wire_15984)
    );

    bfr new_Jinkela_buffer_3047 (
        .din(new_Jinkela_wire_4128),
        .dout(new_Jinkela_wire_4129)
    );

    spl2 new_Jinkela_splitter_1173 (
        .a(_0149_),
        .b(new_Jinkela_wire_16203),
        .c(new_Jinkela_wire_16204)
    );

    bfr new_Jinkela_buffer_2992 (
        .din(new_Jinkela_wire_4063),
        .dout(new_Jinkela_wire_4064)
    );

    bfr new_Jinkela_buffer_13383 (
        .din(new_Jinkela_wire_15984),
        .dout(new_Jinkela_wire_15985)
    );

    bfr new_Jinkela_buffer_3096 (
        .din(new_Jinkela_wire_4185),
        .dout(new_Jinkela_wire_4186)
    );

    bfr new_Jinkela_buffer_13428 (
        .din(new_Jinkela_wire_16041),
        .dout(new_Jinkela_wire_16042)
    );

    bfr new_Jinkela_buffer_2993 (
        .din(new_Jinkela_wire_4064),
        .dout(new_Jinkela_wire_4065)
    );

    bfr new_Jinkela_buffer_13384 (
        .din(new_Jinkela_wire_15985),
        .dout(new_Jinkela_wire_15986)
    );

    bfr new_Jinkela_buffer_3048 (
        .din(new_Jinkela_wire_4129),
        .dout(new_Jinkela_wire_4130)
    );

    bfr new_Jinkela_buffer_13499 (
        .din(new_Jinkela_wire_16136),
        .dout(new_Jinkela_wire_16137)
    );

    bfr new_Jinkela_buffer_2994 (
        .din(new_Jinkela_wire_4065),
        .dout(new_Jinkela_wire_4066)
    );

    bfr new_Jinkela_buffer_13385 (
        .din(new_Jinkela_wire_15986),
        .dout(new_Jinkela_wire_15987)
    );

    bfr new_Jinkela_buffer_3155 (
        .din(new_Jinkela_wire_4258),
        .dout(new_Jinkela_wire_4259)
    );

    bfr new_Jinkela_buffer_13429 (
        .din(new_Jinkela_wire_16042),
        .dout(new_Jinkela_wire_16043)
    );

    bfr new_Jinkela_buffer_2995 (
        .din(new_Jinkela_wire_4066),
        .dout(new_Jinkela_wire_4067)
    );

    bfr new_Jinkela_buffer_13386 (
        .din(new_Jinkela_wire_15987),
        .dout(new_Jinkela_wire_15988)
    );

    bfr new_Jinkela_buffer_3049 (
        .din(new_Jinkela_wire_4130),
        .dout(new_Jinkela_wire_4131)
    );

    bfr new_Jinkela_buffer_13551 (
        .din(new_Jinkela_wire_16196),
        .dout(new_Jinkela_wire_16197)
    );

    bfr new_Jinkela_buffer_2996 (
        .din(new_Jinkela_wire_4067),
        .dout(new_Jinkela_wire_4068)
    );

    bfr new_Jinkela_buffer_13387 (
        .din(new_Jinkela_wire_15988),
        .dout(new_Jinkela_wire_15989)
    );

    bfr new_Jinkela_buffer_3097 (
        .din(new_Jinkela_wire_4186),
        .dout(new_Jinkela_wire_4187)
    );

    bfr new_Jinkela_buffer_13430 (
        .din(new_Jinkela_wire_16043),
        .dout(new_Jinkela_wire_16044)
    );

    bfr new_Jinkela_buffer_2997 (
        .din(new_Jinkela_wire_4068),
        .dout(new_Jinkela_wire_4069)
    );

    bfr new_Jinkela_buffer_13388 (
        .din(new_Jinkela_wire_15989),
        .dout(new_Jinkela_wire_15990)
    );

    bfr new_Jinkela_buffer_3050 (
        .din(new_Jinkela_wire_4131),
        .dout(new_Jinkela_wire_4132)
    );

    bfr new_Jinkela_buffer_13500 (
        .din(new_Jinkela_wire_16137),
        .dout(new_Jinkela_wire_16138)
    );

    spl2 new_Jinkela_splitter_385 (
        .a(new_Jinkela_wire_4069),
        .b(new_Jinkela_wire_4070),
        .c(new_Jinkela_wire_4071)
    );

    bfr new_Jinkela_buffer_13389 (
        .din(new_Jinkela_wire_15990),
        .dout(new_Jinkela_wire_15991)
    );

    bfr new_Jinkela_buffer_3051 (
        .din(new_Jinkela_wire_4132),
        .dout(new_Jinkela_wire_4133)
    );

    bfr new_Jinkela_buffer_13431 (
        .din(new_Jinkela_wire_16044),
        .dout(new_Jinkela_wire_16045)
    );

    bfr new_Jinkela_buffer_3181 (
        .din(_0714_),
        .dout(new_Jinkela_wire_4291)
    );

    bfr new_Jinkela_buffer_16817 (
        .din(new_Jinkela_wire_20063),
        .dout(new_Jinkela_wire_20064)
    );

    and_bb _2161_ (
        .a(new_Jinkela_wire_1774),
        .b(new_Jinkela_wire_6845),
        .c(_1201_)
    );

    bfr new_Jinkela_buffer_16773 (
        .din(new_Jinkela_wire_20009),
        .dout(new_Jinkela_wire_20010)
    );

    or_bb _2162_ (
        .a(new_Jinkela_wire_4662),
        .b(new_Jinkela_wire_19117),
        .c(new_net_3954)
    );

    bfr new_Jinkela_buffer_16893 (
        .din(new_Jinkela_wire_20145),
        .dout(new_Jinkela_wire_20146)
    );

    and_bb _2163_ (
        .a(new_Jinkela_wire_20325),
        .b(new_Jinkela_wire_19959),
        .c(_1202_)
    );

    bfr new_Jinkela_buffer_16774 (
        .din(new_Jinkela_wire_20010),
        .dout(new_Jinkela_wire_20011)
    );

    or_bb _2164_ (
        .a(new_Jinkela_wire_5967),
        .b(new_Jinkela_wire_4672),
        .c(new_net_3974)
    );

    bfr new_Jinkela_buffer_16818 (
        .din(new_Jinkela_wire_20064),
        .dout(new_Jinkela_wire_20065)
    );

    and_bb _2165_ (
        .a(new_Jinkela_wire_121),
        .b(new_Jinkela_wire_338),
        .c(_1203_)
    );

    bfr new_Jinkela_buffer_16775 (
        .din(new_Jinkela_wire_20011),
        .dout(new_Jinkela_wire_20012)
    );

    and_bi _2166_ (
        .a(new_Jinkela_wire_6247),
        .b(new_Jinkela_wire_19108),
        .c(_1204_)
    );

    and_bb _2167_ (
        .a(new_Jinkela_wire_88),
        .b(new_Jinkela_wire_13),
        .c(_1205_)
    );

    spl2 new_Jinkela_splitter_1477 (
        .a(_1053_),
        .b(new_Jinkela_wire_20217),
        .c(new_Jinkela_wire_20218)
    );

    bfr new_Jinkela_buffer_16776 (
        .din(new_Jinkela_wire_20012),
        .dout(new_Jinkela_wire_20013)
    );

    and_bi _2168_ (
        .a(new_Jinkela_wire_10956),
        .b(new_Jinkela_wire_7274),
        .c(_1206_)
    );

    bfr new_Jinkela_buffer_16819 (
        .din(new_Jinkela_wire_20065),
        .dout(new_Jinkela_wire_20066)
    );

    and_bb _2169_ (
        .a(new_Jinkela_wire_457),
        .b(new_Jinkela_wire_553),
        .c(_1207_)
    );

    bfr new_Jinkela_buffer_16777 (
        .din(new_Jinkela_wire_20013),
        .dout(new_Jinkela_wire_20014)
    );

    and_bi _2170_ (
        .a(new_Jinkela_wire_13579),
        .b(new_Jinkela_wire_11396),
        .c(_1208_)
    );

    bfr new_Jinkela_buffer_16894 (
        .din(new_Jinkela_wire_20146),
        .dout(new_Jinkela_wire_20147)
    );

    and_bb _2171_ (
        .a(new_Jinkela_wire_283),
        .b(new_Jinkela_wire_258),
        .c(_1209_)
    );

    bfr new_Jinkela_buffer_16778 (
        .din(new_Jinkela_wire_20014),
        .dout(new_Jinkela_wire_20015)
    );

    and_bi _2172_ (
        .a(new_Jinkela_wire_8848),
        .b(new_Jinkela_wire_2459),
        .c(_1210_)
    );

    bfr new_Jinkela_buffer_16820 (
        .din(new_Jinkela_wire_20066),
        .dout(new_Jinkela_wire_20067)
    );

    and_bb _2173_ (
        .a(new_Jinkela_wire_69),
        .b(new_Jinkela_wire_286),
        .c(_1211_)
    );

    bfr new_Jinkela_buffer_16779 (
        .din(new_Jinkela_wire_20015),
        .dout(new_Jinkela_wire_20016)
    );

    and_bi _2174_ (
        .a(new_Jinkela_wire_1008),
        .b(new_Jinkela_wire_10836),
        .c(_1212_)
    );

    bfr new_Jinkela_buffer_16960 (
        .din(_1007_),
        .dout(new_Jinkela_wire_20219)
    );

    and_bb _2175_ (
        .a(new_Jinkela_wire_473),
        .b(new_Jinkela_wire_57),
        .c(_1213_)
    );

    bfr new_Jinkela_buffer_16780 (
        .din(new_Jinkela_wire_20016),
        .dout(new_Jinkela_wire_20017)
    );

    and_bi _2176_ (
        .a(new_Jinkela_wire_17036),
        .b(new_Jinkela_wire_3181),
        .c(_1214_)
    );

    bfr new_Jinkela_buffer_16821 (
        .din(new_Jinkela_wire_20067),
        .dout(new_Jinkela_wire_20068)
    );

    and_bb _2177_ (
        .a(new_Jinkela_wire_370),
        .b(new_Jinkela_wire_651),
        .c(_1215_)
    );

    bfr new_Jinkela_buffer_16781 (
        .din(new_Jinkela_wire_20017),
        .dout(new_Jinkela_wire_20018)
    );

    and_bi _2178_ (
        .a(new_Jinkela_wire_12620),
        .b(new_Jinkela_wire_5996),
        .c(_1216_)
    );

    bfr new_Jinkela_buffer_16895 (
        .din(new_Jinkela_wire_20147),
        .dout(new_Jinkela_wire_20148)
    );

    and_bb _2179_ (
        .a(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_626),
        .c(_1217_)
    );

    bfr new_Jinkela_buffer_16782 (
        .din(new_Jinkela_wire_20018),
        .dout(new_Jinkela_wire_20019)
    );

    and_bi _2180_ (
        .a(new_Jinkela_wire_3708),
        .b(new_Jinkela_wire_18762),
        .c(_1218_)
    );

    bfr new_Jinkela_buffer_16822 (
        .din(new_Jinkela_wire_20068),
        .dout(new_Jinkela_wire_20069)
    );

    and_bb _2181_ (
        .a(new_Jinkela_wire_549),
        .b(new_Jinkela_wire_506),
        .c(_1219_)
    );

    bfr new_Jinkela_buffer_16783 (
        .din(new_Jinkela_wire_20019),
        .dout(new_Jinkela_wire_20020)
    );

    or_ii _2182_ (
        .a(new_Jinkela_wire_182),
        .b(new_Jinkela_wire_321),
        .c(_1220_)
    );

    bfr new_Jinkela_buffer_16956 (
        .din(new_Jinkela_wire_20212),
        .dout(new_Jinkela_wire_20213)
    );

    and_bi _2183_ (
        .a(new_Jinkela_wire_17050),
        .b(new_Jinkela_wire_6516),
        .c(_1221_)
    );

    bfr new_Jinkela_buffer_16784 (
        .din(new_Jinkela_wire_20020),
        .dout(new_Jinkela_wire_20021)
    );

    and_bb _2184_ (
        .a(new_Jinkela_wire_191),
        .b(new_Jinkela_wire_236),
        .c(_1222_)
    );

    bfr new_Jinkela_buffer_16823 (
        .din(new_Jinkela_wire_20069),
        .dout(new_Jinkela_wire_20070)
    );

    and_bi _2185_ (
        .a(new_Jinkela_wire_1569),
        .b(new_Jinkela_wire_1803),
        .c(_1223_)
    );

    bfr new_Jinkela_buffer_16785 (
        .din(new_Jinkela_wire_20021),
        .dout(new_Jinkela_wire_20022)
    );

    and_ii _2186_ (
        .a(new_Jinkela_wire_7714),
        .b(new_Jinkela_wire_15747),
        .c(_1224_)
    );

    bfr new_Jinkela_buffer_16896 (
        .din(new_Jinkela_wire_20148),
        .dout(new_Jinkela_wire_20149)
    );

    or_bb _2187_ (
        .a(new_Jinkela_wire_9740),
        .b(new_Jinkela_wire_3961),
        .c(_1225_)
    );

    bfr new_Jinkela_buffer_16786 (
        .din(new_Jinkela_wire_20022),
        .dout(new_Jinkela_wire_20023)
    );

    or_ii _2188_ (
        .a(new_Jinkela_wire_9741),
        .b(new_Jinkela_wire_3962),
        .c(_1226_)
    );

    bfr new_Jinkela_buffer_16824 (
        .din(new_Jinkela_wire_20070),
        .dout(new_Jinkela_wire_20071)
    );

    or_ii _2189_ (
        .a(new_Jinkela_wire_10061),
        .b(new_Jinkela_wire_6411),
        .c(_1227_)
    );

    bfr new_Jinkela_buffer_16787 (
        .din(new_Jinkela_wire_20023),
        .dout(new_Jinkela_wire_20024)
    );

    and_ii _2190_ (
        .a(new_Jinkela_wire_6010),
        .b(new_Jinkela_wire_19075),
        .c(_1228_)
    );

    bfr new_Jinkela_buffer_16961 (
        .din(_0548_),
        .dout(new_Jinkela_wire_20220)
    );

    and_bb _2191_ (
        .a(new_Jinkela_wire_6011),
        .b(new_Jinkela_wire_19076),
        .c(_1229_)
    );

    bfr new_Jinkela_buffer_16788 (
        .din(new_Jinkela_wire_20024),
        .dout(new_Jinkela_wire_20025)
    );

    or_bb _2192_ (
        .a(new_Jinkela_wire_16532),
        .b(new_Jinkela_wire_3361),
        .c(_1230_)
    );

    bfr new_Jinkela_buffer_16825 (
        .din(new_Jinkela_wire_20071),
        .dout(new_Jinkela_wire_20072)
    );

    or_bb _2193_ (
        .a(new_Jinkela_wire_18526),
        .b(new_Jinkela_wire_17981),
        .c(_1231_)
    );

    bfr new_Jinkela_buffer_16789 (
        .din(new_Jinkela_wire_20025),
        .dout(new_Jinkela_wire_20026)
    );

    or_ii _2194_ (
        .a(new_Jinkela_wire_18527),
        .b(new_Jinkela_wire_17982),
        .c(_1232_)
    );

    bfr new_Jinkela_buffer_16897 (
        .din(new_Jinkela_wire_20149),
        .dout(new_Jinkela_wire_20150)
    );

    or_ii _2195_ (
        .a(new_Jinkela_wire_16200),
        .b(new_Jinkela_wire_4285),
        .c(_1233_)
    );

    bfr new_Jinkela_buffer_16790 (
        .din(new_Jinkela_wire_20026),
        .dout(new_Jinkela_wire_20027)
    );

    and_ii _2196_ (
        .a(new_Jinkela_wire_20576),
        .b(new_Jinkela_wire_14681),
        .c(_1234_)
    );

    bfr new_Jinkela_buffer_16826 (
        .din(new_Jinkela_wire_20072),
        .dout(new_Jinkela_wire_20073)
    );

    and_bb _2197_ (
        .a(new_Jinkela_wire_20577),
        .b(new_Jinkela_wire_14682),
        .c(_1235_)
    );

    bfr new_Jinkela_buffer_16791 (
        .din(new_Jinkela_wire_20027),
        .dout(new_Jinkela_wire_20028)
    );

    or_bb _2198_ (
        .a(new_Jinkela_wire_5447),
        .b(new_Jinkela_wire_7292),
        .c(_1236_)
    );

    bfr new_Jinkela_buffer_16957 (
        .din(new_Jinkela_wire_20213),
        .dout(new_Jinkela_wire_20214)
    );

    or_bb _2199_ (
        .a(new_Jinkela_wire_10278),
        .b(new_Jinkela_wire_11836),
        .c(_1237_)
    );

    bfr new_Jinkela_buffer_16792 (
        .din(new_Jinkela_wire_20028),
        .dout(new_Jinkela_wire_20029)
    );

    or_ii _2200_ (
        .a(new_Jinkela_wire_10279),
        .b(new_Jinkela_wire_11837),
        .c(_1238_)
    );

    bfr new_Jinkela_buffer_16827 (
        .din(new_Jinkela_wire_20073),
        .dout(new_Jinkela_wire_20074)
    );

    or_ii _2201_ (
        .a(new_Jinkela_wire_11390),
        .b(new_Jinkela_wire_18798),
        .c(_1239_)
    );

    bfr new_Jinkela_buffer_16793 (
        .din(new_Jinkela_wire_20029),
        .dout(new_Jinkela_wire_20030)
    );

    and_ii _2202_ (
        .a(new_Jinkela_wire_714),
        .b(new_Jinkela_wire_6403),
        .c(_1240_)
    );

    bfr new_Jinkela_buffer_9908 (
        .din(new_Jinkela_wire_12027),
        .dout(new_Jinkela_wire_12028)
    );

    bfr new_Jinkela_buffer_9954 (
        .din(new_Jinkela_wire_12093),
        .dout(new_Jinkela_wire_12094)
    );

    bfr new_Jinkela_buffer_9909 (
        .din(new_Jinkela_wire_12028),
        .dout(new_Jinkela_wire_12029)
    );

    bfr new_Jinkela_buffer_9975 (
        .din(new_Jinkela_wire_12120),
        .dout(new_Jinkela_wire_12121)
    );

    bfr new_Jinkela_buffer_9910 (
        .din(new_Jinkela_wire_12029),
        .dout(new_Jinkela_wire_12030)
    );

    bfr new_Jinkela_buffer_9955 (
        .din(new_Jinkela_wire_12094),
        .dout(new_Jinkela_wire_12095)
    );

    bfr new_Jinkela_buffer_9911 (
        .din(new_Jinkela_wire_12030),
        .dout(new_Jinkela_wire_12031)
    );

    bfr new_Jinkela_buffer_9912 (
        .din(new_Jinkela_wire_12031),
        .dout(new_Jinkela_wire_12032)
    );

    bfr new_Jinkela_buffer_9956 (
        .din(new_Jinkela_wire_12095),
        .dout(new_Jinkela_wire_12096)
    );

    bfr new_Jinkela_buffer_9913 (
        .din(new_Jinkela_wire_12032),
        .dout(new_Jinkela_wire_12033)
    );

    bfr new_Jinkela_buffer_10030 (
        .din(new_Jinkela_wire_12175),
        .dout(new_Jinkela_wire_12176)
    );

    bfr new_Jinkela_buffer_9976 (
        .din(new_Jinkela_wire_12121),
        .dout(new_Jinkela_wire_12122)
    );

    bfr new_Jinkela_buffer_9914 (
        .din(new_Jinkela_wire_12033),
        .dout(new_Jinkela_wire_12034)
    );

    bfr new_Jinkela_buffer_9957 (
        .din(new_Jinkela_wire_12096),
        .dout(new_Jinkela_wire_12097)
    );

    bfr new_Jinkela_buffer_9915 (
        .din(new_Jinkela_wire_12034),
        .dout(new_Jinkela_wire_12035)
    );

    bfr new_Jinkela_buffer_9916 (
        .din(new_Jinkela_wire_12035),
        .dout(new_Jinkela_wire_12036)
    );

    bfr new_Jinkela_buffer_9958 (
        .din(new_Jinkela_wire_12097),
        .dout(new_Jinkela_wire_12098)
    );

    bfr new_Jinkela_buffer_9917 (
        .din(new_Jinkela_wire_12036),
        .dout(new_Jinkela_wire_12037)
    );

    bfr new_Jinkela_buffer_10075 (
        .din(new_Jinkela_wire_12224),
        .dout(new_Jinkela_wire_12225)
    );

    bfr new_Jinkela_buffer_9977 (
        .din(new_Jinkela_wire_12122),
        .dout(new_Jinkela_wire_12123)
    );

    bfr new_Jinkela_buffer_9918 (
        .din(new_Jinkela_wire_12037),
        .dout(new_Jinkela_wire_12038)
    );

    bfr new_Jinkela_buffer_9959 (
        .din(new_Jinkela_wire_12098),
        .dout(new_Jinkela_wire_12099)
    );

    bfr new_Jinkela_buffer_9919 (
        .din(new_Jinkela_wire_12038),
        .dout(new_Jinkela_wire_12039)
    );

    bfr new_Jinkela_buffer_9920 (
        .din(new_Jinkela_wire_12039),
        .dout(new_Jinkela_wire_12040)
    );

    bfr new_Jinkela_buffer_9960 (
        .din(new_Jinkela_wire_12099),
        .dout(new_Jinkela_wire_12100)
    );

    bfr new_Jinkela_buffer_9921 (
        .din(new_Jinkela_wire_12040),
        .dout(new_Jinkela_wire_12041)
    );

    bfr new_Jinkela_buffer_10031 (
        .din(new_Jinkela_wire_12176),
        .dout(new_Jinkela_wire_12177)
    );

    bfr new_Jinkela_buffer_9978 (
        .din(new_Jinkela_wire_12123),
        .dout(new_Jinkela_wire_12124)
    );

    bfr new_Jinkela_buffer_9922 (
        .din(new_Jinkela_wire_12041),
        .dout(new_Jinkela_wire_12042)
    );

    spl2 new_Jinkela_splitter_919 (
        .a(new_Jinkela_wire_12100),
        .b(new_Jinkela_wire_12101),
        .c(new_Jinkela_wire_12102)
    );

    spl2 new_Jinkela_splitter_909 (
        .a(new_Jinkela_wire_12042),
        .b(new_Jinkela_wire_12043),
        .c(new_Jinkela_wire_12044)
    );

    bfr new_Jinkela_buffer_9979 (
        .din(new_Jinkela_wire_12124),
        .dout(new_Jinkela_wire_12125)
    );

    spl2 new_Jinkela_splitter_927 (
        .a(_1077_),
        .b(new_Jinkela_wire_12337),
        .c(new_Jinkela_wire_12338)
    );

    bfr new_Jinkela_buffer_10032 (
        .din(new_Jinkela_wire_12177),
        .dout(new_Jinkela_wire_12178)
    );

    bfr new_Jinkela_buffer_9980 (
        .din(new_Jinkela_wire_12125),
        .dout(new_Jinkela_wire_12126)
    );

    bfr new_Jinkela_buffer_10076 (
        .din(new_Jinkela_wire_12225),
        .dout(new_Jinkela_wire_12226)
    );

    bfr new_Jinkela_buffer_9981 (
        .din(new_Jinkela_wire_12126),
        .dout(new_Jinkela_wire_12127)
    );

    bfr new_Jinkela_buffer_10033 (
        .din(new_Jinkela_wire_12178),
        .dout(new_Jinkela_wire_12179)
    );

    bfr new_Jinkela_buffer_9982 (
        .din(new_Jinkela_wire_12127),
        .dout(new_Jinkela_wire_12128)
    );

    bfr new_Jinkela_buffer_10177 (
        .din(new_Jinkela_wire_12332),
        .dout(new_Jinkela_wire_12333)
    );

    bfr new_Jinkela_buffer_9983 (
        .din(new_Jinkela_wire_12128),
        .dout(new_Jinkela_wire_12129)
    );

    spl2 new_Jinkela_splitter_928 (
        .a(_1727_),
        .b(new_Jinkela_wire_12339),
        .c(new_Jinkela_wire_12340)
    );

    bfr new_Jinkela_buffer_16898 (
        .din(new_Jinkela_wire_20150),
        .dout(new_Jinkela_wire_20151)
    );

    bfr new_Jinkela_buffer_16794 (
        .din(new_Jinkela_wire_20030),
        .dout(new_Jinkela_wire_20031)
    );

    bfr new_Jinkela_buffer_16828 (
        .din(new_Jinkela_wire_20074),
        .dout(new_Jinkela_wire_20075)
    );

    bfr new_Jinkela_buffer_16795 (
        .din(new_Jinkela_wire_20031),
        .dout(new_Jinkela_wire_20032)
    );

    spl2 new_Jinkela_splitter_1479 (
        .a(_1073_),
        .b(new_Jinkela_wire_20260),
        .c(new_Jinkela_wire_20261)
    );

    bfr new_Jinkela_buffer_16796 (
        .din(new_Jinkela_wire_20032),
        .dout(new_Jinkela_wire_20033)
    );

    bfr new_Jinkela_buffer_16829 (
        .din(new_Jinkela_wire_20075),
        .dout(new_Jinkela_wire_20076)
    );

    bfr new_Jinkela_buffer_16797 (
        .din(new_Jinkela_wire_20033),
        .dout(new_Jinkela_wire_20034)
    );

    bfr new_Jinkela_buffer_16899 (
        .din(new_Jinkela_wire_20151),
        .dout(new_Jinkela_wire_20152)
    );

    bfr new_Jinkela_buffer_16798 (
        .din(new_Jinkela_wire_20034),
        .dout(new_Jinkela_wire_20035)
    );

    bfr new_Jinkela_buffer_16830 (
        .din(new_Jinkela_wire_20076),
        .dout(new_Jinkela_wire_20077)
    );

    bfr new_Jinkela_buffer_16799 (
        .din(new_Jinkela_wire_20035),
        .dout(new_Jinkela_wire_20036)
    );

    bfr new_Jinkela_buffer_16958 (
        .din(new_Jinkela_wire_20214),
        .dout(new_Jinkela_wire_20215)
    );

    spl2 new_Jinkela_splitter_1467 (
        .a(new_Jinkela_wire_20036),
        .b(new_Jinkela_wire_20037),
        .c(new_Jinkela_wire_20038)
    );

    bfr new_Jinkela_buffer_16900 (
        .din(new_Jinkela_wire_20152),
        .dout(new_Jinkela_wire_20153)
    );

    bfr new_Jinkela_buffer_16831 (
        .din(new_Jinkela_wire_20077),
        .dout(new_Jinkela_wire_20078)
    );

    bfr new_Jinkela_buffer_16832 (
        .din(new_Jinkela_wire_20078),
        .dout(new_Jinkela_wire_20079)
    );

    bfr new_Jinkela_buffer_16999 (
        .din(_1327_),
        .dout(new_Jinkela_wire_20262)
    );

    bfr new_Jinkela_buffer_16833 (
        .din(new_Jinkela_wire_20079),
        .dout(new_Jinkela_wire_20080)
    );

    bfr new_Jinkela_buffer_16901 (
        .din(new_Jinkela_wire_20153),
        .dout(new_Jinkela_wire_20154)
    );

    bfr new_Jinkela_buffer_16834 (
        .din(new_Jinkela_wire_20080),
        .dout(new_Jinkela_wire_20081)
    );

    bfr new_Jinkela_buffer_16962 (
        .din(new_Jinkela_wire_20220),
        .dout(new_Jinkela_wire_20221)
    );

    bfr new_Jinkela_buffer_16835 (
        .din(new_Jinkela_wire_20081),
        .dout(new_Jinkela_wire_20082)
    );

    bfr new_Jinkela_buffer_16902 (
        .din(new_Jinkela_wire_20154),
        .dout(new_Jinkela_wire_20155)
    );

    bfr new_Jinkela_buffer_16836 (
        .din(new_Jinkela_wire_20082),
        .dout(new_Jinkela_wire_20083)
    );

    bfr new_Jinkela_buffer_16837 (
        .din(new_Jinkela_wire_20083),
        .dout(new_Jinkela_wire_20084)
    );

    bfr new_Jinkela_buffer_16903 (
        .din(new_Jinkela_wire_20155),
        .dout(new_Jinkela_wire_20156)
    );

    bfr new_Jinkela_buffer_16838 (
        .din(new_Jinkela_wire_20084),
        .dout(new_Jinkela_wire_20085)
    );

    bfr new_Jinkela_buffer_16963 (
        .din(new_Jinkela_wire_20221),
        .dout(new_Jinkela_wire_20222)
    );

    bfr new_Jinkela_buffer_16839 (
        .din(new_Jinkela_wire_20085),
        .dout(new_Jinkela_wire_20086)
    );

    bfr new_Jinkela_buffer_16904 (
        .din(new_Jinkela_wire_20156),
        .dout(new_Jinkela_wire_20157)
    );

    bfr new_Jinkela_buffer_16840 (
        .din(new_Jinkela_wire_20086),
        .dout(new_Jinkela_wire_20087)
    );

    spl2 new_Jinkela_splitter_1481 (
        .a(_1131_),
        .b(new_Jinkela_wire_20265),
        .c(new_Jinkela_wire_20266)
    );

    spl2 new_Jinkela_splitter_1480 (
        .a(_0962_),
        .b(new_Jinkela_wire_20263),
        .c(new_Jinkela_wire_20264)
    );

    bfr new_Jinkela_buffer_16841 (
        .din(new_Jinkela_wire_20087),
        .dout(new_Jinkela_wire_20088)
    );

    bfr new_Jinkela_buffer_16905 (
        .din(new_Jinkela_wire_20157),
        .dout(new_Jinkela_wire_20158)
    );

    bfr new_Jinkela_buffer_16842 (
        .din(new_Jinkela_wire_20088),
        .dout(new_Jinkela_wire_20089)
    );

    bfr new_Jinkela_buffer_16964 (
        .din(new_Jinkela_wire_20222),
        .dout(new_Jinkela_wire_20223)
    );

    bfr new_Jinkela_buffer_16843 (
        .din(new_Jinkela_wire_20089),
        .dout(new_Jinkela_wire_20090)
    );

    bfr new_Jinkela_buffer_16906 (
        .din(new_Jinkela_wire_20158),
        .dout(new_Jinkela_wire_20159)
    );

    bfr new_Jinkela_buffer_16844 (
        .din(new_Jinkela_wire_20090),
        .dout(new_Jinkela_wire_20091)
    );

    spl2 new_Jinkela_splitter_1482 (
        .a(_1343_),
        .b(new_Jinkela_wire_20267),
        .c(new_Jinkela_wire_20268)
    );

    spl2 new_Jinkela_splitter_1150 (
        .a(new_Jinkela_wire_15991),
        .b(new_Jinkela_wire_15992),
        .c(new_Jinkela_wire_15993)
    );

    bfr new_Jinkela_buffer_13432 (
        .din(new_Jinkela_wire_16045),
        .dout(new_Jinkela_wire_16046)
    );

    bfr new_Jinkela_buffer_13556 (
        .din(new_Jinkela_wire_16207),
        .dout(new_Jinkela_wire_16208)
    );

    bfr new_Jinkela_buffer_13501 (
        .din(new_Jinkela_wire_16138),
        .dout(new_Jinkela_wire_16139)
    );

    bfr new_Jinkela_buffer_13433 (
        .din(new_Jinkela_wire_16046),
        .dout(new_Jinkela_wire_16047)
    );

    bfr new_Jinkela_buffer_13552 (
        .din(new_Jinkela_wire_16197),
        .dout(new_Jinkela_wire_16198)
    );

    bfr new_Jinkela_buffer_13434 (
        .din(new_Jinkela_wire_16047),
        .dout(new_Jinkela_wire_16048)
    );

    bfr new_Jinkela_buffer_13502 (
        .din(new_Jinkela_wire_16139),
        .dout(new_Jinkela_wire_16140)
    );

    bfr new_Jinkela_buffer_13435 (
        .din(new_Jinkela_wire_16048),
        .dout(new_Jinkela_wire_16049)
    );

    bfr new_Jinkela_buffer_13555 (
        .din(_1743_),
        .dout(new_Jinkela_wire_16205)
    );

    bfr new_Jinkela_buffer_13436 (
        .din(new_Jinkela_wire_16049),
        .dout(new_Jinkela_wire_16050)
    );

    bfr new_Jinkela_buffer_13503 (
        .din(new_Jinkela_wire_16140),
        .dout(new_Jinkela_wire_16141)
    );

    bfr new_Jinkela_buffer_13437 (
        .din(new_Jinkela_wire_16050),
        .dout(new_Jinkela_wire_16051)
    );

    bfr new_Jinkela_buffer_13553 (
        .din(new_Jinkela_wire_16198),
        .dout(new_Jinkela_wire_16199)
    );

    bfr new_Jinkela_buffer_13438 (
        .din(new_Jinkela_wire_16051),
        .dout(new_Jinkela_wire_16052)
    );

    bfr new_Jinkela_buffer_13504 (
        .din(new_Jinkela_wire_16141),
        .dout(new_Jinkela_wire_16142)
    );

    bfr new_Jinkela_buffer_13439 (
        .din(new_Jinkela_wire_16052),
        .dout(new_Jinkela_wire_16053)
    );

    spl2 new_Jinkela_splitter_1175 (
        .a(_1079_),
        .b(new_Jinkela_wire_16212),
        .c(new_Jinkela_wire_16213)
    );

    spl2 new_Jinkela_splitter_1174 (
        .a(_0563_),
        .b(new_Jinkela_wire_16206),
        .c(new_Jinkela_wire_16207)
    );

    bfr new_Jinkela_buffer_13440 (
        .din(new_Jinkela_wire_16053),
        .dout(new_Jinkela_wire_16054)
    );

    bfr new_Jinkela_buffer_13505 (
        .din(new_Jinkela_wire_16142),
        .dout(new_Jinkela_wire_16143)
    );

    bfr new_Jinkela_buffer_13441 (
        .din(new_Jinkela_wire_16054),
        .dout(new_Jinkela_wire_16055)
    );

    bfr new_Jinkela_buffer_13442 (
        .din(new_Jinkela_wire_16055),
        .dout(new_Jinkela_wire_16056)
    );

    bfr new_Jinkela_buffer_13506 (
        .din(new_Jinkela_wire_16143),
        .dout(new_Jinkela_wire_16144)
    );

    bfr new_Jinkela_buffer_13443 (
        .din(new_Jinkela_wire_16056),
        .dout(new_Jinkela_wire_16057)
    );

    bfr new_Jinkela_buffer_13560 (
        .din(_0581_),
        .dout(new_Jinkela_wire_16214)
    );

    bfr new_Jinkela_buffer_13444 (
        .din(new_Jinkela_wire_16057),
        .dout(new_Jinkela_wire_16058)
    );

    bfr new_Jinkela_buffer_13507 (
        .din(new_Jinkela_wire_16144),
        .dout(new_Jinkela_wire_16145)
    );

    bfr new_Jinkela_buffer_13445 (
        .din(new_Jinkela_wire_16058),
        .dout(new_Jinkela_wire_16059)
    );

    bfr new_Jinkela_buffer_13446 (
        .din(new_Jinkela_wire_16059),
        .dout(new_Jinkela_wire_16060)
    );

    bfr new_Jinkela_buffer_13508 (
        .din(new_Jinkela_wire_16145),
        .dout(new_Jinkela_wire_16146)
    );

    bfr new_Jinkela_buffer_13447 (
        .din(new_Jinkela_wire_16060),
        .dout(new_Jinkela_wire_16061)
    );

    bfr new_Jinkela_buffer_13557 (
        .din(new_Jinkela_wire_16208),
        .dout(new_Jinkela_wire_16209)
    );

    bfr new_Jinkela_buffer_13448 (
        .din(new_Jinkela_wire_16061),
        .dout(new_Jinkela_wire_16062)
    );

    bfr new_Jinkela_buffer_13509 (
        .din(new_Jinkela_wire_16146),
        .dout(new_Jinkela_wire_16147)
    );

    bfr new_Jinkela_buffer_13449 (
        .din(new_Jinkela_wire_16062),
        .dout(new_Jinkela_wire_16063)
    );

    bfr new_Jinkela_buffer_13561 (
        .din(_0326_),
        .dout(new_Jinkela_wire_16217)
    );

    spl2 new_Jinkela_splitter_1176 (
        .a(_0602_),
        .b(new_Jinkela_wire_16215),
        .c(new_Jinkela_wire_16216)
    );

    bfr new_Jinkela_buffer_13450 (
        .din(new_Jinkela_wire_16063),
        .dout(new_Jinkela_wire_16064)
    );

    bfr new_Jinkela_buffer_13510 (
        .din(new_Jinkela_wire_16147),
        .dout(new_Jinkela_wire_16148)
    );

    bfr new_Jinkela_buffer_13451 (
        .din(new_Jinkela_wire_16064),
        .dout(new_Jinkela_wire_16065)
    );

    bfr new_Jinkela_buffer_13558 (
        .din(new_Jinkela_wire_16209),
        .dout(new_Jinkela_wire_16210)
    );

    bfr new_Jinkela_buffer_6450 (
        .din(new_Jinkela_wire_8141),
        .dout(new_Jinkela_wire_8142)
    );

    bfr new_Jinkela_buffer_6451 (
        .din(new_Jinkela_wire_8142),
        .dout(new_Jinkela_wire_8143)
    );

    bfr new_Jinkela_buffer_6575 (
        .din(new_Jinkela_wire_8284),
        .dout(new_Jinkela_wire_8285)
    );

    bfr new_Jinkela_buffer_6505 (
        .din(new_Jinkela_wire_8204),
        .dout(new_Jinkela_wire_8205)
    );

    bfr new_Jinkela_buffer_6452 (
        .din(new_Jinkela_wire_8143),
        .dout(new_Jinkela_wire_8144)
    );

    bfr new_Jinkela_buffer_6453 (
        .din(new_Jinkela_wire_8144),
        .dout(new_Jinkela_wire_8145)
    );

    bfr new_Jinkela_buffer_6517 (
        .din(new_Jinkela_wire_8216),
        .dout(new_Jinkela_wire_8217)
    );

    bfr new_Jinkela_buffer_6506 (
        .din(new_Jinkela_wire_8205),
        .dout(new_Jinkela_wire_8206)
    );

    bfr new_Jinkela_buffer_6454 (
        .din(new_Jinkela_wire_8145),
        .dout(new_Jinkela_wire_8146)
    );

    bfr new_Jinkela_buffer_6455 (
        .din(new_Jinkela_wire_8146),
        .dout(new_Jinkela_wire_8147)
    );

    bfr new_Jinkela_buffer_6456 (
        .din(new_Jinkela_wire_8147),
        .dout(new_Jinkela_wire_8148)
    );

    bfr new_Jinkela_buffer_6518 (
        .din(new_Jinkela_wire_8217),
        .dout(new_Jinkela_wire_8218)
    );

    bfr new_Jinkela_buffer_6457 (
        .din(new_Jinkela_wire_8148),
        .dout(new_Jinkela_wire_8149)
    );

    bfr new_Jinkela_buffer_6576 (
        .din(new_Jinkela_wire_8285),
        .dout(new_Jinkela_wire_8286)
    );

    bfr new_Jinkela_buffer_6458 (
        .din(new_Jinkela_wire_8149),
        .dout(new_Jinkela_wire_8150)
    );

    bfr new_Jinkela_buffer_6519 (
        .din(new_Jinkela_wire_8218),
        .dout(new_Jinkela_wire_8219)
    );

    bfr new_Jinkela_buffer_6459 (
        .din(new_Jinkela_wire_8150),
        .dout(new_Jinkela_wire_8151)
    );

    bfr new_Jinkela_buffer_6578 (
        .din(_0036_),
        .dout(new_Jinkela_wire_8294)
    );

    bfr new_Jinkela_buffer_6460 (
        .din(new_Jinkela_wire_8151),
        .dout(new_Jinkela_wire_8152)
    );

    bfr new_Jinkela_buffer_6520 (
        .din(new_Jinkela_wire_8219),
        .dout(new_Jinkela_wire_8220)
    );

    bfr new_Jinkela_buffer_6461 (
        .din(new_Jinkela_wire_8152),
        .dout(new_Jinkela_wire_8153)
    );

    bfr new_Jinkela_buffer_6577 (
        .din(new_Jinkela_wire_8286),
        .dout(new_Jinkela_wire_8287)
    );

    bfr new_Jinkela_buffer_6462 (
        .din(new_Jinkela_wire_8153),
        .dout(new_Jinkela_wire_8154)
    );

    bfr new_Jinkela_buffer_6521 (
        .din(new_Jinkela_wire_8220),
        .dout(new_Jinkela_wire_8221)
    );

    bfr new_Jinkela_buffer_6463 (
        .din(new_Jinkela_wire_8154),
        .dout(new_Jinkela_wire_8155)
    );

    bfr new_Jinkela_buffer_6579 (
        .din(_0853_),
        .dout(new_Jinkela_wire_8297)
    );

    spl2 new_Jinkela_splitter_707 (
        .a(_1692_),
        .b(new_Jinkela_wire_8295),
        .c(new_Jinkela_wire_8296)
    );

    bfr new_Jinkela_buffer_6464 (
        .din(new_Jinkela_wire_8155),
        .dout(new_Jinkela_wire_8156)
    );

    bfr new_Jinkela_buffer_6522 (
        .din(new_Jinkela_wire_8221),
        .dout(new_Jinkela_wire_8222)
    );

    bfr new_Jinkela_buffer_6465 (
        .din(new_Jinkela_wire_8156),
        .dout(new_Jinkela_wire_8157)
    );

    spl2 new_Jinkela_splitter_710 (
        .a(_0298_),
        .b(new_Jinkela_wire_8361),
        .c(new_Jinkela_wire_8362)
    );

    bfr new_Jinkela_buffer_6466 (
        .din(new_Jinkela_wire_8157),
        .dout(new_Jinkela_wire_8158)
    );

    bfr new_Jinkela_buffer_6523 (
        .din(new_Jinkela_wire_8222),
        .dout(new_Jinkela_wire_8223)
    );

    bfr new_Jinkela_buffer_6467 (
        .din(new_Jinkela_wire_8158),
        .dout(new_Jinkela_wire_8159)
    );

    bfr new_Jinkela_buffer_6581 (
        .din(_1008_),
        .dout(new_Jinkela_wire_8301)
    );

    bfr new_Jinkela_buffer_6468 (
        .din(new_Jinkela_wire_8159),
        .dout(new_Jinkela_wire_8160)
    );

    bfr new_Jinkela_buffer_6524 (
        .din(new_Jinkela_wire_8223),
        .dout(new_Jinkela_wire_8224)
    );

    bfr new_Jinkela_buffer_6469 (
        .din(new_Jinkela_wire_8160),
        .dout(new_Jinkela_wire_8161)
    );

    bfr new_Jinkela_buffer_6580 (
        .din(new_Jinkela_wire_8297),
        .dout(new_Jinkela_wire_8298)
    );

    bfr new_Jinkela_buffer_6470 (
        .din(new_Jinkela_wire_8161),
        .dout(new_Jinkela_wire_8162)
    );

    bfr new_Jinkela_buffer_6525 (
        .din(new_Jinkela_wire_8224),
        .dout(new_Jinkela_wire_8225)
    );

    bfr new_Jinkela_buffer_3098 (
        .din(new_Jinkela_wire_4187),
        .dout(new_Jinkela_wire_4188)
    );

    and_bb _2203_ (
        .a(new_Jinkela_wire_715),
        .b(new_Jinkela_wire_6404),
        .c(_1241_)
    );

    bfr new_Jinkela_buffer_3052 (
        .din(new_Jinkela_wire_4133),
        .dout(new_Jinkela_wire_4134)
    );

    or_bb _2204_ (
        .a(new_Jinkela_wire_20046),
        .b(new_Jinkela_wire_716),
        .c(_1242_)
    );

    bfr new_Jinkela_buffer_3164 (
        .din(new_Jinkela_wire_4267),
        .dout(new_Jinkela_wire_4268)
    );

    or_bb _2205_ (
        .a(new_Jinkela_wire_5880),
        .b(new_Jinkela_wire_14663),
        .c(_1243_)
    );

    bfr new_Jinkela_buffer_3156 (
        .din(new_Jinkela_wire_4259),
        .dout(new_Jinkela_wire_4260)
    );

    bfr new_Jinkela_buffer_3053 (
        .din(new_Jinkela_wire_4134),
        .dout(new_Jinkela_wire_4135)
    );

    or_ii _2206_ (
        .a(new_Jinkela_wire_5881),
        .b(new_Jinkela_wire_14664),
        .c(_1244_)
    );

    bfr new_Jinkela_buffer_3099 (
        .din(new_Jinkela_wire_4188),
        .dout(new_Jinkela_wire_4189)
    );

    or_ii _2207_ (
        .a(new_Jinkela_wire_8588),
        .b(new_Jinkela_wire_13972),
        .c(_1245_)
    );

    bfr new_Jinkela_buffer_3054 (
        .din(new_Jinkela_wire_4135),
        .dout(new_Jinkela_wire_4136)
    );

    and_ii _2208_ (
        .a(new_Jinkela_wire_14281),
        .b(new_Jinkela_wire_6802),
        .c(_1246_)
    );

    and_bb _2209_ (
        .a(new_Jinkela_wire_14282),
        .b(new_Jinkela_wire_6803),
        .c(_1247_)
    );

    bfr new_Jinkela_buffer_3055 (
        .din(new_Jinkela_wire_4136),
        .dout(new_Jinkela_wire_4137)
    );

    or_bb _2210_ (
        .a(new_Jinkela_wire_3552),
        .b(new_Jinkela_wire_5147),
        .c(_1248_)
    );

    bfr new_Jinkela_buffer_3100 (
        .din(new_Jinkela_wire_4189),
        .dout(new_Jinkela_wire_4190)
    );

    or_bb _2211_ (
        .a(new_Jinkela_wire_11342),
        .b(new_Jinkela_wire_13314),
        .c(_1249_)
    );

    bfr new_Jinkela_buffer_3056 (
        .din(new_Jinkela_wire_4137),
        .dout(new_Jinkela_wire_4138)
    );

    or_ii _2212_ (
        .a(new_Jinkela_wire_11343),
        .b(new_Jinkela_wire_13315),
        .c(_1250_)
    );

    or_ii _2213_ (
        .a(new_Jinkela_wire_15729),
        .b(new_Jinkela_wire_16002),
        .c(_1251_)
    );

    bfr new_Jinkela_buffer_3157 (
        .din(new_Jinkela_wire_4260),
        .dout(new_Jinkela_wire_4261)
    );

    bfr new_Jinkela_buffer_3057 (
        .din(new_Jinkela_wire_4138),
        .dout(new_Jinkela_wire_4139)
    );

    and_ii _2214_ (
        .a(new_Jinkela_wire_17975),
        .b(new_Jinkela_wire_11016),
        .c(_1252_)
    );

    bfr new_Jinkela_buffer_3101 (
        .din(new_Jinkela_wire_4190),
        .dout(new_Jinkela_wire_4191)
    );

    and_bb _2215_ (
        .a(new_Jinkela_wire_17976),
        .b(new_Jinkela_wire_11017),
        .c(_1253_)
    );

    bfr new_Jinkela_buffer_3058 (
        .din(new_Jinkela_wire_4139),
        .dout(new_Jinkela_wire_4140)
    );

    or_bb _2216_ (
        .a(new_Jinkela_wire_10681),
        .b(new_Jinkela_wire_17671),
        .c(_1254_)
    );

    or_bb _2217_ (
        .a(new_Jinkela_wire_3255),
        .b(new_Jinkela_wire_2789),
        .c(_1255_)
    );

    bfr new_Jinkela_buffer_3182 (
        .din(_1274_),
        .dout(new_Jinkela_wire_4292)
    );

    bfr new_Jinkela_buffer_3059 (
        .din(new_Jinkela_wire_4140),
        .dout(new_Jinkela_wire_4141)
    );

    or_ii _2218_ (
        .a(new_Jinkela_wire_3256),
        .b(new_Jinkela_wire_2790),
        .c(_1256_)
    );

    bfr new_Jinkela_buffer_3102 (
        .din(new_Jinkela_wire_4191),
        .dout(new_Jinkela_wire_4192)
    );

    or_ii _2219_ (
        .a(new_Jinkela_wire_20133),
        .b(new_Jinkela_wire_20277),
        .c(_1257_)
    );

    bfr new_Jinkela_buffer_3060 (
        .din(new_Jinkela_wire_4141),
        .dout(new_Jinkela_wire_4142)
    );

    and_ii _2220_ (
        .a(new_Jinkela_wire_7289),
        .b(new_Jinkela_wire_9857),
        .c(_1258_)
    );

    bfr new_Jinkela_buffer_3165 (
        .din(new_Jinkela_wire_4268),
        .dout(new_Jinkela_wire_4269)
    );

    and_bb _2221_ (
        .a(new_Jinkela_wire_7290),
        .b(new_Jinkela_wire_9858),
        .c(_1259_)
    );

    bfr new_Jinkela_buffer_3158 (
        .din(new_Jinkela_wire_4261),
        .dout(new_Jinkela_wire_4262)
    );

    bfr new_Jinkela_buffer_3061 (
        .din(new_Jinkela_wire_4142),
        .dout(new_Jinkela_wire_4143)
    );

    or_bb _2222_ (
        .a(new_Jinkela_wire_11020),
        .b(new_Jinkela_wire_8025),
        .c(_1260_)
    );

    bfr new_Jinkela_buffer_3103 (
        .din(new_Jinkela_wire_4192),
        .dout(new_Jinkela_wire_4193)
    );

    or_bb _2223_ (
        .a(new_Jinkela_wire_10205),
        .b(new_Jinkela_wire_2317),
        .c(_1261_)
    );

    bfr new_Jinkela_buffer_3062 (
        .din(new_Jinkela_wire_4143),
        .dout(new_Jinkela_wire_4144)
    );

    or_ii _2224_ (
        .a(new_Jinkela_wire_10206),
        .b(new_Jinkela_wire_2318),
        .c(_1262_)
    );

    or_ii _2225_ (
        .a(new_Jinkela_wire_7736),
        .b(new_Jinkela_wire_846),
        .c(_1263_)
    );

    bfr new_Jinkela_buffer_3063 (
        .din(new_Jinkela_wire_4144),
        .dout(new_Jinkela_wire_4145)
    );

    and_ii _2226_ (
        .a(new_Jinkela_wire_20383),
        .b(new_Jinkela_wire_7051),
        .c(_1264_)
    );

    bfr new_Jinkela_buffer_3104 (
        .din(new_Jinkela_wire_4193),
        .dout(new_Jinkela_wire_4194)
    );

    and_bb _2227_ (
        .a(new_Jinkela_wire_20384),
        .b(new_Jinkela_wire_7052),
        .c(_1265_)
    );

    bfr new_Jinkela_buffer_3064 (
        .din(new_Jinkela_wire_4145),
        .dout(new_Jinkela_wire_4146)
    );

    or_bb _2228_ (
        .a(new_Jinkela_wire_21194),
        .b(new_Jinkela_wire_13323),
        .c(_1266_)
    );

    or_bb _2229_ (
        .a(new_Jinkela_wire_17992),
        .b(new_Jinkela_wire_19786),
        .c(_1267_)
    );

    bfr new_Jinkela_buffer_3159 (
        .din(new_Jinkela_wire_4262),
        .dout(new_Jinkela_wire_4263)
    );

    bfr new_Jinkela_buffer_3065 (
        .din(new_Jinkela_wire_4146),
        .dout(new_Jinkela_wire_4147)
    );

    or_ii _2230_ (
        .a(new_Jinkela_wire_17993),
        .b(new_Jinkela_wire_19787),
        .c(_1268_)
    );

    bfr new_Jinkela_buffer_3105 (
        .din(new_Jinkela_wire_4194),
        .dout(new_Jinkela_wire_4195)
    );

    or_ii _2231_ (
        .a(new_Jinkela_wire_6523),
        .b(new_Jinkela_wire_17788),
        .c(_1269_)
    );

    bfr new_Jinkela_buffer_3066 (
        .din(new_Jinkela_wire_4147),
        .dout(new_Jinkela_wire_4148)
    );

    and_ii _2232_ (
        .a(new_Jinkela_wire_12520),
        .b(new_Jinkela_wire_16599),
        .c(_1270_)
    );

    and_bb _2233_ (
        .a(new_Jinkela_wire_12521),
        .b(new_Jinkela_wire_16600),
        .c(_1271_)
    );

    bfr new_Jinkela_buffer_3183 (
        .din(_1445_),
        .dout(new_Jinkela_wire_4293)
    );

    bfr new_Jinkela_buffer_3067 (
        .din(new_Jinkela_wire_4148),
        .dout(new_Jinkela_wire_4149)
    );

    or_bb _2234_ (
        .a(new_Jinkela_wire_9019),
        .b(new_Jinkela_wire_3553),
        .c(_1272_)
    );

    bfr new_Jinkela_buffer_3106 (
        .din(new_Jinkela_wire_4195),
        .dout(new_Jinkela_wire_4196)
    );

    or_bb _2235_ (
        .a(new_Jinkela_wire_11440),
        .b(new_Jinkela_wire_21216),
        .c(_1273_)
    );

    bfr new_Jinkela_buffer_3068 (
        .din(new_Jinkela_wire_4149),
        .dout(new_Jinkela_wire_4150)
    );

    and_bb _2236_ (
        .a(new_Jinkela_wire_11441),
        .b(new_Jinkela_wire_21217),
        .c(_1274_)
    );

    bfr new_Jinkela_buffer_3166 (
        .din(new_Jinkela_wire_4269),
        .dout(new_Jinkela_wire_4270)
    );

    or_bi _2237_ (
        .a(new_Jinkela_wire_4292),
        .b(new_Jinkela_wire_1261),
        .c(_1275_)
    );

    bfr new_Jinkela_buffer_3160 (
        .din(new_Jinkela_wire_4263),
        .dout(new_Jinkela_wire_4264)
    );

    bfr new_Jinkela_buffer_3069 (
        .din(new_Jinkela_wire_4150),
        .dout(new_Jinkela_wire_4151)
    );

    and_ii _2238_ (
        .a(new_Jinkela_wire_19077),
        .b(new_Jinkela_wire_2785),
        .c(_1276_)
    );

    bfr new_Jinkela_buffer_3107 (
        .din(new_Jinkela_wire_4196),
        .dout(new_Jinkela_wire_4197)
    );

    and_bb _2239_ (
        .a(new_Jinkela_wire_19078),
        .b(new_Jinkela_wire_2786),
        .c(_1277_)
    );

    bfr new_Jinkela_buffer_3070 (
        .din(new_Jinkela_wire_4151),
        .dout(new_Jinkela_wire_4152)
    );

    or_bb _2240_ (
        .a(new_Jinkela_wire_8693),
        .b(new_Jinkela_wire_7298),
        .c(new_net_3922)
    );

    and_bb _2241_ (
        .a(new_Jinkela_wire_585),
        .b(new_Jinkela_wire_347),
        .c(_1278_)
    );

    bfr new_Jinkela_buffer_3071 (
        .din(new_Jinkela_wire_4152),
        .dout(new_Jinkela_wire_4153)
    );

    and_bi _2242_ (
        .a(new_Jinkela_wire_1266),
        .b(new_Jinkela_wire_7299),
        .c(_1279_)
    );

    bfr new_Jinkela_buffer_3108 (
        .din(new_Jinkela_wire_4197),
        .dout(new_Jinkela_wire_4198)
    );

    and_bb _2243_ (
        .a(new_Jinkela_wire_103),
        .b(new_Jinkela_wire_123),
        .c(_1280_)
    );

    bfr new_Jinkela_buffer_3072 (
        .din(new_Jinkela_wire_4153),
        .dout(new_Jinkela_wire_4154)
    );

    and_bi _2244_ (
        .a(new_Jinkela_wire_17793),
        .b(new_Jinkela_wire_3554),
        .c(_1281_)
    );

    bfr new_Jinkela_buffer_6471 (
        .din(new_Jinkela_wire_8162),
        .dout(new_Jinkela_wire_8163)
    );

    bfr new_Jinkela_buffer_16845 (
        .din(new_Jinkela_wire_20091),
        .dout(new_Jinkela_wire_20092)
    );

    bfr new_Jinkela_buffer_16907 (
        .din(new_Jinkela_wire_20159),
        .dout(new_Jinkela_wire_20160)
    );

    bfr new_Jinkela_buffer_6639 (
        .din(_0519_),
        .dout(new_Jinkela_wire_8363)
    );

    bfr new_Jinkela_buffer_6472 (
        .din(new_Jinkela_wire_8163),
        .dout(new_Jinkela_wire_8164)
    );

    bfr new_Jinkela_buffer_16846 (
        .din(new_Jinkela_wire_20092),
        .dout(new_Jinkela_wire_20093)
    );

    bfr new_Jinkela_buffer_6526 (
        .din(new_Jinkela_wire_8225),
        .dout(new_Jinkela_wire_8226)
    );

    bfr new_Jinkela_buffer_16965 (
        .din(new_Jinkela_wire_20223),
        .dout(new_Jinkela_wire_20224)
    );

    bfr new_Jinkela_buffer_6473 (
        .din(new_Jinkela_wire_8164),
        .dout(new_Jinkela_wire_8165)
    );

    bfr new_Jinkela_buffer_16847 (
        .din(new_Jinkela_wire_20093),
        .dout(new_Jinkela_wire_20094)
    );

    spl2 new_Jinkela_splitter_708 (
        .a(new_Jinkela_wire_8298),
        .b(new_Jinkela_wire_8299),
        .c(new_Jinkela_wire_8300)
    );

    bfr new_Jinkela_buffer_16908 (
        .din(new_Jinkela_wire_20160),
        .dout(new_Jinkela_wire_20161)
    );

    bfr new_Jinkela_buffer_6474 (
        .din(new_Jinkela_wire_8165),
        .dout(new_Jinkela_wire_8166)
    );

    bfr new_Jinkela_buffer_16848 (
        .din(new_Jinkela_wire_20094),
        .dout(new_Jinkela_wire_20095)
    );

    bfr new_Jinkela_buffer_6527 (
        .din(new_Jinkela_wire_8226),
        .dout(new_Jinkela_wire_8227)
    );

    bfr new_Jinkela_buffer_6475 (
        .din(new_Jinkela_wire_8166),
        .dout(new_Jinkela_wire_8167)
    );

    bfr new_Jinkela_buffer_16849 (
        .din(new_Jinkela_wire_20095),
        .dout(new_Jinkela_wire_20096)
    );

    bfr new_Jinkela_buffer_16909 (
        .din(new_Jinkela_wire_20161),
        .dout(new_Jinkela_wire_20162)
    );

    bfr new_Jinkela_buffer_6476 (
        .din(new_Jinkela_wire_8167),
        .dout(new_Jinkela_wire_8168)
    );

    bfr new_Jinkela_buffer_16850 (
        .din(new_Jinkela_wire_20096),
        .dout(new_Jinkela_wire_20097)
    );

    bfr new_Jinkela_buffer_6528 (
        .din(new_Jinkela_wire_8227),
        .dout(new_Jinkela_wire_8228)
    );

    bfr new_Jinkela_buffer_16966 (
        .din(new_Jinkela_wire_20224),
        .dout(new_Jinkela_wire_20225)
    );

    bfr new_Jinkela_buffer_6477 (
        .din(new_Jinkela_wire_8168),
        .dout(new_Jinkela_wire_8169)
    );

    bfr new_Jinkela_buffer_16851 (
        .din(new_Jinkela_wire_20097),
        .dout(new_Jinkela_wire_20098)
    );

    bfr new_Jinkela_buffer_6582 (
        .din(new_Jinkela_wire_8301),
        .dout(new_Jinkela_wire_8302)
    );

    bfr new_Jinkela_buffer_16910 (
        .din(new_Jinkela_wire_20162),
        .dout(new_Jinkela_wire_20163)
    );

    bfr new_Jinkela_buffer_6478 (
        .din(new_Jinkela_wire_8169),
        .dout(new_Jinkela_wire_8170)
    );

    bfr new_Jinkela_buffer_16852 (
        .din(new_Jinkela_wire_20098),
        .dout(new_Jinkela_wire_20099)
    );

    bfr new_Jinkela_buffer_6529 (
        .din(new_Jinkela_wire_8228),
        .dout(new_Jinkela_wire_8229)
    );

    spl2 new_Jinkela_splitter_1483 (
        .a(_0478_),
        .b(new_Jinkela_wire_20269),
        .c(new_Jinkela_wire_20270)
    );

    bfr new_Jinkela_buffer_6479 (
        .din(new_Jinkela_wire_8170),
        .dout(new_Jinkela_wire_8171)
    );

    bfr new_Jinkela_buffer_16853 (
        .din(new_Jinkela_wire_20099),
        .dout(new_Jinkela_wire_20100)
    );

    bfr new_Jinkela_buffer_6583 (
        .din(new_Jinkela_wire_8302),
        .dout(new_Jinkela_wire_8303)
    );

    bfr new_Jinkela_buffer_16911 (
        .din(new_Jinkela_wire_20163),
        .dout(new_Jinkela_wire_20164)
    );

    bfr new_Jinkela_buffer_6480 (
        .din(new_Jinkela_wire_8171),
        .dout(new_Jinkela_wire_8172)
    );

    bfr new_Jinkela_buffer_16854 (
        .din(new_Jinkela_wire_20100),
        .dout(new_Jinkela_wire_20101)
    );

    bfr new_Jinkela_buffer_6530 (
        .din(new_Jinkela_wire_8229),
        .dout(new_Jinkela_wire_8230)
    );

    bfr new_Jinkela_buffer_16967 (
        .din(new_Jinkela_wire_20225),
        .dout(new_Jinkela_wire_20226)
    );

    bfr new_Jinkela_buffer_6481 (
        .din(new_Jinkela_wire_8172),
        .dout(new_Jinkela_wire_8173)
    );

    bfr new_Jinkela_buffer_16855 (
        .din(new_Jinkela_wire_20101),
        .dout(new_Jinkela_wire_20102)
    );

    bfr new_Jinkela_buffer_6736 (
        .din(_0011_),
        .dout(new_Jinkela_wire_8462)
    );

    bfr new_Jinkela_buffer_16912 (
        .din(new_Jinkela_wire_20164),
        .dout(new_Jinkela_wire_20165)
    );

    bfr new_Jinkela_buffer_6640 (
        .din(_0533_),
        .dout(new_Jinkela_wire_8364)
    );

    bfr new_Jinkela_buffer_6482 (
        .din(new_Jinkela_wire_8173),
        .dout(new_Jinkela_wire_8174)
    );

    bfr new_Jinkela_buffer_16856 (
        .din(new_Jinkela_wire_20102),
        .dout(new_Jinkela_wire_20103)
    );

    bfr new_Jinkela_buffer_6531 (
        .din(new_Jinkela_wire_8230),
        .dout(new_Jinkela_wire_8231)
    );

    spl2 new_Jinkela_splitter_1486 (
        .a(_1255_),
        .b(new_Jinkela_wire_20277),
        .c(new_Jinkela_wire_20278)
    );

    bfr new_Jinkela_buffer_17000 (
        .din(_0004_),
        .dout(new_Jinkela_wire_20271)
    );

    spl2 new_Jinkela_splitter_695 (
        .a(new_Jinkela_wire_8174),
        .b(new_Jinkela_wire_8175),
        .c(new_Jinkela_wire_8176)
    );

    bfr new_Jinkela_buffer_16857 (
        .din(new_Jinkela_wire_20103),
        .dout(new_Jinkela_wire_20104)
    );

    bfr new_Jinkela_buffer_6532 (
        .din(new_Jinkela_wire_8231),
        .dout(new_Jinkela_wire_8232)
    );

    bfr new_Jinkela_buffer_16913 (
        .din(new_Jinkela_wire_20165),
        .dout(new_Jinkela_wire_20166)
    );

    bfr new_Jinkela_buffer_6584 (
        .din(new_Jinkela_wire_8303),
        .dout(new_Jinkela_wire_8304)
    );

    bfr new_Jinkela_buffer_16858 (
        .din(new_Jinkela_wire_20104),
        .dout(new_Jinkela_wire_20105)
    );

    bfr new_Jinkela_buffer_16968 (
        .din(new_Jinkela_wire_20226),
        .dout(new_Jinkela_wire_20227)
    );

    spl2 new_Jinkela_splitter_713 (
        .a(_0094_),
        .b(new_Jinkela_wire_8480),
        .c(new_Jinkela_wire_8481)
    );

    bfr new_Jinkela_buffer_6533 (
        .din(new_Jinkela_wire_8232),
        .dout(new_Jinkela_wire_8233)
    );

    bfr new_Jinkela_buffer_16859 (
        .din(new_Jinkela_wire_20105),
        .dout(new_Jinkela_wire_20106)
    );

    bfr new_Jinkela_buffer_6585 (
        .din(new_Jinkela_wire_8304),
        .dout(new_Jinkela_wire_8305)
    );

    bfr new_Jinkela_buffer_16914 (
        .din(new_Jinkela_wire_20166),
        .dout(new_Jinkela_wire_20167)
    );

    bfr new_Jinkela_buffer_6534 (
        .din(new_Jinkela_wire_8233),
        .dout(new_Jinkela_wire_8234)
    );

    bfr new_Jinkela_buffer_16860 (
        .din(new_Jinkela_wire_20106),
        .dout(new_Jinkela_wire_20107)
    );

    bfr new_Jinkela_buffer_6641 (
        .din(new_Jinkela_wire_8364),
        .dout(new_Jinkela_wire_8365)
    );

    spl2 new_Jinkela_splitter_1485 (
        .a(_1386_),
        .b(new_Jinkela_wire_20275),
        .c(new_Jinkela_wire_20276)
    );

    bfr new_Jinkela_buffer_6535 (
        .din(new_Jinkela_wire_8234),
        .dout(new_Jinkela_wire_8235)
    );

    bfr new_Jinkela_buffer_16861 (
        .din(new_Jinkela_wire_20107),
        .dout(new_Jinkela_wire_20108)
    );

    bfr new_Jinkela_buffer_6586 (
        .din(new_Jinkela_wire_8305),
        .dout(new_Jinkela_wire_8306)
    );

    bfr new_Jinkela_buffer_16915 (
        .din(new_Jinkela_wire_20167),
        .dout(new_Jinkela_wire_20168)
    );

    bfr new_Jinkela_buffer_6536 (
        .din(new_Jinkela_wire_8235),
        .dout(new_Jinkela_wire_8236)
    );

    bfr new_Jinkela_buffer_16862 (
        .din(new_Jinkela_wire_20108),
        .dout(new_Jinkela_wire_20109)
    );

    bfr new_Jinkela_buffer_16969 (
        .din(new_Jinkela_wire_20227),
        .dout(new_Jinkela_wire_20228)
    );

    spl2 new_Jinkela_splitter_714 (
        .a(_0057_),
        .b(new_Jinkela_wire_8482),
        .c(new_Jinkela_wire_8483)
    );

    bfr new_Jinkela_buffer_6537 (
        .din(new_Jinkela_wire_8236),
        .dout(new_Jinkela_wire_8237)
    );

    bfr new_Jinkela_buffer_16863 (
        .din(new_Jinkela_wire_20109),
        .dout(new_Jinkela_wire_20110)
    );

    bfr new_Jinkela_buffer_6587 (
        .din(new_Jinkela_wire_8306),
        .dout(new_Jinkela_wire_8307)
    );

    bfr new_Jinkela_buffer_16916 (
        .din(new_Jinkela_wire_20168),
        .dout(new_Jinkela_wire_20169)
    );

    bfr new_Jinkela_buffer_6538 (
        .din(new_Jinkela_wire_8237),
        .dout(new_Jinkela_wire_8238)
    );

    bfr new_Jinkela_buffer_16864 (
        .din(new_Jinkela_wire_20110),
        .dout(new_Jinkela_wire_20111)
    );

    bfr new_Jinkela_buffer_6642 (
        .din(new_Jinkela_wire_8365),
        .dout(new_Jinkela_wire_8366)
    );

    bfr new_Jinkela_buffer_17001 (
        .din(new_Jinkela_wire_20271),
        .dout(new_Jinkela_wire_20272)
    );

    bfr new_Jinkela_buffer_6539 (
        .din(new_Jinkela_wire_8238),
        .dout(new_Jinkela_wire_8239)
    );

    bfr new_Jinkela_buffer_16865 (
        .din(new_Jinkela_wire_20111),
        .dout(new_Jinkela_wire_20112)
    );

    bfr new_Jinkela_buffer_6588 (
        .din(new_Jinkela_wire_8307),
        .dout(new_Jinkela_wire_8308)
    );

    bfr new_Jinkela_buffer_16917 (
        .din(new_Jinkela_wire_20169),
        .dout(new_Jinkela_wire_20170)
    );

    bfr new_Jinkela_buffer_3178 (
        .din(new_Jinkela_wire_4287),
        .dout(new_Jinkela_wire_4288)
    );

    bfr new_Jinkela_buffer_10034 (
        .din(new_Jinkela_wire_12179),
        .dout(new_Jinkela_wire_12180)
    );

    bfr new_Jinkela_buffer_13452 (
        .din(new_Jinkela_wire_16065),
        .dout(new_Jinkela_wire_16066)
    );

    bfr new_Jinkela_buffer_9984 (
        .din(new_Jinkela_wire_12129),
        .dout(new_Jinkela_wire_12130)
    );

    bfr new_Jinkela_buffer_3073 (
        .din(new_Jinkela_wire_4154),
        .dout(new_Jinkela_wire_4155)
    );

    bfr new_Jinkela_buffer_13511 (
        .din(new_Jinkela_wire_16148),
        .dout(new_Jinkela_wire_16149)
    );

    bfr new_Jinkela_buffer_3109 (
        .din(new_Jinkela_wire_4198),
        .dout(new_Jinkela_wire_4199)
    );

    bfr new_Jinkela_buffer_10077 (
        .din(new_Jinkela_wire_12226),
        .dout(new_Jinkela_wire_12227)
    );

    bfr new_Jinkela_buffer_13453 (
        .din(new_Jinkela_wire_16066),
        .dout(new_Jinkela_wire_16067)
    );

    bfr new_Jinkela_buffer_9985 (
        .din(new_Jinkela_wire_12130),
        .dout(new_Jinkela_wire_12131)
    );

    bfr new_Jinkela_buffer_3074 (
        .din(new_Jinkela_wire_4155),
        .dout(new_Jinkela_wire_4156)
    );

    bfr new_Jinkela_buffer_13675 (
        .din(_1540_),
        .dout(new_Jinkela_wire_16333)
    );

    bfr new_Jinkela_buffer_3167 (
        .din(new_Jinkela_wire_4270),
        .dout(new_Jinkela_wire_4271)
    );

    bfr new_Jinkela_buffer_10035 (
        .din(new_Jinkela_wire_12180),
        .dout(new_Jinkela_wire_12181)
    );

    bfr new_Jinkela_buffer_13454 (
        .din(new_Jinkela_wire_16067),
        .dout(new_Jinkela_wire_16068)
    );

    bfr new_Jinkela_buffer_9986 (
        .din(new_Jinkela_wire_12131),
        .dout(new_Jinkela_wire_12132)
    );

    spl2 new_Jinkela_splitter_390 (
        .a(new_Jinkela_wire_4156),
        .b(new_Jinkela_wire_4157),
        .c(new_Jinkela_wire_4158)
    );

    bfr new_Jinkela_buffer_13512 (
        .din(new_Jinkela_wire_16149),
        .dout(new_Jinkela_wire_16150)
    );

    bfr new_Jinkela_buffer_13455 (
        .din(new_Jinkela_wire_16068),
        .dout(new_Jinkela_wire_16069)
    );

    spl2 new_Jinkela_splitter_404 (
        .a(_1831_),
        .b(new_Jinkela_wire_4294),
        .c(new_Jinkela_wire_4295)
    );

    bfr new_Jinkela_buffer_9987 (
        .din(new_Jinkela_wire_12132),
        .dout(new_Jinkela_wire_12133)
    );

    bfr new_Jinkela_buffer_3110 (
        .din(new_Jinkela_wire_4199),
        .dout(new_Jinkela_wire_4200)
    );

    bfr new_Jinkela_buffer_13559 (
        .din(new_Jinkela_wire_16210),
        .dout(new_Jinkela_wire_16211)
    );

    bfr new_Jinkela_buffer_3111 (
        .din(new_Jinkela_wire_4200),
        .dout(new_Jinkela_wire_4201)
    );

    bfr new_Jinkela_buffer_10036 (
        .din(new_Jinkela_wire_12181),
        .dout(new_Jinkela_wire_12182)
    );

    bfr new_Jinkela_buffer_13456 (
        .din(new_Jinkela_wire_16069),
        .dout(new_Jinkela_wire_16070)
    );

    bfr new_Jinkela_buffer_9988 (
        .din(new_Jinkela_wire_12133),
        .dout(new_Jinkela_wire_12134)
    );

    bfr new_Jinkela_buffer_3168 (
        .din(new_Jinkela_wire_4271),
        .dout(new_Jinkela_wire_4272)
    );

    bfr new_Jinkela_buffer_13513 (
        .din(new_Jinkela_wire_16150),
        .dout(new_Jinkela_wire_16151)
    );

    bfr new_Jinkela_buffer_3112 (
        .din(new_Jinkela_wire_4201),
        .dout(new_Jinkela_wire_4202)
    );

    bfr new_Jinkela_buffer_10078 (
        .din(new_Jinkela_wire_12227),
        .dout(new_Jinkela_wire_12228)
    );

    bfr new_Jinkela_buffer_13457 (
        .din(new_Jinkela_wire_16070),
        .dout(new_Jinkela_wire_16071)
    );

    bfr new_Jinkela_buffer_9989 (
        .din(new_Jinkela_wire_12134),
        .dout(new_Jinkela_wire_12135)
    );

    bfr new_Jinkela_buffer_3179 (
        .din(new_Jinkela_wire_4288),
        .dout(new_Jinkela_wire_4289)
    );

    bfr new_Jinkela_buffer_13674 (
        .din(_0469_),
        .dout(new_Jinkela_wire_16332)
    );

    bfr new_Jinkela_buffer_3113 (
        .din(new_Jinkela_wire_4202),
        .dout(new_Jinkela_wire_4203)
    );

    bfr new_Jinkela_buffer_10037 (
        .din(new_Jinkela_wire_12182),
        .dout(new_Jinkela_wire_12183)
    );

    bfr new_Jinkela_buffer_13458 (
        .din(new_Jinkela_wire_16071),
        .dout(new_Jinkela_wire_16072)
    );

    bfr new_Jinkela_buffer_9990 (
        .din(new_Jinkela_wire_12135),
        .dout(new_Jinkela_wire_12136)
    );

    bfr new_Jinkela_buffer_3169 (
        .din(new_Jinkela_wire_4272),
        .dout(new_Jinkela_wire_4273)
    );

    bfr new_Jinkela_buffer_13514 (
        .din(new_Jinkela_wire_16151),
        .dout(new_Jinkela_wire_16152)
    );

    bfr new_Jinkela_buffer_3114 (
        .din(new_Jinkela_wire_4203),
        .dout(new_Jinkela_wire_4204)
    );

    bfr new_Jinkela_buffer_10178 (
        .din(new_Jinkela_wire_12333),
        .dout(new_Jinkela_wire_12334)
    );

    bfr new_Jinkela_buffer_13459 (
        .din(new_Jinkela_wire_16072),
        .dout(new_Jinkela_wire_16073)
    );

    bfr new_Jinkela_buffer_9991 (
        .din(new_Jinkela_wire_12136),
        .dout(new_Jinkela_wire_12137)
    );

    bfr new_Jinkela_buffer_3184 (
        .din(_0141_),
        .dout(new_Jinkela_wire_4296)
    );

    bfr new_Jinkela_buffer_13562 (
        .din(new_Jinkela_wire_16217),
        .dout(new_Jinkela_wire_16218)
    );

    bfr new_Jinkela_buffer_3115 (
        .din(new_Jinkela_wire_4204),
        .dout(new_Jinkela_wire_4205)
    );

    bfr new_Jinkela_buffer_10038 (
        .din(new_Jinkela_wire_12183),
        .dout(new_Jinkela_wire_12184)
    );

    bfr new_Jinkela_buffer_13460 (
        .din(new_Jinkela_wire_16073),
        .dout(new_Jinkela_wire_16074)
    );

    bfr new_Jinkela_buffer_9992 (
        .din(new_Jinkela_wire_12137),
        .dout(new_Jinkela_wire_12138)
    );

    bfr new_Jinkela_buffer_3170 (
        .din(new_Jinkela_wire_4273),
        .dout(new_Jinkela_wire_4274)
    );

    bfr new_Jinkela_buffer_13515 (
        .din(new_Jinkela_wire_16152),
        .dout(new_Jinkela_wire_16153)
    );

    bfr new_Jinkela_buffer_3116 (
        .din(new_Jinkela_wire_4205),
        .dout(new_Jinkela_wire_4206)
    );

    bfr new_Jinkela_buffer_10079 (
        .din(new_Jinkela_wire_12228),
        .dout(new_Jinkela_wire_12229)
    );

    bfr new_Jinkela_buffer_13461 (
        .din(new_Jinkela_wire_16074),
        .dout(new_Jinkela_wire_16075)
    );

    bfr new_Jinkela_buffer_9993 (
        .din(new_Jinkela_wire_12138),
        .dout(new_Jinkela_wire_12139)
    );

    bfr new_Jinkela_buffer_3180 (
        .din(new_Jinkela_wire_4289),
        .dout(new_Jinkela_wire_4290)
    );

    bfr new_Jinkela_buffer_13676 (
        .din(_1823_),
        .dout(new_Jinkela_wire_16334)
    );

    bfr new_Jinkela_buffer_3117 (
        .din(new_Jinkela_wire_4206),
        .dout(new_Jinkela_wire_4207)
    );

    bfr new_Jinkela_buffer_10039 (
        .din(new_Jinkela_wire_12184),
        .dout(new_Jinkela_wire_12185)
    );

    bfr new_Jinkela_buffer_13462 (
        .din(new_Jinkela_wire_16075),
        .dout(new_Jinkela_wire_16076)
    );

    bfr new_Jinkela_buffer_9994 (
        .din(new_Jinkela_wire_12139),
        .dout(new_Jinkela_wire_12140)
    );

    bfr new_Jinkela_buffer_3171 (
        .din(new_Jinkela_wire_4274),
        .dout(new_Jinkela_wire_4275)
    );

    bfr new_Jinkela_buffer_13516 (
        .din(new_Jinkela_wire_16153),
        .dout(new_Jinkela_wire_16154)
    );

    bfr new_Jinkela_buffer_3118 (
        .din(new_Jinkela_wire_4207),
        .dout(new_Jinkela_wire_4208)
    );

    bfr new_Jinkela_buffer_13463 (
        .din(new_Jinkela_wire_16076),
        .dout(new_Jinkela_wire_16077)
    );

    bfr new_Jinkela_buffer_9995 (
        .din(new_Jinkela_wire_12140),
        .dout(new_Jinkela_wire_12141)
    );

    spl2 new_Jinkela_splitter_405 (
        .a(_1084_),
        .b(new_Jinkela_wire_4298),
        .c(new_Jinkela_wire_4299)
    );

    bfr new_Jinkela_buffer_13563 (
        .din(new_Jinkela_wire_16218),
        .dout(new_Jinkela_wire_16219)
    );

    spl2 new_Jinkela_splitter_929 (
        .a(_1656_),
        .b(new_Jinkela_wire_12341),
        .c(new_Jinkela_wire_12342)
    );

    bfr new_Jinkela_buffer_3119 (
        .din(new_Jinkela_wire_4208),
        .dout(new_Jinkela_wire_4209)
    );

    bfr new_Jinkela_buffer_10040 (
        .din(new_Jinkela_wire_12185),
        .dout(new_Jinkela_wire_12186)
    );

    bfr new_Jinkela_buffer_13464 (
        .din(new_Jinkela_wire_16077),
        .dout(new_Jinkela_wire_16078)
    );

    bfr new_Jinkela_buffer_9996 (
        .din(new_Jinkela_wire_12141),
        .dout(new_Jinkela_wire_12142)
    );

    bfr new_Jinkela_buffer_3172 (
        .din(new_Jinkela_wire_4275),
        .dout(new_Jinkela_wire_4276)
    );

    bfr new_Jinkela_buffer_13517 (
        .din(new_Jinkela_wire_16154),
        .dout(new_Jinkela_wire_16155)
    );

    bfr new_Jinkela_buffer_3120 (
        .din(new_Jinkela_wire_4209),
        .dout(new_Jinkela_wire_4210)
    );

    bfr new_Jinkela_buffer_10080 (
        .din(new_Jinkela_wire_12229),
        .dout(new_Jinkela_wire_12230)
    );

    bfr new_Jinkela_buffer_13465 (
        .din(new_Jinkela_wire_16078),
        .dout(new_Jinkela_wire_16079)
    );

    bfr new_Jinkela_buffer_9997 (
        .din(new_Jinkela_wire_12142),
        .dout(new_Jinkela_wire_12143)
    );

    bfr new_Jinkela_buffer_13708 (
        .din(_1726_),
        .dout(new_Jinkela_wire_16368)
    );

    bfr new_Jinkela_buffer_3185 (
        .din(_0799_),
        .dout(new_Jinkela_wire_4297)
    );

    bfr new_Jinkela_buffer_3121 (
        .din(new_Jinkela_wire_4210),
        .dout(new_Jinkela_wire_4211)
    );

    bfr new_Jinkela_buffer_10041 (
        .din(new_Jinkela_wire_12186),
        .dout(new_Jinkela_wire_12187)
    );

    bfr new_Jinkela_buffer_13466 (
        .din(new_Jinkela_wire_16079),
        .dout(new_Jinkela_wire_16080)
    );

    bfr new_Jinkela_buffer_9998 (
        .din(new_Jinkela_wire_12143),
        .dout(new_Jinkela_wire_12144)
    );

    bfr new_Jinkela_buffer_3173 (
        .din(new_Jinkela_wire_4276),
        .dout(new_Jinkela_wire_4277)
    );

    bfr new_Jinkela_buffer_13518 (
        .din(new_Jinkela_wire_16155),
        .dout(new_Jinkela_wire_16156)
    );

    bfr new_Jinkela_buffer_3122 (
        .din(new_Jinkela_wire_4211),
        .dout(new_Jinkela_wire_4212)
    );

    bfr new_Jinkela_buffer_10179 (
        .din(new_Jinkela_wire_12334),
        .dout(new_Jinkela_wire_12335)
    );

    bfr new_Jinkela_buffer_13467 (
        .din(new_Jinkela_wire_16080),
        .dout(new_Jinkela_wire_16081)
    );

    bfr new_Jinkela_buffer_9999 (
        .din(new_Jinkela_wire_12144),
        .dout(new_Jinkela_wire_12145)
    );

    spl2 new_Jinkela_splitter_407 (
        .a(_0521_),
        .b(new_Jinkela_wire_4303),
        .c(new_Jinkela_wire_4304)
    );

    bfr new_Jinkela_buffer_13564 (
        .din(new_Jinkela_wire_16219),
        .dout(new_Jinkela_wire_16220)
    );

    bfr new_Jinkela_buffer_3123 (
        .din(new_Jinkela_wire_4212),
        .dout(new_Jinkela_wire_4213)
    );

    bfr new_Jinkela_buffer_10042 (
        .din(new_Jinkela_wire_12187),
        .dout(new_Jinkela_wire_12188)
    );

    bfr new_Jinkela_buffer_13468 (
        .din(new_Jinkela_wire_16081),
        .dout(new_Jinkela_wire_16082)
    );

    bfr new_Jinkela_buffer_10000 (
        .din(new_Jinkela_wire_12145),
        .dout(new_Jinkela_wire_12146)
    );

    bfr new_Jinkela_buffer_3174 (
        .din(new_Jinkela_wire_4277),
        .dout(new_Jinkela_wire_4278)
    );

    bfr new_Jinkela_buffer_13519 (
        .din(new_Jinkela_wire_16156),
        .dout(new_Jinkela_wire_16157)
    );

    bfr new_Jinkela_buffer_3124 (
        .din(new_Jinkela_wire_4213),
        .dout(new_Jinkela_wire_4214)
    );

    bfr new_Jinkela_buffer_10081 (
        .din(new_Jinkela_wire_12230),
        .dout(new_Jinkela_wire_12231)
    );

    bfr new_Jinkela_buffer_13469 (
        .din(new_Jinkela_wire_16082),
        .dout(new_Jinkela_wire_16083)
    );

    bfr new_Jinkela_buffer_10001 (
        .din(new_Jinkela_wire_12146),
        .dout(new_Jinkela_wire_12147)
    );

    bfr new_Jinkela_buffer_13709 (
        .din(_1667_),
        .dout(new_Jinkela_wire_16369)
    );

    bfr new_Jinkela_buffer_3125 (
        .din(new_Jinkela_wire_4214),
        .dout(new_Jinkela_wire_4215)
    );

    bfr new_Jinkela_buffer_10043 (
        .din(new_Jinkela_wire_12188),
        .dout(new_Jinkela_wire_12189)
    );

    bfr new_Jinkela_buffer_13470 (
        .din(new_Jinkela_wire_16083),
        .dout(new_Jinkela_wire_16084)
    );

    bfr new_Jinkela_buffer_10002 (
        .din(new_Jinkela_wire_12147),
        .dout(new_Jinkela_wire_12148)
    );

    bfr new_Jinkela_buffer_3175 (
        .din(new_Jinkela_wire_4278),
        .dout(new_Jinkela_wire_4279)
    );

    bfr new_Jinkela_buffer_13520 (
        .din(new_Jinkela_wire_16157),
        .dout(new_Jinkela_wire_16158)
    );

    bfr new_Jinkela_buffer_3126 (
        .din(new_Jinkela_wire_4215),
        .dout(new_Jinkela_wire_4216)
    );

    spl2 new_Jinkela_splitter_931 (
        .a(_1269_),
        .b(new_Jinkela_wire_12520),
        .c(new_Jinkela_wire_12521)
    );

    bfr new_Jinkela_buffer_13471 (
        .din(new_Jinkela_wire_16084),
        .dout(new_Jinkela_wire_16085)
    );

    bfr new_Jinkela_buffer_10003 (
        .din(new_Jinkela_wire_12148),
        .dout(new_Jinkela_wire_12149)
    );

    bfr new_Jinkela_buffer_3187 (
        .din(new_Jinkela_wire_4304),
        .dout(new_Jinkela_wire_4305)
    );

    bfr new_Jinkela_buffer_13565 (
        .din(new_Jinkela_wire_16220),
        .dout(new_Jinkela_wire_16221)
    );

    bfr new_Jinkela_buffer_3186 (
        .din(new_Jinkela_wire_4299),
        .dout(new_Jinkela_wire_4300)
    );

    spl2 new_Jinkela_splitter_930 (
        .a(new_net_0),
        .b(new_Jinkela_wire_12343),
        .c(new_Jinkela_wire_12344)
    );

    bfr new_Jinkela_buffer_3127 (
        .din(new_Jinkela_wire_4216),
        .dout(new_Jinkela_wire_4217)
    );

    bfr new_Jinkela_buffer_10044 (
        .din(new_Jinkela_wire_12189),
        .dout(new_Jinkela_wire_12190)
    );

    bfr new_Jinkela_buffer_13472 (
        .din(new_Jinkela_wire_16085),
        .dout(new_Jinkela_wire_16086)
    );

    bfr new_Jinkela_buffer_10004 (
        .din(new_Jinkela_wire_12149),
        .dout(new_Jinkela_wire_12150)
    );

    bfr new_Jinkela_buffer_3176 (
        .din(new_Jinkela_wire_4279),
        .dout(new_Jinkela_wire_4280)
    );

    bfr new_Jinkela_buffer_13521 (
        .din(new_Jinkela_wire_16158),
        .dout(new_Jinkela_wire_16159)
    );

    bfr new_Jinkela_buffer_16866 (
        .din(new_Jinkela_wire_20112),
        .dout(new_Jinkela_wire_20113)
    );

    bfr new_Jinkela_buffer_10082 (
        .din(new_Jinkela_wire_12231),
        .dout(new_Jinkela_wire_12232)
    );

    and_bb _2245_ (
        .a(new_Jinkela_wire_11),
        .b(new_Jinkela_wire_554),
        .c(_1282_)
    );

    bfr new_Jinkela_buffer_10005 (
        .din(new_Jinkela_wire_12150),
        .dout(new_Jinkela_wire_12151)
    );

    bfr new_Jinkela_buffer_16970 (
        .din(new_Jinkela_wire_20228),
        .dout(new_Jinkela_wire_20229)
    );

    and_bi _2246_ (
        .a(new_Jinkela_wire_851),
        .b(new_Jinkela_wire_13324),
        .c(_1283_)
    );

    bfr new_Jinkela_buffer_16867 (
        .din(new_Jinkela_wire_20113),
        .dout(new_Jinkela_wire_20114)
    );

    bfr new_Jinkela_buffer_10045 (
        .din(new_Jinkela_wire_12190),
        .dout(new_Jinkela_wire_12191)
    );

    and_bb _2247_ (
        .a(new_Jinkela_wire_284),
        .b(new_Jinkela_wire_449),
        .c(_1284_)
    );

    bfr new_Jinkela_buffer_10006 (
        .din(new_Jinkela_wire_12151),
        .dout(new_Jinkela_wire_12152)
    );

    bfr new_Jinkela_buffer_16918 (
        .din(new_Jinkela_wire_20170),
        .dout(new_Jinkela_wire_20171)
    );

    and_bi _2248_ (
        .a(new_Jinkela_wire_20282),
        .b(new_Jinkela_wire_8026),
        .c(_1285_)
    );

    bfr new_Jinkela_buffer_16868 (
        .din(new_Jinkela_wire_20114),
        .dout(new_Jinkela_wire_20115)
    );

    bfr new_Jinkela_buffer_10180 (
        .din(new_Jinkela_wire_12335),
        .dout(new_Jinkela_wire_12336)
    );

    and_bb _2249_ (
        .a(new_Jinkela_wire_68),
        .b(new_Jinkela_wire_243),
        .c(_1286_)
    );

    bfr new_Jinkela_buffer_10007 (
        .din(new_Jinkela_wire_12152),
        .dout(new_Jinkela_wire_12153)
    );

    and_bi _2250_ (
        .a(new_Jinkela_wire_16007),
        .b(new_Jinkela_wire_17672),
        .c(_1287_)
    );

    bfr new_Jinkela_buffer_16869 (
        .din(new_Jinkela_wire_20115),
        .dout(new_Jinkela_wire_20116)
    );

    bfr new_Jinkela_buffer_10046 (
        .din(new_Jinkela_wire_12191),
        .dout(new_Jinkela_wire_12192)
    );

    and_bb _2251_ (
        .a(new_Jinkela_wire_480),
        .b(new_Jinkela_wire_294),
        .c(_1288_)
    );

    bfr new_Jinkela_buffer_10008 (
        .din(new_Jinkela_wire_12153),
        .dout(new_Jinkela_wire_12154)
    );

    bfr new_Jinkela_buffer_16919 (
        .din(new_Jinkela_wire_20171),
        .dout(new_Jinkela_wire_20172)
    );

    and_bi _2252_ (
        .a(new_Jinkela_wire_13977),
        .b(new_Jinkela_wire_5148),
        .c(_1289_)
    );

    bfr new_Jinkela_buffer_16870 (
        .din(new_Jinkela_wire_20116),
        .dout(new_Jinkela_wire_20117)
    );

    bfr new_Jinkela_buffer_10083 (
        .din(new_Jinkela_wire_12232),
        .dout(new_Jinkela_wire_12233)
    );

    and_bb _2253_ (
        .a(new_Jinkela_wire_359),
        .b(new_Jinkela_wire_58),
        .c(_1290_)
    );

    bfr new_Jinkela_buffer_10009 (
        .din(new_Jinkela_wire_12154),
        .dout(new_Jinkela_wire_12155)
    );

    bfr new_Jinkela_buffer_16971 (
        .din(new_Jinkela_wire_20229),
        .dout(new_Jinkela_wire_20230)
    );

    and_bi _2254_ (
        .a(new_Jinkela_wire_18803),
        .b(new_Jinkela_wire_717),
        .c(_1291_)
    );

    bfr new_Jinkela_buffer_16871 (
        .din(new_Jinkela_wire_20117),
        .dout(new_Jinkela_wire_20118)
    );

    bfr new_Jinkela_buffer_10047 (
        .din(new_Jinkela_wire_12192),
        .dout(new_Jinkela_wire_12193)
    );

    and_bb _2255_ (
        .a(new_Jinkela_wire_690),
        .b(new_Jinkela_wire_647),
        .c(_1292_)
    );

    bfr new_Jinkela_buffer_10010 (
        .din(new_Jinkela_wire_12155),
        .dout(new_Jinkela_wire_12156)
    );

    bfr new_Jinkela_buffer_16920 (
        .din(new_Jinkela_wire_20172),
        .dout(new_Jinkela_wire_20173)
    );

    and_bi _2256_ (
        .a(new_Jinkela_wire_4290),
        .b(new_Jinkela_wire_7293),
        .c(_1293_)
    );

    bfr new_Jinkela_buffer_16872 (
        .din(new_Jinkela_wire_20118),
        .dout(new_Jinkela_wire_20119)
    );

    bfr new_Jinkela_buffer_10181 (
        .din(new_Jinkela_wire_12344),
        .dout(new_Jinkela_wire_12345)
    );

    and_bb _2257_ (
        .a(new_Jinkela_wire_621),
        .b(new_Jinkela_wire_493),
        .c(_1294_)
    );

    bfr new_Jinkela_buffer_10011 (
        .din(new_Jinkela_wire_12156),
        .dout(new_Jinkela_wire_12157)
    );

    spl2 new_Jinkela_splitter_1484 (
        .a(new_Jinkela_wire_20272),
        .b(new_Jinkela_wire_20273),
        .c(new_Jinkela_wire_20274)
    );

    and_bi _2258_ (
        .a(new_Jinkela_wire_6416),
        .b(new_Jinkela_wire_3362),
        .c(_1295_)
    );

    bfr new_Jinkela_buffer_16873 (
        .din(new_Jinkela_wire_20119),
        .dout(new_Jinkela_wire_20120)
    );

    bfr new_Jinkela_buffer_10048 (
        .din(new_Jinkela_wire_12193),
        .dout(new_Jinkela_wire_12194)
    );

    and_bb _2259_ (
        .a(new_Jinkela_wire_550),
        .b(new_Jinkela_wire_38),
        .c(_1296_)
    );

    bfr new_Jinkela_buffer_10012 (
        .din(new_Jinkela_wire_12157),
        .dout(new_Jinkela_wire_12158)
    );

    bfr new_Jinkela_buffer_16921 (
        .din(new_Jinkela_wire_20173),
        .dout(new_Jinkela_wire_20174)
    );

    or_ii _2260_ (
        .a(new_Jinkela_wire_376),
        .b(new_Jinkela_wire_317),
        .c(_1297_)
    );

    bfr new_Jinkela_buffer_16874 (
        .din(new_Jinkela_wire_20120),
        .dout(new_Jinkela_wire_20121)
    );

    bfr new_Jinkela_buffer_10084 (
        .din(new_Jinkela_wire_12233),
        .dout(new_Jinkela_wire_12234)
    );

    and_bi _2261_ (
        .a(new_Jinkela_wire_1804),
        .b(new_Jinkela_wire_18523),
        .c(_1298_)
    );

    bfr new_Jinkela_buffer_10013 (
        .din(new_Jinkela_wire_12158),
        .dout(new_Jinkela_wire_12159)
    );

    bfr new_Jinkela_buffer_16972 (
        .din(new_Jinkela_wire_20230),
        .dout(new_Jinkela_wire_20231)
    );

    and_bb _2262_ (
        .a(new_Jinkela_wire_391),
        .b(new_Jinkela_wire_241),
        .c(_1299_)
    );

    bfr new_Jinkela_buffer_16875 (
        .din(new_Jinkela_wire_20121),
        .dout(new_Jinkela_wire_20122)
    );

    bfr new_Jinkela_buffer_10049 (
        .din(new_Jinkela_wire_12194),
        .dout(new_Jinkela_wire_12195)
    );

    and_bi _2263_ (
        .a(new_Jinkela_wire_6517),
        .b(new_Jinkela_wire_1621),
        .c(_1300_)
    );

    bfr new_Jinkela_buffer_10014 (
        .din(new_Jinkela_wire_12159),
        .dout(new_Jinkela_wire_12160)
    );

    bfr new_Jinkela_buffer_16922 (
        .din(new_Jinkela_wire_20174),
        .dout(new_Jinkela_wire_20175)
    );

    and_ii _2264_ (
        .a(new_Jinkela_wire_21198),
        .b(new_Jinkela_wire_20041),
        .c(_1301_)
    );

    bfr new_Jinkela_buffer_16876 (
        .din(new_Jinkela_wire_20122),
        .dout(new_Jinkela_wire_20123)
    );

    or_bb _2265_ (
        .a(new_Jinkela_wire_14192),
        .b(new_Jinkela_wire_15751),
        .c(_1302_)
    );

    bfr new_Jinkela_buffer_10015 (
        .din(new_Jinkela_wire_12160),
        .dout(new_Jinkela_wire_12161)
    );

    bfr new_Jinkela_buffer_17002 (
        .din(new_Jinkela_wire_20278),
        .dout(new_Jinkela_wire_20279)
    );

    or_ii _2266_ (
        .a(new_Jinkela_wire_14193),
        .b(new_Jinkela_wire_15750),
        .c(_1303_)
    );

    spl2 new_Jinkela_splitter_932 (
        .a(_0355_),
        .b(new_Jinkela_wire_12522),
        .c(new_Jinkela_wire_12523)
    );

    spl2 new_Jinkela_splitter_1488 (
        .a(_0203_),
        .b(new_Jinkela_wire_20285),
        .c(new_Jinkela_wire_20286)
    );

    bfr new_Jinkela_buffer_16877 (
        .din(new_Jinkela_wire_20123),
        .dout(new_Jinkela_wire_20124)
    );

    bfr new_Jinkela_buffer_10050 (
        .din(new_Jinkela_wire_12195),
        .dout(new_Jinkela_wire_12196)
    );

    or_ii _2267_ (
        .a(new_Jinkela_wire_3879),
        .b(new_Jinkela_wire_13141),
        .c(_1304_)
    );

    bfr new_Jinkela_buffer_10016 (
        .din(new_Jinkela_wire_12161),
        .dout(new_Jinkela_wire_12162)
    );

    bfr new_Jinkela_buffer_16923 (
        .din(new_Jinkela_wire_20175),
        .dout(new_Jinkela_wire_20176)
    );

    and_ii _2268_ (
        .a(new_Jinkela_wire_9556),
        .b(new_Jinkela_wire_14297),
        .c(_1305_)
    );

    bfr new_Jinkela_buffer_16878 (
        .din(new_Jinkela_wire_20124),
        .dout(new_Jinkela_wire_20125)
    );

    bfr new_Jinkela_buffer_10085 (
        .din(new_Jinkela_wire_12234),
        .dout(new_Jinkela_wire_12235)
    );

    and_bb _2269_ (
        .a(new_Jinkela_wire_9557),
        .b(new_Jinkela_wire_14298),
        .c(_1306_)
    );

    bfr new_Jinkela_buffer_10017 (
        .din(new_Jinkela_wire_12162),
        .dout(new_Jinkela_wire_12163)
    );

    bfr new_Jinkela_buffer_16973 (
        .din(new_Jinkela_wire_20231),
        .dout(new_Jinkela_wire_20232)
    );

    or_bb _2270_ (
        .a(new_Jinkela_wire_10394),
        .b(new_Jinkela_wire_4726),
        .c(_1307_)
    );

    bfr new_Jinkela_buffer_16879 (
        .din(new_Jinkela_wire_20125),
        .dout(new_Jinkela_wire_20126)
    );

    bfr new_Jinkela_buffer_10051 (
        .din(new_Jinkela_wire_12196),
        .dout(new_Jinkela_wire_12197)
    );

    or_bb _2271_ (
        .a(new_Jinkela_wire_9177),
        .b(new_Jinkela_wire_19930),
        .c(_1308_)
    );

    bfr new_Jinkela_buffer_10018 (
        .din(new_Jinkela_wire_12163),
        .dout(new_Jinkela_wire_12164)
    );

    bfr new_Jinkela_buffer_16924 (
        .din(new_Jinkela_wire_20176),
        .dout(new_Jinkela_wire_20177)
    );

    or_ii _2272_ (
        .a(new_Jinkela_wire_9178),
        .b(new_Jinkela_wire_19931),
        .c(_1309_)
    );

    bfr new_Jinkela_buffer_16880 (
        .din(new_Jinkela_wire_20126),
        .dout(new_Jinkela_wire_20127)
    );

    bfr new_Jinkela_buffer_10356 (
        .din(_0546_),
        .dout(new_Jinkela_wire_12524)
    );

    or_ii _2273_ (
        .a(new_Jinkela_wire_17030),
        .b(new_Jinkela_wire_5422),
        .c(_1310_)
    );

    bfr new_Jinkela_buffer_10019 (
        .din(new_Jinkela_wire_12164),
        .dout(new_Jinkela_wire_12165)
    );

    and_ii _2274_ (
        .a(new_Jinkela_wire_16010),
        .b(new_Jinkela_wire_17106),
        .c(_1311_)
    );

    spl2 new_Jinkela_splitter_1487 (
        .a(_0324_),
        .b(new_Jinkela_wire_20283),
        .c(new_Jinkela_wire_20284)
    );

    bfr new_Jinkela_buffer_16881 (
        .din(new_Jinkela_wire_20127),
        .dout(new_Jinkela_wire_20128)
    );

    bfr new_Jinkela_buffer_10052 (
        .din(new_Jinkela_wire_12197),
        .dout(new_Jinkela_wire_12198)
    );

    and_bb _2275_ (
        .a(new_Jinkela_wire_16011),
        .b(new_Jinkela_wire_17107),
        .c(_1312_)
    );

    bfr new_Jinkela_buffer_10020 (
        .din(new_Jinkela_wire_12165),
        .dout(new_Jinkela_wire_12166)
    );

    bfr new_Jinkela_buffer_16925 (
        .din(new_Jinkela_wire_20177),
        .dout(new_Jinkela_wire_20178)
    );

    or_bb _2276_ (
        .a(new_Jinkela_wire_11829),
        .b(new_Jinkela_wire_7316),
        .c(_1313_)
    );

    bfr new_Jinkela_buffer_16882 (
        .din(new_Jinkela_wire_20128),
        .dout(new_Jinkela_wire_20129)
    );

    bfr new_Jinkela_buffer_10086 (
        .din(new_Jinkela_wire_12235),
        .dout(new_Jinkela_wire_12236)
    );

    or_bb _2277_ (
        .a(new_Jinkela_wire_17534),
        .b(new_Jinkela_wire_14036),
        .c(_1314_)
    );

    bfr new_Jinkela_buffer_10021 (
        .din(new_Jinkela_wire_12166),
        .dout(new_Jinkela_wire_12167)
    );

    bfr new_Jinkela_buffer_16974 (
        .din(new_Jinkela_wire_20232),
        .dout(new_Jinkela_wire_20233)
    );

    or_ii _2278_ (
        .a(new_Jinkela_wire_17535),
        .b(new_Jinkela_wire_14037),
        .c(_1315_)
    );

    bfr new_Jinkela_buffer_16883 (
        .din(new_Jinkela_wire_20129),
        .dout(new_Jinkela_wire_20130)
    );

    bfr new_Jinkela_buffer_10053 (
        .din(new_Jinkela_wire_12198),
        .dout(new_Jinkela_wire_12199)
    );

    or_ii _2279_ (
        .a(new_Jinkela_wire_5998),
        .b(new_Jinkela_wire_11434),
        .c(_1316_)
    );

    bfr new_Jinkela_buffer_10022 (
        .din(new_Jinkela_wire_12167),
        .dout(new_Jinkela_wire_12168)
    );

    bfr new_Jinkela_buffer_16926 (
        .din(new_Jinkela_wire_20178),
        .dout(new_Jinkela_wire_20179)
    );

    and_ii _2280_ (
        .a(new_Jinkela_wire_15779),
        .b(new_Jinkela_wire_20319),
        .c(_1317_)
    );

    spl2 new_Jinkela_splitter_1472 (
        .a(new_Jinkela_wire_20130),
        .b(new_Jinkela_wire_20131),
        .c(new_Jinkela_wire_20132)
    );

    bfr new_Jinkela_buffer_10182 (
        .din(new_Jinkela_wire_12345),
        .dout(new_Jinkela_wire_12346)
    );

    and_bb _2281_ (
        .a(new_Jinkela_wire_15780),
        .b(new_Jinkela_wire_20320),
        .c(_1318_)
    );

    bfr new_Jinkela_buffer_10023 (
        .din(new_Jinkela_wire_12168),
        .dout(new_Jinkela_wire_12169)
    );

    bfr new_Jinkela_buffer_16927 (
        .din(new_Jinkela_wire_20179),
        .dout(new_Jinkela_wire_20180)
    );

    or_bb _2282_ (
        .a(new_Jinkela_wire_4663),
        .b(new_Jinkela_wire_12715),
        .c(_1319_)
    );

    spl2 new_Jinkela_splitter_1489 (
        .a(_1703_),
        .b(new_Jinkela_wire_20287),
        .c(new_Jinkela_wire_20288)
    );

    bfr new_Jinkela_buffer_10054 (
        .din(new_Jinkela_wire_12199),
        .dout(new_Jinkela_wire_12200)
    );

    or_bb _2283_ (
        .a(new_Jinkela_wire_4072),
        .b(new_Jinkela_wire_14690),
        .c(_1320_)
    );

    bfr new_Jinkela_buffer_10024 (
        .din(new_Jinkela_wire_12169),
        .dout(new_Jinkela_wire_12170)
    );

    bfr new_Jinkela_buffer_16975 (
        .din(new_Jinkela_wire_20233),
        .dout(new_Jinkela_wire_20234)
    );

    or_ii _2284_ (
        .a(new_Jinkela_wire_4073),
        .b(new_Jinkela_wire_14691),
        .c(_1321_)
    );

    bfr new_Jinkela_buffer_16928 (
        .din(new_Jinkela_wire_20180),
        .dout(new_Jinkela_wire_20181)
    );

    bfr new_Jinkela_buffer_10087 (
        .din(new_Jinkela_wire_12236),
        .dout(new_Jinkela_wire_12237)
    );

    or_ii _2285_ (
        .a(new_Jinkela_wire_3441),
        .b(new_Jinkela_wire_18381),
        .c(_1322_)
    );

    bfr new_Jinkela_buffer_17003 (
        .din(new_Jinkela_wire_20279),
        .dout(new_Jinkela_wire_20280)
    );

    bfr new_Jinkela_buffer_10055 (
        .din(new_Jinkela_wire_12200),
        .dout(new_Jinkela_wire_12201)
    );

    and_ii _2286_ (
        .a(new_Jinkela_wire_3195),
        .b(new_Jinkela_wire_10612),
        .c(_1323_)
    );

    bfr new_Jinkela_buffer_13473 (
        .din(new_Jinkela_wire_16086),
        .dout(new_Jinkela_wire_16087)
    );

    bfr new_Jinkela_buffer_13677 (
        .din(new_Jinkela_wire_16334),
        .dout(new_Jinkela_wire_16335)
    );

    bfr new_Jinkela_buffer_13474 (
        .din(new_Jinkela_wire_16087),
        .dout(new_Jinkela_wire_16088)
    );

    bfr new_Jinkela_buffer_13522 (
        .din(new_Jinkela_wire_16159),
        .dout(new_Jinkela_wire_16160)
    );

    bfr new_Jinkela_buffer_13475 (
        .din(new_Jinkela_wire_16088),
        .dout(new_Jinkela_wire_16089)
    );

    bfr new_Jinkela_buffer_13566 (
        .din(new_Jinkela_wire_16221),
        .dout(new_Jinkela_wire_16222)
    );

    bfr new_Jinkela_buffer_13476 (
        .din(new_Jinkela_wire_16089),
        .dout(new_Jinkela_wire_16090)
    );

    bfr new_Jinkela_buffer_13523 (
        .din(new_Jinkela_wire_16160),
        .dout(new_Jinkela_wire_16161)
    );

    bfr new_Jinkela_buffer_13477 (
        .din(new_Jinkela_wire_16090),
        .dout(new_Jinkela_wire_16091)
    );

    bfr new_Jinkela_buffer_13710 (
        .din(_1142_),
        .dout(new_Jinkela_wire_16370)
    );

    bfr new_Jinkela_buffer_13478 (
        .din(new_Jinkela_wire_16091),
        .dout(new_Jinkela_wire_16092)
    );

    bfr new_Jinkela_buffer_13524 (
        .din(new_Jinkela_wire_16161),
        .dout(new_Jinkela_wire_16162)
    );

    bfr new_Jinkela_buffer_13479 (
        .din(new_Jinkela_wire_16092),
        .dout(new_Jinkela_wire_16093)
    );

    bfr new_Jinkela_buffer_13567 (
        .din(new_Jinkela_wire_16222),
        .dout(new_Jinkela_wire_16223)
    );

    bfr new_Jinkela_buffer_13480 (
        .din(new_Jinkela_wire_16093),
        .dout(new_Jinkela_wire_16094)
    );

    bfr new_Jinkela_buffer_13525 (
        .din(new_Jinkela_wire_16162),
        .dout(new_Jinkela_wire_16163)
    );

    bfr new_Jinkela_buffer_13481 (
        .din(new_Jinkela_wire_16094),
        .dout(new_Jinkela_wire_16095)
    );

    bfr new_Jinkela_buffer_13678 (
        .din(new_Jinkela_wire_16335),
        .dout(new_Jinkela_wire_16336)
    );

    bfr new_Jinkela_buffer_13482 (
        .din(new_Jinkela_wire_16095),
        .dout(new_Jinkela_wire_16096)
    );

    bfr new_Jinkela_buffer_13526 (
        .din(new_Jinkela_wire_16163),
        .dout(new_Jinkela_wire_16164)
    );

    bfr new_Jinkela_buffer_13483 (
        .din(new_Jinkela_wire_16096),
        .dout(new_Jinkela_wire_16097)
    );

    bfr new_Jinkela_buffer_13568 (
        .din(new_Jinkela_wire_16223),
        .dout(new_Jinkela_wire_16224)
    );

    bfr new_Jinkela_buffer_13484 (
        .din(new_Jinkela_wire_16097),
        .dout(new_Jinkela_wire_16098)
    );

    bfr new_Jinkela_buffer_13527 (
        .din(new_Jinkela_wire_16164),
        .dout(new_Jinkela_wire_16165)
    );

    bfr new_Jinkela_buffer_13485 (
        .din(new_Jinkela_wire_16098),
        .dout(new_Jinkela_wire_16099)
    );

    bfr new_Jinkela_buffer_13718 (
        .din(_0544_),
        .dout(new_Jinkela_wire_16380)
    );

    spl2 new_Jinkela_splitter_1156 (
        .a(new_Jinkela_wire_16099),
        .b(new_Jinkela_wire_16100),
        .c(new_Jinkela_wire_16101)
    );

    bfr new_Jinkela_buffer_13569 (
        .din(new_Jinkela_wire_16224),
        .dout(new_Jinkela_wire_16225)
    );

    bfr new_Jinkela_buffer_13528 (
        .din(new_Jinkela_wire_16165),
        .dout(new_Jinkela_wire_16166)
    );

    bfr new_Jinkela_buffer_13529 (
        .din(new_Jinkela_wire_16166),
        .dout(new_Jinkela_wire_16167)
    );

    bfr new_Jinkela_buffer_13679 (
        .din(new_Jinkela_wire_16336),
        .dout(new_Jinkela_wire_16337)
    );

    bfr new_Jinkela_buffer_13530 (
        .din(new_Jinkela_wire_16167),
        .dout(new_Jinkela_wire_16168)
    );

    bfr new_Jinkela_buffer_13570 (
        .din(new_Jinkela_wire_16225),
        .dout(new_Jinkela_wire_16226)
    );

    bfr new_Jinkela_buffer_13531 (
        .din(new_Jinkela_wire_16168),
        .dout(new_Jinkela_wire_16169)
    );

    spl2 new_Jinkela_splitter_1181 (
        .a(_0411_),
        .b(new_Jinkela_wire_16436),
        .c(new_Jinkela_wire_16437)
    );

    bfr new_Jinkela_buffer_13532 (
        .din(new_Jinkela_wire_16169),
        .dout(new_Jinkela_wire_16170)
    );

    bfr new_Jinkela_buffer_13571 (
        .din(new_Jinkela_wire_16226),
        .dout(new_Jinkela_wire_16227)
    );

    bfr new_Jinkela_buffer_13533 (
        .din(new_Jinkela_wire_16170),
        .dout(new_Jinkela_wire_16171)
    );

    bfr new_Jinkela_buffer_13680 (
        .din(new_Jinkela_wire_16337),
        .dout(new_Jinkela_wire_16338)
    );

    bfr new_Jinkela_buffer_13534 (
        .din(new_Jinkela_wire_16171),
        .dout(new_Jinkela_wire_16172)
    );

    bfr new_Jinkela_buffer_13572 (
        .din(new_Jinkela_wire_16227),
        .dout(new_Jinkela_wire_16228)
    );

    bfr new_Jinkela_buffer_13535 (
        .din(new_Jinkela_wire_16172),
        .dout(new_Jinkela_wire_16173)
    );

    bfr new_Jinkela_buffer_3128 (
        .din(new_Jinkela_wire_4217),
        .dout(new_Jinkela_wire_4218)
    );

    bfr new_Jinkela_buffer_6540 (
        .din(new_Jinkela_wire_8239),
        .dout(new_Jinkela_wire_8240)
    );

    spl2 new_Jinkela_splitter_408 (
        .a(_0814_),
        .b(new_Jinkela_wire_4321),
        .c(new_Jinkela_wire_4322)
    );

    bfr new_Jinkela_buffer_6737 (
        .din(new_Jinkela_wire_8462),
        .dout(new_Jinkela_wire_8463)
    );

    bfr new_Jinkela_buffer_3207 (
        .din(_0670_),
        .dout(new_Jinkela_wire_4327)
    );

    bfr new_Jinkela_buffer_3129 (
        .din(new_Jinkela_wire_4218),
        .dout(new_Jinkela_wire_4219)
    );

    bfr new_Jinkela_buffer_6541 (
        .din(new_Jinkela_wire_8240),
        .dout(new_Jinkela_wire_8241)
    );

    spl2 new_Jinkela_splitter_401 (
        .a(new_Jinkela_wire_4280),
        .b(new_Jinkela_wire_4281),
        .c(new_Jinkela_wire_4282)
    );

    bfr new_Jinkela_buffer_6589 (
        .din(new_Jinkela_wire_8308),
        .dout(new_Jinkela_wire_8309)
    );

    bfr new_Jinkela_buffer_3130 (
        .din(new_Jinkela_wire_4219),
        .dout(new_Jinkela_wire_4220)
    );

    bfr new_Jinkela_buffer_6542 (
        .din(new_Jinkela_wire_8241),
        .dout(new_Jinkela_wire_8242)
    );

    bfr new_Jinkela_buffer_6643 (
        .din(new_Jinkela_wire_8366),
        .dout(new_Jinkela_wire_8367)
    );

    bfr new_Jinkela_buffer_3131 (
        .din(new_Jinkela_wire_4220),
        .dout(new_Jinkela_wire_4221)
    );

    bfr new_Jinkela_buffer_6543 (
        .din(new_Jinkela_wire_8242),
        .dout(new_Jinkela_wire_8243)
    );

    bfr new_Jinkela_buffer_3203 (
        .din(new_Jinkela_wire_4322),
        .dout(new_Jinkela_wire_4323)
    );

    bfr new_Jinkela_buffer_6590 (
        .din(new_Jinkela_wire_8309),
        .dout(new_Jinkela_wire_8310)
    );

    spl2 new_Jinkela_splitter_406 (
        .a(new_Jinkela_wire_4300),
        .b(new_Jinkela_wire_4301),
        .c(new_Jinkela_wire_4302)
    );

    bfr new_Jinkela_buffer_3132 (
        .din(new_Jinkela_wire_4221),
        .dout(new_Jinkela_wire_4222)
    );

    bfr new_Jinkela_buffer_6544 (
        .din(new_Jinkela_wire_8243),
        .dout(new_Jinkela_wire_8244)
    );

    bfr new_Jinkela_buffer_3188 (
        .din(new_Jinkela_wire_4305),
        .dout(new_Jinkela_wire_4306)
    );

    spl2 new_Jinkela_splitter_718 (
        .a(_0146_),
        .b(new_Jinkela_wire_8584),
        .c(new_Jinkela_wire_8585)
    );

    bfr new_Jinkela_buffer_3133 (
        .din(new_Jinkela_wire_4222),
        .dout(new_Jinkela_wire_4223)
    );

    bfr new_Jinkela_buffer_6545 (
        .din(new_Jinkela_wire_8244),
        .dout(new_Jinkela_wire_8245)
    );

    bfr new_Jinkela_buffer_6591 (
        .din(new_Jinkela_wire_8310),
        .dout(new_Jinkela_wire_8311)
    );

    bfr new_Jinkela_buffer_3134 (
        .din(new_Jinkela_wire_4223),
        .dout(new_Jinkela_wire_4224)
    );

    bfr new_Jinkela_buffer_6546 (
        .din(new_Jinkela_wire_8245),
        .dout(new_Jinkela_wire_8246)
    );

    bfr new_Jinkela_buffer_6644 (
        .din(new_Jinkela_wire_8367),
        .dout(new_Jinkela_wire_8368)
    );

    spl2 new_Jinkela_splitter_409 (
        .a(_1414_),
        .b(new_Jinkela_wire_4328),
        .c(new_Jinkela_wire_4329)
    );

    bfr new_Jinkela_buffer_3135 (
        .din(new_Jinkela_wire_4224),
        .dout(new_Jinkela_wire_4225)
    );

    bfr new_Jinkela_buffer_6547 (
        .din(new_Jinkela_wire_8246),
        .dout(new_Jinkela_wire_8247)
    );

    bfr new_Jinkela_buffer_3189 (
        .din(new_Jinkela_wire_4306),
        .dout(new_Jinkela_wire_4307)
    );

    bfr new_Jinkela_buffer_6592 (
        .din(new_Jinkela_wire_8311),
        .dout(new_Jinkela_wire_8312)
    );

    bfr new_Jinkela_buffer_3136 (
        .din(new_Jinkela_wire_4225),
        .dout(new_Jinkela_wire_4226)
    );

    bfr new_Jinkela_buffer_6548 (
        .din(new_Jinkela_wire_8247),
        .dout(new_Jinkela_wire_8248)
    );

    bfr new_Jinkela_buffer_3208 (
        .din(new_net_3950),
        .dout(new_Jinkela_wire_4330)
    );

    bfr new_Jinkela_buffer_6738 (
        .din(new_Jinkela_wire_8463),
        .dout(new_Jinkela_wire_8464)
    );

    bfr new_Jinkela_buffer_3137 (
        .din(new_Jinkela_wire_4226),
        .dout(new_Jinkela_wire_4227)
    );

    bfr new_Jinkela_buffer_6549 (
        .din(new_Jinkela_wire_8248),
        .dout(new_Jinkela_wire_8249)
    );

    bfr new_Jinkela_buffer_3190 (
        .din(new_Jinkela_wire_4307),
        .dout(new_Jinkela_wire_4308)
    );

    bfr new_Jinkela_buffer_6593 (
        .din(new_Jinkela_wire_8312),
        .dout(new_Jinkela_wire_8313)
    );

    bfr new_Jinkela_buffer_3138 (
        .din(new_Jinkela_wire_4227),
        .dout(new_Jinkela_wire_4228)
    );

    bfr new_Jinkela_buffer_6550 (
        .din(new_Jinkela_wire_8249),
        .dout(new_Jinkela_wire_8250)
    );

    bfr new_Jinkela_buffer_3204 (
        .din(new_Jinkela_wire_4323),
        .dout(new_Jinkela_wire_4324)
    );

    bfr new_Jinkela_buffer_6645 (
        .din(new_Jinkela_wire_8368),
        .dout(new_Jinkela_wire_8369)
    );

    bfr new_Jinkela_buffer_3139 (
        .din(new_Jinkela_wire_4228),
        .dout(new_Jinkela_wire_4229)
    );

    bfr new_Jinkela_buffer_6551 (
        .din(new_Jinkela_wire_8250),
        .dout(new_Jinkela_wire_8251)
    );

    bfr new_Jinkela_buffer_3191 (
        .din(new_Jinkela_wire_4308),
        .dout(new_Jinkela_wire_4309)
    );

    bfr new_Jinkela_buffer_6594 (
        .din(new_Jinkela_wire_8313),
        .dout(new_Jinkela_wire_8314)
    );

    bfr new_Jinkela_buffer_3140 (
        .din(new_Jinkela_wire_4229),
        .dout(new_Jinkela_wire_4230)
    );

    bfr new_Jinkela_buffer_6552 (
        .din(new_Jinkela_wire_8251),
        .dout(new_Jinkela_wire_8252)
    );

    bfr new_Jinkela_buffer_3209 (
        .din(new_Jinkela_wire_4330),
        .dout(new_Jinkela_wire_4331)
    );

    bfr new_Jinkela_buffer_6752 (
        .din(_0964_),
        .dout(new_Jinkela_wire_8484)
    );

    bfr new_Jinkela_buffer_3141 (
        .din(new_Jinkela_wire_4230),
        .dout(new_Jinkela_wire_4231)
    );

    bfr new_Jinkela_buffer_6553 (
        .din(new_Jinkela_wire_8252),
        .dout(new_Jinkela_wire_8253)
    );

    bfr new_Jinkela_buffer_3192 (
        .din(new_Jinkela_wire_4309),
        .dout(new_Jinkela_wire_4310)
    );

    bfr new_Jinkela_buffer_6595 (
        .din(new_Jinkela_wire_8314),
        .dout(new_Jinkela_wire_8315)
    );

    bfr new_Jinkela_buffer_3142 (
        .din(new_Jinkela_wire_4231),
        .dout(new_Jinkela_wire_4232)
    );

    bfr new_Jinkela_buffer_6554 (
        .din(new_Jinkela_wire_8253),
        .dout(new_Jinkela_wire_8254)
    );

    bfr new_Jinkela_buffer_3205 (
        .din(new_Jinkela_wire_4324),
        .dout(new_Jinkela_wire_4325)
    );

    bfr new_Jinkela_buffer_6646 (
        .din(new_Jinkela_wire_8369),
        .dout(new_Jinkela_wire_8370)
    );

    bfr new_Jinkela_buffer_3143 (
        .din(new_Jinkela_wire_4232),
        .dout(new_Jinkela_wire_4233)
    );

    bfr new_Jinkela_buffer_6555 (
        .din(new_Jinkela_wire_8254),
        .dout(new_Jinkela_wire_8255)
    );

    bfr new_Jinkela_buffer_3193 (
        .din(new_Jinkela_wire_4310),
        .dout(new_Jinkela_wire_4311)
    );

    bfr new_Jinkela_buffer_6596 (
        .din(new_Jinkela_wire_8315),
        .dout(new_Jinkela_wire_8316)
    );

    bfr new_Jinkela_buffer_3144 (
        .din(new_Jinkela_wire_4233),
        .dout(new_Jinkela_wire_4234)
    );

    bfr new_Jinkela_buffer_6556 (
        .din(new_Jinkela_wire_8255),
        .dout(new_Jinkela_wire_8256)
    );

    bfr new_Jinkela_buffer_6739 (
        .din(new_Jinkela_wire_8464),
        .dout(new_Jinkela_wire_8465)
    );

    bfr new_Jinkela_buffer_3340 (
        .din(_0571_),
        .dout(new_Jinkela_wire_4462)
    );

    bfr new_Jinkela_buffer_3145 (
        .din(new_Jinkela_wire_4234),
        .dout(new_Jinkela_wire_4235)
    );

    bfr new_Jinkela_buffer_6557 (
        .din(new_Jinkela_wire_8256),
        .dout(new_Jinkela_wire_8257)
    );

    bfr new_Jinkela_buffer_3194 (
        .din(new_Jinkela_wire_4311),
        .dout(new_Jinkela_wire_4312)
    );

    bfr new_Jinkela_buffer_6597 (
        .din(new_Jinkela_wire_8316),
        .dout(new_Jinkela_wire_8317)
    );

    spl2 new_Jinkela_splitter_394 (
        .a(new_Jinkela_wire_4235),
        .b(new_Jinkela_wire_4236),
        .c(new_Jinkela_wire_4237)
    );

    bfr new_Jinkela_buffer_6558 (
        .din(new_Jinkela_wire_8257),
        .dout(new_Jinkela_wire_8258)
    );

    bfr new_Jinkela_buffer_3195 (
        .din(new_Jinkela_wire_4312),
        .dout(new_Jinkela_wire_4313)
    );

    bfr new_Jinkela_buffer_6647 (
        .din(new_Jinkela_wire_8370),
        .dout(new_Jinkela_wire_8371)
    );

    bfr new_Jinkela_buffer_3206 (
        .din(new_Jinkela_wire_4325),
        .dout(new_Jinkela_wire_4326)
    );

    bfr new_Jinkela_buffer_6559 (
        .din(new_Jinkela_wire_8258),
        .dout(new_Jinkela_wire_8259)
    );

    bfr new_Jinkela_buffer_6598 (
        .din(new_Jinkela_wire_8317),
        .dout(new_Jinkela_wire_8318)
    );

    bfr new_Jinkela_buffer_3341 (
        .din(_1082_),
        .dout(new_Jinkela_wire_4463)
    );

    bfr new_Jinkela_buffer_3196 (
        .din(new_Jinkela_wire_4313),
        .dout(new_Jinkela_wire_4314)
    );

    bfr new_Jinkela_buffer_6560 (
        .din(new_Jinkela_wire_8259),
        .dout(new_Jinkela_wire_8260)
    );

    spl2 new_Jinkela_splitter_411 (
        .a(_0917_),
        .b(new_Jinkela_wire_4473),
        .c(new_Jinkela_wire_4474)
    );

    bfr new_Jinkela_buffer_3210 (
        .din(new_Jinkela_wire_4331),
        .dout(new_Jinkela_wire_4332)
    );

    spl2 new_Jinkela_splitter_934 (
        .a(_1154_),
        .b(new_Jinkela_wire_12615),
        .c(new_Jinkela_wire_12616)
    );

    bfr new_Jinkela_buffer_6561 (
        .din(new_Jinkela_wire_8260),
        .dout(new_Jinkela_wire_8261)
    );

    bfr new_Jinkela_buffer_16929 (
        .din(new_Jinkela_wire_20181),
        .dout(new_Jinkela_wire_20182)
    );

    bfr new_Jinkela_buffer_10056 (
        .din(new_Jinkela_wire_12201),
        .dout(new_Jinkela_wire_12202)
    );

    bfr new_Jinkela_buffer_6599 (
        .din(new_Jinkela_wire_8318),
        .dout(new_Jinkela_wire_8319)
    );

    bfr new_Jinkela_buffer_16976 (
        .din(new_Jinkela_wire_20234),
        .dout(new_Jinkela_wire_20235)
    );

    bfr new_Jinkela_buffer_10088 (
        .din(new_Jinkela_wire_12237),
        .dout(new_Jinkela_wire_12238)
    );

    bfr new_Jinkela_buffer_6562 (
        .din(new_Jinkela_wire_8261),
        .dout(new_Jinkela_wire_8262)
    );

    bfr new_Jinkela_buffer_16930 (
        .din(new_Jinkela_wire_20182),
        .dout(new_Jinkela_wire_20183)
    );

    bfr new_Jinkela_buffer_10057 (
        .din(new_Jinkela_wire_12202),
        .dout(new_Jinkela_wire_12203)
    );

    bfr new_Jinkela_buffer_6648 (
        .din(new_Jinkela_wire_8371),
        .dout(new_Jinkela_wire_8372)
    );

    bfr new_Jinkela_buffer_17034 (
        .din(_1504_),
        .dout(new_Jinkela_wire_20321)
    );

    bfr new_Jinkela_buffer_10183 (
        .din(new_Jinkela_wire_12346),
        .dout(new_Jinkela_wire_12347)
    );

    bfr new_Jinkela_buffer_6563 (
        .din(new_Jinkela_wire_8262),
        .dout(new_Jinkela_wire_8263)
    );

    bfr new_Jinkela_buffer_16931 (
        .din(new_Jinkela_wire_20183),
        .dout(new_Jinkela_wire_20184)
    );

    bfr new_Jinkela_buffer_10058 (
        .din(new_Jinkela_wire_12203),
        .dout(new_Jinkela_wire_12204)
    );

    bfr new_Jinkela_buffer_6600 (
        .din(new_Jinkela_wire_8319),
        .dout(new_Jinkela_wire_8320)
    );

    bfr new_Jinkela_buffer_16977 (
        .din(new_Jinkela_wire_20235),
        .dout(new_Jinkela_wire_20236)
    );

    bfr new_Jinkela_buffer_10089 (
        .din(new_Jinkela_wire_12238),
        .dout(new_Jinkela_wire_12239)
    );

    bfr new_Jinkela_buffer_6564 (
        .din(new_Jinkela_wire_8263),
        .dout(new_Jinkela_wire_8264)
    );

    bfr new_Jinkela_buffer_16932 (
        .din(new_Jinkela_wire_20184),
        .dout(new_Jinkela_wire_20185)
    );

    bfr new_Jinkela_buffer_10059 (
        .din(new_Jinkela_wire_12204),
        .dout(new_Jinkela_wire_12205)
    );

    bfr new_Jinkela_buffer_6740 (
        .din(new_Jinkela_wire_8465),
        .dout(new_Jinkela_wire_8466)
    );

    bfr new_Jinkela_buffer_17004 (
        .din(new_Jinkela_wire_20280),
        .dout(new_Jinkela_wire_20281)
    );

    bfr new_Jinkela_buffer_16933 (
        .din(new_Jinkela_wire_20185),
        .dout(new_Jinkela_wire_20186)
    );

    bfr new_Jinkela_buffer_6565 (
        .din(new_Jinkela_wire_8264),
        .dout(new_Jinkela_wire_8265)
    );

    bfr new_Jinkela_buffer_10357 (
        .din(_1454_),
        .dout(new_Jinkela_wire_12525)
    );

    bfr new_Jinkela_buffer_10060 (
        .din(new_Jinkela_wire_12205),
        .dout(new_Jinkela_wire_12206)
    );

    bfr new_Jinkela_buffer_6601 (
        .din(new_Jinkela_wire_8320),
        .dout(new_Jinkela_wire_8321)
    );

    bfr new_Jinkela_buffer_16978 (
        .din(new_Jinkela_wire_20236),
        .dout(new_Jinkela_wire_20237)
    );

    bfr new_Jinkela_buffer_10090 (
        .din(new_Jinkela_wire_12239),
        .dout(new_Jinkela_wire_12240)
    );

    bfr new_Jinkela_buffer_6566 (
        .din(new_Jinkela_wire_8265),
        .dout(new_Jinkela_wire_8266)
    );

    bfr new_Jinkela_buffer_16934 (
        .din(new_Jinkela_wire_20186),
        .dout(new_Jinkela_wire_20187)
    );

    bfr new_Jinkela_buffer_10061 (
        .din(new_Jinkela_wire_12206),
        .dout(new_Jinkela_wire_12207)
    );

    bfr new_Jinkela_buffer_6649 (
        .din(new_Jinkela_wire_8372),
        .dout(new_Jinkela_wire_8373)
    );

    bfr new_Jinkela_buffer_17006 (
        .din(_1835_),
        .dout(new_Jinkela_wire_20289)
    );

    bfr new_Jinkela_buffer_10184 (
        .din(new_Jinkela_wire_12347),
        .dout(new_Jinkela_wire_12348)
    );

    bfr new_Jinkela_buffer_6567 (
        .din(new_Jinkela_wire_8266),
        .dout(new_Jinkela_wire_8267)
    );

    bfr new_Jinkela_buffer_16935 (
        .din(new_Jinkela_wire_20187),
        .dout(new_Jinkela_wire_20188)
    );

    bfr new_Jinkela_buffer_10062 (
        .din(new_Jinkela_wire_12207),
        .dout(new_Jinkela_wire_12208)
    );

    bfr new_Jinkela_buffer_6602 (
        .din(new_Jinkela_wire_8321),
        .dout(new_Jinkela_wire_8322)
    );

    bfr new_Jinkela_buffer_16979 (
        .din(new_Jinkela_wire_20237),
        .dout(new_Jinkela_wire_20238)
    );

    bfr new_Jinkela_buffer_10091 (
        .din(new_Jinkela_wire_12240),
        .dout(new_Jinkela_wire_12241)
    );

    bfr new_Jinkela_buffer_6568 (
        .din(new_Jinkela_wire_8267),
        .dout(new_Jinkela_wire_8268)
    );

    bfr new_Jinkela_buffer_16936 (
        .din(new_Jinkela_wire_20188),
        .dout(new_Jinkela_wire_20189)
    );

    bfr new_Jinkela_buffer_10063 (
        .din(new_Jinkela_wire_12208),
        .dout(new_Jinkela_wire_12209)
    );

    bfr new_Jinkela_buffer_6753 (
        .din(new_Jinkela_wire_8484),
        .dout(new_Jinkela_wire_8485)
    );

    bfr new_Jinkela_buffer_17005 (
        .din(new_Jinkela_wire_20281),
        .dout(new_Jinkela_wire_20282)
    );

    bfr new_Jinkela_buffer_16937 (
        .din(new_Jinkela_wire_20189),
        .dout(new_Jinkela_wire_20190)
    );

    bfr new_Jinkela_buffer_6569 (
        .din(new_Jinkela_wire_8268),
        .dout(new_Jinkela_wire_8269)
    );

    bfr new_Jinkela_buffer_10449 (
        .din(_0356_),
        .dout(new_Jinkela_wire_12621)
    );

    bfr new_Jinkela_buffer_10064 (
        .din(new_Jinkela_wire_12209),
        .dout(new_Jinkela_wire_12210)
    );

    bfr new_Jinkela_buffer_6603 (
        .din(new_Jinkela_wire_8322),
        .dout(new_Jinkela_wire_8323)
    );

    bfr new_Jinkela_buffer_16980 (
        .din(new_Jinkela_wire_20238),
        .dout(new_Jinkela_wire_20239)
    );

    bfr new_Jinkela_buffer_10092 (
        .din(new_Jinkela_wire_12241),
        .dout(new_Jinkela_wire_12242)
    );

    bfr new_Jinkela_buffer_6570 (
        .din(new_Jinkela_wire_8269),
        .dout(new_Jinkela_wire_8270)
    );

    bfr new_Jinkela_buffer_16938 (
        .din(new_Jinkela_wire_20190),
        .dout(new_Jinkela_wire_20191)
    );

    bfr new_Jinkela_buffer_10065 (
        .din(new_Jinkela_wire_12210),
        .dout(new_Jinkela_wire_12211)
    );

    bfr new_Jinkela_buffer_6650 (
        .din(new_Jinkela_wire_8373),
        .dout(new_Jinkela_wire_8374)
    );

    spl2 new_Jinkela_splitter_1492 (
        .a(_0487_),
        .b(new_Jinkela_wire_20322),
        .c(new_Jinkela_wire_20323)
    );

    bfr new_Jinkela_buffer_17010 (
        .din(_1292_),
        .dout(new_Jinkela_wire_20295)
    );

    bfr new_Jinkela_buffer_10185 (
        .din(new_Jinkela_wire_12348),
        .dout(new_Jinkela_wire_12349)
    );

    bfr new_Jinkela_buffer_6571 (
        .din(new_Jinkela_wire_8270),
        .dout(new_Jinkela_wire_8271)
    );

    bfr new_Jinkela_buffer_16939 (
        .din(new_Jinkela_wire_20191),
        .dout(new_Jinkela_wire_20192)
    );

    bfr new_Jinkela_buffer_10066 (
        .din(new_Jinkela_wire_12211),
        .dout(new_Jinkela_wire_12212)
    );

    bfr new_Jinkela_buffer_6604 (
        .din(new_Jinkela_wire_8323),
        .dout(new_Jinkela_wire_8324)
    );

    bfr new_Jinkela_buffer_16981 (
        .din(new_Jinkela_wire_20239),
        .dout(new_Jinkela_wire_20240)
    );

    bfr new_Jinkela_buffer_10093 (
        .din(new_Jinkela_wire_12242),
        .dout(new_Jinkela_wire_12243)
    );

    bfr new_Jinkela_buffer_6572 (
        .din(new_Jinkela_wire_8271),
        .dout(new_Jinkela_wire_8272)
    );

    bfr new_Jinkela_buffer_16940 (
        .din(new_Jinkela_wire_20192),
        .dout(new_Jinkela_wire_20193)
    );

    bfr new_Jinkela_buffer_10067 (
        .din(new_Jinkela_wire_12212),
        .dout(new_Jinkela_wire_12213)
    );

    bfr new_Jinkela_buffer_6741 (
        .din(new_Jinkela_wire_8466),
        .dout(new_Jinkela_wire_8467)
    );

    bfr new_Jinkela_buffer_17007 (
        .din(new_Jinkela_wire_20289),
        .dout(new_Jinkela_wire_20290)
    );

    bfr new_Jinkela_buffer_10358 (
        .din(new_Jinkela_wire_12525),
        .dout(new_Jinkela_wire_12526)
    );

    bfr new_Jinkela_buffer_6573 (
        .din(new_Jinkela_wire_8272),
        .dout(new_Jinkela_wire_8273)
    );

    bfr new_Jinkela_buffer_16941 (
        .din(new_Jinkela_wire_20193),
        .dout(new_Jinkela_wire_20194)
    );

    bfr new_Jinkela_buffer_10068 (
        .din(new_Jinkela_wire_12213),
        .dout(new_Jinkela_wire_12214)
    );

    bfr new_Jinkela_buffer_6605 (
        .din(new_Jinkela_wire_8324),
        .dout(new_Jinkela_wire_8325)
    );

    bfr new_Jinkela_buffer_16982 (
        .din(new_Jinkela_wire_20240),
        .dout(new_Jinkela_wire_20241)
    );

    bfr new_Jinkela_buffer_10094 (
        .din(new_Jinkela_wire_12243),
        .dout(new_Jinkela_wire_12244)
    );

    spl2 new_Jinkela_splitter_699 (
        .a(new_Jinkela_wire_8273),
        .b(new_Jinkela_wire_8274),
        .c(new_Jinkela_wire_8275)
    );

    bfr new_Jinkela_buffer_16942 (
        .din(new_Jinkela_wire_20194),
        .dout(new_Jinkela_wire_20195)
    );

    bfr new_Jinkela_buffer_10069 (
        .din(new_Jinkela_wire_12214),
        .dout(new_Jinkela_wire_12215)
    );

    bfr new_Jinkela_buffer_6606 (
        .din(new_Jinkela_wire_8325),
        .dout(new_Jinkela_wire_8326)
    );

    bfr new_Jinkela_buffer_17008 (
        .din(new_Jinkela_wire_20290),
        .dout(new_Jinkela_wire_20291)
    );

    bfr new_Jinkela_buffer_10186 (
        .din(new_Jinkela_wire_12349),
        .dout(new_Jinkela_wire_12350)
    );

    bfr new_Jinkela_buffer_6651 (
        .din(new_Jinkela_wire_8374),
        .dout(new_Jinkela_wire_8375)
    );

    bfr new_Jinkela_buffer_16943 (
        .din(new_Jinkela_wire_20195),
        .dout(new_Jinkela_wire_20196)
    );

    bfr new_Jinkela_buffer_10070 (
        .din(new_Jinkela_wire_12215),
        .dout(new_Jinkela_wire_12216)
    );

    spl2 new_Jinkela_splitter_717 (
        .a(_0454_),
        .b(new_Jinkela_wire_8582),
        .c(new_Jinkela_wire_8583)
    );

    bfr new_Jinkela_buffer_16983 (
        .din(new_Jinkela_wire_20241),
        .dout(new_Jinkela_wire_20242)
    );

    spl2 new_Jinkela_splitter_716 (
        .a(_0665_),
        .b(new_Jinkela_wire_8580),
        .c(new_Jinkela_wire_8581)
    );

    bfr new_Jinkela_buffer_10095 (
        .din(new_Jinkela_wire_12244),
        .dout(new_Jinkela_wire_12245)
    );

    bfr new_Jinkela_buffer_6607 (
        .din(new_Jinkela_wire_8326),
        .dout(new_Jinkela_wire_8327)
    );

    bfr new_Jinkela_buffer_16944 (
        .din(new_Jinkela_wire_20196),
        .dout(new_Jinkela_wire_20197)
    );

    bfr new_Jinkela_buffer_10071 (
        .din(new_Jinkela_wire_12216),
        .dout(new_Jinkela_wire_12217)
    );

    bfr new_Jinkela_buffer_6652 (
        .din(new_Jinkela_wire_8375),
        .dout(new_Jinkela_wire_8376)
    );

    bfr new_Jinkela_buffer_16945 (
        .din(new_Jinkela_wire_20197),
        .dout(new_Jinkela_wire_20198)
    );

    bfr new_Jinkela_buffer_6608 (
        .din(new_Jinkela_wire_8327),
        .dout(new_Jinkela_wire_8328)
    );

    bfr new_Jinkela_buffer_10445 (
        .din(new_Jinkela_wire_12616),
        .dout(new_Jinkela_wire_12617)
    );

    bfr new_Jinkela_buffer_10072 (
        .din(new_Jinkela_wire_12217),
        .dout(new_Jinkela_wire_12218)
    );

    bfr new_Jinkela_buffer_6742 (
        .din(new_Jinkela_wire_8467),
        .dout(new_Jinkela_wire_8468)
    );

    bfr new_Jinkela_buffer_16984 (
        .din(new_Jinkela_wire_20242),
        .dout(new_Jinkela_wire_20243)
    );

    bfr new_Jinkela_buffer_10096 (
        .din(new_Jinkela_wire_12245),
        .dout(new_Jinkela_wire_12246)
    );

    bfr new_Jinkela_buffer_6609 (
        .din(new_Jinkela_wire_8328),
        .dout(new_Jinkela_wire_8329)
    );

    bfr new_Jinkela_buffer_16946 (
        .din(new_Jinkela_wire_20198),
        .dout(new_Jinkela_wire_20199)
    );

    spl2 new_Jinkela_splitter_922 (
        .a(new_Jinkela_wire_12218),
        .b(new_Jinkela_wire_12219),
        .c(new_Jinkela_wire_12220)
    );

    bfr new_Jinkela_buffer_6653 (
        .din(new_Jinkela_wire_8376),
        .dout(new_Jinkela_wire_8377)
    );

    bfr new_Jinkela_buffer_17011 (
        .din(new_Jinkela_wire_20295),
        .dout(new_Jinkela_wire_20296)
    );

    bfr new_Jinkela_buffer_10097 (
        .din(new_Jinkela_wire_12246),
        .dout(new_Jinkela_wire_12247)
    );

    bfr new_Jinkela_buffer_6610 (
        .din(new_Jinkela_wire_8329),
        .dout(new_Jinkela_wire_8330)
    );

    bfr new_Jinkela_buffer_16947 (
        .din(new_Jinkela_wire_20199),
        .dout(new_Jinkela_wire_20200)
    );

    bfr new_Jinkela_buffer_10187 (
        .din(new_Jinkela_wire_12350),
        .dout(new_Jinkela_wire_12351)
    );

    bfr new_Jinkela_buffer_6754 (
        .din(new_Jinkela_wire_8485),
        .dout(new_Jinkela_wire_8486)
    );

    bfr new_Jinkela_buffer_16985 (
        .din(new_Jinkela_wire_20243),
        .dout(new_Jinkela_wire_20244)
    );

    bfr new_Jinkela_buffer_10359 (
        .din(new_Jinkela_wire_12526),
        .dout(new_Jinkela_wire_12527)
    );

    bfr new_Jinkela_buffer_6611 (
        .din(new_Jinkela_wire_8330),
        .dout(new_Jinkela_wire_8331)
    );

    bfr new_Jinkela_buffer_16948 (
        .din(new_Jinkela_wire_20200),
        .dout(new_Jinkela_wire_20201)
    );

    bfr new_Jinkela_buffer_10098 (
        .din(new_Jinkela_wire_12247),
        .dout(new_Jinkela_wire_12248)
    );

    bfr new_Jinkela_buffer_6654 (
        .din(new_Jinkela_wire_8377),
        .dout(new_Jinkela_wire_8378)
    );

    bfr new_Jinkela_buffer_17009 (
        .din(new_Jinkela_wire_20291),
        .dout(new_Jinkela_wire_20292)
    );

    bfr new_Jinkela_buffer_10188 (
        .din(new_Jinkela_wire_12351),
        .dout(new_Jinkela_wire_12352)
    );

    bfr new_Jinkela_buffer_6612 (
        .din(new_Jinkela_wire_8331),
        .dout(new_Jinkela_wire_8332)
    );

    bfr new_Jinkela_buffer_16949 (
        .din(new_Jinkela_wire_20201),
        .dout(new_Jinkela_wire_20202)
    );

    bfr new_Jinkela_buffer_10099 (
        .din(new_Jinkela_wire_12248),
        .dout(new_Jinkela_wire_12249)
    );

    bfr new_Jinkela_buffer_6743 (
        .din(new_Jinkela_wire_8468),
        .dout(new_Jinkela_wire_8469)
    );

    bfr new_Jinkela_buffer_16986 (
        .din(new_Jinkela_wire_20244),
        .dout(new_Jinkela_wire_20245)
    );

    and_bb _2287_ (
        .a(new_Jinkela_wire_3196),
        .b(new_Jinkela_wire_10613),
        .c(_1324_)
    );

    or_bb _2288_ (
        .a(new_Jinkela_wire_4484),
        .b(new_Jinkela_wire_5731),
        .c(_1325_)
    );

    or_bb _2289_ (
        .a(new_Jinkela_wire_17543),
        .b(new_Jinkela_wire_5968),
        .c(_1326_)
    );

    or_ii _2290_ (
        .a(new_Jinkela_wire_17544),
        .b(new_Jinkela_wire_5969),
        .c(_1327_)
    );

    or_ii _2291_ (
        .a(new_Jinkela_wire_20262),
        .b(new_Jinkela_wire_1906),
        .c(_1328_)
    );

    and_ii _2292_ (
        .a(new_Jinkela_wire_3701),
        .b(new_Jinkela_wire_3427),
        .c(_1329_)
    );

    and_bb _2293_ (
        .a(new_Jinkela_wire_3702),
        .b(new_Jinkela_wire_3428),
        .c(_1330_)
    );

    or_bb _2294_ (
        .a(new_Jinkela_wire_5730),
        .b(new_Jinkela_wire_8278),
        .c(_1331_)
    );

    or_bb _2295_ (
        .a(new_Jinkela_wire_17681),
        .b(new_Jinkela_wire_5435),
        .c(_1332_)
    );

    or_ii _2296_ (
        .a(new_Jinkela_wire_17682),
        .b(new_Jinkela_wire_5436),
        .c(_1333_)
    );

    or_ii _2297_ (
        .a(new_Jinkela_wire_11406),
        .b(new_Jinkela_wire_18963),
        .c(_1334_)
    );

    and_ii _2298_ (
        .a(new_Jinkela_wire_19347),
        .b(new_Jinkela_wire_1385),
        .c(_1335_)
    );

    and_bb _2299_ (
        .a(new_Jinkela_wire_19348),
        .b(new_Jinkela_wire_1386),
        .c(_1336_)
    );

    or_bb _2300_ (
        .a(new_Jinkela_wire_2483),
        .b(new_Jinkela_wire_13065),
        .c(_1337_)
    );

    or_bb _2301_ (
        .a(new_Jinkela_wire_21214),
        .b(new_Jinkela_wire_4475),
        .c(_1338_)
    );

    or_ii _2302_ (
        .a(new_Jinkela_wire_21215),
        .b(new_Jinkela_wire_4476),
        .c(_1339_)
    );

    or_ii _2303_ (
        .a(new_Jinkela_wire_18379),
        .b(new_Jinkela_wire_19144),
        .c(_1340_)
    );

    and_ii _2304_ (
        .a(new_Jinkela_wire_15758),
        .b(new_Jinkela_wire_17782),
        .c(_1341_)
    );

    and_bb _2305_ (
        .a(new_Jinkela_wire_15759),
        .b(new_Jinkela_wire_17783),
        .c(_1342_)
    );

    or_bb _2306_ (
        .a(new_Jinkela_wire_20902),
        .b(new_Jinkela_wire_2462),
        .c(_1343_)
    );

    or_bb _2307_ (
        .a(new_Jinkela_wire_20267),
        .b(new_Jinkela_wire_6194),
        .c(_1344_)
    );

    or_ii _2308_ (
        .a(new_Jinkela_wire_20268),
        .b(new_Jinkela_wire_6195),
        .c(_1345_)
    );

    or_ii _2309_ (
        .a(new_Jinkela_wire_21096),
        .b(new_Jinkela_wire_10085),
        .c(_1346_)
    );

    and_ii _2310_ (
        .a(new_Jinkela_wire_6855),
        .b(new_Jinkela_wire_8758),
        .c(_1347_)
    );

    and_bb _2311_ (
        .a(new_Jinkela_wire_6856),
        .b(new_Jinkela_wire_8759),
        .c(_1348_)
    );

    or_bb _2312_ (
        .a(new_Jinkela_wire_10066),
        .b(new_Jinkela_wire_20394),
        .c(_1349_)
    );

    or_bb _2313_ (
        .a(new_Jinkela_wire_16008),
        .b(new_Jinkela_wire_3269),
        .c(_1350_)
    );

    or_ii _2314_ (
        .a(new_Jinkela_wire_16009),
        .b(new_Jinkela_wire_3270),
        .c(_1351_)
    );

    or_ii _2315_ (
        .a(new_Jinkela_wire_8180),
        .b(new_Jinkela_wire_7136),
        .c(_1352_)
    );

    and_ii _2316_ (
        .a(new_Jinkela_wire_18393),
        .b(new_Jinkela_wire_4157),
        .c(_1353_)
    );

    and_bb _2317_ (
        .a(new_Jinkela_wire_18394),
        .b(new_Jinkela_wire_4158),
        .c(_1354_)
    );

    or_bb _2318_ (
        .a(new_Jinkela_wire_2956),
        .b(new_Jinkela_wire_20049),
        .c(_1355_)
    );

    or_bb _2319_ (
        .a(new_Jinkela_wire_16118),
        .b(new_Jinkela_wire_20398),
        .c(_1356_)
    );

    and_bb _2320_ (
        .a(new_Jinkela_wire_16119),
        .b(new_Jinkela_wire_20399),
        .c(_1357_)
    );

    or_bi _2321_ (
        .a(new_Jinkela_wire_1811),
        .b(new_Jinkela_wire_4690),
        .c(_1358_)
    );

    and_ii _2322_ (
        .a(new_Jinkela_wire_17083),
        .b(new_Jinkela_wire_14776),
        .c(_1359_)
    );

    and_bb _2323_ (
        .a(new_Jinkela_wire_17084),
        .b(new_Jinkela_wire_14777),
        .c(_1360_)
    );

    or_bb _2324_ (
        .a(new_Jinkela_wire_16601),
        .b(new_Jinkela_wire_9599),
        .c(new_net_3926)
    );

    and_bb _2325_ (
        .a(new_Jinkela_wire_217),
        .b(new_Jinkela_wire_334),
        .c(_1361_)
    );

    and_bi _2326_ (
        .a(new_Jinkela_wire_4695),
        .b(new_Jinkela_wire_9600),
        .c(_1362_)
    );

    and_bb _2327_ (
        .a(new_Jinkela_wire_96),
        .b(new_Jinkela_wire_587),
        .c(_1363_)
    );

    and_bi _2328_ (
        .a(new_Jinkela_wire_7141),
        .b(new_Jinkela_wire_20050),
        .c(_1364_)
    );

    bfr new_Jinkela_buffer_13711 (
        .din(new_Jinkela_wire_16370),
        .dout(new_Jinkela_wire_16371)
    );

    bfr new_Jinkela_buffer_13536 (
        .din(new_Jinkela_wire_16173),
        .dout(new_Jinkela_wire_16174)
    );

    bfr new_Jinkela_buffer_13573 (
        .din(new_Jinkela_wire_16228),
        .dout(new_Jinkela_wire_16229)
    );

    bfr new_Jinkela_buffer_13537 (
        .din(new_Jinkela_wire_16174),
        .dout(new_Jinkela_wire_16175)
    );

    bfr new_Jinkela_buffer_13681 (
        .din(new_Jinkela_wire_16338),
        .dout(new_Jinkela_wire_16339)
    );

    bfr new_Jinkela_buffer_13538 (
        .din(new_Jinkela_wire_16175),
        .dout(new_Jinkela_wire_16176)
    );

    bfr new_Jinkela_buffer_13574 (
        .din(new_Jinkela_wire_16229),
        .dout(new_Jinkela_wire_16230)
    );

    bfr new_Jinkela_buffer_13539 (
        .din(new_Jinkela_wire_16176),
        .dout(new_Jinkela_wire_16177)
    );

    bfr new_Jinkela_buffer_13776 (
        .din(_0445_),
        .dout(new_Jinkela_wire_16442)
    );

    bfr new_Jinkela_buffer_13540 (
        .din(new_Jinkela_wire_16177),
        .dout(new_Jinkela_wire_16178)
    );

    bfr new_Jinkela_buffer_13575 (
        .din(new_Jinkela_wire_16230),
        .dout(new_Jinkela_wire_16231)
    );

    bfr new_Jinkela_buffer_13541 (
        .din(new_Jinkela_wire_16178),
        .dout(new_Jinkela_wire_16179)
    );

    bfr new_Jinkela_buffer_13682 (
        .din(new_Jinkela_wire_16339),
        .dout(new_Jinkela_wire_16340)
    );

    bfr new_Jinkela_buffer_13542 (
        .din(new_Jinkela_wire_16179),
        .dout(new_Jinkela_wire_16180)
    );

    bfr new_Jinkela_buffer_13576 (
        .din(new_Jinkela_wire_16231),
        .dout(new_Jinkela_wire_16232)
    );

    bfr new_Jinkela_buffer_13543 (
        .din(new_Jinkela_wire_16180),
        .dout(new_Jinkela_wire_16181)
    );

    bfr new_Jinkela_buffer_13712 (
        .din(new_Jinkela_wire_16371),
        .dout(new_Jinkela_wire_16372)
    );

    bfr new_Jinkela_buffer_13544 (
        .din(new_Jinkela_wire_16181),
        .dout(new_Jinkela_wire_16182)
    );

    bfr new_Jinkela_buffer_13577 (
        .din(new_Jinkela_wire_16232),
        .dout(new_Jinkela_wire_16233)
    );

    bfr new_Jinkela_buffer_13545 (
        .din(new_Jinkela_wire_16182),
        .dout(new_Jinkela_wire_16183)
    );

    bfr new_Jinkela_buffer_13683 (
        .din(new_Jinkela_wire_16340),
        .dout(new_Jinkela_wire_16341)
    );

    bfr new_Jinkela_buffer_13546 (
        .din(new_Jinkela_wire_16183),
        .dout(new_Jinkela_wire_16184)
    );

    bfr new_Jinkela_buffer_13578 (
        .din(new_Jinkela_wire_16233),
        .dout(new_Jinkela_wire_16234)
    );

    bfr new_Jinkela_buffer_13547 (
        .din(new_Jinkela_wire_16184),
        .dout(new_Jinkela_wire_16185)
    );

    bfr new_Jinkela_buffer_13719 (
        .din(new_Jinkela_wire_16380),
        .dout(new_Jinkela_wire_16381)
    );

    bfr new_Jinkela_buffer_13548 (
        .din(new_Jinkela_wire_16185),
        .dout(new_Jinkela_wire_16186)
    );

    bfr new_Jinkela_buffer_13579 (
        .din(new_Jinkela_wire_16234),
        .dout(new_Jinkela_wire_16235)
    );

    bfr new_Jinkela_buffer_13549 (
        .din(new_Jinkela_wire_16186),
        .dout(new_Jinkela_wire_16187)
    );

    bfr new_Jinkela_buffer_13684 (
        .din(new_Jinkela_wire_16341),
        .dout(new_Jinkela_wire_16342)
    );

    spl2 new_Jinkela_splitter_1168 (
        .a(new_Jinkela_wire_16187),
        .b(new_Jinkela_wire_16188),
        .c(new_Jinkela_wire_16189)
    );

    bfr new_Jinkela_buffer_13713 (
        .din(new_Jinkela_wire_16372),
        .dout(new_Jinkela_wire_16373)
    );

    bfr new_Jinkela_buffer_13580 (
        .din(new_Jinkela_wire_16235),
        .dout(new_Jinkela_wire_16236)
    );

    bfr new_Jinkela_buffer_13581 (
        .din(new_Jinkela_wire_16236),
        .dout(new_Jinkela_wire_16237)
    );

    bfr new_Jinkela_buffer_13685 (
        .din(new_Jinkela_wire_16342),
        .dout(new_Jinkela_wire_16343)
    );

    bfr new_Jinkela_buffer_13582 (
        .din(new_Jinkela_wire_16237),
        .dout(new_Jinkela_wire_16238)
    );

    bfr new_Jinkela_buffer_13772 (
        .din(new_Jinkela_wire_16437),
        .dout(new_Jinkela_wire_16438)
    );

    bfr new_Jinkela_buffer_13583 (
        .din(new_Jinkela_wire_16238),
        .dout(new_Jinkela_wire_16239)
    );

    bfr new_Jinkela_buffer_13686 (
        .din(new_Jinkela_wire_16343),
        .dout(new_Jinkela_wire_16344)
    );

    bfr new_Jinkela_buffer_13584 (
        .din(new_Jinkela_wire_16239),
        .dout(new_Jinkela_wire_16240)
    );

    bfr new_Jinkela_buffer_13714 (
        .din(new_Jinkela_wire_16373),
        .dout(new_Jinkela_wire_16374)
    );

    bfr new_Jinkela_buffer_13585 (
        .din(new_Jinkela_wire_16240),
        .dout(new_Jinkela_wire_16241)
    );

    bfr new_Jinkela_buffer_13687 (
        .din(new_Jinkela_wire_16344),
        .dout(new_Jinkela_wire_16345)
    );

    bfr new_Jinkela_buffer_9333 (
        .din(new_Jinkela_wire_11362),
        .dout(new_Jinkela_wire_11363)
    );

    bfr new_Jinkela_buffer_12709 (
        .din(new_Jinkela_wire_15230),
        .dout(new_Jinkela_wire_15231)
    );

    bfr new_Jinkela_buffer_9193 (
        .din(new_Jinkela_wire_11212),
        .dout(new_Jinkela_wire_11213)
    );

    bfr new_Jinkela_buffer_12663 (
        .din(new_Jinkela_wire_15178),
        .dout(new_Jinkela_wire_15179)
    );

    bfr new_Jinkela_buffer_9245 (
        .din(new_Jinkela_wire_11268),
        .dout(new_Jinkela_wire_11269)
    );

    bfr new_Jinkela_buffer_12869 (
        .din(new_Jinkela_wire_15390),
        .dout(new_Jinkela_wire_15391)
    );

    bfr new_Jinkela_buffer_9194 (
        .din(new_Jinkela_wire_11213),
        .dout(new_Jinkela_wire_11214)
    );

    bfr new_Jinkela_buffer_12664 (
        .din(new_Jinkela_wire_15179),
        .dout(new_Jinkela_wire_15180)
    );

    spl2 new_Jinkela_splitter_874 (
        .a(_0105_),
        .b(new_Jinkela_wire_11409),
        .c(new_Jinkela_wire_11410)
    );

    bfr new_Jinkela_buffer_9360 (
        .din(new_Jinkela_wire_11417),
        .dout(new_Jinkela_wire_11418)
    );

    bfr new_Jinkela_buffer_12710 (
        .din(new_Jinkela_wire_15231),
        .dout(new_Jinkela_wire_15232)
    );

    bfr new_Jinkela_buffer_9195 (
        .din(new_Jinkela_wire_11214),
        .dout(new_Jinkela_wire_11215)
    );

    bfr new_Jinkela_buffer_12665 (
        .din(new_Jinkela_wire_15180),
        .dout(new_Jinkela_wire_15181)
    );

    bfr new_Jinkela_buffer_9246 (
        .din(new_Jinkela_wire_11269),
        .dout(new_Jinkela_wire_11270)
    );

    bfr new_Jinkela_buffer_12948 (
        .din(new_Jinkela_wire_15471),
        .dout(new_Jinkela_wire_15472)
    );

    bfr new_Jinkela_buffer_9196 (
        .din(new_Jinkela_wire_11215),
        .dout(new_Jinkela_wire_11216)
    );

    bfr new_Jinkela_buffer_12666 (
        .din(new_Jinkela_wire_15181),
        .dout(new_Jinkela_wire_15182)
    );

    bfr new_Jinkela_buffer_9334 (
        .din(new_Jinkela_wire_11363),
        .dout(new_Jinkela_wire_11364)
    );

    bfr new_Jinkela_buffer_12879 (
        .din(new_Jinkela_wire_15400),
        .dout(new_Jinkela_wire_15401)
    );

    bfr new_Jinkela_buffer_12711 (
        .din(new_Jinkela_wire_15232),
        .dout(new_Jinkela_wire_15233)
    );

    bfr new_Jinkela_buffer_9197 (
        .din(new_Jinkela_wire_11216),
        .dout(new_Jinkela_wire_11217)
    );

    bfr new_Jinkela_buffer_12667 (
        .din(new_Jinkela_wire_15182),
        .dout(new_Jinkela_wire_15183)
    );

    bfr new_Jinkela_buffer_9247 (
        .din(new_Jinkela_wire_11270),
        .dout(new_Jinkela_wire_11271)
    );

    bfr new_Jinkela_buffer_12870 (
        .din(new_Jinkela_wire_15391),
        .dout(new_Jinkela_wire_15392)
    );

    bfr new_Jinkela_buffer_9198 (
        .din(new_Jinkela_wire_11217),
        .dout(new_Jinkela_wire_11218)
    );

    bfr new_Jinkela_buffer_12668 (
        .din(new_Jinkela_wire_15183),
        .dout(new_Jinkela_wire_15184)
    );

    bfr new_Jinkela_buffer_12712 (
        .din(new_Jinkela_wire_15233),
        .dout(new_Jinkela_wire_15234)
    );

    bfr new_Jinkela_buffer_9199 (
        .din(new_Jinkela_wire_11218),
        .dout(new_Jinkela_wire_11219)
    );

    bfr new_Jinkela_buffer_12669 (
        .din(new_Jinkela_wire_15184),
        .dout(new_Jinkela_wire_15185)
    );

    bfr new_Jinkela_buffer_9248 (
        .din(new_Jinkela_wire_11271),
        .dout(new_Jinkela_wire_11272)
    );

    bfr new_Jinkela_buffer_9200 (
        .din(new_Jinkela_wire_11219),
        .dout(new_Jinkela_wire_11220)
    );

    bfr new_Jinkela_buffer_12670 (
        .din(new_Jinkela_wire_15185),
        .dout(new_Jinkela_wire_15186)
    );

    bfr new_Jinkela_buffer_9335 (
        .din(new_Jinkela_wire_11364),
        .dout(new_Jinkela_wire_11365)
    );

    bfr new_Jinkela_buffer_12713 (
        .din(new_Jinkela_wire_15234),
        .dout(new_Jinkela_wire_15235)
    );

    bfr new_Jinkela_buffer_9201 (
        .din(new_Jinkela_wire_11220),
        .dout(new_Jinkela_wire_11221)
    );

    bfr new_Jinkela_buffer_12671 (
        .din(new_Jinkela_wire_15186),
        .dout(new_Jinkela_wire_15187)
    );

    bfr new_Jinkela_buffer_9249 (
        .din(new_Jinkela_wire_11272),
        .dout(new_Jinkela_wire_11273)
    );

    bfr new_Jinkela_buffer_12871 (
        .din(new_Jinkela_wire_15392),
        .dout(new_Jinkela_wire_15393)
    );

    bfr new_Jinkela_buffer_9202 (
        .din(new_Jinkela_wire_11221),
        .dout(new_Jinkela_wire_11222)
    );

    bfr new_Jinkela_buffer_12672 (
        .din(new_Jinkela_wire_15187),
        .dout(new_Jinkela_wire_15188)
    );

    bfr new_Jinkela_buffer_9359 (
        .din(_0297_),
        .dout(new_Jinkela_wire_11411)
    );

    bfr new_Jinkela_buffer_12714 (
        .din(new_Jinkela_wire_15235),
        .dout(new_Jinkela_wire_15236)
    );

    bfr new_Jinkela_buffer_9203 (
        .din(new_Jinkela_wire_11222),
        .dout(new_Jinkela_wire_11223)
    );

    bfr new_Jinkela_buffer_12673 (
        .din(new_Jinkela_wire_15188),
        .dout(new_Jinkela_wire_15189)
    );

    bfr new_Jinkela_buffer_9250 (
        .din(new_Jinkela_wire_11273),
        .dout(new_Jinkela_wire_11274)
    );

    bfr new_Jinkela_buffer_12993 (
        .din(new_Jinkela_wire_15522),
        .dout(new_Jinkela_wire_15523)
    );

    bfr new_Jinkela_buffer_9204 (
        .din(new_Jinkela_wire_11223),
        .dout(new_Jinkela_wire_11224)
    );

    bfr new_Jinkela_buffer_12674 (
        .din(new_Jinkela_wire_15189),
        .dout(new_Jinkela_wire_15190)
    );

    bfr new_Jinkela_buffer_9336 (
        .din(new_Jinkela_wire_11365),
        .dout(new_Jinkela_wire_11366)
    );

    bfr new_Jinkela_buffer_12880 (
        .din(new_Jinkela_wire_15401),
        .dout(new_Jinkela_wire_15402)
    );

    bfr new_Jinkela_buffer_12715 (
        .din(new_Jinkela_wire_15236),
        .dout(new_Jinkela_wire_15237)
    );

    bfr new_Jinkela_buffer_9205 (
        .din(new_Jinkela_wire_11224),
        .dout(new_Jinkela_wire_11225)
    );

    bfr new_Jinkela_buffer_12675 (
        .din(new_Jinkela_wire_15190),
        .dout(new_Jinkela_wire_15191)
    );

    bfr new_Jinkela_buffer_9251 (
        .din(new_Jinkela_wire_11274),
        .dout(new_Jinkela_wire_11275)
    );

    bfr new_Jinkela_buffer_12872 (
        .din(new_Jinkela_wire_15393),
        .dout(new_Jinkela_wire_15394)
    );

    spl2 new_Jinkela_splitter_859 (
        .a(new_Jinkela_wire_11225),
        .b(new_Jinkela_wire_11226),
        .c(new_Jinkela_wire_11227)
    );

    bfr new_Jinkela_buffer_12676 (
        .din(new_Jinkela_wire_15191),
        .dout(new_Jinkela_wire_15192)
    );

    bfr new_Jinkela_buffer_9252 (
        .din(new_Jinkela_wire_11275),
        .dout(new_Jinkela_wire_11276)
    );

    bfr new_Jinkela_buffer_12716 (
        .din(new_Jinkela_wire_15237),
        .dout(new_Jinkela_wire_15238)
    );

    spl2 new_Jinkela_splitter_876 (
        .a(_0413_),
        .b(new_Jinkela_wire_11414),
        .c(new_Jinkela_wire_11415)
    );

    bfr new_Jinkela_buffer_12677 (
        .din(new_Jinkela_wire_15192),
        .dout(new_Jinkela_wire_15193)
    );

    spl2 new_Jinkela_splitter_875 (
        .a(_0345_),
        .b(new_Jinkela_wire_11412),
        .c(new_Jinkela_wire_11413)
    );

    bfr new_Jinkela_buffer_9337 (
        .din(new_Jinkela_wire_11366),
        .dout(new_Jinkela_wire_11367)
    );

    bfr new_Jinkela_buffer_9253 (
        .din(new_Jinkela_wire_11276),
        .dout(new_Jinkela_wire_11277)
    );

    bfr new_Jinkela_buffer_12678 (
        .din(new_Jinkela_wire_15193),
        .dout(new_Jinkela_wire_15194)
    );

    bfr new_Jinkela_buffer_12717 (
        .din(new_Jinkela_wire_15238),
        .dout(new_Jinkela_wire_15239)
    );

    bfr new_Jinkela_buffer_9254 (
        .din(new_Jinkela_wire_11277),
        .dout(new_Jinkela_wire_11278)
    );

    bfr new_Jinkela_buffer_12679 (
        .din(new_Jinkela_wire_15194),
        .dout(new_Jinkela_wire_15195)
    );

    bfr new_Jinkela_buffer_9338 (
        .din(new_Jinkela_wire_11367),
        .dout(new_Jinkela_wire_11368)
    );

    bfr new_Jinkela_buffer_12949 (
        .din(new_Jinkela_wire_15472),
        .dout(new_Jinkela_wire_15473)
    );

    bfr new_Jinkela_buffer_9255 (
        .din(new_Jinkela_wire_11278),
        .dout(new_Jinkela_wire_11279)
    );

    bfr new_Jinkela_buffer_12680 (
        .din(new_Jinkela_wire_15195),
        .dout(new_Jinkela_wire_15196)
    );

    bfr new_Jinkela_buffer_12881 (
        .din(new_Jinkela_wire_15402),
        .dout(new_Jinkela_wire_15403)
    );

    spl2 new_Jinkela_splitter_877 (
        .a(_0682_),
        .b(new_Jinkela_wire_11416),
        .c(new_Jinkela_wire_11417)
    );

    bfr new_Jinkela_buffer_12718 (
        .din(new_Jinkela_wire_15239),
        .dout(new_Jinkela_wire_15240)
    );

    bfr new_Jinkela_buffer_9256 (
        .din(new_Jinkela_wire_11279),
        .dout(new_Jinkela_wire_11280)
    );

    bfr new_Jinkela_buffer_12681 (
        .din(new_Jinkela_wire_15196),
        .dout(new_Jinkela_wire_15197)
    );

    bfr new_Jinkela_buffer_9339 (
        .din(new_Jinkela_wire_11368),
        .dout(new_Jinkela_wire_11369)
    );

    bfr new_Jinkela_buffer_9257 (
        .din(new_Jinkela_wire_11280),
        .dout(new_Jinkela_wire_11281)
    );

    spl2 new_Jinkela_splitter_1107 (
        .a(new_Jinkela_wire_15197),
        .b(new_Jinkela_wire_15198),
        .c(new_Jinkela_wire_15199)
    );

    spl2 new_Jinkela_splitter_878 (
        .a(_0266_),
        .b(new_Jinkela_wire_11422),
        .c(new_Jinkela_wire_11423)
    );

    bfr new_Jinkela_buffer_12997 (
        .din(_0296_),
        .dout(new_Jinkela_wire_15527)
    );

    bfr new_Jinkela_buffer_9258 (
        .din(new_Jinkela_wire_11281),
        .dout(new_Jinkela_wire_11282)
    );

    bfr new_Jinkela_buffer_12719 (
        .din(new_Jinkela_wire_15240),
        .dout(new_Jinkela_wire_15241)
    );

    bfr new_Jinkela_buffer_2282 (
        .din(new_Jinkela_wire_3263),
        .dout(new_Jinkela_wire_3264)
    );

    bfr new_Jinkela_buffer_2136 (
        .din(new_Jinkela_wire_3077),
        .dout(new_Jinkela_wire_3078)
    );

    bfr new_Jinkela_buffer_2226 (
        .din(new_Jinkela_wire_3175),
        .dout(new_Jinkela_wire_3176)
    );

    bfr new_Jinkela_buffer_2137 (
        .din(new_Jinkela_wire_3078),
        .dout(new_Jinkela_wire_3079)
    );

    bfr new_Jinkela_buffer_2253 (
        .din(new_Jinkela_wire_3218),
        .dout(new_Jinkela_wire_3219)
    );

    bfr new_Jinkela_buffer_2138 (
        .din(new_Jinkela_wire_3079),
        .dout(new_Jinkela_wire_3080)
    );

    bfr new_Jinkela_buffer_2227 (
        .din(new_Jinkela_wire_3176),
        .dout(new_Jinkela_wire_3177)
    );

    bfr new_Jinkela_buffer_2139 (
        .din(new_Jinkela_wire_3080),
        .dout(new_Jinkela_wire_3081)
    );

    bfr new_Jinkela_buffer_2140 (
        .din(new_Jinkela_wire_3081),
        .dout(new_Jinkela_wire_3082)
    );

    bfr new_Jinkela_buffer_2371 (
        .din(_0108_),
        .dout(new_Jinkela_wire_3363)
    );

    spl2 new_Jinkela_splitter_324 (
        .a(new_Jinkela_wire_3177),
        .b(new_Jinkela_wire_3178),
        .c(new_Jinkela_wire_3179)
    );

    bfr new_Jinkela_buffer_2141 (
        .din(new_Jinkela_wire_3082),
        .dout(new_Jinkela_wire_3083)
    );

    bfr new_Jinkela_buffer_2283 (
        .din(new_Jinkela_wire_3264),
        .dout(new_Jinkela_wire_3265)
    );

    bfr new_Jinkela_buffer_2142 (
        .din(new_Jinkela_wire_3083),
        .dout(new_Jinkela_wire_3084)
    );

    bfr new_Jinkela_buffer_2254 (
        .din(new_Jinkela_wire_3219),
        .dout(new_Jinkela_wire_3220)
    );

    bfr new_Jinkela_buffer_2143 (
        .din(new_Jinkela_wire_3084),
        .dout(new_Jinkela_wire_3085)
    );

    bfr new_Jinkela_buffer_2255 (
        .din(new_Jinkela_wire_3220),
        .dout(new_Jinkela_wire_3221)
    );

    bfr new_Jinkela_buffer_2144 (
        .din(new_Jinkela_wire_3085),
        .dout(new_Jinkela_wire_3086)
    );

    bfr new_Jinkela_buffer_2286 (
        .din(new_Jinkela_wire_3273),
        .dout(new_Jinkela_wire_3274)
    );

    bfr new_Jinkela_buffer_2145 (
        .din(new_Jinkela_wire_3086),
        .dout(new_Jinkela_wire_3087)
    );

    bfr new_Jinkela_buffer_2256 (
        .din(new_Jinkela_wire_3221),
        .dout(new_Jinkela_wire_3222)
    );

    bfr new_Jinkela_buffer_2146 (
        .din(new_Jinkela_wire_3087),
        .dout(new_Jinkela_wire_3088)
    );

    bfr new_Jinkela_buffer_2284 (
        .din(new_Jinkela_wire_3265),
        .dout(new_Jinkela_wire_3266)
    );

    bfr new_Jinkela_buffer_2147 (
        .din(new_Jinkela_wire_3088),
        .dout(new_Jinkela_wire_3089)
    );

    bfr new_Jinkela_buffer_2257 (
        .din(new_Jinkela_wire_3222),
        .dout(new_Jinkela_wire_3223)
    );

    bfr new_Jinkela_buffer_2148 (
        .din(new_Jinkela_wire_3089),
        .dout(new_Jinkela_wire_3090)
    );

    spl2 new_Jinkela_splitter_347 (
        .a(_1542_),
        .b(new_Jinkela_wire_3429),
        .c(new_Jinkela_wire_3430)
    );

    bfr new_Jinkela_buffer_2149 (
        .din(new_Jinkela_wire_3090),
        .dout(new_Jinkela_wire_3091)
    );

    bfr new_Jinkela_buffer_2258 (
        .din(new_Jinkela_wire_3223),
        .dout(new_Jinkela_wire_3224)
    );

    bfr new_Jinkela_buffer_2150 (
        .din(new_Jinkela_wire_3091),
        .dout(new_Jinkela_wire_3092)
    );

    spl2 new_Jinkela_splitter_340 (
        .a(new_Jinkela_wire_3266),
        .b(new_Jinkela_wire_3267),
        .c(new_Jinkela_wire_3268)
    );

    bfr new_Jinkela_buffer_2151 (
        .din(new_Jinkela_wire_3092),
        .dout(new_Jinkela_wire_3093)
    );

    bfr new_Jinkela_buffer_2259 (
        .din(new_Jinkela_wire_3224),
        .dout(new_Jinkela_wire_3225)
    );

    bfr new_Jinkela_buffer_2152 (
        .din(new_Jinkela_wire_3093),
        .dout(new_Jinkela_wire_3094)
    );

    bfr new_Jinkela_buffer_2153 (
        .din(new_Jinkela_wire_3094),
        .dout(new_Jinkela_wire_3095)
    );

    bfr new_Jinkela_buffer_2393 (
        .din(_1288_),
        .dout(new_Jinkela_wire_3387)
    );

    bfr new_Jinkela_buffer_2260 (
        .din(new_Jinkela_wire_3225),
        .dout(new_Jinkela_wire_3226)
    );

    bfr new_Jinkela_buffer_2154 (
        .din(new_Jinkela_wire_3095),
        .dout(new_Jinkela_wire_3096)
    );

    bfr new_Jinkela_buffer_2287 (
        .din(new_Jinkela_wire_3274),
        .dout(new_Jinkela_wire_3275)
    );

    bfr new_Jinkela_buffer_2155 (
        .din(new_Jinkela_wire_3096),
        .dout(new_Jinkela_wire_3097)
    );

    bfr new_Jinkela_buffer_2261 (
        .din(new_Jinkela_wire_3226),
        .dout(new_Jinkela_wire_3227)
    );

    bfr new_Jinkela_buffer_2156 (
        .din(new_Jinkela_wire_3097),
        .dout(new_Jinkela_wire_3098)
    );

    and_bb _3214_ (
        .a(new_Jinkela_wire_13309),
        .b(new_Jinkela_wire_1897),
        .c(_0483_)
    );

    or_bb _3215_ (
        .a(new_Jinkela_wire_18289),
        .b(new_Jinkela_wire_16961),
        .c(_0484_)
    );

    and_ii _3216_ (
        .a(new_Jinkela_wire_15695),
        .b(new_Jinkela_wire_15198),
        .c(_0485_)
    );

    and_bb _3217_ (
        .a(new_Jinkela_wire_15696),
        .b(new_Jinkela_wire_15199),
        .c(_0486_)
    );

    or_bb _3218_ (
        .a(new_Jinkela_wire_15745),
        .b(new_Jinkela_wire_4711),
        .c(_0487_)
    );

    and_ii _3219_ (
        .a(new_Jinkela_wire_20322),
        .b(new_Jinkela_wire_2016),
        .c(_0488_)
    );

    and_bb _3220_ (
        .a(new_Jinkela_wire_20323),
        .b(new_Jinkela_wire_2017),
        .c(_0489_)
    );

    or_bb _3221_ (
        .a(new_Jinkela_wire_14274),
        .b(new_Jinkela_wire_18111),
        .c(_0490_)
    );

    and_ii _3222_ (
        .a(new_Jinkela_wire_14028),
        .b(new_Jinkela_wire_20131),
        .c(_0491_)
    );

    and_bb _3223_ (
        .a(new_Jinkela_wire_14029),
        .b(new_Jinkela_wire_20132),
        .c(_0493_)
    );

    or_bb _3224_ (
        .a(new_Jinkela_wire_15121),
        .b(new_Jinkela_wire_19542),
        .c(_0494_)
    );

    and_ii _3225_ (
        .a(new_Jinkela_wire_7833),
        .b(new_Jinkela_wire_8178),
        .c(_0495_)
    );

    and_bb _3226_ (
        .a(new_Jinkela_wire_7834),
        .b(new_Jinkela_wire_8179),
        .c(_0496_)
    );

    or_bb _3227_ (
        .a(new_Jinkela_wire_21180),
        .b(new_Jinkela_wire_12717),
        .c(_0497_)
    );

    and_ii _3228_ (
        .a(new_Jinkela_wire_10099),
        .b(new_Jinkela_wire_5416),
        .c(_0498_)
    );

    and_bb _3229_ (
        .a(new_Jinkela_wire_10100),
        .b(new_Jinkela_wire_5417),
        .c(_0499_)
    );

    or_bb _3230_ (
        .a(new_Jinkela_wire_18833),
        .b(new_Jinkela_wire_14214),
        .c(_0500_)
    );

    and_ii _3231_ (
        .a(new_Jinkela_wire_4999),
        .b(new_Jinkela_wire_19556),
        .c(_0501_)
    );

    and_bb _3232_ (
        .a(new_Jinkela_wire_5000),
        .b(new_Jinkela_wire_19557),
        .c(_0502_)
    );

    or_bb _3233_ (
        .a(new_Jinkela_wire_5802),
        .b(new_Jinkela_wire_9558),
        .c(_0504_)
    );

    and_ii _3234_ (
        .a(new_Jinkela_wire_17051),
        .b(new_Jinkela_wire_11823),
        .c(_0505_)
    );

    and_bb _3235_ (
        .a(new_Jinkela_wire_17052),
        .b(new_Jinkela_wire_11824),
        .c(_0506_)
    );

    or_bb _3236_ (
        .a(new_Jinkela_wire_12051),
        .b(new_Jinkela_wire_15683),
        .c(_0507_)
    );

    and_ii _3237_ (
        .a(new_Jinkela_wire_1136),
        .b(new_Jinkela_wire_10397),
        .c(_0508_)
    );

    and_bb _3238_ (
        .a(new_Jinkela_wire_1137),
        .b(new_Jinkela_wire_10398),
        .c(_0509_)
    );

    or_bb _3239_ (
        .a(new_Jinkela_wire_11839),
        .b(new_Jinkela_wire_13984),
        .c(_0510_)
    );

    and_ii _3240_ (
        .a(new_Jinkela_wire_14199),
        .b(new_Jinkela_wire_18101),
        .c(_0511_)
    );

    and_bb _3241_ (
        .a(new_Jinkela_wire_14200),
        .b(new_Jinkela_wire_18102),
        .c(_0512_)
    );

    or_bb _3242_ (
        .a(new_Jinkela_wire_1618),
        .b(new_Jinkela_wire_2960),
        .c(_0513_)
    );

    and_ii _3243_ (
        .a(new_Jinkela_wire_10259),
        .b(new_Jinkela_wire_11136),
        .c(_0515_)
    );

    and_bb _3244_ (
        .a(new_Jinkela_wire_10260),
        .b(new_Jinkela_wire_11137),
        .c(_0516_)
    );

    or_bb _3245_ (
        .a(new_Jinkela_wire_18534),
        .b(new_Jinkela_wire_18573),
        .c(_0517_)
    );

    and_ii _3246_ (
        .a(new_Jinkela_wire_5465),
        .b(new_Jinkela_wire_19906),
        .c(_0518_)
    );

    and_bb _3247_ (
        .a(new_Jinkela_wire_5466),
        .b(new_Jinkela_wire_19907),
        .c(_0519_)
    );

    or_bb _3248_ (
        .a(new_Jinkela_wire_8363),
        .b(new_Jinkela_wire_4675),
        .c(_0520_)
    );

    and_ii _3249_ (
        .a(new_Jinkela_wire_3886),
        .b(new_Jinkela_wire_1763),
        .c(_0521_)
    );

    and_bb _3250_ (
        .a(new_Jinkela_wire_3887),
        .b(new_Jinkela_wire_1764),
        .c(_0522_)
    );

    and_ii _3251_ (
        .a(new_Jinkela_wire_7287),
        .b(new_Jinkela_wire_4303),
        .c(_0523_)
    );

    and_bb _3252_ (
        .a(new_Jinkela_wire_9362),
        .b(new_Jinkela_wire_9099),
        .c(_0524_)
    );

    and_ii _3253_ (
        .a(new_Jinkela_wire_9363),
        .b(new_Jinkela_wire_9100),
        .c(_0526_)
    );

    or_bb _3254_ (
        .a(new_Jinkela_wire_20048),
        .b(new_Jinkela_wire_10079),
        .c(new_net_3970)
    );

    or_bb _3255_ (
        .a(new_Jinkela_wire_10080),
        .b(new_Jinkela_wire_4320),
        .c(_0527_)
    );

    bfr new_Jinkela_buffer_16108 (
        .din(new_Jinkela_wire_19232),
        .dout(new_Jinkela_wire_19233)
    );

    bfr new_Jinkela_buffer_16182 (
        .din(new_Jinkela_wire_19330),
        .dout(new_Jinkela_wire_19331)
    );

    bfr new_Jinkela_buffer_16109 (
        .din(new_Jinkela_wire_19233),
        .dout(new_Jinkela_wire_19234)
    );

    bfr new_Jinkela_buffer_16171 (
        .din(new_Jinkela_wire_19309),
        .dout(new_Jinkela_wire_19310)
    );

    bfr new_Jinkela_buffer_16110 (
        .din(new_Jinkela_wire_19234),
        .dout(new_Jinkela_wire_19235)
    );

    bfr new_Jinkela_buffer_16186 (
        .din(new_Jinkela_wire_19336),
        .dout(new_Jinkela_wire_19337)
    );

    bfr new_Jinkela_buffer_16111 (
        .din(new_Jinkela_wire_19235),
        .dout(new_Jinkela_wire_19236)
    );

    bfr new_Jinkela_buffer_16172 (
        .din(new_Jinkela_wire_19310),
        .dout(new_Jinkela_wire_19311)
    );

    bfr new_Jinkela_buffer_16112 (
        .din(new_Jinkela_wire_19236),
        .dout(new_Jinkela_wire_19237)
    );

    bfr new_Jinkela_buffer_16183 (
        .din(new_Jinkela_wire_19331),
        .dout(new_Jinkela_wire_19332)
    );

    bfr new_Jinkela_buffer_16113 (
        .din(new_Jinkela_wire_19237),
        .dout(new_Jinkela_wire_19238)
    );

    bfr new_Jinkela_buffer_16173 (
        .din(new_Jinkela_wire_19311),
        .dout(new_Jinkela_wire_19312)
    );

    bfr new_Jinkela_buffer_16114 (
        .din(new_Jinkela_wire_19238),
        .dout(new_Jinkela_wire_19239)
    );

    spl2 new_Jinkela_splitter_1424 (
        .a(_1051_),
        .b(new_Jinkela_wire_19342),
        .c(new_Jinkela_wire_19343)
    );

    bfr new_Jinkela_buffer_16115 (
        .din(new_Jinkela_wire_19239),
        .dout(new_Jinkela_wire_19240)
    );

    bfr new_Jinkela_buffer_16174 (
        .din(new_Jinkela_wire_19312),
        .dout(new_Jinkela_wire_19313)
    );

    bfr new_Jinkela_buffer_16116 (
        .din(new_Jinkela_wire_19240),
        .dout(new_Jinkela_wire_19241)
    );

    bfr new_Jinkela_buffer_16184 (
        .din(new_Jinkela_wire_19332),
        .dout(new_Jinkela_wire_19333)
    );

    bfr new_Jinkela_buffer_16117 (
        .din(new_Jinkela_wire_19241),
        .dout(new_Jinkela_wire_19242)
    );

    bfr new_Jinkela_buffer_16175 (
        .din(new_Jinkela_wire_19313),
        .dout(new_Jinkela_wire_19314)
    );

    bfr new_Jinkela_buffer_16118 (
        .din(new_Jinkela_wire_19242),
        .dout(new_Jinkela_wire_19243)
    );

    spl2 new_Jinkela_splitter_1425 (
        .a(_0098_),
        .b(new_Jinkela_wire_19344),
        .c(new_Jinkela_wire_19345)
    );

    bfr new_Jinkela_buffer_16192 (
        .din(_0346_),
        .dout(new_Jinkela_wire_19353)
    );

    bfr new_Jinkela_buffer_16119 (
        .din(new_Jinkela_wire_19243),
        .dout(new_Jinkela_wire_19244)
    );

    bfr new_Jinkela_buffer_16176 (
        .din(new_Jinkela_wire_19314),
        .dout(new_Jinkela_wire_19315)
    );

    bfr new_Jinkela_buffer_16120 (
        .din(new_Jinkela_wire_19244),
        .dout(new_Jinkela_wire_19245)
    );

    bfr new_Jinkela_buffer_16187 (
        .din(new_Jinkela_wire_19337),
        .dout(new_Jinkela_wire_19338)
    );

    bfr new_Jinkela_buffer_16121 (
        .din(new_Jinkela_wire_19245),
        .dout(new_Jinkela_wire_19246)
    );

    spl2 new_Jinkela_splitter_1418 (
        .a(new_Jinkela_wire_19315),
        .b(new_Jinkela_wire_19316),
        .c(new_Jinkela_wire_19317)
    );

    bfr new_Jinkela_buffer_16122 (
        .din(new_Jinkela_wire_19246),
        .dout(new_Jinkela_wire_19247)
    );

    bfr new_Jinkela_buffer_16188 (
        .din(new_Jinkela_wire_19338),
        .dout(new_Jinkela_wire_19339)
    );

    bfr new_Jinkela_buffer_16123 (
        .din(new_Jinkela_wire_19247),
        .dout(new_Jinkela_wire_19248)
    );

    bfr new_Jinkela_buffer_16124 (
        .din(new_Jinkela_wire_19248),
        .dout(new_Jinkela_wire_19249)
    );

    bfr new_Jinkela_buffer_16191 (
        .din(_0479_),
        .dout(new_Jinkela_wire_19346)
    );

    bfr new_Jinkela_buffer_16125 (
        .din(new_Jinkela_wire_19249),
        .dout(new_Jinkela_wire_19250)
    );

    bfr new_Jinkela_buffer_16189 (
        .din(new_Jinkela_wire_19339),
        .dout(new_Jinkela_wire_19340)
    );

    bfr new_Jinkela_buffer_16126 (
        .din(new_Jinkela_wire_19250),
        .dout(new_Jinkela_wire_19251)
    );

    spl2 new_Jinkela_splitter_1427 (
        .a(_0464_),
        .b(new_Jinkela_wire_19349),
        .c(new_Jinkela_wire_19350)
    );

    spl2 new_Jinkela_splitter_1426 (
        .a(_1334_),
        .b(new_Jinkela_wire_19347),
        .c(new_Jinkela_wire_19348)
    );

    bfr new_Jinkela_buffer_16127 (
        .din(new_Jinkela_wire_19251),
        .dout(new_Jinkela_wire_19252)
    );

    bfr new_Jinkela_buffer_16128 (
        .din(new_Jinkela_wire_19252),
        .dout(new_Jinkela_wire_19253)
    );

    spl2 new_Jinkela_splitter_1428 (
        .a(_0813_),
        .b(new_Jinkela_wire_19351),
        .c(new_Jinkela_wire_19352)
    );

    and_bb _2329_ (
        .a(new_Jinkela_wire_115),
        .b(new_Jinkela_wire_563),
        .c(_1365_)
    );

    bfr new_Jinkela_buffer_2288 (
        .din(new_Jinkela_wire_3275),
        .dout(new_Jinkela_wire_3276)
    );

    and_bi _2330_ (
        .a(new_Jinkela_wire_10090),
        .b(new_Jinkela_wire_20395),
        .c(_1366_)
    );

    bfr new_Jinkela_buffer_2157 (
        .din(new_Jinkela_wire_3098),
        .dout(new_Jinkela_wire_3099)
    );

    and_bb _2331_ (
        .a(new_Jinkela_wire_282),
        .b(new_Jinkela_wire_14),
        .c(_1367_)
    );

    bfr new_Jinkela_buffer_2262 (
        .din(new_Jinkela_wire_3227),
        .dout(new_Jinkela_wire_3228)
    );

    and_bi _2332_ (
        .a(new_Jinkela_wire_19149),
        .b(new_Jinkela_wire_2463),
        .c(_1368_)
    );

    bfr new_Jinkela_buffer_2158 (
        .din(new_Jinkela_wire_3099),
        .dout(new_Jinkela_wire_3100)
    );

    and_bb _2333_ (
        .a(new_Jinkela_wire_70),
        .b(new_Jinkela_wire_444),
        .c(_1369_)
    );

    bfr new_Jinkela_buffer_2372 (
        .din(new_Jinkela_wire_3363),
        .dout(new_Jinkela_wire_3364)
    );

    and_bi _2334_ (
        .a(new_Jinkela_wire_18968),
        .b(new_Jinkela_wire_13066),
        .c(_1370_)
    );

    bfr new_Jinkela_buffer_2159 (
        .din(new_Jinkela_wire_3100),
        .dout(new_Jinkela_wire_3101)
    );

    and_bb _2335_ (
        .a(new_Jinkela_wire_484),
        .b(new_Jinkela_wire_246),
        .c(_1371_)
    );

    bfr new_Jinkela_buffer_2263 (
        .din(new_Jinkela_wire_3228),
        .dout(new_Jinkela_wire_3229)
    );

    and_bi _2336_ (
        .a(new_Jinkela_wire_1911),
        .b(new_Jinkela_wire_8279),
        .c(_1372_)
    );

    bfr new_Jinkela_buffer_2160 (
        .din(new_Jinkela_wire_3101),
        .dout(new_Jinkela_wire_3102)
    );

    and_bb _2337_ (
        .a(new_Jinkela_wire_358),
        .b(new_Jinkela_wire_289),
        .c(_1373_)
    );

    bfr new_Jinkela_buffer_2289 (
        .din(new_Jinkela_wire_3276),
        .dout(new_Jinkela_wire_3277)
    );

    and_bi _2338_ (
        .a(new_Jinkela_wire_18386),
        .b(new_Jinkela_wire_5732),
        .c(_1374_)
    );

    bfr new_Jinkela_buffer_2161 (
        .din(new_Jinkela_wire_3102),
        .dout(new_Jinkela_wire_3103)
    );

    and_bb _2339_ (
        .a(new_Jinkela_wire_700),
        .b(new_Jinkela_wire_64),
        .c(_1375_)
    );

    bfr new_Jinkela_buffer_2264 (
        .din(new_Jinkela_wire_3229),
        .dout(new_Jinkela_wire_3230)
    );

    and_bi _2340_ (
        .a(new_Jinkela_wire_11439),
        .b(new_Jinkela_wire_12716),
        .c(_1376_)
    );

    bfr new_Jinkela_buffer_2162 (
        .din(new_Jinkela_wire_3103),
        .dout(new_Jinkela_wire_3104)
    );

    and_bb _2341_ (
        .a(new_Jinkela_wire_657),
        .b(new_Jinkela_wire_488),
        .c(_1377_)
    );

    and_bi _2342_ (
        .a(new_Jinkela_wire_5427),
        .b(new_Jinkela_wire_7317),
        .c(_1378_)
    );

    bfr new_Jinkela_buffer_2163 (
        .din(new_Jinkela_wire_3104),
        .dout(new_Jinkela_wire_3105)
    );

    and_bb _2343_ (
        .a(new_Jinkela_wire_628),
        .b(new_Jinkela_wire_36),
        .c(_1379_)
    );

    spl2 new_Jinkela_splitter_348 (
        .a(_0692_),
        .b(new_Jinkela_wire_3435),
        .c(new_Jinkela_wire_3436)
    );

    bfr new_Jinkela_buffer_2265 (
        .din(new_Jinkela_wire_3230),
        .dout(new_Jinkela_wire_3231)
    );

    and_bi _2344_ (
        .a(new_Jinkela_wire_13146),
        .b(new_Jinkela_wire_4727),
        .c(_1380_)
    );

    bfr new_Jinkela_buffer_2164 (
        .din(new_Jinkela_wire_3105),
        .dout(new_Jinkela_wire_3106)
    );

    and_bb _2345_ (
        .a(new_Jinkela_wire_185),
        .b(new_Jinkela_wire_540),
        .c(_1381_)
    );

    bfr new_Jinkela_buffer_2290 (
        .din(new_Jinkela_wire_3277),
        .dout(new_Jinkela_wire_3278)
    );

    or_ii _2346_ (
        .a(new_Jinkela_wire_395),
        .b(new_Jinkela_wire_313),
        .c(_1382_)
    );

    bfr new_Jinkela_buffer_2165 (
        .din(new_Jinkela_wire_3106),
        .dout(new_Jinkela_wire_3107)
    );

    and_bi _2347_ (
        .a(new_Jinkela_wire_1622),
        .b(new_Jinkela_wire_4831),
        .c(_1383_)
    );

    bfr new_Jinkela_buffer_2266 (
        .din(new_Jinkela_wire_3231),
        .dout(new_Jinkela_wire_3232)
    );

    and_bb _2348_ (
        .a(new_Jinkela_wire_410),
        .b(new_Jinkela_wire_228),
        .c(_1384_)
    );

    bfr new_Jinkela_buffer_2166 (
        .din(new_Jinkela_wire_3107),
        .dout(new_Jinkela_wire_3108)
    );

    and_bi _2349_ (
        .a(new_Jinkela_wire_18524),
        .b(new_Jinkela_wire_15669),
        .c(_1385_)
    );

    bfr new_Jinkela_buffer_2373 (
        .din(new_Jinkela_wire_3364),
        .dout(new_Jinkela_wire_3365)
    );

    and_ii _2350_ (
        .a(new_Jinkela_wire_1623),
        .b(new_Jinkela_wire_9012),
        .c(_1386_)
    );

    bfr new_Jinkela_buffer_2167 (
        .din(new_Jinkela_wire_3108),
        .dout(new_Jinkela_wire_3109)
    );

    or_bb _2351_ (
        .a(new_Jinkela_wire_20275),
        .b(new_Jinkela_wire_20045),
        .c(_1387_)
    );

    bfr new_Jinkela_buffer_2267 (
        .din(new_Jinkela_wire_3232),
        .dout(new_Jinkela_wire_3233)
    );

    or_ii _2352_ (
        .a(new_Jinkela_wire_20276),
        .b(new_Jinkela_wire_20044),
        .c(_1388_)
    );

    bfr new_Jinkela_buffer_2168 (
        .din(new_Jinkela_wire_3109),
        .dout(new_Jinkela_wire_3110)
    );

    or_ii _2353_ (
        .a(new_Jinkela_wire_14085),
        .b(new_Jinkela_wire_5161),
        .c(_1389_)
    );

    bfr new_Jinkela_buffer_2291 (
        .din(new_Jinkela_wire_3278),
        .dout(new_Jinkela_wire_3279)
    );

    and_ii _2354_ (
        .a(new_Jinkela_wire_836),
        .b(new_Jinkela_wire_20803),
        .c(_1390_)
    );

    bfr new_Jinkela_buffer_2169 (
        .din(new_Jinkela_wire_3110),
        .dout(new_Jinkela_wire_3111)
    );

    and_bb _2355_ (
        .a(new_Jinkela_wire_837),
        .b(new_Jinkela_wire_20804),
        .c(_1391_)
    );

    bfr new_Jinkela_buffer_2268 (
        .din(new_Jinkela_wire_3233),
        .dout(new_Jinkela_wire_3234)
    );

    or_bb _2356_ (
        .a(new_Jinkela_wire_17062),
        .b(new_Jinkela_wire_6857),
        .c(_1392_)
    );

    bfr new_Jinkela_buffer_2170 (
        .din(new_Jinkela_wire_3111),
        .dout(new_Jinkela_wire_3112)
    );

    or_bb _2357_ (
        .a(new_Jinkela_wire_5104),
        .b(new_Jinkela_wire_1788),
        .c(_1393_)
    );

    bfr new_Jinkela_buffer_2394 (
        .din(new_Jinkela_wire_3387),
        .dout(new_Jinkela_wire_3388)
    );

    or_ii _2358_ (
        .a(new_Jinkela_wire_5105),
        .b(new_Jinkela_wire_1789),
        .c(_1394_)
    );

    bfr new_Jinkela_buffer_2171 (
        .din(new_Jinkela_wire_3112),
        .dout(new_Jinkela_wire_3113)
    );

    or_ii _2359_ (
        .a(new_Jinkela_wire_7717),
        .b(new_Jinkela_wire_3880),
        .c(_1395_)
    );

    bfr new_Jinkela_buffer_2269 (
        .din(new_Jinkela_wire_3234),
        .dout(new_Jinkela_wire_3235)
    );

    and_ii _2360_ (
        .a(new_Jinkela_wire_13201),
        .b(new_Jinkela_wire_5124),
        .c(_1396_)
    );

    bfr new_Jinkela_buffer_2292 (
        .din(new_Jinkela_wire_3279),
        .dout(new_Jinkela_wire_3280)
    );

    and_bb _2361_ (
        .a(new_Jinkela_wire_13202),
        .b(new_Jinkela_wire_5125),
        .c(_1397_)
    );

    bfr new_Jinkela_buffer_2270 (
        .din(new_Jinkela_wire_3235),
        .dout(new_Jinkela_wire_3236)
    );

    or_bb _2362_ (
        .a(new_Jinkela_wire_4661),
        .b(new_Jinkela_wire_4080),
        .c(_1398_)
    );

    bfr new_Jinkela_buffer_2374 (
        .din(new_Jinkela_wire_3365),
        .dout(new_Jinkela_wire_3366)
    );

    or_bb _2363_ (
        .a(new_Jinkela_wire_841),
        .b(new_Jinkela_wire_19554),
        .c(_1399_)
    );

    spl2 new_Jinkela_splitter_332 (
        .a(new_Jinkela_wire_3236),
        .b(new_Jinkela_wire_3237),
        .c(new_Jinkela_wire_3238)
    );

    or_ii _2364_ (
        .a(new_Jinkela_wire_842),
        .b(new_Jinkela_wire_19555),
        .c(_1400_)
    );

    or_ii _2365_ (
        .a(new_Jinkela_wire_13306),
        .b(new_Jinkela_wire_15521),
        .c(_1401_)
    );

    bfr new_Jinkela_buffer_2433 (
        .din(new_Jinkela_wire_3430),
        .dout(new_Jinkela_wire_3431)
    );

    bfr new_Jinkela_buffer_2293 (
        .din(new_Jinkela_wire_3280),
        .dout(new_Jinkela_wire_3281)
    );

    and_ii _2366_ (
        .a(new_Jinkela_wire_6407),
        .b(new_Jinkela_wire_13717),
        .c(_1402_)
    );

    bfr new_Jinkela_buffer_2294 (
        .din(new_Jinkela_wire_3281),
        .dout(new_Jinkela_wire_3282)
    );

    and_bb _2367_ (
        .a(new_Jinkela_wire_6408),
        .b(new_Jinkela_wire_13718),
        .c(_1403_)
    );

    bfr new_Jinkela_buffer_2375 (
        .din(new_Jinkela_wire_3366),
        .dout(new_Jinkela_wire_3367)
    );

    or_bb _2368_ (
        .a(new_Jinkela_wire_11726),
        .b(new_Jinkela_wire_16514),
        .c(_1404_)
    );

    bfr new_Jinkela_buffer_2295 (
        .din(new_Jinkela_wire_3282),
        .dout(new_Jinkela_wire_3283)
    );

    or_bb _2369_ (
        .a(new_Jinkela_wire_17658),
        .b(new_Jinkela_wire_14024),
        .c(_1405_)
    );

    bfr new_Jinkela_buffer_2395 (
        .din(new_Jinkela_wire_3388),
        .dout(new_Jinkela_wire_3389)
    );

    or_ii _2370_ (
        .a(new_Jinkela_wire_17659),
        .b(new_Jinkela_wire_14025),
        .c(_1406_)
    );

    bfr new_Jinkela_buffer_5761 (
        .din(new_Jinkela_wire_7350),
        .dout(new_Jinkela_wire_7351)
    );

    bfr new_Jinkela_buffer_5862 (
        .din(new_Jinkela_wire_7459),
        .dout(new_Jinkela_wire_7460)
    );

    bfr new_Jinkela_buffer_5762 (
        .din(new_Jinkela_wire_7351),
        .dout(new_Jinkela_wire_7352)
    );

    bfr new_Jinkela_buffer_5973 (
        .din(_1723_),
        .dout(new_Jinkela_wire_7583)
    );

    bfr new_Jinkela_buffer_5763 (
        .din(new_Jinkela_wire_7352),
        .dout(new_Jinkela_wire_7353)
    );

    bfr new_Jinkela_buffer_5863 (
        .din(new_Jinkela_wire_7460),
        .dout(new_Jinkela_wire_7461)
    );

    bfr new_Jinkela_buffer_5764 (
        .din(new_Jinkela_wire_7353),
        .dout(new_Jinkela_wire_7354)
    );

    bfr new_Jinkela_buffer_5906 (
        .din(new_Jinkela_wire_7509),
        .dout(new_Jinkela_wire_7510)
    );

    bfr new_Jinkela_buffer_5765 (
        .din(new_Jinkela_wire_7354),
        .dout(new_Jinkela_wire_7355)
    );

    bfr new_Jinkela_buffer_5864 (
        .din(new_Jinkela_wire_7461),
        .dout(new_Jinkela_wire_7462)
    );

    bfr new_Jinkela_buffer_5766 (
        .din(new_Jinkela_wire_7355),
        .dout(new_Jinkela_wire_7356)
    );

    bfr new_Jinkela_buffer_5972 (
        .din(_0514_),
        .dout(new_Jinkela_wire_7582)
    );

    bfr new_Jinkela_buffer_5767 (
        .din(new_Jinkela_wire_7356),
        .dout(new_Jinkela_wire_7357)
    );

    bfr new_Jinkela_buffer_5865 (
        .din(new_Jinkela_wire_7462),
        .dout(new_Jinkela_wire_7463)
    );

    bfr new_Jinkela_buffer_5768 (
        .din(new_Jinkela_wire_7357),
        .dout(new_Jinkela_wire_7358)
    );

    bfr new_Jinkela_buffer_5907 (
        .din(new_Jinkela_wire_7510),
        .dout(new_Jinkela_wire_7511)
    );

    bfr new_Jinkela_buffer_5769 (
        .din(new_Jinkela_wire_7358),
        .dout(new_Jinkela_wire_7359)
    );

    bfr new_Jinkela_buffer_5866 (
        .din(new_Jinkela_wire_7463),
        .dout(new_Jinkela_wire_7464)
    );

    bfr new_Jinkela_buffer_5770 (
        .din(new_Jinkela_wire_7359),
        .dout(new_Jinkela_wire_7360)
    );

    bfr new_Jinkela_buffer_5909 (
        .din(new_Jinkela_wire_7516),
        .dout(new_Jinkela_wire_7517)
    );

    bfr new_Jinkela_buffer_5771 (
        .din(new_Jinkela_wire_7360),
        .dout(new_Jinkela_wire_7361)
    );

    bfr new_Jinkela_buffer_5867 (
        .din(new_Jinkela_wire_7464),
        .dout(new_Jinkela_wire_7465)
    );

    bfr new_Jinkela_buffer_5772 (
        .din(new_Jinkela_wire_7361),
        .dout(new_Jinkela_wire_7362)
    );

    spl2 new_Jinkela_splitter_654 (
        .a(_1115_),
        .b(new_Jinkela_wire_7584),
        .c(new_Jinkela_wire_7585)
    );

    bfr new_Jinkela_buffer_5773 (
        .din(new_Jinkela_wire_7362),
        .dout(new_Jinkela_wire_7363)
    );

    bfr new_Jinkela_buffer_5868 (
        .din(new_Jinkela_wire_7465),
        .dout(new_Jinkela_wire_7466)
    );

    bfr new_Jinkela_buffer_5774 (
        .din(new_Jinkela_wire_7363),
        .dout(new_Jinkela_wire_7364)
    );

    bfr new_Jinkela_buffer_5910 (
        .din(new_Jinkela_wire_7517),
        .dout(new_Jinkela_wire_7518)
    );

    bfr new_Jinkela_buffer_5775 (
        .din(new_Jinkela_wire_7364),
        .dout(new_Jinkela_wire_7365)
    );

    bfr new_Jinkela_buffer_5869 (
        .din(new_Jinkela_wire_7466),
        .dout(new_Jinkela_wire_7467)
    );

    bfr new_Jinkela_buffer_5776 (
        .din(new_Jinkela_wire_7365),
        .dout(new_Jinkela_wire_7366)
    );

    spl2 new_Jinkela_splitter_655 (
        .a(_0780_),
        .b(new_Jinkela_wire_7586),
        .c(new_Jinkela_wire_7587)
    );

    bfr new_Jinkela_buffer_5777 (
        .din(new_Jinkela_wire_7366),
        .dout(new_Jinkela_wire_7367)
    );

    bfr new_Jinkela_buffer_5870 (
        .din(new_Jinkela_wire_7467),
        .dout(new_Jinkela_wire_7468)
    );

    bfr new_Jinkela_buffer_5778 (
        .din(new_Jinkela_wire_7367),
        .dout(new_Jinkela_wire_7368)
    );

    bfr new_Jinkela_buffer_5911 (
        .din(new_Jinkela_wire_7518),
        .dout(new_Jinkela_wire_7519)
    );

    bfr new_Jinkela_buffer_5779 (
        .din(new_Jinkela_wire_7368),
        .dout(new_Jinkela_wire_7369)
    );

    bfr new_Jinkela_buffer_5871 (
        .din(new_Jinkela_wire_7468),
        .dout(new_Jinkela_wire_7469)
    );

    bfr new_Jinkela_buffer_5780 (
        .din(new_Jinkela_wire_7369),
        .dout(new_Jinkela_wire_7370)
    );

    bfr new_Jinkela_buffer_5974 (
        .din(_1552_),
        .dout(new_Jinkela_wire_7588)
    );

    bfr new_Jinkela_buffer_5781 (
        .din(new_Jinkela_wire_7370),
        .dout(new_Jinkela_wire_7371)
    );

    bfr new_Jinkela_buffer_5872 (
        .din(new_Jinkela_wire_7469),
        .dout(new_Jinkela_wire_7470)
    );

    bfr new_Jinkela_buffer_12882 (
        .din(new_Jinkela_wire_15403),
        .dout(new_Jinkela_wire_15404)
    );

    bfr new_Jinkela_buffer_16129 (
        .din(new_Jinkela_wire_19253),
        .dout(new_Jinkela_wire_19254)
    );

    bfr new_Jinkela_buffer_12720 (
        .din(new_Jinkela_wire_15241),
        .dout(new_Jinkela_wire_15242)
    );

    spl2 new_Jinkela_splitter_1431 (
        .a(_0847_),
        .b(new_Jinkela_wire_19468),
        .c(new_Jinkela_wire_19469)
    );

    bfr new_Jinkela_buffer_16130 (
        .din(new_Jinkela_wire_19254),
        .dout(new_Jinkela_wire_19255)
    );

    bfr new_Jinkela_buffer_12721 (
        .din(new_Jinkela_wire_15242),
        .dout(new_Jinkela_wire_15243)
    );

    bfr new_Jinkela_buffer_12950 (
        .din(new_Jinkela_wire_15473),
        .dout(new_Jinkela_wire_15474)
    );

    bfr new_Jinkela_buffer_16230 (
        .din(_1569_),
        .dout(new_Jinkela_wire_19393)
    );

    bfr new_Jinkela_buffer_12883 (
        .din(new_Jinkela_wire_15404),
        .dout(new_Jinkela_wire_15405)
    );

    bfr new_Jinkela_buffer_16131 (
        .din(new_Jinkela_wire_19255),
        .dout(new_Jinkela_wire_19256)
    );

    bfr new_Jinkela_buffer_12722 (
        .din(new_Jinkela_wire_15243),
        .dout(new_Jinkela_wire_15244)
    );

    bfr new_Jinkela_buffer_16193 (
        .din(new_Jinkela_wire_19353),
        .dout(new_Jinkela_wire_19354)
    );

    bfr new_Jinkela_buffer_16132 (
        .din(new_Jinkela_wire_19256),
        .dout(new_Jinkela_wire_19257)
    );

    bfr new_Jinkela_buffer_12723 (
        .din(new_Jinkela_wire_15244),
        .dout(new_Jinkela_wire_15245)
    );

    bfr new_Jinkela_buffer_13021 (
        .din(_0686_),
        .dout(new_Jinkela_wire_15553)
    );

    bfr new_Jinkela_buffer_16307 (
        .din(_1827_),
        .dout(new_Jinkela_wire_19474)
    );

    bfr new_Jinkela_buffer_12884 (
        .din(new_Jinkela_wire_15405),
        .dout(new_Jinkela_wire_15406)
    );

    bfr new_Jinkela_buffer_16133 (
        .din(new_Jinkela_wire_19257),
        .dout(new_Jinkela_wire_19258)
    );

    bfr new_Jinkela_buffer_12724 (
        .din(new_Jinkela_wire_15245),
        .dout(new_Jinkela_wire_15246)
    );

    bfr new_Jinkela_buffer_16194 (
        .din(new_Jinkela_wire_19354),
        .dout(new_Jinkela_wire_19355)
    );

    bfr new_Jinkela_buffer_16134 (
        .din(new_Jinkela_wire_19258),
        .dout(new_Jinkela_wire_19259)
    );

    bfr new_Jinkela_buffer_12725 (
        .din(new_Jinkela_wire_15246),
        .dout(new_Jinkela_wire_15247)
    );

    bfr new_Jinkela_buffer_16231 (
        .din(new_Jinkela_wire_19393),
        .dout(new_Jinkela_wire_19394)
    );

    bfr new_Jinkela_buffer_12951 (
        .din(new_Jinkela_wire_15474),
        .dout(new_Jinkela_wire_15475)
    );

    bfr new_Jinkela_buffer_12885 (
        .din(new_Jinkela_wire_15406),
        .dout(new_Jinkela_wire_15407)
    );

    bfr new_Jinkela_buffer_16135 (
        .din(new_Jinkela_wire_19259),
        .dout(new_Jinkela_wire_19260)
    );

    bfr new_Jinkela_buffer_12726 (
        .din(new_Jinkela_wire_15247),
        .dout(new_Jinkela_wire_15248)
    );

    bfr new_Jinkela_buffer_16195 (
        .din(new_Jinkela_wire_19355),
        .dout(new_Jinkela_wire_19356)
    );

    bfr new_Jinkela_buffer_16136 (
        .din(new_Jinkela_wire_19260),
        .dout(new_Jinkela_wire_19261)
    );

    bfr new_Jinkela_buffer_12727 (
        .din(new_Jinkela_wire_15248),
        .dout(new_Jinkela_wire_15249)
    );

    spl2 new_Jinkela_splitter_1115 (
        .a(_1625_),
        .b(new_Jinkela_wire_15554),
        .c(new_Jinkela_wire_15555)
    );

    bfr new_Jinkela_buffer_12886 (
        .din(new_Jinkela_wire_15407),
        .dout(new_Jinkela_wire_15408)
    );

    bfr new_Jinkela_buffer_16137 (
        .din(new_Jinkela_wire_19261),
        .dout(new_Jinkela_wire_19262)
    );

    bfr new_Jinkela_buffer_12728 (
        .din(new_Jinkela_wire_15249),
        .dout(new_Jinkela_wire_15250)
    );

    bfr new_Jinkela_buffer_16196 (
        .din(new_Jinkela_wire_19356),
        .dout(new_Jinkela_wire_19357)
    );

    bfr new_Jinkela_buffer_12994 (
        .din(new_Jinkela_wire_15523),
        .dout(new_Jinkela_wire_15524)
    );

    bfr new_Jinkela_buffer_16138 (
        .din(new_Jinkela_wire_19262),
        .dout(new_Jinkela_wire_19263)
    );

    bfr new_Jinkela_buffer_12729 (
        .din(new_Jinkela_wire_15250),
        .dout(new_Jinkela_wire_15251)
    );

    bfr new_Jinkela_buffer_16232 (
        .din(new_Jinkela_wire_19394),
        .dout(new_Jinkela_wire_19395)
    );

    bfr new_Jinkela_buffer_12952 (
        .din(new_Jinkela_wire_15475),
        .dout(new_Jinkela_wire_15476)
    );

    bfr new_Jinkela_buffer_12887 (
        .din(new_Jinkela_wire_15408),
        .dout(new_Jinkela_wire_15409)
    );

    bfr new_Jinkela_buffer_16139 (
        .din(new_Jinkela_wire_19263),
        .dout(new_Jinkela_wire_19264)
    );

    bfr new_Jinkela_buffer_12730 (
        .din(new_Jinkela_wire_15251),
        .dout(new_Jinkela_wire_15252)
    );

    bfr new_Jinkela_buffer_16197 (
        .din(new_Jinkela_wire_19357),
        .dout(new_Jinkela_wire_19358)
    );

    bfr new_Jinkela_buffer_16140 (
        .din(new_Jinkela_wire_19264),
        .dout(new_Jinkela_wire_19265)
    );

    bfr new_Jinkela_buffer_12731 (
        .din(new_Jinkela_wire_15252),
        .dout(new_Jinkela_wire_15253)
    );

    bfr new_Jinkela_buffer_16303 (
        .din(new_Jinkela_wire_19469),
        .dout(new_Jinkela_wire_19470)
    );

    spl2 new_Jinkela_splitter_1433 (
        .a(_1479_),
        .b(new_Jinkela_wire_19540),
        .c(new_Jinkela_wire_19541)
    );

    bfr new_Jinkela_buffer_12888 (
        .din(new_Jinkela_wire_15409),
        .dout(new_Jinkela_wire_15410)
    );

    bfr new_Jinkela_buffer_16141 (
        .din(new_Jinkela_wire_19265),
        .dout(new_Jinkela_wire_19266)
    );

    bfr new_Jinkela_buffer_12732 (
        .din(new_Jinkela_wire_15253),
        .dout(new_Jinkela_wire_15254)
    );

    bfr new_Jinkela_buffer_16198 (
        .din(new_Jinkela_wire_19358),
        .dout(new_Jinkela_wire_19359)
    );

    bfr new_Jinkela_buffer_12998 (
        .din(new_Jinkela_wire_15527),
        .dout(new_Jinkela_wire_15528)
    );

    bfr new_Jinkela_buffer_16142 (
        .din(new_Jinkela_wire_19266),
        .dout(new_Jinkela_wire_19267)
    );

    bfr new_Jinkela_buffer_12733 (
        .din(new_Jinkela_wire_15254),
        .dout(new_Jinkela_wire_15255)
    );

    bfr new_Jinkela_buffer_16233 (
        .din(new_Jinkela_wire_19395),
        .dout(new_Jinkela_wire_19396)
    );

    bfr new_Jinkela_buffer_12953 (
        .din(new_Jinkela_wire_15476),
        .dout(new_Jinkela_wire_15477)
    );

    bfr new_Jinkela_buffer_12889 (
        .din(new_Jinkela_wire_15410),
        .dout(new_Jinkela_wire_15411)
    );

    bfr new_Jinkela_buffer_16143 (
        .din(new_Jinkela_wire_19267),
        .dout(new_Jinkela_wire_19268)
    );

    bfr new_Jinkela_buffer_12734 (
        .din(new_Jinkela_wire_15255),
        .dout(new_Jinkela_wire_15256)
    );

    bfr new_Jinkela_buffer_16199 (
        .din(new_Jinkela_wire_19359),
        .dout(new_Jinkela_wire_19360)
    );

    bfr new_Jinkela_buffer_16144 (
        .din(new_Jinkela_wire_19268),
        .dout(new_Jinkela_wire_19269)
    );

    bfr new_Jinkela_buffer_12735 (
        .din(new_Jinkela_wire_15256),
        .dout(new_Jinkela_wire_15257)
    );

    spl2 new_Jinkela_splitter_1434 (
        .a(_0491_),
        .b(new_Jinkela_wire_19542),
        .c(new_Jinkela_wire_19543)
    );

    bfr new_Jinkela_buffer_12890 (
        .din(new_Jinkela_wire_15411),
        .dout(new_Jinkela_wire_15412)
    );

    bfr new_Jinkela_buffer_16145 (
        .din(new_Jinkela_wire_19269),
        .dout(new_Jinkela_wire_19270)
    );

    bfr new_Jinkela_buffer_12736 (
        .din(new_Jinkela_wire_15257),
        .dout(new_Jinkela_wire_15258)
    );

    bfr new_Jinkela_buffer_16200 (
        .din(new_Jinkela_wire_19360),
        .dout(new_Jinkela_wire_19361)
    );

    bfr new_Jinkela_buffer_12995 (
        .din(new_Jinkela_wire_15524),
        .dout(new_Jinkela_wire_15525)
    );

    bfr new_Jinkela_buffer_16146 (
        .din(new_Jinkela_wire_19270),
        .dout(new_Jinkela_wire_19271)
    );

    bfr new_Jinkela_buffer_12737 (
        .din(new_Jinkela_wire_15258),
        .dout(new_Jinkela_wire_15259)
    );

    bfr new_Jinkela_buffer_16234 (
        .din(new_Jinkela_wire_19396),
        .dout(new_Jinkela_wire_19397)
    );

    bfr new_Jinkela_buffer_12954 (
        .din(new_Jinkela_wire_15477),
        .dout(new_Jinkela_wire_15478)
    );

    bfr new_Jinkela_buffer_12891 (
        .din(new_Jinkela_wire_15412),
        .dout(new_Jinkela_wire_15413)
    );

    spl2 new_Jinkela_splitter_1411 (
        .a(new_Jinkela_wire_19271),
        .b(new_Jinkela_wire_19272),
        .c(new_Jinkela_wire_19273)
    );

    bfr new_Jinkela_buffer_12738 (
        .din(new_Jinkela_wire_15259),
        .dout(new_Jinkela_wire_15260)
    );

    bfr new_Jinkela_buffer_16304 (
        .din(new_Jinkela_wire_19470),
        .dout(new_Jinkela_wire_19471)
    );

    bfr new_Jinkela_buffer_16201 (
        .din(new_Jinkela_wire_19361),
        .dout(new_Jinkela_wire_19362)
    );

    bfr new_Jinkela_buffer_12739 (
        .din(new_Jinkela_wire_15260),
        .dout(new_Jinkela_wire_15261)
    );

    bfr new_Jinkela_buffer_16202 (
        .din(new_Jinkela_wire_19362),
        .dout(new_Jinkela_wire_19363)
    );

    bfr new_Jinkela_buffer_16235 (
        .din(new_Jinkela_wire_19397),
        .dout(new_Jinkela_wire_19398)
    );

    bfr new_Jinkela_buffer_12892 (
        .din(new_Jinkela_wire_15413),
        .dout(new_Jinkela_wire_15414)
    );

    bfr new_Jinkela_buffer_12740 (
        .din(new_Jinkela_wire_15261),
        .dout(new_Jinkela_wire_15262)
    );

    bfr new_Jinkela_buffer_16203 (
        .din(new_Jinkela_wire_19363),
        .dout(new_Jinkela_wire_19364)
    );

    bfr new_Jinkela_buffer_9340 (
        .din(new_Jinkela_wire_11369),
        .dout(new_Jinkela_wire_11370)
    );

    bfr new_Jinkela_buffer_9259 (
        .din(new_Jinkela_wire_11282),
        .dout(new_Jinkela_wire_11283)
    );

    bfr new_Jinkela_buffer_9368 (
        .din(_0897_),
        .dout(new_Jinkela_wire_11428)
    );

    bfr new_Jinkela_buffer_9260 (
        .din(new_Jinkela_wire_11283),
        .dout(new_Jinkela_wire_11284)
    );

    bfr new_Jinkela_buffer_9341 (
        .din(new_Jinkela_wire_11370),
        .dout(new_Jinkela_wire_11371)
    );

    bfr new_Jinkela_buffer_9261 (
        .din(new_Jinkela_wire_11284),
        .dout(new_Jinkela_wire_11285)
    );

    bfr new_Jinkela_buffer_9262 (
        .din(new_Jinkela_wire_11285),
        .dout(new_Jinkela_wire_11286)
    );

    bfr new_Jinkela_buffer_9342 (
        .din(new_Jinkela_wire_11371),
        .dout(new_Jinkela_wire_11372)
    );

    bfr new_Jinkela_buffer_9263 (
        .din(new_Jinkela_wire_11286),
        .dout(new_Jinkela_wire_11287)
    );

    bfr new_Jinkela_buffer_9361 (
        .din(new_Jinkela_wire_11418),
        .dout(new_Jinkela_wire_11419)
    );

    bfr new_Jinkela_buffer_9264 (
        .din(new_Jinkela_wire_11287),
        .dout(new_Jinkela_wire_11288)
    );

    bfr new_Jinkela_buffer_9343 (
        .din(new_Jinkela_wire_11372),
        .dout(new_Jinkela_wire_11373)
    );

    bfr new_Jinkela_buffer_9265 (
        .din(new_Jinkela_wire_11288),
        .dout(new_Jinkela_wire_11289)
    );

    bfr new_Jinkela_buffer_9364 (
        .din(new_Jinkela_wire_11423),
        .dout(new_Jinkela_wire_11424)
    );

    spl2 new_Jinkela_splitter_880 (
        .a(_1314_),
        .b(new_Jinkela_wire_11434),
        .c(new_Jinkela_wire_11435)
    );

    bfr new_Jinkela_buffer_9266 (
        .din(new_Jinkela_wire_11289),
        .dout(new_Jinkela_wire_11290)
    );

    bfr new_Jinkela_buffer_9344 (
        .din(new_Jinkela_wire_11373),
        .dout(new_Jinkela_wire_11374)
    );

    bfr new_Jinkela_buffer_9267 (
        .din(new_Jinkela_wire_11290),
        .dout(new_Jinkela_wire_11291)
    );

    bfr new_Jinkela_buffer_9362 (
        .din(new_Jinkela_wire_11419),
        .dout(new_Jinkela_wire_11420)
    );

    bfr new_Jinkela_buffer_9268 (
        .din(new_Jinkela_wire_11291),
        .dout(new_Jinkela_wire_11292)
    );

    bfr new_Jinkela_buffer_9345 (
        .din(new_Jinkela_wire_11374),
        .dout(new_Jinkela_wire_11375)
    );

    bfr new_Jinkela_buffer_9269 (
        .din(new_Jinkela_wire_11292),
        .dout(new_Jinkela_wire_11293)
    );

    spl2 new_Jinkela_splitter_881 (
        .a(_1272_),
        .b(new_Jinkela_wire_11440),
        .c(new_Jinkela_wire_11441)
    );

    bfr new_Jinkela_buffer_9270 (
        .din(new_Jinkela_wire_11293),
        .dout(new_Jinkela_wire_11294)
    );

    bfr new_Jinkela_buffer_9346 (
        .din(new_Jinkela_wire_11375),
        .dout(new_Jinkela_wire_11376)
    );

    bfr new_Jinkela_buffer_9271 (
        .din(new_Jinkela_wire_11294),
        .dout(new_Jinkela_wire_11295)
    );

    bfr new_Jinkela_buffer_9363 (
        .din(new_Jinkela_wire_11420),
        .dout(new_Jinkela_wire_11421)
    );

    bfr new_Jinkela_buffer_9272 (
        .din(new_Jinkela_wire_11295),
        .dout(new_Jinkela_wire_11296)
    );

    bfr new_Jinkela_buffer_9347 (
        .din(new_Jinkela_wire_11376),
        .dout(new_Jinkela_wire_11377)
    );

    bfr new_Jinkela_buffer_9273 (
        .din(new_Jinkela_wire_11296),
        .dout(new_Jinkela_wire_11297)
    );

    bfr new_Jinkela_buffer_9365 (
        .din(new_Jinkela_wire_11424),
        .dout(new_Jinkela_wire_11425)
    );

    bfr new_Jinkela_buffer_9274 (
        .din(new_Jinkela_wire_11297),
        .dout(new_Jinkela_wire_11298)
    );

    bfr new_Jinkela_buffer_9348 (
        .din(new_Jinkela_wire_11377),
        .dout(new_Jinkela_wire_11378)
    );

    bfr new_Jinkela_buffer_9275 (
        .din(new_Jinkela_wire_11298),
        .dout(new_Jinkela_wire_11299)
    );

    bfr new_Jinkela_buffer_9369 (
        .din(new_Jinkela_wire_11428),
        .dout(new_Jinkela_wire_11429)
    );

    bfr new_Jinkela_buffer_9276 (
        .din(new_Jinkela_wire_11299),
        .dout(new_Jinkela_wire_11300)
    );

    bfr new_Jinkela_buffer_9349 (
        .din(new_Jinkela_wire_11378),
        .dout(new_Jinkela_wire_11379)
    );

    bfr new_Jinkela_buffer_9277 (
        .din(new_Jinkela_wire_11300),
        .dout(new_Jinkela_wire_11301)
    );

    bfr new_Jinkela_buffer_9366 (
        .din(new_Jinkela_wire_11425),
        .dout(new_Jinkela_wire_11426)
    );

    bfr new_Jinkela_buffer_9278 (
        .din(new_Jinkela_wire_11301),
        .dout(new_Jinkela_wire_11302)
    );

    bfr new_Jinkela_buffer_9350 (
        .din(new_Jinkela_wire_11379),
        .dout(new_Jinkela_wire_11380)
    );

    bfr new_Jinkela_buffer_9279 (
        .din(new_Jinkela_wire_11302),
        .dout(new_Jinkela_wire_11303)
    );

    and_ii _3256_ (
        .a(new_Jinkela_wire_4676),
        .b(new_Jinkela_wire_18578),
        .c(_0528_)
    );

    bfr new_Jinkela_buffer_5782 (
        .din(new_Jinkela_wire_7371),
        .dout(new_Jinkela_wire_7372)
    );

    and_bb _3257_ (
        .a(new_Jinkela_wire_371),
        .b(new_Jinkela_wire_679),
        .c(_0529_)
    );

    bfr new_Jinkela_buffer_5912 (
        .din(new_Jinkela_wire_7519),
        .dout(new_Jinkela_wire_7520)
    );

    and_ii _3258_ (
        .a(new_Jinkela_wire_2961),
        .b(new_Jinkela_wire_13989),
        .c(_0530_)
    );

    bfr new_Jinkela_buffer_5783 (
        .din(new_Jinkela_wire_7372),
        .dout(new_Jinkela_wire_7373)
    );

    and_bb _3259_ (
        .a(new_Jinkela_wire_693),
        .b(new_Jinkela_wire_520),
        .c(_0531_)
    );

    bfr new_Jinkela_buffer_5873 (
        .din(new_Jinkela_wire_7470),
        .dout(new_Jinkela_wire_7471)
    );

    and_ii _3260_ (
        .a(new_Jinkela_wire_15684),
        .b(new_Jinkela_wire_9563),
        .c(_0532_)
    );

    bfr new_Jinkela_buffer_5784 (
        .din(new_Jinkela_wire_7373),
        .dout(new_Jinkela_wire_7374)
    );

    and_bb _3261_ (
        .a(new_Jinkela_wire_147),
        .b(new_Jinkela_wire_491),
        .c(_0533_)
    );

    bfr new_Jinkela_buffer_5975 (
        .din(_0963_),
        .dout(new_Jinkela_wire_7591)
    );

    and_ii _3262_ (
        .a(new_Jinkela_wire_14215),
        .b(new_Jinkela_wire_12722),
        .c(_0534_)
    );

    bfr new_Jinkela_buffer_5785 (
        .din(new_Jinkela_wire_7374),
        .dout(new_Jinkela_wire_7375)
    );

    and_bb _3263_ (
        .a(new_Jinkela_wire_26),
        .b(new_Jinkela_wire_216),
        .c(_0536_)
    );

    bfr new_Jinkela_buffer_5874 (
        .din(new_Jinkela_wire_7471),
        .dout(new_Jinkela_wire_7472)
    );

    and_ii _3264_ (
        .a(new_Jinkela_wire_19543),
        .b(new_Jinkela_wire_18116),
        .c(_0537_)
    );

    bfr new_Jinkela_buffer_5786 (
        .din(new_Jinkela_wire_7375),
        .dout(new_Jinkela_wire_7376)
    );

    and_bb _3265_ (
        .a(new_Jinkela_wire_190),
        .b(new_Jinkela_wire_578),
        .c(_0538_)
    );

    bfr new_Jinkela_buffer_5913 (
        .din(new_Jinkela_wire_7520),
        .dout(new_Jinkela_wire_7521)
    );

    and_ii _3266_ (
        .a(new_Jinkela_wire_4712),
        .b(new_Jinkela_wire_16966),
        .c(_0539_)
    );

    bfr new_Jinkela_buffer_5787 (
        .din(new_Jinkela_wire_7376),
        .dout(new_Jinkela_wire_7377)
    );

    and_bb _3267_ (
        .a(new_Jinkela_wire_386),
        .b(new_Jinkela_wire_127),
        .c(_0540_)
    );

    bfr new_Jinkela_buffer_5875 (
        .din(new_Jinkela_wire_7472),
        .dout(new_Jinkela_wire_7473)
    );

    and_ii _3268_ (
        .a(new_Jinkela_wire_20270),
        .b(new_Jinkela_wire_20967),
        .c(_0541_)
    );

    bfr new_Jinkela_buffer_5788 (
        .din(new_Jinkela_wire_7377),
        .dout(new_Jinkela_wire_7378)
    );

    and_bb _3269_ (
        .a(new_Jinkela_wire_406),
        .b(new_Jinkela_wire_16),
        .c(_0542_)
    );

    spl2 new_Jinkela_splitter_656 (
        .a(_0217_),
        .b(new_Jinkela_wire_7589),
        .c(new_Jinkela_wire_7590)
    );

    and_ii _3270_ (
        .a(new_Jinkela_wire_3259),
        .b(new_Jinkela_wire_11349),
        .c(_0543_)
    );

    bfr new_Jinkela_buffer_5789 (
        .din(new_Jinkela_wire_7378),
        .dout(new_Jinkela_wire_7379)
    );

    and_bb _3271_ (
        .a(new_Jinkela_wire_166),
        .b(new_Jinkela_wire_456),
        .c(_0544_)
    );

    bfr new_Jinkela_buffer_5876 (
        .din(new_Jinkela_wire_7473),
        .dout(new_Jinkela_wire_7474)
    );

    and_ii _3272_ (
        .a(new_Jinkela_wire_14688),
        .b(new_Jinkela_wire_17322),
        .c(_0545_)
    );

    bfr new_Jinkela_buffer_5790 (
        .din(new_Jinkela_wire_7379),
        .dout(new_Jinkela_wire_7380)
    );

    and_bb _3273_ (
        .a(new_Jinkela_wire_606),
        .b(new_Jinkela_wire_263),
        .c(_0547_)
    );

    bfr new_Jinkela_buffer_5914 (
        .din(new_Jinkela_wire_7521),
        .dout(new_Jinkela_wire_7522)
    );

    and_bb _3274_ (
        .a(new_Jinkela_wire_434),
        .b(new_Jinkela_wire_300),
        .c(_0548_)
    );

    bfr new_Jinkela_buffer_5791 (
        .din(new_Jinkela_wire_7380),
        .dout(new_Jinkela_wire_7381)
    );

    and_ii _3275_ (
        .a(new_Jinkela_wire_20358),
        .b(new_Jinkela_wire_1802),
        .c(_0549_)
    );

    bfr new_Jinkela_buffer_5877 (
        .din(new_Jinkela_wire_7474),
        .dout(new_Jinkela_wire_7475)
    );

    and_ii _3276_ (
        .a(new_Jinkela_wire_12729),
        .b(new_Jinkela_wire_20258),
        .c(_0550_)
    );

    bfr new_Jinkela_buffer_5792 (
        .din(new_Jinkela_wire_7381),
        .dout(new_Jinkela_wire_7382)
    );

    and_bb _3277_ (
        .a(new_Jinkela_wire_12730),
        .b(new_Jinkela_wire_20259),
        .c(_0551_)
    );

    spl2 new_Jinkela_splitter_659 (
        .a(_1475_),
        .b(new_Jinkela_wire_7693),
        .c(new_Jinkela_wire_7694)
    );

    or_bb _3278_ (
        .a(new_Jinkela_wire_5803),
        .b(new_Jinkela_wire_14301),
        .c(_0552_)
    );

    bfr new_Jinkela_buffer_5793 (
        .din(new_Jinkela_wire_7382),
        .dout(new_Jinkela_wire_7383)
    );

    and_ii _3279_ (
        .a(new_Jinkela_wire_7296),
        .b(new_Jinkela_wire_18492),
        .c(_0553_)
    );

    bfr new_Jinkela_buffer_5878 (
        .din(new_Jinkela_wire_7475),
        .dout(new_Jinkela_wire_7476)
    );

    and_bb _3280_ (
        .a(new_Jinkela_wire_7297),
        .b(new_Jinkela_wire_18493),
        .c(_0554_)
    );

    bfr new_Jinkela_buffer_5794 (
        .din(new_Jinkela_wire_7383),
        .dout(new_Jinkela_wire_7384)
    );

    or_bb _3281_ (
        .a(new_Jinkela_wire_10204),
        .b(new_Jinkela_wire_15517),
        .c(_0555_)
    );

    bfr new_Jinkela_buffer_5915 (
        .din(new_Jinkela_wire_7522),
        .dout(new_Jinkela_wire_7523)
    );

    and_ii _3282_ (
        .a(new_Jinkela_wire_1786),
        .b(new_Jinkela_wire_5665),
        .c(_0556_)
    );

    bfr new_Jinkela_buffer_5795 (
        .din(new_Jinkela_wire_7384),
        .dout(new_Jinkela_wire_7385)
    );

    and_bb _3283_ (
        .a(new_Jinkela_wire_1787),
        .b(new_Jinkela_wire_5666),
        .c(_0558_)
    );

    bfr new_Jinkela_buffer_5879 (
        .din(new_Jinkela_wire_7476),
        .dout(new_Jinkela_wire_7477)
    );

    or_bb _3284_ (
        .a(new_Jinkela_wire_13957),
        .b(new_Jinkela_wire_5448),
        .c(_0559_)
    );

    bfr new_Jinkela_buffer_5796 (
        .din(new_Jinkela_wire_7385),
        .dout(new_Jinkela_wire_7386)
    );

    and_ii _3285_ (
        .a(new_Jinkela_wire_3442),
        .b(new_Jinkela_wire_16434),
        .c(_0560_)
    );

    spl2 new_Jinkela_splitter_658 (
        .a(_1121_),
        .b(new_Jinkela_wire_7691),
        .c(new_Jinkela_wire_7692)
    );

    and_bb _3286_ (
        .a(new_Jinkela_wire_3443),
        .b(new_Jinkela_wire_16435),
        .c(_0561_)
    );

    bfr new_Jinkela_buffer_5797 (
        .din(new_Jinkela_wire_7386),
        .dout(new_Jinkela_wire_7387)
    );

    or_bb _3287_ (
        .a(new_Jinkela_wire_18532),
        .b(new_Jinkela_wire_18117),
        .c(_0562_)
    );

    bfr new_Jinkela_buffer_5880 (
        .din(new_Jinkela_wire_7477),
        .dout(new_Jinkela_wire_7478)
    );

    and_ii _3288_ (
        .a(new_Jinkela_wire_4984),
        .b(new_Jinkela_wire_4709),
        .c(_0563_)
    );

    bfr new_Jinkela_buffer_5798 (
        .din(new_Jinkela_wire_7387),
        .dout(new_Jinkela_wire_7388)
    );

    and_bb _3289_ (
        .a(new_Jinkela_wire_4985),
        .b(new_Jinkela_wire_4710),
        .c(_0564_)
    );

    bfr new_Jinkela_buffer_5916 (
        .din(new_Jinkela_wire_7523),
        .dout(new_Jinkela_wire_7524)
    );

    or_bb _3290_ (
        .a(new_Jinkela_wire_840),
        .b(new_Jinkela_wire_16206),
        .c(_0565_)
    );

    bfr new_Jinkela_buffer_5799 (
        .din(new_Jinkela_wire_7388),
        .dout(new_Jinkela_wire_7389)
    );

    and_ii _3291_ (
        .a(new_Jinkela_wire_11393),
        .b(new_Jinkela_wire_5878),
        .c(_0566_)
    );

    bfr new_Jinkela_buffer_5881 (
        .din(new_Jinkela_wire_7478),
        .dout(new_Jinkela_wire_7479)
    );

    and_bb _3292_ (
        .a(new_Jinkela_wire_11394),
        .b(new_Jinkela_wire_5879),
        .c(_0567_)
    );

    bfr new_Jinkela_buffer_5800 (
        .din(new_Jinkela_wire_7389),
        .dout(new_Jinkela_wire_7390)
    );

    or_bb _3293_ (
        .a(new_Jinkela_wire_5990),
        .b(new_Jinkela_wire_2943),
        .c(_0569_)
    );

    bfr new_Jinkela_buffer_5976 (
        .din(new_Jinkela_wire_7591),
        .dout(new_Jinkela_wire_7592)
    );

    and_ii _3294_ (
        .a(new_Jinkela_wire_5158),
        .b(new_Jinkela_wire_6372),
        .c(_0570_)
    );

    bfr new_Jinkela_buffer_5801 (
        .din(new_Jinkela_wire_7390),
        .dout(new_Jinkela_wire_7391)
    );

    and_bb _3295_ (
        .a(new_Jinkela_wire_5159),
        .b(new_Jinkela_wire_6373),
        .c(_0571_)
    );

    bfr new_Jinkela_buffer_5882 (
        .din(new_Jinkela_wire_7479),
        .dout(new_Jinkela_wire_7480)
    );

    or_bb _3296_ (
        .a(new_Jinkela_wire_4462),
        .b(new_Jinkela_wire_6685),
        .c(_0572_)
    );

    bfr new_Jinkela_buffer_5802 (
        .din(new_Jinkela_wire_7391),
        .dout(new_Jinkela_wire_7392)
    );

    and_ii _3297_ (
        .a(new_Jinkela_wire_17989),
        .b(new_Jinkela_wire_9092),
        .c(_0573_)
    );

    bfr new_Jinkela_buffer_5917 (
        .din(new_Jinkela_wire_7524),
        .dout(new_Jinkela_wire_7525)
    );

    bfr new_Jinkela_buffer_13022 (
        .din(_0329_),
        .dout(new_Jinkela_wire_15556)
    );

    bfr new_Jinkela_buffer_12741 (
        .din(new_Jinkela_wire_15262),
        .dout(new_Jinkela_wire_15263)
    );

    bfr new_Jinkela_buffer_12955 (
        .din(new_Jinkela_wire_15478),
        .dout(new_Jinkela_wire_15479)
    );

    bfr new_Jinkela_buffer_12893 (
        .din(new_Jinkela_wire_15414),
        .dout(new_Jinkela_wire_15415)
    );

    bfr new_Jinkela_buffer_12742 (
        .din(new_Jinkela_wire_15263),
        .dout(new_Jinkela_wire_15264)
    );

    bfr new_Jinkela_buffer_12743 (
        .din(new_Jinkela_wire_15264),
        .dout(new_Jinkela_wire_15265)
    );

    spl2 new_Jinkela_splitter_1117 (
        .a(_1103_),
        .b(new_Jinkela_wire_15662),
        .c(new_Jinkela_wire_15663)
    );

    bfr new_Jinkela_buffer_12894 (
        .din(new_Jinkela_wire_15415),
        .dout(new_Jinkela_wire_15416)
    );

    bfr new_Jinkela_buffer_12744 (
        .din(new_Jinkela_wire_15265),
        .dout(new_Jinkela_wire_15266)
    );

    bfr new_Jinkela_buffer_12996 (
        .din(new_Jinkela_wire_15525),
        .dout(new_Jinkela_wire_15526)
    );

    bfr new_Jinkela_buffer_12745 (
        .din(new_Jinkela_wire_15266),
        .dout(new_Jinkela_wire_15267)
    );

    bfr new_Jinkela_buffer_12956 (
        .din(new_Jinkela_wire_15479),
        .dout(new_Jinkela_wire_15480)
    );

    bfr new_Jinkela_buffer_12895 (
        .din(new_Jinkela_wire_15416),
        .dout(new_Jinkela_wire_15417)
    );

    bfr new_Jinkela_buffer_12746 (
        .din(new_Jinkela_wire_15267),
        .dout(new_Jinkela_wire_15268)
    );

    bfr new_Jinkela_buffer_12747 (
        .din(new_Jinkela_wire_15268),
        .dout(new_Jinkela_wire_15269)
    );

    bfr new_Jinkela_buffer_12896 (
        .din(new_Jinkela_wire_15417),
        .dout(new_Jinkela_wire_15418)
    );

    bfr new_Jinkela_buffer_12748 (
        .din(new_Jinkela_wire_15269),
        .dout(new_Jinkela_wire_15270)
    );

    bfr new_Jinkela_buffer_12999 (
        .din(new_Jinkela_wire_15528),
        .dout(new_Jinkela_wire_15529)
    );

    bfr new_Jinkela_buffer_12749 (
        .din(new_Jinkela_wire_15270),
        .dout(new_Jinkela_wire_15271)
    );

    bfr new_Jinkela_buffer_12957 (
        .din(new_Jinkela_wire_15480),
        .dout(new_Jinkela_wire_15481)
    );

    bfr new_Jinkela_buffer_12897 (
        .din(new_Jinkela_wire_15418),
        .dout(new_Jinkela_wire_15419)
    );

    bfr new_Jinkela_buffer_12750 (
        .din(new_Jinkela_wire_15271),
        .dout(new_Jinkela_wire_15272)
    );

    bfr new_Jinkela_buffer_12751 (
        .din(new_Jinkela_wire_15272),
        .dout(new_Jinkela_wire_15273)
    );

    bfr new_Jinkela_buffer_12898 (
        .din(new_Jinkela_wire_15419),
        .dout(new_Jinkela_wire_15420)
    );

    bfr new_Jinkela_buffer_12752 (
        .din(new_Jinkela_wire_15273),
        .dout(new_Jinkela_wire_15274)
    );

    bfr new_Jinkela_buffer_12753 (
        .din(new_Jinkela_wire_15274),
        .dout(new_Jinkela_wire_15275)
    );

    bfr new_Jinkela_buffer_12958 (
        .din(new_Jinkela_wire_15481),
        .dout(new_Jinkela_wire_15482)
    );

    bfr new_Jinkela_buffer_12899 (
        .din(new_Jinkela_wire_15420),
        .dout(new_Jinkela_wire_15421)
    );

    bfr new_Jinkela_buffer_12754 (
        .din(new_Jinkela_wire_15275),
        .dout(new_Jinkela_wire_15276)
    );

    bfr new_Jinkela_buffer_12755 (
        .din(new_Jinkela_wire_15276),
        .dout(new_Jinkela_wire_15277)
    );

    bfr new_Jinkela_buffer_12900 (
        .din(new_Jinkela_wire_15421),
        .dout(new_Jinkela_wire_15422)
    );

    bfr new_Jinkela_buffer_12756 (
        .din(new_Jinkela_wire_15277),
        .dout(new_Jinkela_wire_15278)
    );

    bfr new_Jinkela_buffer_13000 (
        .din(new_Jinkela_wire_15529),
        .dout(new_Jinkela_wire_15530)
    );

    bfr new_Jinkela_buffer_12757 (
        .din(new_Jinkela_wire_15278),
        .dout(new_Jinkela_wire_15279)
    );

    bfr new_Jinkela_buffer_12959 (
        .din(new_Jinkela_wire_15482),
        .dout(new_Jinkela_wire_15483)
    );

    bfr new_Jinkela_buffer_12901 (
        .din(new_Jinkela_wire_15422),
        .dout(new_Jinkela_wire_15423)
    );

    bfr new_Jinkela_buffer_12758 (
        .din(new_Jinkela_wire_15279),
        .dout(new_Jinkela_wire_15280)
    );

    bfr new_Jinkela_buffer_12759 (
        .din(new_Jinkela_wire_15280),
        .dout(new_Jinkela_wire_15281)
    );

    bfr new_Jinkela_buffer_12902 (
        .din(new_Jinkela_wire_15423),
        .dout(new_Jinkela_wire_15424)
    );

    bfr new_Jinkela_buffer_12760 (
        .din(new_Jinkela_wire_15281),
        .dout(new_Jinkela_wire_15282)
    );

    bfr new_Jinkela_buffer_12761 (
        .din(new_Jinkela_wire_15282),
        .dout(new_Jinkela_wire_15283)
    );

    bfr new_Jinkela_buffer_12960 (
        .din(new_Jinkela_wire_15483),
        .dout(new_Jinkela_wire_15484)
    );

    bfr new_Jinkela_buffer_9372 (
        .din(new_Jinkela_wire_11435),
        .dout(new_Jinkela_wire_11436)
    );

    or_ii _2371_ (
        .a(new_Jinkela_wire_14990),
        .b(new_Jinkela_wire_1765),
        .c(_1407_)
    );

    bfr new_Jinkela_buffer_9280 (
        .din(new_Jinkela_wire_11303),
        .dout(new_Jinkela_wire_11304)
    );

    and_ii _2372_ (
        .a(new_Jinkela_wire_9541),
        .b(new_Jinkela_wire_14076),
        .c(_1408_)
    );

    bfr new_Jinkela_buffer_9351 (
        .din(new_Jinkela_wire_11380),
        .dout(new_Jinkela_wire_11381)
    );

    and_bb _2373_ (
        .a(new_Jinkela_wire_9542),
        .b(new_Jinkela_wire_14077),
        .c(_1409_)
    );

    bfr new_Jinkela_buffer_9281 (
        .din(new_Jinkela_wire_11304),
        .dout(new_Jinkela_wire_11305)
    );

    or_bb _2374_ (
        .a(new_Jinkela_wire_8186),
        .b(new_Jinkela_wire_15519),
        .c(_1410_)
    );

    bfr new_Jinkela_buffer_9367 (
        .din(new_Jinkela_wire_11426),
        .dout(new_Jinkela_wire_11427)
    );

    or_bb _2375_ (
        .a(new_Jinkela_wire_9183),
        .b(new_Jinkela_wire_18528),
        .c(_1411_)
    );

    bfr new_Jinkela_buffer_9282 (
        .din(new_Jinkela_wire_11305),
        .dout(new_Jinkela_wire_11306)
    );

    or_ii _2376_ (
        .a(new_Jinkela_wire_9184),
        .b(new_Jinkela_wire_18529),
        .c(_1412_)
    );

    bfr new_Jinkela_buffer_9352 (
        .din(new_Jinkela_wire_11381),
        .dout(new_Jinkela_wire_11382)
    );

    or_ii _2377_ (
        .a(new_Jinkela_wire_18563),
        .b(new_Jinkela_wire_14319),
        .c(_1413_)
    );

    bfr new_Jinkela_buffer_9283 (
        .din(new_Jinkela_wire_11306),
        .dout(new_Jinkela_wire_11307)
    );

    and_ii _2378_ (
        .a(new_Jinkela_wire_19282),
        .b(new_Jinkela_wire_17724),
        .c(_1414_)
    );

    bfr new_Jinkela_buffer_9370 (
        .din(new_Jinkela_wire_11429),
        .dout(new_Jinkela_wire_11430)
    );

    and_bb _2379_ (
        .a(new_Jinkela_wire_19283),
        .b(new_Jinkela_wire_17725),
        .c(_1415_)
    );

    bfr new_Jinkela_buffer_9284 (
        .din(new_Jinkela_wire_11307),
        .dout(new_Jinkela_wire_11308)
    );

    or_bb _2380_ (
        .a(new_Jinkela_wire_13014),
        .b(new_Jinkela_wire_4328),
        .c(_1416_)
    );

    bfr new_Jinkela_buffer_9353 (
        .din(new_Jinkela_wire_11382),
        .dout(new_Jinkela_wire_11383)
    );

    or_bb _2381_ (
        .a(new_Jinkela_wire_7443),
        .b(new_Jinkela_wire_15743),
        .c(_1417_)
    );

    bfr new_Jinkela_buffer_9285 (
        .din(new_Jinkela_wire_11308),
        .dout(new_Jinkela_wire_11309)
    );

    or_ii _2382_ (
        .a(new_Jinkela_wire_7444),
        .b(new_Jinkela_wire_15744),
        .c(_1418_)
    );

    or_ii _2383_ (
        .a(new_Jinkela_wire_20339),
        .b(new_Jinkela_wire_10091),
        .c(_1419_)
    );

    spl2 new_Jinkela_splitter_882 (
        .a(_1585_),
        .b(new_Jinkela_wire_11442),
        .c(new_Jinkela_wire_11443)
    );

    bfr new_Jinkela_buffer_9286 (
        .din(new_Jinkela_wire_11309),
        .dout(new_Jinkela_wire_11310)
    );

    and_ii _2384_ (
        .a(new_Jinkela_wire_19783),
        .b(new_Jinkela_wire_17915),
        .c(_1420_)
    );

    spl2 new_Jinkela_splitter_864 (
        .a(new_Jinkela_wire_11383),
        .b(new_Jinkela_wire_11384),
        .c(new_Jinkela_wire_11385)
    );

    and_bb _2385_ (
        .a(new_Jinkela_wire_19784),
        .b(new_Jinkela_wire_17916),
        .c(_1421_)
    );

    bfr new_Jinkela_buffer_9287 (
        .din(new_Jinkela_wire_11310),
        .dout(new_Jinkela_wire_11311)
    );

    or_bb _2386_ (
        .a(new_Jinkela_wire_3963),
        .b(new_Jinkela_wire_2259),
        .c(_1422_)
    );

    or_bb _2387_ (
        .a(new_Jinkela_wire_4164),
        .b(new_Jinkela_wire_9860),
        .c(_1423_)
    );

    bfr new_Jinkela_buffer_9288 (
        .din(new_Jinkela_wire_11311),
        .dout(new_Jinkela_wire_11312)
    );

    or_ii _2388_ (
        .a(new_Jinkela_wire_4165),
        .b(new_Jinkela_wire_9861),
        .c(_1424_)
    );

    bfr new_Jinkela_buffer_9371 (
        .din(new_Jinkela_wire_11430),
        .dout(new_Jinkela_wire_11431)
    );

    or_ii _2389_ (
        .a(new_Jinkela_wire_13586),
        .b(new_Jinkela_wire_6196),
        .c(_1425_)
    );

    bfr new_Jinkela_buffer_9289 (
        .din(new_Jinkela_wire_11312),
        .dout(new_Jinkela_wire_11313)
    );

    and_ii _2390_ (
        .a(new_Jinkela_wire_5683),
        .b(new_Jinkela_wire_16188),
        .c(_1426_)
    );

    spl2 new_Jinkela_splitter_879 (
        .a(new_Jinkela_wire_11431),
        .b(new_Jinkela_wire_11432),
        .c(new_Jinkela_wire_11433)
    );

    and_bb _2391_ (
        .a(new_Jinkela_wire_5684),
        .b(new_Jinkela_wire_16189),
        .c(_1427_)
    );

    bfr new_Jinkela_buffer_9290 (
        .din(new_Jinkela_wire_11313),
        .dout(new_Jinkela_wire_11314)
    );

    or_bb _2392_ (
        .a(new_Jinkela_wire_13011),
        .b(new_Jinkela_wire_13730),
        .c(_1428_)
    );

    spl2 new_Jinkela_splitter_885 (
        .a(_1628_),
        .b(new_Jinkela_wire_11454),
        .c(new_Jinkela_wire_11455)
    );

    or_bb _2393_ (
        .a(new_Jinkela_wire_16959),
        .b(new_Jinkela_wire_5681),
        .c(_1429_)
    );

    bfr new_Jinkela_buffer_9376 (
        .din(_0842_),
        .dout(new_Jinkela_wire_11444)
    );

    bfr new_Jinkela_buffer_9291 (
        .din(new_Jinkela_wire_11314),
        .dout(new_Jinkela_wire_11315)
    );

    or_ii _2394_ (
        .a(new_Jinkela_wire_16960),
        .b(new_Jinkela_wire_5682),
        .c(_1430_)
    );

    bfr new_Jinkela_buffer_9373 (
        .din(new_Jinkela_wire_11436),
        .dout(new_Jinkela_wire_11437)
    );

    or_ii _2395_ (
        .a(new_Jinkela_wire_2018),
        .b(new_Jinkela_wire_21208),
        .c(_1431_)
    );

    bfr new_Jinkela_buffer_9292 (
        .din(new_Jinkela_wire_11315),
        .dout(new_Jinkela_wire_11316)
    );

    and_ii _2396_ (
        .a(new_Jinkela_wire_18697),
        .b(new_Jinkela_wire_11523),
        .c(_1432_)
    );

    bfr new_Jinkela_buffer_9374 (
        .din(new_Jinkela_wire_11437),
        .dout(new_Jinkela_wire_11438)
    );

    and_bb _2397_ (
        .a(new_Jinkela_wire_18698),
        .b(new_Jinkela_wire_11524),
        .c(_1433_)
    );

    bfr new_Jinkela_buffer_9293 (
        .din(new_Jinkela_wire_11316),
        .dout(new_Jinkela_wire_11317)
    );

    or_bb _2398_ (
        .a(new_Jinkela_wire_21167),
        .b(new_Jinkela_wire_5544),
        .c(_1434_)
    );

    bfr new_Jinkela_buffer_9377 (
        .din(_0591_),
        .dout(new_Jinkela_wire_11447)
    );

    or_bb _2399_ (
        .a(new_Jinkela_wire_13400),
        .b(new_Jinkela_wire_18104),
        .c(_1435_)
    );

    spl2 new_Jinkela_splitter_883 (
        .a(_0015_),
        .b(new_Jinkela_wire_11445),
        .c(new_Jinkela_wire_11446)
    );

    bfr new_Jinkela_buffer_9294 (
        .din(new_Jinkela_wire_11317),
        .dout(new_Jinkela_wire_11318)
    );

    or_ii _2400_ (
        .a(new_Jinkela_wire_13401),
        .b(new_Jinkela_wire_18105),
        .c(_1436_)
    );

    bfr new_Jinkela_buffer_9375 (
        .din(new_Jinkela_wire_11438),
        .dout(new_Jinkela_wire_11439)
    );

    or_ii _2401_ (
        .a(new_Jinkela_wire_17797),
        .b(new_Jinkela_wire_19548),
        .c(_1437_)
    );

    bfr new_Jinkela_buffer_9295 (
        .din(new_Jinkela_wire_11318),
        .dout(new_Jinkela_wire_11319)
    );

    and_ii _2402_ (
        .a(new_Jinkela_wire_5723),
        .b(new_Jinkela_wire_11612),
        .c(_1438_)
    );

    bfr new_Jinkela_buffer_9378 (
        .din(new_Jinkela_wire_11449),
        .dout(new_Jinkela_wire_11450)
    );

    and_bb _2403_ (
        .a(new_Jinkela_wire_5724),
        .b(new_Jinkela_wire_11613),
        .c(_1439_)
    );

    bfr new_Jinkela_buffer_9296 (
        .din(new_Jinkela_wire_11319),
        .dout(new_Jinkela_wire_11320)
    );

    or_bb _2404_ (
        .a(new_Jinkela_wire_7269),
        .b(new_Jinkela_wire_17043),
        .c(_1440_)
    );

    or_bb _2405_ (
        .a(new_Jinkela_wire_12735),
        .b(new_Jinkela_wire_9747),
        .c(_1441_)
    );

    spl2 new_Jinkela_splitter_884 (
        .a(_1118_),
        .b(new_Jinkela_wire_11448),
        .c(new_Jinkela_wire_11449)
    );

    bfr new_Jinkela_buffer_9297 (
        .din(new_Jinkela_wire_11320),
        .dout(new_Jinkela_wire_11321)
    );

    or_ii _2406_ (
        .a(new_Jinkela_wire_12736),
        .b(new_Jinkela_wire_9748),
        .c(_1442_)
    );

    or_ii _2407_ (
        .a(new_Jinkela_wire_6738),
        .b(new_Jinkela_wire_9601),
        .c(_1443_)
    );

    bfr new_Jinkela_buffer_9298 (
        .din(new_Jinkela_wire_11321),
        .dout(new_Jinkela_wire_11322)
    );

    and_ii _2408_ (
        .a(new_Jinkela_wire_6519),
        .b(new_Jinkela_wire_12709),
        .c(_1444_)
    );

    and_bb _2409_ (
        .a(new_Jinkela_wire_6520),
        .b(new_Jinkela_wire_12710),
        .c(_1445_)
    );

    spl2 new_Jinkela_splitter_886 (
        .a(_1589_),
        .b(new_Jinkela_wire_11456),
        .c(new_Jinkela_wire_11457)
    );

    bfr new_Jinkela_buffer_9299 (
        .din(new_Jinkela_wire_11322),
        .dout(new_Jinkela_wire_11323)
    );

    or_bb _2410_ (
        .a(new_Jinkela_wire_4293),
        .b(new_Jinkela_wire_14026),
        .c(_1446_)
    );

    bfr new_Jinkela_buffer_9383 (
        .din(_1367_),
        .dout(new_Jinkela_wire_11459)
    );

    or_bb _2411_ (
        .a(new_Jinkela_wire_2312),
        .b(new_Jinkela_wire_13058),
        .c(_1447_)
    );

    bfr new_Jinkela_buffer_9300 (
        .din(new_Jinkela_wire_11323),
        .dout(new_Jinkela_wire_11324)
    );

    and_bb _2412_ (
        .a(new_Jinkela_wire_2313),
        .b(new_Jinkela_wire_13059),
        .c(_1448_)
    );

    bfr new_Jinkela_buffer_5803 (
        .din(new_Jinkela_wire_7392),
        .dout(new_Jinkela_wire_7393)
    );

    bfr new_Jinkela_buffer_5883 (
        .din(new_Jinkela_wire_7480),
        .dout(new_Jinkela_wire_7481)
    );

    bfr new_Jinkela_buffer_5804 (
        .din(new_Jinkela_wire_7393),
        .dout(new_Jinkela_wire_7394)
    );

    bfr new_Jinkela_buffer_6073 (
        .din(new_Jinkela_wire_7696),
        .dout(new_Jinkela_wire_7697)
    );

    bfr new_Jinkela_buffer_5805 (
        .din(new_Jinkela_wire_7394),
        .dout(new_Jinkela_wire_7395)
    );

    bfr new_Jinkela_buffer_5884 (
        .din(new_Jinkela_wire_7481),
        .dout(new_Jinkela_wire_7482)
    );

    bfr new_Jinkela_buffer_5806 (
        .din(new_Jinkela_wire_7395),
        .dout(new_Jinkela_wire_7396)
    );

    bfr new_Jinkela_buffer_5918 (
        .din(new_Jinkela_wire_7525),
        .dout(new_Jinkela_wire_7526)
    );

    bfr new_Jinkela_buffer_5807 (
        .din(new_Jinkela_wire_7396),
        .dout(new_Jinkela_wire_7397)
    );

    bfr new_Jinkela_buffer_5885 (
        .din(new_Jinkela_wire_7482),
        .dout(new_Jinkela_wire_7483)
    );

    bfr new_Jinkela_buffer_5808 (
        .din(new_Jinkela_wire_7397),
        .dout(new_Jinkela_wire_7398)
    );

    bfr new_Jinkela_buffer_5977 (
        .din(new_Jinkela_wire_7592),
        .dout(new_Jinkela_wire_7593)
    );

    bfr new_Jinkela_buffer_5809 (
        .din(new_Jinkela_wire_7398),
        .dout(new_Jinkela_wire_7399)
    );

    bfr new_Jinkela_buffer_5886 (
        .din(new_Jinkela_wire_7483),
        .dout(new_Jinkela_wire_7484)
    );

    bfr new_Jinkela_buffer_5810 (
        .din(new_Jinkela_wire_7399),
        .dout(new_Jinkela_wire_7400)
    );

    bfr new_Jinkela_buffer_5919 (
        .din(new_Jinkela_wire_7526),
        .dout(new_Jinkela_wire_7527)
    );

    bfr new_Jinkela_buffer_5811 (
        .din(new_Jinkela_wire_7400),
        .dout(new_Jinkela_wire_7401)
    );

    bfr new_Jinkela_buffer_5887 (
        .din(new_Jinkela_wire_7484),
        .dout(new_Jinkela_wire_7485)
    );

    bfr new_Jinkela_buffer_5812 (
        .din(new_Jinkela_wire_7401),
        .dout(new_Jinkela_wire_7402)
    );

    spl2 new_Jinkela_splitter_660 (
        .a(_0596_),
        .b(new_Jinkela_wire_7695),
        .c(new_Jinkela_wire_7696)
    );

    bfr new_Jinkela_buffer_5813 (
        .din(new_Jinkela_wire_7402),
        .dout(new_Jinkela_wire_7403)
    );

    bfr new_Jinkela_buffer_5888 (
        .din(new_Jinkela_wire_7485),
        .dout(new_Jinkela_wire_7486)
    );

    bfr new_Jinkela_buffer_5814 (
        .din(new_Jinkela_wire_7403),
        .dout(new_Jinkela_wire_7404)
    );

    bfr new_Jinkela_buffer_5920 (
        .din(new_Jinkela_wire_7527),
        .dout(new_Jinkela_wire_7528)
    );

    bfr new_Jinkela_buffer_5815 (
        .din(new_Jinkela_wire_7404),
        .dout(new_Jinkela_wire_7405)
    );

    bfr new_Jinkela_buffer_5889 (
        .din(new_Jinkela_wire_7486),
        .dout(new_Jinkela_wire_7487)
    );

    bfr new_Jinkela_buffer_5816 (
        .din(new_Jinkela_wire_7405),
        .dout(new_Jinkela_wire_7406)
    );

    bfr new_Jinkela_buffer_5978 (
        .din(new_Jinkela_wire_7593),
        .dout(new_Jinkela_wire_7594)
    );

    bfr new_Jinkela_buffer_5817 (
        .din(new_Jinkela_wire_7406),
        .dout(new_Jinkela_wire_7407)
    );

    bfr new_Jinkela_buffer_5890 (
        .din(new_Jinkela_wire_7487),
        .dout(new_Jinkela_wire_7488)
    );

    bfr new_Jinkela_buffer_5818 (
        .din(new_Jinkela_wire_7407),
        .dout(new_Jinkela_wire_7408)
    );

    bfr new_Jinkela_buffer_5921 (
        .din(new_Jinkela_wire_7528),
        .dout(new_Jinkela_wire_7529)
    );

    bfr new_Jinkela_buffer_5819 (
        .din(new_Jinkela_wire_7408),
        .dout(new_Jinkela_wire_7409)
    );

    bfr new_Jinkela_buffer_5891 (
        .din(new_Jinkela_wire_7488),
        .dout(new_Jinkela_wire_7489)
    );

    bfr new_Jinkela_buffer_5820 (
        .din(new_Jinkela_wire_7409),
        .dout(new_Jinkela_wire_7410)
    );

    spl2 new_Jinkela_splitter_661 (
        .a(_0785_),
        .b(new_Jinkela_wire_7701),
        .c(new_Jinkela_wire_7702)
    );

    bfr new_Jinkela_buffer_5821 (
        .din(new_Jinkela_wire_7410),
        .dout(new_Jinkela_wire_7411)
    );

    bfr new_Jinkela_buffer_5892 (
        .din(new_Jinkela_wire_7489),
        .dout(new_Jinkela_wire_7490)
    );

    bfr new_Jinkela_buffer_5822 (
        .din(new_Jinkela_wire_7411),
        .dout(new_Jinkela_wire_7412)
    );

    bfr new_Jinkela_buffer_5922 (
        .din(new_Jinkela_wire_7529),
        .dout(new_Jinkela_wire_7530)
    );

    bfr new_Jinkela_buffer_5823 (
        .din(new_Jinkela_wire_7412),
        .dout(new_Jinkela_wire_7413)
    );

    bfr new_Jinkela_buffer_5893 (
        .din(new_Jinkela_wire_7490),
        .dout(new_Jinkela_wire_7491)
    );

    bfr new_Jinkela_buffer_2296 (
        .din(new_Jinkela_wire_3283),
        .dout(new_Jinkela_wire_3284)
    );

    bfr new_Jinkela_buffer_2376 (
        .din(new_Jinkela_wire_3367),
        .dout(new_Jinkela_wire_3368)
    );

    bfr new_Jinkela_buffer_2297 (
        .din(new_Jinkela_wire_3284),
        .dout(new_Jinkela_wire_3285)
    );

    spl2 new_Jinkela_splitter_349 (
        .a(_0879_),
        .b(new_Jinkela_wire_3437),
        .c(new_Jinkela_wire_3438)
    );

    bfr new_Jinkela_buffer_2298 (
        .din(new_Jinkela_wire_3285),
        .dout(new_Jinkela_wire_3286)
    );

    bfr new_Jinkela_buffer_2377 (
        .din(new_Jinkela_wire_3368),
        .dout(new_Jinkela_wire_3369)
    );

    bfr new_Jinkela_buffer_2299 (
        .din(new_Jinkela_wire_3286),
        .dout(new_Jinkela_wire_3287)
    );

    bfr new_Jinkela_buffer_2396 (
        .din(new_Jinkela_wire_3389),
        .dout(new_Jinkela_wire_3390)
    );

    bfr new_Jinkela_buffer_2300 (
        .din(new_Jinkela_wire_3287),
        .dout(new_Jinkela_wire_3288)
    );

    bfr new_Jinkela_buffer_2378 (
        .din(new_Jinkela_wire_3369),
        .dout(new_Jinkela_wire_3370)
    );

    bfr new_Jinkela_buffer_2301 (
        .din(new_Jinkela_wire_3288),
        .dout(new_Jinkela_wire_3289)
    );

    bfr new_Jinkela_buffer_2302 (
        .din(new_Jinkela_wire_3289),
        .dout(new_Jinkela_wire_3290)
    );

    bfr new_Jinkela_buffer_2379 (
        .din(new_Jinkela_wire_3370),
        .dout(new_Jinkela_wire_3371)
    );

    bfr new_Jinkela_buffer_2303 (
        .din(new_Jinkela_wire_3290),
        .dout(new_Jinkela_wire_3291)
    );

    bfr new_Jinkela_buffer_2397 (
        .din(new_Jinkela_wire_3390),
        .dout(new_Jinkela_wire_3391)
    );

    bfr new_Jinkela_buffer_2304 (
        .din(new_Jinkela_wire_3291),
        .dout(new_Jinkela_wire_3292)
    );

    bfr new_Jinkela_buffer_2380 (
        .din(new_Jinkela_wire_3371),
        .dout(new_Jinkela_wire_3372)
    );

    bfr new_Jinkela_buffer_2305 (
        .din(new_Jinkela_wire_3292),
        .dout(new_Jinkela_wire_3293)
    );

    bfr new_Jinkela_buffer_2434 (
        .din(new_Jinkela_wire_3431),
        .dout(new_Jinkela_wire_3432)
    );

    bfr new_Jinkela_buffer_2306 (
        .din(new_Jinkela_wire_3293),
        .dout(new_Jinkela_wire_3294)
    );

    bfr new_Jinkela_buffer_2381 (
        .din(new_Jinkela_wire_3372),
        .dout(new_Jinkela_wire_3373)
    );

    bfr new_Jinkela_buffer_2307 (
        .din(new_Jinkela_wire_3294),
        .dout(new_Jinkela_wire_3295)
    );

    bfr new_Jinkela_buffer_2398 (
        .din(new_Jinkela_wire_3391),
        .dout(new_Jinkela_wire_3392)
    );

    bfr new_Jinkela_buffer_2308 (
        .din(new_Jinkela_wire_3295),
        .dout(new_Jinkela_wire_3296)
    );

    bfr new_Jinkela_buffer_2382 (
        .din(new_Jinkela_wire_3373),
        .dout(new_Jinkela_wire_3374)
    );

    bfr new_Jinkela_buffer_2309 (
        .din(new_Jinkela_wire_3296),
        .dout(new_Jinkela_wire_3297)
    );

    bfr new_Jinkela_buffer_2437 (
        .din(_1321_),
        .dout(new_Jinkela_wire_3441)
    );

    spl2 new_Jinkela_splitter_350 (
        .a(_1156_),
        .b(new_Jinkela_wire_3439),
        .c(new_Jinkela_wire_3440)
    );

    bfr new_Jinkela_buffer_2310 (
        .din(new_Jinkela_wire_3297),
        .dout(new_Jinkela_wire_3298)
    );

    bfr new_Jinkela_buffer_2383 (
        .din(new_Jinkela_wire_3374),
        .dout(new_Jinkela_wire_3375)
    );

    bfr new_Jinkela_buffer_2311 (
        .din(new_Jinkela_wire_3298),
        .dout(new_Jinkela_wire_3299)
    );

    bfr new_Jinkela_buffer_2399 (
        .din(new_Jinkela_wire_3392),
        .dout(new_Jinkela_wire_3393)
    );

    bfr new_Jinkela_buffer_2312 (
        .din(new_Jinkela_wire_3299),
        .dout(new_Jinkela_wire_3300)
    );

    bfr new_Jinkela_buffer_2384 (
        .din(new_Jinkela_wire_3375),
        .dout(new_Jinkela_wire_3376)
    );

    bfr new_Jinkela_buffer_2313 (
        .din(new_Jinkela_wire_3300),
        .dout(new_Jinkela_wire_3301)
    );

    bfr new_Jinkela_buffer_2435 (
        .din(new_Jinkela_wire_3432),
        .dout(new_Jinkela_wire_3433)
    );

    bfr new_Jinkela_buffer_2314 (
        .din(new_Jinkela_wire_3301),
        .dout(new_Jinkela_wire_3302)
    );

    bfr new_Jinkela_buffer_2385 (
        .din(new_Jinkela_wire_3376),
        .dout(new_Jinkela_wire_3377)
    );

    bfr new_Jinkela_buffer_2315 (
        .din(new_Jinkela_wire_3302),
        .dout(new_Jinkela_wire_3303)
    );

    bfr new_Jinkela_buffer_2400 (
        .din(new_Jinkela_wire_3393),
        .dout(new_Jinkela_wire_3394)
    );

    bfr new_Jinkela_buffer_2316 (
        .din(new_Jinkela_wire_3303),
        .dout(new_Jinkela_wire_3304)
    );

    bfr new_Jinkela_buffer_2386 (
        .din(new_Jinkela_wire_3377),
        .dout(new_Jinkela_wire_3378)
    );

    bfr new_Jinkela_buffer_2317 (
        .din(new_Jinkela_wire_3304),
        .dout(new_Jinkela_wire_3305)
    );

    bfr new_Jinkela_buffer_9379 (
        .din(new_Jinkela_wire_11450),
        .dout(new_Jinkela_wire_11451)
    );

    bfr new_Jinkela_buffer_12903 (
        .din(new_Jinkela_wire_15424),
        .dout(new_Jinkela_wire_15425)
    );

    bfr new_Jinkela_buffer_12762 (
        .din(new_Jinkela_wire_15283),
        .dout(new_Jinkela_wire_15284)
    );

    spl2 new_Jinkela_splitter_352 (
        .a(_0437_),
        .b(new_Jinkela_wire_3444),
        .c(new_Jinkela_wire_3445)
    );

    bfr new_Jinkela_buffer_9301 (
        .din(new_Jinkela_wire_11324),
        .dout(new_Jinkela_wire_11325)
    );

    bfr new_Jinkela_buffer_2318 (
        .din(new_Jinkela_wire_3305),
        .dout(new_Jinkela_wire_3306)
    );

    bfr new_Jinkela_buffer_9382 (
        .din(new_Jinkela_wire_11457),
        .dout(new_Jinkela_wire_11458)
    );

    bfr new_Jinkela_buffer_12763 (
        .din(new_Jinkela_wire_15284),
        .dout(new_Jinkela_wire_15285)
    );

    bfr new_Jinkela_buffer_2387 (
        .din(new_Jinkela_wire_3378),
        .dout(new_Jinkela_wire_3379)
    );

    bfr new_Jinkela_buffer_9302 (
        .din(new_Jinkela_wire_11325),
        .dout(new_Jinkela_wire_11326)
    );

    spl2 new_Jinkela_splitter_1118 (
        .a(_1797_),
        .b(new_Jinkela_wire_15664),
        .c(new_Jinkela_wire_15665)
    );

    bfr new_Jinkela_buffer_2319 (
        .din(new_Jinkela_wire_3306),
        .dout(new_Jinkela_wire_3307)
    );

    bfr new_Jinkela_buffer_9380 (
        .din(new_Jinkela_wire_11451),
        .dout(new_Jinkela_wire_11452)
    );

    bfr new_Jinkela_buffer_12904 (
        .din(new_Jinkela_wire_15425),
        .dout(new_Jinkela_wire_15426)
    );

    bfr new_Jinkela_buffer_12764 (
        .din(new_Jinkela_wire_15285),
        .dout(new_Jinkela_wire_15286)
    );

    bfr new_Jinkela_buffer_2401 (
        .din(new_Jinkela_wire_3394),
        .dout(new_Jinkela_wire_3395)
    );

    bfr new_Jinkela_buffer_9303 (
        .din(new_Jinkela_wire_11326),
        .dout(new_Jinkela_wire_11327)
    );

    bfr new_Jinkela_buffer_2320 (
        .din(new_Jinkela_wire_3307),
        .dout(new_Jinkela_wire_3308)
    );

    bfr new_Jinkela_buffer_13001 (
        .din(new_Jinkela_wire_15530),
        .dout(new_Jinkela_wire_15531)
    );

    spl2 new_Jinkela_splitter_888 (
        .a(_0022_),
        .b(new_Jinkela_wire_11525),
        .c(new_Jinkela_wire_11526)
    );

    bfr new_Jinkela_buffer_12765 (
        .din(new_Jinkela_wire_15286),
        .dout(new_Jinkela_wire_15287)
    );

    bfr new_Jinkela_buffer_2388 (
        .din(new_Jinkela_wire_3379),
        .dout(new_Jinkela_wire_3380)
    );

    bfr new_Jinkela_buffer_9304 (
        .din(new_Jinkela_wire_11327),
        .dout(new_Jinkela_wire_11328)
    );

    bfr new_Jinkela_buffer_12961 (
        .din(new_Jinkela_wire_15484),
        .dout(new_Jinkela_wire_15485)
    );

    bfr new_Jinkela_buffer_2321 (
        .din(new_Jinkela_wire_3308),
        .dout(new_Jinkela_wire_3309)
    );

    bfr new_Jinkela_buffer_9381 (
        .din(new_Jinkela_wire_11452),
        .dout(new_Jinkela_wire_11453)
    );

    bfr new_Jinkela_buffer_12905 (
        .din(new_Jinkela_wire_15426),
        .dout(new_Jinkela_wire_15427)
    );

    bfr new_Jinkela_buffer_12766 (
        .din(new_Jinkela_wire_15287),
        .dout(new_Jinkela_wire_15288)
    );

    bfr new_Jinkela_buffer_2436 (
        .din(new_Jinkela_wire_3433),
        .dout(new_Jinkela_wire_3434)
    );

    bfr new_Jinkela_buffer_9305 (
        .din(new_Jinkela_wire_11328),
        .dout(new_Jinkela_wire_11329)
    );

    bfr new_Jinkela_buffer_2322 (
        .din(new_Jinkela_wire_3309),
        .dout(new_Jinkela_wire_3310)
    );

    spl2 new_Jinkela_splitter_889 (
        .a(_0816_),
        .b(new_Jinkela_wire_11527),
        .c(new_Jinkela_wire_11528)
    );

    bfr new_Jinkela_buffer_12767 (
        .din(new_Jinkela_wire_15288),
        .dout(new_Jinkela_wire_15289)
    );

    bfr new_Jinkela_buffer_2389 (
        .din(new_Jinkela_wire_3380),
        .dout(new_Jinkela_wire_3381)
    );

    bfr new_Jinkela_buffer_9306 (
        .din(new_Jinkela_wire_11329),
        .dout(new_Jinkela_wire_11330)
    );

    bfr new_Jinkela_buffer_2323 (
        .din(new_Jinkela_wire_3310),
        .dout(new_Jinkela_wire_3311)
    );

    bfr new_Jinkela_buffer_9384 (
        .din(new_Jinkela_wire_11459),
        .dout(new_Jinkela_wire_11460)
    );

    bfr new_Jinkela_buffer_12906 (
        .din(new_Jinkela_wire_15427),
        .dout(new_Jinkela_wire_15428)
    );

    bfr new_Jinkela_buffer_12768 (
        .din(new_Jinkela_wire_15289),
        .dout(new_Jinkela_wire_15290)
    );

    bfr new_Jinkela_buffer_2402 (
        .din(new_Jinkela_wire_3395),
        .dout(new_Jinkela_wire_3396)
    );

    bfr new_Jinkela_buffer_9307 (
        .din(new_Jinkela_wire_11330),
        .dout(new_Jinkela_wire_11331)
    );

    bfr new_Jinkela_buffer_2324 (
        .din(new_Jinkela_wire_3311),
        .dout(new_Jinkela_wire_3312)
    );

    bfr new_Jinkela_buffer_13023 (
        .din(new_Jinkela_wire_15556),
        .dout(new_Jinkela_wire_15557)
    );

    bfr new_Jinkela_buffer_12769 (
        .din(new_Jinkela_wire_15290),
        .dout(new_Jinkela_wire_15291)
    );

    bfr new_Jinkela_buffer_2390 (
        .din(new_Jinkela_wire_3381),
        .dout(new_Jinkela_wire_3382)
    );

    bfr new_Jinkela_buffer_9308 (
        .din(new_Jinkela_wire_11331),
        .dout(new_Jinkela_wire_11332)
    );

    bfr new_Jinkela_buffer_12962 (
        .din(new_Jinkela_wire_15485),
        .dout(new_Jinkela_wire_15486)
    );

    bfr new_Jinkela_buffer_2325 (
        .din(new_Jinkela_wire_3312),
        .dout(new_Jinkela_wire_3313)
    );

    bfr new_Jinkela_buffer_9385 (
        .din(new_Jinkela_wire_11460),
        .dout(new_Jinkela_wire_11461)
    );

    bfr new_Jinkela_buffer_12907 (
        .din(new_Jinkela_wire_15428),
        .dout(new_Jinkela_wire_15429)
    );

    bfr new_Jinkela_buffer_12770 (
        .din(new_Jinkela_wire_15291),
        .dout(new_Jinkela_wire_15292)
    );

    bfr new_Jinkela_buffer_9309 (
        .din(new_Jinkela_wire_11332),
        .dout(new_Jinkela_wire_11333)
    );

    spl2 new_Jinkela_splitter_351 (
        .a(_0559_),
        .b(new_Jinkela_wire_3442),
        .c(new_Jinkela_wire_3443)
    );

    bfr new_Jinkela_buffer_2326 (
        .din(new_Jinkela_wire_3313),
        .dout(new_Jinkela_wire_3314)
    );

    spl2 new_Jinkela_splitter_890 (
        .a(_1735_),
        .b(new_Jinkela_wire_11529),
        .c(new_Jinkela_wire_11530)
    );

    bfr new_Jinkela_buffer_12771 (
        .din(new_Jinkela_wire_15292),
        .dout(new_Jinkela_wire_15293)
    );

    bfr new_Jinkela_buffer_2391 (
        .din(new_Jinkela_wire_3382),
        .dout(new_Jinkela_wire_3383)
    );

    bfr new_Jinkela_buffer_9310 (
        .din(new_Jinkela_wire_11333),
        .dout(new_Jinkela_wire_11334)
    );

    bfr new_Jinkela_buffer_2327 (
        .din(new_Jinkela_wire_3314),
        .dout(new_Jinkela_wire_3315)
    );

    bfr new_Jinkela_buffer_9386 (
        .din(new_Jinkela_wire_11461),
        .dout(new_Jinkela_wire_11462)
    );

    bfr new_Jinkela_buffer_12908 (
        .din(new_Jinkela_wire_15429),
        .dout(new_Jinkela_wire_15430)
    );

    bfr new_Jinkela_buffer_12772 (
        .din(new_Jinkela_wire_15293),
        .dout(new_Jinkela_wire_15294)
    );

    bfr new_Jinkela_buffer_2403 (
        .din(new_Jinkela_wire_3396),
        .dout(new_Jinkela_wire_3397)
    );

    bfr new_Jinkela_buffer_9311 (
        .din(new_Jinkela_wire_11334),
        .dout(new_Jinkela_wire_11335)
    );

    bfr new_Jinkela_buffer_2328 (
        .din(new_Jinkela_wire_3315),
        .dout(new_Jinkela_wire_3316)
    );

    bfr new_Jinkela_buffer_13002 (
        .din(new_Jinkela_wire_15531),
        .dout(new_Jinkela_wire_15532)
    );

    spl2 new_Jinkela_splitter_891 (
        .a(_0330_),
        .b(new_Jinkela_wire_11531),
        .c(new_Jinkela_wire_11532)
    );

    bfr new_Jinkela_buffer_12773 (
        .din(new_Jinkela_wire_15294),
        .dout(new_Jinkela_wire_15295)
    );

    bfr new_Jinkela_buffer_2392 (
        .din(new_Jinkela_wire_3383),
        .dout(new_Jinkela_wire_3384)
    );

    bfr new_Jinkela_buffer_9312 (
        .din(new_Jinkela_wire_11335),
        .dout(new_Jinkela_wire_11336)
    );

    bfr new_Jinkela_buffer_12963 (
        .din(new_Jinkela_wire_15486),
        .dout(new_Jinkela_wire_15487)
    );

    bfr new_Jinkela_buffer_2329 (
        .din(new_Jinkela_wire_3316),
        .dout(new_Jinkela_wire_3317)
    );

    bfr new_Jinkela_buffer_9387 (
        .din(new_Jinkela_wire_11462),
        .dout(new_Jinkela_wire_11463)
    );

    bfr new_Jinkela_buffer_12909 (
        .din(new_Jinkela_wire_15430),
        .dout(new_Jinkela_wire_15431)
    );

    bfr new_Jinkela_buffer_12774 (
        .din(new_Jinkela_wire_15295),
        .dout(new_Jinkela_wire_15296)
    );

    bfr new_Jinkela_buffer_9313 (
        .din(new_Jinkela_wire_11336),
        .dout(new_Jinkela_wire_11337)
    );

    bfr new_Jinkela_buffer_2330 (
        .din(new_Jinkela_wire_3317),
        .dout(new_Jinkela_wire_3318)
    );

    bfr new_Jinkela_buffer_9448 (
        .din(new_Jinkela_wire_11535),
        .dout(new_Jinkela_wire_11536)
    );

    bfr new_Jinkela_buffer_9447 (
        .din(_0188_),
        .dout(new_Jinkela_wire_11533)
    );

    bfr new_Jinkela_buffer_12775 (
        .din(new_Jinkela_wire_15296),
        .dout(new_Jinkela_wire_15297)
    );

    spl2 new_Jinkela_splitter_345 (
        .a(new_Jinkela_wire_3384),
        .b(new_Jinkela_wire_3385),
        .c(new_Jinkela_wire_3386)
    );

    spl2 new_Jinkela_splitter_861 (
        .a(new_Jinkela_wire_11337),
        .b(new_Jinkela_wire_11338),
        .c(new_Jinkela_wire_11339)
    );

    bfr new_Jinkela_buffer_2331 (
        .din(new_Jinkela_wire_3318),
        .dout(new_Jinkela_wire_3319)
    );

    bfr new_Jinkela_buffer_9452 (
        .din(_1365_),
        .dout(new_Jinkela_wire_11540)
    );

    bfr new_Jinkela_buffer_12910 (
        .din(new_Jinkela_wire_15431),
        .dout(new_Jinkela_wire_15432)
    );

    spl2 new_Jinkela_splitter_892 (
        .a(_0675_),
        .b(new_Jinkela_wire_11534),
        .c(new_Jinkela_wire_11535)
    );

    bfr new_Jinkela_buffer_12776 (
        .din(new_Jinkela_wire_15297),
        .dout(new_Jinkela_wire_15298)
    );

    bfr new_Jinkela_buffer_9388 (
        .din(new_Jinkela_wire_11463),
        .dout(new_Jinkela_wire_11464)
    );

    bfr new_Jinkela_buffer_2438 (
        .din(_0734_),
        .dout(new_Jinkela_wire_3446)
    );

    bfr new_Jinkela_buffer_2332 (
        .din(new_Jinkela_wire_3319),
        .dout(new_Jinkela_wire_3320)
    );

    bfr new_Jinkela_buffer_9389 (
        .din(new_Jinkela_wire_11464),
        .dout(new_Jinkela_wire_11465)
    );

    bfr new_Jinkela_buffer_12777 (
        .din(new_Jinkela_wire_15298),
        .dout(new_Jinkela_wire_15299)
    );

    bfr new_Jinkela_buffer_2404 (
        .din(new_Jinkela_wire_3397),
        .dout(new_Jinkela_wire_3398)
    );

    bfr new_Jinkela_buffer_12964 (
        .din(new_Jinkela_wire_15487),
        .dout(new_Jinkela_wire_15488)
    );

    bfr new_Jinkela_buffer_2333 (
        .din(new_Jinkela_wire_3320),
        .dout(new_Jinkela_wire_3321)
    );

    bfr new_Jinkela_buffer_9390 (
        .din(new_Jinkela_wire_11465),
        .dout(new_Jinkela_wire_11466)
    );

    bfr new_Jinkela_buffer_12911 (
        .din(new_Jinkela_wire_15432),
        .dout(new_Jinkela_wire_15433)
    );

    bfr new_Jinkela_buffer_12778 (
        .din(new_Jinkela_wire_15299),
        .dout(new_Jinkela_wire_15300)
    );

    bfr new_Jinkela_buffer_2405 (
        .din(new_Jinkela_wire_3398),
        .dout(new_Jinkela_wire_3399)
    );

    spl2 new_Jinkela_splitter_894 (
        .a(_0060_),
        .b(new_Jinkela_wire_11614),
        .c(new_Jinkela_wire_11615)
    );

    bfr new_Jinkela_buffer_2334 (
        .din(new_Jinkela_wire_3321),
        .dout(new_Jinkela_wire_3322)
    );

    bfr new_Jinkela_buffer_9391 (
        .din(new_Jinkela_wire_11466),
        .dout(new_Jinkela_wire_11467)
    );

    bfr new_Jinkela_buffer_12779 (
        .din(new_Jinkela_wire_15300),
        .dout(new_Jinkela_wire_15301)
    );

    bfr new_Jinkela_buffer_2439 (
        .din(_0106_),
        .dout(new_Jinkela_wire_3449)
    );

    spl2 new_Jinkela_splitter_353 (
        .a(_0798_),
        .b(new_Jinkela_wire_3447),
        .c(new_Jinkela_wire_3448)
    );

    spl2 new_Jinkela_splitter_895 (
        .a(_1189_),
        .b(new_Jinkela_wire_11616),
        .c(new_Jinkela_wire_11617)
    );

    bfr new_Jinkela_buffer_13126 (
        .din(_0389_),
        .dout(new_Jinkela_wire_15666)
    );

    bfr new_Jinkela_buffer_2335 (
        .din(new_Jinkela_wire_3322),
        .dout(new_Jinkela_wire_3323)
    );

    bfr new_Jinkela_buffer_9392 (
        .din(new_Jinkela_wire_11467),
        .dout(new_Jinkela_wire_11468)
    );

    bfr new_Jinkela_buffer_12912 (
        .din(new_Jinkela_wire_15433),
        .dout(new_Jinkela_wire_15434)
    );

    bfr new_Jinkela_buffer_12780 (
        .din(new_Jinkela_wire_15301),
        .dout(new_Jinkela_wire_15302)
    );

    bfr new_Jinkela_buffer_2406 (
        .din(new_Jinkela_wire_3399),
        .dout(new_Jinkela_wire_3400)
    );

    bfr new_Jinkela_buffer_9449 (
        .din(new_Jinkela_wire_11536),
        .dout(new_Jinkela_wire_11537)
    );

    bfr new_Jinkela_buffer_2336 (
        .din(new_Jinkela_wire_3323),
        .dout(new_Jinkela_wire_3324)
    );

    bfr new_Jinkela_buffer_9393 (
        .din(new_Jinkela_wire_11468),
        .dout(new_Jinkela_wire_11469)
    );

    bfr new_Jinkela_buffer_13003 (
        .din(new_Jinkela_wire_15532),
        .dout(new_Jinkela_wire_15533)
    );

    bfr new_Jinkela_buffer_12781 (
        .din(new_Jinkela_wire_15302),
        .dout(new_Jinkela_wire_15303)
    );

    spl2 new_Jinkela_splitter_355 (
        .a(_0937_),
        .b(new_Jinkela_wire_3483),
        .c(new_Jinkela_wire_3484)
    );

    bfr new_Jinkela_buffer_9453 (
        .din(new_Jinkela_wire_11540),
        .dout(new_Jinkela_wire_11541)
    );

    bfr new_Jinkela_buffer_12965 (
        .din(new_Jinkela_wire_15488),
        .dout(new_Jinkela_wire_15489)
    );

    bfr new_Jinkela_buffer_2337 (
        .din(new_Jinkela_wire_3324),
        .dout(new_Jinkela_wire_3325)
    );

    bfr new_Jinkela_buffer_9394 (
        .din(new_Jinkela_wire_11469),
        .dout(new_Jinkela_wire_11470)
    );

    bfr new_Jinkela_buffer_12913 (
        .din(new_Jinkela_wire_15434),
        .dout(new_Jinkela_wire_15435)
    );

    bfr new_Jinkela_buffer_12782 (
        .din(new_Jinkela_wire_15303),
        .dout(new_Jinkela_wire_15304)
    );

    bfr new_Jinkela_buffer_2407 (
        .din(new_Jinkela_wire_3400),
        .dout(new_Jinkela_wire_3401)
    );

    bfr new_Jinkela_buffer_9450 (
        .din(new_Jinkela_wire_11537),
        .dout(new_Jinkela_wire_11538)
    );

    and_bb _3298_ (
        .a(new_Jinkela_wire_17990),
        .b(new_Jinkela_wire_9093),
        .c(_0574_)
    );

    or_bb _3299_ (
        .a(new_Jinkela_wire_10694),
        .b(new_Jinkela_wire_8589),
        .c(_0575_)
    );

    and_ii _3300_ (
        .a(new_Jinkela_wire_2460),
        .b(new_Jinkela_wire_17636),
        .c(_0576_)
    );

    and_bb _3301_ (
        .a(new_Jinkela_wire_2461),
        .b(new_Jinkela_wire_17637),
        .c(_0577_)
    );

    or_bb _3302_ (
        .a(new_Jinkela_wire_15025),
        .b(new_Jinkela_wire_4477),
        .c(_0578_)
    );

    and_ii _3303_ (
        .a(new_Jinkela_wire_6368),
        .b(new_Jinkela_wire_13673),
        .c(_0580_)
    );

    and_bb _3304_ (
        .a(new_Jinkela_wire_6369),
        .b(new_Jinkela_wire_13674),
        .c(_0581_)
    );

    or_bb _3305_ (
        .a(new_Jinkela_wire_16214),
        .b(new_Jinkela_wire_6409),
        .c(_0582_)
    );

    and_ii _3306_ (
        .a(new_Jinkela_wire_21108),
        .b(new_Jinkela_wire_1904),
        .c(_0583_)
    );

    and_bb _3307_ (
        .a(new_Jinkela_wire_21109),
        .b(new_Jinkela_wire_1905),
        .c(_0584_)
    );

    or_bb _3308_ (
        .a(new_Jinkela_wire_2819),
        .b(new_Jinkela_wire_9101),
        .c(_0585_)
    );

    and_ii _3309_ (
        .a(new_Jinkela_wire_5144),
        .b(new_Jinkela_wire_15117),
        .c(_0586_)
    );

    and_bb _3310_ (
        .a(new_Jinkela_wire_5145),
        .b(new_Jinkela_wire_15118),
        .c(_0587_)
    );

    or_bb _3311_ (
        .a(new_Jinkela_wire_18797),
        .b(new_Jinkela_wire_4678),
        .c(_0588_)
    );

    and_ii _3312_ (
        .a(new_Jinkela_wire_12731),
        .b(new_Jinkela_wire_16957),
        .c(_0589_)
    );

    and_bb _3313_ (
        .a(new_Jinkela_wire_12732),
        .b(new_Jinkela_wire_16958),
        .c(_0591_)
    );

    or_bb _3314_ (
        .a(new_Jinkela_wire_11447),
        .b(new_Jinkela_wire_10574),
        .c(_0592_)
    );

    and_ii _3315_ (
        .a(new_Jinkela_wire_18448),
        .b(new_Jinkela_wire_8460),
        .c(_0593_)
    );

    and_bb _3316_ (
        .a(new_Jinkela_wire_18449),
        .b(new_Jinkela_wire_8461),
        .c(_0594_)
    );

    or_bb _3317_ (
        .a(new_Jinkela_wire_20216),
        .b(new_Jinkela_wire_13683),
        .c(_0595_)
    );

    and_ii _3318_ (
        .a(new_Jinkela_wire_5142),
        .b(new_Jinkela_wire_4907),
        .c(_0596_)
    );

    and_bb _3319_ (
        .a(new_Jinkela_wire_5143),
        .b(new_Jinkela_wire_4908),
        .c(_0597_)
    );

    or_bb _3320_ (
        .a(new_Jinkela_wire_7718),
        .b(new_Jinkela_wire_7695),
        .c(_0598_)
    );

    and_ii _3321_ (
        .a(new_Jinkela_wire_19737),
        .b(new_Jinkela_wire_13570),
        .c(_0599_)
    );

    and_bb _3322_ (
        .a(new_Jinkela_wire_19738),
        .b(new_Jinkela_wire_13571),
        .c(_0600_)
    );

    or_bb _3323_ (
        .a(new_Jinkela_wire_18808),
        .b(new_Jinkela_wire_12060),
        .c(_0602_)
    );

    and_ii _3324_ (
        .a(new_Jinkela_wire_16215),
        .b(new_Jinkela_wire_19055),
        .c(_0603_)
    );

    and_bb _3325_ (
        .a(new_Jinkela_wire_16216),
        .b(new_Jinkela_wire_19056),
        .c(_0604_)
    );

    or_bb _3326_ (
        .a(new_Jinkela_wire_2464),
        .b(new_Jinkela_wire_15734),
        .c(_0605_)
    );

    and_ii _3327_ (
        .a(new_Jinkela_wire_9807),
        .b(new_Jinkela_wire_2932),
        .c(_0606_)
    );

    and_bb _3328_ (
        .a(new_Jinkela_wire_9808),
        .b(new_Jinkela_wire_2933),
        .c(_0607_)
    );

    or_bb _3329_ (
        .a(new_Jinkela_wire_9349),
        .b(new_Jinkela_wire_14086),
        .c(_0608_)
    );

    and_ii _3330_ (
        .a(new_Jinkela_wire_10614),
        .b(new_Jinkela_wire_13402),
        .c(_0609_)
    );

    and_bb _3331_ (
        .a(new_Jinkela_wire_10615),
        .b(new_Jinkela_wire_13403),
        .c(_0610_)
    );

    and_ii _3332_ (
        .a(new_Jinkela_wire_3260),
        .b(new_Jinkela_wire_21124),
        .c(_0611_)
    );

    and_bb _3333_ (
        .a(new_Jinkela_wire_5986),
        .b(new_Jinkela_wire_2481),
        .c(_0613_)
    );

    and_ii _3334_ (
        .a(new_Jinkela_wire_5987),
        .b(new_Jinkela_wire_2482),
        .c(_0614_)
    );

    or_bb _3335_ (
        .a(new_Jinkela_wire_14283),
        .b(new_Jinkela_wire_1775),
        .c(new_net_3966)
    );

    or_bb _3336_ (
        .a(new_Jinkela_wire_1776),
        .b(new_Jinkela_wire_21145),
        .c(_0615_)
    );

    and_ii _3337_ (
        .a(new_Jinkela_wire_14087),
        .b(new_Jinkela_wire_15739),
        .c(_0616_)
    );

    and_bb _3338_ (
        .a(new_Jinkela_wire_695),
        .b(new_Jinkela_wire_668),
        .c(_0617_)
    );

    and_ii _3339_ (
        .a(new_Jinkela_wire_12061),
        .b(new_Jinkela_wire_7700),
        .c(_0618_)
    );

    bfr new_Jinkela_buffer_5824 (
        .din(new_Jinkela_wire_7413),
        .dout(new_Jinkela_wire_7414)
    );

    bfr new_Jinkela_buffer_2338 (
        .din(new_Jinkela_wire_3325),
        .dout(new_Jinkela_wire_3326)
    );

    bfr new_Jinkela_buffer_16308 (
        .din(new_Jinkela_wire_19474),
        .dout(new_Jinkela_wire_19475)
    );

    bfr new_Jinkela_buffer_16204 (
        .din(new_Jinkela_wire_19364),
        .dout(new_Jinkela_wire_19365)
    );

    bfr new_Jinkela_buffer_5979 (
        .din(new_Jinkela_wire_7594),
        .dout(new_Jinkela_wire_7595)
    );

    bfr new_Jinkela_buffer_2471 (
        .din(_0340_),
        .dout(new_Jinkela_wire_3485)
    );

    bfr new_Jinkela_buffer_5825 (
        .din(new_Jinkela_wire_7414),
        .dout(new_Jinkela_wire_7415)
    );

    bfr new_Jinkela_buffer_2339 (
        .din(new_Jinkela_wire_3326),
        .dout(new_Jinkela_wire_3327)
    );

    bfr new_Jinkela_buffer_16236 (
        .din(new_Jinkela_wire_19398),
        .dout(new_Jinkela_wire_19399)
    );

    bfr new_Jinkela_buffer_5894 (
        .din(new_Jinkela_wire_7491),
        .dout(new_Jinkela_wire_7492)
    );

    bfr new_Jinkela_buffer_2408 (
        .din(new_Jinkela_wire_3401),
        .dout(new_Jinkela_wire_3402)
    );

    bfr new_Jinkela_buffer_16205 (
        .din(new_Jinkela_wire_19365),
        .dout(new_Jinkela_wire_19366)
    );

    bfr new_Jinkela_buffer_5826 (
        .din(new_Jinkela_wire_7415),
        .dout(new_Jinkela_wire_7416)
    );

    bfr new_Jinkela_buffer_2340 (
        .din(new_Jinkela_wire_3327),
        .dout(new_Jinkela_wire_3328)
    );

    bfr new_Jinkela_buffer_16305 (
        .din(new_Jinkela_wire_19471),
        .dout(new_Jinkela_wire_19472)
    );

    bfr new_Jinkela_buffer_5923 (
        .din(new_Jinkela_wire_7530),
        .dout(new_Jinkela_wire_7531)
    );

    bfr new_Jinkela_buffer_2440 (
        .din(new_Jinkela_wire_3449),
        .dout(new_Jinkela_wire_3450)
    );

    bfr new_Jinkela_buffer_16206 (
        .din(new_Jinkela_wire_19366),
        .dout(new_Jinkela_wire_19367)
    );

    bfr new_Jinkela_buffer_5827 (
        .din(new_Jinkela_wire_7416),
        .dout(new_Jinkela_wire_7417)
    );

    bfr new_Jinkela_buffer_2341 (
        .din(new_Jinkela_wire_3328),
        .dout(new_Jinkela_wire_3329)
    );

    bfr new_Jinkela_buffer_16237 (
        .din(new_Jinkela_wire_19399),
        .dout(new_Jinkela_wire_19400)
    );

    bfr new_Jinkela_buffer_5895 (
        .din(new_Jinkela_wire_7492),
        .dout(new_Jinkela_wire_7493)
    );

    bfr new_Jinkela_buffer_2409 (
        .din(new_Jinkela_wire_3402),
        .dout(new_Jinkela_wire_3403)
    );

    bfr new_Jinkela_buffer_16207 (
        .din(new_Jinkela_wire_19367),
        .dout(new_Jinkela_wire_19368)
    );

    bfr new_Jinkela_buffer_5828 (
        .din(new_Jinkela_wire_7417),
        .dout(new_Jinkela_wire_7418)
    );

    bfr new_Jinkela_buffer_2342 (
        .din(new_Jinkela_wire_3329),
        .dout(new_Jinkela_wire_3330)
    );

    bfr new_Jinkela_buffer_16208 (
        .din(new_Jinkela_wire_19368),
        .dout(new_Jinkela_wire_19369)
    );

    bfr new_Jinkela_buffer_2536 (
        .din(_1247_),
        .dout(new_Jinkela_wire_3552)
    );

    spl2 new_Jinkela_splitter_662 (
        .a(_0024_),
        .b(new_Jinkela_wire_7703),
        .c(new_Jinkela_wire_7704)
    );

    bfr new_Jinkela_buffer_5829 (
        .din(new_Jinkela_wire_7418),
        .dout(new_Jinkela_wire_7419)
    );

    bfr new_Jinkela_buffer_2343 (
        .din(new_Jinkela_wire_3330),
        .dout(new_Jinkela_wire_3331)
    );

    bfr new_Jinkela_buffer_16238 (
        .din(new_Jinkela_wire_19400),
        .dout(new_Jinkela_wire_19401)
    );

    bfr new_Jinkela_buffer_5896 (
        .din(new_Jinkela_wire_7493),
        .dout(new_Jinkela_wire_7494)
    );

    bfr new_Jinkela_buffer_2410 (
        .din(new_Jinkela_wire_3403),
        .dout(new_Jinkela_wire_3404)
    );

    bfr new_Jinkela_buffer_16209 (
        .din(new_Jinkela_wire_19369),
        .dout(new_Jinkela_wire_19370)
    );

    bfr new_Jinkela_buffer_5830 (
        .din(new_Jinkela_wire_7419),
        .dout(new_Jinkela_wire_7420)
    );

    bfr new_Jinkela_buffer_2344 (
        .din(new_Jinkela_wire_3331),
        .dout(new_Jinkela_wire_3332)
    );

    bfr new_Jinkela_buffer_16306 (
        .din(new_Jinkela_wire_19472),
        .dout(new_Jinkela_wire_19473)
    );

    bfr new_Jinkela_buffer_5924 (
        .din(new_Jinkela_wire_7531),
        .dout(new_Jinkela_wire_7532)
    );

    bfr new_Jinkela_buffer_2441 (
        .din(new_Jinkela_wire_3450),
        .dout(new_Jinkela_wire_3451)
    );

    bfr new_Jinkela_buffer_16210 (
        .din(new_Jinkela_wire_19370),
        .dout(new_Jinkela_wire_19371)
    );

    bfr new_Jinkela_buffer_5831 (
        .din(new_Jinkela_wire_7420),
        .dout(new_Jinkela_wire_7421)
    );

    bfr new_Jinkela_buffer_2345 (
        .din(new_Jinkela_wire_3332),
        .dout(new_Jinkela_wire_3333)
    );

    bfr new_Jinkela_buffer_16239 (
        .din(new_Jinkela_wire_19401),
        .dout(new_Jinkela_wire_19402)
    );

    bfr new_Jinkela_buffer_5897 (
        .din(new_Jinkela_wire_7494),
        .dout(new_Jinkela_wire_7495)
    );

    bfr new_Jinkela_buffer_2411 (
        .din(new_Jinkela_wire_3404),
        .dout(new_Jinkela_wire_3405)
    );

    bfr new_Jinkela_buffer_16211 (
        .din(new_Jinkela_wire_19371),
        .dout(new_Jinkela_wire_19372)
    );

    bfr new_Jinkela_buffer_5832 (
        .din(new_Jinkela_wire_7421),
        .dout(new_Jinkela_wire_7422)
    );

    bfr new_Jinkela_buffer_2346 (
        .din(new_Jinkela_wire_3333),
        .dout(new_Jinkela_wire_3334)
    );

    bfr new_Jinkela_buffer_16309 (
        .din(new_Jinkela_wire_19475),
        .dout(new_Jinkela_wire_19476)
    );

    bfr new_Jinkela_buffer_16212 (
        .din(new_Jinkela_wire_19372),
        .dout(new_Jinkela_wire_19373)
    );

    bfr new_Jinkela_buffer_5980 (
        .din(new_Jinkela_wire_7595),
        .dout(new_Jinkela_wire_7596)
    );

    bfr new_Jinkela_buffer_2535 (
        .din(_0310_),
        .dout(new_Jinkela_wire_3551)
    );

    bfr new_Jinkela_buffer_5833 (
        .din(new_Jinkela_wire_7422),
        .dout(new_Jinkela_wire_7423)
    );

    bfr new_Jinkela_buffer_2347 (
        .din(new_Jinkela_wire_3334),
        .dout(new_Jinkela_wire_3335)
    );

    bfr new_Jinkela_buffer_16240 (
        .din(new_Jinkela_wire_19402),
        .dout(new_Jinkela_wire_19403)
    );

    bfr new_Jinkela_buffer_5898 (
        .din(new_Jinkela_wire_7495),
        .dout(new_Jinkela_wire_7496)
    );

    bfr new_Jinkela_buffer_2412 (
        .din(new_Jinkela_wire_3405),
        .dout(new_Jinkela_wire_3406)
    );

    bfr new_Jinkela_buffer_16213 (
        .din(new_Jinkela_wire_19373),
        .dout(new_Jinkela_wire_19374)
    );

    bfr new_Jinkela_buffer_5834 (
        .din(new_Jinkela_wire_7423),
        .dout(new_Jinkela_wire_7424)
    );

    bfr new_Jinkela_buffer_2348 (
        .din(new_Jinkela_wire_3335),
        .dout(new_Jinkela_wire_3336)
    );

    spl2 new_Jinkela_splitter_1435 (
        .a(_1528_),
        .b(new_Jinkela_wire_19544),
        .c(new_Jinkela_wire_19545)
    );

    bfr new_Jinkela_buffer_5925 (
        .din(new_Jinkela_wire_7532),
        .dout(new_Jinkela_wire_7533)
    );

    bfr new_Jinkela_buffer_2442 (
        .din(new_Jinkela_wire_3451),
        .dout(new_Jinkela_wire_3452)
    );

    bfr new_Jinkela_buffer_16214 (
        .din(new_Jinkela_wire_19374),
        .dout(new_Jinkela_wire_19375)
    );

    bfr new_Jinkela_buffer_5835 (
        .din(new_Jinkela_wire_7424),
        .dout(new_Jinkela_wire_7425)
    );

    bfr new_Jinkela_buffer_2349 (
        .din(new_Jinkela_wire_3336),
        .dout(new_Jinkela_wire_3337)
    );

    bfr new_Jinkela_buffer_16241 (
        .din(new_Jinkela_wire_19403),
        .dout(new_Jinkela_wire_19404)
    );

    bfr new_Jinkela_buffer_5899 (
        .din(new_Jinkela_wire_7496),
        .dout(new_Jinkela_wire_7497)
    );

    bfr new_Jinkela_buffer_2413 (
        .din(new_Jinkela_wire_3406),
        .dout(new_Jinkela_wire_3407)
    );

    bfr new_Jinkela_buffer_16215 (
        .din(new_Jinkela_wire_19375),
        .dout(new_Jinkela_wire_19376)
    );

    bfr new_Jinkela_buffer_5836 (
        .din(new_Jinkela_wire_7425),
        .dout(new_Jinkela_wire_7426)
    );

    bfr new_Jinkela_buffer_2350 (
        .din(new_Jinkela_wire_3337),
        .dout(new_Jinkela_wire_3338)
    );

    bfr new_Jinkela_buffer_16310 (
        .din(new_Jinkela_wire_19476),
        .dout(new_Jinkela_wire_19477)
    );

    spl2 new_Jinkela_splitter_663 (
        .a(_1032_),
        .b(new_Jinkela_wire_7705),
        .c(new_Jinkela_wire_7706)
    );

    bfr new_Jinkela_buffer_2472 (
        .din(new_Jinkela_wire_3485),
        .dout(new_Jinkela_wire_3486)
    );

    bfr new_Jinkela_buffer_16216 (
        .din(new_Jinkela_wire_19376),
        .dout(new_Jinkela_wire_19377)
    );

    bfr new_Jinkela_buffer_5837 (
        .din(new_Jinkela_wire_7426),
        .dout(new_Jinkela_wire_7427)
    );

    bfr new_Jinkela_buffer_2351 (
        .din(new_Jinkela_wire_3338),
        .dout(new_Jinkela_wire_3339)
    );

    bfr new_Jinkela_buffer_16242 (
        .din(new_Jinkela_wire_19404),
        .dout(new_Jinkela_wire_19405)
    );

    bfr new_Jinkela_buffer_5900 (
        .din(new_Jinkela_wire_7497),
        .dout(new_Jinkela_wire_7498)
    );

    bfr new_Jinkela_buffer_2414 (
        .din(new_Jinkela_wire_3407),
        .dout(new_Jinkela_wire_3408)
    );

    bfr new_Jinkela_buffer_16217 (
        .din(new_Jinkela_wire_19377),
        .dout(new_Jinkela_wire_19378)
    );

    bfr new_Jinkela_buffer_5838 (
        .din(new_Jinkela_wire_7427),
        .dout(new_Jinkela_wire_7428)
    );

    bfr new_Jinkela_buffer_2352 (
        .din(new_Jinkela_wire_3339),
        .dout(new_Jinkela_wire_3340)
    );

    spl2 new_Jinkela_splitter_1436 (
        .a(_1099_),
        .b(new_Jinkela_wire_19546),
        .c(new_Jinkela_wire_19547)
    );

    bfr new_Jinkela_buffer_5926 (
        .din(new_Jinkela_wire_7533),
        .dout(new_Jinkela_wire_7534)
    );

    bfr new_Jinkela_buffer_2443 (
        .din(new_Jinkela_wire_3452),
        .dout(new_Jinkela_wire_3453)
    );

    bfr new_Jinkela_buffer_16218 (
        .din(new_Jinkela_wire_19378),
        .dout(new_Jinkela_wire_19379)
    );

    bfr new_Jinkela_buffer_5839 (
        .din(new_Jinkela_wire_7428),
        .dout(new_Jinkela_wire_7429)
    );

    bfr new_Jinkela_buffer_2353 (
        .din(new_Jinkela_wire_3340),
        .dout(new_Jinkela_wire_3341)
    );

    bfr new_Jinkela_buffer_16243 (
        .din(new_Jinkela_wire_19405),
        .dout(new_Jinkela_wire_19406)
    );

    bfr new_Jinkela_buffer_5901 (
        .din(new_Jinkela_wire_7498),
        .dout(new_Jinkela_wire_7499)
    );

    bfr new_Jinkela_buffer_2415 (
        .din(new_Jinkela_wire_3408),
        .dout(new_Jinkela_wire_3409)
    );

    bfr new_Jinkela_buffer_16219 (
        .din(new_Jinkela_wire_19379),
        .dout(new_Jinkela_wire_19380)
    );

    bfr new_Jinkela_buffer_5840 (
        .din(new_Jinkela_wire_7429),
        .dout(new_Jinkela_wire_7430)
    );

    bfr new_Jinkela_buffer_2354 (
        .din(new_Jinkela_wire_3341),
        .dout(new_Jinkela_wire_3342)
    );

    bfr new_Jinkela_buffer_16311 (
        .din(new_Jinkela_wire_19477),
        .dout(new_Jinkela_wire_19478)
    );

    bfr new_Jinkela_buffer_16220 (
        .din(new_Jinkela_wire_19380),
        .dout(new_Jinkela_wire_19381)
    );

    bfr new_Jinkela_buffer_5981 (
        .din(new_Jinkela_wire_7596),
        .dout(new_Jinkela_wire_7597)
    );

    spl2 new_Jinkela_splitter_357 (
        .a(_1270_),
        .b(new_Jinkela_wire_3553),
        .c(new_Jinkela_wire_3554)
    );

    bfr new_Jinkela_buffer_5841 (
        .din(new_Jinkela_wire_7430),
        .dout(new_Jinkela_wire_7431)
    );

    bfr new_Jinkela_buffer_2355 (
        .din(new_Jinkela_wire_3342),
        .dout(new_Jinkela_wire_3343)
    );

    bfr new_Jinkela_buffer_16244 (
        .din(new_Jinkela_wire_19406),
        .dout(new_Jinkela_wire_19407)
    );

    spl2 new_Jinkela_splitter_648 (
        .a(new_Jinkela_wire_7499),
        .b(new_Jinkela_wire_7500),
        .c(new_Jinkela_wire_7501)
    );

    bfr new_Jinkela_buffer_2416 (
        .din(new_Jinkela_wire_3409),
        .dout(new_Jinkela_wire_3410)
    );

    bfr new_Jinkela_buffer_16221 (
        .din(new_Jinkela_wire_19381),
        .dout(new_Jinkela_wire_19382)
    );

    bfr new_Jinkela_buffer_5842 (
        .din(new_Jinkela_wire_7431),
        .dout(new_Jinkela_wire_7432)
    );

    bfr new_Jinkela_buffer_2356 (
        .din(new_Jinkela_wire_3343),
        .dout(new_Jinkela_wire_3344)
    );

    spl2 new_Jinkela_splitter_1438 (
        .a(_1378_),
        .b(new_Jinkela_wire_19554),
        .c(new_Jinkela_wire_19555)
    );

    spl2 new_Jinkela_splitter_1437 (
        .a(_1435_),
        .b(new_Jinkela_wire_19548),
        .c(new_Jinkela_wire_19549)
    );

    bfr new_Jinkela_buffer_6074 (
        .din(new_Jinkela_wire_7697),
        .dout(new_Jinkela_wire_7698)
    );

    bfr new_Jinkela_buffer_2444 (
        .din(new_Jinkela_wire_3453),
        .dout(new_Jinkela_wire_3454)
    );

    bfr new_Jinkela_buffer_16222 (
        .din(new_Jinkela_wire_19382),
        .dout(new_Jinkela_wire_19383)
    );

    bfr new_Jinkela_buffer_5843 (
        .din(new_Jinkela_wire_7432),
        .dout(new_Jinkela_wire_7433)
    );

    bfr new_Jinkela_buffer_2357 (
        .din(new_Jinkela_wire_3344),
        .dout(new_Jinkela_wire_3345)
    );

    bfr new_Jinkela_buffer_16245 (
        .din(new_Jinkela_wire_19407),
        .dout(new_Jinkela_wire_19408)
    );

    bfr new_Jinkela_buffer_5927 (
        .din(new_Jinkela_wire_7534),
        .dout(new_Jinkela_wire_7535)
    );

    bfr new_Jinkela_buffer_2417 (
        .din(new_Jinkela_wire_3410),
        .dout(new_Jinkela_wire_3411)
    );

    bfr new_Jinkela_buffer_16223 (
        .din(new_Jinkela_wire_19383),
        .dout(new_Jinkela_wire_19384)
    );

    bfr new_Jinkela_buffer_5844 (
        .din(new_Jinkela_wire_7433),
        .dout(new_Jinkela_wire_7434)
    );

    bfr new_Jinkela_buffer_2358 (
        .din(new_Jinkela_wire_3345),
        .dout(new_Jinkela_wire_3346)
    );

    bfr new_Jinkela_buffer_16312 (
        .din(new_Jinkela_wire_19478),
        .dout(new_Jinkela_wire_19479)
    );

    bfr new_Jinkela_buffer_5928 (
        .din(new_Jinkela_wire_7535),
        .dout(new_Jinkela_wire_7536)
    );

    bfr new_Jinkela_buffer_2473 (
        .din(new_Jinkela_wire_3486),
        .dout(new_Jinkela_wire_3487)
    );

    bfr new_Jinkela_buffer_16224 (
        .din(new_Jinkela_wire_19384),
        .dout(new_Jinkela_wire_19385)
    );

    bfr new_Jinkela_buffer_16246 (
        .din(new_Jinkela_wire_19408),
        .dout(new_Jinkela_wire_19409)
    );

    or_bi _2413_ (
        .a(new_Jinkela_wire_10276),
        .b(new_Jinkela_wire_9544),
        .c(_1449_)
    );

    bfr new_Jinkela_buffer_12783 (
        .din(new_Jinkela_wire_15304),
        .dout(new_Jinkela_wire_15305)
    );

    bfr new_Jinkela_buffer_16225 (
        .din(new_Jinkela_wire_19385),
        .dout(new_Jinkela_wire_19386)
    );

    and_ii _2414_ (
        .a(new_Jinkela_wire_5133),
        .b(new_Jinkela_wire_1761),
        .c(_1450_)
    );

    bfr new_Jinkela_buffer_12914 (
        .din(new_Jinkela_wire_15435),
        .dout(new_Jinkela_wire_15436)
    );

    bfr new_Jinkela_buffer_16371 (
        .din(new_Jinkela_wire_19549),
        .dout(new_Jinkela_wire_19550)
    );

    and_bb _2415_ (
        .a(new_Jinkela_wire_5134),
        .b(new_Jinkela_wire_1762),
        .c(_1451_)
    );

    bfr new_Jinkela_buffer_12784 (
        .din(new_Jinkela_wire_15305),
        .dout(new_Jinkela_wire_15306)
    );

    bfr new_Jinkela_buffer_16226 (
        .din(new_Jinkela_wire_19386),
        .dout(new_Jinkela_wire_19387)
    );

    or_bb _2416_ (
        .a(new_Jinkela_wire_15730),
        .b(new_Jinkela_wire_8839),
        .c(new_net_3952)
    );

    bfr new_Jinkela_buffer_13024 (
        .din(new_Jinkela_wire_15557),
        .dout(new_Jinkela_wire_15558)
    );

    bfr new_Jinkela_buffer_16247 (
        .din(new_Jinkela_wire_19409),
        .dout(new_Jinkela_wire_19410)
    );

    and_bb _2417_ (
        .a(new_Jinkela_wire_140),
        .b(new_Jinkela_wire_342),
        .c(_1452_)
    );

    bfr new_Jinkela_buffer_12785 (
        .din(new_Jinkela_wire_15306),
        .dout(new_Jinkela_wire_15307)
    );

    bfr new_Jinkela_buffer_16227 (
        .din(new_Jinkela_wire_19387),
        .dout(new_Jinkela_wire_19388)
    );

    and_bi _2418_ (
        .a(new_Jinkela_wire_9549),
        .b(new_Jinkela_wire_8840),
        .c(_1453_)
    );

    bfr new_Jinkela_buffer_12966 (
        .din(new_Jinkela_wire_15489),
        .dout(new_Jinkela_wire_15490)
    );

    bfr new_Jinkela_buffer_12915 (
        .din(new_Jinkela_wire_15436),
        .dout(new_Jinkela_wire_15437)
    );

    bfr new_Jinkela_buffer_16313 (
        .din(new_Jinkela_wire_19479),
        .dout(new_Jinkela_wire_19480)
    );

    and_bb _2419_ (
        .a(new_Jinkela_wire_90),
        .b(new_Jinkela_wire_213),
        .c(_1454_)
    );

    bfr new_Jinkela_buffer_12786 (
        .din(new_Jinkela_wire_15307),
        .dout(new_Jinkela_wire_15308)
    );

    bfr new_Jinkela_buffer_16228 (
        .din(new_Jinkela_wire_19388),
        .dout(new_Jinkela_wire_19389)
    );

    and_bi _2420_ (
        .a(new_Jinkela_wire_9606),
        .b(new_Jinkela_wire_14027),
        .c(_1455_)
    );

    bfr new_Jinkela_buffer_16248 (
        .din(new_Jinkela_wire_19410),
        .dout(new_Jinkela_wire_19411)
    );

    and_bb _2421_ (
        .a(new_Jinkela_wire_588),
        .b(new_Jinkela_wire_560),
        .c(_1456_)
    );

    bfr new_Jinkela_buffer_12787 (
        .din(new_Jinkela_wire_15308),
        .dout(new_Jinkela_wire_15309)
    );

    bfr new_Jinkela_buffer_16229 (
        .din(new_Jinkela_wire_19389),
        .dout(new_Jinkela_wire_19390)
    );

    and_bi _2422_ (
        .a(new_Jinkela_wire_19553),
        .b(new_Jinkela_wire_17044),
        .c(_1457_)
    );

    bfr new_Jinkela_buffer_12916 (
        .din(new_Jinkela_wire_15437),
        .dout(new_Jinkela_wire_15438)
    );

    and_bb _2423_ (
        .a(new_Jinkela_wire_274),
        .b(new_Jinkela_wire_117),
        .c(_1459_)
    );

    bfr new_Jinkela_buffer_12788 (
        .din(new_Jinkela_wire_15309),
        .dout(new_Jinkela_wire_15310)
    );

    spl2 new_Jinkela_splitter_1439 (
        .a(_0438_),
        .b(new_Jinkela_wire_19556),
        .c(new_Jinkela_wire_19557)
    );

    spl2 new_Jinkela_splitter_1429 (
        .a(new_Jinkela_wire_19390),
        .b(new_Jinkela_wire_19391),
        .c(new_Jinkela_wire_19392)
    );

    and_bi _2424_ (
        .a(new_Jinkela_wire_21213),
        .b(new_Jinkela_wire_5545),
        .c(_1460_)
    );

    bfr new_Jinkela_buffer_13004 (
        .din(new_Jinkela_wire_15533),
        .dout(new_Jinkela_wire_15534)
    );

    bfr new_Jinkela_buffer_16314 (
        .din(new_Jinkela_wire_19480),
        .dout(new_Jinkela_wire_19481)
    );

    and_bb _2425_ (
        .a(new_Jinkela_wire_75),
        .b(new_Jinkela_wire_1),
        .c(_1461_)
    );

    bfr new_Jinkela_buffer_12789 (
        .din(new_Jinkela_wire_15310),
        .dout(new_Jinkela_wire_15311)
    );

    bfr new_Jinkela_buffer_16249 (
        .din(new_Jinkela_wire_19411),
        .dout(new_Jinkela_wire_19412)
    );

    and_bi _2426_ (
        .a(new_Jinkela_wire_6201),
        .b(new_Jinkela_wire_13731),
        .c(_1462_)
    );

    bfr new_Jinkela_buffer_12967 (
        .din(new_Jinkela_wire_15490),
        .dout(new_Jinkela_wire_15491)
    );

    bfr new_Jinkela_buffer_12917 (
        .din(new_Jinkela_wire_15438),
        .dout(new_Jinkela_wire_15439)
    );

    bfr new_Jinkela_buffer_16250 (
        .din(new_Jinkela_wire_19412),
        .dout(new_Jinkela_wire_19413)
    );

    and_bb _2427_ (
        .a(new_Jinkela_wire_467),
        .b(new_Jinkela_wire_453),
        .c(_1463_)
    );

    bfr new_Jinkela_buffer_12790 (
        .din(new_Jinkela_wire_15311),
        .dout(new_Jinkela_wire_15312)
    );

    and_bi _2428_ (
        .a(new_Jinkela_wire_10096),
        .b(new_Jinkela_wire_2260),
        .c(_1464_)
    );

    bfr new_Jinkela_buffer_16251 (
        .din(new_Jinkela_wire_19413),
        .dout(new_Jinkela_wire_19414)
    );

    and_bb _2429_ (
        .a(new_Jinkela_wire_356),
        .b(new_Jinkela_wire_255),
        .c(_1465_)
    );

    bfr new_Jinkela_buffer_12791 (
        .din(new_Jinkela_wire_15312),
        .dout(new_Jinkela_wire_15313)
    );

    bfr new_Jinkela_buffer_16315 (
        .din(new_Jinkela_wire_19481),
        .dout(new_Jinkela_wire_19482)
    );

    and_bi _2430_ (
        .a(new_Jinkela_wire_14324),
        .b(new_Jinkela_wire_4329),
        .c(_1466_)
    );

    bfr new_Jinkela_buffer_12918 (
        .din(new_Jinkela_wire_15439),
        .dout(new_Jinkela_wire_15440)
    );

    bfr new_Jinkela_buffer_16252 (
        .din(new_Jinkela_wire_19414),
        .dout(new_Jinkela_wire_19415)
    );

    and_bb _2431_ (
        .a(new_Jinkela_wire_698),
        .b(new_Jinkela_wire_296),
        .c(_1467_)
    );

    bfr new_Jinkela_buffer_12792 (
        .din(new_Jinkela_wire_15313),
        .dout(new_Jinkela_wire_15314)
    );

    bfr new_Jinkela_buffer_16372 (
        .din(new_Jinkela_wire_19550),
        .dout(new_Jinkela_wire_19551)
    );

    and_bi _2432_ (
        .a(new_Jinkela_wire_1770),
        .b(new_Jinkela_wire_15520),
        .c(_1468_)
    );

    spl2 new_Jinkela_splitter_1120 (
        .a(_1384_),
        .b(new_Jinkela_wire_15669),
        .c(new_Jinkela_wire_15670)
    );

    bfr new_Jinkela_buffer_16253 (
        .din(new_Jinkela_wire_19415),
        .dout(new_Jinkela_wire_19416)
    );

    and_bb _2433_ (
        .a(new_Jinkela_wire_65),
        .b(new_Jinkela_wire_489),
        .c(_1470_)
    );

    bfr new_Jinkela_buffer_12793 (
        .din(new_Jinkela_wire_15314),
        .dout(new_Jinkela_wire_15315)
    );

    bfr new_Jinkela_buffer_16316 (
        .din(new_Jinkela_wire_19482),
        .dout(new_Jinkela_wire_19483)
    );

    and_bi _2434_ (
        .a(new_Jinkela_wire_15526),
        .b(new_Jinkela_wire_16515),
        .c(_1471_)
    );

    bfr new_Jinkela_buffer_12968 (
        .din(new_Jinkela_wire_15491),
        .dout(new_Jinkela_wire_15492)
    );

    bfr new_Jinkela_buffer_12919 (
        .din(new_Jinkela_wire_15440),
        .dout(new_Jinkela_wire_15441)
    );

    bfr new_Jinkela_buffer_16254 (
        .din(new_Jinkela_wire_19416),
        .dout(new_Jinkela_wire_19417)
    );

    and_bb _2435_ (
        .a(new_Jinkela_wire_37),
        .b(new_Jinkela_wire_648),
        .c(_1472_)
    );

    bfr new_Jinkela_buffer_12794 (
        .din(new_Jinkela_wire_15315),
        .dout(new_Jinkela_wire_15316)
    );

    and_bi _2436_ (
        .a(new_Jinkela_wire_3885),
        .b(new_Jinkela_wire_4081),
        .c(_1473_)
    );

    spl2 new_Jinkela_splitter_1440 (
        .a(_0914_),
        .b(new_Jinkela_wire_19558),
        .c(new_Jinkela_wire_19559)
    );

    bfr new_Jinkela_buffer_16255 (
        .din(new_Jinkela_wire_19417),
        .dout(new_Jinkela_wire_19418)
    );

    and_bb _2437_ (
        .a(new_Jinkela_wire_189),
        .b(new_Jinkela_wire_635),
        .c(_1474_)
    );

    bfr new_Jinkela_buffer_12795 (
        .din(new_Jinkela_wire_15316),
        .dout(new_Jinkela_wire_15317)
    );

    bfr new_Jinkela_buffer_16317 (
        .din(new_Jinkela_wire_19483),
        .dout(new_Jinkela_wire_19484)
    );

    and_bi _2438_ (
        .a(new_Jinkela_wire_5166),
        .b(new_Jinkela_wire_6858),
        .c(_1475_)
    );

    bfr new_Jinkela_buffer_12920 (
        .din(new_Jinkela_wire_15441),
        .dout(new_Jinkela_wire_15442)
    );

    bfr new_Jinkela_buffer_16256 (
        .din(new_Jinkela_wire_19418),
        .dout(new_Jinkela_wire_19419)
    );

    and_bb _2439_ (
        .a(new_Jinkela_wire_381),
        .b(new_Jinkela_wire_548),
        .c(_1476_)
    );

    bfr new_Jinkela_buffer_12796 (
        .din(new_Jinkela_wire_15317),
        .dout(new_Jinkela_wire_15318)
    );

    bfr new_Jinkela_buffer_16373 (
        .din(new_Jinkela_wire_19551),
        .dout(new_Jinkela_wire_19552)
    );

    or_ii _2440_ (
        .a(new_Jinkela_wire_162),
        .b(new_Jinkela_wire_315),
        .c(_1477_)
    );

    bfr new_Jinkela_buffer_13005 (
        .din(new_Jinkela_wire_15534),
        .dout(new_Jinkela_wire_15535)
    );

    bfr new_Jinkela_buffer_16257 (
        .din(new_Jinkela_wire_19419),
        .dout(new_Jinkela_wire_19420)
    );

    and_bi _2441_ (
        .a(new_Jinkela_wire_15670),
        .b(new_Jinkela_wire_17087),
        .c(_1478_)
    );

    bfr new_Jinkela_buffer_12797 (
        .din(new_Jinkela_wire_15318),
        .dout(new_Jinkela_wire_15319)
    );

    bfr new_Jinkela_buffer_16318 (
        .din(new_Jinkela_wire_19484),
        .dout(new_Jinkela_wire_19485)
    );

    or_ii _2442_ (
        .a(new_Jinkela_wire_163),
        .b(new_Jinkela_wire_240),
        .c(_1479_)
    );

    bfr new_Jinkela_buffer_12969 (
        .din(new_Jinkela_wire_15492),
        .dout(new_Jinkela_wire_15493)
    );

    bfr new_Jinkela_buffer_12921 (
        .din(new_Jinkela_wire_15442),
        .dout(new_Jinkela_wire_15443)
    );

    bfr new_Jinkela_buffer_16258 (
        .din(new_Jinkela_wire_19420),
        .dout(new_Jinkela_wire_19421)
    );

    and_bb _2443_ (
        .a(new_Jinkela_wire_19540),
        .b(new_Jinkela_wire_4832),
        .c(_1481_)
    );

    bfr new_Jinkela_buffer_12798 (
        .din(new_Jinkela_wire_15319),
        .dout(new_Jinkela_wire_15320)
    );

    bfr new_Jinkela_buffer_16375 (
        .din(new_Jinkela_wire_19561),
        .dout(new_Jinkela_wire_19562)
    );

    and_ii _2444_ (
        .a(new_Jinkela_wire_8866),
        .b(new_Jinkela_wire_19925),
        .c(_1482_)
    );

    spl2 new_Jinkela_splitter_1441 (
        .a(_0193_),
        .b(new_Jinkela_wire_19560),
        .c(new_Jinkela_wire_19561)
    );

    bfr new_Jinkela_buffer_16259 (
        .din(new_Jinkela_wire_19421),
        .dout(new_Jinkela_wire_19422)
    );

    or_bb _2445_ (
        .a(new_Jinkela_wire_718),
        .b(new_Jinkela_wire_9015),
        .c(_1483_)
    );

    bfr new_Jinkela_buffer_12799 (
        .din(new_Jinkela_wire_15320),
        .dout(new_Jinkela_wire_15321)
    );

    bfr new_Jinkela_buffer_16319 (
        .din(new_Jinkela_wire_19485),
        .dout(new_Jinkela_wire_19486)
    );

    or_ii _2446_ (
        .a(new_Jinkela_wire_719),
        .b(new_Jinkela_wire_9016),
        .c(_1484_)
    );

    bfr new_Jinkela_buffer_12922 (
        .din(new_Jinkela_wire_15443),
        .dout(new_Jinkela_wire_15444)
    );

    bfr new_Jinkela_buffer_16260 (
        .din(new_Jinkela_wire_19422),
        .dout(new_Jinkela_wire_19423)
    );

    or_ii _2447_ (
        .a(new_Jinkela_wire_21199),
        .b(new_Jinkela_wire_18763),
        .c(_1485_)
    );

    bfr new_Jinkela_buffer_12800 (
        .din(new_Jinkela_wire_15321),
        .dout(new_Jinkela_wire_15322)
    );

    bfr new_Jinkela_buffer_16374 (
        .din(new_Jinkela_wire_19552),
        .dout(new_Jinkela_wire_19553)
    );

    and_ii _2448_ (
        .a(new_Jinkela_wire_5714),
        .b(new_Jinkela_wire_2340),
        .c(_1486_)
    );

    bfr new_Jinkela_buffer_13025 (
        .din(new_Jinkela_wire_15558),
        .dout(new_Jinkela_wire_15559)
    );

    bfr new_Jinkela_buffer_16261 (
        .din(new_Jinkela_wire_19423),
        .dout(new_Jinkela_wire_19424)
    );

    and_bb _2449_ (
        .a(new_Jinkela_wire_5715),
        .b(new_Jinkela_wire_2341),
        .c(_1487_)
    );

    bfr new_Jinkela_buffer_12801 (
        .din(new_Jinkela_wire_15322),
        .dout(new_Jinkela_wire_15323)
    );

    bfr new_Jinkela_buffer_16320 (
        .din(new_Jinkela_wire_19486),
        .dout(new_Jinkela_wire_19487)
    );

    or_bb _2450_ (
        .a(new_Jinkela_wire_16511),
        .b(new_Jinkela_wire_19156),
        .c(_1488_)
    );

    bfr new_Jinkela_buffer_12970 (
        .din(new_Jinkela_wire_15493),
        .dout(new_Jinkela_wire_15494)
    );

    bfr new_Jinkela_buffer_12923 (
        .din(new_Jinkela_wire_15444),
        .dout(new_Jinkela_wire_15445)
    );

    bfr new_Jinkela_buffer_16262 (
        .din(new_Jinkela_wire_19424),
        .dout(new_Jinkela_wire_19425)
    );

    or_bb _2451_ (
        .a(new_Jinkela_wire_7128),
        .b(new_Jinkela_wire_7693),
        .c(_1489_)
    );

    bfr new_Jinkela_buffer_12802 (
        .din(new_Jinkela_wire_15323),
        .dout(new_Jinkela_wire_15324)
    );

    or_ii _2452_ (
        .a(new_Jinkela_wire_7129),
        .b(new_Jinkela_wire_7694),
        .c(_1490_)
    );

    bfr new_Jinkela_buffer_16379 (
        .din(_1779_),
        .dout(new_Jinkela_wire_19566)
    );

    bfr new_Jinkela_buffer_16263 (
        .din(new_Jinkela_wire_19425),
        .dout(new_Jinkela_wire_19426)
    );

    or_ii _2453_ (
        .a(new_Jinkela_wire_14016),
        .b(new_Jinkela_wire_18791),
        .c(_1492_)
    );

    bfr new_Jinkela_buffer_12803 (
        .din(new_Jinkela_wire_15324),
        .dout(new_Jinkela_wire_15325)
    );

    bfr new_Jinkela_buffer_16321 (
        .din(new_Jinkela_wire_19487),
        .dout(new_Jinkela_wire_19488)
    );

    and_ii _2454_ (
        .a(new_Jinkela_wire_13203),
        .b(new_Jinkela_wire_11038),
        .c(_1493_)
    );

    bfr new_Jinkela_buffer_2359 (
        .din(new_Jinkela_wire_3346),
        .dout(new_Jinkela_wire_3347)
    );

    bfr new_Jinkela_buffer_2418 (
        .din(new_Jinkela_wire_3411),
        .dout(new_Jinkela_wire_3412)
    );

    bfr new_Jinkela_buffer_2360 (
        .din(new_Jinkela_wire_3347),
        .dout(new_Jinkela_wire_3348)
    );

    bfr new_Jinkela_buffer_2445 (
        .din(new_Jinkela_wire_3454),
        .dout(new_Jinkela_wire_3455)
    );

    bfr new_Jinkela_buffer_2361 (
        .din(new_Jinkela_wire_3348),
        .dout(new_Jinkela_wire_3349)
    );

    bfr new_Jinkela_buffer_2419 (
        .din(new_Jinkela_wire_3412),
        .dout(new_Jinkela_wire_3413)
    );

    bfr new_Jinkela_buffer_2362 (
        .din(new_Jinkela_wire_3349),
        .dout(new_Jinkela_wire_3350)
    );

    spl2 new_Jinkela_splitter_358 (
        .a(_0652_),
        .b(new_Jinkela_wire_3555),
        .c(new_Jinkela_wire_3556)
    );

    bfr new_Jinkela_buffer_2676 (
        .din(_0176_),
        .dout(new_Jinkela_wire_3720)
    );

    bfr new_Jinkela_buffer_2363 (
        .din(new_Jinkela_wire_3350),
        .dout(new_Jinkela_wire_3351)
    );

    bfr new_Jinkela_buffer_2420 (
        .din(new_Jinkela_wire_3413),
        .dout(new_Jinkela_wire_3414)
    );

    bfr new_Jinkela_buffer_2364 (
        .din(new_Jinkela_wire_3351),
        .dout(new_Jinkela_wire_3352)
    );

    bfr new_Jinkela_buffer_2446 (
        .din(new_Jinkela_wire_3455),
        .dout(new_Jinkela_wire_3456)
    );

    bfr new_Jinkela_buffer_2365 (
        .din(new_Jinkela_wire_3352),
        .dout(new_Jinkela_wire_3353)
    );

    bfr new_Jinkela_buffer_2421 (
        .din(new_Jinkela_wire_3414),
        .dout(new_Jinkela_wire_3415)
    );

    bfr new_Jinkela_buffer_2366 (
        .din(new_Jinkela_wire_3353),
        .dout(new_Jinkela_wire_3354)
    );

    bfr new_Jinkela_buffer_2474 (
        .din(new_Jinkela_wire_3487),
        .dout(new_Jinkela_wire_3488)
    );

    bfr new_Jinkela_buffer_2367 (
        .din(new_Jinkela_wire_3354),
        .dout(new_Jinkela_wire_3355)
    );

    bfr new_Jinkela_buffer_2422 (
        .din(new_Jinkela_wire_3415),
        .dout(new_Jinkela_wire_3416)
    );

    bfr new_Jinkela_buffer_2368 (
        .din(new_Jinkela_wire_3355),
        .dout(new_Jinkela_wire_3356)
    );

    bfr new_Jinkela_buffer_2447 (
        .din(new_Jinkela_wire_3456),
        .dout(new_Jinkela_wire_3457)
    );

    bfr new_Jinkela_buffer_2369 (
        .din(new_Jinkela_wire_3356),
        .dout(new_Jinkela_wire_3357)
    );

    bfr new_Jinkela_buffer_2423 (
        .din(new_Jinkela_wire_3416),
        .dout(new_Jinkela_wire_3417)
    );

    bfr new_Jinkela_buffer_2370 (
        .din(new_Jinkela_wire_3357),
        .dout(new_Jinkela_wire_3358)
    );

    bfr new_Jinkela_buffer_2563 (
        .din(new_Jinkela_wire_3582),
        .dout(new_Jinkela_wire_3583)
    );

    spl2 new_Jinkela_splitter_343 (
        .a(new_Jinkela_wire_3358),
        .b(new_Jinkela_wire_3359),
        .c(new_Jinkela_wire_3360)
    );

    bfr new_Jinkela_buffer_2448 (
        .din(new_Jinkela_wire_3457),
        .dout(new_Jinkela_wire_3458)
    );

    bfr new_Jinkela_buffer_2424 (
        .din(new_Jinkela_wire_3417),
        .dout(new_Jinkela_wire_3418)
    );

    bfr new_Jinkela_buffer_2425 (
        .din(new_Jinkela_wire_3418),
        .dout(new_Jinkela_wire_3419)
    );

    bfr new_Jinkela_buffer_2475 (
        .din(new_Jinkela_wire_3488),
        .dout(new_Jinkela_wire_3489)
    );

    bfr new_Jinkela_buffer_2426 (
        .din(new_Jinkela_wire_3419),
        .dout(new_Jinkela_wire_3420)
    );

    bfr new_Jinkela_buffer_2449 (
        .din(new_Jinkela_wire_3458),
        .dout(new_Jinkela_wire_3459)
    );

    bfr new_Jinkela_buffer_2427 (
        .din(new_Jinkela_wire_3420),
        .dout(new_Jinkela_wire_3421)
    );

    bfr new_Jinkela_buffer_2428 (
        .din(new_Jinkela_wire_3421),
        .dout(new_Jinkela_wire_3422)
    );

    bfr new_Jinkela_buffer_2450 (
        .din(new_Jinkela_wire_3459),
        .dout(new_Jinkela_wire_3460)
    );

    bfr new_Jinkela_buffer_2429 (
        .din(new_Jinkela_wire_3422),
        .dout(new_Jinkela_wire_3423)
    );

    bfr new_Jinkela_buffer_2476 (
        .din(new_Jinkela_wire_3489),
        .dout(new_Jinkela_wire_3490)
    );

    bfr new_Jinkela_buffer_2430 (
        .din(new_Jinkela_wire_3423),
        .dout(new_Jinkela_wire_3424)
    );

    bfr new_Jinkela_buffer_2451 (
        .din(new_Jinkela_wire_3460),
        .dout(new_Jinkela_wire_3461)
    );

    bfr new_Jinkela_buffer_2431 (
        .din(new_Jinkela_wire_3424),
        .dout(new_Jinkela_wire_3425)
    );

    bfr new_Jinkela_buffer_2432 (
        .din(new_Jinkela_wire_3425),
        .dout(new_Jinkela_wire_3426)
    );

    bfr new_Jinkela_buffer_5845 (
        .din(new_Jinkela_wire_7434),
        .dout(new_Jinkela_wire_7435)
    );

    bfr new_Jinkela_buffer_5982 (
        .din(new_Jinkela_wire_7597),
        .dout(new_Jinkela_wire_7598)
    );

    bfr new_Jinkela_buffer_5846 (
        .din(new_Jinkela_wire_7435),
        .dout(new_Jinkela_wire_7436)
    );

    bfr new_Jinkela_buffer_5929 (
        .din(new_Jinkela_wire_7536),
        .dout(new_Jinkela_wire_7537)
    );

    bfr new_Jinkela_buffer_5847 (
        .din(new_Jinkela_wire_7436),
        .dout(new_Jinkela_wire_7437)
    );

    spl2 new_Jinkela_splitter_644 (
        .a(new_Jinkela_wire_7437),
        .b(new_Jinkela_wire_7438),
        .c(new_Jinkela_wire_7439)
    );

    bfr new_Jinkela_buffer_5983 (
        .din(new_Jinkela_wire_7598),
        .dout(new_Jinkela_wire_7599)
    );

    bfr new_Jinkela_buffer_5930 (
        .din(new_Jinkela_wire_7537),
        .dout(new_Jinkela_wire_7538)
    );

    bfr new_Jinkela_buffer_5931 (
        .din(new_Jinkela_wire_7538),
        .dout(new_Jinkela_wire_7539)
    );

    bfr new_Jinkela_buffer_6075 (
        .din(new_Jinkela_wire_7698),
        .dout(new_Jinkela_wire_7699)
    );

    bfr new_Jinkela_buffer_5932 (
        .din(new_Jinkela_wire_7539),
        .dout(new_Jinkela_wire_7540)
    );

    bfr new_Jinkela_buffer_5984 (
        .din(new_Jinkela_wire_7599),
        .dout(new_Jinkela_wire_7600)
    );

    bfr new_Jinkela_buffer_5933 (
        .din(new_Jinkela_wire_7540),
        .dout(new_Jinkela_wire_7541)
    );

    spl2 new_Jinkela_splitter_665 (
        .a(_1455_),
        .b(new_Jinkela_wire_7710),
        .c(new_Jinkela_wire_7711)
    );

    bfr new_Jinkela_buffer_5934 (
        .din(new_Jinkela_wire_7541),
        .dout(new_Jinkela_wire_7542)
    );

    bfr new_Jinkela_buffer_5985 (
        .din(new_Jinkela_wire_7600),
        .dout(new_Jinkela_wire_7601)
    );

    bfr new_Jinkela_buffer_5935 (
        .din(new_Jinkela_wire_7542),
        .dout(new_Jinkela_wire_7543)
    );

    bfr new_Jinkela_buffer_6076 (
        .din(new_Jinkela_wire_7699),
        .dout(new_Jinkela_wire_7700)
    );

    bfr new_Jinkela_buffer_5936 (
        .din(new_Jinkela_wire_7543),
        .dout(new_Jinkela_wire_7544)
    );

    bfr new_Jinkela_buffer_5986 (
        .din(new_Jinkela_wire_7601),
        .dout(new_Jinkela_wire_7602)
    );

    bfr new_Jinkela_buffer_5937 (
        .din(new_Jinkela_wire_7544),
        .dout(new_Jinkela_wire_7545)
    );

    bfr new_Jinkela_buffer_6077 (
        .din(new_Jinkela_wire_7706),
        .dout(new_Jinkela_wire_7707)
    );

    spl2 new_Jinkela_splitter_666 (
        .a(_0196_),
        .b(new_Jinkela_wire_7712),
        .c(new_Jinkela_wire_7713)
    );

    bfr new_Jinkela_buffer_5938 (
        .din(new_Jinkela_wire_7545),
        .dout(new_Jinkela_wire_7546)
    );

    bfr new_Jinkela_buffer_5987 (
        .din(new_Jinkela_wire_7602),
        .dout(new_Jinkela_wire_7603)
    );

    bfr new_Jinkela_buffer_5939 (
        .din(new_Jinkela_wire_7546),
        .dout(new_Jinkela_wire_7547)
    );

    bfr new_Jinkela_buffer_6078 (
        .din(_1223_),
        .dout(new_Jinkela_wire_7714)
    );

    bfr new_Jinkela_buffer_5940 (
        .din(new_Jinkela_wire_7547),
        .dout(new_Jinkela_wire_7548)
    );

    bfr new_Jinkela_buffer_5988 (
        .din(new_Jinkela_wire_7603),
        .dout(new_Jinkela_wire_7604)
    );

    bfr new_Jinkela_buffer_5941 (
        .din(new_Jinkela_wire_7548),
        .dout(new_Jinkela_wire_7549)
    );

    spl2 new_Jinkela_splitter_664 (
        .a(new_Jinkela_wire_7707),
        .b(new_Jinkela_wire_7708),
        .c(new_Jinkela_wire_7709)
    );

    bfr new_Jinkela_buffer_5942 (
        .din(new_Jinkela_wire_7549),
        .dout(new_Jinkela_wire_7550)
    );

    bfr new_Jinkela_buffer_5989 (
        .din(new_Jinkela_wire_7604),
        .dout(new_Jinkela_wire_7605)
    );

    bfr new_Jinkela_buffer_5943 (
        .din(new_Jinkela_wire_7550),
        .dout(new_Jinkela_wire_7551)
    );

    bfr new_Jinkela_buffer_6079 (
        .din(_1394_),
        .dout(new_Jinkela_wire_7717)
    );

    bfr new_Jinkela_buffer_5944 (
        .din(new_Jinkela_wire_7551),
        .dout(new_Jinkela_wire_7552)
    );

    bfr new_Jinkela_buffer_5990 (
        .din(new_Jinkela_wire_7605),
        .dout(new_Jinkela_wire_7606)
    );

    bfr new_Jinkela_buffer_5945 (
        .din(new_Jinkela_wire_7552),
        .dout(new_Jinkela_wire_7553)
    );

    spl2 new_Jinkela_splitter_667 (
        .a(_0777_),
        .b(new_Jinkela_wire_7715),
        .c(new_Jinkela_wire_7716)
    );

    bfr new_Jinkela_buffer_5946 (
        .din(new_Jinkela_wire_7553),
        .dout(new_Jinkela_wire_7554)
    );

    bfr new_Jinkela_buffer_5991 (
        .din(new_Jinkela_wire_7606),
        .dout(new_Jinkela_wire_7607)
    );

    bfr new_Jinkela_buffer_5947 (
        .din(new_Jinkela_wire_7554),
        .dout(new_Jinkela_wire_7555)
    );

    bfr new_Jinkela_buffer_12924 (
        .din(new_Jinkela_wire_15445),
        .dout(new_Jinkela_wire_15446)
    );

    bfr new_Jinkela_buffer_12804 (
        .din(new_Jinkela_wire_15325),
        .dout(new_Jinkela_wire_15326)
    );

    bfr new_Jinkela_buffer_13006 (
        .din(new_Jinkela_wire_15535),
        .dout(new_Jinkela_wire_15536)
    );

    bfr new_Jinkela_buffer_12805 (
        .din(new_Jinkela_wire_15326),
        .dout(new_Jinkela_wire_15327)
    );

    bfr new_Jinkela_buffer_12971 (
        .din(new_Jinkela_wire_15494),
        .dout(new_Jinkela_wire_15495)
    );

    bfr new_Jinkela_buffer_12925 (
        .din(new_Jinkela_wire_15446),
        .dout(new_Jinkela_wire_15447)
    );

    bfr new_Jinkela_buffer_12806 (
        .din(new_Jinkela_wire_15327),
        .dout(new_Jinkela_wire_15328)
    );

    bfr new_Jinkela_buffer_12807 (
        .din(new_Jinkela_wire_15328),
        .dout(new_Jinkela_wire_15329)
    );

    bfr new_Jinkela_buffer_12926 (
        .din(new_Jinkela_wire_15447),
        .dout(new_Jinkela_wire_15448)
    );

    bfr new_Jinkela_buffer_12808 (
        .din(new_Jinkela_wire_15329),
        .dout(new_Jinkela_wire_15330)
    );

    bfr new_Jinkela_buffer_12809 (
        .din(new_Jinkela_wire_15330),
        .dout(new_Jinkela_wire_15331)
    );

    bfr new_Jinkela_buffer_12972 (
        .din(new_Jinkela_wire_15495),
        .dout(new_Jinkela_wire_15496)
    );

    bfr new_Jinkela_buffer_12927 (
        .din(new_Jinkela_wire_15448),
        .dout(new_Jinkela_wire_15449)
    );

    bfr new_Jinkela_buffer_12810 (
        .din(new_Jinkela_wire_15331),
        .dout(new_Jinkela_wire_15332)
    );

    bfr new_Jinkela_buffer_12811 (
        .din(new_Jinkela_wire_15332),
        .dout(new_Jinkela_wire_15333)
    );

    spl2 new_Jinkela_splitter_1119 (
        .a(_0101_),
        .b(new_Jinkela_wire_15667),
        .c(new_Jinkela_wire_15668)
    );

    bfr new_Jinkela_buffer_12928 (
        .din(new_Jinkela_wire_15449),
        .dout(new_Jinkela_wire_15450)
    );

    bfr new_Jinkela_buffer_12812 (
        .din(new_Jinkela_wire_15333),
        .dout(new_Jinkela_wire_15334)
    );

    bfr new_Jinkela_buffer_13007 (
        .din(new_Jinkela_wire_15536),
        .dout(new_Jinkela_wire_15537)
    );

    bfr new_Jinkela_buffer_12813 (
        .din(new_Jinkela_wire_15334),
        .dout(new_Jinkela_wire_15335)
    );

    bfr new_Jinkela_buffer_12973 (
        .din(new_Jinkela_wire_15496),
        .dout(new_Jinkela_wire_15497)
    );

    bfr new_Jinkela_buffer_12929 (
        .din(new_Jinkela_wire_15450),
        .dout(new_Jinkela_wire_15451)
    );

    bfr new_Jinkela_buffer_12814 (
        .din(new_Jinkela_wire_15335),
        .dout(new_Jinkela_wire_15336)
    );

    bfr new_Jinkela_buffer_12815 (
        .din(new_Jinkela_wire_15336),
        .dout(new_Jinkela_wire_15337)
    );

    bfr new_Jinkela_buffer_12930 (
        .din(new_Jinkela_wire_15451),
        .dout(new_Jinkela_wire_15452)
    );

    bfr new_Jinkela_buffer_12816 (
        .din(new_Jinkela_wire_15337),
        .dout(new_Jinkela_wire_15338)
    );

    bfr new_Jinkela_buffer_13026 (
        .din(new_Jinkela_wire_15559),
        .dout(new_Jinkela_wire_15560)
    );

    bfr new_Jinkela_buffer_12817 (
        .din(new_Jinkela_wire_15338),
        .dout(new_Jinkela_wire_15339)
    );

    bfr new_Jinkela_buffer_12974 (
        .din(new_Jinkela_wire_15497),
        .dout(new_Jinkela_wire_15498)
    );

    bfr new_Jinkela_buffer_12931 (
        .din(new_Jinkela_wire_15452),
        .dout(new_Jinkela_wire_15453)
    );

    bfr new_Jinkela_buffer_12818 (
        .din(new_Jinkela_wire_15339),
        .dout(new_Jinkela_wire_15340)
    );

    bfr new_Jinkela_buffer_12819 (
        .din(new_Jinkela_wire_15340),
        .dout(new_Jinkela_wire_15341)
    );

    bfr new_Jinkela_buffer_12932 (
        .din(new_Jinkela_wire_15453),
        .dout(new_Jinkela_wire_15454)
    );

    bfr new_Jinkela_buffer_12820 (
        .din(new_Jinkela_wire_15341),
        .dout(new_Jinkela_wire_15342)
    );

    bfr new_Jinkela_buffer_13008 (
        .din(new_Jinkela_wire_15537),
        .dout(new_Jinkela_wire_15538)
    );

    bfr new_Jinkela_buffer_12821 (
        .din(new_Jinkela_wire_15342),
        .dout(new_Jinkela_wire_15343)
    );

    bfr new_Jinkela_buffer_12975 (
        .din(new_Jinkela_wire_15498),
        .dout(new_Jinkela_wire_15499)
    );

    bfr new_Jinkela_buffer_12933 (
        .din(new_Jinkela_wire_15454),
        .dout(new_Jinkela_wire_15455)
    );

    bfr new_Jinkela_buffer_12822 (
        .din(new_Jinkela_wire_15343),
        .dout(new_Jinkela_wire_15344)
    );

    bfr new_Jinkela_buffer_12823 (
        .din(new_Jinkela_wire_15344),
        .dout(new_Jinkela_wire_15345)
    );

    bfr new_Jinkela_buffer_12934 (
        .din(new_Jinkela_wire_15455),
        .dout(new_Jinkela_wire_15456)
    );

    bfr new_Jinkela_buffer_12824 (
        .din(new_Jinkela_wire_15345),
        .dout(new_Jinkela_wire_15346)
    );

    and_bb _3340_ (
        .a(new_Jinkela_wire_503),
        .b(new_Jinkela_wire_516),
        .c(_0619_)
    );

    bfr new_Jinkela_buffer_16264 (
        .din(new_Jinkela_wire_19426),
        .dout(new_Jinkela_wire_19427)
    );

    and_ii _3341_ (
        .a(new_Jinkela_wire_13684),
        .b(new_Jinkela_wire_10579),
        .c(_0620_)
    );

    spl2 new_Jinkela_splitter_1442 (
        .a(_0070_),
        .b(new_Jinkela_wire_19567),
        .c(new_Jinkela_wire_19568)
    );

    and_bb _3342_ (
        .a(new_Jinkela_wire_143),
        .b(new_Jinkela_wire_35),
        .c(_0621_)
    );

    bfr new_Jinkela_buffer_16265 (
        .din(new_Jinkela_wire_19427),
        .dout(new_Jinkela_wire_19428)
    );

    and_ii _3343_ (
        .a(new_Jinkela_wire_4679),
        .b(new_Jinkela_wire_9106),
        .c(_0622_)
    );

    bfr new_Jinkela_buffer_16322 (
        .din(new_Jinkela_wire_19488),
        .dout(new_Jinkela_wire_19489)
    );

    and_bb _3344_ (
        .a(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_203),
        .c(_0623_)
    );

    bfr new_Jinkela_buffer_16266 (
        .din(new_Jinkela_wire_19428),
        .dout(new_Jinkela_wire_19429)
    );

    and_ii _3345_ (
        .a(new_Jinkela_wire_6410),
        .b(new_Jinkela_wire_4482),
        .c(_0624_)
    );

    bfr new_Jinkela_buffer_16380 (
        .din(new_net_3928),
        .dout(new_Jinkela_wire_19569)
    );

    bfr new_Jinkela_buffer_16540 (
        .din(_0754_),
        .dout(new_Jinkela_wire_19731)
    );

    and_bb _3346_ (
        .a(new_Jinkela_wire_392),
        .b(new_Jinkela_wire_590),
        .c(_0625_)
    );

    bfr new_Jinkela_buffer_16267 (
        .din(new_Jinkela_wire_19429),
        .dout(new_Jinkela_wire_19430)
    );

    and_ii _3347_ (
        .a(new_Jinkela_wire_8590),
        .b(new_Jinkela_wire_6690),
        .c(_0626_)
    );

    bfr new_Jinkela_buffer_16323 (
        .din(new_Jinkela_wire_19489),
        .dout(new_Jinkela_wire_19490)
    );

    and_bb _3348_ (
        .a(new_Jinkela_wire_396),
        .b(new_Jinkela_wire_126),
        .c(_0627_)
    );

    bfr new_Jinkela_buffer_16268 (
        .din(new_Jinkela_wire_19430),
        .dout(new_Jinkela_wire_19431)
    );

    and_ii _3349_ (
        .a(new_Jinkela_wire_2944),
        .b(new_Jinkela_wire_16211),
        .c(_0628_)
    );

    bfr new_Jinkela_buffer_16376 (
        .din(new_Jinkela_wire_19562),
        .dout(new_Jinkela_wire_19563)
    );

    and_bb _3350_ (
        .a(new_Jinkela_wire_169),
        .b(new_Jinkela_wire_4),
        .c(_0629_)
    );

    bfr new_Jinkela_buffer_16269 (
        .din(new_Jinkela_wire_19431),
        .dout(new_Jinkela_wire_19432)
    );

    and_ii _3351_ (
        .a(new_Jinkela_wire_18118),
        .b(new_Jinkela_wire_5453),
        .c(_0630_)
    );

    bfr new_Jinkela_buffer_16324 (
        .din(new_Jinkela_wire_19490),
        .dout(new_Jinkela_wire_19491)
    );

    and_bb _3352_ (
        .a(new_Jinkela_wire_597),
        .b(new_Jinkela_wire_464),
        .c(_0631_)
    );

    bfr new_Jinkela_buffer_16270 (
        .din(new_Jinkela_wire_19432),
        .dout(new_Jinkela_wire_19433)
    );

    and_bb _3353_ (
        .a(new_Jinkela_wire_435),
        .b(new_Jinkela_wire_260),
        .c(_0634_)
    );

    bfr new_Jinkela_buffer_16381 (
        .din(new_Jinkela_wire_19569),
        .dout(new_Jinkela_wire_19570)
    );

    and_ii _3354_ (
        .a(new_Jinkela_wire_15518),
        .b(new_Jinkela_wire_14306),
        .c(_0635_)
    );

    bfr new_Jinkela_buffer_16271 (
        .din(new_Jinkela_wire_19433),
        .dout(new_Jinkela_wire_19434)
    );

    and_ii _3355_ (
        .a(new_Jinkela_wire_5988),
        .b(new_Jinkela_wire_20624),
        .c(_0636_)
    );

    bfr new_Jinkela_buffer_16325 (
        .din(new_Jinkela_wire_19491),
        .dout(new_Jinkela_wire_19492)
    );

    and_bb _3356_ (
        .a(new_Jinkela_wire_5989),
        .b(new_Jinkela_wire_20625),
        .c(_0637_)
    );

    bfr new_Jinkela_buffer_16272 (
        .din(new_Jinkela_wire_19434),
        .dout(new_Jinkela_wire_19435)
    );

    or_bb _3357_ (
        .a(new_Jinkela_wire_21116),
        .b(new_Jinkela_wire_14038),
        .c(_0638_)
    );

    bfr new_Jinkela_buffer_16377 (
        .din(new_Jinkela_wire_19563),
        .dout(new_Jinkela_wire_19564)
    );

    and_ii _3358_ (
        .a(new_Jinkela_wire_4899),
        .b(new_Jinkela_wire_20958),
        .c(_0639_)
    );

    bfr new_Jinkela_buffer_16273 (
        .din(new_Jinkela_wire_19435),
        .dout(new_Jinkela_wire_19436)
    );

    and_bb _3359_ (
        .a(new_Jinkela_wire_4900),
        .b(new_Jinkela_wire_20959),
        .c(_0640_)
    );

    bfr new_Jinkela_buffer_16326 (
        .din(new_Jinkela_wire_19492),
        .dout(new_Jinkela_wire_19493)
    );

    or_bb _3360_ (
        .a(new_Jinkela_wire_13341),
        .b(new_Jinkela_wire_20362),
        .c(_0641_)
    );

    bfr new_Jinkela_buffer_16274 (
        .din(new_Jinkela_wire_19436),
        .dout(new_Jinkela_wire_19437)
    );

    and_ii _3361_ (
        .a(new_Jinkela_wire_10967),
        .b(new_Jinkela_wire_8183),
        .c(_0642_)
    );

    spl2 new_Jinkela_splitter_1443 (
        .a(_0953_),
        .b(new_Jinkela_wire_19685),
        .c(new_Jinkela_wire_19686)
    );

    and_bb _3362_ (
        .a(new_Jinkela_wire_10968),
        .b(new_Jinkela_wire_8184),
        .c(_0643_)
    );

    bfr new_Jinkela_buffer_16275 (
        .din(new_Jinkela_wire_19437),
        .dout(new_Jinkela_wire_19438)
    );

    or_bb _3363_ (
        .a(new_Jinkela_wire_13461),
        .b(new_Jinkela_wire_20136),
        .c(_0645_)
    );

    bfr new_Jinkela_buffer_16327 (
        .din(new_Jinkela_wire_19493),
        .dout(new_Jinkela_wire_19494)
    );

    and_ii _3364_ (
        .a(new_Jinkela_wire_17554),
        .b(new_Jinkela_wire_19043),
        .c(_0646_)
    );

    bfr new_Jinkela_buffer_16276 (
        .din(new_Jinkela_wire_19438),
        .dout(new_Jinkela_wire_19439)
    );

    and_bb _3365_ (
        .a(new_Jinkela_wire_17555),
        .b(new_Jinkela_wire_19044),
        .c(_0647_)
    );

    bfr new_Jinkela_buffer_16378 (
        .din(new_Jinkela_wire_19564),
        .dout(new_Jinkela_wire_19565)
    );

    or_bb _3366_ (
        .a(new_Jinkela_wire_4483),
        .b(new_Jinkela_wire_6682),
        .c(_0648_)
    );

    bfr new_Jinkela_buffer_16277 (
        .din(new_Jinkela_wire_19439),
        .dout(new_Jinkela_wire_19440)
    );

    and_ii _3367_ (
        .a(new_Jinkela_wire_13982),
        .b(new_Jinkela_wire_14007),
        .c(_0649_)
    );

    bfr new_Jinkela_buffer_16328 (
        .din(new_Jinkela_wire_19494),
        .dout(new_Jinkela_wire_19495)
    );

    and_bb _3368_ (
        .a(new_Jinkela_wire_13983),
        .b(new_Jinkela_wire_14008),
        .c(_0650_)
    );

    bfr new_Jinkela_buffer_16278 (
        .din(new_Jinkela_wire_19440),
        .dout(new_Jinkela_wire_19441)
    );

    or_bb _3369_ (
        .a(new_Jinkela_wire_16872),
        .b(new_Jinkela_wire_18955),
        .c(_0651_)
    );

    bfr new_Jinkela_buffer_16496 (
        .din(new_Jinkela_wire_19686),
        .dout(new_Jinkela_wire_19687)
    );

    and_ii _3370_ (
        .a(new_Jinkela_wire_19962),
        .b(new_Jinkela_wire_7126),
        .c(_0652_)
    );

    bfr new_Jinkela_buffer_16279 (
        .din(new_Jinkela_wire_19441),
        .dout(new_Jinkela_wire_19442)
    );

    and_bb _3371_ (
        .a(new_Jinkela_wire_19963),
        .b(new_Jinkela_wire_7127),
        .c(_0653_)
    );

    bfr new_Jinkela_buffer_16329 (
        .din(new_Jinkela_wire_19495),
        .dout(new_Jinkela_wire_19496)
    );

    or_bb _3372_ (
        .a(new_Jinkela_wire_1781),
        .b(new_Jinkela_wire_3555),
        .c(_0654_)
    );

    bfr new_Jinkela_buffer_16280 (
        .din(new_Jinkela_wire_19442),
        .dout(new_Jinkela_wire_19443)
    );

    and_ii _3373_ (
        .a(new_Jinkela_wire_6374),
        .b(new_Jinkela_wire_13060),
        .c(_0656_)
    );

    bfr new_Jinkela_buffer_16382 (
        .din(new_Jinkela_wire_19570),
        .dout(new_Jinkela_wire_19571)
    );

    and_bb _3374_ (
        .a(new_Jinkela_wire_6375),
        .b(new_Jinkela_wire_13061),
        .c(_0657_)
    );

    bfr new_Jinkela_buffer_16281 (
        .din(new_Jinkela_wire_19443),
        .dout(new_Jinkela_wire_19444)
    );

    or_bb _3375_ (
        .a(new_Jinkela_wire_17864),
        .b(new_Jinkela_wire_5697),
        .c(_0658_)
    );

    bfr new_Jinkela_buffer_16330 (
        .din(new_Jinkela_wire_19496),
        .dout(new_Jinkela_wire_19497)
    );

    and_ii _3376_ (
        .a(new_Jinkela_wire_10116),
        .b(new_Jinkela_wire_15992),
        .c(_0659_)
    );

    bfr new_Jinkela_buffer_16282 (
        .din(new_Jinkela_wire_19444),
        .dout(new_Jinkela_wire_19445)
    );

    and_bb _3377_ (
        .a(new_Jinkela_wire_10117),
        .b(new_Jinkela_wire_15993),
        .c(_0660_)
    );

    or_bb _3378_ (
        .a(new_Jinkela_wire_5135),
        .b(new_Jinkela_wire_12221),
        .c(_0661_)
    );

    bfr new_Jinkela_buffer_16283 (
        .din(new_Jinkela_wire_19445),
        .dout(new_Jinkela_wire_19446)
    );

    and_ii _3379_ (
        .a(new_Jinkela_wire_19061),
        .b(new_Jinkela_wire_4541),
        .c(_0662_)
    );

    bfr new_Jinkela_buffer_16331 (
        .din(new_Jinkela_wire_19497),
        .dout(new_Jinkela_wire_19498)
    );

    and_bb _3380_ (
        .a(new_Jinkela_wire_19062),
        .b(new_Jinkela_wire_4542),
        .c(_0663_)
    );

    bfr new_Jinkela_buffer_16284 (
        .din(new_Jinkela_wire_19446),
        .dout(new_Jinkela_wire_19447)
    );

    or_bb _3381_ (
        .a(new_Jinkela_wire_16970),
        .b(new_Jinkela_wire_6248),
        .c(_0664_)
    );

    bfr new_Jinkela_buffer_16383 (
        .din(new_Jinkela_wire_19571),
        .dout(new_Jinkela_wire_19572)
    );

    bfr new_Jinkela_buffer_2452 (
        .din(new_Jinkela_wire_3461),
        .dout(new_Jinkela_wire_3462)
    );

    spl2 new_Jinkela_splitter_346 (
        .a(new_Jinkela_wire_3426),
        .b(new_Jinkela_wire_3427),
        .c(new_Jinkela_wire_3428)
    );

    bfr new_Jinkela_buffer_2453 (
        .din(new_Jinkela_wire_3462),
        .dout(new_Jinkela_wire_3463)
    );

    bfr new_Jinkela_buffer_2477 (
        .din(new_Jinkela_wire_3490),
        .dout(new_Jinkela_wire_3491)
    );

    spl2 new_Jinkela_splitter_360 (
        .a(_0751_),
        .b(new_Jinkela_wire_3663),
        .c(new_Jinkela_wire_3664)
    );

    bfr new_Jinkela_buffer_2454 (
        .din(new_Jinkela_wire_3463),
        .dout(new_Jinkela_wire_3464)
    );

    bfr new_Jinkela_buffer_2478 (
        .din(new_Jinkela_wire_3491),
        .dout(new_Jinkela_wire_3492)
    );

    bfr new_Jinkela_buffer_2455 (
        .din(new_Jinkela_wire_3464),
        .dout(new_Jinkela_wire_3465)
    );

    spl2 new_Jinkela_splitter_361 (
        .a(_0723_),
        .b(new_Jinkela_wire_3665),
        .c(new_Jinkela_wire_3666)
    );

    bfr new_Jinkela_buffer_2456 (
        .din(new_Jinkela_wire_3465),
        .dout(new_Jinkela_wire_3466)
    );

    bfr new_Jinkela_buffer_2479 (
        .din(new_Jinkela_wire_3492),
        .dout(new_Jinkela_wire_3493)
    );

    bfr new_Jinkela_buffer_2457 (
        .din(new_Jinkela_wire_3466),
        .dout(new_Jinkela_wire_3467)
    );

    bfr new_Jinkela_buffer_2538 (
        .din(new_Jinkela_wire_3557),
        .dout(new_Jinkela_wire_3558)
    );

    bfr new_Jinkela_buffer_2458 (
        .din(new_Jinkela_wire_3467),
        .dout(new_Jinkela_wire_3468)
    );

    bfr new_Jinkela_buffer_2480 (
        .din(new_Jinkela_wire_3493),
        .dout(new_Jinkela_wire_3494)
    );

    bfr new_Jinkela_buffer_2459 (
        .din(new_Jinkela_wire_3468),
        .dout(new_Jinkela_wire_3469)
    );

    bfr new_Jinkela_buffer_2460 (
        .din(new_Jinkela_wire_3469),
        .dout(new_Jinkela_wire_3470)
    );

    bfr new_Jinkela_buffer_2481 (
        .din(new_Jinkela_wire_3494),
        .dout(new_Jinkela_wire_3495)
    );

    bfr new_Jinkela_buffer_2461 (
        .din(new_Jinkela_wire_3470),
        .dout(new_Jinkela_wire_3471)
    );

    bfr new_Jinkela_buffer_2539 (
        .din(new_Jinkela_wire_3558),
        .dout(new_Jinkela_wire_3559)
    );

    bfr new_Jinkela_buffer_2462 (
        .din(new_Jinkela_wire_3471),
        .dout(new_Jinkela_wire_3472)
    );

    bfr new_Jinkela_buffer_2482 (
        .din(new_Jinkela_wire_3495),
        .dout(new_Jinkela_wire_3496)
    );

    bfr new_Jinkela_buffer_2463 (
        .din(new_Jinkela_wire_3472),
        .dout(new_Jinkela_wire_3473)
    );

    spl2 new_Jinkela_splitter_362 (
        .a(_0170_),
        .b(new_Jinkela_wire_3667),
        .c(new_Jinkela_wire_3668)
    );

    bfr new_Jinkela_buffer_2464 (
        .din(new_Jinkela_wire_3473),
        .dout(new_Jinkela_wire_3474)
    );

    bfr new_Jinkela_buffer_2483 (
        .din(new_Jinkela_wire_3496),
        .dout(new_Jinkela_wire_3497)
    );

    bfr new_Jinkela_buffer_2465 (
        .din(new_Jinkela_wire_3474),
        .dout(new_Jinkela_wire_3475)
    );

    bfr new_Jinkela_buffer_2540 (
        .din(new_Jinkela_wire_3559),
        .dout(new_Jinkela_wire_3560)
    );

    bfr new_Jinkela_buffer_2466 (
        .din(new_Jinkela_wire_3475),
        .dout(new_Jinkela_wire_3476)
    );

    bfr new_Jinkela_buffer_2484 (
        .din(new_Jinkela_wire_3497),
        .dout(new_Jinkela_wire_3498)
    );

    bfr new_Jinkela_buffer_2467 (
        .din(new_Jinkela_wire_3476),
        .dout(new_Jinkela_wire_3477)
    );

    bfr new_Jinkela_buffer_2641 (
        .din(_0453_),
        .dout(new_Jinkela_wire_3669)
    );

    bfr new_Jinkela_buffer_2468 (
        .din(new_Jinkela_wire_3477),
        .dout(new_Jinkela_wire_3478)
    );

    bfr new_Jinkela_buffer_2485 (
        .din(new_Jinkela_wire_3498),
        .dout(new_Jinkela_wire_3499)
    );

    bfr new_Jinkela_buffer_2469 (
        .din(new_Jinkela_wire_3478),
        .dout(new_Jinkela_wire_3479)
    );

    bfr new_Jinkela_buffer_2541 (
        .din(new_Jinkela_wire_3560),
        .dout(new_Jinkela_wire_3561)
    );

    bfr new_Jinkela_buffer_2470 (
        .din(new_Jinkela_wire_3479),
        .dout(new_Jinkela_wire_3480)
    );

    bfr new_Jinkela_buffer_2486 (
        .din(new_Jinkela_wire_3499),
        .dout(new_Jinkela_wire_3500)
    );

    spl2 new_Jinkela_splitter_354 (
        .a(new_Jinkela_wire_3480),
        .b(new_Jinkela_wire_3481),
        .c(new_Jinkela_wire_3482)
    );

    bfr new_Jinkela_buffer_2487 (
        .din(new_Jinkela_wire_3500),
        .dout(new_Jinkela_wire_3501)
    );

    spl2 new_Jinkela_splitter_364 (
        .a(_1328_),
        .b(new_Jinkela_wire_3701),
        .c(new_Jinkela_wire_3702)
    );

    bfr new_Jinkela_buffer_2537 (
        .din(_1560_),
        .dout(new_Jinkela_wire_3557)
    );

    and_bb _2455_ (
        .a(new_Jinkela_wire_13204),
        .b(new_Jinkela_wire_11039),
        .c(_1494_)
    );

    or_bb _2456_ (
        .a(new_Jinkela_wire_14695),
        .b(new_Jinkela_wire_17979),
        .c(_1495_)
    );

    or_bb _2457_ (
        .a(new_Jinkela_wire_7318),
        .b(new_Jinkela_wire_15687),
        .c(_1496_)
    );

    or_ii _2458_ (
        .a(new_Jinkela_wire_7319),
        .b(new_Jinkela_wire_15688),
        .c(_1497_)
    );

    or_ii _2459_ (
        .a(new_Jinkela_wire_14662),
        .b(new_Jinkela_wire_11228),
        .c(_1498_)
    );

    and_ii _2460_ (
        .a(new_Jinkela_wire_3888),
        .b(new_Jinkela_wire_18732),
        .c(_1499_)
    );

    and_bb _2461_ (
        .a(new_Jinkela_wire_3889),
        .b(new_Jinkela_wire_18733),
        .c(_1500_)
    );

    or_bb _2462_ (
        .a(new_Jinkela_wire_6518),
        .b(new_Jinkela_wire_6363),
        .c(_1501_)
    );

    or_bb _2463_ (
        .a(new_Jinkela_wire_17063),
        .b(new_Jinkela_wire_20386),
        .c(_1503_)
    );

    or_ii _2464_ (
        .a(new_Jinkela_wire_17064),
        .b(new_Jinkela_wire_20387),
        .c(_1504_)
    );

    or_ii _2465_ (
        .a(new_Jinkela_wire_20321),
        .b(new_Jinkela_wire_13990),
        .c(_1505_)
    );

    and_ii _2466_ (
        .a(new_Jinkela_wire_21195),
        .b(new_Jinkela_wire_15023),
        .c(_1506_)
    );

    and_bb _2467_ (
        .a(new_Jinkela_wire_21196),
        .b(new_Jinkela_wire_15024),
        .c(_1507_)
    );

    or_bb _2468_ (
        .a(new_Jinkela_wire_3814),
        .b(new_Jinkela_wire_6735),
        .c(_1508_)
    );

    or_bb _2469_ (
        .a(new_Jinkela_wire_4664),
        .b(new_Jinkela_wire_13387),
        .c(_1509_)
    );

    or_ii _2470_ (
        .a(new_Jinkela_wire_4665),
        .b(new_Jinkela_wire_13388),
        .c(_1510_)
    );

    or_ii _2471_ (
        .a(new_Jinkela_wire_1258),
        .b(new_Jinkela_wire_1577),
        .c(_1511_)
    );

    and_ii _2472_ (
        .a(new_Jinkela_wire_6768),
        .b(new_Jinkela_wire_9906),
        .c(_1512_)
    );

    and_bb _2473_ (
        .a(new_Jinkela_wire_6769),
        .b(new_Jinkela_wire_9907),
        .c(_1514_)
    );

    or_bb _2474_ (
        .a(new_Jinkela_wire_19079),
        .b(new_Jinkela_wire_13214),
        .c(_1515_)
    );

    or_bb _2475_ (
        .a(new_Jinkela_wire_10257),
        .b(new_Jinkela_wire_5727),
        .c(_1516_)
    );

    or_ii _2476_ (
        .a(new_Jinkela_wire_10258),
        .b(new_Jinkela_wire_5728),
        .c(_1517_)
    );

    or_ii _2477_ (
        .a(new_Jinkela_wire_18688),
        .b(new_Jinkela_wire_4074),
        .c(_1518_)
    );

    and_ii _2478_ (
        .a(new_Jinkela_wire_5733),
        .b(new_Jinkela_wire_2310),
        .c(_1519_)
    );

    and_bb _2479_ (
        .a(new_Jinkela_wire_5734),
        .b(new_Jinkela_wire_2311),
        .c(_1520_)
    );

    or_bb _2480_ (
        .a(new_Jinkela_wire_7504),
        .b(new_Jinkela_wire_19296),
        .c(_1521_)
    );

    or_bb _2481_ (
        .a(new_Jinkela_wire_15775),
        .b(new_Jinkela_wire_1777),
        .c(_1522_)
    );

    or_ii _2482_ (
        .a(new_Jinkela_wire_15776),
        .b(new_Jinkela_wire_1778),
        .c(_1523_)
    );

    or_ii _2483_ (
        .a(new_Jinkela_wire_20359),
        .b(new_Jinkela_wire_16999),
        .c(_1525_)
    );

    and_ii _2484_ (
        .a(new_Jinkela_wire_5687),
        .b(new_Jinkela_wire_5798),
        .c(_1526_)
    );

    and_bb _2485_ (
        .a(new_Jinkela_wire_5688),
        .b(new_Jinkela_wire_5799),
        .c(_1527_)
    );

    or_bb _2486_ (
        .a(new_Jinkela_wire_19734),
        .b(new_Jinkela_wire_9521),
        .c(_1528_)
    );

    or_bb _2487_ (
        .a(new_Jinkela_wire_19544),
        .b(new_Jinkela_wire_13055),
        .c(_1529_)
    );

    or_ii _2488_ (
        .a(new_Jinkela_wire_19545),
        .b(new_Jinkela_wire_13056),
        .c(_1530_)
    );

    or_ii _2489_ (
        .a(new_Jinkela_wire_720),
        .b(new_Jinkela_wire_8867),
        .c(_1531_)
    );

    and_ii _2490_ (
        .a(new_Jinkela_wire_1281),
        .b(new_Jinkela_wire_8274),
        .c(_1532_)
    );

    and_bb _2491_ (
        .a(new_Jinkela_wire_1282),
        .b(new_Jinkela_wire_8275),
        .c(_1533_)
    );

    or_bb _2492_ (
        .a(new_Jinkela_wire_2422),
        .b(new_Jinkela_wire_4688),
        .c(_1534_)
    );

    or_bb _2493_ (
        .a(new_Jinkela_wire_18969),
        .b(new_Jinkela_wire_4901),
        .c(_1536_)
    );

    or_ii _2494_ (
        .a(new_Jinkela_wire_18970),
        .b(new_Jinkela_wire_4902),
        .c(_1537_)
    );

    or_ii _2495_ (
        .a(new_Jinkela_wire_8963),
        .b(new_Jinkela_wire_13685),
        .c(_1538_)
    );

    and_ii _2496_ (
        .a(new_Jinkela_wire_13199),
        .b(new_Jinkela_wire_12903),
        .c(_1539_)
    );

    spl2 new_Jinkela_splitter_1121 (
        .a(_0027_),
        .b(new_Jinkela_wire_15672),
        .c(new_Jinkela_wire_15673)
    );

    bfr new_Jinkela_buffer_12825 (
        .din(new_Jinkela_wire_15346),
        .dout(new_Jinkela_wire_15347)
    );

    bfr new_Jinkela_buffer_12976 (
        .din(new_Jinkela_wire_15499),
        .dout(new_Jinkela_wire_15500)
    );

    bfr new_Jinkela_buffer_12935 (
        .din(new_Jinkela_wire_15456),
        .dout(new_Jinkela_wire_15457)
    );

    bfr new_Jinkela_buffer_12826 (
        .din(new_Jinkela_wire_15347),
        .dout(new_Jinkela_wire_15348)
    );

    bfr new_Jinkela_buffer_12827 (
        .din(new_Jinkela_wire_15348),
        .dout(new_Jinkela_wire_15349)
    );

    bfr new_Jinkela_buffer_12936 (
        .din(new_Jinkela_wire_15457),
        .dout(new_Jinkela_wire_15458)
    );

    bfr new_Jinkela_buffer_12828 (
        .din(new_Jinkela_wire_15349),
        .dout(new_Jinkela_wire_15350)
    );

    bfr new_Jinkela_buffer_13009 (
        .din(new_Jinkela_wire_15538),
        .dout(new_Jinkela_wire_15539)
    );

    bfr new_Jinkela_buffer_12829 (
        .din(new_Jinkela_wire_15350),
        .dout(new_Jinkela_wire_15351)
    );

    bfr new_Jinkela_buffer_12977 (
        .din(new_Jinkela_wire_15500),
        .dout(new_Jinkela_wire_15501)
    );

    bfr new_Jinkela_buffer_12937 (
        .din(new_Jinkela_wire_15458),
        .dout(new_Jinkela_wire_15459)
    );

    bfr new_Jinkela_buffer_12830 (
        .din(new_Jinkela_wire_15351),
        .dout(new_Jinkela_wire_15352)
    );

    bfr new_Jinkela_buffer_12831 (
        .din(new_Jinkela_wire_15352),
        .dout(new_Jinkela_wire_15353)
    );

    bfr new_Jinkela_buffer_12938 (
        .din(new_Jinkela_wire_15459),
        .dout(new_Jinkela_wire_15460)
    );

    bfr new_Jinkela_buffer_12832 (
        .din(new_Jinkela_wire_15353),
        .dout(new_Jinkela_wire_15354)
    );

    bfr new_Jinkela_buffer_13027 (
        .din(new_Jinkela_wire_15560),
        .dout(new_Jinkela_wire_15561)
    );

    bfr new_Jinkela_buffer_12833 (
        .din(new_Jinkela_wire_15354),
        .dout(new_Jinkela_wire_15355)
    );

    bfr new_Jinkela_buffer_12978 (
        .din(new_Jinkela_wire_15501),
        .dout(new_Jinkela_wire_15502)
    );

    bfr new_Jinkela_buffer_12939 (
        .din(new_Jinkela_wire_15460),
        .dout(new_Jinkela_wire_15461)
    );

    bfr new_Jinkela_buffer_12834 (
        .din(new_Jinkela_wire_15355),
        .dout(new_Jinkela_wire_15356)
    );

    bfr new_Jinkela_buffer_12835 (
        .din(new_Jinkela_wire_15356),
        .dout(new_Jinkela_wire_15357)
    );

    bfr new_Jinkela_buffer_12940 (
        .din(new_Jinkela_wire_15461),
        .dout(new_Jinkela_wire_15462)
    );

    bfr new_Jinkela_buffer_12836 (
        .din(new_Jinkela_wire_15357),
        .dout(new_Jinkela_wire_15358)
    );

    bfr new_Jinkela_buffer_13010 (
        .din(new_Jinkela_wire_15539),
        .dout(new_Jinkela_wire_15540)
    );

    bfr new_Jinkela_buffer_12837 (
        .din(new_Jinkela_wire_15358),
        .dout(new_Jinkela_wire_15359)
    );

    bfr new_Jinkela_buffer_12979 (
        .din(new_Jinkela_wire_15502),
        .dout(new_Jinkela_wire_15503)
    );

    bfr new_Jinkela_buffer_12941 (
        .din(new_Jinkela_wire_15462),
        .dout(new_Jinkela_wire_15463)
    );

    bfr new_Jinkela_buffer_12838 (
        .din(new_Jinkela_wire_15359),
        .dout(new_Jinkela_wire_15360)
    );

    bfr new_Jinkela_buffer_12839 (
        .din(new_Jinkela_wire_15360),
        .dout(new_Jinkela_wire_15361)
    );

    bfr new_Jinkela_buffer_12942 (
        .din(new_Jinkela_wire_15463),
        .dout(new_Jinkela_wire_15464)
    );

    bfr new_Jinkela_buffer_12840 (
        .din(new_Jinkela_wire_15361),
        .dout(new_Jinkela_wire_15362)
    );

    bfr new_Jinkela_buffer_12841 (
        .din(new_Jinkela_wire_15362),
        .dout(new_Jinkela_wire_15363)
    );

    bfr new_Jinkela_buffer_12980 (
        .din(new_Jinkela_wire_15503),
        .dout(new_Jinkela_wire_15504)
    );

    bfr new_Jinkela_buffer_12943 (
        .din(new_Jinkela_wire_15464),
        .dout(new_Jinkela_wire_15465)
    );

    bfr new_Jinkela_buffer_12842 (
        .din(new_Jinkela_wire_15363),
        .dout(new_Jinkela_wire_15364)
    );

    bfr new_Jinkela_buffer_12843 (
        .din(new_Jinkela_wire_15364),
        .dout(new_Jinkela_wire_15365)
    );

    bfr new_Jinkela_buffer_13127 (
        .din(_0922_),
        .dout(new_Jinkela_wire_15671)
    );

    bfr new_Jinkela_buffer_12944 (
        .din(new_Jinkela_wire_15465),
        .dout(new_Jinkela_wire_15466)
    );

    bfr new_Jinkela_buffer_12844 (
        .din(new_Jinkela_wire_15365),
        .dout(new_Jinkela_wire_15366)
    );

    bfr new_Jinkela_buffer_13011 (
        .din(new_Jinkela_wire_15540),
        .dout(new_Jinkela_wire_15541)
    );

    bfr new_Jinkela_buffer_12845 (
        .din(new_Jinkela_wire_15366),
        .dout(new_Jinkela_wire_15367)
    );

    bfr new_Jinkela_buffer_12981 (
        .din(new_Jinkela_wire_15504),
        .dout(new_Jinkela_wire_15505)
    );

    bfr new_Jinkela_buffer_2542 (
        .din(new_Jinkela_wire_3561),
        .dout(new_Jinkela_wire_3562)
    );

    bfr new_Jinkela_buffer_9395 (
        .din(new_Jinkela_wire_11470),
        .dout(new_Jinkela_wire_11471)
    );

    bfr new_Jinkela_buffer_16285 (
        .din(new_Jinkela_wire_19447),
        .dout(new_Jinkela_wire_19448)
    );

    bfr new_Jinkela_buffer_2488 (
        .din(new_Jinkela_wire_3501),
        .dout(new_Jinkela_wire_3502)
    );

    spl2 new_Jinkela_splitter_898 (
        .a(_1629_),
        .b(new_Jinkela_wire_11724),
        .c(new_Jinkela_wire_11725)
    );

    bfr new_Jinkela_buffer_16332 (
        .din(new_Jinkela_wire_19498),
        .dout(new_Jinkela_wire_19499)
    );

    bfr new_Jinkela_buffer_2642 (
        .din(new_Jinkela_wire_3669),
        .dout(new_Jinkela_wire_3670)
    );

    bfr new_Jinkela_buffer_9396 (
        .din(new_Jinkela_wire_11471),
        .dout(new_Jinkela_wire_11472)
    );

    bfr new_Jinkela_buffer_16286 (
        .din(new_Jinkela_wire_19448),
        .dout(new_Jinkela_wire_19449)
    );

    bfr new_Jinkela_buffer_2489 (
        .din(new_Jinkela_wire_3502),
        .dout(new_Jinkela_wire_3503)
    );

    bfr new_Jinkela_buffer_9451 (
        .din(new_Jinkela_wire_11538),
        .dout(new_Jinkela_wire_11539)
    );

    spl2 new_Jinkela_splitter_1444 (
        .a(_0811_),
        .b(new_Jinkela_wire_19732),
        .c(new_Jinkela_wire_19733)
    );

    bfr new_Jinkela_buffer_2543 (
        .din(new_Jinkela_wire_3562),
        .dout(new_Jinkela_wire_3563)
    );

    bfr new_Jinkela_buffer_9397 (
        .din(new_Jinkela_wire_11472),
        .dout(new_Jinkela_wire_11473)
    );

    bfr new_Jinkela_buffer_16287 (
        .din(new_Jinkela_wire_19449),
        .dout(new_Jinkela_wire_19450)
    );

    bfr new_Jinkela_buffer_2490 (
        .din(new_Jinkela_wire_3503),
        .dout(new_Jinkela_wire_3504)
    );

    bfr new_Jinkela_buffer_9454 (
        .din(new_Jinkela_wire_11541),
        .dout(new_Jinkela_wire_11542)
    );

    bfr new_Jinkela_buffer_16333 (
        .din(new_Jinkela_wire_19499),
        .dout(new_Jinkela_wire_19500)
    );

    bfr new_Jinkela_buffer_9398 (
        .din(new_Jinkela_wire_11473),
        .dout(new_Jinkela_wire_11474)
    );

    bfr new_Jinkela_buffer_16288 (
        .din(new_Jinkela_wire_19450),
        .dout(new_Jinkela_wire_19451)
    );

    bfr new_Jinkela_buffer_2491 (
        .din(new_Jinkela_wire_3504),
        .dout(new_Jinkela_wire_3505)
    );

    bfr new_Jinkela_buffer_16541 (
        .din(_1527_),
        .dout(new_Jinkela_wire_19734)
    );

    bfr new_Jinkela_buffer_9524 (
        .din(_0988_),
        .dout(new_Jinkela_wire_11618)
    );

    bfr new_Jinkela_buffer_16384 (
        .din(new_Jinkela_wire_19572),
        .dout(new_Jinkela_wire_19573)
    );

    bfr new_Jinkela_buffer_2544 (
        .din(new_Jinkela_wire_3563),
        .dout(new_Jinkela_wire_3564)
    );

    bfr new_Jinkela_buffer_9399 (
        .din(new_Jinkela_wire_11474),
        .dout(new_Jinkela_wire_11475)
    );

    bfr new_Jinkela_buffer_16289 (
        .din(new_Jinkela_wire_19451),
        .dout(new_Jinkela_wire_19452)
    );

    bfr new_Jinkela_buffer_2492 (
        .din(new_Jinkela_wire_3505),
        .dout(new_Jinkela_wire_3506)
    );

    bfr new_Jinkela_buffer_9455 (
        .din(new_Jinkela_wire_11542),
        .dout(new_Jinkela_wire_11543)
    );

    bfr new_Jinkela_buffer_16334 (
        .din(new_Jinkela_wire_19500),
        .dout(new_Jinkela_wire_19501)
    );

    bfr new_Jinkela_buffer_2643 (
        .din(new_Jinkela_wire_3670),
        .dout(new_Jinkela_wire_3671)
    );

    bfr new_Jinkela_buffer_9400 (
        .din(new_Jinkela_wire_11475),
        .dout(new_Jinkela_wire_11476)
    );

    bfr new_Jinkela_buffer_16290 (
        .din(new_Jinkela_wire_19452),
        .dout(new_Jinkela_wire_19453)
    );

    bfr new_Jinkela_buffer_2493 (
        .din(new_Jinkela_wire_3506),
        .dout(new_Jinkela_wire_3507)
    );

    spl2 new_Jinkela_splitter_897 (
        .a(_0702_),
        .b(new_Jinkela_wire_11722),
        .c(new_Jinkela_wire_11723)
    );

    spl2 new_Jinkela_splitter_1446 (
        .a(_0598_),
        .b(new_Jinkela_wire_19737),
        .c(new_Jinkela_wire_19738)
    );

    bfr new_Jinkela_buffer_2545 (
        .din(new_Jinkela_wire_3564),
        .dout(new_Jinkela_wire_3565)
    );

    bfr new_Jinkela_buffer_9401 (
        .din(new_Jinkela_wire_11476),
        .dout(new_Jinkela_wire_11477)
    );

    bfr new_Jinkela_buffer_16291 (
        .din(new_Jinkela_wire_19453),
        .dout(new_Jinkela_wire_19454)
    );

    bfr new_Jinkela_buffer_2494 (
        .din(new_Jinkela_wire_3507),
        .dout(new_Jinkela_wire_3508)
    );

    bfr new_Jinkela_buffer_9456 (
        .din(new_Jinkela_wire_11543),
        .dout(new_Jinkela_wire_11544)
    );

    bfr new_Jinkela_buffer_16335 (
        .din(new_Jinkela_wire_19501),
        .dout(new_Jinkela_wire_19502)
    );

    bfr new_Jinkela_buffer_9402 (
        .din(new_Jinkela_wire_11477),
        .dout(new_Jinkela_wire_11478)
    );

    bfr new_Jinkela_buffer_16292 (
        .din(new_Jinkela_wire_19454),
        .dout(new_Jinkela_wire_19455)
    );

    spl2 new_Jinkela_splitter_366 (
        .a(_0362_),
        .b(new_Jinkela_wire_3709),
        .c(new_Jinkela_wire_3710)
    );

    bfr new_Jinkela_buffer_2495 (
        .din(new_Jinkela_wire_3508),
        .dout(new_Jinkela_wire_3509)
    );

    bfr new_Jinkela_buffer_9525 (
        .din(new_Jinkela_wire_11618),
        .dout(new_Jinkela_wire_11619)
    );

    bfr new_Jinkela_buffer_16497 (
        .din(new_Jinkela_wire_19687),
        .dout(new_Jinkela_wire_19688)
    );

    bfr new_Jinkela_buffer_16385 (
        .din(new_Jinkela_wire_19573),
        .dout(new_Jinkela_wire_19574)
    );

    bfr new_Jinkela_buffer_2546 (
        .din(new_Jinkela_wire_3565),
        .dout(new_Jinkela_wire_3566)
    );

    bfr new_Jinkela_buffer_9403 (
        .din(new_Jinkela_wire_11478),
        .dout(new_Jinkela_wire_11479)
    );

    bfr new_Jinkela_buffer_16293 (
        .din(new_Jinkela_wire_19455),
        .dout(new_Jinkela_wire_19456)
    );

    bfr new_Jinkela_buffer_2496 (
        .din(new_Jinkela_wire_3509),
        .dout(new_Jinkela_wire_3510)
    );

    bfr new_Jinkela_buffer_9457 (
        .din(new_Jinkela_wire_11544),
        .dout(new_Jinkela_wire_11545)
    );

    bfr new_Jinkela_buffer_16336 (
        .din(new_Jinkela_wire_19502),
        .dout(new_Jinkela_wire_19503)
    );

    bfr new_Jinkela_buffer_2644 (
        .din(new_Jinkela_wire_3671),
        .dout(new_Jinkela_wire_3672)
    );

    bfr new_Jinkela_buffer_9404 (
        .din(new_Jinkela_wire_11479),
        .dout(new_Jinkela_wire_11480)
    );

    bfr new_Jinkela_buffer_16294 (
        .din(new_Jinkela_wire_19456),
        .dout(new_Jinkela_wire_19457)
    );

    bfr new_Jinkela_buffer_2497 (
        .din(new_Jinkela_wire_3510),
        .dout(new_Jinkela_wire_3511)
    );

    bfr new_Jinkela_buffer_2547 (
        .din(new_Jinkela_wire_3566),
        .dout(new_Jinkela_wire_3567)
    );

    bfr new_Jinkela_buffer_9405 (
        .din(new_Jinkela_wire_11480),
        .dout(new_Jinkela_wire_11481)
    );

    bfr new_Jinkela_buffer_16295 (
        .din(new_Jinkela_wire_19457),
        .dout(new_Jinkela_wire_19458)
    );

    bfr new_Jinkela_buffer_2498 (
        .din(new_Jinkela_wire_3511),
        .dout(new_Jinkela_wire_3512)
    );

    bfr new_Jinkela_buffer_9458 (
        .din(new_Jinkela_wire_11545),
        .dout(new_Jinkela_wire_11546)
    );

    bfr new_Jinkela_buffer_16337 (
        .din(new_Jinkela_wire_19503),
        .dout(new_Jinkela_wire_19504)
    );

    bfr new_Jinkela_buffer_2671 (
        .din(new_Jinkela_wire_3704),
        .dout(new_Jinkela_wire_3705)
    );

    bfr new_Jinkela_buffer_9406 (
        .din(new_Jinkela_wire_11481),
        .dout(new_Jinkela_wire_11482)
    );

    bfr new_Jinkela_buffer_16296 (
        .din(new_Jinkela_wire_19458),
        .dout(new_Jinkela_wire_19459)
    );

    spl2 new_Jinkela_splitter_367 (
        .a(_0921_),
        .b(new_Jinkela_wire_3711),
        .c(new_Jinkela_wire_3712)
    );

    bfr new_Jinkela_buffer_2499 (
        .din(new_Jinkela_wire_3512),
        .dout(new_Jinkela_wire_3513)
    );

    bfr new_Jinkela_buffer_9526 (
        .din(new_Jinkela_wire_11619),
        .dout(new_Jinkela_wire_11620)
    );

    bfr new_Jinkela_buffer_16386 (
        .din(new_Jinkela_wire_19574),
        .dout(new_Jinkela_wire_19575)
    );

    bfr new_Jinkela_buffer_2548 (
        .din(new_Jinkela_wire_3567),
        .dout(new_Jinkela_wire_3568)
    );

    bfr new_Jinkela_buffer_9407 (
        .din(new_Jinkela_wire_11482),
        .dout(new_Jinkela_wire_11483)
    );

    bfr new_Jinkela_buffer_16297 (
        .din(new_Jinkela_wire_19459),
        .dout(new_Jinkela_wire_19460)
    );

    bfr new_Jinkela_buffer_2500 (
        .din(new_Jinkela_wire_3513),
        .dout(new_Jinkela_wire_3514)
    );

    bfr new_Jinkela_buffer_9459 (
        .din(new_Jinkela_wire_11546),
        .dout(new_Jinkela_wire_11547)
    );

    bfr new_Jinkela_buffer_16338 (
        .din(new_Jinkela_wire_19504),
        .dout(new_Jinkela_wire_19505)
    );

    bfr new_Jinkela_buffer_2645 (
        .din(new_Jinkela_wire_3672),
        .dout(new_Jinkela_wire_3673)
    );

    bfr new_Jinkela_buffer_9408 (
        .din(new_Jinkela_wire_11483),
        .dout(new_Jinkela_wire_11484)
    );

    bfr new_Jinkela_buffer_16298 (
        .din(new_Jinkela_wire_19460),
        .dout(new_Jinkela_wire_19461)
    );

    bfr new_Jinkela_buffer_2501 (
        .din(new_Jinkela_wire_3514),
        .dout(new_Jinkela_wire_3515)
    );

    bfr new_Jinkela_buffer_9626 (
        .din(_1403_),
        .dout(new_Jinkela_wire_11726)
    );

    bfr new_Jinkela_buffer_2549 (
        .din(new_Jinkela_wire_3568),
        .dout(new_Jinkela_wire_3569)
    );

    bfr new_Jinkela_buffer_9409 (
        .din(new_Jinkela_wire_11484),
        .dout(new_Jinkela_wire_11485)
    );

    bfr new_Jinkela_buffer_16299 (
        .din(new_Jinkela_wire_19461),
        .dout(new_Jinkela_wire_19462)
    );

    bfr new_Jinkela_buffer_2502 (
        .din(new_Jinkela_wire_3515),
        .dout(new_Jinkela_wire_3516)
    );

    bfr new_Jinkela_buffer_9460 (
        .din(new_Jinkela_wire_11547),
        .dout(new_Jinkela_wire_11548)
    );

    bfr new_Jinkela_buffer_16339 (
        .din(new_Jinkela_wire_19505),
        .dout(new_Jinkela_wire_19506)
    );

    spl2 new_Jinkela_splitter_368 (
        .a(_1568_),
        .b(new_Jinkela_wire_3713),
        .c(new_Jinkela_wire_3714)
    );

    bfr new_Jinkela_buffer_9410 (
        .din(new_Jinkela_wire_11485),
        .dout(new_Jinkela_wire_11486)
    );

    bfr new_Jinkela_buffer_16300 (
        .din(new_Jinkela_wire_19462),
        .dout(new_Jinkela_wire_19463)
    );

    bfr new_Jinkela_buffer_2503 (
        .din(new_Jinkela_wire_3516),
        .dout(new_Jinkela_wire_3517)
    );

    bfr new_Jinkela_buffer_9527 (
        .din(new_Jinkela_wire_11620),
        .dout(new_Jinkela_wire_11621)
    );

    bfr new_Jinkela_buffer_16498 (
        .din(new_Jinkela_wire_19688),
        .dout(new_Jinkela_wire_19689)
    );

    bfr new_Jinkela_buffer_16387 (
        .din(new_Jinkela_wire_19575),
        .dout(new_Jinkela_wire_19576)
    );

    bfr new_Jinkela_buffer_2550 (
        .din(new_Jinkela_wire_3569),
        .dout(new_Jinkela_wire_3570)
    );

    bfr new_Jinkela_buffer_9411 (
        .din(new_Jinkela_wire_11486),
        .dout(new_Jinkela_wire_11487)
    );

    bfr new_Jinkela_buffer_16301 (
        .din(new_Jinkela_wire_19463),
        .dout(new_Jinkela_wire_19464)
    );

    bfr new_Jinkela_buffer_2504 (
        .din(new_Jinkela_wire_3517),
        .dout(new_Jinkela_wire_3518)
    );

    bfr new_Jinkela_buffer_9461 (
        .din(new_Jinkela_wire_11548),
        .dout(new_Jinkela_wire_11549)
    );

    bfr new_Jinkela_buffer_16340 (
        .din(new_Jinkela_wire_19506),
        .dout(new_Jinkela_wire_19507)
    );

    bfr new_Jinkela_buffer_2646 (
        .din(new_Jinkela_wire_3673),
        .dout(new_Jinkela_wire_3674)
    );

    bfr new_Jinkela_buffer_9412 (
        .din(new_Jinkela_wire_11487),
        .dout(new_Jinkela_wire_11488)
    );

    bfr new_Jinkela_buffer_16302 (
        .din(new_Jinkela_wire_19464),
        .dout(new_Jinkela_wire_19465)
    );

    bfr new_Jinkela_buffer_2505 (
        .din(new_Jinkela_wire_3518),
        .dout(new_Jinkela_wire_3519)
    );

    spl2 new_Jinkela_splitter_900 (
        .a(_0144_),
        .b(new_Jinkela_wire_11825),
        .c(new_Jinkela_wire_11826)
    );

    bfr new_Jinkela_buffer_9627 (
        .din(_0436_),
        .dout(new_Jinkela_wire_11727)
    );

    bfr new_Jinkela_buffer_2551 (
        .din(new_Jinkela_wire_3570),
        .dout(new_Jinkela_wire_3571)
    );

    bfr new_Jinkela_buffer_9413 (
        .din(new_Jinkela_wire_11488),
        .dout(new_Jinkela_wire_11489)
    );

    spl2 new_Jinkela_splitter_1430 (
        .a(new_Jinkela_wire_19465),
        .b(new_Jinkela_wire_19466),
        .c(new_Jinkela_wire_19467)
    );

    bfr new_Jinkela_buffer_2506 (
        .din(new_Jinkela_wire_3519),
        .dout(new_Jinkela_wire_3520)
    );

    bfr new_Jinkela_buffer_9462 (
        .din(new_Jinkela_wire_11549),
        .dout(new_Jinkela_wire_11550)
    );

    bfr new_Jinkela_buffer_16388 (
        .din(new_Jinkela_wire_19576),
        .dout(new_Jinkela_wire_19577)
    );

    bfr new_Jinkela_buffer_2672 (
        .din(new_Jinkela_wire_3705),
        .dout(new_Jinkela_wire_3706)
    );

    bfr new_Jinkela_buffer_9414 (
        .din(new_Jinkela_wire_11489),
        .dout(new_Jinkela_wire_11490)
    );

    bfr new_Jinkela_buffer_16341 (
        .din(new_Jinkela_wire_19507),
        .dout(new_Jinkela_wire_19508)
    );

    bfr new_Jinkela_buffer_2507 (
        .din(new_Jinkela_wire_3520),
        .dout(new_Jinkela_wire_3521)
    );

    bfr new_Jinkela_buffer_9528 (
        .din(new_Jinkela_wire_11621),
        .dout(new_Jinkela_wire_11622)
    );

    bfr new_Jinkela_buffer_16342 (
        .din(new_Jinkela_wire_19508),
        .dout(new_Jinkela_wire_19509)
    );

    bfr new_Jinkela_buffer_2552 (
        .din(new_Jinkela_wire_3571),
        .dout(new_Jinkela_wire_3572)
    );

    bfr new_Jinkela_buffer_9415 (
        .din(new_Jinkela_wire_11490),
        .dout(new_Jinkela_wire_11491)
    );

    spl2 new_Jinkela_splitter_365 (
        .a(_1148_),
        .b(new_Jinkela_wire_3703),
        .c(new_Jinkela_wire_3704)
    );

    spl2 new_Jinkela_splitter_1445 (
        .a(_0684_),
        .b(new_Jinkela_wire_19735),
        .c(new_Jinkela_wire_19736)
    );

    bfr new_Jinkela_buffer_2508 (
        .din(new_Jinkela_wire_3521),
        .dout(new_Jinkela_wire_3522)
    );

    bfr new_Jinkela_buffer_9463 (
        .din(new_Jinkela_wire_11550),
        .dout(new_Jinkela_wire_11551)
    );

    bfr new_Jinkela_buffer_16343 (
        .din(new_Jinkela_wire_19509),
        .dout(new_Jinkela_wire_19510)
    );

    bfr new_Jinkela_buffer_9416 (
        .din(new_Jinkela_wire_11491),
        .dout(new_Jinkela_wire_11492)
    );

    spl2 new_Jinkela_splitter_901 (
        .a(_0393_),
        .b(new_Jinkela_wire_11827),
        .c(new_Jinkela_wire_11828)
    );

    bfr new_Jinkela_buffer_9417 (
        .din(new_Jinkela_wire_11492),
        .dout(new_Jinkela_wire_11493)
    );

    bfr new_Jinkela_buffer_9464 (
        .din(new_Jinkela_wire_11551),
        .dout(new_Jinkela_wire_11552)
    );

    bfr new_Jinkela_buffer_9418 (
        .din(new_Jinkela_wire_11493),
        .dout(new_Jinkela_wire_11494)
    );

    bfr new_Jinkela_buffer_9529 (
        .din(new_Jinkela_wire_11622),
        .dout(new_Jinkela_wire_11623)
    );

    bfr new_Jinkela_buffer_9419 (
        .din(new_Jinkela_wire_11494),
        .dout(new_Jinkela_wire_11495)
    );

    bfr new_Jinkela_buffer_9465 (
        .din(new_Jinkela_wire_11552),
        .dout(new_Jinkela_wire_11553)
    );

    bfr new_Jinkela_buffer_9420 (
        .din(new_Jinkela_wire_11495),
        .dout(new_Jinkela_wire_11496)
    );

    bfr new_Jinkela_buffer_9628 (
        .din(new_Jinkela_wire_11727),
        .dout(new_Jinkela_wire_11728)
    );

    bfr new_Jinkela_buffer_9421 (
        .din(new_Jinkela_wire_11496),
        .dout(new_Jinkela_wire_11497)
    );

    bfr new_Jinkela_buffer_9466 (
        .din(new_Jinkela_wire_11553),
        .dout(new_Jinkela_wire_11554)
    );

    bfr new_Jinkela_buffer_9422 (
        .din(new_Jinkela_wire_11497),
        .dout(new_Jinkela_wire_11498)
    );

    bfr new_Jinkela_buffer_9530 (
        .din(new_Jinkela_wire_11623),
        .dout(new_Jinkela_wire_11624)
    );

    bfr new_Jinkela_buffer_9423 (
        .din(new_Jinkela_wire_11498),
        .dout(new_Jinkela_wire_11499)
    );

    bfr new_Jinkela_buffer_9467 (
        .din(new_Jinkela_wire_11554),
        .dout(new_Jinkela_wire_11555)
    );

    bfr new_Jinkela_buffer_9424 (
        .din(new_Jinkela_wire_11499),
        .dout(new_Jinkela_wire_11500)
    );

    bfr new_Jinkela_buffer_9425 (
        .din(new_Jinkela_wire_11500),
        .dout(new_Jinkela_wire_11501)
    );

    bfr new_Jinkela_buffer_9468 (
        .din(new_Jinkela_wire_11555),
        .dout(new_Jinkela_wire_11556)
    );

    bfr new_Jinkela_buffer_9426 (
        .din(new_Jinkela_wire_11501),
        .dout(new_Jinkela_wire_11502)
    );

    bfr new_Jinkela_buffer_9531 (
        .din(new_Jinkela_wire_11624),
        .dout(new_Jinkela_wire_11625)
    );

    bfr new_Jinkela_buffer_9427 (
        .din(new_Jinkela_wire_11502),
        .dout(new_Jinkela_wire_11503)
    );

    bfr new_Jinkela_buffer_9469 (
        .din(new_Jinkela_wire_11556),
        .dout(new_Jinkela_wire_11557)
    );

    bfr new_Jinkela_buffer_9428 (
        .din(new_Jinkela_wire_11503),
        .dout(new_Jinkela_wire_11504)
    );

    bfr new_Jinkela_buffer_9629 (
        .din(new_Jinkela_wire_11728),
        .dout(new_Jinkela_wire_11729)
    );

    bfr new_Jinkela_buffer_9429 (
        .din(new_Jinkela_wire_11504),
        .dout(new_Jinkela_wire_11505)
    );

    bfr new_Jinkela_buffer_9470 (
        .din(new_Jinkela_wire_11557),
        .dout(new_Jinkela_wire_11558)
    );

    bfr new_Jinkela_buffer_9430 (
        .din(new_Jinkela_wire_11505),
        .dout(new_Jinkela_wire_11506)
    );

    bfr new_Jinkela_buffer_9532 (
        .din(new_Jinkela_wire_11625),
        .dout(new_Jinkela_wire_11626)
    );

    bfr new_Jinkela_buffer_9431 (
        .din(new_Jinkela_wire_11506),
        .dout(new_Jinkela_wire_11507)
    );

    bfr new_Jinkela_buffer_9471 (
        .din(new_Jinkela_wire_11558),
        .dout(new_Jinkela_wire_11559)
    );

    bfr new_Jinkela_buffer_9432 (
        .din(new_Jinkela_wire_11507),
        .dout(new_Jinkela_wire_11508)
    );

    spl2 new_Jinkela_splitter_902 (
        .a(_1751_),
        .b(new_Jinkela_wire_11830),
        .c(new_Jinkela_wire_11831)
    );

    bfr new_Jinkela_buffer_9723 (
        .din(_1312_),
        .dout(new_Jinkela_wire_11829)
    );

    bfr new_Jinkela_buffer_9433 (
        .din(new_Jinkela_wire_11508),
        .dout(new_Jinkela_wire_11509)
    );

    bfr new_Jinkela_buffer_9472 (
        .din(new_Jinkela_wire_11559),
        .dout(new_Jinkela_wire_11560)
    );

    bfr new_Jinkela_buffer_9434 (
        .din(new_Jinkela_wire_11509),
        .dout(new_Jinkela_wire_11510)
    );

    bfr new_Jinkela_buffer_9533 (
        .din(new_Jinkela_wire_11626),
        .dout(new_Jinkela_wire_11627)
    );

    bfr new_Jinkela_buffer_9435 (
        .din(new_Jinkela_wire_11510),
        .dout(new_Jinkela_wire_11511)
    );

    bfr new_Jinkela_buffer_9473 (
        .din(new_Jinkela_wire_11560),
        .dout(new_Jinkela_wire_11561)
    );

    bfr new_Jinkela_buffer_9436 (
        .din(new_Jinkela_wire_11511),
        .dout(new_Jinkela_wire_11512)
    );

    bfr new_Jinkela_buffer_9630 (
        .din(new_Jinkela_wire_11729),
        .dout(new_Jinkela_wire_11730)
    );

    and_ii _3382_ (
        .a(new_Jinkela_wire_12058),
        .b(new_Jinkela_wire_4659),
        .c(_0665_)
    );

    and_bb _3383_ (
        .a(new_Jinkela_wire_12059),
        .b(new_Jinkela_wire_4660),
        .c(_0667_)
    );

    or_bb _3384_ (
        .a(new_Jinkela_wire_2591),
        .b(new_Jinkela_wire_8580),
        .c(_0668_)
    );

    and_ii _3385_ (
        .a(new_Jinkela_wire_21218),
        .b(new_Jinkela_wire_15731),
        .c(_0669_)
    );

    and_bb _3386_ (
        .a(new_Jinkela_wire_21219),
        .b(new_Jinkela_wire_15732),
        .c(_0670_)
    );

    or_bb _3387_ (
        .a(new_Jinkela_wire_4327),
        .b(new_Jinkela_wire_7263),
        .c(_0671_)
    );

    and_ii _3388_ (
        .a(new_Jinkela_wire_2147),
        .b(new_Jinkela_wire_2115),
        .c(_0672_)
    );

    and_bb _3389_ (
        .a(new_Jinkela_wire_2148),
        .b(new_Jinkela_wire_2116),
        .c(_0673_)
    );

    or_bb _3390_ (
        .a(new_Jinkela_wire_21179),
        .b(new_Jinkela_wire_5467),
        .c(_0674_)
    );

    and_ii _3391_ (
        .a(new_Jinkela_wire_15771),
        .b(new_Jinkela_wire_6759),
        .c(_0675_)
    );

    and_bb _3392_ (
        .a(new_Jinkela_wire_15772),
        .b(new_Jinkela_wire_6760),
        .c(_0676_)
    );

    or_bb _3393_ (
        .a(new_Jinkela_wire_14006),
        .b(new_Jinkela_wire_11534),
        .c(_0678_)
    );

    and_ii _3394_ (
        .a(new_Jinkela_wire_5538),
        .b(new_Jinkela_wire_10556),
        .c(_0679_)
    );

    and_bb _3395_ (
        .a(new_Jinkela_wire_5539),
        .b(new_Jinkela_wire_10557),
        .c(_0680_)
    );

    or_bb _3396_ (
        .a(new_Jinkela_wire_5456),
        .b(new_Jinkela_wire_14277),
        .c(_0681_)
    );

    and_ii _3397_ (
        .a(new_Jinkela_wire_14279),
        .b(new_Jinkela_wire_15122),
        .c(_0682_)
    );

    and_bb _3398_ (
        .a(new_Jinkela_wire_14280),
        .b(new_Jinkela_wire_15123),
        .c(_0683_)
    );

    or_bb _3399_ (
        .a(new_Jinkela_wire_12738),
        .b(new_Jinkela_wire_11416),
        .c(_0684_)
    );

    and_ii _3400_ (
        .a(new_Jinkela_wire_19735),
        .b(new_Jinkela_wire_14890),
        .c(_0685_)
    );

    and_bb _3401_ (
        .a(new_Jinkela_wire_19736),
        .b(new_Jinkela_wire_14891),
        .c(_0686_)
    );

    or_bb _3402_ (
        .a(new_Jinkela_wire_15553),
        .b(new_Jinkela_wire_16104),
        .c(_0687_)
    );

    and_ii _3403_ (
        .a(new_Jinkela_wire_3716),
        .b(new_Jinkela_wire_8027),
        .c(_0689_)
    );

    and_bb _3404_ (
        .a(new_Jinkela_wire_3717),
        .b(new_Jinkela_wire_8028),
        .c(_0690_)
    );

    and_ii _3405_ (
        .a(new_Jinkela_wire_13996),
        .b(new_Jinkela_wire_18537),
        .c(_0691_)
    );

    and_bb _3406_ (
        .a(new_Jinkela_wire_18514),
        .b(new_Jinkela_wire_7738),
        .c(_0692_)
    );

    and_ii _3407_ (
        .a(new_Jinkela_wire_18515),
        .b(new_Jinkela_wire_7739),
        .c(_0693_)
    );

    or_bb _3408_ (
        .a(new_Jinkela_wire_5997),
        .b(new_Jinkela_wire_3435),
        .c(new_net_3944)
    );

    or_bb _3409_ (
        .a(new_Jinkela_wire_3436),
        .b(new_Jinkela_wire_18562),
        .c(_0694_)
    );

    and_ii _3410_ (
        .a(new_Jinkela_wire_16105),
        .b(new_Jinkela_wire_11421),
        .c(_0695_)
    );

    and_bb _3411_ (
        .a(new_Jinkela_wire_677),
        .b(new_Jinkela_wire_501),
        .c(_0696_)
    );

    and_ii _3412_ (
        .a(new_Jinkela_wire_14278),
        .b(new_Jinkela_wire_11539),
        .c(_0697_)
    );

    and_bb _3413_ (
        .a(new_Jinkela_wire_28),
        .b(new_Jinkela_wire_522),
        .c(_0699_)
    );

    and_ii _3414_ (
        .a(new_Jinkela_wire_5468),
        .b(new_Jinkela_wire_7268),
        .c(_0700_)
    );

    and_bb _3415_ (
        .a(new_Jinkela_wire_187),
        .b(new_Jinkela_wire_144),
        .c(_0701_)
    );

    and_ii _3416_ (
        .a(new_Jinkela_wire_8581),
        .b(new_Jinkela_wire_6253),
        .c(_0702_)
    );

    and_bb _3417_ (
        .a(new_Jinkela_wire_390),
        .b(new_Jinkela_wire_208),
        .c(_0703_)
    );

    and_ii _3418_ (
        .a(new_Jinkela_wire_12222),
        .b(new_Jinkela_wire_5702),
        .c(_0704_)
    );

    and_bb _3419_ (
        .a(new_Jinkela_wire_412),
        .b(new_Jinkela_wire_592),
        .c(_0705_)
    );

    and_ii _3420_ (
        .a(new_Jinkela_wire_3556),
        .b(new_Jinkela_wire_18960),
        .c(_0706_)
    );

    and_bb _3421_ (
        .a(new_Jinkela_wire_156),
        .b(new_Jinkela_wire_120),
        .c(_0707_)
    );

    and_ii _3422_ (
        .a(new_Jinkela_wire_6683),
        .b(new_Jinkela_wire_20141),
        .c(_0708_)
    );

    and_bb _3423_ (
        .a(new_Jinkela_wire_596),
        .b(new_Jinkela_wire_5),
        .c(_0710_)
    );

    bfr new_Jinkela_buffer_2647 (
        .din(new_Jinkela_wire_3674),
        .dout(new_Jinkela_wire_3675)
    );

    spl2 new_Jinkela_splitter_1110 (
        .a(new_Jinkela_wire_15466),
        .b(new_Jinkela_wire_15467),
        .c(new_Jinkela_wire_15468)
    );

    bfr new_Jinkela_buffer_6081 (
        .din(_0919_),
        .dout(new_Jinkela_wire_7719)
    );

    bfr new_Jinkela_buffer_12846 (
        .din(new_Jinkela_wire_15367),
        .dout(new_Jinkela_wire_15368)
    );

    bfr new_Jinkela_buffer_2509 (
        .din(new_Jinkela_wire_3522),
        .dout(new_Jinkela_wire_3523)
    );

    bfr new_Jinkela_buffer_5948 (
        .din(new_Jinkela_wire_7555),
        .dout(new_Jinkela_wire_7556)
    );

    bfr new_Jinkela_buffer_2553 (
        .din(new_Jinkela_wire_3572),
        .dout(new_Jinkela_wire_3573)
    );

    bfr new_Jinkela_buffer_5992 (
        .din(new_Jinkela_wire_7607),
        .dout(new_Jinkela_wire_7608)
    );

    bfr new_Jinkela_buffer_13028 (
        .din(new_Jinkela_wire_15561),
        .dout(new_Jinkela_wire_15562)
    );

    bfr new_Jinkela_buffer_12847 (
        .din(new_Jinkela_wire_15368),
        .dout(new_Jinkela_wire_15369)
    );

    bfr new_Jinkela_buffer_2510 (
        .din(new_Jinkela_wire_3523),
        .dout(new_Jinkela_wire_3524)
    );

    bfr new_Jinkela_buffer_5949 (
        .din(new_Jinkela_wire_7556),
        .dout(new_Jinkela_wire_7557)
    );

    bfr new_Jinkela_buffer_12982 (
        .din(new_Jinkela_wire_15505),
        .dout(new_Jinkela_wire_15506)
    );

    bfr new_Jinkela_buffer_6080 (
        .din(_0597_),
        .dout(new_Jinkela_wire_7718)
    );

    bfr new_Jinkela_buffer_12848 (
        .din(new_Jinkela_wire_15369),
        .dout(new_Jinkela_wire_15370)
    );

    bfr new_Jinkela_buffer_2511 (
        .din(new_Jinkela_wire_3524),
        .dout(new_Jinkela_wire_3525)
    );

    bfr new_Jinkela_buffer_5950 (
        .din(new_Jinkela_wire_7557),
        .dout(new_Jinkela_wire_7558)
    );

    bfr new_Jinkela_buffer_2554 (
        .din(new_Jinkela_wire_3573),
        .dout(new_Jinkela_wire_3574)
    );

    bfr new_Jinkela_buffer_5993 (
        .din(new_Jinkela_wire_7608),
        .dout(new_Jinkela_wire_7609)
    );

    bfr new_Jinkela_buffer_12849 (
        .din(new_Jinkela_wire_15370),
        .dout(new_Jinkela_wire_15371)
    );

    bfr new_Jinkela_buffer_2512 (
        .din(new_Jinkela_wire_3525),
        .dout(new_Jinkela_wire_3526)
    );

    bfr new_Jinkela_buffer_5951 (
        .din(new_Jinkela_wire_7558),
        .dout(new_Jinkela_wire_7559)
    );

    bfr new_Jinkela_buffer_2648 (
        .din(new_Jinkela_wire_3675),
        .dout(new_Jinkela_wire_3676)
    );

    bfr new_Jinkela_buffer_13012 (
        .din(new_Jinkela_wire_15541),
        .dout(new_Jinkela_wire_15542)
    );

    spl2 new_Jinkela_splitter_668 (
        .a(_0134_),
        .b(new_Jinkela_wire_7720),
        .c(new_Jinkela_wire_7721)
    );

    bfr new_Jinkela_buffer_12850 (
        .din(new_Jinkela_wire_15371),
        .dout(new_Jinkela_wire_15372)
    );

    bfr new_Jinkela_buffer_2513 (
        .din(new_Jinkela_wire_3526),
        .dout(new_Jinkela_wire_3527)
    );

    bfr new_Jinkela_buffer_5952 (
        .din(new_Jinkela_wire_7559),
        .dout(new_Jinkela_wire_7560)
    );

    bfr new_Jinkela_buffer_12983 (
        .din(new_Jinkela_wire_15506),
        .dout(new_Jinkela_wire_15507)
    );

    bfr new_Jinkela_buffer_2555 (
        .din(new_Jinkela_wire_3574),
        .dout(new_Jinkela_wire_3575)
    );

    bfr new_Jinkela_buffer_5994 (
        .din(new_Jinkela_wire_7609),
        .dout(new_Jinkela_wire_7610)
    );

    bfr new_Jinkela_buffer_12851 (
        .din(new_Jinkela_wire_15372),
        .dout(new_Jinkela_wire_15373)
    );

    bfr new_Jinkela_buffer_2514 (
        .din(new_Jinkela_wire_3527),
        .dout(new_Jinkela_wire_3528)
    );

    bfr new_Jinkela_buffer_5953 (
        .din(new_Jinkela_wire_7560),
        .dout(new_Jinkela_wire_7561)
    );

    bfr new_Jinkela_buffer_2673 (
        .din(new_Jinkela_wire_3706),
        .dout(new_Jinkela_wire_3707)
    );

    spl2 new_Jinkela_splitter_669 (
        .a(_0764_),
        .b(new_Jinkela_wire_7726),
        .c(new_Jinkela_wire_7727)
    );

    spl2 new_Jinkela_splitter_1122 (
        .a(_0910_),
        .b(new_Jinkela_wire_15674),
        .c(new_Jinkela_wire_15675)
    );

    bfr new_Jinkela_buffer_6082 (
        .din(new_Jinkela_wire_7721),
        .dout(new_Jinkela_wire_7722)
    );

    bfr new_Jinkela_buffer_12852 (
        .din(new_Jinkela_wire_15373),
        .dout(new_Jinkela_wire_15374)
    );

    bfr new_Jinkela_buffer_2515 (
        .din(new_Jinkela_wire_3528),
        .dout(new_Jinkela_wire_3529)
    );

    bfr new_Jinkela_buffer_5954 (
        .din(new_Jinkela_wire_7561),
        .dout(new_Jinkela_wire_7562)
    );

    bfr new_Jinkela_buffer_12984 (
        .din(new_Jinkela_wire_15507),
        .dout(new_Jinkela_wire_15508)
    );

    bfr new_Jinkela_buffer_2556 (
        .din(new_Jinkela_wire_3575),
        .dout(new_Jinkela_wire_3576)
    );

    bfr new_Jinkela_buffer_5995 (
        .din(new_Jinkela_wire_7610),
        .dout(new_Jinkela_wire_7611)
    );

    bfr new_Jinkela_buffer_12853 (
        .din(new_Jinkela_wire_15374),
        .dout(new_Jinkela_wire_15375)
    );

    bfr new_Jinkela_buffer_2516 (
        .din(new_Jinkela_wire_3529),
        .dout(new_Jinkela_wire_3530)
    );

    bfr new_Jinkela_buffer_5955 (
        .din(new_Jinkela_wire_7562),
        .dout(new_Jinkela_wire_7563)
    );

    bfr new_Jinkela_buffer_13128 (
        .din(new_Jinkela_wire_15677),
        .dout(new_Jinkela_wire_15678)
    );

    bfr new_Jinkela_buffer_2649 (
        .din(new_Jinkela_wire_3676),
        .dout(new_Jinkela_wire_3677)
    );

    bfr new_Jinkela_buffer_13013 (
        .din(new_Jinkela_wire_15542),
        .dout(new_Jinkela_wire_15543)
    );

    bfr new_Jinkela_buffer_12854 (
        .din(new_Jinkela_wire_15375),
        .dout(new_Jinkela_wire_15376)
    );

    bfr new_Jinkela_buffer_2517 (
        .din(new_Jinkela_wire_3530),
        .dout(new_Jinkela_wire_3531)
    );

    bfr new_Jinkela_buffer_5956 (
        .din(new_Jinkela_wire_7563),
        .dout(new_Jinkela_wire_7564)
    );

    bfr new_Jinkela_buffer_12985 (
        .din(new_Jinkela_wire_15508),
        .dout(new_Jinkela_wire_15509)
    );

    bfr new_Jinkela_buffer_2557 (
        .din(new_Jinkela_wire_3576),
        .dout(new_Jinkela_wire_3577)
    );

    bfr new_Jinkela_buffer_5996 (
        .din(new_Jinkela_wire_7611),
        .dout(new_Jinkela_wire_7612)
    );

    bfr new_Jinkela_buffer_12855 (
        .din(new_Jinkela_wire_15376),
        .dout(new_Jinkela_wire_15377)
    );

    bfr new_Jinkela_buffer_2518 (
        .din(new_Jinkela_wire_3531),
        .dout(new_Jinkela_wire_3532)
    );

    bfr new_Jinkela_buffer_5957 (
        .din(new_Jinkela_wire_7564),
        .dout(new_Jinkela_wire_7565)
    );

    bfr new_Jinkela_buffer_13029 (
        .din(new_Jinkela_wire_15562),
        .dout(new_Jinkela_wire_15563)
    );

    bfr new_Jinkela_buffer_2675 (
        .din(_0115_),
        .dout(new_Jinkela_wire_3715)
    );

    bfr new_Jinkela_buffer_6086 (
        .din(_1555_),
        .dout(new_Jinkela_wire_7728)
    );

    bfr new_Jinkela_buffer_12856 (
        .din(new_Jinkela_wire_15377),
        .dout(new_Jinkela_wire_15378)
    );

    bfr new_Jinkela_buffer_2519 (
        .din(new_Jinkela_wire_3532),
        .dout(new_Jinkela_wire_3533)
    );

    bfr new_Jinkela_buffer_5958 (
        .din(new_Jinkela_wire_7565),
        .dout(new_Jinkela_wire_7566)
    );

    bfr new_Jinkela_buffer_12986 (
        .din(new_Jinkela_wire_15509),
        .dout(new_Jinkela_wire_15510)
    );

    bfr new_Jinkela_buffer_2558 (
        .din(new_Jinkela_wire_3577),
        .dout(new_Jinkela_wire_3578)
    );

    bfr new_Jinkela_buffer_5997 (
        .din(new_Jinkela_wire_7612),
        .dout(new_Jinkela_wire_7613)
    );

    bfr new_Jinkela_buffer_2520 (
        .din(new_Jinkela_wire_3533),
        .dout(new_Jinkela_wire_3534)
    );

    bfr new_Jinkela_buffer_5959 (
        .din(new_Jinkela_wire_7566),
        .dout(new_Jinkela_wire_7567)
    );

    bfr new_Jinkela_buffer_13014 (
        .din(new_Jinkela_wire_15543),
        .dout(new_Jinkela_wire_15544)
    );

    bfr new_Jinkela_buffer_12987 (
        .din(new_Jinkela_wire_15510),
        .dout(new_Jinkela_wire_15511)
    );

    bfr new_Jinkela_buffer_2650 (
        .din(new_Jinkela_wire_3677),
        .dout(new_Jinkela_wire_3678)
    );

    bfr new_Jinkela_buffer_2521 (
        .din(new_Jinkela_wire_3534),
        .dout(new_Jinkela_wire_3535)
    );

    bfr new_Jinkela_buffer_5960 (
        .din(new_Jinkela_wire_7567),
        .dout(new_Jinkela_wire_7568)
    );

    bfr new_Jinkela_buffer_12988 (
        .din(new_Jinkela_wire_15511),
        .dout(new_Jinkela_wire_15512)
    );

    bfr new_Jinkela_buffer_2559 (
        .din(new_Jinkela_wire_3578),
        .dout(new_Jinkela_wire_3579)
    );

    bfr new_Jinkela_buffer_5998 (
        .din(new_Jinkela_wire_7613),
        .dout(new_Jinkela_wire_7614)
    );

    bfr new_Jinkela_buffer_2522 (
        .din(new_Jinkela_wire_3535),
        .dout(new_Jinkela_wire_3536)
    );

    bfr new_Jinkela_buffer_5961 (
        .din(new_Jinkela_wire_7568),
        .dout(new_Jinkela_wire_7569)
    );

    bfr new_Jinkela_buffer_13015 (
        .din(new_Jinkela_wire_15544),
        .dout(new_Jinkela_wire_15545)
    );

    bfr new_Jinkela_buffer_12989 (
        .din(new_Jinkela_wire_15512),
        .dout(new_Jinkela_wire_15513)
    );

    bfr new_Jinkela_buffer_2674 (
        .din(new_Jinkela_wire_3707),
        .dout(new_Jinkela_wire_3708)
    );

    bfr new_Jinkela_buffer_6083 (
        .din(new_Jinkela_wire_7722),
        .dout(new_Jinkela_wire_7723)
    );

    bfr new_Jinkela_buffer_2523 (
        .din(new_Jinkela_wire_3536),
        .dout(new_Jinkela_wire_3537)
    );

    bfr new_Jinkela_buffer_5962 (
        .din(new_Jinkela_wire_7569),
        .dout(new_Jinkela_wire_7570)
    );

    bfr new_Jinkela_buffer_13030 (
        .din(new_Jinkela_wire_15563),
        .dout(new_Jinkela_wire_15564)
    );

    bfr new_Jinkela_buffer_12990 (
        .din(new_Jinkela_wire_15513),
        .dout(new_Jinkela_wire_15514)
    );

    bfr new_Jinkela_buffer_2560 (
        .din(new_Jinkela_wire_3579),
        .dout(new_Jinkela_wire_3580)
    );

    bfr new_Jinkela_buffer_5999 (
        .din(new_Jinkela_wire_7614),
        .dout(new_Jinkela_wire_7615)
    );

    bfr new_Jinkela_buffer_2524 (
        .din(new_Jinkela_wire_3537),
        .dout(new_Jinkela_wire_3538)
    );

    bfr new_Jinkela_buffer_5963 (
        .din(new_Jinkela_wire_7570),
        .dout(new_Jinkela_wire_7571)
    );

    bfr new_Jinkela_buffer_13016 (
        .din(new_Jinkela_wire_15545),
        .dout(new_Jinkela_wire_15546)
    );

    bfr new_Jinkela_buffer_12991 (
        .din(new_Jinkela_wire_15514),
        .dout(new_Jinkela_wire_15515)
    );

    bfr new_Jinkela_buffer_2651 (
        .din(new_Jinkela_wire_3678),
        .dout(new_Jinkela_wire_3679)
    );

    spl2 new_Jinkela_splitter_672 (
        .a(_1794_),
        .b(new_Jinkela_wire_7734),
        .c(new_Jinkela_wire_7735)
    );

    spl2 new_Jinkela_splitter_670 (
        .a(_1491_),
        .b(new_Jinkela_wire_7729),
        .c(new_Jinkela_wire_7730)
    );

    bfr new_Jinkela_buffer_2525 (
        .din(new_Jinkela_wire_3538),
        .dout(new_Jinkela_wire_3539)
    );

    bfr new_Jinkela_buffer_5964 (
        .din(new_Jinkela_wire_7571),
        .dout(new_Jinkela_wire_7572)
    );

    bfr new_Jinkela_buffer_12992 (
        .din(new_Jinkela_wire_15515),
        .dout(new_Jinkela_wire_15516)
    );

    bfr new_Jinkela_buffer_2561 (
        .din(new_Jinkela_wire_3580),
        .dout(new_Jinkela_wire_3581)
    );

    bfr new_Jinkela_buffer_6000 (
        .din(new_Jinkela_wire_7615),
        .dout(new_Jinkela_wire_7616)
    );

    spl2 new_Jinkela_splitter_1123 (
        .a(_0991_),
        .b(new_Jinkela_wire_15676),
        .c(new_Jinkela_wire_15677)
    );

    bfr new_Jinkela_buffer_2526 (
        .din(new_Jinkela_wire_3539),
        .dout(new_Jinkela_wire_3540)
    );

    bfr new_Jinkela_buffer_5965 (
        .din(new_Jinkela_wire_7572),
        .dout(new_Jinkela_wire_7573)
    );

    bfr new_Jinkela_buffer_13017 (
        .din(new_Jinkela_wire_15546),
        .dout(new_Jinkela_wire_15547)
    );

    spl2 new_Jinkela_splitter_370 (
        .a(_0942_),
        .b(new_Jinkela_wire_3718),
        .c(new_Jinkela_wire_3719)
    );

    bfr new_Jinkela_buffer_6084 (
        .din(new_Jinkela_wire_7723),
        .dout(new_Jinkela_wire_7724)
    );

    bfr new_Jinkela_buffer_13031 (
        .din(new_Jinkela_wire_15564),
        .dout(new_Jinkela_wire_15565)
    );

    spl2 new_Jinkela_splitter_369 (
        .a(_0687_),
        .b(new_Jinkela_wire_3716),
        .c(new_Jinkela_wire_3717)
    );

    bfr new_Jinkela_buffer_2527 (
        .din(new_Jinkela_wire_3540),
        .dout(new_Jinkela_wire_3541)
    );

    bfr new_Jinkela_buffer_5966 (
        .din(new_Jinkela_wire_7573),
        .dout(new_Jinkela_wire_7574)
    );

    bfr new_Jinkela_buffer_13018 (
        .din(new_Jinkela_wire_15547),
        .dout(new_Jinkela_wire_15548)
    );

    bfr new_Jinkela_buffer_2562 (
        .din(new_Jinkela_wire_3581),
        .dout(new_Jinkela_wire_3582)
    );

    bfr new_Jinkela_buffer_6001 (
        .din(new_Jinkela_wire_7616),
        .dout(new_Jinkela_wire_7617)
    );

    bfr new_Jinkela_buffer_13132 (
        .din(_0892_),
        .dout(new_Jinkela_wire_15682)
    );

    bfr new_Jinkela_buffer_2528 (
        .din(new_Jinkela_wire_3541),
        .dout(new_Jinkela_wire_3542)
    );

    bfr new_Jinkela_buffer_5967 (
        .din(new_Jinkela_wire_7574),
        .dout(new_Jinkela_wire_7575)
    );

    bfr new_Jinkela_buffer_13019 (
        .din(new_Jinkela_wire_15548),
        .dout(new_Jinkela_wire_15549)
    );

    bfr new_Jinkela_buffer_2652 (
        .din(new_Jinkela_wire_3679),
        .dout(new_Jinkela_wire_3680)
    );

    bfr new_Jinkela_buffer_6087 (
        .din(new_Jinkela_wire_7730),
        .dout(new_Jinkela_wire_7731)
    );

    bfr new_Jinkela_buffer_13032 (
        .din(new_Jinkela_wire_15565),
        .dout(new_Jinkela_wire_15566)
    );

    bfr new_Jinkela_buffer_2529 (
        .din(new_Jinkela_wire_3542),
        .dout(new_Jinkela_wire_3543)
    );

    bfr new_Jinkela_buffer_5968 (
        .din(new_Jinkela_wire_7575),
        .dout(new_Jinkela_wire_7576)
    );

    bfr new_Jinkela_buffer_13020 (
        .din(new_Jinkela_wire_15549),
        .dout(new_Jinkela_wire_15550)
    );

    bfr new_Jinkela_buffer_9437 (
        .din(new_Jinkela_wire_11512),
        .dout(new_Jinkela_wire_11513)
    );

    bfr new_Jinkela_buffer_9474 (
        .din(new_Jinkela_wire_11561),
        .dout(new_Jinkela_wire_11562)
    );

    bfr new_Jinkela_buffer_9438 (
        .din(new_Jinkela_wire_11513),
        .dout(new_Jinkela_wire_11514)
    );

    bfr new_Jinkela_buffer_9534 (
        .din(new_Jinkela_wire_11627),
        .dout(new_Jinkela_wire_11628)
    );

    bfr new_Jinkela_buffer_9439 (
        .din(new_Jinkela_wire_11514),
        .dout(new_Jinkela_wire_11515)
    );

    bfr new_Jinkela_buffer_9475 (
        .din(new_Jinkela_wire_11562),
        .dout(new_Jinkela_wire_11563)
    );

    bfr new_Jinkela_buffer_9440 (
        .din(new_Jinkela_wire_11515),
        .dout(new_Jinkela_wire_11516)
    );

    spl2 new_Jinkela_splitter_903 (
        .a(_1216_),
        .b(new_Jinkela_wire_11836),
        .c(new_Jinkela_wire_11837)
    );

    bfr new_Jinkela_buffer_9724 (
        .din(new_Jinkela_wire_11831),
        .dout(new_Jinkela_wire_11832)
    );

    bfr new_Jinkela_buffer_9441 (
        .din(new_Jinkela_wire_11516),
        .dout(new_Jinkela_wire_11517)
    );

    bfr new_Jinkela_buffer_9476 (
        .din(new_Jinkela_wire_11563),
        .dout(new_Jinkela_wire_11564)
    );

    bfr new_Jinkela_buffer_9442 (
        .din(new_Jinkela_wire_11517),
        .dout(new_Jinkela_wire_11518)
    );

    bfr new_Jinkela_buffer_9535 (
        .din(new_Jinkela_wire_11628),
        .dout(new_Jinkela_wire_11629)
    );

    bfr new_Jinkela_buffer_9443 (
        .din(new_Jinkela_wire_11518),
        .dout(new_Jinkela_wire_11519)
    );

    bfr new_Jinkela_buffer_9477 (
        .din(new_Jinkela_wire_11564),
        .dout(new_Jinkela_wire_11565)
    );

    bfr new_Jinkela_buffer_9444 (
        .din(new_Jinkela_wire_11519),
        .dout(new_Jinkela_wire_11520)
    );

    bfr new_Jinkela_buffer_9631 (
        .din(new_Jinkela_wire_11730),
        .dout(new_Jinkela_wire_11731)
    );

    bfr new_Jinkela_buffer_9445 (
        .din(new_Jinkela_wire_11520),
        .dout(new_Jinkela_wire_11521)
    );

    bfr new_Jinkela_buffer_9478 (
        .din(new_Jinkela_wire_11565),
        .dout(new_Jinkela_wire_11566)
    );

    bfr new_Jinkela_buffer_9446 (
        .din(new_Jinkela_wire_11521),
        .dout(new_Jinkela_wire_11522)
    );

    bfr new_Jinkela_buffer_9536 (
        .din(new_Jinkela_wire_11629),
        .dout(new_Jinkela_wire_11630)
    );

    spl2 new_Jinkela_splitter_887 (
        .a(new_Jinkela_wire_11522),
        .b(new_Jinkela_wire_11523),
        .c(new_Jinkela_wire_11524)
    );

    bfr new_Jinkela_buffer_9479 (
        .din(new_Jinkela_wire_11566),
        .dout(new_Jinkela_wire_11567)
    );

    bfr new_Jinkela_buffer_9480 (
        .din(new_Jinkela_wire_11567),
        .dout(new_Jinkela_wire_11568)
    );

    bfr new_Jinkela_buffer_9537 (
        .din(new_Jinkela_wire_11630),
        .dout(new_Jinkela_wire_11631)
    );

    bfr new_Jinkela_buffer_9481 (
        .din(new_Jinkela_wire_11568),
        .dout(new_Jinkela_wire_11569)
    );

    bfr new_Jinkela_buffer_9632 (
        .din(new_Jinkela_wire_11731),
        .dout(new_Jinkela_wire_11732)
    );

    bfr new_Jinkela_buffer_9482 (
        .din(new_Jinkela_wire_11569),
        .dout(new_Jinkela_wire_11570)
    );

    bfr new_Jinkela_buffer_9538 (
        .din(new_Jinkela_wire_11631),
        .dout(new_Jinkela_wire_11632)
    );

    bfr new_Jinkela_buffer_9483 (
        .din(new_Jinkela_wire_11570),
        .dout(new_Jinkela_wire_11571)
    );

    bfr new_Jinkela_buffer_9728 (
        .din(_1789_),
        .dout(new_Jinkela_wire_11838)
    );

    bfr new_Jinkela_buffer_9484 (
        .din(new_Jinkela_wire_11571),
        .dout(new_Jinkela_wire_11572)
    );

    bfr new_Jinkela_buffer_9539 (
        .din(new_Jinkela_wire_11632),
        .dout(new_Jinkela_wire_11633)
    );

    bfr new_Jinkela_buffer_9485 (
        .din(new_Jinkela_wire_11572),
        .dout(new_Jinkela_wire_11573)
    );

    bfr new_Jinkela_buffer_9633 (
        .din(new_Jinkela_wire_11732),
        .dout(new_Jinkela_wire_11733)
    );

    bfr new_Jinkela_buffer_9486 (
        .din(new_Jinkela_wire_11573),
        .dout(new_Jinkela_wire_11574)
    );

    bfr new_Jinkela_buffer_9540 (
        .din(new_Jinkela_wire_11633),
        .dout(new_Jinkela_wire_11634)
    );

    bfr new_Jinkela_buffer_9487 (
        .din(new_Jinkela_wire_11574),
        .dout(new_Jinkela_wire_11575)
    );

    bfr new_Jinkela_buffer_9729 (
        .din(_0509_),
        .dout(new_Jinkela_wire_11839)
    );

    bfr new_Jinkela_buffer_9488 (
        .din(new_Jinkela_wire_11575),
        .dout(new_Jinkela_wire_11576)
    );

    bfr new_Jinkela_buffer_9541 (
        .din(new_Jinkela_wire_11634),
        .dout(new_Jinkela_wire_11635)
    );

    bfr new_Jinkela_buffer_9489 (
        .din(new_Jinkela_wire_11576),
        .dout(new_Jinkela_wire_11577)
    );

    bfr new_Jinkela_buffer_6002 (
        .din(new_Jinkela_wire_7617),
        .dout(new_Jinkela_wire_7618)
    );

    bfr new_Jinkela_buffer_16499 (
        .din(new_Jinkela_wire_19689),
        .dout(new_Jinkela_wire_19690)
    );

    bfr new_Jinkela_buffer_16389 (
        .din(new_Jinkela_wire_19577),
        .dout(new_Jinkela_wire_19578)
    );

    bfr new_Jinkela_buffer_5969 (
        .din(new_Jinkela_wire_7576),
        .dout(new_Jinkela_wire_7577)
    );

    bfr new_Jinkela_buffer_16344 (
        .din(new_Jinkela_wire_19510),
        .dout(new_Jinkela_wire_19511)
    );

    bfr new_Jinkela_buffer_6085 (
        .din(new_Jinkela_wire_7724),
        .dout(new_Jinkela_wire_7725)
    );

    bfr new_Jinkela_buffer_5970 (
        .din(new_Jinkela_wire_7577),
        .dout(new_Jinkela_wire_7578)
    );

    bfr new_Jinkela_buffer_16345 (
        .din(new_Jinkela_wire_19511),
        .dout(new_Jinkela_wire_19512)
    );

    bfr new_Jinkela_buffer_6003 (
        .din(new_Jinkela_wire_7618),
        .dout(new_Jinkela_wire_7619)
    );

    bfr new_Jinkela_buffer_16586 (
        .din(new_Jinkela_wire_19794),
        .dout(new_Jinkela_wire_19795)
    );

    bfr new_Jinkela_buffer_16390 (
        .din(new_Jinkela_wire_19578),
        .dout(new_Jinkela_wire_19579)
    );

    bfr new_Jinkela_buffer_5971 (
        .din(new_Jinkela_wire_7578),
        .dout(new_Jinkela_wire_7579)
    );

    bfr new_Jinkela_buffer_16346 (
        .din(new_Jinkela_wire_19512),
        .dout(new_Jinkela_wire_19513)
    );

    spl2 new_Jinkela_splitter_653 (
        .a(new_Jinkela_wire_7579),
        .b(new_Jinkela_wire_7580),
        .c(new_Jinkela_wire_7581)
    );

    bfr new_Jinkela_buffer_16347 (
        .din(new_Jinkela_wire_19513),
        .dout(new_Jinkela_wire_19514)
    );

    bfr new_Jinkela_buffer_6088 (
        .din(_1262_),
        .dout(new_Jinkela_wire_7736)
    );

    bfr new_Jinkela_buffer_16500 (
        .din(new_Jinkela_wire_19690),
        .dout(new_Jinkela_wire_19691)
    );

    bfr new_Jinkela_buffer_16391 (
        .din(new_Jinkela_wire_19579),
        .dout(new_Jinkela_wire_19580)
    );

    bfr new_Jinkela_buffer_6004 (
        .din(new_Jinkela_wire_7619),
        .dout(new_Jinkela_wire_7620)
    );

    bfr new_Jinkela_buffer_16348 (
        .din(new_Jinkela_wire_19514),
        .dout(new_Jinkela_wire_19515)
    );

    bfr new_Jinkela_buffer_6005 (
        .din(new_Jinkela_wire_7620),
        .dout(new_Jinkela_wire_7621)
    );

    bfr new_Jinkela_buffer_6089 (
        .din(_0257_),
        .dout(new_Jinkela_wire_7737)
    );

    bfr new_Jinkela_buffer_16349 (
        .din(new_Jinkela_wire_19515),
        .dout(new_Jinkela_wire_19516)
    );

    spl2 new_Jinkela_splitter_671 (
        .a(new_Jinkela_wire_7731),
        .b(new_Jinkela_wire_7732),
        .c(new_Jinkela_wire_7733)
    );

    bfr new_Jinkela_buffer_6006 (
        .din(new_Jinkela_wire_7621),
        .dout(new_Jinkela_wire_7622)
    );

    bfr new_Jinkela_buffer_16392 (
        .din(new_Jinkela_wire_19580),
        .dout(new_Jinkela_wire_19581)
    );

    bfr new_Jinkela_buffer_16350 (
        .din(new_Jinkela_wire_19516),
        .dout(new_Jinkela_wire_19517)
    );

    bfr new_Jinkela_buffer_6007 (
        .din(new_Jinkela_wire_7622),
        .dout(new_Jinkela_wire_7623)
    );

    spl2 new_Jinkela_splitter_1447 (
        .a(_1135_),
        .b(new_Jinkela_wire_19739),
        .c(new_Jinkela_wire_19740)
    );

    spl2 new_Jinkela_splitter_674 (
        .a(_0124_),
        .b(new_Jinkela_wire_7742),
        .c(new_Jinkela_wire_7743)
    );

    bfr new_Jinkela_buffer_16351 (
        .din(new_Jinkela_wire_19517),
        .dout(new_Jinkela_wire_19518)
    );

    spl2 new_Jinkela_splitter_673 (
        .a(_0615_),
        .b(new_Jinkela_wire_7738),
        .c(new_Jinkela_wire_7739)
    );

    bfr new_Jinkela_buffer_6008 (
        .din(new_Jinkela_wire_7623),
        .dout(new_Jinkela_wire_7624)
    );

    bfr new_Jinkela_buffer_16501 (
        .din(new_Jinkela_wire_19691),
        .dout(new_Jinkela_wire_19692)
    );

    bfr new_Jinkela_buffer_16393 (
        .din(new_Jinkela_wire_19581),
        .dout(new_Jinkela_wire_19582)
    );

    bfr new_Jinkela_buffer_6090 (
        .din(_0872_),
        .dout(new_Jinkela_wire_7740)
    );

    bfr new_Jinkela_buffer_16352 (
        .din(new_Jinkela_wire_19518),
        .dout(new_Jinkela_wire_19519)
    );

    bfr new_Jinkela_buffer_6009 (
        .din(new_Jinkela_wire_7624),
        .dout(new_Jinkela_wire_7625)
    );

    bfr new_Jinkela_buffer_16353 (
        .din(new_Jinkela_wire_19519),
        .dout(new_Jinkela_wire_19520)
    );

    bfr new_Jinkela_buffer_6091 (
        .din(_1630_),
        .dout(new_Jinkela_wire_7741)
    );

    bfr new_Jinkela_buffer_6010 (
        .din(new_Jinkela_wire_7625),
        .dout(new_Jinkela_wire_7626)
    );

    bfr new_Jinkela_buffer_16552 (
        .din(new_Jinkela_wire_19750),
        .dout(new_Jinkela_wire_19751)
    );

    bfr new_Jinkela_buffer_16394 (
        .din(new_Jinkela_wire_19582),
        .dout(new_Jinkela_wire_19583)
    );

    spl2 new_Jinkela_splitter_675 (
        .a(_0824_),
        .b(new_Jinkela_wire_7744),
        .c(new_Jinkela_wire_7745)
    );

    bfr new_Jinkela_buffer_16354 (
        .din(new_Jinkela_wire_19520),
        .dout(new_Jinkela_wire_19521)
    );

    bfr new_Jinkela_buffer_6011 (
        .din(new_Jinkela_wire_7626),
        .dout(new_Jinkela_wire_7627)
    );

    bfr new_Jinkela_buffer_16355 (
        .din(new_Jinkela_wire_19521),
        .dout(new_Jinkela_wire_19522)
    );

    bfr new_Jinkela_buffer_6012 (
        .din(new_Jinkela_wire_7627),
        .dout(new_Jinkela_wire_7628)
    );

    bfr new_Jinkela_buffer_16502 (
        .din(new_Jinkela_wire_19692),
        .dout(new_Jinkela_wire_19693)
    );

    bfr new_Jinkela_buffer_16395 (
        .din(new_Jinkela_wire_19583),
        .dout(new_Jinkela_wire_19584)
    );

    bfr new_Jinkela_buffer_16356 (
        .din(new_Jinkela_wire_19522),
        .dout(new_Jinkela_wire_19523)
    );

    spl2 new_Jinkela_splitter_676 (
        .a(_0423_),
        .b(new_Jinkela_wire_7746),
        .c(new_Jinkela_wire_7747)
    );

    bfr new_Jinkela_buffer_6013 (
        .din(new_Jinkela_wire_7628),
        .dout(new_Jinkela_wire_7629)
    );

    bfr new_Jinkela_buffer_16357 (
        .din(new_Jinkela_wire_19523),
        .dout(new_Jinkela_wire_19524)
    );

    spl2 new_Jinkela_splitter_677 (
        .a(_0844_),
        .b(new_Jinkela_wire_7748),
        .c(new_Jinkela_wire_7749)
    );

    bfr new_Jinkela_buffer_6014 (
        .din(new_Jinkela_wire_7629),
        .dout(new_Jinkela_wire_7630)
    );

    spl2 new_Jinkela_splitter_1454 (
        .a(_1183_),
        .b(new_Jinkela_wire_19908),
        .c(new_Jinkela_wire_19909)
    );

    bfr new_Jinkela_buffer_16396 (
        .din(new_Jinkela_wire_19584),
        .dout(new_Jinkela_wire_19585)
    );

    bfr new_Jinkela_buffer_16358 (
        .din(new_Jinkela_wire_19524),
        .dout(new_Jinkela_wire_19525)
    );

    bfr new_Jinkela_buffer_6092 (
        .din(_0957_),
        .dout(new_Jinkela_wire_7750)
    );

    bfr new_Jinkela_buffer_6015 (
        .din(new_Jinkela_wire_7630),
        .dout(new_Jinkela_wire_7631)
    );

    spl2 new_Jinkela_splitter_679 (
        .a(_0494_),
        .b(new_Jinkela_wire_7833),
        .c(new_Jinkela_wire_7834)
    );

    bfr new_Jinkela_buffer_16359 (
        .din(new_Jinkela_wire_19525),
        .dout(new_Jinkela_wire_19526)
    );

    bfr new_Jinkela_buffer_6093 (
        .din(_0093_),
        .dout(new_Jinkela_wire_7751)
    );

    bfr new_Jinkela_buffer_6016 (
        .din(new_Jinkela_wire_7631),
        .dout(new_Jinkela_wire_7632)
    );

    bfr new_Jinkela_buffer_16503 (
        .din(new_Jinkela_wire_19693),
        .dout(new_Jinkela_wire_19694)
    );

    bfr new_Jinkela_buffer_16397 (
        .din(new_Jinkela_wire_19585),
        .dout(new_Jinkela_wire_19586)
    );

    bfr new_Jinkela_buffer_16360 (
        .din(new_Jinkela_wire_19526),
        .dout(new_Jinkela_wire_19527)
    );

    bfr new_Jinkela_buffer_6173 (
        .din(_1653_),
        .dout(new_Jinkela_wire_7835)
    );

    bfr new_Jinkela_buffer_6017 (
        .din(new_Jinkela_wire_7632),
        .dout(new_Jinkela_wire_7633)
    );

    bfr new_Jinkela_buffer_6094 (
        .din(new_Jinkela_wire_7751),
        .dout(new_Jinkela_wire_7752)
    );

    bfr new_Jinkela_buffer_16361 (
        .din(new_Jinkela_wire_19527),
        .dout(new_Jinkela_wire_19528)
    );

    bfr new_Jinkela_buffer_6018 (
        .din(new_Jinkela_wire_7633),
        .dout(new_Jinkela_wire_7634)
    );

    bfr new_Jinkela_buffer_16398 (
        .din(new_Jinkela_wire_19586),
        .dout(new_Jinkela_wire_19587)
    );

    bfr new_Jinkela_buffer_16362 (
        .din(new_Jinkela_wire_19528),
        .dout(new_Jinkela_wire_19529)
    );

    bfr new_Jinkela_buffer_6019 (
        .din(new_Jinkela_wire_7634),
        .dout(new_Jinkela_wire_7635)
    );

    bfr new_Jinkela_buffer_16697 (
        .din(_1614_),
        .dout(new_Jinkela_wire_19910)
    );

    bfr new_Jinkela_buffer_6095 (
        .din(new_Jinkela_wire_7752),
        .dout(new_Jinkela_wire_7753)
    );

    bfr new_Jinkela_buffer_16363 (
        .din(new_Jinkela_wire_19529),
        .dout(new_Jinkela_wire_19530)
    );

    bfr new_Jinkela_buffer_6020 (
        .din(new_Jinkela_wire_7635),
        .dout(new_Jinkela_wire_7636)
    );

    bfr new_Jinkela_buffer_16504 (
        .din(new_Jinkela_wire_19694),
        .dout(new_Jinkela_wire_19695)
    );

    bfr new_Jinkela_buffer_16399 (
        .din(new_Jinkela_wire_19587),
        .dout(new_Jinkela_wire_19588)
    );

    spl2 new_Jinkela_splitter_681 (
        .a(_0211_),
        .b(new_Jinkela_wire_7842),
        .c(new_Jinkela_wire_7843)
    );

    bfr new_Jinkela_buffer_16364 (
        .din(new_Jinkela_wire_19530),
        .dout(new_Jinkela_wire_19531)
    );

    spl2 new_Jinkela_splitter_680 (
        .a(_1048_),
        .b(new_Jinkela_wire_7836),
        .c(new_Jinkela_wire_7837)
    );

    bfr new_Jinkela_buffer_2564 (
        .din(new_Jinkela_wire_3583),
        .dout(new_Jinkela_wire_3584)
    );

    bfr new_Jinkela_buffer_2530 (
        .din(new_Jinkela_wire_3543),
        .dout(new_Jinkela_wire_3544)
    );

    bfr new_Jinkela_buffer_2653 (
        .din(new_Jinkela_wire_3680),
        .dout(new_Jinkela_wire_3681)
    );

    bfr new_Jinkela_buffer_2531 (
        .din(new_Jinkela_wire_3544),
        .dout(new_Jinkela_wire_3545)
    );

    bfr new_Jinkela_buffer_2565 (
        .din(new_Jinkela_wire_3584),
        .dout(new_Jinkela_wire_3585)
    );

    bfr new_Jinkela_buffer_2532 (
        .din(new_Jinkela_wire_3545),
        .dout(new_Jinkela_wire_3546)
    );

    bfr new_Jinkela_buffer_2678 (
        .din(_0930_),
        .dout(new_Jinkela_wire_3722)
    );

    bfr new_Jinkela_buffer_2533 (
        .din(new_Jinkela_wire_3546),
        .dout(new_Jinkela_wire_3547)
    );

    bfr new_Jinkela_buffer_2566 (
        .din(new_Jinkela_wire_3585),
        .dout(new_Jinkela_wire_3586)
    );

    bfr new_Jinkela_buffer_2534 (
        .din(new_Jinkela_wire_3547),
        .dout(new_Jinkela_wire_3548)
    );

    bfr new_Jinkela_buffer_2654 (
        .din(new_Jinkela_wire_3681),
        .dout(new_Jinkela_wire_3682)
    );

    spl2 new_Jinkela_splitter_356 (
        .a(new_Jinkela_wire_3548),
        .b(new_Jinkela_wire_3549),
        .c(new_Jinkela_wire_3550)
    );

    bfr new_Jinkela_buffer_2677 (
        .din(_0948_),
        .dout(new_Jinkela_wire_3721)
    );

    bfr new_Jinkela_buffer_2567 (
        .din(new_Jinkela_wire_3586),
        .dout(new_Jinkela_wire_3587)
    );

    bfr new_Jinkela_buffer_2568 (
        .din(new_Jinkela_wire_3587),
        .dout(new_Jinkela_wire_3588)
    );

    bfr new_Jinkela_buffer_2655 (
        .din(new_Jinkela_wire_3682),
        .dout(new_Jinkela_wire_3683)
    );

    bfr new_Jinkela_buffer_2569 (
        .din(new_Jinkela_wire_3588),
        .dout(new_Jinkela_wire_3589)
    );

    bfr new_Jinkela_buffer_2768 (
        .din(_1507_),
        .dout(new_Jinkela_wire_3814)
    );

    bfr new_Jinkela_buffer_2570 (
        .din(new_Jinkela_wire_3589),
        .dout(new_Jinkela_wire_3590)
    );

    bfr new_Jinkela_buffer_2656 (
        .din(new_Jinkela_wire_3683),
        .dout(new_Jinkela_wire_3684)
    );

    bfr new_Jinkela_buffer_2571 (
        .din(new_Jinkela_wire_3590),
        .dout(new_Jinkela_wire_3591)
    );

    bfr new_Jinkela_buffer_2769 (
        .din(_1769_),
        .dout(new_Jinkela_wire_3815)
    );

    bfr new_Jinkela_buffer_2572 (
        .din(new_Jinkela_wire_3591),
        .dout(new_Jinkela_wire_3592)
    );

    bfr new_Jinkela_buffer_2657 (
        .din(new_Jinkela_wire_3684),
        .dout(new_Jinkela_wire_3685)
    );

    bfr new_Jinkela_buffer_2573 (
        .din(new_Jinkela_wire_3592),
        .dout(new_Jinkela_wire_3593)
    );

    bfr new_Jinkela_buffer_2679 (
        .din(new_Jinkela_wire_3722),
        .dout(new_Jinkela_wire_3723)
    );

    bfr new_Jinkela_buffer_2574 (
        .din(new_Jinkela_wire_3593),
        .dout(new_Jinkela_wire_3594)
    );

    bfr new_Jinkela_buffer_2658 (
        .din(new_Jinkela_wire_3685),
        .dout(new_Jinkela_wire_3686)
    );

    bfr new_Jinkela_buffer_2575 (
        .din(new_Jinkela_wire_3594),
        .dout(new_Jinkela_wire_3595)
    );

    bfr new_Jinkela_buffer_2770 (
        .din(_0422_),
        .dout(new_Jinkela_wire_3816)
    );

    bfr new_Jinkela_buffer_2576 (
        .din(new_Jinkela_wire_3595),
        .dout(new_Jinkela_wire_3596)
    );

    bfr new_Jinkela_buffer_2659 (
        .din(new_Jinkela_wire_3686),
        .dout(new_Jinkela_wire_3687)
    );

    bfr new_Jinkela_buffer_2577 (
        .din(new_Jinkela_wire_3596),
        .dout(new_Jinkela_wire_3597)
    );

    bfr new_Jinkela_buffer_2680 (
        .din(new_Jinkela_wire_3723),
        .dout(new_Jinkela_wire_3724)
    );

    bfr new_Jinkela_buffer_2578 (
        .din(new_Jinkela_wire_3597),
        .dout(new_Jinkela_wire_3598)
    );

    bfr new_Jinkela_buffer_2660 (
        .din(new_Jinkela_wire_3687),
        .dout(new_Jinkela_wire_3688)
    );

    bfr new_Jinkela_buffer_2579 (
        .din(new_Jinkela_wire_3598),
        .dout(new_Jinkela_wire_3599)
    );

    spl2 new_Jinkela_splitter_372 (
        .a(_0338_),
        .b(new_Jinkela_wire_3817),
        .c(new_Jinkela_wire_3818)
    );

    bfr new_Jinkela_buffer_2580 (
        .din(new_Jinkela_wire_3599),
        .dout(new_Jinkela_wire_3600)
    );

    bfr new_Jinkela_buffer_2661 (
        .din(new_Jinkela_wire_3688),
        .dout(new_Jinkela_wire_3689)
    );

    bfr new_Jinkela_buffer_2581 (
        .din(new_Jinkela_wire_3600),
        .dout(new_Jinkela_wire_3601)
    );

    bfr new_Jinkela_buffer_2681 (
        .din(new_Jinkela_wire_3724),
        .dout(new_Jinkela_wire_3725)
    );

    and_bb _3424_ (
        .a(new_Jinkela_wire_436),
        .b(new_Jinkela_wire_448),
        .c(_0711_)
    );

    and_ii _3425_ (
        .a(new_Jinkela_wire_20363),
        .b(new_Jinkela_wire_14043),
        .c(_0712_)
    );

    and_ii _3426_ (
        .a(new_Jinkela_wire_19318),
        .b(new_Jinkela_wire_6674),
        .c(_0713_)
    );

    and_bb _3427_ (
        .a(new_Jinkela_wire_19319),
        .b(new_Jinkela_wire_6675),
        .c(_0714_)
    );

    or_bb _3428_ (
        .a(new_Jinkela_wire_4291),
        .b(new_Jinkela_wire_14538),
        .c(_0715_)
    );

    and_ii _3429_ (
        .a(new_Jinkela_wire_10083),
        .b(new_Jinkela_wire_18373),
        .c(_0716_)
    );

    and_bb _3430_ (
        .a(new_Jinkela_wire_10084),
        .b(new_Jinkela_wire_18374),
        .c(_0717_)
    );

    or_bb _3431_ (
        .a(new_Jinkela_wire_20901),
        .b(new_Jinkela_wire_10062),
        .c(_0718_)
    );

    and_ii _3432_ (
        .a(new_Jinkela_wire_5708),
        .b(new_Jinkela_wire_2324),
        .c(_0719_)
    );

    and_bb _3433_ (
        .a(new_Jinkela_wire_5709),
        .b(new_Jinkela_wire_2325),
        .c(_0721_)
    );

    or_bb _3434_ (
        .a(new_Jinkela_wire_6617),
        .b(new_Jinkela_wire_18283),
        .c(_0722_)
    );

    and_ii _3435_ (
        .a(new_Jinkela_wire_10692),
        .b(new_Jinkela_wire_4236),
        .c(_0723_)
    );

    and_bb _3436_ (
        .a(new_Jinkela_wire_10693),
        .b(new_Jinkela_wire_4237),
        .c(_0724_)
    );

    or_bb _3437_ (
        .a(new_Jinkela_wire_13678),
        .b(new_Jinkela_wire_3665),
        .c(_0725_)
    );

    and_ii _3438_ (
        .a(new_Jinkela_wire_19059),
        .b(new_Jinkela_wire_16533),
        .c(_0726_)
    );

    and_bb _3439_ (
        .a(new_Jinkela_wire_19060),
        .b(new_Jinkela_wire_16534),
        .c(_0727_)
    );

    or_bb _3440_ (
        .a(new_Jinkela_wire_13064),
        .b(new_Jinkela_wire_20677),
        .c(_0728_)
    );

    and_ii _3441_ (
        .a(new_Jinkela_wire_5721),
        .b(new_Jinkela_wire_12043),
        .c(_0729_)
    );

    and_bb _3442_ (
        .a(new_Jinkela_wire_5722),
        .b(new_Jinkela_wire_12044),
        .c(_0730_)
    );

    or_bb _3443_ (
        .a(new_Jinkela_wire_7291),
        .b(new_Jinkela_wire_10263),
        .c(_0732_)
    );

    and_ii _3444_ (
        .a(new_Jinkela_wire_18291),
        .b(new_Jinkela_wire_5149),
        .c(_0733_)
    );

    and_bb _3445_ (
        .a(new_Jinkela_wire_18292),
        .b(new_Jinkela_wire_5150),
        .c(_0734_)
    );

    or_bb _3446_ (
        .a(new_Jinkela_wire_3446),
        .b(new_Jinkela_wire_16524),
        .c(_0735_)
    );

    and_ii _3447_ (
        .a(new_Jinkela_wire_15994),
        .b(new_Jinkela_wire_12829),
        .c(_0736_)
    );

    and_bb _3448_ (
        .a(new_Jinkela_wire_15995),
        .b(new_Jinkela_wire_12830),
        .c(_0737_)
    );

    or_bb _3449_ (
        .a(new_Jinkela_wire_14309),
        .b(new_Jinkela_wire_1334),
        .c(_0738_)
    );

    and_ii _3450_ (
        .a(new_Jinkela_wire_5430),
        .b(new_Jinkela_wire_11722),
        .c(_0739_)
    );

    and_bb _3451_ (
        .a(new_Jinkela_wire_5431),
        .b(new_Jinkela_wire_11723),
        .c(_0740_)
    );

    or_bb _3452_ (
        .a(new_Jinkela_wire_14273),
        .b(new_Jinkela_wire_19335),
        .c(_0741_)
    );

    and_ii _3453_ (
        .a(new_Jinkela_wire_18223),
        .b(new_Jinkela_wire_18220),
        .c(_0743_)
    );

    and_bb _3454_ (
        .a(new_Jinkela_wire_18224),
        .b(new_Jinkela_wire_18221),
        .c(_0744_)
    );

    or_bb _3455_ (
        .a(new_Jinkela_wire_11021),
        .b(new_Jinkela_wire_16522),
        .c(_0745_)
    );

    and_ii _3456_ (
        .a(new_Jinkela_wire_16941),
        .b(new_Jinkela_wire_843),
        .c(_0746_)
    );

    and_bb _3457_ (
        .a(new_Jinkela_wire_16942),
        .b(new_Jinkela_wire_844),
        .c(_0747_)
    );

    or_bb _3458_ (
        .a(new_Jinkela_wire_15206),
        .b(new_Jinkela_wire_10106),
        .c(_0748_)
    );

    and_ii _3459_ (
        .a(new_Jinkela_wire_2964),
        .b(new_Jinkela_wire_13952),
        .c(_0749_)
    );

    and_bb _3460_ (
        .a(new_Jinkela_wire_2965),
        .b(new_Jinkela_wire_13953),
        .c(_0750_)
    );

    or_bb _3461_ (
        .a(new_Jinkela_wire_9695),
        .b(new_Jinkela_wire_18685),
        .c(_0751_)
    );

    and_ii _3462_ (
        .a(new_Jinkela_wire_3663),
        .b(new_Jinkela_wire_20364),
        .c(_0752_)
    );

    and_bb _3463_ (
        .a(new_Jinkela_wire_3664),
        .b(new_Jinkela_wire_20365),
        .c(_0754_)
    );

    or_bb _3464_ (
        .a(new_Jinkela_wire_19731),
        .b(new_Jinkela_wire_7301),
        .c(_0755_)
    );

    and_ii _3465_ (
        .a(new_Jinkela_wire_13679),
        .b(new_Jinkela_wire_10949),
        .c(_0756_)
    );

    bfr new_Jinkela_buffer_16365 (
        .din(new_Jinkela_wire_19531),
        .dout(new_Jinkela_wire_19532)
    );

    spl2 new_Jinkela_splitter_1449 (
        .a(_1419_),
        .b(new_Jinkela_wire_19783),
        .c(new_Jinkela_wire_19784)
    );

    bfr new_Jinkela_buffer_16400 (
        .din(new_Jinkela_wire_19588),
        .dout(new_Jinkela_wire_19589)
    );

    bfr new_Jinkela_buffer_16366 (
        .din(new_Jinkela_wire_19532),
        .dout(new_Jinkela_wire_19533)
    );

    bfr new_Jinkela_buffer_16367 (
        .din(new_Jinkela_wire_19533),
        .dout(new_Jinkela_wire_19534)
    );

    bfr new_Jinkela_buffer_16505 (
        .din(new_Jinkela_wire_19695),
        .dout(new_Jinkela_wire_19696)
    );

    bfr new_Jinkela_buffer_16401 (
        .din(new_Jinkela_wire_19589),
        .dout(new_Jinkela_wire_19590)
    );

    bfr new_Jinkela_buffer_16368 (
        .din(new_Jinkela_wire_19534),
        .dout(new_Jinkela_wire_19535)
    );

    bfr new_Jinkela_buffer_16369 (
        .din(new_Jinkela_wire_19535),
        .dout(new_Jinkela_wire_19536)
    );

    bfr new_Jinkela_buffer_16402 (
        .din(new_Jinkela_wire_19590),
        .dout(new_Jinkela_wire_19591)
    );

    bfr new_Jinkela_buffer_16370 (
        .din(new_Jinkela_wire_19536),
        .dout(new_Jinkela_wire_19537)
    );

    bfr new_Jinkela_buffer_16582 (
        .din(_0062_),
        .dout(new_Jinkela_wire_19785)
    );

    spl2 new_Jinkela_splitter_1432 (
        .a(new_Jinkela_wire_19537),
        .b(new_Jinkela_wire_19538),
        .c(new_Jinkela_wire_19539)
    );

    bfr new_Jinkela_buffer_16506 (
        .din(new_Jinkela_wire_19696),
        .dout(new_Jinkela_wire_19697)
    );

    bfr new_Jinkela_buffer_16403 (
        .din(new_Jinkela_wire_19591),
        .dout(new_Jinkela_wire_19592)
    );

    bfr new_Jinkela_buffer_16543 (
        .din(new_Jinkela_wire_19741),
        .dout(new_Jinkela_wire_19742)
    );

    bfr new_Jinkela_buffer_16404 (
        .din(new_Jinkela_wire_19592),
        .dout(new_Jinkela_wire_19593)
    );

    bfr new_Jinkela_buffer_16507 (
        .din(new_Jinkela_wire_19697),
        .dout(new_Jinkela_wire_19698)
    );

    bfr new_Jinkela_buffer_16405 (
        .din(new_Jinkela_wire_19593),
        .dout(new_Jinkela_wire_19594)
    );

    bfr new_Jinkela_buffer_16406 (
        .din(new_Jinkela_wire_19594),
        .dout(new_Jinkela_wire_19595)
    );

    bfr new_Jinkela_buffer_16508 (
        .din(new_Jinkela_wire_19698),
        .dout(new_Jinkela_wire_19699)
    );

    bfr new_Jinkela_buffer_16407 (
        .din(new_Jinkela_wire_19595),
        .dout(new_Jinkela_wire_19596)
    );

    bfr new_Jinkela_buffer_16544 (
        .din(new_Jinkela_wire_19742),
        .dout(new_Jinkela_wire_19743)
    );

    bfr new_Jinkela_buffer_16408 (
        .din(new_Jinkela_wire_19596),
        .dout(new_Jinkela_wire_19597)
    );

    bfr new_Jinkela_buffer_16509 (
        .din(new_Jinkela_wire_19699),
        .dout(new_Jinkela_wire_19700)
    );

    bfr new_Jinkela_buffer_16409 (
        .din(new_Jinkela_wire_19597),
        .dout(new_Jinkela_wire_19598)
    );

    spl2 new_Jinkela_splitter_1451 (
        .a(_1754_),
        .b(new_Jinkela_wire_19788),
        .c(new_Jinkela_wire_19789)
    );

    bfr new_Jinkela_buffer_16410 (
        .din(new_Jinkela_wire_19598),
        .dout(new_Jinkela_wire_19599)
    );

    spl2 new_Jinkela_splitter_1450 (
        .a(_1206_),
        .b(new_Jinkela_wire_19786),
        .c(new_Jinkela_wire_19787)
    );

    bfr new_Jinkela_buffer_16510 (
        .din(new_Jinkela_wire_19700),
        .dout(new_Jinkela_wire_19701)
    );

    bfr new_Jinkela_buffer_16411 (
        .din(new_Jinkela_wire_19599),
        .dout(new_Jinkela_wire_19600)
    );

    bfr new_Jinkela_buffer_16545 (
        .din(new_Jinkela_wire_19743),
        .dout(new_Jinkela_wire_19744)
    );

    bfr new_Jinkela_buffer_16412 (
        .din(new_Jinkela_wire_19600),
        .dout(new_Jinkela_wire_19601)
    );

    bfr new_Jinkela_buffer_16511 (
        .din(new_Jinkela_wire_19701),
        .dout(new_Jinkela_wire_19702)
    );

    bfr new_Jinkela_buffer_16413 (
        .din(new_Jinkela_wire_19601),
        .dout(new_Jinkela_wire_19602)
    );

    bfr new_Jinkela_buffer_16583 (
        .din(_0476_),
        .dout(new_Jinkela_wire_19790)
    );

    bfr new_Jinkela_buffer_16414 (
        .din(new_Jinkela_wire_19602),
        .dout(new_Jinkela_wire_19603)
    );

    bfr new_Jinkela_buffer_16512 (
        .din(new_Jinkela_wire_19702),
        .dout(new_Jinkela_wire_19703)
    );

    bfr new_Jinkela_buffer_16415 (
        .din(new_Jinkela_wire_19603),
        .dout(new_Jinkela_wire_19604)
    );

    bfr new_Jinkela_buffer_16546 (
        .din(new_Jinkela_wire_19744),
        .dout(new_Jinkela_wire_19745)
    );

    bfr new_Jinkela_buffer_16416 (
        .din(new_Jinkela_wire_19604),
        .dout(new_Jinkela_wire_19605)
    );

    bfr new_Jinkela_buffer_16542 (
        .din(_1698_),
        .dout(new_Jinkela_wire_19741)
    );

    bfr new_Jinkela_buffer_2582 (
        .din(new_Jinkela_wire_3601),
        .dout(new_Jinkela_wire_3602)
    );

    bfr new_Jinkela_buffer_9634 (
        .din(new_Jinkela_wire_11733),
        .dout(new_Jinkela_wire_11734)
    );

    bfr new_Jinkela_buffer_2662 (
        .din(new_Jinkela_wire_3689),
        .dout(new_Jinkela_wire_3690)
    );

    bfr new_Jinkela_buffer_9490 (
        .din(new_Jinkela_wire_11577),
        .dout(new_Jinkela_wire_11578)
    );

    bfr new_Jinkela_buffer_2583 (
        .din(new_Jinkela_wire_3602),
        .dout(new_Jinkela_wire_3603)
    );

    bfr new_Jinkela_buffer_9542 (
        .din(new_Jinkela_wire_11635),
        .dout(new_Jinkela_wire_11636)
    );

    spl2 new_Jinkela_splitter_373 (
        .a(_0826_),
        .b(new_Jinkela_wire_3819),
        .c(new_Jinkela_wire_3820)
    );

    bfr new_Jinkela_buffer_9491 (
        .din(new_Jinkela_wire_11578),
        .dout(new_Jinkela_wire_11579)
    );

    spl2 new_Jinkela_splitter_375 (
        .a(_1393_),
        .b(new_Jinkela_wire_3880),
        .c(new_Jinkela_wire_3881)
    );

    bfr new_Jinkela_buffer_2584 (
        .din(new_Jinkela_wire_3603),
        .dout(new_Jinkela_wire_3604)
    );

    bfr new_Jinkela_buffer_9725 (
        .din(new_Jinkela_wire_11832),
        .dout(new_Jinkela_wire_11833)
    );

    bfr new_Jinkela_buffer_2663 (
        .din(new_Jinkela_wire_3690),
        .dout(new_Jinkela_wire_3691)
    );

    bfr new_Jinkela_buffer_9492 (
        .din(new_Jinkela_wire_11579),
        .dout(new_Jinkela_wire_11580)
    );

    bfr new_Jinkela_buffer_2585 (
        .din(new_Jinkela_wire_3604),
        .dout(new_Jinkela_wire_3605)
    );

    bfr new_Jinkela_buffer_9543 (
        .din(new_Jinkela_wire_11636),
        .dout(new_Jinkela_wire_11637)
    );

    bfr new_Jinkela_buffer_2682 (
        .din(new_Jinkela_wire_3725),
        .dout(new_Jinkela_wire_3726)
    );

    bfr new_Jinkela_buffer_9493 (
        .din(new_Jinkela_wire_11580),
        .dout(new_Jinkela_wire_11581)
    );

    bfr new_Jinkela_buffer_2586 (
        .din(new_Jinkela_wire_3605),
        .dout(new_Jinkela_wire_3606)
    );

    bfr new_Jinkela_buffer_9635 (
        .din(new_Jinkela_wire_11734),
        .dout(new_Jinkela_wire_11735)
    );

    bfr new_Jinkela_buffer_2664 (
        .din(new_Jinkela_wire_3691),
        .dout(new_Jinkela_wire_3692)
    );

    bfr new_Jinkela_buffer_9494 (
        .din(new_Jinkela_wire_11581),
        .dout(new_Jinkela_wire_11582)
    );

    bfr new_Jinkela_buffer_2587 (
        .din(new_Jinkela_wire_3606),
        .dout(new_Jinkela_wire_3607)
    );

    bfr new_Jinkela_buffer_9544 (
        .din(new_Jinkela_wire_11637),
        .dout(new_Jinkela_wire_11638)
    );

    bfr new_Jinkela_buffer_9495 (
        .din(new_Jinkela_wire_11582),
        .dout(new_Jinkela_wire_11583)
    );

    bfr new_Jinkela_buffer_2588 (
        .din(new_Jinkela_wire_3607),
        .dout(new_Jinkela_wire_3608)
    );

    bfr new_Jinkela_buffer_9730 (
        .din(_0767_),
        .dout(new_Jinkela_wire_11840)
    );

    bfr new_Jinkela_buffer_2665 (
        .din(new_Jinkela_wire_3692),
        .dout(new_Jinkela_wire_3693)
    );

    bfr new_Jinkela_buffer_9496 (
        .din(new_Jinkela_wire_11583),
        .dout(new_Jinkela_wire_11584)
    );

    bfr new_Jinkela_buffer_2589 (
        .din(new_Jinkela_wire_3608),
        .dout(new_Jinkela_wire_3609)
    );

    bfr new_Jinkela_buffer_9545 (
        .din(new_Jinkela_wire_11638),
        .dout(new_Jinkela_wire_11639)
    );

    bfr new_Jinkela_buffer_2683 (
        .din(new_Jinkela_wire_3726),
        .dout(new_Jinkela_wire_3727)
    );

    bfr new_Jinkela_buffer_9497 (
        .din(new_Jinkela_wire_11584),
        .dout(new_Jinkela_wire_11585)
    );

    bfr new_Jinkela_buffer_2590 (
        .din(new_Jinkela_wire_3609),
        .dout(new_Jinkela_wire_3610)
    );

    bfr new_Jinkela_buffer_9636 (
        .din(new_Jinkela_wire_11735),
        .dout(new_Jinkela_wire_11736)
    );

    bfr new_Jinkela_buffer_2666 (
        .din(new_Jinkela_wire_3693),
        .dout(new_Jinkela_wire_3694)
    );

    bfr new_Jinkela_buffer_9498 (
        .din(new_Jinkela_wire_11585),
        .dout(new_Jinkela_wire_11586)
    );

    bfr new_Jinkela_buffer_2591 (
        .din(new_Jinkela_wire_3610),
        .dout(new_Jinkela_wire_3611)
    );

    bfr new_Jinkela_buffer_9546 (
        .din(new_Jinkela_wire_11639),
        .dout(new_Jinkela_wire_11640)
    );

    bfr new_Jinkela_buffer_9499 (
        .din(new_Jinkela_wire_11586),
        .dout(new_Jinkela_wire_11587)
    );

    bfr new_Jinkela_buffer_2771 (
        .din(_0447_),
        .dout(new_Jinkela_wire_3821)
    );

    bfr new_Jinkela_buffer_2592 (
        .din(new_Jinkela_wire_3611),
        .dout(new_Jinkela_wire_3612)
    );

    bfr new_Jinkela_buffer_9726 (
        .din(new_Jinkela_wire_11833),
        .dout(new_Jinkela_wire_11834)
    );

    bfr new_Jinkela_buffer_2667 (
        .din(new_Jinkela_wire_3694),
        .dout(new_Jinkela_wire_3695)
    );

    bfr new_Jinkela_buffer_9500 (
        .din(new_Jinkela_wire_11587),
        .dout(new_Jinkela_wire_11588)
    );

    bfr new_Jinkela_buffer_2593 (
        .din(new_Jinkela_wire_3612),
        .dout(new_Jinkela_wire_3613)
    );

    bfr new_Jinkela_buffer_9547 (
        .din(new_Jinkela_wire_11640),
        .dout(new_Jinkela_wire_11641)
    );

    bfr new_Jinkela_buffer_2684 (
        .din(new_Jinkela_wire_3727),
        .dout(new_Jinkela_wire_3728)
    );

    bfr new_Jinkela_buffer_9501 (
        .din(new_Jinkela_wire_11588),
        .dout(new_Jinkela_wire_11589)
    );

    bfr new_Jinkela_buffer_2594 (
        .din(new_Jinkela_wire_3613),
        .dout(new_Jinkela_wire_3614)
    );

    bfr new_Jinkela_buffer_9637 (
        .din(new_Jinkela_wire_11736),
        .dout(new_Jinkela_wire_11737)
    );

    bfr new_Jinkela_buffer_2668 (
        .din(new_Jinkela_wire_3695),
        .dout(new_Jinkela_wire_3696)
    );

    bfr new_Jinkela_buffer_9502 (
        .din(new_Jinkela_wire_11589),
        .dout(new_Jinkela_wire_11590)
    );

    bfr new_Jinkela_buffer_2595 (
        .din(new_Jinkela_wire_3614),
        .dout(new_Jinkela_wire_3615)
    );

    bfr new_Jinkela_buffer_9548 (
        .din(new_Jinkela_wire_11641),
        .dout(new_Jinkela_wire_11642)
    );

    bfr new_Jinkela_buffer_9503 (
        .din(new_Jinkela_wire_11590),
        .dout(new_Jinkela_wire_11591)
    );

    bfr new_Jinkela_buffer_2827 (
        .din(_1303_),
        .dout(new_Jinkela_wire_3879)
    );

    bfr new_Jinkela_buffer_2596 (
        .din(new_Jinkela_wire_3615),
        .dout(new_Jinkela_wire_3616)
    );

    bfr new_Jinkela_buffer_9842 (
        .din(_1650_),
        .dout(new_Jinkela_wire_11954)
    );

    bfr new_Jinkela_buffer_2669 (
        .din(new_Jinkela_wire_3696),
        .dout(new_Jinkela_wire_3697)
    );

    bfr new_Jinkela_buffer_9504 (
        .din(new_Jinkela_wire_11591),
        .dout(new_Jinkela_wire_11592)
    );

    bfr new_Jinkela_buffer_2597 (
        .din(new_Jinkela_wire_3616),
        .dout(new_Jinkela_wire_3617)
    );

    bfr new_Jinkela_buffer_9549 (
        .din(new_Jinkela_wire_11642),
        .dout(new_Jinkela_wire_11643)
    );

    bfr new_Jinkela_buffer_2685 (
        .din(new_Jinkela_wire_3728),
        .dout(new_Jinkela_wire_3729)
    );

    bfr new_Jinkela_buffer_9505 (
        .din(new_Jinkela_wire_11592),
        .dout(new_Jinkela_wire_11593)
    );

    bfr new_Jinkela_buffer_2598 (
        .din(new_Jinkela_wire_3617),
        .dout(new_Jinkela_wire_3618)
    );

    bfr new_Jinkela_buffer_9638 (
        .din(new_Jinkela_wire_11737),
        .dout(new_Jinkela_wire_11738)
    );

    bfr new_Jinkela_buffer_2670 (
        .din(new_Jinkela_wire_3697),
        .dout(new_Jinkela_wire_3698)
    );

    bfr new_Jinkela_buffer_9506 (
        .din(new_Jinkela_wire_11593),
        .dout(new_Jinkela_wire_11594)
    );

    bfr new_Jinkela_buffer_2599 (
        .din(new_Jinkela_wire_3618),
        .dout(new_Jinkela_wire_3619)
    );

    bfr new_Jinkela_buffer_9550 (
        .din(new_Jinkela_wire_11643),
        .dout(new_Jinkela_wire_11644)
    );

    bfr new_Jinkela_buffer_2772 (
        .din(new_Jinkela_wire_3821),
        .dout(new_Jinkela_wire_3822)
    );

    bfr new_Jinkela_buffer_9507 (
        .din(new_Jinkela_wire_11594),
        .dout(new_Jinkela_wire_11595)
    );

    bfr new_Jinkela_buffer_2600 (
        .din(new_Jinkela_wire_3619),
        .dout(new_Jinkela_wire_3620)
    );

    bfr new_Jinkela_buffer_9727 (
        .din(new_Jinkela_wire_11834),
        .dout(new_Jinkela_wire_11835)
    );

    spl2 new_Jinkela_splitter_363 (
        .a(new_Jinkela_wire_3698),
        .b(new_Jinkela_wire_3699),
        .c(new_Jinkela_wire_3700)
    );

    bfr new_Jinkela_buffer_9508 (
        .din(new_Jinkela_wire_11595),
        .dout(new_Jinkela_wire_11596)
    );

    bfr new_Jinkela_buffer_2601 (
        .din(new_Jinkela_wire_3620),
        .dout(new_Jinkela_wire_3621)
    );

    bfr new_Jinkela_buffer_9551 (
        .din(new_Jinkela_wire_11644),
        .dout(new_Jinkela_wire_11645)
    );

    spl2 new_Jinkela_splitter_376 (
        .a(_0520_),
        .b(new_Jinkela_wire_3886),
        .c(new_Jinkela_wire_3887)
    );

    bfr new_Jinkela_buffer_9509 (
        .din(new_Jinkela_wire_11596),
        .dout(new_Jinkela_wire_11597)
    );

    bfr new_Jinkela_buffer_2602 (
        .din(new_Jinkela_wire_3621),
        .dout(new_Jinkela_wire_3622)
    );

    bfr new_Jinkela_buffer_9639 (
        .din(new_Jinkela_wire_11738),
        .dout(new_Jinkela_wire_11739)
    );

    bfr new_Jinkela_buffer_2686 (
        .din(new_Jinkela_wire_3729),
        .dout(new_Jinkela_wire_3730)
    );

    bfr new_Jinkela_buffer_9510 (
        .din(new_Jinkela_wire_11597),
        .dout(new_Jinkela_wire_11598)
    );

    bfr new_Jinkela_buffer_6021 (
        .din(new_Jinkela_wire_7636),
        .dout(new_Jinkela_wire_7637)
    );

    bfr new_Jinkela_buffer_6096 (
        .din(new_Jinkela_wire_7753),
        .dout(new_Jinkela_wire_7754)
    );

    bfr new_Jinkela_buffer_6022 (
        .din(new_Jinkela_wire_7637),
        .dout(new_Jinkela_wire_7638)
    );

    bfr new_Jinkela_buffer_6174 (
        .din(new_Jinkela_wire_7837),
        .dout(new_Jinkela_wire_7838)
    );

    bfr new_Jinkela_buffer_6023 (
        .din(new_Jinkela_wire_7638),
        .dout(new_Jinkela_wire_7639)
    );

    bfr new_Jinkela_buffer_6097 (
        .din(new_Jinkela_wire_7754),
        .dout(new_Jinkela_wire_7755)
    );

    bfr new_Jinkela_buffer_6024 (
        .din(new_Jinkela_wire_7639),
        .dout(new_Jinkela_wire_7640)
    );

    bfr new_Jinkela_buffer_6178 (
        .din(_0080_),
        .dout(new_Jinkela_wire_7844)
    );

    bfr new_Jinkela_buffer_6025 (
        .din(new_Jinkela_wire_7640),
        .dout(new_Jinkela_wire_7641)
    );

    bfr new_Jinkela_buffer_6098 (
        .din(new_Jinkela_wire_7755),
        .dout(new_Jinkela_wire_7756)
    );

    bfr new_Jinkela_buffer_6026 (
        .din(new_Jinkela_wire_7641),
        .dout(new_Jinkela_wire_7642)
    );

    bfr new_Jinkela_buffer_6200 (
        .din(_0886_),
        .dout(new_Jinkela_wire_7874)
    );

    bfr new_Jinkela_buffer_6027 (
        .din(new_Jinkela_wire_7642),
        .dout(new_Jinkela_wire_7643)
    );

    bfr new_Jinkela_buffer_6099 (
        .din(new_Jinkela_wire_7756),
        .dout(new_Jinkela_wire_7757)
    );

    bfr new_Jinkela_buffer_6028 (
        .din(new_Jinkela_wire_7643),
        .dout(new_Jinkela_wire_7644)
    );

    bfr new_Jinkela_buffer_6175 (
        .din(new_Jinkela_wire_7838),
        .dout(new_Jinkela_wire_7839)
    );

    bfr new_Jinkela_buffer_6029 (
        .din(new_Jinkela_wire_7644),
        .dout(new_Jinkela_wire_7645)
    );

    bfr new_Jinkela_buffer_6100 (
        .din(new_Jinkela_wire_7757),
        .dout(new_Jinkela_wire_7758)
    );

    bfr new_Jinkela_buffer_6030 (
        .din(new_Jinkela_wire_7645),
        .dout(new_Jinkela_wire_7646)
    );

    spl2 new_Jinkela_splitter_683 (
        .a(_1788_),
        .b(new_Jinkela_wire_7847),
        .c(new_Jinkela_wire_7848)
    );

    spl2 new_Jinkela_splitter_682 (
        .a(_0175_),
        .b(new_Jinkela_wire_7845),
        .c(new_Jinkela_wire_7846)
    );

    bfr new_Jinkela_buffer_6031 (
        .din(new_Jinkela_wire_7646),
        .dout(new_Jinkela_wire_7647)
    );

    bfr new_Jinkela_buffer_6101 (
        .din(new_Jinkela_wire_7758),
        .dout(new_Jinkela_wire_7759)
    );

    bfr new_Jinkela_buffer_6032 (
        .din(new_Jinkela_wire_7647),
        .dout(new_Jinkela_wire_7648)
    );

    bfr new_Jinkela_buffer_6176 (
        .din(new_Jinkela_wire_7839),
        .dout(new_Jinkela_wire_7840)
    );

    bfr new_Jinkela_buffer_6033 (
        .din(new_Jinkela_wire_7648),
        .dout(new_Jinkela_wire_7649)
    );

    bfr new_Jinkela_buffer_6102 (
        .din(new_Jinkela_wire_7759),
        .dout(new_Jinkela_wire_7760)
    );

    bfr new_Jinkela_buffer_6034 (
        .din(new_Jinkela_wire_7649),
        .dout(new_Jinkela_wire_7650)
    );

    bfr new_Jinkela_buffer_6035 (
        .din(new_Jinkela_wire_7650),
        .dout(new_Jinkela_wire_7651)
    );

    bfr new_Jinkela_buffer_6103 (
        .din(new_Jinkela_wire_7760),
        .dout(new_Jinkela_wire_7761)
    );

    bfr new_Jinkela_buffer_6036 (
        .din(new_Jinkela_wire_7651),
        .dout(new_Jinkela_wire_7652)
    );

    bfr new_Jinkela_buffer_6177 (
        .din(new_Jinkela_wire_7840),
        .dout(new_Jinkela_wire_7841)
    );

    bfr new_Jinkela_buffer_6037 (
        .din(new_Jinkela_wire_7652),
        .dout(new_Jinkela_wire_7653)
    );

    bfr new_Jinkela_buffer_6104 (
        .din(new_Jinkela_wire_7761),
        .dout(new_Jinkela_wire_7762)
    );

    bfr new_Jinkela_buffer_6038 (
        .din(new_Jinkela_wire_7653),
        .dout(new_Jinkela_wire_7654)
    );

    bfr new_Jinkela_buffer_6179 (
        .din(_1028_),
        .dout(new_Jinkela_wire_7849)
    );

    bfr new_Jinkela_buffer_6039 (
        .din(new_Jinkela_wire_7654),
        .dout(new_Jinkela_wire_7655)
    );

    bfr new_Jinkela_buffer_6105 (
        .din(new_Jinkela_wire_7762),
        .dout(new_Jinkela_wire_7763)
    );

    bfr new_Jinkela_buffer_6040 (
        .din(new_Jinkela_wire_7655),
        .dout(new_Jinkela_wire_7656)
    );

    spl2 new_Jinkela_splitter_685 (
        .a(_1784_),
        .b(new_Jinkela_wire_7868),
        .c(new_Jinkela_wire_7869)
    );

    bfr new_Jinkela_buffer_6041 (
        .din(new_Jinkela_wire_7656),
        .dout(new_Jinkela_wire_7657)
    );

    bfr new_Jinkela_buffer_6106 (
        .din(new_Jinkela_wire_7763),
        .dout(new_Jinkela_wire_7764)
    );

    bfr new_Jinkela_buffer_2603 (
        .din(new_Jinkela_wire_3622),
        .dout(new_Jinkela_wire_3623)
    );

    bfr new_Jinkela_buffer_2687 (
        .din(new_Jinkela_wire_3730),
        .dout(new_Jinkela_wire_3731)
    );

    bfr new_Jinkela_buffer_2604 (
        .din(new_Jinkela_wire_3623),
        .dout(new_Jinkela_wire_3624)
    );

    bfr new_Jinkela_buffer_2773 (
        .din(new_Jinkela_wire_3822),
        .dout(new_Jinkela_wire_3823)
    );

    bfr new_Jinkela_buffer_2605 (
        .din(new_Jinkela_wire_3624),
        .dout(new_Jinkela_wire_3625)
    );

    bfr new_Jinkela_buffer_2688 (
        .din(new_Jinkela_wire_3731),
        .dout(new_Jinkela_wire_3732)
    );

    bfr new_Jinkela_buffer_2606 (
        .din(new_Jinkela_wire_3625),
        .dout(new_Jinkela_wire_3626)
    );

    bfr new_Jinkela_buffer_2828 (
        .din(new_Jinkela_wire_3881),
        .dout(new_Jinkela_wire_3882)
    );

    bfr new_Jinkela_buffer_2607 (
        .din(new_Jinkela_wire_3626),
        .dout(new_Jinkela_wire_3627)
    );

    bfr new_Jinkela_buffer_2689 (
        .din(new_Jinkela_wire_3732),
        .dout(new_Jinkela_wire_3733)
    );

    bfr new_Jinkela_buffer_2608 (
        .din(new_Jinkela_wire_3627),
        .dout(new_Jinkela_wire_3628)
    );

    bfr new_Jinkela_buffer_2774 (
        .din(new_Jinkela_wire_3823),
        .dout(new_Jinkela_wire_3824)
    );

    bfr new_Jinkela_buffer_2609 (
        .din(new_Jinkela_wire_3628),
        .dout(new_Jinkela_wire_3629)
    );

    bfr new_Jinkela_buffer_2690 (
        .din(new_Jinkela_wire_3733),
        .dout(new_Jinkela_wire_3734)
    );

    bfr new_Jinkela_buffer_2610 (
        .din(new_Jinkela_wire_3629),
        .dout(new_Jinkela_wire_3630)
    );

    spl2 new_Jinkela_splitter_377 (
        .a(_1498_),
        .b(new_Jinkela_wire_3888),
        .c(new_Jinkela_wire_3889)
    );

    bfr new_Jinkela_buffer_2611 (
        .din(new_Jinkela_wire_3630),
        .dout(new_Jinkela_wire_3631)
    );

    bfr new_Jinkela_buffer_2691 (
        .din(new_Jinkela_wire_3734),
        .dout(new_Jinkela_wire_3735)
    );

    bfr new_Jinkela_buffer_2612 (
        .din(new_Jinkela_wire_3631),
        .dout(new_Jinkela_wire_3632)
    );

    bfr new_Jinkela_buffer_2775 (
        .din(new_Jinkela_wire_3824),
        .dout(new_Jinkela_wire_3825)
    );

    bfr new_Jinkela_buffer_2613 (
        .din(new_Jinkela_wire_3632),
        .dout(new_Jinkela_wire_3633)
    );

    bfr new_Jinkela_buffer_2692 (
        .din(new_Jinkela_wire_3735),
        .dout(new_Jinkela_wire_3736)
    );

    bfr new_Jinkela_buffer_2614 (
        .din(new_Jinkela_wire_3633),
        .dout(new_Jinkela_wire_3634)
    );

    bfr new_Jinkela_buffer_2615 (
        .din(new_Jinkela_wire_3634),
        .dout(new_Jinkela_wire_3635)
    );

    bfr new_Jinkela_buffer_2693 (
        .din(new_Jinkela_wire_3736),
        .dout(new_Jinkela_wire_3737)
    );

    bfr new_Jinkela_buffer_2616 (
        .din(new_Jinkela_wire_3635),
        .dout(new_Jinkela_wire_3636)
    );

    bfr new_Jinkela_buffer_2776 (
        .din(new_Jinkela_wire_3825),
        .dout(new_Jinkela_wire_3826)
    );

    bfr new_Jinkela_buffer_2617 (
        .din(new_Jinkela_wire_3636),
        .dout(new_Jinkela_wire_3637)
    );

    bfr new_Jinkela_buffer_2694 (
        .din(new_Jinkela_wire_3737),
        .dout(new_Jinkela_wire_3738)
    );

    bfr new_Jinkela_buffer_2618 (
        .din(new_Jinkela_wire_3637),
        .dout(new_Jinkela_wire_3638)
    );

    bfr new_Jinkela_buffer_2829 (
        .din(new_Jinkela_wire_3882),
        .dout(new_Jinkela_wire_3883)
    );

    bfr new_Jinkela_buffer_2619 (
        .din(new_Jinkela_wire_3638),
        .dout(new_Jinkela_wire_3639)
    );

    bfr new_Jinkela_buffer_2695 (
        .din(new_Jinkela_wire_3738),
        .dout(new_Jinkela_wire_3739)
    );

    bfr new_Jinkela_buffer_2620 (
        .din(new_Jinkela_wire_3639),
        .dout(new_Jinkela_wire_3640)
    );

    bfr new_Jinkela_buffer_2777 (
        .din(new_Jinkela_wire_3826),
        .dout(new_Jinkela_wire_3827)
    );

    bfr new_Jinkela_buffer_2621 (
        .din(new_Jinkela_wire_3640),
        .dout(new_Jinkela_wire_3641)
    );

    bfr new_Jinkela_buffer_2696 (
        .din(new_Jinkela_wire_3739),
        .dout(new_Jinkela_wire_3740)
    );

    bfr new_Jinkela_buffer_2622 (
        .din(new_Jinkela_wire_3641),
        .dout(new_Jinkela_wire_3642)
    );

    spl2 new_Jinkela_splitter_379 (
        .a(_0030_),
        .b(new_Jinkela_wire_3892),
        .c(new_Jinkela_wire_3893)
    );

    spl2 new_Jinkela_splitter_378 (
        .a(_1091_),
        .b(new_Jinkela_wire_3890),
        .c(new_Jinkela_wire_3891)
    );

    bfr new_Jinkela_buffer_2623 (
        .din(new_Jinkela_wire_3642),
        .dout(new_Jinkela_wire_3643)
    );

    bfr new_Jinkela_buffer_2697 (
        .din(new_Jinkela_wire_3740),
        .dout(new_Jinkela_wire_3741)
    );

    and_bb _3466_ (
        .a(new_Jinkela_wire_13680),
        .b(new_Jinkela_wire_10950),
        .c(_0757_)
    );

    bfr new_Jinkela_buffer_9552 (
        .din(new_Jinkela_wire_11645),
        .dout(new_Jinkela_wire_11646)
    );

    or_bb _3467_ (
        .a(new_Jinkela_wire_9543),
        .b(new_Jinkela_wire_17860),
        .c(_0758_)
    );

    bfr new_Jinkela_buffer_9511 (
        .din(new_Jinkela_wire_11598),
        .dout(new_Jinkela_wire_11599)
    );

    and_ii _3468_ (
        .a(new_Jinkela_wire_14658),
        .b(new_Jinkela_wire_13681),
        .c(_0759_)
    );

    spl2 new_Jinkela_splitter_905 (
        .a(_0403_),
        .b(new_Jinkela_wire_11955),
        .c(new_Jinkela_wire_11956)
    );

    and_bb _3469_ (
        .a(new_Jinkela_wire_14659),
        .b(new_Jinkela_wire_13682),
        .c(_0760_)
    );

    bfr new_Jinkela_buffer_9512 (
        .din(new_Jinkela_wire_11599),
        .dout(new_Jinkela_wire_11600)
    );

    and_ii _3470_ (
        .a(new_Jinkela_wire_2457),
        .b(new_Jinkela_wire_16874),
        .c(_0761_)
    );

    bfr new_Jinkela_buffer_9553 (
        .din(new_Jinkela_wire_11646),
        .dout(new_Jinkela_wire_11647)
    );

    and_bb _3471_ (
        .a(new_Jinkela_wire_6990),
        .b(new_Jinkela_wire_19120),
        .c(_0762_)
    );

    bfr new_Jinkela_buffer_9513 (
        .din(new_Jinkela_wire_11600),
        .dout(new_Jinkela_wire_11601)
    );

    and_ii _3472_ (
        .a(new_Jinkela_wire_6991),
        .b(new_Jinkela_wire_19121),
        .c(_0763_)
    );

    bfr new_Jinkela_buffer_9640 (
        .din(new_Jinkela_wire_11739),
        .dout(new_Jinkela_wire_11740)
    );

    or_bb _3473_ (
        .a(new_Jinkela_wire_839),
        .b(new_Jinkela_wire_17549),
        .c(new_net_3918)
    );

    bfr new_Jinkela_buffer_9514 (
        .din(new_Jinkela_wire_11601),
        .dout(new_Jinkela_wire_11602)
    );

    or_bb _3474_ (
        .a(new_Jinkela_wire_17550),
        .b(new_Jinkela_wire_16903),
        .c(_0765_)
    );

    bfr new_Jinkela_buffer_9554 (
        .din(new_Jinkela_wire_11647),
        .dout(new_Jinkela_wire_11648)
    );

    and_ii _3475_ (
        .a(new_Jinkela_wire_17861),
        .b(new_Jinkela_wire_7306),
        .c(_0766_)
    );

    bfr new_Jinkela_buffer_9515 (
        .din(new_Jinkela_wire_11602),
        .dout(new_Jinkela_wire_11603)
    );

    and_bb _3476_ (
        .a(new_Jinkela_wire_670),
        .b(new_Jinkela_wire_41),
        .c(_0767_)
    );

    bfr new_Jinkela_buffer_9731 (
        .din(new_Jinkela_wire_11840),
        .dout(new_Jinkela_wire_11841)
    );

    and_ii _3477_ (
        .a(new_Jinkela_wire_18686),
        .b(new_Jinkela_wire_10111),
        .c(_0768_)
    );

    bfr new_Jinkela_buffer_9516 (
        .din(new_Jinkela_wire_11603),
        .dout(new_Jinkela_wire_11604)
    );

    and_bb _3478_ (
        .a(new_Jinkela_wire_197),
        .b(new_Jinkela_wire_528),
        .c(_0769_)
    );

    bfr new_Jinkela_buffer_9555 (
        .din(new_Jinkela_wire_11648),
        .dout(new_Jinkela_wire_11649)
    );

    and_ii _3479_ (
        .a(new_Jinkela_wire_16523),
        .b(new_Jinkela_wire_19340),
        .c(_0770_)
    );

    bfr new_Jinkela_buffer_9517 (
        .din(new_Jinkela_wire_11604),
        .dout(new_Jinkela_wire_11605)
    );

    and_bb _3480_ (
        .a(new_Jinkela_wire_389),
        .b(new_Jinkela_wire_145),
        .c(_0771_)
    );

    bfr new_Jinkela_buffer_9641 (
        .din(new_Jinkela_wire_11740),
        .dout(new_Jinkela_wire_11741)
    );

    and_ii _3481_ (
        .a(new_Jinkela_wire_1335),
        .b(new_Jinkela_wire_16529),
        .c(_0772_)
    );

    bfr new_Jinkela_buffer_9518 (
        .din(new_Jinkela_wire_11605),
        .dout(new_Jinkela_wire_11606)
    );

    and_bb _3482_ (
        .a(new_Jinkela_wire_401),
        .b(new_Jinkela_wire_212),
        .c(_0773_)
    );

    bfr new_Jinkela_buffer_9556 (
        .din(new_Jinkela_wire_11649),
        .dout(new_Jinkela_wire_11650)
    );

    and_ii _3483_ (
        .a(new_Jinkela_wire_10264),
        .b(new_Jinkela_wire_20682),
        .c(_0775_)
    );

    bfr new_Jinkela_buffer_9519 (
        .din(new_Jinkela_wire_11606),
        .dout(new_Jinkela_wire_11607)
    );

    and_bb _3484_ (
        .a(new_Jinkela_wire_168),
        .b(new_Jinkela_wire_583),
        .c(_0776_)
    );

    spl2 new_Jinkela_splitter_906 (
        .a(_1658_),
        .b(new_Jinkela_wire_11957),
        .c(new_Jinkela_wire_11958)
    );

    spl2 new_Jinkela_splitter_908 (
        .a(_1683_),
        .b(new_Jinkela_wire_11961),
        .c(new_Jinkela_wire_11962)
    );

    and_ii _3485_ (
        .a(new_Jinkela_wire_3666),
        .b(new_Jinkela_wire_18288),
        .c(_0777_)
    );

    bfr new_Jinkela_buffer_9520 (
        .din(new_Jinkela_wire_11607),
        .dout(new_Jinkela_wire_11608)
    );

    and_bb _3486_ (
        .a(new_Jinkela_wire_602),
        .b(new_Jinkela_wire_113),
        .c(_0778_)
    );

    bfr new_Jinkela_buffer_9557 (
        .din(new_Jinkela_wire_11650),
        .dout(new_Jinkela_wire_11651)
    );

    and_bb _3487_ (
        .a(new_Jinkela_wire_424),
        .b(new_Jinkela_wire_20),
        .c(_0779_)
    );

    bfr new_Jinkela_buffer_9521 (
        .din(new_Jinkela_wire_11608),
        .dout(new_Jinkela_wire_11609)
    );

    and_ii _3488_ (
        .a(new_Jinkela_wire_10063),
        .b(new_Jinkela_wire_14543),
        .c(_0780_)
    );

    bfr new_Jinkela_buffer_9642 (
        .din(new_Jinkela_wire_11741),
        .dout(new_Jinkela_wire_11742)
    );

    and_ii _3489_ (
        .a(new_Jinkela_wire_7586),
        .b(new_Jinkela_wire_20037),
        .c(_0781_)
    );

    bfr new_Jinkela_buffer_9522 (
        .din(new_Jinkela_wire_11609),
        .dout(new_Jinkela_wire_11610)
    );

    and_bb _3490_ (
        .a(new_Jinkela_wire_7587),
        .b(new_Jinkela_wire_20038),
        .c(_0782_)
    );

    bfr new_Jinkela_buffer_9558 (
        .din(new_Jinkela_wire_11651),
        .dout(new_Jinkela_wire_11652)
    );

    or_bb _3491_ (
        .a(new_Jinkela_wire_18533),
        .b(new_Jinkela_wire_2326),
        .c(_0783_)
    );

    bfr new_Jinkela_buffer_9523 (
        .din(new_Jinkela_wire_11610),
        .dout(new_Jinkela_wire_11611)
    );

    and_ii _3492_ (
        .a(new_Jinkela_wire_21092),
        .b(new_Jinkela_wire_4980),
        .c(_0784_)
    );

    bfr new_Jinkela_buffer_9732 (
        .din(new_Jinkela_wire_11841),
        .dout(new_Jinkela_wire_11842)
    );

    and_bb _3493_ (
        .a(new_Jinkela_wire_21093),
        .b(new_Jinkela_wire_4981),
        .c(_0786_)
    );

    spl2 new_Jinkela_splitter_893 (
        .a(new_Jinkela_wire_11611),
        .b(new_Jinkela_wire_11612),
        .c(new_Jinkela_wire_11613)
    );

    or_bb _3494_ (
        .a(new_Jinkela_wire_2122),
        .b(new_Jinkela_wire_19063),
        .c(_0787_)
    );

    bfr new_Jinkela_buffer_9643 (
        .din(new_Jinkela_wire_11742),
        .dout(new_Jinkela_wire_11743)
    );

    and_ii _3495_ (
        .a(new_Jinkela_wire_5695),
        .b(new_Jinkela_wire_7715),
        .c(_0788_)
    );

    bfr new_Jinkela_buffer_9559 (
        .din(new_Jinkela_wire_11652),
        .dout(new_Jinkela_wire_11653)
    );

    and_bb _3496_ (
        .a(new_Jinkela_wire_5696),
        .b(new_Jinkela_wire_7716),
        .c(_0789_)
    );

    bfr new_Jinkela_buffer_9560 (
        .din(new_Jinkela_wire_11653),
        .dout(new_Jinkela_wire_11654)
    );

    or_bb _3497_ (
        .a(new_Jinkela_wire_4998),
        .b(new_Jinkela_wire_10686),
        .c(_0790_)
    );

    and_ii _3498_ (
        .a(new_Jinkela_wire_5718),
        .b(new_Jinkela_wire_5965),
        .c(_0791_)
    );

    bfr new_Jinkela_buffer_9561 (
        .din(new_Jinkela_wire_11654),
        .dout(new_Jinkela_wire_11655)
    );

    and_bb _3499_ (
        .a(new_Jinkela_wire_5719),
        .b(new_Jinkela_wire_5966),
        .c(_0792_)
    );

    bfr new_Jinkela_buffer_9644 (
        .din(new_Jinkela_wire_11743),
        .dout(new_Jinkela_wire_11744)
    );

    or_bb _3500_ (
        .a(new_Jinkela_wire_1077),
        .b(new_Jinkela_wire_18695),
        .c(_0793_)
    );

    bfr new_Jinkela_buffer_9562 (
        .din(new_Jinkela_wire_11655),
        .dout(new_Jinkela_wire_11656)
    );

    and_ii _3501_ (
        .a(new_Jinkela_wire_5712),
        .b(new_Jinkela_wire_16870),
        .c(_0794_)
    );

    bfr new_Jinkela_buffer_9733 (
        .din(new_Jinkela_wire_11842),
        .dout(new_Jinkela_wire_11843)
    );

    and_bb _3502_ (
        .a(new_Jinkela_wire_5713),
        .b(new_Jinkela_wire_16871),
        .c(_0795_)
    );

    bfr new_Jinkela_buffer_9563 (
        .din(new_Jinkela_wire_11656),
        .dout(new_Jinkela_wire_11657)
    );

    or_bb _3503_ (
        .a(new_Jinkela_wire_1914),
        .b(new_Jinkela_wire_7176),
        .c(_0797_)
    );

    bfr new_Jinkela_buffer_9645 (
        .din(new_Jinkela_wire_11744),
        .dout(new_Jinkela_wire_11745)
    );

    and_ii _3504_ (
        .a(new_Jinkela_wire_14317),
        .b(new_Jinkela_wire_20899),
        .c(_0798_)
    );

    bfr new_Jinkela_buffer_9564 (
        .din(new_Jinkela_wire_11657),
        .dout(new_Jinkela_wire_11658)
    );

    and_bb _3505_ (
        .a(new_Jinkela_wire_14318),
        .b(new_Jinkela_wire_20900),
        .c(_0799_)
    );

    spl2 new_Jinkela_splitter_907 (
        .a(_0172_),
        .b(new_Jinkela_wire_11959),
        .c(new_Jinkela_wire_11960)
    );

    or_bb _3506_ (
        .a(new_Jinkela_wire_4297),
        .b(new_Jinkela_wire_3447),
        .c(_0800_)
    );

    bfr new_Jinkela_buffer_9565 (
        .din(new_Jinkela_wire_11658),
        .dout(new_Jinkela_wire_11659)
    );

    and_ii _3507_ (
        .a(new_Jinkela_wire_19182),
        .b(new_Jinkela_wire_21114),
        .c(_0801_)
    );

    bfr new_Jinkela_buffer_9646 (
        .din(new_Jinkela_wire_11745),
        .dout(new_Jinkela_wire_11746)
    );

    bfr new_Jinkela_buffer_6042 (
        .din(new_Jinkela_wire_7657),
        .dout(new_Jinkela_wire_7658)
    );

    bfr new_Jinkela_buffer_6180 (
        .din(new_Jinkela_wire_7849),
        .dout(new_Jinkela_wire_7850)
    );

    bfr new_Jinkela_buffer_6043 (
        .din(new_Jinkela_wire_7658),
        .dout(new_Jinkela_wire_7659)
    );

    bfr new_Jinkela_buffer_6107 (
        .din(new_Jinkela_wire_7764),
        .dout(new_Jinkela_wire_7765)
    );

    bfr new_Jinkela_buffer_6044 (
        .din(new_Jinkela_wire_7659),
        .dout(new_Jinkela_wire_7660)
    );

    bfr new_Jinkela_buffer_6196 (
        .din(new_Jinkela_wire_7869),
        .dout(new_Jinkela_wire_7870)
    );

    bfr new_Jinkela_buffer_6045 (
        .din(new_Jinkela_wire_7660),
        .dout(new_Jinkela_wire_7661)
    );

    bfr new_Jinkela_buffer_6108 (
        .din(new_Jinkela_wire_7765),
        .dout(new_Jinkela_wire_7766)
    );

    bfr new_Jinkela_buffer_6046 (
        .din(new_Jinkela_wire_7661),
        .dout(new_Jinkela_wire_7662)
    );

    bfr new_Jinkela_buffer_6181 (
        .din(new_Jinkela_wire_7850),
        .dout(new_Jinkela_wire_7851)
    );

    bfr new_Jinkela_buffer_6047 (
        .din(new_Jinkela_wire_7662),
        .dout(new_Jinkela_wire_7663)
    );

    bfr new_Jinkela_buffer_6109 (
        .din(new_Jinkela_wire_7766),
        .dout(new_Jinkela_wire_7767)
    );

    bfr new_Jinkela_buffer_6048 (
        .din(new_Jinkela_wire_7663),
        .dout(new_Jinkela_wire_7664)
    );

    bfr new_Jinkela_buffer_6294 (
        .din(_0460_),
        .dout(new_Jinkela_wire_7970)
    );

    bfr new_Jinkela_buffer_6049 (
        .din(new_Jinkela_wire_7664),
        .dout(new_Jinkela_wire_7665)
    );

    bfr new_Jinkela_buffer_6110 (
        .din(new_Jinkela_wire_7767),
        .dout(new_Jinkela_wire_7768)
    );

    bfr new_Jinkela_buffer_6050 (
        .din(new_Jinkela_wire_7665),
        .dout(new_Jinkela_wire_7666)
    );

    bfr new_Jinkela_buffer_6182 (
        .din(new_Jinkela_wire_7851),
        .dout(new_Jinkela_wire_7852)
    );

    bfr new_Jinkela_buffer_6051 (
        .din(new_Jinkela_wire_7666),
        .dout(new_Jinkela_wire_7667)
    );

    bfr new_Jinkela_buffer_6111 (
        .din(new_Jinkela_wire_7768),
        .dout(new_Jinkela_wire_7769)
    );

    bfr new_Jinkela_buffer_6052 (
        .din(new_Jinkela_wire_7667),
        .dout(new_Jinkela_wire_7668)
    );

    bfr new_Jinkela_buffer_6295 (
        .din(_1772_),
        .dout(new_Jinkela_wire_7971)
    );

    bfr new_Jinkela_buffer_6053 (
        .din(new_Jinkela_wire_7668),
        .dout(new_Jinkela_wire_7669)
    );

    bfr new_Jinkela_buffer_6112 (
        .din(new_Jinkela_wire_7769),
        .dout(new_Jinkela_wire_7770)
    );

    bfr new_Jinkela_buffer_6054 (
        .din(new_Jinkela_wire_7669),
        .dout(new_Jinkela_wire_7670)
    );

    bfr new_Jinkela_buffer_6183 (
        .din(new_Jinkela_wire_7852),
        .dout(new_Jinkela_wire_7853)
    );

    bfr new_Jinkela_buffer_6055 (
        .din(new_Jinkela_wire_7670),
        .dout(new_Jinkela_wire_7671)
    );

    bfr new_Jinkela_buffer_6113 (
        .din(new_Jinkela_wire_7770),
        .dout(new_Jinkela_wire_7771)
    );

    bfr new_Jinkela_buffer_6056 (
        .din(new_Jinkela_wire_7671),
        .dout(new_Jinkela_wire_7672)
    );

    bfr new_Jinkela_buffer_6197 (
        .din(new_Jinkela_wire_7870),
        .dout(new_Jinkela_wire_7871)
    );

    bfr new_Jinkela_buffer_6057 (
        .din(new_Jinkela_wire_7672),
        .dout(new_Jinkela_wire_7673)
    );

    bfr new_Jinkela_buffer_6114 (
        .din(new_Jinkela_wire_7771),
        .dout(new_Jinkela_wire_7772)
    );

    bfr new_Jinkela_buffer_6058 (
        .din(new_Jinkela_wire_7673),
        .dout(new_Jinkela_wire_7674)
    );

    bfr new_Jinkela_buffer_6184 (
        .din(new_Jinkela_wire_7853),
        .dout(new_Jinkela_wire_7854)
    );

    bfr new_Jinkela_buffer_6059 (
        .din(new_Jinkela_wire_7674),
        .dout(new_Jinkela_wire_7675)
    );

    bfr new_Jinkela_buffer_6115 (
        .din(new_Jinkela_wire_7772),
        .dout(new_Jinkela_wire_7773)
    );

    bfr new_Jinkela_buffer_6060 (
        .din(new_Jinkela_wire_7675),
        .dout(new_Jinkela_wire_7676)
    );

    bfr new_Jinkela_buffer_6201 (
        .din(new_Jinkela_wire_7874),
        .dout(new_Jinkela_wire_7875)
    );

    bfr new_Jinkela_buffer_6061 (
        .din(new_Jinkela_wire_7676),
        .dout(new_Jinkela_wire_7677)
    );

    bfr new_Jinkela_buffer_6116 (
        .din(new_Jinkela_wire_7773),
        .dout(new_Jinkela_wire_7774)
    );

    bfr new_Jinkela_buffer_6062 (
        .din(new_Jinkela_wire_7677),
        .dout(new_Jinkela_wire_7678)
    );

    bfr new_Jinkela_buffer_6185 (
        .din(new_Jinkela_wire_7854),
        .dout(new_Jinkela_wire_7855)
    );

    bfr new_Jinkela_buffer_2624 (
        .din(new_Jinkela_wire_3643),
        .dout(new_Jinkela_wire_3644)
    );

    bfr new_Jinkela_buffer_16513 (
        .din(new_Jinkela_wire_19703),
        .dout(new_Jinkela_wire_19704)
    );

    and_bb _1864_ (
        .a(new_Jinkela_wire_5107),
        .b(new_Jinkela_wire_8864),
        .c(_1741_)
    );

    bfr new_Jinkela_buffer_16417 (
        .din(new_Jinkela_wire_19605),
        .dout(new_Jinkela_wire_19606)
    );

    bfr new_Jinkela_buffer_2778 (
        .din(new_Jinkela_wire_3827),
        .dout(new_Jinkela_wire_3828)
    );

    or_bb _1865_ (
        .a(new_Jinkela_wire_4833),
        .b(new_Jinkela_wire_6618),
        .c(_1752_)
    );

    bfr new_Jinkela_buffer_2625 (
        .din(new_Jinkela_wire_3644),
        .dout(new_Jinkela_wire_3645)
    );

    bfr new_Jinkela_buffer_16584 (
        .din(_1052_),
        .dout(new_Jinkela_wire_19793)
    );

    or_bb _1866_ (
        .a(new_Jinkela_wire_4667),
        .b(new_Jinkela_wire_5043),
        .c(_1763_)
    );

    bfr new_Jinkela_buffer_16418 (
        .din(new_Jinkela_wire_19606),
        .dout(new_Jinkela_wire_19607)
    );

    bfr new_Jinkela_buffer_2698 (
        .din(new_Jinkela_wire_3741),
        .dout(new_Jinkela_wire_3742)
    );

    and_bb _1867_ (
        .a(new_Jinkela_wire_4668),
        .b(new_Jinkela_wire_5044),
        .c(_1774_)
    );

    bfr new_Jinkela_buffer_2626 (
        .din(new_Jinkela_wire_3645),
        .dout(new_Jinkela_wire_3646)
    );

    bfr new_Jinkela_buffer_16514 (
        .din(new_Jinkela_wire_19704),
        .dout(new_Jinkela_wire_19705)
    );

    or_bi _1868_ (
        .a(new_Jinkela_wire_8208),
        .b(new_Jinkela_wire_10067),
        .c(_1785_)
    );

    bfr new_Jinkela_buffer_16419 (
        .din(new_Jinkela_wire_19607),
        .dout(new_Jinkela_wire_19608)
    );

    bfr new_Jinkela_buffer_2830 (
        .din(new_Jinkela_wire_3883),
        .dout(new_Jinkela_wire_3884)
    );

    and_ii _1869_ (
        .a(new_Jinkela_wire_7980),
        .b(new_Jinkela_wire_15910),
        .c(_1796_)
    );

    bfr new_Jinkela_buffer_2627 (
        .din(new_Jinkela_wire_3646),
        .dout(new_Jinkela_wire_3647)
    );

    bfr new_Jinkela_buffer_16547 (
        .din(new_Jinkela_wire_19745),
        .dout(new_Jinkela_wire_19746)
    );

    and_bb _1870_ (
        .a(new_Jinkela_wire_7981),
        .b(new_Jinkela_wire_15911),
        .c(_1806_)
    );

    bfr new_Jinkela_buffer_16420 (
        .din(new_Jinkela_wire_19608),
        .dout(new_Jinkela_wire_19609)
    );

    bfr new_Jinkela_buffer_2699 (
        .din(new_Jinkela_wire_3742),
        .dout(new_Jinkela_wire_3743)
    );

    or_bb _1871_ (
        .a(new_Jinkela_wire_16789),
        .b(new_Jinkela_wire_14275),
        .c(new_net_3968)
    );

    bfr new_Jinkela_buffer_2628 (
        .din(new_Jinkela_wire_3647),
        .dout(new_Jinkela_wire_3648)
    );

    bfr new_Jinkela_buffer_16515 (
        .din(new_Jinkela_wire_19705),
        .dout(new_Jinkela_wire_19706)
    );

    and_bb _1872_ (
        .a(new_Jinkela_wire_345),
        .b(new_Jinkela_wire_21),
        .c(_1827_)
    );

    bfr new_Jinkela_buffer_16421 (
        .din(new_Jinkela_wire_19609),
        .dout(new_Jinkela_wire_19610)
    );

    bfr new_Jinkela_buffer_2779 (
        .din(new_Jinkela_wire_3828),
        .dout(new_Jinkela_wire_3829)
    );

    and_bi _1873_ (
        .a(new_Jinkela_wire_10072),
        .b(new_Jinkela_wire_14276),
        .c(_0000_)
    );

    bfr new_Jinkela_buffer_2629 (
        .din(new_Jinkela_wire_3648),
        .dout(new_Jinkela_wire_3649)
    );

    and_bb _1874_ (
        .a(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_631),
        .c(_0011_)
    );

    bfr new_Jinkela_buffer_16422 (
        .din(new_Jinkela_wire_19610),
        .dout(new_Jinkela_wire_19611)
    );

    bfr new_Jinkela_buffer_2700 (
        .din(new_Jinkela_wire_3743),
        .dout(new_Jinkela_wire_3744)
    );

    and_bi _1875_ (
        .a(new_Jinkela_wire_5156),
        .b(new_Jinkela_wire_6619),
        .c(_0022_)
    );

    spl2 new_Jinkela_splitter_1452 (
        .a(_1192_),
        .b(new_Jinkela_wire_19791),
        .c(new_Jinkela_wire_19792)
    );

    bfr new_Jinkela_buffer_2630 (
        .din(new_Jinkela_wire_3649),
        .dout(new_Jinkela_wire_3650)
    );

    bfr new_Jinkela_buffer_16516 (
        .din(new_Jinkela_wire_19706),
        .dout(new_Jinkela_wire_19707)
    );

    and_bb _1876_ (
        .a(new_Jinkela_wire_535),
        .b(new_Jinkela_wire_570),
        .c(_0033_)
    );

    bfr new_Jinkela_buffer_16423 (
        .din(new_Jinkela_wire_19611),
        .dout(new_Jinkela_wire_19612)
    );

    spl2 new_Jinkela_splitter_382 (
        .a(_1144_),
        .b(new_Jinkela_wire_3958),
        .c(new_Jinkela_wire_3959)
    );

    or_ii _1877_ (
        .a(new_Jinkela_wire_79),
        .b(new_Jinkela_wire_309),
        .c(_0044_)
    );

    bfr new_Jinkela_buffer_2631 (
        .din(new_Jinkela_wire_3650),
        .dout(new_Jinkela_wire_3651)
    );

    bfr new_Jinkela_buffer_16548 (
        .din(new_Jinkela_wire_19746),
        .dout(new_Jinkela_wire_19747)
    );

    and_bi _1878_ (
        .a(new_Jinkela_wire_5738),
        .b(new_Jinkela_wire_1286),
        .c(_0055_)
    );

    bfr new_Jinkela_buffer_16424 (
        .din(new_Jinkela_wire_19612),
        .dout(new_Jinkela_wire_19613)
    );

    bfr new_Jinkela_buffer_2701 (
        .din(new_Jinkela_wire_3744),
        .dout(new_Jinkela_wire_3745)
    );

    and_bb _1879_ (
        .a(new_Jinkela_wire_83),
        .b(new_Jinkela_wire_221),
        .c(_0066_)
    );

    bfr new_Jinkela_buffer_2632 (
        .din(new_Jinkela_wire_3651),
        .dout(new_Jinkela_wire_3652)
    );

    bfr new_Jinkela_buffer_16517 (
        .din(new_Jinkela_wire_19707),
        .dout(new_Jinkela_wire_19708)
    );

    and_bi _1880_ (
        .a(new_Jinkela_wire_4714),
        .b(new_Jinkela_wire_10077),
        .c(_0077_)
    );

    bfr new_Jinkela_buffer_16425 (
        .din(new_Jinkela_wire_19613),
        .dout(new_Jinkela_wire_19614)
    );

    bfr new_Jinkela_buffer_2780 (
        .din(new_Jinkela_wire_3829),
        .dout(new_Jinkela_wire_3830)
    );

    and_ii _1881_ (
        .a(new_Jinkela_wire_14429),
        .b(new_Jinkela_wire_8686),
        .c(_0088_)
    );

    bfr new_Jinkela_buffer_2633 (
        .din(new_Jinkela_wire_3652),
        .dout(new_Jinkela_wire_3653)
    );

    or_bb _1882_ (
        .a(new_Jinkela_wire_14202),
        .b(new_Jinkela_wire_6766),
        .c(_0099_)
    );

    bfr new_Jinkela_buffer_16426 (
        .din(new_Jinkela_wire_19614),
        .dout(new_Jinkela_wire_19615)
    );

    bfr new_Jinkela_buffer_2702 (
        .din(new_Jinkela_wire_3745),
        .dout(new_Jinkela_wire_3746)
    );

    or_ii _1883_ (
        .a(new_Jinkela_wire_14203),
        .b(new_Jinkela_wire_6767),
        .c(_0110_)
    );

    bfr new_Jinkela_buffer_2634 (
        .din(new_Jinkela_wire_3653),
        .dout(new_Jinkela_wire_3654)
    );

    bfr new_Jinkela_buffer_16518 (
        .din(new_Jinkela_wire_19708),
        .dout(new_Jinkela_wire_19709)
    );

    or_bb _1887_ (
        .a(new_Jinkela_wire_15028),
        .b(new_Jinkela_wire_3187),
        .c(_0154_)
    );

    bfr new_Jinkela_buffer_16427 (
        .din(new_Jinkela_wire_19615),
        .dout(new_Jinkela_wire_19616)
    );

    bfr new_Jinkela_buffer_2831 (
        .din(new_Jinkela_wire_3884),
        .dout(new_Jinkela_wire_3885)
    );

    or_bb _1888_ (
        .a(new_Jinkela_wire_21206),
        .b(new_Jinkela_wire_11525),
        .c(_0165_)
    );

    bfr new_Jinkela_buffer_2635 (
        .din(new_Jinkela_wire_3654),
        .dout(new_Jinkela_wire_3655)
    );

    bfr new_Jinkela_buffer_16549 (
        .din(new_Jinkela_wire_19747),
        .dout(new_Jinkela_wire_19748)
    );

    or_ii _1889_ (
        .a(new_Jinkela_wire_21207),
        .b(new_Jinkela_wire_11526),
        .c(_0176_)
    );

    bfr new_Jinkela_buffer_16428 (
        .din(new_Jinkela_wire_19616),
        .dout(new_Jinkela_wire_19617)
    );

    bfr new_Jinkela_buffer_2703 (
        .din(new_Jinkela_wire_3746),
        .dout(new_Jinkela_wire_3747)
    );

    or_ii _1890_ (
        .a(new_Jinkela_wire_3720),
        .b(new_Jinkela_wire_17037),
        .c(_0187_)
    );

    bfr new_Jinkela_buffer_2636 (
        .din(new_Jinkela_wire_3655),
        .dout(new_Jinkela_wire_3656)
    );

    bfr new_Jinkela_buffer_16519 (
        .din(new_Jinkela_wire_19709),
        .dout(new_Jinkela_wire_19710)
    );

    and_ii _1891_ (
        .a(new_Jinkela_wire_16906),
        .b(new_Jinkela_wire_8478),
        .c(_0198_)
    );

    bfr new_Jinkela_buffer_16429 (
        .din(new_Jinkela_wire_19617),
        .dout(new_Jinkela_wire_19618)
    );

    bfr new_Jinkela_buffer_2781 (
        .din(new_Jinkela_wire_3830),
        .dout(new_Jinkela_wire_3831)
    );

    and_bb _1892_ (
        .a(new_Jinkela_wire_16907),
        .b(new_Jinkela_wire_8479),
        .c(_0209_)
    );

    bfr new_Jinkela_buffer_2637 (
        .din(new_Jinkela_wire_3656),
        .dout(new_Jinkela_wire_3657)
    );

    or_bb _1893_ (
        .a(new_Jinkela_wire_6362),
        .b(new_Jinkela_wire_14328),
        .c(_0219_)
    );

    bfr new_Jinkela_buffer_16430 (
        .din(new_Jinkela_wire_19618),
        .dout(new_Jinkela_wire_19619)
    );

    bfr new_Jinkela_buffer_2704 (
        .din(new_Jinkela_wire_3747),
        .dout(new_Jinkela_wire_3748)
    );

    or_bb _1894_ (
        .a(new_Jinkela_wire_1275),
        .b(new_Jinkela_wire_4241),
        .c(_0230_)
    );

    bfr new_Jinkela_buffer_16585 (
        .din(_0432_),
        .dout(new_Jinkela_wire_19794)
    );

    bfr new_Jinkela_buffer_2638 (
        .din(new_Jinkela_wire_3657),
        .dout(new_Jinkela_wire_3658)
    );

    bfr new_Jinkela_buffer_16520 (
        .din(new_Jinkela_wire_19710),
        .dout(new_Jinkela_wire_19711)
    );

    and_bb _1895_ (
        .a(new_Jinkela_wire_339),
        .b(new_Jinkela_wire_645),
        .c(_0241_)
    );

    bfr new_Jinkela_buffer_16431 (
        .din(new_Jinkela_wire_19619),
        .dout(new_Jinkela_wire_19620)
    );

    and_bb _1896_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_4242),
        .c(_0252_)
    );

    bfr new_Jinkela_buffer_2832 (
        .din(_1130_),
        .dout(new_Jinkela_wire_3894)
    );

    bfr new_Jinkela_buffer_2639 (
        .din(new_Jinkela_wire_3658),
        .dout(new_Jinkela_wire_3659)
    );

    bfr new_Jinkela_buffer_16550 (
        .din(new_Jinkela_wire_19748),
        .dout(new_Jinkela_wire_19749)
    );

    or_bi _1897_ (
        .a(new_Jinkela_wire_10677),
        .b(new_Jinkela_wire_7275),
        .c(_0263_)
    );

    bfr new_Jinkela_buffer_16432 (
        .din(new_Jinkela_wire_19620),
        .dout(new_Jinkela_wire_19621)
    );

    bfr new_Jinkela_buffer_2705 (
        .din(new_Jinkela_wire_3748),
        .dout(new_Jinkela_wire_3749)
    );

    and_ii _1898_ (
        .a(new_Jinkela_wire_20324),
        .b(new_Jinkela_wire_19958),
        .c(_0274_)
    );

    bfr new_Jinkela_buffer_2640 (
        .din(new_Jinkela_wire_3659),
        .dout(new_Jinkela_wire_3660)
    );

    bfr new_Jinkela_buffer_16521 (
        .din(new_Jinkela_wire_19711),
        .dout(new_Jinkela_wire_19712)
    );

    and_bi _1899_ (
        .a(new_Jinkela_wire_7280),
        .b(new_Jinkela_wire_4671),
        .c(_0285_)
    );

    bfr new_Jinkela_buffer_16433 (
        .din(new_Jinkela_wire_19621),
        .dout(new_Jinkela_wire_19622)
    );

    bfr new_Jinkela_buffer_2782 (
        .din(new_Jinkela_wire_3831),
        .dout(new_Jinkela_wire_3832)
    );

    and_bb _1900_ (
        .a(new_Jinkela_wire_93),
        .b(new_Jinkela_wire_652),
        .c(_0296_)
    );

    spl2 new_Jinkela_splitter_359 (
        .a(new_Jinkela_wire_3660),
        .b(new_Jinkela_wire_3661),
        .c(new_Jinkela_wire_3662)
    );

    and_bi _1901_ (
        .a(new_Jinkela_wire_17042),
        .b(new_Jinkela_wire_14329),
        .c(_0307_)
    );

    bfr new_Jinkela_buffer_16434 (
        .din(new_Jinkela_wire_19622),
        .dout(new_Jinkela_wire_19623)
    );

    and_bb _1902_ (
        .a(new_Jinkela_wire_636),
        .b(new_Jinkela_wire_558),
        .c(_0318_)
    );

    spl2 new_Jinkela_splitter_381 (
        .a(_1798_),
        .b(new_Jinkela_wire_3952),
        .c(new_Jinkela_wire_3953)
    );

    spl2 new_Jinkela_splitter_1455 (
        .a(_0898_),
        .b(new_Jinkela_wire_19911),
        .c(new_Jinkela_wire_19912)
    );

    bfr new_Jinkela_buffer_2706 (
        .din(new_Jinkela_wire_3749),
        .dout(new_Jinkela_wire_3750)
    );

    bfr new_Jinkela_buffer_16522 (
        .din(new_Jinkela_wire_19712),
        .dout(new_Jinkela_wire_19713)
    );

    and_bi _1903_ (
        .a(new_Jinkela_wire_14209),
        .b(new_Jinkela_wire_3188),
        .c(_0328_)
    );

    bfr new_Jinkela_buffer_16435 (
        .din(new_Jinkela_wire_19623),
        .dout(new_Jinkela_wire_19624)
    );

    bfr new_Jinkela_buffer_2707 (
        .din(new_Jinkela_wire_3750),
        .dout(new_Jinkela_wire_3751)
    );

    and_bb _1904_ (
        .a(new_Jinkela_wire_281),
        .b(new_Jinkela_wire_544),
        .c(_0339_)
    );

    bfr new_Jinkela_buffer_2783 (
        .din(new_Jinkela_wire_3832),
        .dout(new_Jinkela_wire_3833)
    );

    bfr new_Jinkela_buffer_16551 (
        .din(new_Jinkela_wire_19749),
        .dout(new_Jinkela_wire_19750)
    );

    or_ii _1905_ (
        .a(new_Jinkela_wire_478),
        .b(new_Jinkela_wire_323),
        .c(_0350_)
    );

    bfr new_Jinkela_buffer_16436 (
        .din(new_Jinkela_wire_19624),
        .dout(new_Jinkela_wire_19625)
    );

    bfr new_Jinkela_buffer_2708 (
        .din(new_Jinkela_wire_3751),
        .dout(new_Jinkela_wire_3752)
    );

    and_bi _1906_ (
        .a(new_Jinkela_wire_10078),
        .b(new_Jinkela_wire_2962),
        .c(_0361_)
    );

    bfr new_Jinkela_buffer_2833 (
        .din(new_Jinkela_wire_3894),
        .dout(new_Jinkela_wire_3895)
    );

    bfr new_Jinkela_buffer_16523 (
        .din(new_Jinkela_wire_19713),
        .dout(new_Jinkela_wire_19714)
    );

    and_bb _1907_ (
        .a(new_Jinkela_wire_482),
        .b(new_Jinkela_wire_226),
        .c(_0372_)
    );

    bfr new_Jinkela_buffer_16437 (
        .din(new_Jinkela_wire_19625),
        .dout(new_Jinkela_wire_19626)
    );

    bfr new_Jinkela_buffer_2709 (
        .din(new_Jinkela_wire_3752),
        .dout(new_Jinkela_wire_3753)
    );

    and_bi _1908_ (
        .a(new_Jinkela_wire_1287),
        .b(new_Jinkela_wire_16116),
        .c(_0383_)
    );

    spl2 new_Jinkela_splitter_1124 (
        .a(_0505_),
        .b(new_Jinkela_wire_15683),
        .c(new_Jinkela_wire_15684)
    );

    spl2 new_Jinkela_splitter_1114 (
        .a(new_Jinkela_wire_15550),
        .b(new_Jinkela_wire_15551),
        .c(new_Jinkela_wire_15552)
    );

    spl2 new_Jinkela_splitter_1125 (
        .a(_0139_),
        .b(new_Jinkela_wire_15685),
        .c(new_Jinkela_wire_15686)
    );

    bfr new_Jinkela_buffer_13033 (
        .din(new_Jinkela_wire_15566),
        .dout(new_Jinkela_wire_15567)
    );

    bfr new_Jinkela_buffer_13034 (
        .din(new_Jinkela_wire_15567),
        .dout(new_Jinkela_wire_15568)
    );

    bfr new_Jinkela_buffer_13129 (
        .din(new_Jinkela_wire_15678),
        .dout(new_Jinkela_wire_15679)
    );

    bfr new_Jinkela_buffer_13035 (
        .din(new_Jinkela_wire_15568),
        .dout(new_Jinkela_wire_15569)
    );

    bfr new_Jinkela_buffer_13036 (
        .din(new_Jinkela_wire_15569),
        .dout(new_Jinkela_wire_15570)
    );

    bfr new_Jinkela_buffer_13130 (
        .din(new_Jinkela_wire_15679),
        .dout(new_Jinkela_wire_15680)
    );

    bfr new_Jinkela_buffer_13037 (
        .din(new_Jinkela_wire_15570),
        .dout(new_Jinkela_wire_15571)
    );

    spl2 new_Jinkela_splitter_1126 (
        .a(_1473_),
        .b(new_Jinkela_wire_15687),
        .c(new_Jinkela_wire_15688)
    );

    bfr new_Jinkela_buffer_13038 (
        .din(new_Jinkela_wire_15571),
        .dout(new_Jinkela_wire_15572)
    );

    bfr new_Jinkela_buffer_13131 (
        .din(new_Jinkela_wire_15680),
        .dout(new_Jinkela_wire_15681)
    );

    bfr new_Jinkela_buffer_13039 (
        .din(new_Jinkela_wire_15572),
        .dout(new_Jinkela_wire_15573)
    );

    spl2 new_Jinkela_splitter_1127 (
        .a(_1713_),
        .b(new_Jinkela_wire_15689),
        .c(new_Jinkela_wire_15690)
    );

    bfr new_Jinkela_buffer_13040 (
        .din(new_Jinkela_wire_15573),
        .dout(new_Jinkela_wire_15574)
    );

    spl2 new_Jinkela_splitter_1128 (
        .a(_0484_),
        .b(new_Jinkela_wire_15695),
        .c(new_Jinkela_wire_15696)
    );

    bfr new_Jinkela_buffer_13041 (
        .din(new_Jinkela_wire_15574),
        .dout(new_Jinkela_wire_15575)
    );

    bfr new_Jinkela_buffer_13133 (
        .din(new_Jinkela_wire_15690),
        .dout(new_Jinkela_wire_15691)
    );

    spl2 new_Jinkela_splitter_1129 (
        .a(_0157_),
        .b(new_Jinkela_wire_15697),
        .c(new_Jinkela_wire_15698)
    );

    bfr new_Jinkela_buffer_13042 (
        .din(new_Jinkela_wire_15575),
        .dout(new_Jinkela_wire_15576)
    );

    bfr new_Jinkela_buffer_13043 (
        .din(new_Jinkela_wire_15576),
        .dout(new_Jinkela_wire_15577)
    );

    bfr new_Jinkela_buffer_13134 (
        .din(new_Jinkela_wire_15691),
        .dout(new_Jinkela_wire_15692)
    );

    bfr new_Jinkela_buffer_13044 (
        .din(new_Jinkela_wire_15577),
        .dout(new_Jinkela_wire_15578)
    );

    bfr new_Jinkela_buffer_13166 (
        .din(_1451_),
        .dout(new_Jinkela_wire_15730)
    );

    bfr new_Jinkela_buffer_13137 (
        .din(_0823_),
        .dout(new_Jinkela_wire_15699)
    );

    bfr new_Jinkela_buffer_13045 (
        .din(new_Jinkela_wire_15578),
        .dout(new_Jinkela_wire_15579)
    );

    bfr new_Jinkela_buffer_13135 (
        .din(new_Jinkela_wire_15692),
        .dout(new_Jinkela_wire_15693)
    );

    bfr new_Jinkela_buffer_13046 (
        .din(new_Jinkela_wire_15579),
        .dout(new_Jinkela_wire_15580)
    );

    bfr new_Jinkela_buffer_13165 (
        .din(_1250_),
        .dout(new_Jinkela_wire_15729)
    );

    bfr new_Jinkela_buffer_13047 (
        .din(new_Jinkela_wire_15580),
        .dout(new_Jinkela_wire_15581)
    );

    bfr new_Jinkela_buffer_13136 (
        .din(new_Jinkela_wire_15693),
        .dout(new_Jinkela_wire_15694)
    );

    bfr new_Jinkela_buffer_13048 (
        .din(new_Jinkela_wire_15581),
        .dout(new_Jinkela_wire_15582)
    );

    bfr new_Jinkela_buffer_13138 (
        .din(new_Jinkela_wire_15699),
        .dout(new_Jinkela_wire_15700)
    );

    bfr new_Jinkela_buffer_13049 (
        .din(new_Jinkela_wire_15582),
        .dout(new_Jinkela_wire_15583)
    );

    spl2 new_Jinkela_splitter_1131 (
        .a(_0622_),
        .b(new_Jinkela_wire_15731),
        .c(new_Jinkela_wire_15732)
    );

    bfr new_Jinkela_buffer_13050 (
        .din(new_Jinkela_wire_15583),
        .dout(new_Jinkela_wire_15584)
    );

    bfr new_Jinkela_buffer_13139 (
        .din(new_Jinkela_wire_15700),
        .dout(new_Jinkela_wire_15701)
    );

    bfr new_Jinkela_buffer_13051 (
        .din(new_Jinkela_wire_15584),
        .dout(new_Jinkela_wire_15585)
    );

    bfr new_Jinkela_buffer_13167 (
        .din(_1543_),
        .dout(new_Jinkela_wire_15733)
    );

    bfr new_Jinkela_buffer_13052 (
        .din(new_Jinkela_wire_15585),
        .dout(new_Jinkela_wire_15586)
    );

    bfr new_Jinkela_buffer_13140 (
        .din(new_Jinkela_wire_15701),
        .dout(new_Jinkela_wire_15702)
    );

    bfr new_Jinkela_buffer_6063 (
        .din(new_Jinkela_wire_7678),
        .dout(new_Jinkela_wire_7679)
    );

    bfr new_Jinkela_buffer_6117 (
        .din(new_Jinkela_wire_7774),
        .dout(new_Jinkela_wire_7775)
    );

    bfr new_Jinkela_buffer_6064 (
        .din(new_Jinkela_wire_7679),
        .dout(new_Jinkela_wire_7680)
    );

    bfr new_Jinkela_buffer_6198 (
        .din(new_Jinkela_wire_7871),
        .dout(new_Jinkela_wire_7872)
    );

    bfr new_Jinkela_buffer_6065 (
        .din(new_Jinkela_wire_7680),
        .dout(new_Jinkela_wire_7681)
    );

    bfr new_Jinkela_buffer_6118 (
        .din(new_Jinkela_wire_7775),
        .dout(new_Jinkela_wire_7776)
    );

    bfr new_Jinkela_buffer_6066 (
        .din(new_Jinkela_wire_7681),
        .dout(new_Jinkela_wire_7682)
    );

    bfr new_Jinkela_buffer_6186 (
        .din(new_Jinkela_wire_7855),
        .dout(new_Jinkela_wire_7856)
    );

    bfr new_Jinkela_buffer_6067 (
        .din(new_Jinkela_wire_7682),
        .dout(new_Jinkela_wire_7683)
    );

    bfr new_Jinkela_buffer_6119 (
        .din(new_Jinkela_wire_7776),
        .dout(new_Jinkela_wire_7777)
    );

    bfr new_Jinkela_buffer_6068 (
        .din(new_Jinkela_wire_7683),
        .dout(new_Jinkela_wire_7684)
    );

    bfr new_Jinkela_buffer_6296 (
        .din(_0912_),
        .dout(new_Jinkela_wire_7972)
    );

    bfr new_Jinkela_buffer_6069 (
        .din(new_Jinkela_wire_7684),
        .dout(new_Jinkela_wire_7685)
    );

    bfr new_Jinkela_buffer_6120 (
        .din(new_Jinkela_wire_7777),
        .dout(new_Jinkela_wire_7778)
    );

    bfr new_Jinkela_buffer_6070 (
        .din(new_Jinkela_wire_7685),
        .dout(new_Jinkela_wire_7686)
    );

    bfr new_Jinkela_buffer_6187 (
        .din(new_Jinkela_wire_7856),
        .dout(new_Jinkela_wire_7857)
    );

    bfr new_Jinkela_buffer_6071 (
        .din(new_Jinkela_wire_7686),
        .dout(new_Jinkela_wire_7687)
    );

    bfr new_Jinkela_buffer_6121 (
        .din(new_Jinkela_wire_7778),
        .dout(new_Jinkela_wire_7779)
    );

    bfr new_Jinkela_buffer_6072 (
        .din(new_Jinkela_wire_7687),
        .dout(new_Jinkela_wire_7688)
    );

    bfr new_Jinkela_buffer_6199 (
        .din(new_Jinkela_wire_7872),
        .dout(new_Jinkela_wire_7873)
    );

    spl2 new_Jinkela_splitter_657 (
        .a(new_Jinkela_wire_7688),
        .b(new_Jinkela_wire_7689),
        .c(new_Jinkela_wire_7690)
    );

    bfr new_Jinkela_buffer_6188 (
        .din(new_Jinkela_wire_7857),
        .dout(new_Jinkela_wire_7858)
    );

    bfr new_Jinkela_buffer_6122 (
        .din(new_Jinkela_wire_7779),
        .dout(new_Jinkela_wire_7780)
    );

    bfr new_Jinkela_buffer_6123 (
        .din(new_Jinkela_wire_7780),
        .dout(new_Jinkela_wire_7781)
    );

    bfr new_Jinkela_buffer_6202 (
        .din(new_Jinkela_wire_7875),
        .dout(new_Jinkela_wire_7876)
    );

    bfr new_Jinkela_buffer_6124 (
        .din(new_Jinkela_wire_7781),
        .dout(new_Jinkela_wire_7782)
    );

    bfr new_Jinkela_buffer_6189 (
        .din(new_Jinkela_wire_7858),
        .dout(new_Jinkela_wire_7859)
    );

    bfr new_Jinkela_buffer_6125 (
        .din(new_Jinkela_wire_7782),
        .dout(new_Jinkela_wire_7783)
    );

    spl2 new_Jinkela_splitter_687 (
        .a(_0078_),
        .b(new_Jinkela_wire_7973),
        .c(new_Jinkela_wire_7974)
    );

    bfr new_Jinkela_buffer_6126 (
        .din(new_Jinkela_wire_7783),
        .dout(new_Jinkela_wire_7784)
    );

    bfr new_Jinkela_buffer_6190 (
        .din(new_Jinkela_wire_7859),
        .dout(new_Jinkela_wire_7860)
    );

    bfr new_Jinkela_buffer_6127 (
        .din(new_Jinkela_wire_7784),
        .dout(new_Jinkela_wire_7785)
    );

    bfr new_Jinkela_buffer_6203 (
        .din(new_Jinkela_wire_7876),
        .dout(new_Jinkela_wire_7877)
    );

    bfr new_Jinkela_buffer_6128 (
        .din(new_Jinkela_wire_7785),
        .dout(new_Jinkela_wire_7786)
    );

    bfr new_Jinkela_buffer_6191 (
        .din(new_Jinkela_wire_7860),
        .dout(new_Jinkela_wire_7861)
    );

    bfr new_Jinkela_buffer_6129 (
        .din(new_Jinkela_wire_7786),
        .dout(new_Jinkela_wire_7787)
    );

    bfr new_Jinkela_buffer_6301 (
        .din(_1037_),
        .dout(new_Jinkela_wire_7979)
    );

    bfr new_Jinkela_buffer_6130 (
        .din(new_Jinkela_wire_7787),
        .dout(new_Jinkela_wire_7788)
    );

    bfr new_Jinkela_buffer_6192 (
        .din(new_Jinkela_wire_7861),
        .dout(new_Jinkela_wire_7862)
    );

    bfr new_Jinkela_buffer_6131 (
        .din(new_Jinkela_wire_7788),
        .dout(new_Jinkela_wire_7789)
    );

    bfr new_Jinkela_buffer_6204 (
        .din(new_Jinkela_wire_7877),
        .dout(new_Jinkela_wire_7878)
    );

    bfr new_Jinkela_buffer_6132 (
        .din(new_Jinkela_wire_7789),
        .dout(new_Jinkela_wire_7790)
    );

    bfr new_Jinkela_buffer_9566 (
        .din(new_Jinkela_wire_11659),
        .dout(new_Jinkela_wire_11660)
    );

    bfr new_Jinkela_buffer_16553 (
        .din(new_Jinkela_wire_19751),
        .dout(new_Jinkela_wire_19752)
    );

    bfr new_Jinkela_buffer_16438 (
        .din(new_Jinkela_wire_19626),
        .dout(new_Jinkela_wire_19627)
    );

    bfr new_Jinkela_buffer_9734 (
        .din(new_Jinkela_wire_11843),
        .dout(new_Jinkela_wire_11844)
    );

    bfr new_Jinkela_buffer_9567 (
        .din(new_Jinkela_wire_11660),
        .dout(new_Jinkela_wire_11661)
    );

    bfr new_Jinkela_buffer_16524 (
        .din(new_Jinkela_wire_19714),
        .dout(new_Jinkela_wire_19715)
    );

    bfr new_Jinkela_buffer_16439 (
        .din(new_Jinkela_wire_19627),
        .dout(new_Jinkela_wire_19628)
    );

    bfr new_Jinkela_buffer_9647 (
        .din(new_Jinkela_wire_11746),
        .dout(new_Jinkela_wire_11747)
    );

    bfr new_Jinkela_buffer_9568 (
        .din(new_Jinkela_wire_11661),
        .dout(new_Jinkela_wire_11662)
    );

    bfr new_Jinkela_buffer_16587 (
        .din(new_Jinkela_wire_19795),
        .dout(new_Jinkela_wire_19796)
    );

    bfr new_Jinkela_buffer_16440 (
        .din(new_Jinkela_wire_19628),
        .dout(new_Jinkela_wire_19629)
    );

    bfr new_Jinkela_buffer_9927 (
        .din(_0506_),
        .dout(new_Jinkela_wire_12051)
    );

    bfr new_Jinkela_buffer_9569 (
        .din(new_Jinkela_wire_11662),
        .dout(new_Jinkela_wire_11663)
    );

    bfr new_Jinkela_buffer_16525 (
        .din(new_Jinkela_wire_19715),
        .dout(new_Jinkela_wire_19716)
    );

    bfr new_Jinkela_buffer_16441 (
        .din(new_Jinkela_wire_19629),
        .dout(new_Jinkela_wire_19630)
    );

    bfr new_Jinkela_buffer_9648 (
        .din(new_Jinkela_wire_11747),
        .dout(new_Jinkela_wire_11748)
    );

    bfr new_Jinkela_buffer_9570 (
        .din(new_Jinkela_wire_11663),
        .dout(new_Jinkela_wire_11664)
    );

    bfr new_Jinkela_buffer_16554 (
        .din(new_Jinkela_wire_19752),
        .dout(new_Jinkela_wire_19753)
    );

    bfr new_Jinkela_buffer_16442 (
        .din(new_Jinkela_wire_19630),
        .dout(new_Jinkela_wire_19631)
    );

    bfr new_Jinkela_buffer_9735 (
        .din(new_Jinkela_wire_11844),
        .dout(new_Jinkela_wire_11845)
    );

    bfr new_Jinkela_buffer_9571 (
        .din(new_Jinkela_wire_11664),
        .dout(new_Jinkela_wire_11665)
    );

    bfr new_Jinkela_buffer_16526 (
        .din(new_Jinkela_wire_19716),
        .dout(new_Jinkela_wire_19717)
    );

    bfr new_Jinkela_buffer_16443 (
        .din(new_Jinkela_wire_19631),
        .dout(new_Jinkela_wire_19632)
    );

    bfr new_Jinkela_buffer_9649 (
        .din(new_Jinkela_wire_11748),
        .dout(new_Jinkela_wire_11749)
    );

    bfr new_Jinkela_buffer_9572 (
        .din(new_Jinkela_wire_11665),
        .dout(new_Jinkela_wire_11666)
    );

    bfr new_Jinkela_buffer_16702 (
        .din(_0135_),
        .dout(new_Jinkela_wire_19917)
    );

    bfr new_Jinkela_buffer_16444 (
        .din(new_Jinkela_wire_19632),
        .dout(new_Jinkela_wire_19633)
    );

    bfr new_Jinkela_buffer_9843 (
        .din(_0705_),
        .dout(new_Jinkela_wire_11963)
    );

    bfr new_Jinkela_buffer_16698 (
        .din(new_Jinkela_wire_19912),
        .dout(new_Jinkela_wire_19913)
    );

    bfr new_Jinkela_buffer_9573 (
        .din(new_Jinkela_wire_11666),
        .dout(new_Jinkela_wire_11667)
    );

    bfr new_Jinkela_buffer_16527 (
        .din(new_Jinkela_wire_19717),
        .dout(new_Jinkela_wire_19718)
    );

    bfr new_Jinkela_buffer_16445 (
        .din(new_Jinkela_wire_19633),
        .dout(new_Jinkela_wire_19634)
    );

    bfr new_Jinkela_buffer_9650 (
        .din(new_Jinkela_wire_11749),
        .dout(new_Jinkela_wire_11750)
    );

    bfr new_Jinkela_buffer_9574 (
        .din(new_Jinkela_wire_11667),
        .dout(new_Jinkela_wire_11668)
    );

    bfr new_Jinkela_buffer_16555 (
        .din(new_Jinkela_wire_19753),
        .dout(new_Jinkela_wire_19754)
    );

    bfr new_Jinkela_buffer_16446 (
        .din(new_Jinkela_wire_19634),
        .dout(new_Jinkela_wire_19635)
    );

    bfr new_Jinkela_buffer_9736 (
        .din(new_Jinkela_wire_11845),
        .dout(new_Jinkela_wire_11846)
    );

    bfr new_Jinkela_buffer_9575 (
        .din(new_Jinkela_wire_11668),
        .dout(new_Jinkela_wire_11669)
    );

    bfr new_Jinkela_buffer_16528 (
        .din(new_Jinkela_wire_19718),
        .dout(new_Jinkela_wire_19719)
    );

    bfr new_Jinkela_buffer_16447 (
        .din(new_Jinkela_wire_19635),
        .dout(new_Jinkela_wire_19636)
    );

    bfr new_Jinkela_buffer_9651 (
        .din(new_Jinkela_wire_11750),
        .dout(new_Jinkela_wire_11751)
    );

    bfr new_Jinkela_buffer_9576 (
        .din(new_Jinkela_wire_11669),
        .dout(new_Jinkela_wire_11670)
    );

    bfr new_Jinkela_buffer_16588 (
        .din(new_Jinkela_wire_19796),
        .dout(new_Jinkela_wire_19797)
    );

    bfr new_Jinkela_buffer_16448 (
        .din(new_Jinkela_wire_19636),
        .dout(new_Jinkela_wire_19637)
    );

    spl2 new_Jinkela_splitter_910 (
        .a(_1659_),
        .b(new_Jinkela_wire_12045),
        .c(new_Jinkela_wire_12046)
    );

    bfr new_Jinkela_buffer_9577 (
        .din(new_Jinkela_wire_11670),
        .dout(new_Jinkela_wire_11671)
    );

    bfr new_Jinkela_buffer_16529 (
        .din(new_Jinkela_wire_19719),
        .dout(new_Jinkela_wire_19720)
    );

    bfr new_Jinkela_buffer_16449 (
        .din(new_Jinkela_wire_19637),
        .dout(new_Jinkela_wire_19638)
    );

    bfr new_Jinkela_buffer_9652 (
        .din(new_Jinkela_wire_11751),
        .dout(new_Jinkela_wire_11752)
    );

    bfr new_Jinkela_buffer_9578 (
        .din(new_Jinkela_wire_11671),
        .dout(new_Jinkela_wire_11672)
    );

    bfr new_Jinkela_buffer_16556 (
        .din(new_Jinkela_wire_19754),
        .dout(new_Jinkela_wire_19755)
    );

    bfr new_Jinkela_buffer_16450 (
        .din(new_Jinkela_wire_19638),
        .dout(new_Jinkela_wire_19639)
    );

    bfr new_Jinkela_buffer_9737 (
        .din(new_Jinkela_wire_11846),
        .dout(new_Jinkela_wire_11847)
    );

    bfr new_Jinkela_buffer_9579 (
        .din(new_Jinkela_wire_11672),
        .dout(new_Jinkela_wire_11673)
    );

    bfr new_Jinkela_buffer_16530 (
        .din(new_Jinkela_wire_19720),
        .dout(new_Jinkela_wire_19721)
    );

    bfr new_Jinkela_buffer_16451 (
        .din(new_Jinkela_wire_19639),
        .dout(new_Jinkela_wire_19640)
    );

    bfr new_Jinkela_buffer_9653 (
        .din(new_Jinkela_wire_11752),
        .dout(new_Jinkela_wire_11753)
    );

    bfr new_Jinkela_buffer_9580 (
        .din(new_Jinkela_wire_11673),
        .dout(new_Jinkela_wire_11674)
    );

    bfr new_Jinkela_buffer_16452 (
        .din(new_Jinkela_wire_19640),
        .dout(new_Jinkela_wire_19641)
    );

    bfr new_Jinkela_buffer_9844 (
        .din(new_Jinkela_wire_11963),
        .dout(new_Jinkela_wire_11964)
    );

    bfr new_Jinkela_buffer_9581 (
        .din(new_Jinkela_wire_11674),
        .dout(new_Jinkela_wire_11675)
    );

    bfr new_Jinkela_buffer_16531 (
        .din(new_Jinkela_wire_19721),
        .dout(new_Jinkela_wire_19722)
    );

    bfr new_Jinkela_buffer_16453 (
        .din(new_Jinkela_wire_19641),
        .dout(new_Jinkela_wire_19642)
    );

    bfr new_Jinkela_buffer_9654 (
        .din(new_Jinkela_wire_11753),
        .dout(new_Jinkela_wire_11754)
    );

    bfr new_Jinkela_buffer_9582 (
        .din(new_Jinkela_wire_11675),
        .dout(new_Jinkela_wire_11676)
    );

    bfr new_Jinkela_buffer_16557 (
        .din(new_Jinkela_wire_19755),
        .dout(new_Jinkela_wire_19756)
    );

    bfr new_Jinkela_buffer_16454 (
        .din(new_Jinkela_wire_19642),
        .dout(new_Jinkela_wire_19643)
    );

    bfr new_Jinkela_buffer_9738 (
        .din(new_Jinkela_wire_11847),
        .dout(new_Jinkela_wire_11848)
    );

    bfr new_Jinkela_buffer_9583 (
        .din(new_Jinkela_wire_11676),
        .dout(new_Jinkela_wire_11677)
    );

    bfr new_Jinkela_buffer_16532 (
        .din(new_Jinkela_wire_19722),
        .dout(new_Jinkela_wire_19723)
    );

    bfr new_Jinkela_buffer_16455 (
        .din(new_Jinkela_wire_19643),
        .dout(new_Jinkela_wire_19644)
    );

    bfr new_Jinkela_buffer_9655 (
        .din(new_Jinkela_wire_11754),
        .dout(new_Jinkela_wire_11755)
    );

    bfr new_Jinkela_buffer_9584 (
        .din(new_Jinkela_wire_11677),
        .dout(new_Jinkela_wire_11678)
    );

    bfr new_Jinkela_buffer_16589 (
        .din(new_Jinkela_wire_19797),
        .dout(new_Jinkela_wire_19798)
    );

    bfr new_Jinkela_buffer_16456 (
        .din(new_Jinkela_wire_19644),
        .dout(new_Jinkela_wire_19645)
    );

    bfr new_Jinkela_buffer_9923 (
        .din(new_Jinkela_wire_12046),
        .dout(new_Jinkela_wire_12047)
    );

    bfr new_Jinkela_buffer_9585 (
        .din(new_Jinkela_wire_11678),
        .dout(new_Jinkela_wire_11679)
    );

    bfr new_Jinkela_buffer_16533 (
        .din(new_Jinkela_wire_19723),
        .dout(new_Jinkela_wire_19724)
    );

    bfr new_Jinkela_buffer_16457 (
        .din(new_Jinkela_wire_19645),
        .dout(new_Jinkela_wire_19646)
    );

    bfr new_Jinkela_buffer_9656 (
        .din(new_Jinkela_wire_11755),
        .dout(new_Jinkela_wire_11756)
    );

    bfr new_Jinkela_buffer_9586 (
        .din(new_Jinkela_wire_11679),
        .dout(new_Jinkela_wire_11680)
    );

    bfr new_Jinkela_buffer_16558 (
        .din(new_Jinkela_wire_19756),
        .dout(new_Jinkela_wire_19757)
    );

    bfr new_Jinkela_buffer_16458 (
        .din(new_Jinkela_wire_19646),
        .dout(new_Jinkela_wire_19647)
    );

    bfr new_Jinkela_buffer_9739 (
        .din(new_Jinkela_wire_11848),
        .dout(new_Jinkela_wire_11849)
    );

    and_bb _3508_ (
        .a(new_Jinkela_wire_19183),
        .b(new_Jinkela_wire_21115),
        .c(_0802_)
    );

    bfr new_Jinkela_buffer_13053 (
        .din(new_Jinkela_wire_15586),
        .dout(new_Jinkela_wire_15587)
    );

    or_bb _3509_ (
        .a(new_Jinkela_wire_8685),
        .b(new_Jinkela_wire_16790),
        .c(_0803_)
    );

    bfr new_Jinkela_buffer_13172 (
        .din(_1110_),
        .dout(new_Jinkela_wire_15740)
    );

    bfr new_Jinkela_buffer_13168 (
        .din(new_Jinkela_wire_15735),
        .dout(new_Jinkela_wire_15736)
    );

    and_ii _3510_ (
        .a(new_Jinkela_wire_12622),
        .b(new_Jinkela_wire_2011),
        .c(_0804_)
    );

    bfr new_Jinkela_buffer_13054 (
        .din(new_Jinkela_wire_15587),
        .dout(new_Jinkela_wire_15588)
    );

    and_bb _3511_ (
        .a(new_Jinkela_wire_12623),
        .b(new_Jinkela_wire_2012),
        .c(_0805_)
    );

    bfr new_Jinkela_buffer_13141 (
        .din(new_Jinkela_wire_15702),
        .dout(new_Jinkela_wire_15703)
    );

    or_bb _3512_ (
        .a(new_Jinkela_wire_19189),
        .b(new_Jinkela_wire_17024),
        .c(_0806_)
    );

    bfr new_Jinkela_buffer_13055 (
        .din(new_Jinkela_wire_15588),
        .dout(new_Jinkela_wire_15589)
    );

    and_ii _3513_ (
        .a(new_Jinkela_wire_21200),
        .b(new_Jinkela_wire_14190),
        .c(_0808_)
    );

    spl2 new_Jinkela_splitter_1132 (
        .a(_0603_),
        .b(new_Jinkela_wire_15734),
        .c(new_Jinkela_wire_15735)
    );

    and_bb _3514_ (
        .a(new_Jinkela_wire_21201),
        .b(new_Jinkela_wire_14191),
        .c(_0809_)
    );

    bfr new_Jinkela_buffer_13056 (
        .din(new_Jinkela_wire_15589),
        .dout(new_Jinkela_wire_15590)
    );

    or_bb _3515_ (
        .a(new_Jinkela_wire_14088),
        .b(new_Jinkela_wire_7320),
        .c(_0810_)
    );

    bfr new_Jinkela_buffer_13142 (
        .din(new_Jinkela_wire_15703),
        .dout(new_Jinkela_wire_15704)
    );

    and_ii _3516_ (
        .a(new_Jinkela_wire_11046),
        .b(new_Jinkela_wire_12327),
        .c(_0811_)
    );

    bfr new_Jinkela_buffer_13057 (
        .din(new_Jinkela_wire_15590),
        .dout(new_Jinkela_wire_15591)
    );

    and_bb _3517_ (
        .a(new_Jinkela_wire_11047),
        .b(new_Jinkela_wire_12328),
        .c(_0812_)
    );

    or_bb _3518_ (
        .a(new_Jinkela_wire_10075),
        .b(new_Jinkela_wire_19732),
        .c(_0813_)
    );

    bfr new_Jinkela_buffer_13058 (
        .din(new_Jinkela_wire_15591),
        .dout(new_Jinkela_wire_15592)
    );

    and_ii _3519_ (
        .a(new_Jinkela_wire_19351),
        .b(new_Jinkela_wire_7514),
        .c(_0814_)
    );

    bfr new_Jinkela_buffer_13143 (
        .din(new_Jinkela_wire_15704),
        .dout(new_Jinkela_wire_15705)
    );

    and_bb _3520_ (
        .a(new_Jinkela_wire_19352),
        .b(new_Jinkela_wire_7515),
        .c(_0815_)
    );

    bfr new_Jinkela_buffer_13059 (
        .din(new_Jinkela_wire_15592),
        .dout(new_Jinkela_wire_15593)
    );

    or_bb _3521_ (
        .a(new_Jinkela_wire_4248),
        .b(new_Jinkela_wire_4321),
        .c(_0816_)
    );

    spl2 new_Jinkela_splitter_1133 (
        .a(_0076_),
        .b(new_Jinkela_wire_15741),
        .c(new_Jinkela_wire_15742)
    );

    and_ii _3522_ (
        .a(new_Jinkela_wire_11527),
        .b(new_Jinkela_wire_11952),
        .c(_0817_)
    );

    bfr new_Jinkela_buffer_13060 (
        .din(new_Jinkela_wire_15593),
        .dout(new_Jinkela_wire_15594)
    );

    and_bb _3523_ (
        .a(new_Jinkela_wire_11528),
        .b(new_Jinkela_wire_11953),
        .c(_0819_)
    );

    bfr new_Jinkela_buffer_13144 (
        .din(new_Jinkela_wire_15705),
        .dout(new_Jinkela_wire_15706)
    );

    or_bb _3524_ (
        .a(new_Jinkela_wire_13954),
        .b(new_Jinkela_wire_16201),
        .c(_0820_)
    );

    bfr new_Jinkela_buffer_13061 (
        .din(new_Jinkela_wire_15594),
        .dout(new_Jinkela_wire_15595)
    );

    and_ii _3525_ (
        .a(new_Jinkela_wire_2150),
        .b(new_Jinkela_wire_13691),
        .c(_0821_)
    );

    spl2 new_Jinkela_splitter_1134 (
        .a(_1372_),
        .b(new_Jinkela_wire_15743),
        .c(new_Jinkela_wire_15744)
    );

    spl2 new_Jinkela_splitter_1135 (
        .a(_1221_),
        .b(new_Jinkela_wire_15747),
        .c(new_Jinkela_wire_15748)
    );

    and_bb _3526_ (
        .a(new_Jinkela_wire_2151),
        .b(new_Jinkela_wire_13692),
        .c(_0822_)
    );

    bfr new_Jinkela_buffer_13062 (
        .din(new_Jinkela_wire_15595),
        .dout(new_Jinkela_wire_15596)
    );

    and_ii _3527_ (
        .a(new_Jinkela_wire_8177),
        .b(new_Jinkela_wire_6204),
        .c(_0823_)
    );

    bfr new_Jinkela_buffer_13145 (
        .din(new_Jinkela_wire_15706),
        .dout(new_Jinkela_wire_15707)
    );

    and_bb _3528_ (
        .a(new_Jinkela_wire_15727),
        .b(new_Jinkela_wire_5548),
        .c(_0824_)
    );

    bfr new_Jinkela_buffer_13063 (
        .din(new_Jinkela_wire_15596),
        .dout(new_Jinkela_wire_15597)
    );

    and_ii _3529_ (
        .a(new_Jinkela_wire_15728),
        .b(new_Jinkela_wire_5549),
        .c(_0825_)
    );

    bfr new_Jinkela_buffer_13169 (
        .din(new_Jinkela_wire_15736),
        .dout(new_Jinkela_wire_15737)
    );

    or_bb _3530_ (
        .a(new_Jinkela_wire_5421),
        .b(new_Jinkela_wire_7744),
        .c(new_net_3946)
    );

    bfr new_Jinkela_buffer_13064 (
        .din(new_Jinkela_wire_15597),
        .dout(new_Jinkela_wire_15598)
    );

    or_bb _3531_ (
        .a(new_Jinkela_wire_7745),
        .b(new_Jinkela_wire_6237),
        .c(_0826_)
    );

    bfr new_Jinkela_buffer_13146 (
        .din(new_Jinkela_wire_15707),
        .dout(new_Jinkela_wire_15708)
    );

    and_ii _3532_ (
        .a(new_Jinkela_wire_16202),
        .b(new_Jinkela_wire_4326),
        .c(_0827_)
    );

    bfr new_Jinkela_buffer_13065 (
        .din(new_Jinkela_wire_15598),
        .dout(new_Jinkela_wire_15599)
    );

    and_bb _3533_ (
        .a(new_Jinkela_wire_184),
        .b(new_Jinkela_wire_665),
        .c(_0829_)
    );

    and_ii _3534_ (
        .a(new_Jinkela_wire_19733),
        .b(new_Jinkela_wire_7325),
        .c(_0830_)
    );

    bfr new_Jinkela_buffer_13066 (
        .din(new_Jinkela_wire_15599),
        .dout(new_Jinkela_wire_15600)
    );

    and_bb _3535_ (
        .a(new_Jinkela_wire_380),
        .b(new_Jinkela_wire_511),
        .c(_0831_)
    );

    bfr new_Jinkela_buffer_13147 (
        .din(new_Jinkela_wire_15708),
        .dout(new_Jinkela_wire_15709)
    );

    and_ii _3536_ (
        .a(new_Jinkela_wire_17025),
        .b(new_Jinkela_wire_16795),
        .c(_0832_)
    );

    bfr new_Jinkela_buffer_13067 (
        .din(new_Jinkela_wire_15600),
        .dout(new_Jinkela_wire_15601)
    );

    and_bb _3537_ (
        .a(new_Jinkela_wire_398),
        .b(new_Jinkela_wire_150),
        .c(_0833_)
    );

    bfr new_Jinkela_buffer_13170 (
        .din(new_Jinkela_wire_15737),
        .dout(new_Jinkela_wire_15738)
    );

    and_ii _3538_ (
        .a(new_Jinkela_wire_3448),
        .b(new_Jinkela_wire_7181),
        .c(_0834_)
    );

    bfr new_Jinkela_buffer_13068 (
        .din(new_Jinkela_wire_15601),
        .dout(new_Jinkela_wire_15602)
    );

    and_bb _3539_ (
        .a(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_218),
        .c(_0835_)
    );

    bfr new_Jinkela_buffer_13148 (
        .din(new_Jinkela_wire_15709),
        .dout(new_Jinkela_wire_15710)
    );

    and_ii _3540_ (
        .a(new_Jinkela_wire_18696),
        .b(new_Jinkela_wire_10691),
        .c(_0836_)
    );

    bfr new_Jinkela_buffer_13069 (
        .din(new_Jinkela_wire_15602),
        .dout(new_Jinkela_wire_15603)
    );

    and_bb _3541_ (
        .a(new_Jinkela_wire_613),
        .b(new_Jinkela_wire_581),
        .c(_0837_)
    );

    bfr new_Jinkela_buffer_13173 (
        .din(_0486_),
        .dout(new_Jinkela_wire_15745)
    );

    and_bb _3542_ (
        .a(new_Jinkela_wire_422),
        .b(new_Jinkela_wire_128),
        .c(_0838_)
    );

    bfr new_Jinkela_buffer_13070 (
        .din(new_Jinkela_wire_15603),
        .dout(new_Jinkela_wire_15604)
    );

    and_ii _3543_ (
        .a(new_Jinkela_wire_19064),
        .b(new_Jinkela_wire_2331),
        .c(_0840_)
    );

    bfr new_Jinkela_buffer_13149 (
        .din(new_Jinkela_wire_15710),
        .dout(new_Jinkela_wire_15711)
    );

    and_ii _3544_ (
        .a(new_Jinkela_wire_21175),
        .b(new_Jinkela_wire_8836),
        .c(_0841_)
    );

    bfr new_Jinkela_buffer_13071 (
        .din(new_Jinkela_wire_15604),
        .dout(new_Jinkela_wire_15605)
    );

    and_bb _3545_ (
        .a(new_Jinkela_wire_21176),
        .b(new_Jinkela_wire_8837),
        .c(_0842_)
    );

    bfr new_Jinkela_buffer_13171 (
        .din(new_Jinkela_wire_15738),
        .dout(new_Jinkela_wire_15739)
    );

    or_bb _3546_ (
        .a(new_Jinkela_wire_11444),
        .b(new_Jinkela_wire_1608),
        .c(_0843_)
    );

    bfr new_Jinkela_buffer_13072 (
        .din(new_Jinkela_wire_15605),
        .dout(new_Jinkela_wire_15606)
    );

    and_ii _3547_ (
        .a(new_Jinkela_wire_2126),
        .b(new_Jinkela_wire_8175),
        .c(_0844_)
    );

    bfr new_Jinkela_buffer_13150 (
        .din(new_Jinkela_wire_15711),
        .dout(new_Jinkela_wire_15712)
    );

    and_bb _3548_ (
        .a(new_Jinkela_wire_2127),
        .b(new_Jinkela_wire_8176),
        .c(_0845_)
    );

    bfr new_Jinkela_buffer_13073 (
        .din(new_Jinkela_wire_15606),
        .dout(new_Jinkela_wire_15607)
    );

    or_bb _3549_ (
        .a(new_Jinkela_wire_18525),
        .b(new_Jinkela_wire_7748),
        .c(_0846_)
    );

    bfr new_Jinkela_buffer_13174 (
        .din(_0868_),
        .dout(new_Jinkela_wire_15746)
    );

    bfr new_Jinkela_buffer_13074 (
        .din(new_Jinkela_wire_15607),
        .dout(new_Jinkela_wire_15608)
    );

    bfr new_Jinkela_buffer_16534 (
        .din(new_Jinkela_wire_19724),
        .dout(new_Jinkela_wire_19725)
    );

    and_ii _1909_ (
        .a(new_Jinkela_wire_1790),
        .b(new_Jinkela_wire_21146),
        .c(_0394_)
    );

    bfr new_Jinkela_buffer_16459 (
        .din(new_Jinkela_wire_19647),
        .dout(new_Jinkela_wire_19648)
    );

    bfr new_Jinkela_buffer_13151 (
        .din(new_Jinkela_wire_15712),
        .dout(new_Jinkela_wire_15713)
    );

    or_bb _1910_ (
        .a(new_Jinkela_wire_13462),
        .b(new_Jinkela_wire_8690),
        .c(_0405_)
    );

    bfr new_Jinkela_buffer_13075 (
        .din(new_Jinkela_wire_15608),
        .dout(new_Jinkela_wire_15609)
    );

    or_ii _1911_ (
        .a(new_Jinkela_wire_13463),
        .b(new_Jinkela_wire_8689),
        .c(_0416_)
    );

    bfr new_Jinkela_buffer_16460 (
        .din(new_Jinkela_wire_19648),
        .dout(new_Jinkela_wire_19649)
    );

    bfr new_Jinkela_buffer_13176 (
        .din(_0273_),
        .dout(new_Jinkela_wire_15752)
    );

    or_ii _1912_ (
        .a(new_Jinkela_wire_15760),
        .b(new_Jinkela_wire_18387),
        .c(_0427_)
    );

    bfr new_Jinkela_buffer_16703 (
        .din(_1759_),
        .dout(new_Jinkela_wire_19918)
    );

    bfr new_Jinkela_buffer_13076 (
        .din(new_Jinkela_wire_15609),
        .dout(new_Jinkela_wire_15610)
    );

    bfr new_Jinkela_buffer_16535 (
        .din(new_Jinkela_wire_19725),
        .dout(new_Jinkela_wire_19726)
    );

    and_ii _1913_ (
        .a(new_Jinkela_wire_20905),
        .b(new_Jinkela_wire_17371),
        .c(_0437_)
    );

    bfr new_Jinkela_buffer_16461 (
        .din(new_Jinkela_wire_19649),
        .dout(new_Jinkela_wire_19650)
    );

    bfr new_Jinkela_buffer_13152 (
        .din(new_Jinkela_wire_15713),
        .dout(new_Jinkela_wire_15714)
    );

    and_bb _1914_ (
        .a(new_Jinkela_wire_20906),
        .b(new_Jinkela_wire_17372),
        .c(_0448_)
    );

    bfr new_Jinkela_buffer_13077 (
        .din(new_Jinkela_wire_15610),
        .dout(new_Jinkela_wire_15611)
    );

    bfr new_Jinkela_buffer_16559 (
        .din(new_Jinkela_wire_19757),
        .dout(new_Jinkela_wire_19758)
    );

    or_bb _1915_ (
        .a(new_Jinkela_wire_16908),
        .b(new_Jinkela_wire_3444),
        .c(_0459_)
    );

    bfr new_Jinkela_buffer_16462 (
        .din(new_Jinkela_wire_19650),
        .dout(new_Jinkela_wire_19651)
    );

    or_bb _1916_ (
        .a(new_Jinkela_wire_10675),
        .b(new_Jinkela_wire_10558),
        .c(_0470_)
    );

    bfr new_Jinkela_buffer_13078 (
        .din(new_Jinkela_wire_15611),
        .dout(new_Jinkela_wire_15612)
    );

    bfr new_Jinkela_buffer_16536 (
        .din(new_Jinkela_wire_19726),
        .dout(new_Jinkela_wire_19727)
    );

    or_ii _1917_ (
        .a(new_Jinkela_wire_10676),
        .b(new_Jinkela_wire_10559),
        .c(_0481_)
    );

    bfr new_Jinkela_buffer_16463 (
        .din(new_Jinkela_wire_19651),
        .dout(new_Jinkela_wire_19652)
    );

    bfr new_Jinkela_buffer_13153 (
        .din(new_Jinkela_wire_15714),
        .dout(new_Jinkela_wire_15715)
    );

    or_ii _1918_ (
        .a(new_Jinkela_wire_702),
        .b(new_Jinkela_wire_4989),
        .c(_0492_)
    );

    bfr new_Jinkela_buffer_13079 (
        .din(new_Jinkela_wire_15612),
        .dout(new_Jinkela_wire_15613)
    );

    bfr new_Jinkela_buffer_16590 (
        .din(new_Jinkela_wire_19798),
        .dout(new_Jinkela_wire_19799)
    );

    and_ii _1919_ (
        .a(new_Jinkela_wire_4911),
        .b(new_Jinkela_wire_19180),
        .c(_0503_)
    );

    bfr new_Jinkela_buffer_16464 (
        .din(new_Jinkela_wire_19652),
        .dout(new_Jinkela_wire_19653)
    );

    bfr new_Jinkela_buffer_13177 (
        .din(_0072_),
        .dout(new_Jinkela_wire_15753)
    );

    and_bb _1920_ (
        .a(new_Jinkela_wire_4912),
        .b(new_Jinkela_wire_19181),
        .c(_0514_)
    );

    bfr new_Jinkela_buffer_13175 (
        .din(new_Jinkela_wire_15748),
        .dout(new_Jinkela_wire_15749)
    );

    bfr new_Jinkela_buffer_13080 (
        .din(new_Jinkela_wire_15613),
        .dout(new_Jinkela_wire_15614)
    );

    bfr new_Jinkela_buffer_16537 (
        .din(new_Jinkela_wire_19727),
        .dout(new_Jinkela_wire_19728)
    );

    or_bb _1921_ (
        .a(new_Jinkela_wire_7582),
        .b(new_Jinkela_wire_4249),
        .c(_0525_)
    );

    bfr new_Jinkela_buffer_16465 (
        .din(new_Jinkela_wire_19653),
        .dout(new_Jinkela_wire_19654)
    );

    bfr new_Jinkela_buffer_13154 (
        .din(new_Jinkela_wire_15715),
        .dout(new_Jinkela_wire_15716)
    );

    or_bb _1922_ (
        .a(new_Jinkela_wire_2013),
        .b(new_Jinkela_wire_14022),
        .c(_0535_)
    );

    bfr new_Jinkela_buffer_13081 (
        .din(new_Jinkela_wire_15614),
        .dout(new_Jinkela_wire_15615)
    );

    bfr new_Jinkela_buffer_16560 (
        .din(new_Jinkela_wire_19758),
        .dout(new_Jinkela_wire_19759)
    );

    or_ii _1923_ (
        .a(new_Jinkela_wire_2014),
        .b(new_Jinkela_wire_14023),
        .c(_0546_)
    );

    bfr new_Jinkela_buffer_16466 (
        .din(new_Jinkela_wire_19654),
        .dout(new_Jinkela_wire_19655)
    );

    spl2 new_Jinkela_splitter_1137 (
        .a(_1147_),
        .b(new_Jinkela_wire_15754),
        .c(new_Jinkela_wire_15755)
    );

    or_ii _1924_ (
        .a(new_Jinkela_wire_12524),
        .b(new_Jinkela_wire_19320),
        .c(_0557_)
    );

    bfr new_Jinkela_buffer_13082 (
        .din(new_Jinkela_wire_15615),
        .dout(new_Jinkela_wire_15616)
    );

    bfr new_Jinkela_buffer_16538 (
        .din(new_Jinkela_wire_19728),
        .dout(new_Jinkela_wire_19729)
    );

    and_ii _1925_ (
        .a(new_Jinkela_wire_7294),
        .b(new_Jinkela_wire_15551),
        .c(_0568_)
    );

    bfr new_Jinkela_buffer_16467 (
        .din(new_Jinkela_wire_19655),
        .dout(new_Jinkela_wire_19656)
    );

    bfr new_Jinkela_buffer_13155 (
        .din(new_Jinkela_wire_15716),
        .dout(new_Jinkela_wire_15717)
    );

    and_bb _1926_ (
        .a(new_Jinkela_wire_7295),
        .b(new_Jinkela_wire_15552),
        .c(_0579_)
    );

    bfr new_Jinkela_buffer_13083 (
        .din(new_Jinkela_wire_15616),
        .dout(new_Jinkela_wire_15617)
    );

    or_bb _1927_ (
        .a(new_Jinkela_wire_19163),
        .b(new_Jinkela_wire_14014),
        .c(_0590_)
    );

    bfr new_Jinkela_buffer_16468 (
        .din(new_Jinkela_wire_19656),
        .dout(new_Jinkela_wire_19657)
    );

    spl2 new_Jinkela_splitter_1138 (
        .a(_0068_),
        .b(new_Jinkela_wire_15756),
        .c(new_Jinkela_wire_15757)
    );

    or_bb _1928_ (
        .a(new_Jinkela_wire_20369),
        .b(new_Jinkela_wire_13958),
        .c(_0601_)
    );

    spl2 new_Jinkela_splitter_1136 (
        .a(new_Jinkela_wire_15749),
        .b(new_Jinkela_wire_15750),
        .c(new_Jinkela_wire_15751)
    );

    spl2 new_Jinkela_splitter_1456 (
        .a(_0925_),
        .b(new_Jinkela_wire_19919),
        .c(new_Jinkela_wire_19920)
    );

    bfr new_Jinkela_buffer_13084 (
        .din(new_Jinkela_wire_15617),
        .dout(new_Jinkela_wire_15618)
    );

    bfr new_Jinkela_buffer_16539 (
        .din(new_Jinkela_wire_19729),
        .dout(new_Jinkela_wire_19730)
    );

    and_bb _1929_ (
        .a(new_Jinkela_wire_53),
        .b(new_Jinkela_wire_344),
        .c(_0612_)
    );

    bfr new_Jinkela_buffer_16469 (
        .din(new_Jinkela_wire_19657),
        .dout(new_Jinkela_wire_19658)
    );

    bfr new_Jinkela_buffer_13156 (
        .din(new_Jinkela_wire_15717),
        .dout(new_Jinkela_wire_15718)
    );

    and_bb _1930_ (
        .a(new_Jinkela_wire_20370),
        .b(new_Jinkela_wire_13959),
        .c(_0632_)
    );

    bfr new_Jinkela_buffer_13085 (
        .din(new_Jinkela_wire_15618),
        .dout(new_Jinkela_wire_15619)
    );

    bfr new_Jinkela_buffer_16561 (
        .din(new_Jinkela_wire_19759),
        .dout(new_Jinkela_wire_19760)
    );

    or_bi _1931_ (
        .a(new_Jinkela_wire_14009),
        .b(new_Jinkela_wire_18277),
        .c(_0633_)
    );

    bfr new_Jinkela_buffer_16470 (
        .din(new_Jinkela_wire_19658),
        .dout(new_Jinkela_wire_19659)
    );

    and_ii _1932_ (
        .a(new_Jinkela_wire_1773),
        .b(new_Jinkela_wire_6844),
        .c(_0644_)
    );

    bfr new_Jinkela_buffer_13086 (
        .din(new_Jinkela_wire_15619),
        .dout(new_Jinkela_wire_15620)
    );

    bfr new_Jinkela_buffer_16591 (
        .din(new_Jinkela_wire_19799),
        .dout(new_Jinkela_wire_19800)
    );

    and_bi _1933_ (
        .a(new_Jinkela_wire_18282),
        .b(new_Jinkela_wire_19116),
        .c(_0655_)
    );

    bfr new_Jinkela_buffer_16471 (
        .din(new_Jinkela_wire_19659),
        .dout(new_Jinkela_wire_19660)
    );

    bfr new_Jinkela_buffer_13157 (
        .din(new_Jinkela_wire_15718),
        .dout(new_Jinkela_wire_15719)
    );

    and_bb _1934_ (
        .a(new_Jinkela_wire_99),
        .b(new_Jinkela_wire_60),
        .c(_0666_)
    );

    bfr new_Jinkela_buffer_13087 (
        .din(new_Jinkela_wire_15620),
        .dout(new_Jinkela_wire_15621)
    );

    bfr new_Jinkela_buffer_16562 (
        .din(new_Jinkela_wire_19760),
        .dout(new_Jinkela_wire_19761)
    );

    and_bi _1935_ (
        .a(new_Jinkela_wire_19325),
        .b(new_Jinkela_wire_14015),
        .c(_0677_)
    );

    bfr new_Jinkela_buffer_16472 (
        .din(new_Jinkela_wire_19660),
        .dout(new_Jinkela_wire_19661)
    );

    and_bb _1936_ (
        .a(new_Jinkela_wire_653),
        .b(new_Jinkela_wire_569),
        .c(_0688_)
    );

    bfr new_Jinkela_buffer_13088 (
        .din(new_Jinkela_wire_15621),
        .dout(new_Jinkela_wire_15622)
    );

    bfr new_Jinkela_buffer_16699 (
        .din(new_Jinkela_wire_19913),
        .dout(new_Jinkela_wire_19914)
    );

    and_bi _1937_ (
        .a(new_Jinkela_wire_4994),
        .b(new_Jinkela_wire_4250),
        .c(_0698_)
    );

    bfr new_Jinkela_buffer_16473 (
        .din(new_Jinkela_wire_19661),
        .dout(new_Jinkela_wire_19662)
    );

    bfr new_Jinkela_buffer_13158 (
        .din(new_Jinkela_wire_15719),
        .dout(new_Jinkela_wire_15720)
    );

    and_bb _1938_ (
        .a(new_Jinkela_wire_266),
        .b(new_Jinkela_wire_623),
        .c(_0709_)
    );

    bfr new_Jinkela_buffer_13089 (
        .din(new_Jinkela_wire_15622),
        .dout(new_Jinkela_wire_15623)
    );

    bfr new_Jinkela_buffer_16563 (
        .din(new_Jinkela_wire_19761),
        .dout(new_Jinkela_wire_19762)
    );

    and_bi _1939_ (
        .a(new_Jinkela_wire_18392),
        .b(new_Jinkela_wire_3445),
        .c(_0720_)
    );

    bfr new_Jinkela_buffer_16474 (
        .din(new_Jinkela_wire_19662),
        .dout(new_Jinkela_wire_19663)
    );

    and_bb _1940_ (
        .a(new_Jinkela_wire_85),
        .b(new_Jinkela_wire_530),
        .c(_0731_)
    );

    spl2 new_Jinkela_splitter_1139 (
        .a(_1340_),
        .b(new_Jinkela_wire_15758),
        .c(new_Jinkela_wire_15759)
    );

    bfr new_Jinkela_buffer_13090 (
        .din(new_Jinkela_wire_15623),
        .dout(new_Jinkela_wire_15624)
    );

    bfr new_Jinkela_buffer_16592 (
        .din(new_Jinkela_wire_19800),
        .dout(new_Jinkela_wire_19801)
    );

    or_ii _1941_ (
        .a(new_Jinkela_wire_365),
        .b(new_Jinkela_wire_326),
        .c(_0742_)
    );

    bfr new_Jinkela_buffer_16475 (
        .din(new_Jinkela_wire_19663),
        .dout(new_Jinkela_wire_19664)
    );

    bfr new_Jinkela_buffer_13159 (
        .din(new_Jinkela_wire_15720),
        .dout(new_Jinkela_wire_15721)
    );

    and_bi _1942_ (
        .a(new_Jinkela_wire_16117),
        .b(new_Jinkela_wire_15777),
        .c(_0753_)
    );

    bfr new_Jinkela_buffer_13091 (
        .din(new_Jinkela_wire_15624),
        .dout(new_Jinkela_wire_15625)
    );

    bfr new_Jinkela_buffer_16564 (
        .din(new_Jinkela_wire_19762),
        .dout(new_Jinkela_wire_19763)
    );

    and_bb _1943_ (
        .a(new_Jinkela_wire_366),
        .b(new_Jinkela_wire_235),
        .c(_0764_)
    );

    bfr new_Jinkela_buffer_16476 (
        .din(new_Jinkela_wire_19664),
        .dout(new_Jinkela_wire_19665)
    );

    and_bi _1944_ (
        .a(new_Jinkela_wire_2963),
        .b(new_Jinkela_wire_7726),
        .c(_0774_)
    );

    bfr new_Jinkela_buffer_13178 (
        .din(_0416_),
        .dout(new_Jinkela_wire_15760)
    );

    bfr new_Jinkela_buffer_13092 (
        .din(new_Jinkela_wire_15625),
        .dout(new_Jinkela_wire_15626)
    );

    spl2 new_Jinkela_splitter_1457 (
        .a(_1478_),
        .b(new_Jinkela_wire_19925),
        .c(new_Jinkela_wire_19926)
    );

    and_ii _1945_ (
        .a(new_Jinkela_wire_10451),
        .b(new_Jinkela_wire_5045),
        .c(_0785_)
    );

    bfr new_Jinkela_buffer_16477 (
        .din(new_Jinkela_wire_19665),
        .dout(new_Jinkela_wire_19666)
    );

    bfr new_Jinkela_buffer_13160 (
        .din(new_Jinkela_wire_15721),
        .dout(new_Jinkela_wire_15722)
    );

    or_bb _1946_ (
        .a(new_Jinkela_wire_7701),
        .b(new_Jinkela_wire_21149),
        .c(_0796_)
    );

    bfr new_Jinkela_buffer_13093 (
        .din(new_Jinkela_wire_15626),
        .dout(new_Jinkela_wire_15627)
    );

    bfr new_Jinkela_buffer_16565 (
        .din(new_Jinkela_wire_19763),
        .dout(new_Jinkela_wire_19764)
    );

    or_ii _1947_ (
        .a(new_Jinkela_wire_7702),
        .b(new_Jinkela_wire_21150),
        .c(_0807_)
    );

    bfr new_Jinkela_buffer_16478 (
        .din(new_Jinkela_wire_19666),
        .dout(new_Jinkela_wire_19667)
    );

    spl2 new_Jinkela_splitter_1141 (
        .a(_0674_),
        .b(new_Jinkela_wire_15771),
        .c(new_Jinkela_wire_15772)
    );

    or_ii _1948_ (
        .a(new_Jinkela_wire_705),
        .b(new_Jinkela_wire_21184),
        .c(_0818_)
    );

    bfr new_Jinkela_buffer_13179 (
        .din(_1030_),
        .dout(new_Jinkela_wire_15761)
    );

    bfr new_Jinkela_buffer_13094 (
        .din(new_Jinkela_wire_15627),
        .dout(new_Jinkela_wire_15628)
    );

    bfr new_Jinkela_buffer_16593 (
        .din(new_Jinkela_wire_19801),
        .dout(new_Jinkela_wire_19802)
    );

    and_ii _1949_ (
        .a(new_Jinkela_wire_16190),
        .b(new_Jinkela_wire_6533),
        .c(_0828_)
    );

    bfr new_Jinkela_buffer_16479 (
        .din(new_Jinkela_wire_19667),
        .dout(new_Jinkela_wire_19668)
    );

    bfr new_Jinkela_buffer_13161 (
        .din(new_Jinkela_wire_15722),
        .dout(new_Jinkela_wire_15723)
    );

    and_bb _1950_ (
        .a(new_Jinkela_wire_16191),
        .b(new_Jinkela_wire_6534),
        .c(_0839_)
    );

    bfr new_Jinkela_buffer_9587 (
        .din(new_Jinkela_wire_11680),
        .dout(new_Jinkela_wire_11681)
    );

    bfr new_Jinkela_buffer_9657 (
        .din(new_Jinkela_wire_11756),
        .dout(new_Jinkela_wire_11757)
    );

    bfr new_Jinkela_buffer_9588 (
        .din(new_Jinkela_wire_11681),
        .dout(new_Jinkela_wire_11682)
    );

    bfr new_Jinkela_buffer_9845 (
        .din(new_Jinkela_wire_11964),
        .dout(new_Jinkela_wire_11965)
    );

    bfr new_Jinkela_buffer_9589 (
        .din(new_Jinkela_wire_11682),
        .dout(new_Jinkela_wire_11683)
    );

    bfr new_Jinkela_buffer_9658 (
        .din(new_Jinkela_wire_11757),
        .dout(new_Jinkela_wire_11758)
    );

    bfr new_Jinkela_buffer_9590 (
        .din(new_Jinkela_wire_11683),
        .dout(new_Jinkela_wire_11684)
    );

    bfr new_Jinkela_buffer_9740 (
        .din(new_Jinkela_wire_11849),
        .dout(new_Jinkela_wire_11850)
    );

    bfr new_Jinkela_buffer_9591 (
        .din(new_Jinkela_wire_11684),
        .dout(new_Jinkela_wire_11685)
    );

    bfr new_Jinkela_buffer_9659 (
        .din(new_Jinkela_wire_11758),
        .dout(new_Jinkela_wire_11759)
    );

    bfr new_Jinkela_buffer_9592 (
        .din(new_Jinkela_wire_11685),
        .dout(new_Jinkela_wire_11686)
    );

    spl2 new_Jinkela_splitter_911 (
        .a(_0341_),
        .b(new_Jinkela_wire_12052),
        .c(new_Jinkela_wire_12053)
    );

    bfr new_Jinkela_buffer_9593 (
        .din(new_Jinkela_wire_11686),
        .dout(new_Jinkela_wire_11687)
    );

    bfr new_Jinkela_buffer_9660 (
        .din(new_Jinkela_wire_11759),
        .dout(new_Jinkela_wire_11760)
    );

    bfr new_Jinkela_buffer_9594 (
        .din(new_Jinkela_wire_11687),
        .dout(new_Jinkela_wire_11688)
    );

    bfr new_Jinkela_buffer_9741 (
        .din(new_Jinkela_wire_11850),
        .dout(new_Jinkela_wire_11851)
    );

    bfr new_Jinkela_buffer_9595 (
        .din(new_Jinkela_wire_11688),
        .dout(new_Jinkela_wire_11689)
    );

    bfr new_Jinkela_buffer_9661 (
        .din(new_Jinkela_wire_11760),
        .dout(new_Jinkela_wire_11761)
    );

    bfr new_Jinkela_buffer_9596 (
        .din(new_Jinkela_wire_11689),
        .dout(new_Jinkela_wire_11690)
    );

    bfr new_Jinkela_buffer_9846 (
        .din(new_Jinkela_wire_11965),
        .dout(new_Jinkela_wire_11966)
    );

    bfr new_Jinkela_buffer_9597 (
        .din(new_Jinkela_wire_11690),
        .dout(new_Jinkela_wire_11691)
    );

    bfr new_Jinkela_buffer_9662 (
        .din(new_Jinkela_wire_11761),
        .dout(new_Jinkela_wire_11762)
    );

    bfr new_Jinkela_buffer_9598 (
        .din(new_Jinkela_wire_11691),
        .dout(new_Jinkela_wire_11692)
    );

    bfr new_Jinkela_buffer_9742 (
        .din(new_Jinkela_wire_11851),
        .dout(new_Jinkela_wire_11852)
    );

    bfr new_Jinkela_buffer_9599 (
        .din(new_Jinkela_wire_11692),
        .dout(new_Jinkela_wire_11693)
    );

    bfr new_Jinkela_buffer_9663 (
        .din(new_Jinkela_wire_11762),
        .dout(new_Jinkela_wire_11763)
    );

    bfr new_Jinkela_buffer_9600 (
        .din(new_Jinkela_wire_11693),
        .dout(new_Jinkela_wire_11694)
    );

    spl2 new_Jinkela_splitter_912 (
        .a(_0417_),
        .b(new_Jinkela_wire_12054),
        .c(new_Jinkela_wire_12055)
    );

    bfr new_Jinkela_buffer_9601 (
        .din(new_Jinkela_wire_11694),
        .dout(new_Jinkela_wire_11695)
    );

    bfr new_Jinkela_buffer_9664 (
        .din(new_Jinkela_wire_11763),
        .dout(new_Jinkela_wire_11764)
    );

    bfr new_Jinkela_buffer_9602 (
        .din(new_Jinkela_wire_11695),
        .dout(new_Jinkela_wire_11696)
    );

    bfr new_Jinkela_buffer_9743 (
        .din(new_Jinkela_wire_11852),
        .dout(new_Jinkela_wire_11853)
    );

    bfr new_Jinkela_buffer_9603 (
        .din(new_Jinkela_wire_11696),
        .dout(new_Jinkela_wire_11697)
    );

    bfr new_Jinkela_buffer_9665 (
        .din(new_Jinkela_wire_11764),
        .dout(new_Jinkela_wire_11765)
    );

    bfr new_Jinkela_buffer_9604 (
        .din(new_Jinkela_wire_11697),
        .dout(new_Jinkela_wire_11698)
    );

    bfr new_Jinkela_buffer_9847 (
        .din(new_Jinkela_wire_11966),
        .dout(new_Jinkela_wire_11967)
    );

    bfr new_Jinkela_buffer_9605 (
        .din(new_Jinkela_wire_11698),
        .dout(new_Jinkela_wire_11699)
    );

    bfr new_Jinkela_buffer_9666 (
        .din(new_Jinkela_wire_11765),
        .dout(new_Jinkela_wire_11766)
    );

    bfr new_Jinkela_buffer_9606 (
        .din(new_Jinkela_wire_11699),
        .dout(new_Jinkela_wire_11700)
    );

    bfr new_Jinkela_buffer_9744 (
        .din(new_Jinkela_wire_11853),
        .dout(new_Jinkela_wire_11854)
    );

    bfr new_Jinkela_buffer_9607 (
        .din(new_Jinkela_wire_11700),
        .dout(new_Jinkela_wire_11701)
    );

    bfr new_Jinkela_buffer_9667 (
        .din(new_Jinkela_wire_11766),
        .dout(new_Jinkela_wire_11767)
    );

    bfr new_Jinkela_buffer_2784 (
        .din(new_Jinkela_wire_3833),
        .dout(new_Jinkela_wire_3834)
    );

    bfr new_Jinkela_buffer_2710 (
        .din(new_Jinkela_wire_3753),
        .dout(new_Jinkela_wire_3754)
    );

    bfr new_Jinkela_buffer_2888 (
        .din(new_Jinkela_wire_3953),
        .dout(new_Jinkela_wire_3954)
    );

    bfr new_Jinkela_buffer_2711 (
        .din(new_Jinkela_wire_3754),
        .dout(new_Jinkela_wire_3755)
    );

    bfr new_Jinkela_buffer_2785 (
        .din(new_Jinkela_wire_3834),
        .dout(new_Jinkela_wire_3835)
    );

    bfr new_Jinkela_buffer_2712 (
        .din(new_Jinkela_wire_3755),
        .dout(new_Jinkela_wire_3756)
    );

    bfr new_Jinkela_buffer_2834 (
        .din(new_Jinkela_wire_3895),
        .dout(new_Jinkela_wire_3896)
    );

    bfr new_Jinkela_buffer_2713 (
        .din(new_Jinkela_wire_3756),
        .dout(new_Jinkela_wire_3757)
    );

    bfr new_Jinkela_buffer_2786 (
        .din(new_Jinkela_wire_3835),
        .dout(new_Jinkela_wire_3836)
    );

    bfr new_Jinkela_buffer_2714 (
        .din(new_Jinkela_wire_3757),
        .dout(new_Jinkela_wire_3758)
    );

    bfr new_Jinkela_buffer_2893 (
        .din(_1421_),
        .dout(new_Jinkela_wire_3963)
    );

    bfr new_Jinkela_buffer_2715 (
        .din(new_Jinkela_wire_3758),
        .dout(new_Jinkela_wire_3759)
    );

    bfr new_Jinkela_buffer_2787 (
        .din(new_Jinkela_wire_3836),
        .dout(new_Jinkela_wire_3837)
    );

    bfr new_Jinkela_buffer_2716 (
        .din(new_Jinkela_wire_3759),
        .dout(new_Jinkela_wire_3760)
    );

    bfr new_Jinkela_buffer_2835 (
        .din(new_Jinkela_wire_3896),
        .dout(new_Jinkela_wire_3897)
    );

    bfr new_Jinkela_buffer_2717 (
        .din(new_Jinkela_wire_3760),
        .dout(new_Jinkela_wire_3761)
    );

    bfr new_Jinkela_buffer_2788 (
        .din(new_Jinkela_wire_3837),
        .dout(new_Jinkela_wire_3838)
    );

    bfr new_Jinkela_buffer_2718 (
        .din(new_Jinkela_wire_3761),
        .dout(new_Jinkela_wire_3762)
    );

    bfr new_Jinkela_buffer_2719 (
        .din(new_Jinkela_wire_3762),
        .dout(new_Jinkela_wire_3763)
    );

    bfr new_Jinkela_buffer_2789 (
        .din(new_Jinkela_wire_3838),
        .dout(new_Jinkela_wire_3839)
    );

    bfr new_Jinkela_buffer_2720 (
        .din(new_Jinkela_wire_3763),
        .dout(new_Jinkela_wire_3764)
    );

    bfr new_Jinkela_buffer_2836 (
        .din(new_Jinkela_wire_3897),
        .dout(new_Jinkela_wire_3898)
    );

    bfr new_Jinkela_buffer_2721 (
        .din(new_Jinkela_wire_3764),
        .dout(new_Jinkela_wire_3765)
    );

    bfr new_Jinkela_buffer_2790 (
        .din(new_Jinkela_wire_3839),
        .dout(new_Jinkela_wire_3840)
    );

    bfr new_Jinkela_buffer_2722 (
        .din(new_Jinkela_wire_3765),
        .dout(new_Jinkela_wire_3766)
    );

    bfr new_Jinkela_buffer_2889 (
        .din(new_Jinkela_wire_3954),
        .dout(new_Jinkela_wire_3955)
    );

    bfr new_Jinkela_buffer_2723 (
        .din(new_Jinkela_wire_3766),
        .dout(new_Jinkela_wire_3767)
    );

    bfr new_Jinkela_buffer_2791 (
        .din(new_Jinkela_wire_3840),
        .dout(new_Jinkela_wire_3841)
    );

    bfr new_Jinkela_buffer_2724 (
        .din(new_Jinkela_wire_3767),
        .dout(new_Jinkela_wire_3768)
    );

    bfr new_Jinkela_buffer_2837 (
        .din(new_Jinkela_wire_3898),
        .dout(new_Jinkela_wire_3899)
    );

    bfr new_Jinkela_buffer_2725 (
        .din(new_Jinkela_wire_3768),
        .dout(new_Jinkela_wire_3769)
    );

    bfr new_Jinkela_buffer_2792 (
        .din(new_Jinkela_wire_3841),
        .dout(new_Jinkela_wire_3842)
    );

    bfr new_Jinkela_buffer_2726 (
        .din(new_Jinkela_wire_3769),
        .dout(new_Jinkela_wire_3770)
    );

    bfr new_Jinkela_buffer_2892 (
        .din(new_Jinkela_wire_3959),
        .dout(new_Jinkela_wire_3960)
    );

    spl2 new_Jinkela_splitter_384 (
        .a(_0900_),
        .b(new_Jinkela_wire_3964),
        .c(new_Jinkela_wire_3965)
    );

    bfr new_Jinkela_buffer_2727 (
        .din(new_Jinkela_wire_3770),
        .dout(new_Jinkela_wire_3771)
    );

    bfr new_Jinkela_buffer_2793 (
        .din(new_Jinkela_wire_3842),
        .dout(new_Jinkela_wire_3843)
    );

    bfr new_Jinkela_buffer_2728 (
        .din(new_Jinkela_wire_3771),
        .dout(new_Jinkela_wire_3772)
    );

    bfr new_Jinkela_buffer_2838 (
        .din(new_Jinkela_wire_3899),
        .dout(new_Jinkela_wire_3900)
    );

    bfr new_Jinkela_buffer_2729 (
        .din(new_Jinkela_wire_3772),
        .dout(new_Jinkela_wire_3773)
    );

    bfr new_Jinkela_buffer_2794 (
        .din(new_Jinkela_wire_3843),
        .dout(new_Jinkela_wire_3844)
    );

    bfr new_Jinkela_buffer_2730 (
        .din(new_Jinkela_wire_3773),
        .dout(new_Jinkela_wire_3774)
    );

    bfr new_Jinkela_buffer_13095 (
        .din(new_Jinkela_wire_15628),
        .dout(new_Jinkela_wire_15629)
    );

    spl2 new_Jinkela_splitter_1142 (
        .a(_1824_),
        .b(new_Jinkela_wire_15773),
        .c(new_Jinkela_wire_15774)
    );

    bfr new_Jinkela_buffer_13096 (
        .din(new_Jinkela_wire_15629),
        .dout(new_Jinkela_wire_15630)
    );

    bfr new_Jinkela_buffer_13162 (
        .din(new_Jinkela_wire_15723),
        .dout(new_Jinkela_wire_15724)
    );

    bfr new_Jinkela_buffer_13097 (
        .din(new_Jinkela_wire_15630),
        .dout(new_Jinkela_wire_15631)
    );

    bfr new_Jinkela_buffer_13180 (
        .din(new_Jinkela_wire_15761),
        .dout(new_Jinkela_wire_15762)
    );

    bfr new_Jinkela_buffer_13098 (
        .din(new_Jinkela_wire_15631),
        .dout(new_Jinkela_wire_15632)
    );

    bfr new_Jinkela_buffer_13163 (
        .din(new_Jinkela_wire_15724),
        .dout(new_Jinkela_wire_15725)
    );

    bfr new_Jinkela_buffer_13099 (
        .din(new_Jinkela_wire_15632),
        .dout(new_Jinkela_wire_15633)
    );

    bfr new_Jinkela_buffer_13100 (
        .din(new_Jinkela_wire_15633),
        .dout(new_Jinkela_wire_15634)
    );

    bfr new_Jinkela_buffer_13164 (
        .din(new_Jinkela_wire_15725),
        .dout(new_Jinkela_wire_15726)
    );

    bfr new_Jinkela_buffer_13101 (
        .din(new_Jinkela_wire_15634),
        .dout(new_Jinkela_wire_15635)
    );

    bfr new_Jinkela_buffer_13181 (
        .din(new_Jinkela_wire_15762),
        .dout(new_Jinkela_wire_15763)
    );

    bfr new_Jinkela_buffer_13102 (
        .din(new_Jinkela_wire_15635),
        .dout(new_Jinkela_wire_15636)
    );

    spl2 new_Jinkela_splitter_1130 (
        .a(new_Jinkela_wire_15726),
        .b(new_Jinkela_wire_15727),
        .c(new_Jinkela_wire_15728)
    );

    bfr new_Jinkela_buffer_13103 (
        .din(new_Jinkela_wire_15636),
        .dout(new_Jinkela_wire_15637)
    );

    bfr new_Jinkela_buffer_13182 (
        .din(new_Jinkela_wire_15763),
        .dout(new_Jinkela_wire_15764)
    );

    bfr new_Jinkela_buffer_13104 (
        .din(new_Jinkela_wire_15637),
        .dout(new_Jinkela_wire_15638)
    );

    spl2 new_Jinkela_splitter_1143 (
        .a(_1521_),
        .b(new_Jinkela_wire_15775),
        .c(new_Jinkela_wire_15776)
    );

    bfr new_Jinkela_buffer_13105 (
        .din(new_Jinkela_wire_15638),
        .dout(new_Jinkela_wire_15639)
    );

    spl2 new_Jinkela_splitter_1144 (
        .a(_0742_),
        .b(new_Jinkela_wire_15777),
        .c(new_Jinkela_wire_15778)
    );

    bfr new_Jinkela_buffer_13106 (
        .din(new_Jinkela_wire_15639),
        .dout(new_Jinkela_wire_15640)
    );

    bfr new_Jinkela_buffer_13183 (
        .din(new_Jinkela_wire_15764),
        .dout(new_Jinkela_wire_15765)
    );

    bfr new_Jinkela_buffer_13107 (
        .din(new_Jinkela_wire_15640),
        .dout(new_Jinkela_wire_15641)
    );

    spl2 new_Jinkela_splitter_1145 (
        .a(_1316_),
        .b(new_Jinkela_wire_15779),
        .c(new_Jinkela_wire_15780)
    );

    bfr new_Jinkela_buffer_13108 (
        .din(new_Jinkela_wire_15641),
        .dout(new_Jinkela_wire_15642)
    );

    bfr new_Jinkela_buffer_13184 (
        .din(new_Jinkela_wire_15765),
        .dout(new_Jinkela_wire_15766)
    );

    bfr new_Jinkela_buffer_13109 (
        .din(new_Jinkela_wire_15642),
        .dout(new_Jinkela_wire_15643)
    );

    spl2 new_Jinkela_splitter_1146 (
        .a(_0395_),
        .b(new_Jinkela_wire_15781),
        .c(new_Jinkela_wire_15782)
    );

    bfr new_Jinkela_buffer_13110 (
        .din(new_Jinkela_wire_15643),
        .dout(new_Jinkela_wire_15644)
    );

    bfr new_Jinkela_buffer_13185 (
        .din(new_Jinkela_wire_15766),
        .dout(new_Jinkela_wire_15767)
    );

    bfr new_Jinkela_buffer_13111 (
        .din(new_Jinkela_wire_15644),
        .dout(new_Jinkela_wire_15645)
    );

    bfr new_Jinkela_buffer_13238 (
        .din(_1185_),
        .dout(new_Jinkela_wire_15836)
    );

    bfr new_Jinkela_buffer_13187 (
        .din(_0999_),
        .dout(new_Jinkela_wire_15783)
    );

    bfr new_Jinkela_buffer_13112 (
        .din(new_Jinkela_wire_15645),
        .dout(new_Jinkela_wire_15646)
    );

    bfr new_Jinkela_buffer_13186 (
        .din(new_Jinkela_wire_15767),
        .dout(new_Jinkela_wire_15768)
    );

    bfr new_Jinkela_buffer_13113 (
        .din(new_Jinkela_wire_15646),
        .dout(new_Jinkela_wire_15647)
    );

    bfr new_Jinkela_buffer_13237 (
        .din(_0904_),
        .dout(new_Jinkela_wire_15835)
    );

    bfr new_Jinkela_buffer_13114 (
        .din(new_Jinkela_wire_15647),
        .dout(new_Jinkela_wire_15648)
    );

    spl2 new_Jinkela_splitter_1140 (
        .a(new_Jinkela_wire_15768),
        .b(new_Jinkela_wire_15769),
        .c(new_Jinkela_wire_15770)
    );

    bfr new_Jinkela_buffer_13115 (
        .din(new_Jinkela_wire_15648),
        .dout(new_Jinkela_wire_15649)
    );

    bfr new_Jinkela_buffer_13188 (
        .din(new_Jinkela_wire_15783),
        .dout(new_Jinkela_wire_15784)
    );

    and_ii _3550_ (
        .a(new_Jinkela_wire_18583),
        .b(new_Jinkela_wire_13398),
        .c(_0847_)
    );

    and_bb _3551_ (
        .a(new_Jinkela_wire_18584),
        .b(new_Jinkela_wire_13399),
        .c(_0848_)
    );

    or_bb _3552_ (
        .a(new_Jinkela_wire_2342),
        .b(new_Jinkela_wire_19468),
        .c(_0849_)
    );

    and_ii _3553_ (
        .a(new_Jinkela_wire_15026),
        .b(new_Jinkela_wire_3359),
        .c(_0851_)
    );

    and_bb _3554_ (
        .a(new_Jinkela_wire_15027),
        .b(new_Jinkela_wire_3360),
        .c(_0852_)
    );

    or_bb _3555_ (
        .a(new_Jinkela_wire_2015),
        .b(new_Jinkela_wire_19185),
        .c(_0853_)
    );

    and_ii _3556_ (
        .a(new_Jinkela_wire_8299),
        .b(new_Jinkela_wire_1575),
        .c(_0854_)
    );

    and_bb _3557_ (
        .a(new_Jinkela_wire_8300),
        .b(new_Jinkela_wire_1576),
        .c(_0855_)
    );

    or_bb _3558_ (
        .a(new_Jinkela_wire_13677),
        .b(new_Jinkela_wire_14184),
        .c(_0856_)
    );

    and_ii _3559_ (
        .a(new_Jinkela_wire_20367),
        .b(new_Jinkela_wire_21090),
        .c(_0857_)
    );

    and_bb _3560_ (
        .a(new_Jinkela_wire_20368),
        .b(new_Jinkela_wire_21091),
        .c(_0858_)
    );

    or_bb _3561_ (
        .a(new_Jinkela_wire_5050),
        .b(new_Jinkela_wire_6806),
        .c(_0859_)
    );

    and_ii _3562_ (
        .a(new_Jinkela_wire_13390),
        .b(new_Jinkela_wire_16868),
        .c(_0860_)
    );

    and_bb _3563_ (
        .a(new_Jinkela_wire_13391),
        .b(new_Jinkela_wire_16869),
        .c(_0862_)
    );

    or_bb _3564_ (
        .a(new_Jinkela_wire_18804),
        .b(new_Jinkela_wire_16194),
        .c(_0863_)
    );

    and_ii _3565_ (
        .a(new_Jinkela_wire_852),
        .b(new_Jinkela_wire_18940),
        .c(_0864_)
    );

    and_bb _3566_ (
        .a(new_Jinkela_wire_853),
        .b(new_Jinkela_wire_18941),
        .c(_0865_)
    );

    or_bb _3567_ (
        .a(new_Jinkela_wire_4708),
        .b(new_Jinkela_wire_17551),
        .c(_0866_)
    );

    and_ii _3568_ (
        .a(new_Jinkela_wire_10102),
        .b(new_Jinkela_wire_2958),
        .c(_0867_)
    );

    and_bb _3569_ (
        .a(new_Jinkela_wire_10103),
        .b(new_Jinkela_wire_2959),
        .c(_0868_)
    );

    or_bb _3570_ (
        .a(new_Jinkela_wire_15746),
        .b(new_Jinkela_wire_13047),
        .c(_0869_)
    );

    and_ii _3571_ (
        .a(new_Jinkela_wire_13312),
        .b(new_Jinkela_wire_10392),
        .c(_0870_)
    );

    and_bb _3572_ (
        .a(new_Jinkela_wire_13313),
        .b(new_Jinkela_wire_10393),
        .c(_0871_)
    );

    or_bb _3573_ (
        .a(new_Jinkela_wire_4828),
        .b(new_Jinkela_wire_19112),
        .c(_0873_)
    );

    and_ii _3574_ (
        .a(new_Jinkela_wire_4715),
        .b(new_Jinkela_wire_7502),
        .c(_0874_)
    );

    and_bb _3575_ (
        .a(new_Jinkela_wire_4716),
        .b(new_Jinkela_wire_7503),
        .c(_0875_)
    );

    and_ii _3576_ (
        .a(new_Jinkela_wire_2484),
        .b(new_Jinkela_wire_5054),
        .c(_0876_)
    );

    and_bb _3577_ (
        .a(new_Jinkela_wire_7174),
        .b(new_Jinkela_wire_3819),
        .c(_0877_)
    );

    and_ii _3578_ (
        .a(new_Jinkela_wire_7175),
        .b(new_Jinkela_wire_3820),
        .c(_0878_)
    );

    or_bb _3579_ (
        .a(new_Jinkela_wire_4538),
        .b(new_Jinkela_wire_11397),
        .c(new_net_3964)
    );

    or_bb _3580_ (
        .a(new_Jinkela_wire_11398),
        .b(new_Jinkela_wire_5091),
        .c(_0879_)
    );

    and_ii _3581_ (
        .a(new_Jinkela_wire_19113),
        .b(new_Jinkela_wire_13052),
        .c(_0880_)
    );

    and_bb _3582_ (
        .a(new_Jinkela_wire_379),
        .b(new_Jinkela_wire_674),
        .c(_0881_)
    );

    and_ii _3583_ (
        .a(new_Jinkela_wire_17552),
        .b(new_Jinkela_wire_16199),
        .c(_0883_)
    );

    and_bb _3584_ (
        .a(new_Jinkela_wire_407),
        .b(new_Jinkela_wire_513),
        .c(_0884_)
    );

    and_ii _3585_ (
        .a(new_Jinkela_wire_6807),
        .b(new_Jinkela_wire_14189),
        .c(_0885_)
    );

    and_bb _3586_ (
        .a(new_Jinkela_wire_173),
        .b(new_Jinkela_wire_142),
        .c(_0886_)
    );

    and_ii _3587_ (
        .a(new_Jinkela_wire_19186),
        .b(new_Jinkela_wire_19473),
        .c(_0887_)
    );

    and_bb _3588_ (
        .a(new_Jinkela_wire_614),
        .b(new_Jinkela_wire_211),
        .c(_0888_)
    );

    and_bb _3589_ (
        .a(new_Jinkela_wire_419),
        .b(new_Jinkela_wire_586),
        .c(_0889_)
    );

    and_ii _3590_ (
        .a(new_Jinkela_wire_7749),
        .b(new_Jinkela_wire_1613),
        .c(_0890_)
    );

    and_ii _3591_ (
        .a(new_Jinkela_wire_6521),
        .b(new_Jinkela_wire_17634),
        .c(_0891_)
    );

    bfr new_Jinkela_buffer_2890 (
        .din(new_Jinkela_wire_3955),
        .dout(new_Jinkela_wire_3956)
    );

    bfr new_Jinkela_buffer_6193 (
        .din(new_Jinkela_wire_7862),
        .dout(new_Jinkela_wire_7863)
    );

    bfr new_Jinkela_buffer_16566 (
        .din(new_Jinkela_wire_19764),
        .dout(new_Jinkela_wire_19765)
    );

    bfr new_Jinkela_buffer_16480 (
        .din(new_Jinkela_wire_19668),
        .dout(new_Jinkela_wire_19669)
    );

    bfr new_Jinkela_buffer_2731 (
        .din(new_Jinkela_wire_3774),
        .dout(new_Jinkela_wire_3775)
    );

    bfr new_Jinkela_buffer_6133 (
        .din(new_Jinkela_wire_7790),
        .dout(new_Jinkela_wire_7791)
    );

    bfr new_Jinkela_buffer_2795 (
        .din(new_Jinkela_wire_3844),
        .dout(new_Jinkela_wire_3845)
    );

    bfr new_Jinkela_buffer_6297 (
        .din(new_Jinkela_wire_7974),
        .dout(new_Jinkela_wire_7975)
    );

    bfr new_Jinkela_buffer_16700 (
        .din(new_Jinkela_wire_19914),
        .dout(new_Jinkela_wire_19915)
    );

    bfr new_Jinkela_buffer_16481 (
        .din(new_Jinkela_wire_19669),
        .dout(new_Jinkela_wire_19670)
    );

    bfr new_Jinkela_buffer_2732 (
        .din(new_Jinkela_wire_3775),
        .dout(new_Jinkela_wire_3776)
    );

    bfr new_Jinkela_buffer_6134 (
        .din(new_Jinkela_wire_7791),
        .dout(new_Jinkela_wire_7792)
    );

    bfr new_Jinkela_buffer_2839 (
        .din(new_Jinkela_wire_3900),
        .dout(new_Jinkela_wire_3901)
    );

    bfr new_Jinkela_buffer_6194 (
        .din(new_Jinkela_wire_7863),
        .dout(new_Jinkela_wire_7864)
    );

    bfr new_Jinkela_buffer_16567 (
        .din(new_Jinkela_wire_19765),
        .dout(new_Jinkela_wire_19766)
    );

    bfr new_Jinkela_buffer_16482 (
        .din(new_Jinkela_wire_19670),
        .dout(new_Jinkela_wire_19671)
    );

    bfr new_Jinkela_buffer_2733 (
        .din(new_Jinkela_wire_3776),
        .dout(new_Jinkela_wire_3777)
    );

    bfr new_Jinkela_buffer_6135 (
        .din(new_Jinkela_wire_7792),
        .dout(new_Jinkela_wire_7793)
    );

    bfr new_Jinkela_buffer_2796 (
        .din(new_Jinkela_wire_3845),
        .dout(new_Jinkela_wire_3846)
    );

    bfr new_Jinkela_buffer_6205 (
        .din(new_Jinkela_wire_7878),
        .dout(new_Jinkela_wire_7879)
    );

    bfr new_Jinkela_buffer_16594 (
        .din(new_Jinkela_wire_19802),
        .dout(new_Jinkela_wire_19803)
    );

    bfr new_Jinkela_buffer_16483 (
        .din(new_Jinkela_wire_19671),
        .dout(new_Jinkela_wire_19672)
    );

    bfr new_Jinkela_buffer_2734 (
        .din(new_Jinkela_wire_3777),
        .dout(new_Jinkela_wire_3778)
    );

    bfr new_Jinkela_buffer_6136 (
        .din(new_Jinkela_wire_7793),
        .dout(new_Jinkela_wire_7794)
    );

    bfr new_Jinkela_buffer_2894 (
        .din(_1804_),
        .dout(new_Jinkela_wire_3966)
    );

    bfr new_Jinkela_buffer_6195 (
        .din(new_Jinkela_wire_7864),
        .dout(new_Jinkela_wire_7865)
    );

    bfr new_Jinkela_buffer_16568 (
        .din(new_Jinkela_wire_19766),
        .dout(new_Jinkela_wire_19767)
    );

    bfr new_Jinkela_buffer_16484 (
        .din(new_Jinkela_wire_19672),
        .dout(new_Jinkela_wire_19673)
    );

    bfr new_Jinkela_buffer_2735 (
        .din(new_Jinkela_wire_3778),
        .dout(new_Jinkela_wire_3779)
    );

    bfr new_Jinkela_buffer_6137 (
        .din(new_Jinkela_wire_7794),
        .dout(new_Jinkela_wire_7795)
    );

    bfr new_Jinkela_buffer_2797 (
        .din(new_Jinkela_wire_3846),
        .dout(new_Jinkela_wire_3847)
    );

    bfr new_Jinkela_buffer_16704 (
        .din(new_Jinkela_wire_19920),
        .dout(new_Jinkela_wire_19921)
    );

    spl2 new_Jinkela_splitter_688 (
        .a(_1785_),
        .b(new_Jinkela_wire_7980),
        .c(new_Jinkela_wire_7981)
    );

    bfr new_Jinkela_buffer_16485 (
        .din(new_Jinkela_wire_19673),
        .dout(new_Jinkela_wire_19674)
    );

    bfr new_Jinkela_buffer_2736 (
        .din(new_Jinkela_wire_3779),
        .dout(new_Jinkela_wire_3780)
    );

    bfr new_Jinkela_buffer_6138 (
        .din(new_Jinkela_wire_7795),
        .dout(new_Jinkela_wire_7796)
    );

    bfr new_Jinkela_buffer_2840 (
        .din(new_Jinkela_wire_3901),
        .dout(new_Jinkela_wire_3902)
    );

    spl2 new_Jinkela_splitter_684 (
        .a(new_Jinkela_wire_7865),
        .b(new_Jinkela_wire_7866),
        .c(new_Jinkela_wire_7867)
    );

    bfr new_Jinkela_buffer_16569 (
        .din(new_Jinkela_wire_19767),
        .dout(new_Jinkela_wire_19768)
    );

    bfr new_Jinkela_buffer_16486 (
        .din(new_Jinkela_wire_19674),
        .dout(new_Jinkela_wire_19675)
    );

    bfr new_Jinkela_buffer_2737 (
        .din(new_Jinkela_wire_3780),
        .dout(new_Jinkela_wire_3781)
    );

    bfr new_Jinkela_buffer_6139 (
        .din(new_Jinkela_wire_7796),
        .dout(new_Jinkela_wire_7797)
    );

    bfr new_Jinkela_buffer_2798 (
        .din(new_Jinkela_wire_3847),
        .dout(new_Jinkela_wire_3848)
    );

    bfr new_Jinkela_buffer_6302 (
        .din(_0415_),
        .dout(new_Jinkela_wire_7982)
    );

    bfr new_Jinkela_buffer_16595 (
        .din(new_Jinkela_wire_19803),
        .dout(new_Jinkela_wire_19804)
    );

    bfr new_Jinkela_buffer_6336 (
        .din(_1055_),
        .dout(new_Jinkela_wire_8018)
    );

    bfr new_Jinkela_buffer_16487 (
        .din(new_Jinkela_wire_19675),
        .dout(new_Jinkela_wire_19676)
    );

    bfr new_Jinkela_buffer_2738 (
        .din(new_Jinkela_wire_3781),
        .dout(new_Jinkela_wire_3782)
    );

    bfr new_Jinkela_buffer_6140 (
        .din(new_Jinkela_wire_7797),
        .dout(new_Jinkela_wire_7798)
    );

    bfr new_Jinkela_buffer_2891 (
        .din(new_Jinkela_wire_3956),
        .dout(new_Jinkela_wire_3957)
    );

    bfr new_Jinkela_buffer_6206 (
        .din(new_Jinkela_wire_7879),
        .dout(new_Jinkela_wire_7880)
    );

    bfr new_Jinkela_buffer_16570 (
        .din(new_Jinkela_wire_19768),
        .dout(new_Jinkela_wire_19769)
    );

    bfr new_Jinkela_buffer_16488 (
        .din(new_Jinkela_wire_19676),
        .dout(new_Jinkela_wire_19677)
    );

    bfr new_Jinkela_buffer_2739 (
        .din(new_Jinkela_wire_3782),
        .dout(new_Jinkela_wire_3783)
    );

    bfr new_Jinkela_buffer_6141 (
        .din(new_Jinkela_wire_7798),
        .dout(new_Jinkela_wire_7799)
    );

    bfr new_Jinkela_buffer_2799 (
        .din(new_Jinkela_wire_3848),
        .dout(new_Jinkela_wire_3849)
    );

    bfr new_Jinkela_buffer_6207 (
        .din(new_Jinkela_wire_7880),
        .dout(new_Jinkela_wire_7881)
    );

    bfr new_Jinkela_buffer_16701 (
        .din(new_Jinkela_wire_19915),
        .dout(new_Jinkela_wire_19916)
    );

    bfr new_Jinkela_buffer_16489 (
        .din(new_Jinkela_wire_19677),
        .dout(new_Jinkela_wire_19678)
    );

    bfr new_Jinkela_buffer_2740 (
        .din(new_Jinkela_wire_3783),
        .dout(new_Jinkela_wire_3784)
    );

    bfr new_Jinkela_buffer_6142 (
        .din(new_Jinkela_wire_7799),
        .dout(new_Jinkela_wire_7800)
    );

    bfr new_Jinkela_buffer_2841 (
        .din(new_Jinkela_wire_3902),
        .dout(new_Jinkela_wire_3903)
    );

    bfr new_Jinkela_buffer_6298 (
        .din(new_Jinkela_wire_7975),
        .dout(new_Jinkela_wire_7976)
    );

    bfr new_Jinkela_buffer_16571 (
        .din(new_Jinkela_wire_19769),
        .dout(new_Jinkela_wire_19770)
    );

    bfr new_Jinkela_buffer_16490 (
        .din(new_Jinkela_wire_19678),
        .dout(new_Jinkela_wire_19679)
    );

    bfr new_Jinkela_buffer_2741 (
        .din(new_Jinkela_wire_3784),
        .dout(new_Jinkela_wire_3785)
    );

    bfr new_Jinkela_buffer_6143 (
        .din(new_Jinkela_wire_7800),
        .dout(new_Jinkela_wire_7801)
    );

    bfr new_Jinkela_buffer_2800 (
        .din(new_Jinkela_wire_3849),
        .dout(new_Jinkela_wire_3850)
    );

    bfr new_Jinkela_buffer_6208 (
        .din(new_Jinkela_wire_7881),
        .dout(new_Jinkela_wire_7882)
    );

    bfr new_Jinkela_buffer_16596 (
        .din(new_Jinkela_wire_19804),
        .dout(new_Jinkela_wire_19805)
    );

    bfr new_Jinkela_buffer_16491 (
        .din(new_Jinkela_wire_19679),
        .dout(new_Jinkela_wire_19680)
    );

    bfr new_Jinkela_buffer_2742 (
        .din(new_Jinkela_wire_3785),
        .dout(new_Jinkela_wire_3786)
    );

    bfr new_Jinkela_buffer_6144 (
        .din(new_Jinkela_wire_7801),
        .dout(new_Jinkela_wire_7802)
    );

    spl2 new_Jinkela_splitter_387 (
        .a(_1516_),
        .b(new_Jinkela_wire_4074),
        .c(new_Jinkela_wire_4075)
    );

    bfr new_Jinkela_buffer_16572 (
        .din(new_Jinkela_wire_19770),
        .dout(new_Jinkela_wire_19771)
    );

    spl2 new_Jinkela_splitter_383 (
        .a(new_Jinkela_wire_3960),
        .b(new_Jinkela_wire_3961),
        .c(new_Jinkela_wire_3962)
    );

    bfr new_Jinkela_buffer_16492 (
        .din(new_Jinkela_wire_19680),
        .dout(new_Jinkela_wire_19681)
    );

    bfr new_Jinkela_buffer_2743 (
        .din(new_Jinkela_wire_3786),
        .dout(new_Jinkela_wire_3787)
    );

    bfr new_Jinkela_buffer_6145 (
        .din(new_Jinkela_wire_7802),
        .dout(new_Jinkela_wire_7803)
    );

    bfr new_Jinkela_buffer_2801 (
        .din(new_Jinkela_wire_3850),
        .dout(new_Jinkela_wire_3851)
    );

    bfr new_Jinkela_buffer_6209 (
        .din(new_Jinkela_wire_7882),
        .dout(new_Jinkela_wire_7883)
    );

    bfr new_Jinkela_buffer_16493 (
        .din(new_Jinkela_wire_19681),
        .dout(new_Jinkela_wire_19682)
    );

    bfr new_Jinkela_buffer_2744 (
        .din(new_Jinkela_wire_3787),
        .dout(new_Jinkela_wire_3788)
    );

    bfr new_Jinkela_buffer_6146 (
        .din(new_Jinkela_wire_7803),
        .dout(new_Jinkela_wire_7804)
    );

    spl2 new_Jinkela_splitter_1459 (
        .a(_1295_),
        .b(new_Jinkela_wire_19930),
        .c(new_Jinkela_wire_19931)
    );

    bfr new_Jinkela_buffer_2842 (
        .din(new_Jinkela_wire_3903),
        .dout(new_Jinkela_wire_3904)
    );

    bfr new_Jinkela_buffer_6299 (
        .din(new_Jinkela_wire_7976),
        .dout(new_Jinkela_wire_7977)
    );

    bfr new_Jinkela_buffer_16573 (
        .din(new_Jinkela_wire_19771),
        .dout(new_Jinkela_wire_19772)
    );

    bfr new_Jinkela_buffer_16494 (
        .din(new_Jinkela_wire_19682),
        .dout(new_Jinkela_wire_19683)
    );

    bfr new_Jinkela_buffer_2745 (
        .din(new_Jinkela_wire_3788),
        .dout(new_Jinkela_wire_3789)
    );

    bfr new_Jinkela_buffer_6147 (
        .din(new_Jinkela_wire_7804),
        .dout(new_Jinkela_wire_7805)
    );

    bfr new_Jinkela_buffer_2802 (
        .din(new_Jinkela_wire_3851),
        .dout(new_Jinkela_wire_3852)
    );

    bfr new_Jinkela_buffer_6210 (
        .din(new_Jinkela_wire_7883),
        .dout(new_Jinkela_wire_7884)
    );

    bfr new_Jinkela_buffer_16597 (
        .din(new_Jinkela_wire_19805),
        .dout(new_Jinkela_wire_19806)
    );

    bfr new_Jinkela_buffer_16495 (
        .din(new_Jinkela_wire_19683),
        .dout(new_Jinkela_wire_19684)
    );

    bfr new_Jinkela_buffer_2746 (
        .din(new_Jinkela_wire_3789),
        .dout(new_Jinkela_wire_3790)
    );

    bfr new_Jinkela_buffer_6148 (
        .din(new_Jinkela_wire_7805),
        .dout(new_Jinkela_wire_7806)
    );

    bfr new_Jinkela_buffer_16574 (
        .din(new_Jinkela_wire_19772),
        .dout(new_Jinkela_wire_19773)
    );

    bfr new_Jinkela_buffer_6303 (
        .din(_1136_),
        .dout(new_Jinkela_wire_7983)
    );

    bfr new_Jinkela_buffer_2747 (
        .din(new_Jinkela_wire_3790),
        .dout(new_Jinkela_wire_3791)
    );

    bfr new_Jinkela_buffer_6149 (
        .din(new_Jinkela_wire_7806),
        .dout(new_Jinkela_wire_7807)
    );

    bfr new_Jinkela_buffer_2803 (
        .din(new_Jinkela_wire_3852),
        .dout(new_Jinkela_wire_3853)
    );

    bfr new_Jinkela_buffer_6211 (
        .din(new_Jinkela_wire_7884),
        .dout(new_Jinkela_wire_7885)
    );

    bfr new_Jinkela_buffer_16575 (
        .din(new_Jinkela_wire_19773),
        .dout(new_Jinkela_wire_19774)
    );

    bfr new_Jinkela_buffer_2748 (
        .din(new_Jinkela_wire_3791),
        .dout(new_Jinkela_wire_3792)
    );

    bfr new_Jinkela_buffer_6150 (
        .din(new_Jinkela_wire_7807),
        .dout(new_Jinkela_wire_7808)
    );

    bfr new_Jinkela_buffer_16598 (
        .din(new_Jinkela_wire_19806),
        .dout(new_Jinkela_wire_19807)
    );

    bfr new_Jinkela_buffer_2843 (
        .din(new_Jinkela_wire_3904),
        .dout(new_Jinkela_wire_3905)
    );

    bfr new_Jinkela_buffer_6300 (
        .din(new_Jinkela_wire_7977),
        .dout(new_Jinkela_wire_7978)
    );

    bfr new_Jinkela_buffer_16576 (
        .din(new_Jinkela_wire_19774),
        .dout(new_Jinkela_wire_19775)
    );

    bfr new_Jinkela_buffer_2749 (
        .din(new_Jinkela_wire_3792),
        .dout(new_Jinkela_wire_3793)
    );

    bfr new_Jinkela_buffer_6151 (
        .din(new_Jinkela_wire_7808),
        .dout(new_Jinkela_wire_7809)
    );

    bfr new_Jinkela_buffer_16705 (
        .din(new_Jinkela_wire_19921),
        .dout(new_Jinkela_wire_19922)
    );

    bfr new_Jinkela_buffer_2804 (
        .din(new_Jinkela_wire_3853),
        .dout(new_Jinkela_wire_3854)
    );

    bfr new_Jinkela_buffer_6212 (
        .din(new_Jinkela_wire_7885),
        .dout(new_Jinkela_wire_7886)
    );

    bfr new_Jinkela_buffer_16577 (
        .din(new_Jinkela_wire_19775),
        .dout(new_Jinkela_wire_19776)
    );

    bfr new_Jinkela_buffer_2750 (
        .din(new_Jinkela_wire_3793),
        .dout(new_Jinkela_wire_3794)
    );

    bfr new_Jinkela_buffer_6152 (
        .din(new_Jinkela_wire_7809),
        .dout(new_Jinkela_wire_7810)
    );

    bfr new_Jinkela_buffer_16599 (
        .din(new_Jinkela_wire_19807),
        .dout(new_Jinkela_wire_19808)
    );

    spl2 new_Jinkela_splitter_386 (
        .a(_1319_),
        .b(new_Jinkela_wire_4072),
        .c(new_Jinkela_wire_4073)
    );

    bfr new_Jinkela_buffer_16578 (
        .din(new_Jinkela_wire_19776),
        .dout(new_Jinkela_wire_19777)
    );

    spl2 new_Jinkela_splitter_690 (
        .a(_0305_),
        .b(new_Jinkela_wire_8019),
        .c(new_Jinkela_wire_8020)
    );

    bfr new_Jinkela_buffer_2751 (
        .din(new_Jinkela_wire_3794),
        .dout(new_Jinkela_wire_3795)
    );

    bfr new_Jinkela_buffer_6153 (
        .din(new_Jinkela_wire_7810),
        .dout(new_Jinkela_wire_7811)
    );

    bfr new_Jinkela_buffer_16708 (
        .din(new_Jinkela_wire_19926),
        .dout(new_Jinkela_wire_19927)
    );

    spl2 new_Jinkela_splitter_1460 (
        .a(_1041_),
        .b(new_Jinkela_wire_19932),
        .c(new_Jinkela_wire_19933)
    );

    bfr new_Jinkela_buffer_15741 (
        .din(new_Jinkela_wire_18753),
        .dout(new_Jinkela_wire_18754)
    );

    bfr new_Jinkela_buffer_15669 (
        .din(new_Jinkela_wire_18667),
        .dout(new_Jinkela_wire_18668)
    );

    bfr new_Jinkela_buffer_15766 (
        .din(new_Jinkela_wire_18788),
        .dout(new_Jinkela_wire_18789)
    );

    bfr new_Jinkela_buffer_15670 (
        .din(new_Jinkela_wire_18668),
        .dout(new_Jinkela_wire_18669)
    );

    bfr new_Jinkela_buffer_15742 (
        .din(new_Jinkela_wire_18754),
        .dout(new_Jinkela_wire_18755)
    );

    bfr new_Jinkela_buffer_15671 (
        .din(new_Jinkela_wire_18669),
        .dout(new_Jinkela_wire_18670)
    );

    bfr new_Jinkela_buffer_15757 (
        .din(new_Jinkela_wire_18775),
        .dout(new_Jinkela_wire_18776)
    );

    bfr new_Jinkela_buffer_15672 (
        .din(new_Jinkela_wire_18670),
        .dout(new_Jinkela_wire_18671)
    );

    bfr new_Jinkela_buffer_15743 (
        .din(new_Jinkela_wire_18755),
        .dout(new_Jinkela_wire_18756)
    );

    bfr new_Jinkela_buffer_15673 (
        .din(new_Jinkela_wire_18671),
        .dout(new_Jinkela_wire_18672)
    );

    bfr new_Jinkela_buffer_15777 (
        .din(_0862_),
        .dout(new_Jinkela_wire_18804)
    );

    bfr new_Jinkela_buffer_15674 (
        .din(new_Jinkela_wire_18672),
        .dout(new_Jinkela_wire_18673)
    );

    bfr new_Jinkela_buffer_15773 (
        .din(new_Jinkela_wire_18799),
        .dout(new_Jinkela_wire_18800)
    );

    bfr new_Jinkela_buffer_15744 (
        .din(new_Jinkela_wire_18756),
        .dout(new_Jinkela_wire_18757)
    );

    bfr new_Jinkela_buffer_15675 (
        .din(new_Jinkela_wire_18673),
        .dout(new_Jinkela_wire_18674)
    );

    bfr new_Jinkela_buffer_15758 (
        .din(new_Jinkela_wire_18776),
        .dout(new_Jinkela_wire_18777)
    );

    bfr new_Jinkela_buffer_15676 (
        .din(new_Jinkela_wire_18674),
        .dout(new_Jinkela_wire_18675)
    );

    spl2 new_Jinkela_splitter_1355 (
        .a(new_Jinkela_wire_18757),
        .b(new_Jinkela_wire_18758),
        .c(new_Jinkela_wire_18759)
    );

    bfr new_Jinkela_buffer_15677 (
        .din(new_Jinkela_wire_18675),
        .dout(new_Jinkela_wire_18676)
    );

    bfr new_Jinkela_buffer_15759 (
        .din(new_Jinkela_wire_18777),
        .dout(new_Jinkela_wire_18778)
    );

    bfr new_Jinkela_buffer_15678 (
        .din(new_Jinkela_wire_18676),
        .dout(new_Jinkela_wire_18677)
    );

    bfr new_Jinkela_buffer_15767 (
        .din(new_Jinkela_wire_18789),
        .dout(new_Jinkela_wire_18790)
    );

    bfr new_Jinkela_buffer_15679 (
        .din(new_Jinkela_wire_18677),
        .dout(new_Jinkela_wire_18678)
    );

    bfr new_Jinkela_buffer_15769 (
        .din(new_Jinkela_wire_18793),
        .dout(new_Jinkela_wire_18794)
    );

    bfr new_Jinkela_buffer_15680 (
        .din(new_Jinkela_wire_18678),
        .dout(new_Jinkela_wire_18679)
    );

    bfr new_Jinkela_buffer_15760 (
        .din(new_Jinkela_wire_18778),
        .dout(new_Jinkela_wire_18779)
    );

    bfr new_Jinkela_buffer_15681 (
        .din(new_Jinkela_wire_18679),
        .dout(new_Jinkela_wire_18680)
    );

    bfr new_Jinkela_buffer_15682 (
        .din(new_Jinkela_wire_18680),
        .dout(new_Jinkela_wire_18681)
    );

    bfr new_Jinkela_buffer_15761 (
        .din(new_Jinkela_wire_18779),
        .dout(new_Jinkela_wire_18780)
    );

    bfr new_Jinkela_buffer_15683 (
        .din(new_Jinkela_wire_18681),
        .dout(new_Jinkela_wire_18682)
    );

    bfr new_Jinkela_buffer_15770 (
        .din(new_Jinkela_wire_18794),
        .dout(new_Jinkela_wire_18795)
    );

    bfr new_Jinkela_buffer_15684 (
        .din(new_Jinkela_wire_18682),
        .dout(new_Jinkela_wire_18683)
    );

    bfr new_Jinkela_buffer_15762 (
        .din(new_Jinkela_wire_18780),
        .dout(new_Jinkela_wire_18781)
    );

    bfr new_Jinkela_buffer_15685 (
        .din(new_Jinkela_wire_18683),
        .dout(new_Jinkela_wire_18684)
    );

    spl2 new_Jinkela_splitter_1362 (
        .a(_0956_),
        .b(new_Jinkela_wire_18805),
        .c(new_Jinkela_wire_18806)
    );

    bfr new_Jinkela_buffer_15763 (
        .din(new_Jinkela_wire_18781),
        .dout(new_Jinkela_wire_18782)
    );

    bfr new_Jinkela_buffer_15771 (
        .din(new_Jinkela_wire_18795),
        .dout(new_Jinkela_wire_18796)
    );

    spl2 new_Jinkela_splitter_1358 (
        .a(new_Jinkela_wire_18782),
        .b(new_Jinkela_wire_18783),
        .c(new_Jinkela_wire_18784)
    );

    bfr new_Jinkela_buffer_15774 (
        .din(new_Jinkela_wire_18800),
        .dout(new_Jinkela_wire_18801)
    );

    bfr new_Jinkela_buffer_15778 (
        .din(_0429_),
        .dout(new_Jinkela_wire_18807)
    );

    bfr new_Jinkela_buffer_15779 (
        .din(_0600_),
        .dout(new_Jinkela_wire_18808)
    );

    bfr new_Jinkela_buffer_12230 (
        .din(new_Jinkela_wire_14727),
        .dout(new_Jinkela_wire_14728)
    );

    bfr new_Jinkela_buffer_12294 (
        .din(new_Jinkela_wire_14793),
        .dout(new_Jinkela_wire_14794)
    );

    bfr new_Jinkela_buffer_12231 (
        .din(new_Jinkela_wire_14728),
        .dout(new_Jinkela_wire_14729)
    );

    bfr new_Jinkela_buffer_12398 (
        .din(new_Jinkela_wire_14899),
        .dout(new_Jinkela_wire_14900)
    );

    bfr new_Jinkela_buffer_12232 (
        .din(new_Jinkela_wire_14729),
        .dout(new_Jinkela_wire_14730)
    );

    bfr new_Jinkela_buffer_12295 (
        .din(new_Jinkela_wire_14794),
        .dout(new_Jinkela_wire_14795)
    );

    bfr new_Jinkela_buffer_12233 (
        .din(new_Jinkela_wire_14730),
        .dout(new_Jinkela_wire_14731)
    );

    bfr new_Jinkela_buffer_12234 (
        .din(new_Jinkela_wire_14731),
        .dout(new_Jinkela_wire_14732)
    );

    bfr new_Jinkela_buffer_12296 (
        .din(new_Jinkela_wire_14795),
        .dout(new_Jinkela_wire_14796)
    );

    bfr new_Jinkela_buffer_12235 (
        .din(new_Jinkela_wire_14732),
        .dout(new_Jinkela_wire_14733)
    );

    bfr new_Jinkela_buffer_12399 (
        .din(new_Jinkela_wire_14900),
        .dout(new_Jinkela_wire_14901)
    );

    bfr new_Jinkela_buffer_12236 (
        .din(new_Jinkela_wire_14733),
        .dout(new_Jinkela_wire_14734)
    );

    bfr new_Jinkela_buffer_12297 (
        .din(new_Jinkela_wire_14796),
        .dout(new_Jinkela_wire_14797)
    );

    bfr new_Jinkela_buffer_12237 (
        .din(new_Jinkela_wire_14734),
        .dout(new_Jinkela_wire_14735)
    );

    bfr new_Jinkela_buffer_12491 (
        .din(new_Jinkela_wire_14994),
        .dout(new_Jinkela_wire_14995)
    );

    bfr new_Jinkela_buffer_12238 (
        .din(new_Jinkela_wire_14735),
        .dout(new_Jinkela_wire_14736)
    );

    bfr new_Jinkela_buffer_12298 (
        .din(new_Jinkela_wire_14797),
        .dout(new_Jinkela_wire_14798)
    );

    bfr new_Jinkela_buffer_12239 (
        .din(new_Jinkela_wire_14736),
        .dout(new_Jinkela_wire_14737)
    );

    bfr new_Jinkela_buffer_12400 (
        .din(new_Jinkela_wire_14901),
        .dout(new_Jinkela_wire_14902)
    );

    bfr new_Jinkela_buffer_12240 (
        .din(new_Jinkela_wire_14737),
        .dout(new_Jinkela_wire_14738)
    );

    bfr new_Jinkela_buffer_12299 (
        .din(new_Jinkela_wire_14798),
        .dout(new_Jinkela_wire_14799)
    );

    bfr new_Jinkela_buffer_12241 (
        .din(new_Jinkela_wire_14738),
        .dout(new_Jinkela_wire_14739)
    );

    spl2 new_Jinkela_splitter_1105 (
        .a(_0618_),
        .b(new_Jinkela_wire_15122),
        .c(new_Jinkela_wire_15123)
    );

    bfr new_Jinkela_buffer_12242 (
        .din(new_Jinkela_wire_14739),
        .dout(new_Jinkela_wire_14740)
    );

    bfr new_Jinkela_buffer_12300 (
        .din(new_Jinkela_wire_14799),
        .dout(new_Jinkela_wire_14800)
    );

    bfr new_Jinkela_buffer_12243 (
        .din(new_Jinkela_wire_14740),
        .dout(new_Jinkela_wire_14741)
    );

    bfr new_Jinkela_buffer_12401 (
        .din(new_Jinkela_wire_14902),
        .dout(new_Jinkela_wire_14903)
    );

    bfr new_Jinkela_buffer_12244 (
        .din(new_Jinkela_wire_14741),
        .dout(new_Jinkela_wire_14742)
    );

    bfr new_Jinkela_buffer_12301 (
        .din(new_Jinkela_wire_14800),
        .dout(new_Jinkela_wire_14801)
    );

    bfr new_Jinkela_buffer_12245 (
        .din(new_Jinkela_wire_14742),
        .dout(new_Jinkela_wire_14743)
    );

    bfr new_Jinkela_buffer_12492 (
        .din(new_Jinkela_wire_14995),
        .dout(new_Jinkela_wire_14996)
    );

    bfr new_Jinkela_buffer_12246 (
        .din(new_Jinkela_wire_14743),
        .dout(new_Jinkela_wire_14744)
    );

    bfr new_Jinkela_buffer_12302 (
        .din(new_Jinkela_wire_14801),
        .dout(new_Jinkela_wire_14802)
    );

    bfr new_Jinkela_buffer_12247 (
        .din(new_Jinkela_wire_14744),
        .dout(new_Jinkela_wire_14745)
    );

    bfr new_Jinkela_buffer_12402 (
        .din(new_Jinkela_wire_14903),
        .dout(new_Jinkela_wire_14904)
    );

    bfr new_Jinkela_buffer_12248 (
        .din(new_Jinkela_wire_14745),
        .dout(new_Jinkela_wire_14746)
    );

    bfr new_Jinkela_buffer_12303 (
        .din(new_Jinkela_wire_14802),
        .dout(new_Jinkela_wire_14803)
    );

    bfr new_Jinkela_buffer_12249 (
        .din(new_Jinkela_wire_14746),
        .dout(new_Jinkela_wire_14747)
    );

    bfr new_Jinkela_buffer_12522 (
        .din(new_Jinkela_wire_15029),
        .dout(new_Jinkela_wire_15030)
    );

    bfr new_Jinkela_buffer_12250 (
        .din(new_Jinkela_wire_14747),
        .dout(new_Jinkela_wire_14748)
    );

    bfr new_Jinkela_buffer_12304 (
        .din(new_Jinkela_wire_14803),
        .dout(new_Jinkela_wire_14804)
    );

    or_bb _1951_ (
        .a(new_Jinkela_wire_14089),
        .b(new_Jinkela_wire_9862),
        .c(_0850_)
    );

    or_bb _1952_ (
        .a(new_Jinkela_wire_1570),
        .b(new_Jinkela_wire_16123),
        .c(_0861_)
    );

    or_ii _1953_ (
        .a(new_Jinkela_wire_1571),
        .b(new_Jinkela_wire_16124),
        .c(_0872_)
    );

    or_ii _1954_ (
        .a(new_Jinkela_wire_7740),
        .b(new_Jinkela_wire_20210),
        .c(_0882_)
    );

    and_ii _1955_ (
        .a(new_Jinkela_wire_9738),
        .b(new_Jinkela_wire_4281),
        .c(_0893_)
    );

    and_bb _1956_ (
        .a(new_Jinkela_wire_9739),
        .b(new_Jinkela_wire_4282),
        .c(_0904_)
    );

    or_bb _1957_ (
        .a(new_Jinkela_wire_15835),
        .b(new_Jinkela_wire_6514),
        .c(_0915_)
    );

    or_bb _1958_ (
        .a(new_Jinkela_wire_14030),
        .b(new_Jinkela_wire_10114),
        .c(_0925_)
    );

    or_ii _1959_ (
        .a(new_Jinkela_wire_14031),
        .b(new_Jinkela_wire_10115),
        .c(_0936_)
    );

    or_ii _1960_ (
        .a(new_Jinkela_wire_2128),
        .b(new_Jinkela_wire_19919),
        .c(_0947_)
    );

    and_ii _1961_ (
        .a(new_Jinkela_wire_16512),
        .b(new_Jinkela_wire_20992),
        .c(_0958_)
    );

    and_bb _1962_ (
        .a(new_Jinkela_wire_16513),
        .b(new_Jinkela_wire_20993),
        .c(_0968_)
    );

    or_bb _1963_ (
        .a(new_Jinkela_wire_17089),
        .b(new_Jinkela_wire_13062),
        .c(_0979_)
    );

    or_bb _1964_ (
        .a(new_Jinkela_wire_834),
        .b(new_Jinkela_wire_12063),
        .c(_0989_)
    );

    or_ii _1965_ (
        .a(new_Jinkela_wire_835),
        .b(new_Jinkela_wire_12064),
        .c(_1000_)
    );

    or_ii _1966_ (
        .a(new_Jinkela_wire_21112),
        .b(new_Jinkela_wire_21117),
        .c(_1010_)
    );

    and_ii _1967_ (
        .a(new_Jinkela_wire_8290),
        .b(new_Jinkela_wire_20546),
        .c(_1013_)
    );

    and_bb _1968_ (
        .a(new_Jinkela_wire_8291),
        .b(new_Jinkela_wire_20547),
        .c(_1014_)
    );

    or_bb _1969_ (
        .a(new_Jinkela_wire_7261),
        .b(new_Jinkela_wire_8181),
        .c(_1015_)
    );

    or_bb _1970_ (
        .a(new_Jinkela_wire_14299),
        .b(new_Jinkela_wire_18530),
        .c(_1016_)
    );

    and_bb _1971_ (
        .a(new_Jinkela_wire_303),
        .b(new_Jinkela_wire_349),
        .c(_1017_)
    );

    and_bb _1972_ (
        .a(new_Jinkela_wire_14300),
        .b(new_Jinkela_wire_18531),
        .c(_1018_)
    );

    or_bi _1973_ (
        .a(new_Jinkela_wire_13153),
        .b(new_Jinkela_wire_2946),
        .c(_1019_)
    );

    and_ii _1974_ (
        .a(new_Jinkela_wire_17858),
        .b(new_Jinkela_wire_5041),
        .c(_1020_)
    );

    and_bi _1975_ (
        .a(new_Jinkela_wire_2951),
        .b(new_Jinkela_wire_6859),
        .c(_1021_)
    );

    and_bb _1976_ (
        .a(new_Jinkela_wire_95),
        .b(new_Jinkela_wire_305),
        .c(_1022_)
    );

    and_bi _1977_ (
        .a(new_Jinkela_wire_21122),
        .b(new_Jinkela_wire_8182),
        .c(_1023_)
    );

    and_bb _1978_ (
        .a(new_Jinkela_wire_49),
        .b(new_Jinkela_wire_565),
        .c(_1024_)
    );

    and_bi _1979_ (
        .a(new_Jinkela_wire_19924),
        .b(new_Jinkela_wire_13063),
        .c(_1025_)
    );

    and_bb _1980_ (
        .a(new_Jinkela_wire_276),
        .b(new_Jinkela_wire_643),
        .c(_1026_)
    );

    and_bi _1981_ (
        .a(new_Jinkela_wire_20215),
        .b(new_Jinkela_wire_6515),
        .c(_1027_)
    );

    and_bb _1982_ (
        .a(new_Jinkela_wire_78),
        .b(new_Jinkela_wire_616),
        .c(_1028_)
    );

    and_bi _1983_ (
        .a(new_Jinkela_wire_21189),
        .b(new_Jinkela_wire_9863),
        .c(_1029_)
    );

    and_bb _1984_ (
        .a(new_Jinkela_wire_468),
        .b(new_Jinkela_wire_545),
        .c(_1030_)
    );

    or_ii _1985_ (
        .a(new_Jinkela_wire_685),
        .b(new_Jinkela_wire_318),
        .c(_1031_)
    );

    and_bi _1986_ (
        .a(new_Jinkela_wire_7727),
        .b(new_Jinkela_wire_18109),
        .c(_1032_)
    );

    and_bb _1987_ (
        .a(new_Jinkela_wire_683),
        .b(new_Jinkela_wire_234),
        .c(_1033_)
    );

    and_bi _1988_ (
        .a(new_Jinkela_wire_15778),
        .b(new_Jinkela_wire_3114),
        .c(_1034_)
    );

    and_ii _1989_ (
        .a(new_Jinkela_wire_6994),
        .b(new_Jinkela_wire_7705),
        .c(_1035_)
    );

    or_bb _1990_ (
        .a(new_Jinkela_wire_5546),
        .b(new_Jinkela_wire_5048),
        .c(_1036_)
    );

    or_ii _1991_ (
        .a(new_Jinkela_wire_5547),
        .b(new_Jinkela_wire_5049),
        .c(_1037_)
    );

    or_ii _1992_ (
        .a(new_Jinkela_wire_7979),
        .b(new_Jinkela_wire_10568),
        .c(_1038_)
    );

    bfr new_Jinkela_buffer_8793 (
        .din(new_Jinkela_wire_10780),
        .dout(new_Jinkela_wire_10781)
    );

    bfr new_Jinkela_buffer_8964 (
        .din(new_Jinkela_wire_10961),
        .dout(new_Jinkela_wire_10962)
    );

    bfr new_Jinkela_buffer_8794 (
        .din(new_Jinkela_wire_10781),
        .dout(new_Jinkela_wire_10782)
    );

    bfr new_Jinkela_buffer_8859 (
        .din(new_Jinkela_wire_10850),
        .dout(new_Jinkela_wire_10851)
    );

    bfr new_Jinkela_buffer_8795 (
        .din(new_Jinkela_wire_10782),
        .dout(new_Jinkela_wire_10783)
    );

    bfr new_Jinkela_buffer_8967 (
        .din(new_Jinkela_wire_10964),
        .dout(new_Jinkela_wire_10965)
    );

    bfr new_Jinkela_buffer_8796 (
        .din(new_Jinkela_wire_10783),
        .dout(new_Jinkela_wire_10784)
    );

    bfr new_Jinkela_buffer_8860 (
        .din(new_Jinkela_wire_10851),
        .dout(new_Jinkela_wire_10852)
    );

    bfr new_Jinkela_buffer_8797 (
        .din(new_Jinkela_wire_10784),
        .dout(new_Jinkela_wire_10785)
    );

    bfr new_Jinkela_buffer_9010 (
        .din(_1259_),
        .dout(new_Jinkela_wire_11020)
    );

    bfr new_Jinkela_buffer_8798 (
        .din(new_Jinkela_wire_10785),
        .dout(new_Jinkela_wire_10786)
    );

    bfr new_Jinkela_buffer_8861 (
        .din(new_Jinkela_wire_10852),
        .dout(new_Jinkela_wire_10853)
    );

    bfr new_Jinkela_buffer_8799 (
        .din(new_Jinkela_wire_10786),
        .dout(new_Jinkela_wire_10787)
    );

    bfr new_Jinkela_buffer_8968 (
        .din(new_Jinkela_wire_10965),
        .dout(new_Jinkela_wire_10966)
    );

    bfr new_Jinkela_buffer_8800 (
        .din(new_Jinkela_wire_10787),
        .dout(new_Jinkela_wire_10788)
    );

    bfr new_Jinkela_buffer_8862 (
        .din(new_Jinkela_wire_10853),
        .dout(new_Jinkela_wire_10854)
    );

    bfr new_Jinkela_buffer_8801 (
        .din(new_Jinkela_wire_10788),
        .dout(new_Jinkela_wire_10789)
    );

    bfr new_Jinkela_buffer_8969 (
        .din(_1211_),
        .dout(new_Jinkela_wire_10975)
    );

    bfr new_Jinkela_buffer_8802 (
        .din(new_Jinkela_wire_10789),
        .dout(new_Jinkela_wire_10790)
    );

    bfr new_Jinkela_buffer_8863 (
        .din(new_Jinkela_wire_10854),
        .dout(new_Jinkela_wire_10855)
    );

    bfr new_Jinkela_buffer_8803 (
        .din(new_Jinkela_wire_10790),
        .dout(new_Jinkela_wire_10791)
    );

    spl2 new_Jinkela_splitter_848 (
        .a(new_Jinkela_wire_10966),
        .b(new_Jinkela_wire_10967),
        .c(new_Jinkela_wire_10968)
    );

    bfr new_Jinkela_buffer_8804 (
        .din(new_Jinkela_wire_10791),
        .dout(new_Jinkela_wire_10792)
    );

    bfr new_Jinkela_buffer_8864 (
        .din(new_Jinkela_wire_10855),
        .dout(new_Jinkela_wire_10856)
    );

    bfr new_Jinkela_buffer_8805 (
        .din(new_Jinkela_wire_10792),
        .dout(new_Jinkela_wire_10793)
    );

    bfr new_Jinkela_buffer_8970 (
        .din(new_Jinkela_wire_10975),
        .dout(new_Jinkela_wire_10976)
    );

    bfr new_Jinkela_buffer_8806 (
        .din(new_Jinkela_wire_10793),
        .dout(new_Jinkela_wire_10794)
    );

    bfr new_Jinkela_buffer_8865 (
        .din(new_Jinkela_wire_10856),
        .dout(new_Jinkela_wire_10857)
    );

    bfr new_Jinkela_buffer_8807 (
        .din(new_Jinkela_wire_10794),
        .dout(new_Jinkela_wire_10795)
    );

    spl2 new_Jinkela_splitter_853 (
        .a(_1114_),
        .b(new_Jinkela_wire_11018),
        .c(new_Jinkela_wire_11019)
    );

    bfr new_Jinkela_buffer_8808 (
        .din(new_Jinkela_wire_10795),
        .dout(new_Jinkela_wire_10796)
    );

    bfr new_Jinkela_buffer_8866 (
        .din(new_Jinkela_wire_10857),
        .dout(new_Jinkela_wire_10858)
    );

    bfr new_Jinkela_buffer_8809 (
        .din(new_Jinkela_wire_10796),
        .dout(new_Jinkela_wire_10797)
    );

    bfr new_Jinkela_buffer_9012 (
        .din(_1474_),
        .dout(new_Jinkela_wire_11022)
    );

    bfr new_Jinkela_buffer_8810 (
        .din(new_Jinkela_wire_10797),
        .dout(new_Jinkela_wire_10798)
    );

    bfr new_Jinkela_buffer_8867 (
        .din(new_Jinkela_wire_10858),
        .dout(new_Jinkela_wire_10859)
    );

    bfr new_Jinkela_buffer_8811 (
        .din(new_Jinkela_wire_10798),
        .dout(new_Jinkela_wire_10799)
    );

    bfr new_Jinkela_buffer_8971 (
        .din(new_Jinkela_wire_10976),
        .dout(new_Jinkela_wire_10977)
    );

    bfr new_Jinkela_buffer_8812 (
        .din(new_Jinkela_wire_10799),
        .dout(new_Jinkela_wire_10800)
    );

    bfr new_Jinkela_buffer_8868 (
        .din(new_Jinkela_wire_10859),
        .dout(new_Jinkela_wire_10860)
    );

    bfr new_Jinkela_buffer_8813 (
        .din(new_Jinkela_wire_10800),
        .dout(new_Jinkela_wire_10801)
    );

    bfr new_Jinkela_buffer_9011 (
        .din(_0744_),
        .dout(new_Jinkela_wire_11021)
    );

    bfr new_Jinkela_buffer_12251 (
        .din(new_Jinkela_wire_14748),
        .dout(new_Jinkela_wire_14749)
    );

    bfr new_Jinkela_buffer_12403 (
        .din(new_Jinkela_wire_14904),
        .dout(new_Jinkela_wire_14905)
    );

    bfr new_Jinkela_buffer_12252 (
        .din(new_Jinkela_wire_14749),
        .dout(new_Jinkela_wire_14750)
    );

    bfr new_Jinkela_buffer_12305 (
        .din(new_Jinkela_wire_14804),
        .dout(new_Jinkela_wire_14805)
    );

    bfr new_Jinkela_buffer_12253 (
        .din(new_Jinkela_wire_14750),
        .dout(new_Jinkela_wire_14751)
    );

    bfr new_Jinkela_buffer_12493 (
        .din(new_Jinkela_wire_14996),
        .dout(new_Jinkela_wire_14997)
    );

    bfr new_Jinkela_buffer_12254 (
        .din(new_Jinkela_wire_14751),
        .dout(new_Jinkela_wire_14752)
    );

    bfr new_Jinkela_buffer_12306 (
        .din(new_Jinkela_wire_14805),
        .dout(new_Jinkela_wire_14806)
    );

    bfr new_Jinkela_buffer_12255 (
        .din(new_Jinkela_wire_14752),
        .dout(new_Jinkela_wire_14753)
    );

    bfr new_Jinkela_buffer_12404 (
        .din(new_Jinkela_wire_14905),
        .dout(new_Jinkela_wire_14906)
    );

    bfr new_Jinkela_buffer_12256 (
        .din(new_Jinkela_wire_14753),
        .dout(new_Jinkela_wire_14754)
    );

    bfr new_Jinkela_buffer_12307 (
        .din(new_Jinkela_wire_14806),
        .dout(new_Jinkela_wire_14807)
    );

    bfr new_Jinkela_buffer_12257 (
        .din(new_Jinkela_wire_14754),
        .dout(new_Jinkela_wire_14755)
    );

    bfr new_Jinkela_buffer_12609 (
        .din(_0493_),
        .dout(new_Jinkela_wire_15121)
    );

    spl2 new_Jinkela_splitter_1104 (
        .a(_1829_),
        .b(new_Jinkela_wire_15119),
        .c(new_Jinkela_wire_15120)
    );

    bfr new_Jinkela_buffer_12258 (
        .din(new_Jinkela_wire_14755),
        .dout(new_Jinkela_wire_14756)
    );

    bfr new_Jinkela_buffer_12308 (
        .din(new_Jinkela_wire_14807),
        .dout(new_Jinkela_wire_14808)
    );

    bfr new_Jinkela_buffer_12259 (
        .din(new_Jinkela_wire_14756),
        .dout(new_Jinkela_wire_14757)
    );

    bfr new_Jinkela_buffer_12405 (
        .din(new_Jinkela_wire_14906),
        .dout(new_Jinkela_wire_14907)
    );

    bfr new_Jinkela_buffer_12260 (
        .din(new_Jinkela_wire_14757),
        .dout(new_Jinkela_wire_14758)
    );

    bfr new_Jinkela_buffer_12309 (
        .din(new_Jinkela_wire_14808),
        .dout(new_Jinkela_wire_14809)
    );

    bfr new_Jinkela_buffer_12261 (
        .din(new_Jinkela_wire_14758),
        .dout(new_Jinkela_wire_14759)
    );

    bfr new_Jinkela_buffer_12494 (
        .din(new_Jinkela_wire_14997),
        .dout(new_Jinkela_wire_14998)
    );

    bfr new_Jinkela_buffer_12262 (
        .din(new_Jinkela_wire_14759),
        .dout(new_Jinkela_wire_14760)
    );

    bfr new_Jinkela_buffer_12310 (
        .din(new_Jinkela_wire_14809),
        .dout(new_Jinkela_wire_14810)
    );

    bfr new_Jinkela_buffer_12263 (
        .din(new_Jinkela_wire_14760),
        .dout(new_Jinkela_wire_14761)
    );

    bfr new_Jinkela_buffer_12406 (
        .din(new_Jinkela_wire_14907),
        .dout(new_Jinkela_wire_14908)
    );

    bfr new_Jinkela_buffer_12264 (
        .din(new_Jinkela_wire_14761),
        .dout(new_Jinkela_wire_14762)
    );

    bfr new_Jinkela_buffer_12311 (
        .din(new_Jinkela_wire_14810),
        .dout(new_Jinkela_wire_14811)
    );

    bfr new_Jinkela_buffer_12265 (
        .din(new_Jinkela_wire_14762),
        .dout(new_Jinkela_wire_14763)
    );

    bfr new_Jinkela_buffer_12523 (
        .din(new_Jinkela_wire_15030),
        .dout(new_Jinkela_wire_15031)
    );

    bfr new_Jinkela_buffer_12266 (
        .din(new_Jinkela_wire_14763),
        .dout(new_Jinkela_wire_14764)
    );

    bfr new_Jinkela_buffer_12312 (
        .din(new_Jinkela_wire_14811),
        .dout(new_Jinkela_wire_14812)
    );

    bfr new_Jinkela_buffer_12267 (
        .din(new_Jinkela_wire_14764),
        .dout(new_Jinkela_wire_14765)
    );

    bfr new_Jinkela_buffer_12407 (
        .din(new_Jinkela_wire_14908),
        .dout(new_Jinkela_wire_14909)
    );

    bfr new_Jinkela_buffer_12268 (
        .din(new_Jinkela_wire_14765),
        .dout(new_Jinkela_wire_14766)
    );

    bfr new_Jinkela_buffer_12313 (
        .din(new_Jinkela_wire_14812),
        .dout(new_Jinkela_wire_14813)
    );

    bfr new_Jinkela_buffer_12269 (
        .din(new_Jinkela_wire_14766),
        .dout(new_Jinkela_wire_14767)
    );

    bfr new_Jinkela_buffer_12495 (
        .din(new_Jinkela_wire_14998),
        .dout(new_Jinkela_wire_14999)
    );

    bfr new_Jinkela_buffer_12270 (
        .din(new_Jinkela_wire_14767),
        .dout(new_Jinkela_wire_14768)
    );

    bfr new_Jinkela_buffer_12314 (
        .din(new_Jinkela_wire_14813),
        .dout(new_Jinkela_wire_14814)
    );

    bfr new_Jinkela_buffer_12271 (
        .din(new_Jinkela_wire_14768),
        .dout(new_Jinkela_wire_14769)
    );

    bfr new_Jinkela_buffer_12408 (
        .din(new_Jinkela_wire_14909),
        .dout(new_Jinkela_wire_14910)
    );

    bfr new_Jinkela_buffer_5344 (
        .din(new_Jinkela_wire_6871),
        .dout(new_Jinkela_wire_6872)
    );

    and_ii _2875_ (
        .a(new_Jinkela_wire_10105),
        .b(new_Jinkela_wire_14264),
        .c(_0113_)
    );

    bfr new_Jinkela_buffer_5515 (
        .din(_1058_),
        .dout(new_Jinkela_wire_7053)
    );

    and_ii _2876_ (
        .a(new_Jinkela_wire_1624),
        .b(new_Jinkela_wire_13331),
        .c(_0114_)
    );

    bfr new_Jinkela_buffer_5345 (
        .din(new_Jinkela_wire_6872),
        .dout(new_Jinkela_wire_6873)
    );

    and_bb _2877_ (
        .a(new_Jinkela_wire_1625),
        .b(new_Jinkela_wire_13332),
        .c(_0115_)
    );

    bfr new_Jinkela_buffer_5437 (
        .din(new_Jinkela_wire_6968),
        .dout(new_Jinkela_wire_6969)
    );

    or_bb _2878_ (
        .a(new_Jinkela_wire_3715),
        .b(new_Jinkela_wire_13404),
        .c(_0116_)
    );

    bfr new_Jinkela_buffer_5346 (
        .din(new_Jinkela_wire_6873),
        .dout(new_Jinkela_wire_6874)
    );

    and_ii _2879_ (
        .a(new_Jinkela_wire_1401),
        .b(new_Jinkela_wire_10058),
        .c(_0117_)
    );

    and_bb _2880_ (
        .a(new_Jinkela_wire_1402),
        .b(new_Jinkela_wire_10059),
        .c(_0118_)
    );

    bfr new_Jinkela_buffer_5516 (
        .din(_0627_),
        .dout(new_Jinkela_wire_7054)
    );

    bfr new_Jinkela_buffer_5347 (
        .din(new_Jinkela_wire_6874),
        .dout(new_Jinkela_wire_6875)
    );

    or_bb _2881_ (
        .a(new_Jinkela_wire_10277),
        .b(new_Jinkela_wire_5804),
        .c(_0119_)
    );

    bfr new_Jinkela_buffer_5438 (
        .din(new_Jinkela_wire_6969),
        .dout(new_Jinkela_wire_6970)
    );

    or_bb _2882_ (
        .a(new_Jinkela_wire_18977),
        .b(new_Jinkela_wire_19161),
        .c(_0120_)
    );

    bfr new_Jinkela_buffer_5348 (
        .din(new_Jinkela_wire_6875),
        .dout(new_Jinkela_wire_6876)
    );

    or_ii _2883_ (
        .a(new_Jinkela_wire_18978),
        .b(new_Jinkela_wire_19162),
        .c(_0122_)
    );

    bfr new_Jinkela_buffer_5460 (
        .din(new_Jinkela_wire_6995),
        .dout(new_Jinkela_wire_6996)
    );

    or_ii _2884_ (
        .a(new_Jinkela_wire_5729),
        .b(new_Jinkela_wire_17073),
        .c(_0123_)
    );

    bfr new_Jinkela_buffer_5349 (
        .din(new_Jinkela_wire_6876),
        .dout(new_Jinkela_wire_6877)
    );

    and_ii _2885_ (
        .a(new_Jinkela_wire_21162),
        .b(new_Jinkela_wire_3385),
        .c(_0124_)
    );

    bfr new_Jinkela_buffer_5439 (
        .din(new_Jinkela_wire_6970),
        .dout(new_Jinkela_wire_6971)
    );

    and_bb _2886_ (
        .a(new_Jinkela_wire_21163),
        .b(new_Jinkela_wire_3386),
        .c(_0125_)
    );

    bfr new_Jinkela_buffer_5350 (
        .din(new_Jinkela_wire_6877),
        .dout(new_Jinkela_wire_6878)
    );

    or_bb _2887_ (
        .a(new_Jinkela_wire_2600),
        .b(new_Jinkela_wire_7742),
        .c(_0126_)
    );

    spl2 new_Jinkela_splitter_619 (
        .a(_1488_),
        .b(new_Jinkela_wire_7128),
        .c(new_Jinkela_wire_7129)
    );

    or_bb _2888_ (
        .a(new_Jinkela_wire_1590),
        .b(new_Jinkela_wire_16953),
        .c(_0127_)
    );

    bfr new_Jinkela_buffer_5351 (
        .din(new_Jinkela_wire_6878),
        .dout(new_Jinkela_wire_6879)
    );

    or_ii _2889_ (
        .a(new_Jinkela_wire_1591),
        .b(new_Jinkela_wire_16954),
        .c(_0128_)
    );

    bfr new_Jinkela_buffer_5440 (
        .din(new_Jinkela_wire_6971),
        .dout(new_Jinkela_wire_6972)
    );

    or_ii _2890_ (
        .a(new_Jinkela_wire_4485),
        .b(new_Jinkela_wire_13960),
        .c(_0129_)
    );

    bfr new_Jinkela_buffer_5352 (
        .din(new_Jinkela_wire_6879),
        .dout(new_Jinkela_wire_6880)
    );

    and_ii _2891_ (
        .a(new_Jinkela_wire_6417),
        .b(new_Jinkela_wire_3481),
        .c(_0130_)
    );

    bfr new_Jinkela_buffer_5461 (
        .din(new_Jinkela_wire_6996),
        .dout(new_Jinkela_wire_6997)
    );

    and_bb _2892_ (
        .a(new_Jinkela_wire_6418),
        .b(new_Jinkela_wire_3482),
        .c(_0131_)
    );

    bfr new_Jinkela_buffer_5353 (
        .din(new_Jinkela_wire_6880),
        .dout(new_Jinkela_wire_6881)
    );

    or_bb _2893_ (
        .a(new_Jinkela_wire_7288),
        .b(new_Jinkela_wire_21106),
        .c(_0133_)
    );

    bfr new_Jinkela_buffer_5441 (
        .din(new_Jinkela_wire_6972),
        .dout(new_Jinkela_wire_6973)
    );

    or_bb _2894_ (
        .a(new_Jinkela_wire_17047),
        .b(new_Jinkela_wire_11409),
        .c(_0134_)
    );

    bfr new_Jinkela_buffer_5354 (
        .din(new_Jinkela_wire_6881),
        .dout(new_Jinkela_wire_6882)
    );

    or_ii _2895_ (
        .a(new_Jinkela_wire_17048),
        .b(new_Jinkela_wire_11410),
        .c(_0135_)
    );

    or_ii _2896_ (
        .a(new_Jinkela_wire_19917),
        .b(new_Jinkela_wire_7720),
        .c(_0136_)
    );

    spl2 new_Jinkela_splitter_620 (
        .a(_0064_),
        .b(new_Jinkela_wire_7130),
        .c(new_Jinkela_wire_7131)
    );

    bfr new_Jinkela_buffer_5355 (
        .din(new_Jinkela_wire_6882),
        .dout(new_Jinkela_wire_6883)
    );

    and_ii _2897_ (
        .a(new_Jinkela_wire_1254),
        .b(new_Jinkela_wire_9736),
        .c(_0137_)
    );

    bfr new_Jinkela_buffer_5442 (
        .din(new_Jinkela_wire_6973),
        .dout(new_Jinkela_wire_6974)
    );

    and_bb _2898_ (
        .a(new_Jinkela_wire_1255),
        .b(new_Jinkela_wire_9737),
        .c(_0138_)
    );

    bfr new_Jinkela_buffer_5356 (
        .din(new_Jinkela_wire_6883),
        .dout(new_Jinkela_wire_6884)
    );

    or_bb _2899_ (
        .a(new_Jinkela_wire_3189),
        .b(new_Jinkela_wire_1779),
        .c(_0139_)
    );

    bfr new_Jinkela_buffer_5462 (
        .din(new_Jinkela_wire_6997),
        .dout(new_Jinkela_wire_6998)
    );

    or_bb _2900_ (
        .a(new_Jinkela_wire_15685),
        .b(new_Jinkela_wire_3243),
        .c(_0140_)
    );

    bfr new_Jinkela_buffer_5357 (
        .din(new_Jinkela_wire_6884),
        .dout(new_Jinkela_wire_6885)
    );

    or_ii _2901_ (
        .a(new_Jinkela_wire_15686),
        .b(new_Jinkela_wire_3244),
        .c(_0141_)
    );

    bfr new_Jinkela_buffer_5443 (
        .din(new_Jinkela_wire_6974),
        .dout(new_Jinkela_wire_6975)
    );

    or_ii _2902_ (
        .a(new_Jinkela_wire_4296),
        .b(new_Jinkela_wire_2251),
        .c(_0142_)
    );

    bfr new_Jinkela_buffer_5358 (
        .din(new_Jinkela_wire_6885),
        .dout(new_Jinkela_wire_6886)
    );

    and_ii _2903_ (
        .a(new_Jinkela_wire_8853),
        .b(new_Jinkela_wire_10743),
        .c(_0144_)
    );

    bfr new_Jinkela_buffer_5517 (
        .din(new_Jinkela_wire_7054),
        .dout(new_Jinkela_wire_7055)
    );

    and_bb _2904_ (
        .a(new_Jinkela_wire_8854),
        .b(new_Jinkela_wire_10744),
        .c(_0145_)
    );

    bfr new_Jinkela_buffer_5359 (
        .din(new_Jinkela_wire_6886),
        .dout(new_Jinkela_wire_6887)
    );

    or_bb _2905_ (
        .a(new_Jinkela_wire_20134),
        .b(new_Jinkela_wire_11825),
        .c(_0146_)
    );

    bfr new_Jinkela_buffer_5444 (
        .din(new_Jinkela_wire_6975),
        .dout(new_Jinkela_wire_6976)
    );

    or_bb _2906_ (
        .a(new_Jinkela_wire_8584),
        .b(new_Jinkela_wire_15667),
        .c(_0147_)
    );

    bfr new_Jinkela_buffer_5360 (
        .din(new_Jinkela_wire_6887),
        .dout(new_Jinkela_wire_6888)
    );

    or_ii _2907_ (
        .a(new_Jinkela_wire_8585),
        .b(new_Jinkela_wire_15668),
        .c(_0148_)
    );

    bfr new_Jinkela_buffer_5463 (
        .din(new_Jinkela_wire_6998),
        .dout(new_Jinkela_wire_6999)
    );

    or_ii _2908_ (
        .a(new_Jinkela_wire_2953),
        .b(new_Jinkela_wire_1269),
        .c(_0149_)
    );

    bfr new_Jinkela_buffer_5361 (
        .din(new_Jinkela_wire_6888),
        .dout(new_Jinkela_wire_6889)
    );

    and_ii _2909_ (
        .a(new_Jinkela_wire_16203),
        .b(new_Jinkela_wire_4895),
        .c(_0150_)
    );

    bfr new_Jinkela_buffer_5445 (
        .din(new_Jinkela_wire_6976),
        .dout(new_Jinkela_wire_6977)
    );

    and_bb _2910_ (
        .a(new_Jinkela_wire_16204),
        .b(new_Jinkela_wire_4896),
        .c(_0151_)
    );

    bfr new_Jinkela_buffer_5362 (
        .din(new_Jinkela_wire_6889),
        .dout(new_Jinkela_wire_6890)
    );

    or_bb _2911_ (
        .a(new_Jinkela_wire_6684),
        .b(new_Jinkela_wire_7270),
        .c(_0152_)
    );

    spl2 new_Jinkela_splitter_621 (
        .a(_1350_),
        .b(new_Jinkela_wire_7136),
        .c(new_Jinkela_wire_7137)
    );

    or_bb _2912_ (
        .a(new_Jinkela_wire_706),
        .b(new_Jinkela_wire_19344),
        .c(_0153_)
    );

    bfr new_Jinkela_buffer_5363 (
        .din(new_Jinkela_wire_6890),
        .dout(new_Jinkela_wire_6891)
    );

    or_ii _2913_ (
        .a(new_Jinkela_wire_707),
        .b(new_Jinkela_wire_19345),
        .c(_0155_)
    );

    bfr new_Jinkela_buffer_5446 (
        .din(new_Jinkela_wire_6977),
        .dout(new_Jinkela_wire_6978)
    );

    or_ii _2914_ (
        .a(new_Jinkela_wire_13213),
        .b(new_Jinkela_wire_18702),
        .c(_0156_)
    );

    bfr new_Jinkela_buffer_5364 (
        .din(new_Jinkela_wire_6891),
        .dout(new_Jinkela_wire_6892)
    );

    and_ii _2915_ (
        .a(new_Jinkela_wire_17081),
        .b(new_Jinkela_wire_8093),
        .c(_0157_)
    );

    bfr new_Jinkela_buffer_5464 (
        .din(new_Jinkela_wire_6999),
        .dout(new_Jinkela_wire_7000)
    );

    and_bb _2916_ (
        .a(new_Jinkela_wire_17082),
        .b(new_Jinkela_wire_8094),
        .c(_0158_)
    );

    bfr new_Jinkela_buffer_8814 (
        .din(new_Jinkela_wire_10801),
        .dout(new_Jinkela_wire_10802)
    );

    bfr new_Jinkela_buffer_1874 (
        .din(new_Jinkela_wire_2795),
        .dout(new_Jinkela_wire_2796)
    );

    bfr new_Jinkela_buffer_12272 (
        .din(new_Jinkela_wire_14769),
        .dout(new_Jinkela_wire_14770)
    );

    and_ii _1993_ (
        .a(new_Jinkela_wire_14210),
        .b(new_Jinkela_wire_15769),
        .c(_1039_)
    );

    bfr new_Jinkela_buffer_1774 (
        .din(new_Jinkela_wire_2685),
        .dout(new_Jinkela_wire_2686)
    );

    bfr new_Jinkela_buffer_12315 (
        .din(new_Jinkela_wire_14814),
        .dout(new_Jinkela_wire_14815)
    );

    bfr new_Jinkela_buffer_8869 (
        .din(new_Jinkela_wire_10860),
        .dout(new_Jinkela_wire_10861)
    );

    and_bb _1994_ (
        .a(new_Jinkela_wire_14211),
        .b(new_Jinkela_wire_15770),
        .c(_1040_)
    );

    bfr new_Jinkela_buffer_1809 (
        .din(new_Jinkela_wire_2724),
        .dout(new_Jinkela_wire_2725)
    );

    bfr new_Jinkela_buffer_12273 (
        .din(new_Jinkela_wire_14770),
        .dout(new_Jinkela_wire_14771)
    );

    bfr new_Jinkela_buffer_8815 (
        .din(new_Jinkela_wire_10802),
        .dout(new_Jinkela_wire_10803)
    );

    or_bb _1995_ (
        .a(new_Jinkela_wire_13979),
        .b(new_Jinkela_wire_11386),
        .c(_1041_)
    );

    bfr new_Jinkela_buffer_1775 (
        .din(new_Jinkela_wire_2686),
        .dout(new_Jinkela_wire_2687)
    );

    spl2 new_Jinkela_splitter_1106 (
        .a(_0073_),
        .b(new_Jinkela_wire_15124),
        .c(new_Jinkela_wire_15125)
    );

    bfr new_Jinkela_buffer_8972 (
        .din(new_Jinkela_wire_10977),
        .dout(new_Jinkela_wire_10978)
    );

    or_bb _1996_ (
        .a(new_Jinkela_wire_19932),
        .b(new_Jinkela_wire_19970),
        .c(_1042_)
    );

    spl2 new_Jinkela_splitter_1108 (
        .a(_1171_),
        .b(new_Jinkela_wire_15200),
        .c(new_Jinkela_wire_15201)
    );

    bfr new_Jinkela_buffer_12274 (
        .din(new_Jinkela_wire_14771),
        .dout(new_Jinkela_wire_14772)
    );

    bfr new_Jinkela_buffer_8816 (
        .din(new_Jinkela_wire_10803),
        .dout(new_Jinkela_wire_10804)
    );

    or_ii _1997_ (
        .a(new_Jinkela_wire_19933),
        .b(new_Jinkela_wire_19971),
        .c(_1043_)
    );

    bfr new_Jinkela_buffer_1776 (
        .din(new_Jinkela_wire_2687),
        .dout(new_Jinkela_wire_2688)
    );

    bfr new_Jinkela_buffer_12316 (
        .din(new_Jinkela_wire_14815),
        .dout(new_Jinkela_wire_14816)
    );

    bfr new_Jinkela_buffer_8870 (
        .din(new_Jinkela_wire_10861),
        .dout(new_Jinkela_wire_10862)
    );

    or_ii _1998_ (
        .a(new_Jinkela_wire_3186),
        .b(new_Jinkela_wire_20340),
        .c(_1044_)
    );

    bfr new_Jinkela_buffer_1810 (
        .din(new_Jinkela_wire_2725),
        .dout(new_Jinkela_wire_2726)
    );

    bfr new_Jinkela_buffer_12275 (
        .din(new_Jinkela_wire_14772),
        .dout(new_Jinkela_wire_14773)
    );

    bfr new_Jinkela_buffer_8817 (
        .din(new_Jinkela_wire_10804),
        .dout(new_Jinkela_wire_10805)
    );

    and_ii _1999_ (
        .a(new_Jinkela_wire_5454),
        .b(new_Jinkela_wire_7866),
        .c(_1045_)
    );

    bfr new_Jinkela_buffer_1777 (
        .din(new_Jinkela_wire_2688),
        .dout(new_Jinkela_wire_2689)
    );

    bfr new_Jinkela_buffer_12409 (
        .din(new_Jinkela_wire_14910),
        .dout(new_Jinkela_wire_14911)
    );

    bfr new_Jinkela_buffer_9028 (
        .din(_0939_),
        .dout(new_Jinkela_wire_11040)
    );

    and_bb _2000_ (
        .a(new_Jinkela_wire_5455),
        .b(new_Jinkela_wire_7867),
        .c(_1046_)
    );

    bfr new_Jinkela_buffer_1900 (
        .din(new_Jinkela_wire_2821),
        .dout(new_Jinkela_wire_2822)
    );

    bfr new_Jinkela_buffer_8818 (
        .din(new_Jinkela_wire_10805),
        .dout(new_Jinkela_wire_10806)
    );

    bfr new_Jinkela_buffer_1875 (
        .din(new_Jinkela_wire_2796),
        .dout(new_Jinkela_wire_2797)
    );

    bfr new_Jinkela_buffer_12276 (
        .din(new_Jinkela_wire_14773),
        .dout(new_Jinkela_wire_14774)
    );

    or_bb _2001_ (
        .a(new_Jinkela_wire_1583),
        .b(new_Jinkela_wire_21204),
        .c(_1047_)
    );

    bfr new_Jinkela_buffer_1778 (
        .din(new_Jinkela_wire_2689),
        .dout(new_Jinkela_wire_2690)
    );

    bfr new_Jinkela_buffer_12317 (
        .din(new_Jinkela_wire_14816),
        .dout(new_Jinkela_wire_14817)
    );

    bfr new_Jinkela_buffer_8871 (
        .din(new_Jinkela_wire_10862),
        .dout(new_Jinkela_wire_10863)
    );

    or_bb _2002_ (
        .a(new_Jinkela_wire_6007),
        .b(new_Jinkela_wire_17045),
        .c(_1048_)
    );

    bfr new_Jinkela_buffer_1811 (
        .din(new_Jinkela_wire_2726),
        .dout(new_Jinkela_wire_2727)
    );

    bfr new_Jinkela_buffer_12277 (
        .din(new_Jinkela_wire_14774),
        .dout(new_Jinkela_wire_14775)
    );

    bfr new_Jinkela_buffer_8819 (
        .din(new_Jinkela_wire_10806),
        .dout(new_Jinkela_wire_10807)
    );

    or_ii _2003_ (
        .a(new_Jinkela_wire_6008),
        .b(new_Jinkela_wire_17046),
        .c(_1049_)
    );

    bfr new_Jinkela_buffer_1779 (
        .din(new_Jinkela_wire_2690),
        .dout(new_Jinkela_wire_2691)
    );

    bfr new_Jinkela_buffer_12496 (
        .din(new_Jinkela_wire_14999),
        .dout(new_Jinkela_wire_15000)
    );

    bfr new_Jinkela_buffer_8973 (
        .din(new_Jinkela_wire_10978),
        .dout(new_Jinkela_wire_10979)
    );

    or_ii _2004_ (
        .a(new_Jinkela_wire_7300),
        .b(new_Jinkela_wire_7836),
        .c(_1050_)
    );

    spl2 new_Jinkela_splitter_1098 (
        .a(new_Jinkela_wire_14775),
        .b(new_Jinkela_wire_14776),
        .c(new_Jinkela_wire_14777)
    );

    bfr new_Jinkela_buffer_8820 (
        .din(new_Jinkela_wire_10807),
        .dout(new_Jinkela_wire_10808)
    );

    and_ii _2005_ (
        .a(new_Jinkela_wire_18225),
        .b(new_Jinkela_wire_19105),
        .c(_1051_)
    );

    bfr new_Jinkela_buffer_1780 (
        .din(new_Jinkela_wire_2691),
        .dout(new_Jinkela_wire_2692)
    );

    bfr new_Jinkela_buffer_12410 (
        .din(new_Jinkela_wire_14911),
        .dout(new_Jinkela_wire_14912)
    );

    bfr new_Jinkela_buffer_8872 (
        .din(new_Jinkela_wire_10863),
        .dout(new_Jinkela_wire_10864)
    );

    and_bb _2006_ (
        .a(new_Jinkela_wire_18226),
        .b(new_Jinkela_wire_19106),
        .c(_1052_)
    );

    bfr new_Jinkela_buffer_1812 (
        .din(new_Jinkela_wire_2727),
        .dout(new_Jinkela_wire_2728)
    );

    bfr new_Jinkela_buffer_12318 (
        .din(new_Jinkela_wire_14817),
        .dout(new_Jinkela_wire_14818)
    );

    bfr new_Jinkela_buffer_8821 (
        .din(new_Jinkela_wire_10808),
        .dout(new_Jinkela_wire_10809)
    );

    or_bb _2007_ (
        .a(new_Jinkela_wire_19793),
        .b(new_Jinkela_wire_19342),
        .c(_1053_)
    );

    bfr new_Jinkela_buffer_1781 (
        .din(new_Jinkela_wire_2692),
        .dout(new_Jinkela_wire_2693)
    );

    bfr new_Jinkela_buffer_12319 (
        .din(new_Jinkela_wire_14818),
        .dout(new_Jinkela_wire_14819)
    );

    or_bb _2008_ (
        .a(new_Jinkela_wire_20217),
        .b(new_Jinkela_wire_16192),
        .c(_1054_)
    );

    bfr new_Jinkela_buffer_2011 (
        .din(new_Jinkela_wire_2936),
        .dout(new_Jinkela_wire_2937)
    );

    spl2 new_Jinkela_splitter_856 (
        .a(_0810_),
        .b(new_Jinkela_wire_11046),
        .c(new_Jinkela_wire_11047)
    );

    bfr new_Jinkela_buffer_8822 (
        .din(new_Jinkela_wire_10809),
        .dout(new_Jinkela_wire_10810)
    );

    bfr new_Jinkela_buffer_1876 (
        .din(new_Jinkela_wire_2797),
        .dout(new_Jinkela_wire_2798)
    );

    bfr new_Jinkela_buffer_12524 (
        .din(new_Jinkela_wire_15031),
        .dout(new_Jinkela_wire_15032)
    );

    or_ii _2009_ (
        .a(new_Jinkela_wire_20218),
        .b(new_Jinkela_wire_16193),
        .c(_1055_)
    );

    bfr new_Jinkela_buffer_1782 (
        .din(new_Jinkela_wire_2693),
        .dout(new_Jinkela_wire_2694)
    );

    bfr new_Jinkela_buffer_12320 (
        .din(new_Jinkela_wire_14819),
        .dout(new_Jinkela_wire_14820)
    );

    bfr new_Jinkela_buffer_8873 (
        .din(new_Jinkela_wire_10864),
        .dout(new_Jinkela_wire_10865)
    );

    or_ii _2010_ (
        .a(new_Jinkela_wire_8018),
        .b(new_Jinkela_wire_7281),
        .c(_1056_)
    );

    bfr new_Jinkela_buffer_1813 (
        .din(new_Jinkela_wire_2728),
        .dout(new_Jinkela_wire_2729)
    );

    bfr new_Jinkela_buffer_12411 (
        .din(new_Jinkela_wire_14912),
        .dout(new_Jinkela_wire_14913)
    );

    bfr new_Jinkela_buffer_8823 (
        .din(new_Jinkela_wire_10810),
        .dout(new_Jinkela_wire_10811)
    );

    and_ii _2011_ (
        .a(new_Jinkela_wire_9744),
        .b(new_Jinkela_wire_9597),
        .c(_1057_)
    );

    bfr new_Jinkela_buffer_1783 (
        .din(new_Jinkela_wire_2694),
        .dout(new_Jinkela_wire_2695)
    );

    bfr new_Jinkela_buffer_12321 (
        .din(new_Jinkela_wire_14820),
        .dout(new_Jinkela_wire_14821)
    );

    bfr new_Jinkela_buffer_8974 (
        .din(new_Jinkela_wire_10979),
        .dout(new_Jinkela_wire_10980)
    );

    and_bb _2012_ (
        .a(new_Jinkela_wire_9745),
        .b(new_Jinkela_wire_9598),
        .c(_1058_)
    );

    bfr new_Jinkela_buffer_12497 (
        .din(new_Jinkela_wire_15000),
        .dout(new_Jinkela_wire_15001)
    );

    bfr new_Jinkela_buffer_8824 (
        .din(new_Jinkela_wire_10811),
        .dout(new_Jinkela_wire_10812)
    );

    or_bb _2013_ (
        .a(new_Jinkela_wire_7053),
        .b(new_Jinkela_wire_8851),
        .c(_1059_)
    );

    bfr new_Jinkela_buffer_1784 (
        .din(new_Jinkela_wire_2695),
        .dout(new_Jinkela_wire_2696)
    );

    bfr new_Jinkela_buffer_12322 (
        .din(new_Jinkela_wire_14821),
        .dout(new_Jinkela_wire_14822)
    );

    bfr new_Jinkela_buffer_8874 (
        .din(new_Jinkela_wire_10865),
        .dout(new_Jinkela_wire_10866)
    );

    or_bb _2014_ (
        .a(new_Jinkela_wire_18700),
        .b(new_Jinkela_wire_5716),
        .c(_1060_)
    );

    bfr new_Jinkela_buffer_1814 (
        .din(new_Jinkela_wire_2729),
        .dout(new_Jinkela_wire_2730)
    );

    bfr new_Jinkela_buffer_12412 (
        .din(new_Jinkela_wire_14913),
        .dout(new_Jinkela_wire_14914)
    );

    bfr new_Jinkela_buffer_8825 (
        .din(new_Jinkela_wire_10812),
        .dout(new_Jinkela_wire_10813)
    );

    or_ii _2015_ (
        .a(new_Jinkela_wire_18701),
        .b(new_Jinkela_wire_5717),
        .c(_1061_)
    );

    bfr new_Jinkela_buffer_1785 (
        .din(new_Jinkela_wire_2696),
        .dout(new_Jinkela_wire_2697)
    );

    bfr new_Jinkela_buffer_12323 (
        .din(new_Jinkela_wire_14822),
        .dout(new_Jinkela_wire_14823)
    );

    bfr new_Jinkela_buffer_9013 (
        .din(new_Jinkela_wire_11022),
        .dout(new_Jinkela_wire_11023)
    );

    or_ii _2016_ (
        .a(new_Jinkela_wire_21166),
        .b(new_Jinkela_wire_1805),
        .c(_1062_)
    );

    bfr new_Jinkela_buffer_1901 (
        .din(new_Jinkela_wire_2822),
        .dout(new_Jinkela_wire_2823)
    );

    bfr new_Jinkela_buffer_8826 (
        .din(new_Jinkela_wire_10813),
        .dout(new_Jinkela_wire_10814)
    );

    bfr new_Jinkela_buffer_1877 (
        .din(new_Jinkela_wire_2798),
        .dout(new_Jinkela_wire_2799)
    );

    and_ii _2017_ (
        .a(new_Jinkela_wire_5735),
        .b(new_Jinkela_wire_10160),
        .c(_1063_)
    );

    bfr new_Jinkela_buffer_1786 (
        .din(new_Jinkela_wire_2697),
        .dout(new_Jinkela_wire_2698)
    );

    bfr new_Jinkela_buffer_12324 (
        .din(new_Jinkela_wire_14823),
        .dout(new_Jinkela_wire_14824)
    );

    bfr new_Jinkela_buffer_8875 (
        .din(new_Jinkela_wire_10866),
        .dout(new_Jinkela_wire_10867)
    );

    and_bb _2018_ (
        .a(new_Jinkela_wire_5736),
        .b(new_Jinkela_wire_10161),
        .c(_1064_)
    );

    bfr new_Jinkela_buffer_1815 (
        .din(new_Jinkela_wire_2730),
        .dout(new_Jinkela_wire_2731)
    );

    bfr new_Jinkela_buffer_12413 (
        .din(new_Jinkela_wire_14914),
        .dout(new_Jinkela_wire_14915)
    );

    bfr new_Jinkela_buffer_8827 (
        .din(new_Jinkela_wire_10814),
        .dout(new_Jinkela_wire_10815)
    );

    or_bb _2019_ (
        .a(new_Jinkela_wire_5420),
        .b(new_Jinkela_wire_8762),
        .c(_1065_)
    );

    bfr new_Jinkela_buffer_1787 (
        .din(new_Jinkela_wire_2698),
        .dout(new_Jinkela_wire_2699)
    );

    bfr new_Jinkela_buffer_12325 (
        .din(new_Jinkela_wire_14824),
        .dout(new_Jinkela_wire_14825)
    );

    bfr new_Jinkela_buffer_8975 (
        .din(new_Jinkela_wire_10980),
        .dout(new_Jinkela_wire_10981)
    );

    or_bb _2020_ (
        .a(new_Jinkela_wire_1592),
        .b(new_Jinkela_wire_16798),
        .c(_1066_)
    );

    bfr new_Jinkela_buffer_12498 (
        .din(new_Jinkela_wire_15001),
        .dout(new_Jinkela_wire_15002)
    );

    bfr new_Jinkela_buffer_8828 (
        .din(new_Jinkela_wire_10815),
        .dout(new_Jinkela_wire_10816)
    );

    and_bb _2021_ (
        .a(new_Jinkela_wire_252),
        .b(new_Jinkela_wire_333),
        .c(_1067_)
    );

    bfr new_Jinkela_buffer_1788 (
        .din(new_Jinkela_wire_2699),
        .dout(new_Jinkela_wire_2700)
    );

    bfr new_Jinkela_buffer_12326 (
        .din(new_Jinkela_wire_14825),
        .dout(new_Jinkela_wire_14826)
    );

    bfr new_Jinkela_buffer_8876 (
        .din(new_Jinkela_wire_10867),
        .dout(new_Jinkela_wire_10868)
    );

    and_bb _2022_ (
        .a(new_Jinkela_wire_1593),
        .b(new_Jinkela_wire_16799),
        .c(_1068_)
    );

    bfr new_Jinkela_buffer_1816 (
        .din(new_Jinkela_wire_2731),
        .dout(new_Jinkela_wire_2732)
    );

    bfr new_Jinkela_buffer_12414 (
        .din(new_Jinkela_wire_14915),
        .dout(new_Jinkela_wire_14916)
    );

    bfr new_Jinkela_buffer_8829 (
        .din(new_Jinkela_wire_10816),
        .dout(new_Jinkela_wire_10817)
    );

    or_bi _2023_ (
        .a(new_Jinkela_wire_5167),
        .b(new_Jinkela_wire_20326),
        .c(_1069_)
    );

    bfr new_Jinkela_buffer_1789 (
        .din(new_Jinkela_wire_2700),
        .dout(new_Jinkela_wire_2701)
    );

    bfr new_Jinkela_buffer_12327 (
        .din(new_Jinkela_wire_14826),
        .dout(new_Jinkela_wire_14827)
    );

    and_ii _2024_ (
        .a(new_Jinkela_wire_13053),
        .b(new_Jinkela_wire_7500),
        .c(_1070_)
    );

    bfr new_Jinkela_buffer_9032 (
        .din(_0931_),
        .dout(new_Jinkela_wire_11048)
    );

    bfr new_Jinkela_buffer_8830 (
        .din(new_Jinkela_wire_10817),
        .dout(new_Jinkela_wire_10818)
    );

    bfr new_Jinkela_buffer_1878 (
        .din(new_Jinkela_wire_2799),
        .dout(new_Jinkela_wire_2800)
    );

    bfr new_Jinkela_buffer_12525 (
        .din(new_Jinkela_wire_15032),
        .dout(new_Jinkela_wire_15033)
    );

    and_bi _2025_ (
        .a(new_Jinkela_wire_20331),
        .b(new_Jinkela_wire_19326),
        .c(_1071_)
    );

    bfr new_Jinkela_buffer_1790 (
        .din(new_Jinkela_wire_2701),
        .dout(new_Jinkela_wire_2702)
    );

    bfr new_Jinkela_buffer_12328 (
        .din(new_Jinkela_wire_14827),
        .dout(new_Jinkela_wire_14828)
    );

    bfr new_Jinkela_buffer_8877 (
        .din(new_Jinkela_wire_10868),
        .dout(new_Jinkela_wire_10869)
    );

    and_bb _2026_ (
        .a(new_Jinkela_wire_105),
        .b(new_Jinkela_wire_262),
        .c(_1072_)
    );

    bfr new_Jinkela_buffer_1817 (
        .din(new_Jinkela_wire_2732),
        .dout(new_Jinkela_wire_2733)
    );

    bfr new_Jinkela_buffer_12415 (
        .din(new_Jinkela_wire_14916),
        .dout(new_Jinkela_wire_14917)
    );

    bfr new_Jinkela_buffer_8831 (
        .din(new_Jinkela_wire_10818),
        .dout(new_Jinkela_wire_10819)
    );

    and_bi _2027_ (
        .a(new_Jinkela_wire_1810),
        .b(new_Jinkela_wire_8763),
        .c(_1073_)
    );

    bfr new_Jinkela_buffer_1791 (
        .din(new_Jinkela_wire_2702),
        .dout(new_Jinkela_wire_2703)
    );

    bfr new_Jinkela_buffer_12329 (
        .din(new_Jinkela_wire_14828),
        .dout(new_Jinkela_wire_14829)
    );

    bfr new_Jinkela_buffer_8976 (
        .din(new_Jinkela_wire_10981),
        .dout(new_Jinkela_wire_10982)
    );

    and_bb _2028_ (
        .a(new_Jinkela_wire_295),
        .b(new_Jinkela_wire_566),
        .c(_1074_)
    );

    bfr new_Jinkela_buffer_8832 (
        .din(new_Jinkela_wire_10819),
        .dout(new_Jinkela_wire_10820)
    );

    spl2 new_Jinkela_splitter_313 (
        .a(_0566_),
        .b(new_Jinkela_wire_2943),
        .c(new_Jinkela_wire_2944)
    );

    bfr new_Jinkela_buffer_12499 (
        .din(new_Jinkela_wire_15002),
        .dout(new_Jinkela_wire_15003)
    );

    and_bi _2029_ (
        .a(new_Jinkela_wire_7286),
        .b(new_Jinkela_wire_8852),
        .c(_1075_)
    );

    bfr new_Jinkela_buffer_1792 (
        .din(new_Jinkela_wire_2703),
        .dout(new_Jinkela_wire_2704)
    );

    bfr new_Jinkela_buffer_12330 (
        .din(new_Jinkela_wire_14829),
        .dout(new_Jinkela_wire_14830)
    );

    bfr new_Jinkela_buffer_8878 (
        .din(new_Jinkela_wire_10869),
        .dout(new_Jinkela_wire_10870)
    );

    and_bb _2030_ (
        .a(new_Jinkela_wire_268),
        .b(new_Jinkela_wire_62),
        .c(_1076_)
    );

    bfr new_Jinkela_buffer_1818 (
        .din(new_Jinkela_wire_2733),
        .dout(new_Jinkela_wire_2734)
    );

    bfr new_Jinkela_buffer_12416 (
        .din(new_Jinkela_wire_14917),
        .dout(new_Jinkela_wire_14918)
    );

    bfr new_Jinkela_buffer_8833 (
        .din(new_Jinkela_wire_10820),
        .dout(new_Jinkela_wire_10821)
    );

    and_bi _2031_ (
        .a(new_Jinkela_wire_7841),
        .b(new_Jinkela_wire_19343),
        .c(_1077_)
    );

    bfr new_Jinkela_buffer_1793 (
        .din(new_Jinkela_wire_2704),
        .dout(new_Jinkela_wire_2705)
    );

    bfr new_Jinkela_buffer_12331 (
        .din(new_Jinkela_wire_14830),
        .dout(new_Jinkela_wire_14831)
    );

    bfr new_Jinkela_buffer_9014 (
        .din(new_Jinkela_wire_11023),
        .dout(new_Jinkela_wire_11024)
    );

    and_bb _2032_ (
        .a(new_Jinkela_wire_82),
        .b(new_Jinkela_wire_638),
        .c(_1078_)
    );

    bfr new_Jinkela_buffer_1902 (
        .din(new_Jinkela_wire_2823),
        .dout(new_Jinkela_wire_2824)
    );

    bfr new_Jinkela_buffer_8834 (
        .din(new_Jinkela_wire_10821),
        .dout(new_Jinkela_wire_10822)
    );

    bfr new_Jinkela_buffer_1879 (
        .din(new_Jinkela_wire_2800),
        .dout(new_Jinkela_wire_2801)
    );

    and_bi _2033_ (
        .a(new_Jinkela_wire_20345),
        .b(new_Jinkela_wire_21205),
        .c(_1079_)
    );

    bfr new_Jinkela_buffer_1794 (
        .din(new_Jinkela_wire_2705),
        .dout(new_Jinkela_wire_2706)
    );

    bfr new_Jinkela_buffer_12610 (
        .din(_0443_),
        .dout(new_Jinkela_wire_15126)
    );

    bfr new_Jinkela_buffer_12332 (
        .din(new_Jinkela_wire_14831),
        .dout(new_Jinkela_wire_14832)
    );

    bfr new_Jinkela_buffer_8879 (
        .din(new_Jinkela_wire_10870),
        .dout(new_Jinkela_wire_10871)
    );

    and_bb _2034_ (
        .a(new_Jinkela_wire_470),
        .b(new_Jinkela_wire_625),
        .c(_1080_)
    );

    bfr new_Jinkela_buffer_1819 (
        .din(new_Jinkela_wire_2734),
        .dout(new_Jinkela_wire_2735)
    );

    bfr new_Jinkela_buffer_5365 (
        .din(new_Jinkela_wire_6892),
        .dout(new_Jinkela_wire_6893)
    );

    bfr new_Jinkela_buffer_1795 (
        .din(new_Jinkela_wire_2706),
        .dout(new_Jinkela_wire_2707)
    );

    bfr new_Jinkela_buffer_5447 (
        .din(new_Jinkela_wire_6978),
        .dout(new_Jinkela_wire_6979)
    );

    bfr new_Jinkela_buffer_5366 (
        .din(new_Jinkela_wire_6893),
        .dout(new_Jinkela_wire_6894)
    );

    bfr new_Jinkela_buffer_1796 (
        .din(new_Jinkela_wire_2707),
        .dout(new_Jinkela_wire_2708)
    );

    bfr new_Jinkela_buffer_5518 (
        .din(new_Jinkela_wire_7055),
        .dout(new_Jinkela_wire_7056)
    );

    bfr new_Jinkela_buffer_1820 (
        .din(new_Jinkela_wire_2735),
        .dout(new_Jinkela_wire_2736)
    );

    bfr new_Jinkela_buffer_5367 (
        .din(new_Jinkela_wire_6894),
        .dout(new_Jinkela_wire_6895)
    );

    spl2 new_Jinkela_splitter_305 (
        .a(new_Jinkela_wire_2708),
        .b(new_Jinkela_wire_2709),
        .c(new_Jinkela_wire_2710)
    );

    bfr new_Jinkela_buffer_5448 (
        .din(new_Jinkela_wire_6979),
        .dout(new_Jinkela_wire_6980)
    );

    bfr new_Jinkela_buffer_1821 (
        .din(new_Jinkela_wire_2736),
        .dout(new_Jinkela_wire_2737)
    );

    bfr new_Jinkela_buffer_5368 (
        .din(new_Jinkela_wire_6895),
        .dout(new_Jinkela_wire_6896)
    );

    bfr new_Jinkela_buffer_1880 (
        .din(new_Jinkela_wire_2801),
        .dout(new_Jinkela_wire_2802)
    );

    bfr new_Jinkela_buffer_5465 (
        .din(new_Jinkela_wire_7000),
        .dout(new_Jinkela_wire_7001)
    );

    bfr new_Jinkela_buffer_5369 (
        .din(new_Jinkela_wire_6896),
        .dout(new_Jinkela_wire_6897)
    );

    bfr new_Jinkela_buffer_1822 (
        .din(new_Jinkela_wire_2737),
        .dout(new_Jinkela_wire_2738)
    );

    bfr new_Jinkela_buffer_5449 (
        .din(new_Jinkela_wire_6980),
        .dout(new_Jinkela_wire_6981)
    );

    bfr new_Jinkela_buffer_1903 (
        .din(new_Jinkela_wire_2824),
        .dout(new_Jinkela_wire_2825)
    );

    bfr new_Jinkela_buffer_1881 (
        .din(new_Jinkela_wire_2802),
        .dout(new_Jinkela_wire_2803)
    );

    bfr new_Jinkela_buffer_5370 (
        .din(new_Jinkela_wire_6897),
        .dout(new_Jinkela_wire_6898)
    );

    bfr new_Jinkela_buffer_1823 (
        .din(new_Jinkela_wire_2738),
        .dout(new_Jinkela_wire_2739)
    );

    bfr new_Jinkela_buffer_5588 (
        .din(new_Jinkela_wire_7131),
        .dout(new_Jinkela_wire_7132)
    );

    bfr new_Jinkela_buffer_5371 (
        .din(new_Jinkela_wire_6898),
        .dout(new_Jinkela_wire_6899)
    );

    bfr new_Jinkela_buffer_1824 (
        .din(new_Jinkela_wire_2739),
        .dout(new_Jinkela_wire_2740)
    );

    bfr new_Jinkela_buffer_5450 (
        .din(new_Jinkela_wire_6981),
        .dout(new_Jinkela_wire_6982)
    );

    bfr new_Jinkela_buffer_2012 (
        .din(new_Jinkela_wire_2937),
        .dout(new_Jinkela_wire_2938)
    );

    bfr new_Jinkela_buffer_1882 (
        .din(new_Jinkela_wire_2803),
        .dout(new_Jinkela_wire_2804)
    );

    bfr new_Jinkela_buffer_5372 (
        .din(new_Jinkela_wire_6899),
        .dout(new_Jinkela_wire_6900)
    );

    bfr new_Jinkela_buffer_1825 (
        .din(new_Jinkela_wire_2740),
        .dout(new_Jinkela_wire_2741)
    );

    bfr new_Jinkela_buffer_5466 (
        .din(new_Jinkela_wire_7001),
        .dout(new_Jinkela_wire_7002)
    );

    bfr new_Jinkela_buffer_5373 (
        .din(new_Jinkela_wire_6900),
        .dout(new_Jinkela_wire_6901)
    );

    bfr new_Jinkela_buffer_1826 (
        .din(new_Jinkela_wire_2741),
        .dout(new_Jinkela_wire_2742)
    );

    bfr new_Jinkela_buffer_5451 (
        .din(new_Jinkela_wire_6982),
        .dout(new_Jinkela_wire_6983)
    );

    bfr new_Jinkela_buffer_1904 (
        .din(new_Jinkela_wire_2825),
        .dout(new_Jinkela_wire_2826)
    );

    bfr new_Jinkela_buffer_1883 (
        .din(new_Jinkela_wire_2804),
        .dout(new_Jinkela_wire_2805)
    );

    bfr new_Jinkela_buffer_5374 (
        .din(new_Jinkela_wire_6901),
        .dout(new_Jinkela_wire_6902)
    );

    bfr new_Jinkela_buffer_1827 (
        .din(new_Jinkela_wire_2742),
        .dout(new_Jinkela_wire_2743)
    );

    bfr new_Jinkela_buffer_5519 (
        .din(new_Jinkela_wire_7056),
        .dout(new_Jinkela_wire_7057)
    );

    bfr new_Jinkela_buffer_5375 (
        .din(new_Jinkela_wire_6902),
        .dout(new_Jinkela_wire_6903)
    );

    bfr new_Jinkela_buffer_1828 (
        .din(new_Jinkela_wire_2743),
        .dout(new_Jinkela_wire_2744)
    );

    bfr new_Jinkela_buffer_5452 (
        .din(new_Jinkela_wire_6983),
        .dout(new_Jinkela_wire_6984)
    );

    bfr new_Jinkela_buffer_1884 (
        .din(new_Jinkela_wire_2805),
        .dout(new_Jinkela_wire_2806)
    );

    bfr new_Jinkela_buffer_5376 (
        .din(new_Jinkela_wire_6903),
        .dout(new_Jinkela_wire_6904)
    );

    bfr new_Jinkela_buffer_1829 (
        .din(new_Jinkela_wire_2744),
        .dout(new_Jinkela_wire_2745)
    );

    bfr new_Jinkela_buffer_5467 (
        .din(new_Jinkela_wire_7002),
        .dout(new_Jinkela_wire_7003)
    );

    bfr new_Jinkela_buffer_2015 (
        .din(_0267_),
        .dout(new_Jinkela_wire_2945)
    );

    bfr new_Jinkela_buffer_5377 (
        .din(new_Jinkela_wire_6904),
        .dout(new_Jinkela_wire_6905)
    );

    bfr new_Jinkela_buffer_1830 (
        .din(new_Jinkela_wire_2745),
        .dout(new_Jinkela_wire_2746)
    );

    bfr new_Jinkela_buffer_5453 (
        .din(new_Jinkela_wire_6984),
        .dout(new_Jinkela_wire_6985)
    );

    bfr new_Jinkela_buffer_1905 (
        .din(new_Jinkela_wire_2826),
        .dout(new_Jinkela_wire_2827)
    );

    bfr new_Jinkela_buffer_1885 (
        .din(new_Jinkela_wire_2806),
        .dout(new_Jinkela_wire_2807)
    );

    bfr new_Jinkela_buffer_5378 (
        .din(new_Jinkela_wire_6905),
        .dout(new_Jinkela_wire_6906)
    );

    bfr new_Jinkela_buffer_1831 (
        .din(new_Jinkela_wire_2746),
        .dout(new_Jinkela_wire_2747)
    );

    bfr new_Jinkela_buffer_5596 (
        .din(_0876_),
        .dout(new_Jinkela_wire_7142)
    );

    bfr new_Jinkela_buffer_5379 (
        .din(new_Jinkela_wire_6906),
        .dout(new_Jinkela_wire_6907)
    );

    bfr new_Jinkela_buffer_1832 (
        .din(new_Jinkela_wire_2747),
        .dout(new_Jinkela_wire_2748)
    );

    bfr new_Jinkela_buffer_5454 (
        .din(new_Jinkela_wire_6985),
        .dout(new_Jinkela_wire_6986)
    );

    bfr new_Jinkela_buffer_2013 (
        .din(new_Jinkela_wire_2938),
        .dout(new_Jinkela_wire_2939)
    );

    bfr new_Jinkela_buffer_1886 (
        .din(new_Jinkela_wire_2807),
        .dout(new_Jinkela_wire_2808)
    );

    bfr new_Jinkela_buffer_5380 (
        .din(new_Jinkela_wire_6907),
        .dout(new_Jinkela_wire_6908)
    );

    bfr new_Jinkela_buffer_1833 (
        .din(new_Jinkela_wire_2748),
        .dout(new_Jinkela_wire_2749)
    );

    bfr new_Jinkela_buffer_5468 (
        .din(new_Jinkela_wire_7003),
        .dout(new_Jinkela_wire_7004)
    );

    bfr new_Jinkela_buffer_5381 (
        .din(new_Jinkela_wire_6908),
        .dout(new_Jinkela_wire_6909)
    );

    bfr new_Jinkela_buffer_1834 (
        .din(new_Jinkela_wire_2749),
        .dout(new_Jinkela_wire_2750)
    );

    bfr new_Jinkela_buffer_5455 (
        .din(new_Jinkela_wire_6986),
        .dout(new_Jinkela_wire_6987)
    );

    bfr new_Jinkela_buffer_1906 (
        .din(new_Jinkela_wire_2827),
        .dout(new_Jinkela_wire_2828)
    );

    bfr new_Jinkela_buffer_1887 (
        .din(new_Jinkela_wire_2808),
        .dout(new_Jinkela_wire_2809)
    );

    bfr new_Jinkela_buffer_5382 (
        .din(new_Jinkela_wire_6909),
        .dout(new_Jinkela_wire_6910)
    );

    bfr new_Jinkela_buffer_1835 (
        .din(new_Jinkela_wire_2750),
        .dout(new_Jinkela_wire_2751)
    );

    bfr new_Jinkela_buffer_5520 (
        .din(new_Jinkela_wire_7057),
        .dout(new_Jinkela_wire_7058)
    );

    bfr new_Jinkela_buffer_5383 (
        .din(new_Jinkela_wire_6910),
        .dout(new_Jinkela_wire_6911)
    );

    bfr new_Jinkela_buffer_1836 (
        .din(new_Jinkela_wire_2751),
        .dout(new_Jinkela_wire_2752)
    );

    bfr new_Jinkela_buffer_5456 (
        .din(new_Jinkela_wire_6987),
        .dout(new_Jinkela_wire_6988)
    );

    bfr new_Jinkela_buffer_2020 (
        .din(_1627_),
        .dout(new_Jinkela_wire_2952)
    );

    bfr new_Jinkela_buffer_1888 (
        .din(new_Jinkela_wire_2809),
        .dout(new_Jinkela_wire_2810)
    );

    bfr new_Jinkela_buffer_5384 (
        .din(new_Jinkela_wire_6911),
        .dout(new_Jinkela_wire_6912)
    );

    bfr new_Jinkela_buffer_1837 (
        .din(new_Jinkela_wire_2752),
        .dout(new_Jinkela_wire_2753)
    );

    bfr new_Jinkela_buffer_5469 (
        .din(new_Jinkela_wire_7004),
        .dout(new_Jinkela_wire_7005)
    );

    spl2 new_Jinkela_splitter_314 (
        .a(_1016_),
        .b(new_Jinkela_wire_2946),
        .c(new_Jinkela_wire_2947)
    );

    bfr new_Jinkela_buffer_5385 (
        .din(new_Jinkela_wire_6912),
        .dout(new_Jinkela_wire_6913)
    );

    bfr new_Jinkela_buffer_1838 (
        .din(new_Jinkela_wire_2753),
        .dout(new_Jinkela_wire_2754)
    );

    bfr new_Jinkela_buffer_5457 (
        .din(new_Jinkela_wire_6988),
        .dout(new_Jinkela_wire_6989)
    );

    bfr new_Jinkela_buffer_1907 (
        .din(new_Jinkela_wire_2828),
        .dout(new_Jinkela_wire_2829)
    );

    bfr new_Jinkela_buffer_8835 (
        .din(new_Jinkela_wire_10822),
        .dout(new_Jinkela_wire_10823)
    );

    bfr new_Jinkela_buffer_8977 (
        .din(new_Jinkela_wire_10982),
        .dout(new_Jinkela_wire_10983)
    );

    bfr new_Jinkela_buffer_8836 (
        .din(new_Jinkela_wire_10823),
        .dout(new_Jinkela_wire_10824)
    );

    bfr new_Jinkela_buffer_8880 (
        .din(new_Jinkela_wire_10871),
        .dout(new_Jinkela_wire_10872)
    );

    bfr new_Jinkela_buffer_8837 (
        .din(new_Jinkela_wire_10824),
        .dout(new_Jinkela_wire_10825)
    );

    bfr new_Jinkela_buffer_9029 (
        .din(new_Jinkela_wire_11040),
        .dout(new_Jinkela_wire_11041)
    );

    bfr new_Jinkela_buffer_8838 (
        .din(new_Jinkela_wire_10825),
        .dout(new_Jinkela_wire_10826)
    );

    bfr new_Jinkela_buffer_8881 (
        .din(new_Jinkela_wire_10872),
        .dout(new_Jinkela_wire_10873)
    );

    bfr new_Jinkela_buffer_8839 (
        .din(new_Jinkela_wire_10826),
        .dout(new_Jinkela_wire_10827)
    );

    bfr new_Jinkela_buffer_8978 (
        .din(new_Jinkela_wire_10983),
        .dout(new_Jinkela_wire_10984)
    );

    bfr new_Jinkela_buffer_8840 (
        .din(new_Jinkela_wire_10827),
        .dout(new_Jinkela_wire_10828)
    );

    bfr new_Jinkela_buffer_8882 (
        .din(new_Jinkela_wire_10873),
        .dout(new_Jinkela_wire_10874)
    );

    bfr new_Jinkela_buffer_8841 (
        .din(new_Jinkela_wire_10828),
        .dout(new_Jinkela_wire_10829)
    );

    bfr new_Jinkela_buffer_9015 (
        .din(new_Jinkela_wire_11024),
        .dout(new_Jinkela_wire_11025)
    );

    bfr new_Jinkela_buffer_8842 (
        .din(new_Jinkela_wire_10829),
        .dout(new_Jinkela_wire_10830)
    );

    bfr new_Jinkela_buffer_8883 (
        .din(new_Jinkela_wire_10874),
        .dout(new_Jinkela_wire_10875)
    );

    bfr new_Jinkela_buffer_8843 (
        .din(new_Jinkela_wire_10830),
        .dout(new_Jinkela_wire_10831)
    );

    bfr new_Jinkela_buffer_8979 (
        .din(new_Jinkela_wire_10984),
        .dout(new_Jinkela_wire_10985)
    );

    bfr new_Jinkela_buffer_8844 (
        .din(new_Jinkela_wire_10831),
        .dout(new_Jinkela_wire_10832)
    );

    bfr new_Jinkela_buffer_8884 (
        .din(new_Jinkela_wire_10875),
        .dout(new_Jinkela_wire_10876)
    );

    spl2 new_Jinkela_splitter_843 (
        .a(new_Jinkela_wire_10832),
        .b(new_Jinkela_wire_10833),
        .c(new_Jinkela_wire_10834)
    );

    bfr new_Jinkela_buffer_8885 (
        .din(new_Jinkela_wire_10876),
        .dout(new_Jinkela_wire_10877)
    );

    spl2 new_Jinkela_splitter_860 (
        .a(_1496_),
        .b(new_Jinkela_wire_11228),
        .c(new_Jinkela_wire_11229)
    );

    bfr new_Jinkela_buffer_8980 (
        .din(new_Jinkela_wire_10985),
        .dout(new_Jinkela_wire_10986)
    );

    bfr new_Jinkela_buffer_8886 (
        .din(new_Jinkela_wire_10877),
        .dout(new_Jinkela_wire_10878)
    );

    bfr new_Jinkela_buffer_9016 (
        .din(new_Jinkela_wire_11025),
        .dout(new_Jinkela_wire_11026)
    );

    bfr new_Jinkela_buffer_8887 (
        .din(new_Jinkela_wire_10878),
        .dout(new_Jinkela_wire_10879)
    );

    bfr new_Jinkela_buffer_8981 (
        .din(new_Jinkela_wire_10986),
        .dout(new_Jinkela_wire_10987)
    );

    bfr new_Jinkela_buffer_8888 (
        .din(new_Jinkela_wire_10879),
        .dout(new_Jinkela_wire_10880)
    );

    bfr new_Jinkela_buffer_9030 (
        .din(new_Jinkela_wire_11041),
        .dout(new_Jinkela_wire_11042)
    );

    bfr new_Jinkela_buffer_8889 (
        .din(new_Jinkela_wire_10880),
        .dout(new_Jinkela_wire_10881)
    );

    bfr new_Jinkela_buffer_8982 (
        .din(new_Jinkela_wire_10987),
        .dout(new_Jinkela_wire_10988)
    );

    bfr new_Jinkela_buffer_8890 (
        .din(new_Jinkela_wire_10881),
        .dout(new_Jinkela_wire_10882)
    );

    bfr new_Jinkela_buffer_9017 (
        .din(new_Jinkela_wire_11026),
        .dout(new_Jinkela_wire_11027)
    );

    bfr new_Jinkela_buffer_8891 (
        .din(new_Jinkela_wire_10882),
        .dout(new_Jinkela_wire_10883)
    );

    bfr new_Jinkela_buffer_8983 (
        .din(new_Jinkela_wire_10988),
        .dout(new_Jinkela_wire_10989)
    );

    bfr new_Jinkela_buffer_8892 (
        .din(new_Jinkela_wire_10883),
        .dout(new_Jinkela_wire_10884)
    );

    bfr new_Jinkela_buffer_8893 (
        .din(new_Jinkela_wire_10884),
        .dout(new_Jinkela_wire_10885)
    );

    bfr new_Jinkela_buffer_8984 (
        .din(new_Jinkela_wire_10989),
        .dout(new_Jinkela_wire_10990)
    );

    bfr new_Jinkela_buffer_8894 (
        .din(new_Jinkela_wire_10885),
        .dout(new_Jinkela_wire_10886)
    );

    bfr new_Jinkela_buffer_9018 (
        .din(new_Jinkela_wire_11027),
        .dout(new_Jinkela_wire_11028)
    );

    bfr new_Jinkela_buffer_15775 (
        .din(new_Jinkela_wire_18801),
        .dout(new_Jinkela_wire_18802)
    );

    bfr new_Jinkela_buffer_15780 (
        .din(_0349_),
        .dout(new_Jinkela_wire_18809)
    );

    bfr new_Jinkela_buffer_15776 (
        .din(new_Jinkela_wire_18802),
        .dout(new_Jinkela_wire_18803)
    );

    bfr new_Jinkela_buffer_15802 (
        .din(_0499_),
        .dout(new_Jinkela_wire_18833)
    );

    bfr new_Jinkela_buffer_15786 (
        .din(new_Jinkela_wire_18814),
        .dout(new_Jinkela_wire_18815)
    );

    spl2 new_Jinkela_splitter_1364 (
        .a(_1822_),
        .b(new_Jinkela_wire_18834),
        .c(new_Jinkela_wire_18835)
    );

    bfr new_Jinkela_buffer_15781 (
        .din(new_Jinkela_wire_18809),
        .dout(new_Jinkela_wire_18810)
    );

    bfr new_Jinkela_buffer_15803 (
        .din(_0831_),
        .dout(new_Jinkela_wire_18836)
    );

    bfr new_Jinkela_buffer_15782 (
        .din(new_Jinkela_wire_18810),
        .dout(new_Jinkela_wire_18811)
    );

    spl2 new_Jinkela_splitter_1367 (
        .a(_0933_),
        .b(new_Jinkela_wire_18944),
        .c(new_Jinkela_wire_18945)
    );

    bfr new_Jinkela_buffer_15783 (
        .din(new_Jinkela_wire_18811),
        .dout(new_Jinkela_wire_18812)
    );

    spl2 new_Jinkela_splitter_1366 (
        .a(_1612_),
        .b(new_Jinkela_wire_18942),
        .c(new_Jinkela_wire_18943)
    );

    bfr new_Jinkela_buffer_15784 (
        .din(new_Jinkela_wire_18812),
        .dout(new_Jinkela_wire_18813)
    );

    bfr new_Jinkela_buffer_15804 (
        .din(new_Jinkela_wire_18836),
        .dout(new_Jinkela_wire_18837)
    );

    bfr new_Jinkela_buffer_15785 (
        .din(new_Jinkela_wire_18813),
        .dout(new_Jinkela_wire_18814)
    );

    bfr new_Jinkela_buffer_15805 (
        .din(new_Jinkela_wire_18837),
        .dout(new_Jinkela_wire_18838)
    );

    bfr new_Jinkela_buffer_15787 (
        .din(new_Jinkela_wire_18815),
        .dout(new_Jinkela_wire_18816)
    );

    spl2 new_Jinkela_splitter_1368 (
        .a(_1635_),
        .b(new_Jinkela_wire_18950),
        .c(new_Jinkela_wire_18951)
    );

    bfr new_Jinkela_buffer_15788 (
        .din(new_Jinkela_wire_18816),
        .dout(new_Jinkela_wire_18817)
    );

    bfr new_Jinkela_buffer_15806 (
        .din(new_Jinkela_wire_18838),
        .dout(new_Jinkela_wire_18839)
    );

    bfr new_Jinkela_buffer_15789 (
        .din(new_Jinkela_wire_18817),
        .dout(new_Jinkela_wire_18818)
    );

    bfr new_Jinkela_buffer_15907 (
        .din(new_Jinkela_wire_18945),
        .dout(new_Jinkela_wire_18946)
    );

    bfr new_Jinkela_buffer_15911 (
        .din(_1716_),
        .dout(new_Jinkela_wire_18952)
    );

    bfr new_Jinkela_buffer_15790 (
        .din(new_Jinkela_wire_18818),
        .dout(new_Jinkela_wire_18819)
    );

    bfr new_Jinkela_buffer_15807 (
        .din(new_Jinkela_wire_18839),
        .dout(new_Jinkela_wire_18840)
    );

    bfr new_Jinkela_buffer_15791 (
        .din(new_Jinkela_wire_18819),
        .dout(new_Jinkela_wire_18820)
    );

    bfr new_Jinkela_buffer_15792 (
        .din(new_Jinkela_wire_18820),
        .dout(new_Jinkela_wire_18821)
    );

    bfr new_Jinkela_buffer_15808 (
        .din(new_Jinkela_wire_18840),
        .dout(new_Jinkela_wire_18841)
    );

    bfr new_Jinkela_buffer_15793 (
        .din(new_Jinkela_wire_18821),
        .dout(new_Jinkela_wire_18822)
    );

    bfr new_Jinkela_buffer_15908 (
        .din(new_Jinkela_wire_18946),
        .dout(new_Jinkela_wire_18947)
    );

    bfr new_Jinkela_buffer_15794 (
        .din(new_Jinkela_wire_18822),
        .dout(new_Jinkela_wire_18823)
    );

    bfr new_Jinkela_buffer_15809 (
        .din(new_Jinkela_wire_18841),
        .dout(new_Jinkela_wire_18842)
    );

    bfr new_Jinkela_buffer_15795 (
        .din(new_Jinkela_wire_18823),
        .dout(new_Jinkela_wire_18824)
    );

    spl2 new_Jinkela_splitter_1370 (
        .a(_0649_),
        .b(new_Jinkela_wire_18955),
        .c(new_Jinkela_wire_18956)
    );

    spl2 new_Jinkela_splitter_1369 (
        .a(_1688_),
        .b(new_Jinkela_wire_18953),
        .c(new_Jinkela_wire_18954)
    );

    bfr new_Jinkela_buffer_15796 (
        .din(new_Jinkela_wire_18824),
        .dout(new_Jinkela_wire_18825)
    );

    bfr new_Jinkela_buffer_15810 (
        .din(new_Jinkela_wire_18842),
        .dout(new_Jinkela_wire_18843)
    );

    bfr new_Jinkela_buffer_15797 (
        .din(new_Jinkela_wire_18825),
        .dout(new_Jinkela_wire_18826)
    );

    bfr new_Jinkela_buffer_15909 (
        .din(new_Jinkela_wire_18947),
        .dout(new_Jinkela_wire_18948)
    );

    bfr new_Jinkela_buffer_15798 (
        .din(new_Jinkela_wire_18826),
        .dout(new_Jinkela_wire_18827)
    );

    bfr new_Jinkela_buffer_15811 (
        .din(new_Jinkela_wire_18843),
        .dout(new_Jinkela_wire_18844)
    );

    bfr new_Jinkela_buffer_15799 (
        .din(new_Jinkela_wire_18827),
        .dout(new_Jinkela_wire_18828)
    );

    or_bb _2917_ (
        .a(new_Jinkela_wire_8865),
        .b(new_Jinkela_wire_15697),
        .c(_0159_)
    );

    or_bb _2918_ (
        .a(new_Jinkela_wire_4724),
        .b(new_Jinkela_wire_10971),
        .c(_0160_)
    );

    or_ii _2919_ (
        .a(new_Jinkela_wire_4725),
        .b(new_Jinkela_wire_10972),
        .c(_0161_)
    );

    or_ii _2920_ (
        .a(new_Jinkela_wire_5051),
        .b(new_Jinkela_wire_10562),
        .c(_0162_)
    );

    and_ii _2921_ (
        .a(new_Jinkela_wire_1586),
        .b(new_Jinkela_wire_16774),
        .c(_0163_)
    );

    and_bb _2922_ (
        .a(new_Jinkela_wire_1587),
        .b(new_Jinkela_wire_16775),
        .c(_0164_)
    );

    or_bb _2923_ (
        .a(new_Jinkela_wire_9564),
        .b(new_Jinkela_wire_12627),
        .c(_0166_)
    );

    or_bb _2924_ (
        .a(new_Jinkela_wire_12905),
        .b(new_Jinkela_wire_8480),
        .c(_0167_)
    );

    or_ii _2925_ (
        .a(new_Jinkela_wire_12906),
        .b(new_Jinkela_wire_8481),
        .c(_0168_)
    );

    or_ii _2926_ (
        .a(new_Jinkela_wire_21113),
        .b(new_Jinkela_wire_1602),
        .c(_0169_)
    );

    and_ii _2927_ (
        .a(new_Jinkela_wire_6680),
        .b(new_Jinkela_wire_7831),
        .c(_0170_)
    );

    and_bb _2928_ (
        .a(new_Jinkela_wire_6681),
        .b(new_Jinkela_wire_7832),
        .c(_0171_)
    );

    or_bb _2929_ (
        .a(new_Jinkela_wire_13322),
        .b(new_Jinkela_wire_3667),
        .c(_0172_)
    );

    or_bb _2930_ (
        .a(new_Jinkela_wire_11959),
        .b(new_Jinkela_wire_13310),
        .c(_0173_)
    );

    or_ii _2931_ (
        .a(new_Jinkela_wire_11960),
        .b(new_Jinkela_wire_13311),
        .c(_0174_)
    );

    or_ii _2932_ (
        .a(new_Jinkela_wire_19047),
        .b(new_Jinkela_wire_6001),
        .c(_0175_)
    );

    and_ii _2933_ (
        .a(new_Jinkela_wire_7845),
        .b(new_Jinkela_wire_13304),
        .c(_0177_)
    );

    and_bb _2934_ (
        .a(new_Jinkela_wire_7846),
        .b(new_Jinkela_wire_13305),
        .c(_0178_)
    );

    or_bb _2935_ (
        .a(new_Jinkela_wire_14272),
        .b(new_Jinkela_wire_9173),
        .c(_0179_)
    );

    or_bb _2936_ (
        .a(new_Jinkela_wire_5127),
        .b(new_Jinkela_wire_17022),
        .c(_0180_)
    );

    or_ii _2937_ (
        .a(new_Jinkela_wire_5128),
        .b(new_Jinkela_wire_17023),
        .c(_0181_)
    );

    or_ii _2938_ (
        .a(new_Jinkela_wire_14021),
        .b(new_Jinkela_wire_3247),
        .c(_0182_)
    );

    and_ii _2939_ (
        .a(new_Jinkela_wire_13147),
        .b(new_Jinkela_wire_2249),
        .c(_0183_)
    );

    and_bb _2940_ (
        .a(new_Jinkela_wire_13148),
        .b(new_Jinkela_wire_2250),
        .c(_0184_)
    );

    or_bb _2941_ (
        .a(new_Jinkela_wire_5886),
        .b(new_Jinkela_wire_1616),
        .c(_0185_)
    );

    or_bb _2942_ (
        .a(new_Jinkela_wire_16967),
        .b(new_Jinkela_wire_6810),
        .c(_0186_)
    );

    or_ii _2943_ (
        .a(new_Jinkela_wire_16968),
        .b(new_Jinkela_wire_6811),
        .c(_0188_)
    );

    or_ii _2944_ (
        .a(new_Jinkela_wire_11533),
        .b(new_Jinkela_wire_13587),
        .c(_0189_)
    );

    and_ii _2945_ (
        .a(new_Jinkela_wire_17656),
        .b(new_Jinkela_wire_21324),
        .c(_0190_)
    );

    and_bb _2946_ (
        .a(new_Jinkela_wire_17657),
        .b(new_Jinkela_wire_21325),
        .c(_0191_)
    );

    or_bb _2947_ (
        .a(new_Jinkela_wire_14201),
        .b(new_Jinkela_wire_8764),
        .c(_0192_)
    );

    or_bb _2948_ (
        .a(new_Jinkela_wire_19190),
        .b(new_Jinkela_wire_13339),
        .c(_0193_)
    );

    or_ii _2949_ (
        .a(new_Jinkela_wire_19191),
        .b(new_Jinkela_wire_13340),
        .c(_0194_)
    );

    or_ii _2950_ (
        .a(new_Jinkela_wire_2319),
        .b(new_Jinkela_wire_19560),
        .c(_0195_)
    );

    and_ii _2951_ (
        .a(new_Jinkela_wire_4539),
        .b(new_Jinkela_wire_7438),
        .c(_0196_)
    );

    and_bb _2952_ (
        .a(new_Jinkela_wire_4540),
        .b(new_Jinkela_wire_7439),
        .c(_0197_)
    );

    or_bb _2953_ (
        .a(new_Jinkela_wire_17055),
        .b(new_Jinkela_wire_7712),
        .c(_0199_)
    );

    and_ii _2954_ (
        .a(new_Jinkela_wire_12713),
        .b(new_Jinkela_wire_4722),
        .c(_0200_)
    );

    and_bb _2955_ (
        .a(new_Jinkela_wire_12714),
        .b(new_Jinkela_wire_4723),
        .c(_0201_)
    );

    or_bb _2956_ (
        .a(new_Jinkela_wire_16113),
        .b(new_Jinkela_wire_20805),
        .c(_0202_)
    );

    or_bb _2957_ (
        .a(new_Jinkela_wire_2146),
        .b(new_Jinkela_wire_3957),
        .c(_0203_)
    );

    and_bb _2958_ (
        .a(new_Jinkela_wire_16782),
        .b(new_Jinkela_wire_13845),
        .c(_0204_)
    );

    bfr new_Jinkela_buffer_5386 (
        .din(new_Jinkela_wire_6913),
        .dout(new_Jinkela_wire_6914)
    );

    bfr new_Jinkela_buffer_5592 (
        .din(new_Jinkela_wire_7137),
        .dout(new_Jinkela_wire_7138)
    );

    bfr new_Jinkela_buffer_5387 (
        .din(new_Jinkela_wire_6914),
        .dout(new_Jinkela_wire_6915)
    );

    spl2 new_Jinkela_splitter_615 (
        .a(new_Jinkela_wire_6989),
        .b(new_Jinkela_wire_6990),
        .c(new_Jinkela_wire_6991)
    );

    bfr new_Jinkela_buffer_5388 (
        .din(new_Jinkela_wire_6915),
        .dout(new_Jinkela_wire_6916)
    );

    bfr new_Jinkela_buffer_5521 (
        .din(new_Jinkela_wire_7058),
        .dout(new_Jinkela_wire_7059)
    );

    bfr new_Jinkela_buffer_5389 (
        .din(new_Jinkela_wire_6916),
        .dout(new_Jinkela_wire_6917)
    );

    bfr new_Jinkela_buffer_5470 (
        .din(new_Jinkela_wire_7005),
        .dout(new_Jinkela_wire_7006)
    );

    bfr new_Jinkela_buffer_5390 (
        .din(new_Jinkela_wire_6917),
        .dout(new_Jinkela_wire_6918)
    );

    bfr new_Jinkela_buffer_5471 (
        .din(new_Jinkela_wire_7006),
        .dout(new_Jinkela_wire_7007)
    );

    bfr new_Jinkela_buffer_5391 (
        .din(new_Jinkela_wire_6918),
        .dout(new_Jinkela_wire_6919)
    );

    bfr new_Jinkela_buffer_5589 (
        .din(new_Jinkela_wire_7132),
        .dout(new_Jinkela_wire_7133)
    );

    bfr new_Jinkela_buffer_5392 (
        .din(new_Jinkela_wire_6919),
        .dout(new_Jinkela_wire_6920)
    );

    bfr new_Jinkela_buffer_5472 (
        .din(new_Jinkela_wire_7007),
        .dout(new_Jinkela_wire_7008)
    );

    bfr new_Jinkela_buffer_5393 (
        .din(new_Jinkela_wire_6920),
        .dout(new_Jinkela_wire_6921)
    );

    bfr new_Jinkela_buffer_5522 (
        .din(new_Jinkela_wire_7059),
        .dout(new_Jinkela_wire_7060)
    );

    bfr new_Jinkela_buffer_5394 (
        .din(new_Jinkela_wire_6921),
        .dout(new_Jinkela_wire_6922)
    );

    bfr new_Jinkela_buffer_5473 (
        .din(new_Jinkela_wire_7008),
        .dout(new_Jinkela_wire_7009)
    );

    bfr new_Jinkela_buffer_5395 (
        .din(new_Jinkela_wire_6922),
        .dout(new_Jinkela_wire_6923)
    );

    bfr new_Jinkela_buffer_5396 (
        .din(new_Jinkela_wire_6923),
        .dout(new_Jinkela_wire_6924)
    );

    bfr new_Jinkela_buffer_5474 (
        .din(new_Jinkela_wire_7009),
        .dout(new_Jinkela_wire_7010)
    );

    bfr new_Jinkela_buffer_5397 (
        .din(new_Jinkela_wire_6924),
        .dout(new_Jinkela_wire_6925)
    );

    bfr new_Jinkela_buffer_5523 (
        .din(new_Jinkela_wire_7060),
        .dout(new_Jinkela_wire_7061)
    );

    bfr new_Jinkela_buffer_5398 (
        .din(new_Jinkela_wire_6925),
        .dout(new_Jinkela_wire_6926)
    );

    bfr new_Jinkela_buffer_5475 (
        .din(new_Jinkela_wire_7010),
        .dout(new_Jinkela_wire_7011)
    );

    bfr new_Jinkela_buffer_5399 (
        .din(new_Jinkela_wire_6926),
        .dout(new_Jinkela_wire_6927)
    );

    bfr new_Jinkela_buffer_5590 (
        .din(new_Jinkela_wire_7133),
        .dout(new_Jinkela_wire_7134)
    );

    bfr new_Jinkela_buffer_5400 (
        .din(new_Jinkela_wire_6927),
        .dout(new_Jinkela_wire_6928)
    );

    bfr new_Jinkela_buffer_5476 (
        .din(new_Jinkela_wire_7011),
        .dout(new_Jinkela_wire_7012)
    );

    bfr new_Jinkela_buffer_5401 (
        .din(new_Jinkela_wire_6928),
        .dout(new_Jinkela_wire_6929)
    );

    bfr new_Jinkela_buffer_5524 (
        .din(new_Jinkela_wire_7061),
        .dout(new_Jinkela_wire_7062)
    );

    bfr new_Jinkela_buffer_5402 (
        .din(new_Jinkela_wire_6929),
        .dout(new_Jinkela_wire_6930)
    );

    bfr new_Jinkela_buffer_5477 (
        .din(new_Jinkela_wire_7012),
        .dout(new_Jinkela_wire_7013)
    );

    bfr new_Jinkela_buffer_5403 (
        .din(new_Jinkela_wire_6930),
        .dout(new_Jinkela_wire_6931)
    );

    bfr new_Jinkela_buffer_5628 (
        .din(new_Jinkela_wire_7177),
        .dout(new_Jinkela_wire_7178)
    );

    bfr new_Jinkela_buffer_5404 (
        .din(new_Jinkela_wire_6931),
        .dout(new_Jinkela_wire_6932)
    );

    bfr new_Jinkela_buffer_5478 (
        .din(new_Jinkela_wire_7013),
        .dout(new_Jinkela_wire_7014)
    );

    bfr new_Jinkela_buffer_5405 (
        .din(new_Jinkela_wire_6932),
        .dout(new_Jinkela_wire_6933)
    );

    bfr new_Jinkela_buffer_5525 (
        .din(new_Jinkela_wire_7062),
        .dout(new_Jinkela_wire_7063)
    );

    bfr new_Jinkela_buffer_5406 (
        .din(new_Jinkela_wire_6933),
        .dout(new_Jinkela_wire_6934)
    );

    bfr new_Jinkela_buffer_5479 (
        .din(new_Jinkela_wire_7014),
        .dout(new_Jinkela_wire_7015)
    );

    bfr new_Jinkela_buffer_1889 (
        .din(new_Jinkela_wire_2810),
        .dout(new_Jinkela_wire_2811)
    );

    and_bi _2035_ (
        .a(new_Jinkela_wire_10573),
        .b(new_Jinkela_wire_11387),
        .c(_1081_)
    );

    bfr new_Jinkela_buffer_1839 (
        .din(new_Jinkela_wire_2754),
        .dout(new_Jinkela_wire_2755)
    );

    and_bb _2036_ (
        .a(new_Jinkela_wire_368),
        .b(new_Jinkela_wire_542),
        .c(_1082_)
    );

    or_ii _2037_ (
        .a(new_Jinkela_wire_327),
        .b(new_Jinkela_wire_490),
        .c(_1083_)
    );

    bfr new_Jinkela_buffer_1840 (
        .din(new_Jinkela_wire_2755),
        .dout(new_Jinkela_wire_2756)
    );

    and_bi _2038_ (
        .a(new_Jinkela_wire_3115),
        .b(new_Jinkela_wire_5432),
        .c(_1084_)
    );

    bfr new_Jinkela_buffer_2014 (
        .din(new_Jinkela_wire_2939),
        .dout(new_Jinkela_wire_2940)
    );

    bfr new_Jinkela_buffer_1890 (
        .din(new_Jinkela_wire_2811),
        .dout(new_Jinkela_wire_2812)
    );

    and_bb _2039_ (
        .a(new_Jinkela_wire_229),
        .b(new_Jinkela_wire_499),
        .c(_1085_)
    );

    bfr new_Jinkela_buffer_1841 (
        .din(new_Jinkela_wire_2756),
        .dout(new_Jinkela_wire_2757)
    );

    and_bi _2040_ (
        .a(new_Jinkela_wire_18110),
        .b(new_Jinkela_wire_17067),
        .c(_1086_)
    );

    and_ii _2041_ (
        .a(new_Jinkela_wire_838),
        .b(new_Jinkela_wire_4298),
        .c(_1087_)
    );

    bfr new_Jinkela_buffer_1842 (
        .din(new_Jinkela_wire_2757),
        .dout(new_Jinkela_wire_2758)
    );

    or_bb _2042_ (
        .a(new_Jinkela_wire_6365),
        .b(new_Jinkela_wire_7708),
        .c(_1088_)
    );

    bfr new_Jinkela_buffer_1908 (
        .din(new_Jinkela_wire_2829),
        .dout(new_Jinkela_wire_2830)
    );

    bfr new_Jinkela_buffer_1891 (
        .din(new_Jinkela_wire_2812),
        .dout(new_Jinkela_wire_2813)
    );

    or_ii _2043_ (
        .a(new_Jinkela_wire_6366),
        .b(new_Jinkela_wire_7709),
        .c(_1089_)
    );

    bfr new_Jinkela_buffer_1843 (
        .din(new_Jinkela_wire_2758),
        .dout(new_Jinkela_wire_2759)
    );

    or_ii _2044_ (
        .a(new_Jinkela_wire_15205),
        .b(new_Jinkela_wire_8282),
        .c(_1090_)
    );

    and_ii _2045_ (
        .a(new_Jinkela_wire_9017),
        .b(new_Jinkela_wire_4471),
        .c(_1091_)
    );

    bfr new_Jinkela_buffer_1844 (
        .din(new_Jinkela_wire_2759),
        .dout(new_Jinkela_wire_2760)
    );

    and_bb _2046_ (
        .a(new_Jinkela_wire_9018),
        .b(new_Jinkela_wire_4472),
        .c(_1092_)
    );

    bfr new_Jinkela_buffer_2016 (
        .din(new_Jinkela_wire_2947),
        .dout(new_Jinkela_wire_2948)
    );

    bfr new_Jinkela_buffer_1892 (
        .din(new_Jinkela_wire_2813),
        .dout(new_Jinkela_wire_2814)
    );

    or_bb _2047_ (
        .a(new_Jinkela_wire_19974),
        .b(new_Jinkela_wire_3890),
        .c(_1093_)
    );

    bfr new_Jinkela_buffer_1845 (
        .din(new_Jinkela_wire_2760),
        .dout(new_Jinkela_wire_2761)
    );

    or_bb _2048_ (
        .a(new_Jinkela_wire_11388),
        .b(new_Jinkela_wire_4720),
        .c(_1094_)
    );

    or_ii _2049_ (
        .a(new_Jinkela_wire_11389),
        .b(new_Jinkela_wire_4721),
        .c(_1095_)
    );

    bfr new_Jinkela_buffer_1846 (
        .din(new_Jinkela_wire_2761),
        .dout(new_Jinkela_wire_2762)
    );

    or_ii _2050_ (
        .a(new_Jinkela_wire_7451),
        .b(new_Jinkela_wire_5098),
        .c(_1096_)
    );

    bfr new_Jinkela_buffer_1909 (
        .din(new_Jinkela_wire_2830),
        .dout(new_Jinkela_wire_2831)
    );

    bfr new_Jinkela_buffer_1893 (
        .din(new_Jinkela_wire_2814),
        .dout(new_Jinkela_wire_2815)
    );

    and_ii _2051_ (
        .a(new_Jinkela_wire_19159),
        .b(new_Jinkela_wire_9539),
        .c(_1097_)
    );

    bfr new_Jinkela_buffer_1847 (
        .din(new_Jinkela_wire_2762),
        .dout(new_Jinkela_wire_2763)
    );

    and_bb _2052_ (
        .a(new_Jinkela_wire_19160),
        .b(new_Jinkela_wire_9540),
        .c(_1098_)
    );

    or_bb _2053_ (
        .a(new_Jinkela_wire_17794),
        .b(new_Jinkela_wire_20142),
        .c(_1099_)
    );

    bfr new_Jinkela_buffer_1848 (
        .din(new_Jinkela_wire_2763),
        .dout(new_Jinkela_wire_2764)
    );

    or_bb _2054_ (
        .a(new_Jinkela_wire_19546),
        .b(new_Jinkela_wire_16212),
        .c(_1100_)
    );

    bfr new_Jinkela_buffer_1894 (
        .din(new_Jinkela_wire_2815),
        .dout(new_Jinkela_wire_2816)
    );

    or_ii _2055_ (
        .a(new_Jinkela_wire_19547),
        .b(new_Jinkela_wire_16213),
        .c(_1101_)
    );

    bfr new_Jinkela_buffer_1849 (
        .din(new_Jinkela_wire_2764),
        .dout(new_Jinkela_wire_2765)
    );

    or_ii _2056_ (
        .a(new_Jinkela_wire_18293),
        .b(new_Jinkela_wire_20333),
        .c(_1102_)
    );

    bfr new_Jinkela_buffer_2021 (
        .din(_0148_),
        .dout(new_Jinkela_wire_2953)
    );

    and_ii _2057_ (
        .a(new_Jinkela_wire_8849),
        .b(new_Jinkela_wire_20651),
        .c(_1103_)
    );

    bfr new_Jinkela_buffer_1850 (
        .din(new_Jinkela_wire_2765),
        .dout(new_Jinkela_wire_2766)
    );

    and_bb _2058_ (
        .a(new_Jinkela_wire_8850),
        .b(new_Jinkela_wire_20652),
        .c(_1104_)
    );

    bfr new_Jinkela_buffer_1910 (
        .din(new_Jinkela_wire_2831),
        .dout(new_Jinkela_wire_2832)
    );

    bfr new_Jinkela_buffer_1895 (
        .din(new_Jinkela_wire_2816),
        .dout(new_Jinkela_wire_2817)
    );

    or_bb _2059_ (
        .a(new_Jinkela_wire_19341),
        .b(new_Jinkela_wire_15662),
        .c(_1105_)
    );

    bfr new_Jinkela_buffer_1851 (
        .din(new_Jinkela_wire_2766),
        .dout(new_Jinkela_wire_2767)
    );

    or_bb _2060_ (
        .a(new_Jinkela_wire_1614),
        .b(new_Jinkela_wire_12337),
        .c(_1106_)
    );

    or_ii _2061_ (
        .a(new_Jinkela_wire_1615),
        .b(new_Jinkela_wire_12338),
        .c(_1107_)
    );

    bfr new_Jinkela_buffer_1852 (
        .din(new_Jinkela_wire_2767),
        .dout(new_Jinkela_wire_2768)
    );

    or_ii _2062_ (
        .a(new_Jinkela_wire_14101),
        .b(new_Jinkela_wire_18785),
        .c(_1108_)
    );

    bfr new_Jinkela_buffer_1896 (
        .din(new_Jinkela_wire_2817),
        .dout(new_Jinkela_wire_2818)
    );

    and_ii _2063_ (
        .a(new_Jinkela_wire_20371),
        .b(new_Jinkela_wire_2455),
        .c(_1109_)
    );

    bfr new_Jinkela_buffer_1853 (
        .din(new_Jinkela_wire_2768),
        .dout(new_Jinkela_wire_2769)
    );

    and_bb _2064_ (
        .a(new_Jinkela_wire_20372),
        .b(new_Jinkela_wire_2456),
        .c(_1110_)
    );

    spl2 new_Jinkela_splitter_315 (
        .a(_0929_),
        .b(new_Jinkela_wire_2954),
        .c(new_Jinkela_wire_2955)
    );

    or_bb _2065_ (
        .a(new_Jinkela_wire_15740),
        .b(new_Jinkela_wire_3271),
        .c(_1111_)
    );

    bfr new_Jinkela_buffer_1854 (
        .din(new_Jinkela_wire_2769),
        .dout(new_Jinkela_wire_2770)
    );

    or_bb _2066_ (
        .a(new_Jinkela_wire_11407),
        .b(new_Jinkela_wire_16949),
        .c(_1112_)
    );

    bfr new_Jinkela_buffer_1911 (
        .din(new_Jinkela_wire_2832),
        .dout(new_Jinkela_wire_2833)
    );

    or_ii _2067_ (
        .a(new_Jinkela_wire_11408),
        .b(new_Jinkela_wire_16950),
        .c(_1113_)
    );

    bfr new_Jinkela_buffer_1855 (
        .din(new_Jinkela_wire_2770),
        .dout(new_Jinkela_wire_2771)
    );

    or_ii _2068_ (
        .a(new_Jinkela_wire_2314),
        .b(new_Jinkela_wire_9550),
        .c(_1114_)
    );

    bfr new_Jinkela_buffer_2017 (
        .din(new_Jinkela_wire_2948),
        .dout(new_Jinkela_wire_2949)
    );

    and_ii _2069_ (
        .a(new_Jinkela_wire_11018),
        .b(new_Jinkela_wire_5326),
        .c(_1115_)
    );

    bfr new_Jinkela_buffer_1856 (
        .din(new_Jinkela_wire_2771),
        .dout(new_Jinkela_wire_2772)
    );

    and_bb _2070_ (
        .a(new_Jinkela_wire_11019),
        .b(new_Jinkela_wire_5327),
        .c(_1116_)
    );

    bfr new_Jinkela_buffer_1912 (
        .din(new_Jinkela_wire_2833),
        .dout(new_Jinkela_wire_2834)
    );

    or_bb _2071_ (
        .a(new_Jinkela_wire_18294),
        .b(new_Jinkela_wire_7584),
        .c(_1117_)
    );

    bfr new_Jinkela_buffer_1857 (
        .din(new_Jinkela_wire_2772),
        .dout(new_Jinkela_wire_2773)
    );

    or_bb _2072_ (
        .a(new_Jinkela_wire_18295),
        .b(new_Jinkela_wire_20260),
        .c(_1118_)
    );

    bfr new_Jinkela_buffer_2022 (
        .din(_1354_),
        .dout(new_Jinkela_wire_2956)
    );

    or_ii _2073_ (
        .a(new_Jinkela_wire_18296),
        .b(new_Jinkela_wire_20261),
        .c(_1119_)
    );

    bfr new_Jinkela_buffer_1858 (
        .din(new_Jinkela_wire_2773),
        .dout(new_Jinkela_wire_2774)
    );

    or_ii _2074_ (
        .a(new_Jinkela_wire_18297),
        .b(new_Jinkela_wire_11448),
        .c(_1120_)
    );

    bfr new_Jinkela_buffer_1913 (
        .din(new_Jinkela_wire_2834),
        .dout(new_Jinkela_wire_2835)
    );

    and_ii _2075_ (
        .a(new_Jinkela_wire_4836),
        .b(new_Jinkela_wire_17421),
        .c(_1121_)
    );

    bfr new_Jinkela_buffer_1859 (
        .din(new_Jinkela_wire_2774),
        .dout(new_Jinkela_wire_2775)
    );

    and_bb _2076_ (
        .a(new_Jinkela_wire_4837),
        .b(new_Jinkela_wire_17422),
        .c(_1122_)
    );

    bfr new_Jinkela_buffer_2018 (
        .din(new_Jinkela_wire_2949),
        .dout(new_Jinkela_wire_2950)
    );

    bfr new_Jinkela_buffer_12417 (
        .din(new_Jinkela_wire_14918),
        .dout(new_Jinkela_wire_14919)
    );

    bfr new_Jinkela_buffer_12333 (
        .din(new_Jinkela_wire_14832),
        .dout(new_Jinkela_wire_14833)
    );

    bfr new_Jinkela_buffer_15800 (
        .din(new_Jinkela_wire_18828),
        .dout(new_Jinkela_wire_18829)
    );

    bfr new_Jinkela_buffer_12500 (
        .din(new_Jinkela_wire_15003),
        .dout(new_Jinkela_wire_15004)
    );

    bfr new_Jinkela_buffer_15812 (
        .din(new_Jinkela_wire_18844),
        .dout(new_Jinkela_wire_18845)
    );

    bfr new_Jinkela_buffer_12334 (
        .din(new_Jinkela_wire_14833),
        .dout(new_Jinkela_wire_14834)
    );

    bfr new_Jinkela_buffer_15801 (
        .din(new_Jinkela_wire_18829),
        .dout(new_Jinkela_wire_18830)
    );

    bfr new_Jinkela_buffer_12418 (
        .din(new_Jinkela_wire_14919),
        .dout(new_Jinkela_wire_14920)
    );

    bfr new_Jinkela_buffer_15910 (
        .din(new_Jinkela_wire_18948),
        .dout(new_Jinkela_wire_18949)
    );

    bfr new_Jinkela_buffer_12335 (
        .din(new_Jinkela_wire_14834),
        .dout(new_Jinkela_wire_14835)
    );

    spl2 new_Jinkela_splitter_1363 (
        .a(new_Jinkela_wire_18830),
        .b(new_Jinkela_wire_18831),
        .c(new_Jinkela_wire_18832)
    );

    bfr new_Jinkela_buffer_12526 (
        .din(new_Jinkela_wire_15033),
        .dout(new_Jinkela_wire_15034)
    );

    spl2 new_Jinkela_splitter_1371 (
        .a(_0220_),
        .b(new_Jinkela_wire_18961),
        .c(new_Jinkela_wire_18962)
    );

    bfr new_Jinkela_buffer_12336 (
        .din(new_Jinkela_wire_14835),
        .dout(new_Jinkela_wire_14836)
    );

    bfr new_Jinkela_buffer_15813 (
        .din(new_Jinkela_wire_18845),
        .dout(new_Jinkela_wire_18846)
    );

    bfr new_Jinkela_buffer_12419 (
        .din(new_Jinkela_wire_14920),
        .dout(new_Jinkela_wire_14921)
    );

    bfr new_Jinkela_buffer_15814 (
        .din(new_Jinkela_wire_18846),
        .dout(new_Jinkela_wire_18847)
    );

    bfr new_Jinkela_buffer_12337 (
        .din(new_Jinkela_wire_14836),
        .dout(new_Jinkela_wire_14837)
    );

    bfr new_Jinkela_buffer_15912 (
        .din(new_Jinkela_wire_18956),
        .dout(new_Jinkela_wire_18957)
    );

    spl2 new_Jinkela_splitter_1372 (
        .a(_1332_),
        .b(new_Jinkela_wire_18963),
        .c(new_Jinkela_wire_18964)
    );

    bfr new_Jinkela_buffer_12501 (
        .din(new_Jinkela_wire_15004),
        .dout(new_Jinkela_wire_15005)
    );

    bfr new_Jinkela_buffer_15815 (
        .din(new_Jinkela_wire_18847),
        .dout(new_Jinkela_wire_18848)
    );

    bfr new_Jinkela_buffer_12338 (
        .din(new_Jinkela_wire_14837),
        .dout(new_Jinkela_wire_14838)
    );

    bfr new_Jinkela_buffer_12420 (
        .din(new_Jinkela_wire_14921),
        .dout(new_Jinkela_wire_14922)
    );

    bfr new_Jinkela_buffer_15816 (
        .din(new_Jinkela_wire_18848),
        .dout(new_Jinkela_wire_18849)
    );

    bfr new_Jinkela_buffer_12339 (
        .din(new_Jinkela_wire_14838),
        .dout(new_Jinkela_wire_14839)
    );

    bfr new_Jinkela_buffer_15913 (
        .din(new_Jinkela_wire_18957),
        .dout(new_Jinkela_wire_18958)
    );

    bfr new_Jinkela_buffer_15817 (
        .din(new_Jinkela_wire_18849),
        .dout(new_Jinkela_wire_18850)
    );

    bfr new_Jinkela_buffer_12682 (
        .din(_0323_),
        .dout(new_Jinkela_wire_15202)
    );

    bfr new_Jinkela_buffer_12340 (
        .din(new_Jinkela_wire_14839),
        .dout(new_Jinkela_wire_14840)
    );

    spl2 new_Jinkela_splitter_1373 (
        .a(_1534_),
        .b(new_Jinkela_wire_18969),
        .c(new_Jinkela_wire_18970)
    );

    bfr new_Jinkela_buffer_12421 (
        .din(new_Jinkela_wire_14922),
        .dout(new_Jinkela_wire_14923)
    );

    bfr new_Jinkela_buffer_15818 (
        .din(new_Jinkela_wire_18850),
        .dout(new_Jinkela_wire_18851)
    );

    bfr new_Jinkela_buffer_12341 (
        .din(new_Jinkela_wire_14840),
        .dout(new_Jinkela_wire_14841)
    );

    bfr new_Jinkela_buffer_15914 (
        .din(new_Jinkela_wire_18958),
        .dout(new_Jinkela_wire_18959)
    );

    bfr new_Jinkela_buffer_12502 (
        .din(new_Jinkela_wire_15005),
        .dout(new_Jinkela_wire_15006)
    );

    bfr new_Jinkela_buffer_15819 (
        .din(new_Jinkela_wire_18851),
        .dout(new_Jinkela_wire_18852)
    );

    bfr new_Jinkela_buffer_12342 (
        .din(new_Jinkela_wire_14841),
        .dout(new_Jinkela_wire_14842)
    );

    bfr new_Jinkela_buffer_15916 (
        .din(new_Jinkela_wire_18964),
        .dout(new_Jinkela_wire_18965)
    );

    spl2 new_Jinkela_splitter_1374 (
        .a(_1590_),
        .b(new_Jinkela_wire_18971),
        .c(new_Jinkela_wire_18972)
    );

    bfr new_Jinkela_buffer_12422 (
        .din(new_Jinkela_wire_14923),
        .dout(new_Jinkela_wire_14924)
    );

    bfr new_Jinkela_buffer_15820 (
        .din(new_Jinkela_wire_18852),
        .dout(new_Jinkela_wire_18853)
    );

    bfr new_Jinkela_buffer_12343 (
        .din(new_Jinkela_wire_14842),
        .dout(new_Jinkela_wire_14843)
    );

    bfr new_Jinkela_buffer_15915 (
        .din(new_Jinkela_wire_18959),
        .dout(new_Jinkela_wire_18960)
    );

    bfr new_Jinkela_buffer_12527 (
        .din(new_Jinkela_wire_15034),
        .dout(new_Jinkela_wire_15035)
    );

    bfr new_Jinkela_buffer_15821 (
        .din(new_Jinkela_wire_18853),
        .dout(new_Jinkela_wire_18854)
    );

    bfr new_Jinkela_buffer_12344 (
        .din(new_Jinkela_wire_14843),
        .dout(new_Jinkela_wire_14844)
    );

    bfr new_Jinkela_buffer_12423 (
        .din(new_Jinkela_wire_14924),
        .dout(new_Jinkela_wire_14925)
    );

    bfr new_Jinkela_buffer_15822 (
        .din(new_Jinkela_wire_18854),
        .dout(new_Jinkela_wire_18855)
    );

    bfr new_Jinkela_buffer_12345 (
        .din(new_Jinkela_wire_14844),
        .dout(new_Jinkela_wire_14845)
    );

    bfr new_Jinkela_buffer_15917 (
        .din(new_Jinkela_wire_18965),
        .dout(new_Jinkela_wire_18966)
    );

    bfr new_Jinkela_buffer_12503 (
        .din(new_Jinkela_wire_15006),
        .dout(new_Jinkela_wire_15007)
    );

    bfr new_Jinkela_buffer_15823 (
        .din(new_Jinkela_wire_18855),
        .dout(new_Jinkela_wire_18856)
    );

    bfr new_Jinkela_buffer_12346 (
        .din(new_Jinkela_wire_14845),
        .dout(new_Jinkela_wire_14846)
    );

    bfr new_Jinkela_buffer_15924 (
        .din(_0629_),
        .dout(new_Jinkela_wire_18981)
    );

    bfr new_Jinkela_buffer_15920 (
        .din(_0119_),
        .dout(new_Jinkela_wire_18973)
    );

    bfr new_Jinkela_buffer_12424 (
        .din(new_Jinkela_wire_14925),
        .dout(new_Jinkela_wire_14926)
    );

    bfr new_Jinkela_buffer_15824 (
        .din(new_Jinkela_wire_18856),
        .dout(new_Jinkela_wire_18857)
    );

    bfr new_Jinkela_buffer_12347 (
        .din(new_Jinkela_wire_14846),
        .dout(new_Jinkela_wire_14847)
    );

    bfr new_Jinkela_buffer_15918 (
        .din(new_Jinkela_wire_18966),
        .dout(new_Jinkela_wire_18967)
    );

    bfr new_Jinkela_buffer_12611 (
        .din(new_Jinkela_wire_15126),
        .dout(new_Jinkela_wire_15127)
    );

    bfr new_Jinkela_buffer_15825 (
        .din(new_Jinkela_wire_18857),
        .dout(new_Jinkela_wire_18858)
    );

    bfr new_Jinkela_buffer_12348 (
        .din(new_Jinkela_wire_14847),
        .dout(new_Jinkela_wire_14848)
    );

    spl2 new_Jinkela_splitter_1376 (
        .a(_1685_),
        .b(new_Jinkela_wire_18979),
        .c(new_Jinkela_wire_18980)
    );

    bfr new_Jinkela_buffer_12425 (
        .din(new_Jinkela_wire_14926),
        .dout(new_Jinkela_wire_14927)
    );

    bfr new_Jinkela_buffer_15826 (
        .din(new_Jinkela_wire_18858),
        .dout(new_Jinkela_wire_18859)
    );

    bfr new_Jinkela_buffer_12349 (
        .din(new_Jinkela_wire_14848),
        .dout(new_Jinkela_wire_14849)
    );

    bfr new_Jinkela_buffer_15919 (
        .din(new_Jinkela_wire_18967),
        .dout(new_Jinkela_wire_18968)
    );

    bfr new_Jinkela_buffer_12504 (
        .din(new_Jinkela_wire_15007),
        .dout(new_Jinkela_wire_15008)
    );

    bfr new_Jinkela_buffer_15827 (
        .din(new_Jinkela_wire_18859),
        .dout(new_Jinkela_wire_18860)
    );

    bfr new_Jinkela_buffer_12350 (
        .din(new_Jinkela_wire_14849),
        .dout(new_Jinkela_wire_14850)
    );

    bfr new_Jinkela_buffer_15921 (
        .din(new_Jinkela_wire_18973),
        .dout(new_Jinkela_wire_18974)
    );

    bfr new_Jinkela_buffer_12426 (
        .din(new_Jinkela_wire_14927),
        .dout(new_Jinkela_wire_14928)
    );

    bfr new_Jinkela_buffer_15828 (
        .din(new_Jinkela_wire_18860),
        .dout(new_Jinkela_wire_18861)
    );

    bfr new_Jinkela_buffer_12351 (
        .din(new_Jinkela_wire_14850),
        .dout(new_Jinkela_wire_14851)
    );

    bfr new_Jinkela_buffer_15986 (
        .din(_0174_),
        .dout(new_Jinkela_wire_19047)
    );

    bfr new_Jinkela_buffer_15922 (
        .din(new_Jinkela_wire_18974),
        .dout(new_Jinkela_wire_18975)
    );

    bfr new_Jinkela_buffer_12528 (
        .din(new_Jinkela_wire_15035),
        .dout(new_Jinkela_wire_15036)
    );

    bfr new_Jinkela_buffer_15829 (
        .din(new_Jinkela_wire_18861),
        .dout(new_Jinkela_wire_18862)
    );

    bfr new_Jinkela_buffer_12352 (
        .din(new_Jinkela_wire_14851),
        .dout(new_Jinkela_wire_14852)
    );

    bfr new_Jinkela_buffer_12427 (
        .din(new_Jinkela_wire_14928),
        .dout(new_Jinkela_wire_14929)
    );

    bfr new_Jinkela_buffer_15830 (
        .din(new_Jinkela_wire_18862),
        .dout(new_Jinkela_wire_18863)
    );

    bfr new_Jinkela_buffer_12353 (
        .din(new_Jinkela_wire_14852),
        .dout(new_Jinkela_wire_14853)
    );

    spl2 new_Jinkela_splitter_1378 (
        .a(_1816_),
        .b(new_Jinkela_wire_19045),
        .c(new_Jinkela_wire_19046)
    );

    bfr new_Jinkela_buffer_8895 (
        .din(new_Jinkela_wire_10886),
        .dout(new_Jinkela_wire_10887)
    );

    bfr new_Jinkela_buffer_5407 (
        .din(new_Jinkela_wire_6934),
        .dout(new_Jinkela_wire_6935)
    );

    bfr new_Jinkela_buffer_8985 (
        .din(new_Jinkela_wire_10990),
        .dout(new_Jinkela_wire_10991)
    );

    bfr new_Jinkela_buffer_5591 (
        .din(new_Jinkela_wire_7134),
        .dout(new_Jinkela_wire_7135)
    );

    bfr new_Jinkela_buffer_8896 (
        .din(new_Jinkela_wire_10887),
        .dout(new_Jinkela_wire_10888)
    );

    bfr new_Jinkela_buffer_5408 (
        .din(new_Jinkela_wire_6935),
        .dout(new_Jinkela_wire_6936)
    );

    bfr new_Jinkela_buffer_9031 (
        .din(new_Jinkela_wire_11042),
        .dout(new_Jinkela_wire_11043)
    );

    bfr new_Jinkela_buffer_5480 (
        .din(new_Jinkela_wire_7015),
        .dout(new_Jinkela_wire_7016)
    );

    bfr new_Jinkela_buffer_8897 (
        .din(new_Jinkela_wire_10888),
        .dout(new_Jinkela_wire_10889)
    );

    bfr new_Jinkela_buffer_5409 (
        .din(new_Jinkela_wire_6936),
        .dout(new_Jinkela_wire_6937)
    );

    bfr new_Jinkela_buffer_8986 (
        .din(new_Jinkela_wire_10991),
        .dout(new_Jinkela_wire_10992)
    );

    bfr new_Jinkela_buffer_5526 (
        .din(new_Jinkela_wire_7063),
        .dout(new_Jinkela_wire_7064)
    );

    bfr new_Jinkela_buffer_8898 (
        .din(new_Jinkela_wire_10889),
        .dout(new_Jinkela_wire_10890)
    );

    bfr new_Jinkela_buffer_5410 (
        .din(new_Jinkela_wire_6937),
        .dout(new_Jinkela_wire_6938)
    );

    bfr new_Jinkela_buffer_9019 (
        .din(new_Jinkela_wire_11028),
        .dout(new_Jinkela_wire_11029)
    );

    bfr new_Jinkela_buffer_5481 (
        .din(new_Jinkela_wire_7016),
        .dout(new_Jinkela_wire_7017)
    );

    bfr new_Jinkela_buffer_8899 (
        .din(new_Jinkela_wire_10890),
        .dout(new_Jinkela_wire_10891)
    );

    bfr new_Jinkela_buffer_5411 (
        .din(new_Jinkela_wire_6938),
        .dout(new_Jinkela_wire_6939)
    );

    bfr new_Jinkela_buffer_8987 (
        .din(new_Jinkela_wire_10992),
        .dout(new_Jinkela_wire_10993)
    );

    bfr new_Jinkela_buffer_5593 (
        .din(new_Jinkela_wire_7138),
        .dout(new_Jinkela_wire_7139)
    );

    bfr new_Jinkela_buffer_8900 (
        .din(new_Jinkela_wire_10891),
        .dout(new_Jinkela_wire_10892)
    );

    bfr new_Jinkela_buffer_5412 (
        .din(new_Jinkela_wire_6939),
        .dout(new_Jinkela_wire_6940)
    );

    bfr new_Jinkela_buffer_9033 (
        .din(new_Jinkela_wire_11048),
        .dout(new_Jinkela_wire_11049)
    );

    bfr new_Jinkela_buffer_5482 (
        .din(new_Jinkela_wire_7017),
        .dout(new_Jinkela_wire_7018)
    );

    bfr new_Jinkela_buffer_8901 (
        .din(new_Jinkela_wire_10892),
        .dout(new_Jinkela_wire_10893)
    );

    bfr new_Jinkela_buffer_5413 (
        .din(new_Jinkela_wire_6940),
        .dout(new_Jinkela_wire_6941)
    );

    bfr new_Jinkela_buffer_8988 (
        .din(new_Jinkela_wire_10993),
        .dout(new_Jinkela_wire_10994)
    );

    bfr new_Jinkela_buffer_5527 (
        .din(new_Jinkela_wire_7064),
        .dout(new_Jinkela_wire_7065)
    );

    bfr new_Jinkela_buffer_8902 (
        .din(new_Jinkela_wire_10893),
        .dout(new_Jinkela_wire_10894)
    );

    bfr new_Jinkela_buffer_5414 (
        .din(new_Jinkela_wire_6941),
        .dout(new_Jinkela_wire_6942)
    );

    bfr new_Jinkela_buffer_9020 (
        .din(new_Jinkela_wire_11029),
        .dout(new_Jinkela_wire_11030)
    );

    bfr new_Jinkela_buffer_5483 (
        .din(new_Jinkela_wire_7018),
        .dout(new_Jinkela_wire_7019)
    );

    bfr new_Jinkela_buffer_8903 (
        .din(new_Jinkela_wire_10894),
        .dout(new_Jinkela_wire_10895)
    );

    bfr new_Jinkela_buffer_5415 (
        .din(new_Jinkela_wire_6942),
        .dout(new_Jinkela_wire_6943)
    );

    bfr new_Jinkela_buffer_8989 (
        .din(new_Jinkela_wire_10994),
        .dout(new_Jinkela_wire_10995)
    );

    bfr new_Jinkela_buffer_5597 (
        .din(new_Jinkela_wire_7142),
        .dout(new_Jinkela_wire_7143)
    );

    bfr new_Jinkela_buffer_8904 (
        .din(new_Jinkela_wire_10895),
        .dout(new_Jinkela_wire_10896)
    );

    bfr new_Jinkela_buffer_5416 (
        .din(new_Jinkela_wire_6943),
        .dout(new_Jinkela_wire_6944)
    );

    spl2 new_Jinkela_splitter_855 (
        .a(new_Jinkela_wire_11043),
        .b(new_Jinkela_wire_11044),
        .c(new_Jinkela_wire_11045)
    );

    bfr new_Jinkela_buffer_5484 (
        .din(new_Jinkela_wire_7019),
        .dout(new_Jinkela_wire_7020)
    );

    bfr new_Jinkela_buffer_8905 (
        .din(new_Jinkela_wire_10896),
        .dout(new_Jinkela_wire_10897)
    );

    bfr new_Jinkela_buffer_5417 (
        .din(new_Jinkela_wire_6944),
        .dout(new_Jinkela_wire_6945)
    );

    bfr new_Jinkela_buffer_8990 (
        .din(new_Jinkela_wire_10995),
        .dout(new_Jinkela_wire_10996)
    );

    bfr new_Jinkela_buffer_5528 (
        .din(new_Jinkela_wire_7065),
        .dout(new_Jinkela_wire_7066)
    );

    bfr new_Jinkela_buffer_8906 (
        .din(new_Jinkela_wire_10897),
        .dout(new_Jinkela_wire_10898)
    );

    bfr new_Jinkela_buffer_5418 (
        .din(new_Jinkela_wire_6945),
        .dout(new_Jinkela_wire_6946)
    );

    bfr new_Jinkela_buffer_9021 (
        .din(new_Jinkela_wire_11030),
        .dout(new_Jinkela_wire_11031)
    );

    bfr new_Jinkela_buffer_5485 (
        .din(new_Jinkela_wire_7020),
        .dout(new_Jinkela_wire_7021)
    );

    bfr new_Jinkela_buffer_8907 (
        .din(new_Jinkela_wire_10898),
        .dout(new_Jinkela_wire_10899)
    );

    bfr new_Jinkela_buffer_5419 (
        .din(new_Jinkela_wire_6946),
        .dout(new_Jinkela_wire_6947)
    );

    bfr new_Jinkela_buffer_8991 (
        .din(new_Jinkela_wire_10996),
        .dout(new_Jinkela_wire_10997)
    );

    bfr new_Jinkela_buffer_5594 (
        .din(new_Jinkela_wire_7139),
        .dout(new_Jinkela_wire_7140)
    );

    bfr new_Jinkela_buffer_8908 (
        .din(new_Jinkela_wire_10899),
        .dout(new_Jinkela_wire_10900)
    );

    bfr new_Jinkela_buffer_5420 (
        .din(new_Jinkela_wire_6947),
        .dout(new_Jinkela_wire_6948)
    );

    bfr new_Jinkela_buffer_9034 (
        .din(new_Jinkela_wire_11049),
        .dout(new_Jinkela_wire_11050)
    );

    bfr new_Jinkela_buffer_5486 (
        .din(new_Jinkela_wire_7021),
        .dout(new_Jinkela_wire_7022)
    );

    bfr new_Jinkela_buffer_8909 (
        .din(new_Jinkela_wire_10900),
        .dout(new_Jinkela_wire_10901)
    );

    bfr new_Jinkela_buffer_5421 (
        .din(new_Jinkela_wire_6948),
        .dout(new_Jinkela_wire_6949)
    );

    bfr new_Jinkela_buffer_8992 (
        .din(new_Jinkela_wire_10997),
        .dout(new_Jinkela_wire_10998)
    );

    bfr new_Jinkela_buffer_5529 (
        .din(new_Jinkela_wire_7066),
        .dout(new_Jinkela_wire_7067)
    );

    bfr new_Jinkela_buffer_8910 (
        .din(new_Jinkela_wire_10901),
        .dout(new_Jinkela_wire_10902)
    );

    bfr new_Jinkela_buffer_5422 (
        .din(new_Jinkela_wire_6949),
        .dout(new_Jinkela_wire_6950)
    );

    bfr new_Jinkela_buffer_9022 (
        .din(new_Jinkela_wire_11031),
        .dout(new_Jinkela_wire_11032)
    );

    bfr new_Jinkela_buffer_5487 (
        .din(new_Jinkela_wire_7022),
        .dout(new_Jinkela_wire_7023)
    );

    bfr new_Jinkela_buffer_8911 (
        .din(new_Jinkela_wire_10902),
        .dout(new_Jinkela_wire_10903)
    );

    bfr new_Jinkela_buffer_5423 (
        .din(new_Jinkela_wire_6950),
        .dout(new_Jinkela_wire_6951)
    );

    bfr new_Jinkela_buffer_8993 (
        .din(new_Jinkela_wire_10998),
        .dout(new_Jinkela_wire_10999)
    );

    spl2 new_Jinkela_splitter_624 (
        .a(_1803_),
        .b(new_Jinkela_wire_7182),
        .c(new_Jinkela_wire_7183)
    );

    spl2 new_Jinkela_splitter_623 (
        .a(_0794_),
        .b(new_Jinkela_wire_7176),
        .c(new_Jinkela_wire_7177)
    );

    bfr new_Jinkela_buffer_8912 (
        .din(new_Jinkela_wire_10903),
        .dout(new_Jinkela_wire_10904)
    );

    bfr new_Jinkela_buffer_5424 (
        .din(new_Jinkela_wire_6951),
        .dout(new_Jinkela_wire_6952)
    );

    bfr new_Jinkela_buffer_9118 (
        .din(_1564_),
        .dout(new_Jinkela_wire_11138)
    );

    bfr new_Jinkela_buffer_5488 (
        .din(new_Jinkela_wire_7023),
        .dout(new_Jinkela_wire_7024)
    );

    spl2 new_Jinkela_splitter_858 (
        .a(_0433_),
        .b(new_Jinkela_wire_11136),
        .c(new_Jinkela_wire_11137)
    );

    bfr new_Jinkela_buffer_8913 (
        .din(new_Jinkela_wire_10904),
        .dout(new_Jinkela_wire_10905)
    );

    bfr new_Jinkela_buffer_5425 (
        .din(new_Jinkela_wire_6952),
        .dout(new_Jinkela_wire_6953)
    );

    bfr new_Jinkela_buffer_8994 (
        .din(new_Jinkela_wire_10999),
        .dout(new_Jinkela_wire_11000)
    );

    bfr new_Jinkela_buffer_5530 (
        .din(new_Jinkela_wire_7067),
        .dout(new_Jinkela_wire_7068)
    );

    bfr new_Jinkela_buffer_8914 (
        .din(new_Jinkela_wire_10905),
        .dout(new_Jinkela_wire_10906)
    );

    bfr new_Jinkela_buffer_5426 (
        .din(new_Jinkela_wire_6953),
        .dout(new_Jinkela_wire_6954)
    );

    bfr new_Jinkela_buffer_9023 (
        .din(new_Jinkela_wire_11032),
        .dout(new_Jinkela_wire_11033)
    );

    bfr new_Jinkela_buffer_5489 (
        .din(new_Jinkela_wire_7024),
        .dout(new_Jinkela_wire_7025)
    );

    bfr new_Jinkela_buffer_8915 (
        .din(new_Jinkela_wire_10906),
        .dout(new_Jinkela_wire_10907)
    );

    bfr new_Jinkela_buffer_5427 (
        .din(new_Jinkela_wire_6954),
        .dout(new_Jinkela_wire_6955)
    );

    bfr new_Jinkela_buffer_8995 (
        .din(new_Jinkela_wire_11000),
        .dout(new_Jinkela_wire_11001)
    );

    bfr new_Jinkela_buffer_5595 (
        .din(new_Jinkela_wire_7140),
        .dout(new_Jinkela_wire_7141)
    );

    bfr new_Jinkela_buffer_12505 (
        .din(new_Jinkela_wire_15008),
        .dout(new_Jinkela_wire_15009)
    );

    and_ii _2959_ (
        .a(new_Jinkela_wire_7262),
        .b(new_Jinkela_wire_7308),
        .c(_0205_)
    );

    bfr new_Jinkela_buffer_1860 (
        .din(new_Jinkela_wire_2775),
        .dout(new_Jinkela_wire_2776)
    );

    bfr new_Jinkela_buffer_12354 (
        .din(new_Jinkela_wire_14853),
        .dout(new_Jinkela_wire_14854)
    );

    or_bb _2960_ (
        .a(new_Jinkela_wire_9742),
        .b(new_Jinkela_wire_20285),
        .c(_0206_)
    );

    bfr new_Jinkela_buffer_1914 (
        .din(new_Jinkela_wire_2835),
        .dout(new_Jinkela_wire_2836)
    );

    bfr new_Jinkela_buffer_12428 (
        .din(new_Jinkela_wire_14929),
        .dout(new_Jinkela_wire_14930)
    );

    and_bi _2961_ (
        .a(new_Jinkela_wire_4162),
        .b(new_Jinkela_wire_5052),
        .c(_0207_)
    );

    bfr new_Jinkela_buffer_1861 (
        .din(new_Jinkela_wire_2776),
        .dout(new_Jinkela_wire_2777)
    );

    bfr new_Jinkela_buffer_12355 (
        .din(new_Jinkela_wire_14854),
        .dout(new_Jinkela_wire_14855)
    );

    and_bi _2962_ (
        .a(new_Jinkela_wire_5053),
        .b(new_Jinkela_wire_4163),
        .c(_0208_)
    );

    spl2 new_Jinkela_splitter_316 (
        .a(_0830_),
        .b(new_Jinkela_wire_2958),
        .c(new_Jinkela_wire_2959)
    );

    bfr new_Jinkela_buffer_12683 (
        .din(_1089_),
        .dout(new_Jinkela_wire_15205)
    );

    or_bb _2963_ (
        .a(new_Jinkela_wire_12724),
        .b(new_Jinkela_wire_16121),
        .c(new_net_3936)
    );

    bfr new_Jinkela_buffer_1862 (
        .din(new_Jinkela_wire_2777),
        .dout(new_Jinkela_wire_2778)
    );

    bfr new_Jinkela_buffer_12356 (
        .din(new_Jinkela_wire_14855),
        .dout(new_Jinkela_wire_14856)
    );

    or_bb _2964_ (
        .a(new_Jinkela_wire_16122),
        .b(new_Jinkela_wire_20810),
        .c(_0210_)
    );

    bfr new_Jinkela_buffer_1915 (
        .din(new_Jinkela_wire_2836),
        .dout(new_Jinkela_wire_2837)
    );

    bfr new_Jinkela_buffer_12429 (
        .din(new_Jinkela_wire_14930),
        .dout(new_Jinkela_wire_14931)
    );

    and_bi _2965_ (
        .a(new_Jinkela_wire_19565),
        .b(new_Jinkela_wire_7713),
        .c(_0211_)
    );

    bfr new_Jinkela_buffer_1863 (
        .din(new_Jinkela_wire_2778),
        .dout(new_Jinkela_wire_2779)
    );

    bfr new_Jinkela_buffer_12357 (
        .din(new_Jinkela_wire_14856),
        .dout(new_Jinkela_wire_14857)
    );

    and_bb _2966_ (
        .a(new_Jinkela_wire_273),
        .b(new_Jinkela_wire_678),
        .c(_0212_)
    );

    bfr new_Jinkela_buffer_2019 (
        .din(new_Jinkela_wire_2950),
        .dout(new_Jinkela_wire_2951)
    );

    bfr new_Jinkela_buffer_12506 (
        .din(new_Jinkela_wire_15009),
        .dout(new_Jinkela_wire_15010)
    );

    and_bi _2967_ (
        .a(new_Jinkela_wire_13592),
        .b(new_Jinkela_wire_8765),
        .c(_0213_)
    );

    bfr new_Jinkela_buffer_1864 (
        .din(new_Jinkela_wire_2779),
        .dout(new_Jinkela_wire_2780)
    );

    bfr new_Jinkela_buffer_12358 (
        .din(new_Jinkela_wire_14857),
        .dout(new_Jinkela_wire_14858)
    );

    and_bb _2968_ (
        .a(new_Jinkela_wire_74),
        .b(new_Jinkela_wire_508),
        .c(_0214_)
    );

    bfr new_Jinkela_buffer_1916 (
        .din(new_Jinkela_wire_2837),
        .dout(new_Jinkela_wire_2838)
    );

    bfr new_Jinkela_buffer_12430 (
        .din(new_Jinkela_wire_14931),
        .dout(new_Jinkela_wire_14932)
    );

    and_bi _2969_ (
        .a(new_Jinkela_wire_3252),
        .b(new_Jinkela_wire_1617),
        .c(_0215_)
    );

    bfr new_Jinkela_buffer_1865 (
        .din(new_Jinkela_wire_2780),
        .dout(new_Jinkela_wire_2781)
    );

    bfr new_Jinkela_buffer_12359 (
        .din(new_Jinkela_wire_14858),
        .dout(new_Jinkela_wire_14859)
    );

    and_bb _2970_ (
        .a(new_Jinkela_wire_469),
        .b(new_Jinkela_wire_139),
        .c(_0216_)
    );

    bfr new_Jinkela_buffer_2023 (
        .din(_1640_),
        .dout(new_Jinkela_wire_2957)
    );

    bfr new_Jinkela_buffer_12529 (
        .din(new_Jinkela_wire_15036),
        .dout(new_Jinkela_wire_15037)
    );

    and_bi _2971_ (
        .a(new_Jinkela_wire_6006),
        .b(new_Jinkela_wire_9174),
        .c(_0217_)
    );

    bfr new_Jinkela_buffer_1866 (
        .din(new_Jinkela_wire_2781),
        .dout(new_Jinkela_wire_2782)
    );

    bfr new_Jinkela_buffer_12360 (
        .din(new_Jinkela_wire_14859),
        .dout(new_Jinkela_wire_14860)
    );

    and_bb _2972_ (
        .a(new_Jinkela_wire_364),
        .b(new_Jinkela_wire_206),
        .c(_0218_)
    );

    bfr new_Jinkela_buffer_1917 (
        .din(new_Jinkela_wire_2838),
        .dout(new_Jinkela_wire_2839)
    );

    bfr new_Jinkela_buffer_12431 (
        .din(new_Jinkela_wire_14932),
        .dout(new_Jinkela_wire_14933)
    );

    and_bi _2973_ (
        .a(new_Jinkela_wire_1607),
        .b(new_Jinkela_wire_3668),
        .c(_0220_)
    );

    bfr new_Jinkela_buffer_1867 (
        .din(new_Jinkela_wire_2782),
        .dout(new_Jinkela_wire_2783)
    );

    bfr new_Jinkela_buffer_12361 (
        .din(new_Jinkela_wire_14860),
        .dout(new_Jinkela_wire_14861)
    );

    and_bb _2974_ (
        .a(new_Jinkela_wire_686),
        .b(new_Jinkela_wire_580),
        .c(_0221_)
    );

    spl2 new_Jinkela_splitter_317 (
        .a(_0511_),
        .b(new_Jinkela_wire_2960),
        .c(new_Jinkela_wire_2961)
    );

    bfr new_Jinkela_buffer_12507 (
        .din(new_Jinkela_wire_15010),
        .dout(new_Jinkela_wire_15011)
    );

    and_bi _2975_ (
        .a(new_Jinkela_wire_10567),
        .b(new_Jinkela_wire_12628),
        .c(_0222_)
    );

    bfr new_Jinkela_buffer_1868 (
        .din(new_Jinkela_wire_2783),
        .dout(new_Jinkela_wire_2784)
    );

    bfr new_Jinkela_buffer_12362 (
        .din(new_Jinkela_wire_14861),
        .dout(new_Jinkela_wire_14862)
    );

    and_bb _2976_ (
        .a(new_Jinkela_wire_116),
        .b(new_Jinkela_wire_496),
        .c(_0223_)
    );

    bfr new_Jinkela_buffer_1918 (
        .din(new_Jinkela_wire_2839),
        .dout(new_Jinkela_wire_2840)
    );

    bfr new_Jinkela_buffer_12432 (
        .din(new_Jinkela_wire_14933),
        .dout(new_Jinkela_wire_14934)
    );

    and_bi _2977_ (
        .a(new_Jinkela_wire_18707),
        .b(new_Jinkela_wire_15698),
        .c(_0224_)
    );

    spl2 new_Jinkela_splitter_307 (
        .a(new_Jinkela_wire_2784),
        .b(new_Jinkela_wire_2785),
        .c(new_Jinkela_wire_2786)
    );

    bfr new_Jinkela_buffer_12363 (
        .din(new_Jinkela_wire_14862),
        .dout(new_Jinkela_wire_14863)
    );

    and_bb _2978_ (
        .a(new_Jinkela_wire_42),
        .b(new_Jinkela_wire_15),
        .c(_0225_)
    );

    bfr new_Jinkela_buffer_1919 (
        .din(new_Jinkela_wire_2840),
        .dout(new_Jinkela_wire_2841)
    );

    bfr new_Jinkela_buffer_12612 (
        .din(new_Jinkela_wire_15127),
        .dout(new_Jinkela_wire_15128)
    );

    and_bi _2979_ (
        .a(new_Jinkela_wire_1274),
        .b(new_Jinkela_wire_7271),
        .c(_0226_)
    );

    bfr new_Jinkela_buffer_12364 (
        .din(new_Jinkela_wire_14863),
        .dout(new_Jinkela_wire_14864)
    );

    and_bb _2980_ (
        .a(new_Jinkela_wire_196),
        .b(new_Jinkela_wire_447),
        .c(_0227_)
    );

    spl2 new_Jinkela_splitter_318 (
        .a(_0350_),
        .b(new_Jinkela_wire_2962),
        .c(new_Jinkela_wire_2963)
    );

    bfr new_Jinkela_buffer_12433 (
        .din(new_Jinkela_wire_14934),
        .dout(new_Jinkela_wire_14935)
    );

    and_bi _2981_ (
        .a(new_Jinkela_wire_2256),
        .b(new_Jinkela_wire_11826),
        .c(_0228_)
    );

    bfr new_Jinkela_buffer_1920 (
        .din(new_Jinkela_wire_2841),
        .dout(new_Jinkela_wire_2842)
    );

    bfr new_Jinkela_buffer_12365 (
        .din(new_Jinkela_wire_14864),
        .dout(new_Jinkela_wire_14865)
    );

    and_bb _2982_ (
        .a(new_Jinkela_wire_374),
        .b(new_Jinkela_wire_248),
        .c(_0229_)
    );

    spl2 new_Jinkela_splitter_319 (
        .a(_0748_),
        .b(new_Jinkela_wire_2964),
        .c(new_Jinkela_wire_2965)
    );

    bfr new_Jinkela_buffer_12508 (
        .din(new_Jinkela_wire_15011),
        .dout(new_Jinkela_wire_15012)
    );

    and_bi _2983_ (
        .a(new_Jinkela_wire_7725),
        .b(new_Jinkela_wire_1780),
        .c(_0231_)
    );

    bfr new_Jinkela_buffer_1921 (
        .din(new_Jinkela_wire_2842),
        .dout(new_Jinkela_wire_2843)
    );

    bfr new_Jinkela_buffer_12366 (
        .din(new_Jinkela_wire_14865),
        .dout(new_Jinkela_wire_14866)
    );

    and_bb _2984_ (
        .a(new_Jinkela_wire_405),
        .b(new_Jinkela_wire_304),
        .c(_0232_)
    );

    bfr new_Jinkela_buffer_2025 (
        .din(new_Jinkela_wire_2966),
        .dout(new_Jinkela_wire_2967)
    );

    bfr new_Jinkela_buffer_2024 (
        .din(new_net_3974),
        .dout(new_Jinkela_wire_2966)
    );

    bfr new_Jinkela_buffer_12434 (
        .din(new_Jinkela_wire_14935),
        .dout(new_Jinkela_wire_14936)
    );

    and_bi _2985_ (
        .a(new_Jinkela_wire_13965),
        .b(new_Jinkela_wire_21107),
        .c(_0233_)
    );

    bfr new_Jinkela_buffer_1922 (
        .din(new_Jinkela_wire_2843),
        .dout(new_Jinkela_wire_2844)
    );

    bfr new_Jinkela_buffer_12367 (
        .din(new_Jinkela_wire_14866),
        .dout(new_Jinkela_wire_14867)
    );

    and_bb _2986_ (
        .a(new_Jinkela_wire_159),
        .b(new_Jinkela_wire_50),
        .c(_0234_)
    );

    spl2 new_Jinkela_splitter_321 (
        .a(_1690_),
        .b(new_Jinkela_wire_3116),
        .c(new_Jinkela_wire_3117)
    );

    spl2 new_Jinkela_splitter_320 (
        .a(_1033_),
        .b(new_Jinkela_wire_3114),
        .c(new_Jinkela_wire_3115)
    );

    bfr new_Jinkela_buffer_12530 (
        .din(new_Jinkela_wire_15037),
        .dout(new_Jinkela_wire_15038)
    );

    and_bi _2987_ (
        .a(new_Jinkela_wire_17078),
        .b(new_Jinkela_wire_7743),
        .c(_0235_)
    );

    bfr new_Jinkela_buffer_1923 (
        .din(new_Jinkela_wire_2844),
        .dout(new_Jinkela_wire_2845)
    );

    bfr new_Jinkela_buffer_12368 (
        .din(new_Jinkela_wire_14867),
        .dout(new_Jinkela_wire_14868)
    );

    and_bb _2988_ (
        .a(new_Jinkela_wire_612),
        .b(new_Jinkela_wire_658),
        .c(_0236_)
    );

    bfr new_Jinkela_buffer_12435 (
        .din(new_Jinkela_wire_14936),
        .dout(new_Jinkela_wire_14937)
    );

    and_bb _2989_ (
        .a(new_Jinkela_wire_426),
        .b(new_Jinkela_wire_620),
        .c(_0237_)
    );

    bfr new_Jinkela_buffer_1924 (
        .din(new_Jinkela_wire_2845),
        .dout(new_Jinkela_wire_2846)
    );

    bfr new_Jinkela_buffer_12369 (
        .din(new_Jinkela_wire_14868),
        .dout(new_Jinkela_wire_14869)
    );

    and_ii _2990_ (
        .a(new_Jinkela_wire_5805),
        .b(new_Jinkela_wire_13409),
        .c(_0238_)
    );

    bfr new_Jinkela_buffer_2026 (
        .din(new_Jinkela_wire_2967),
        .dout(new_Jinkela_wire_2968)
    );

    bfr new_Jinkela_buffer_12509 (
        .din(new_Jinkela_wire_15012),
        .dout(new_Jinkela_wire_15013)
    );

    and_ii _2991_ (
        .a(new_Jinkela_wire_13580),
        .b(new_Jinkela_wire_2479),
        .c(_0239_)
    );

    bfr new_Jinkela_buffer_1925 (
        .din(new_Jinkela_wire_2846),
        .dout(new_Jinkela_wire_2847)
    );

    bfr new_Jinkela_buffer_12370 (
        .din(new_Jinkela_wire_14869),
        .dout(new_Jinkela_wire_14870)
    );

    and_bb _2992_ (
        .a(new_Jinkela_wire_13581),
        .b(new_Jinkela_wire_2480),
        .c(_0240_)
    );

    bfr new_Jinkela_buffer_12436 (
        .din(new_Jinkela_wire_14937),
        .dout(new_Jinkela_wire_14938)
    );

    or_bb _2993_ (
        .a(new_Jinkela_wire_13456),
        .b(new_Jinkela_wire_10745),
        .c(_0242_)
    );

    bfr new_Jinkela_buffer_1926 (
        .din(new_Jinkela_wire_2847),
        .dout(new_Jinkela_wire_2848)
    );

    bfr new_Jinkela_buffer_12371 (
        .din(new_Jinkela_wire_14870),
        .dout(new_Jinkela_wire_14871)
    );

    and_ii _2994_ (
        .a(new_Jinkela_wire_8288),
        .b(new_Jinkela_wire_19316),
        .c(_0243_)
    );

    bfr new_Jinkela_buffer_2027 (
        .din(new_Jinkela_wire_2968),
        .dout(new_Jinkela_wire_2969)
    );

    and_bb _2995_ (
        .a(new_Jinkela_wire_8289),
        .b(new_Jinkela_wire_19317),
        .c(_0244_)
    );

    bfr new_Jinkela_buffer_1927 (
        .din(new_Jinkela_wire_2848),
        .dout(new_Jinkela_wire_2849)
    );

    spl2 new_Jinkela_splitter_1109 (
        .a(_1168_),
        .b(new_Jinkela_wire_15203),
        .c(new_Jinkela_wire_15204)
    );

    bfr new_Jinkela_buffer_12372 (
        .din(new_Jinkela_wire_14871),
        .dout(new_Jinkela_wire_14872)
    );

    or_bb _2996_ (
        .a(new_Jinkela_wire_12062),
        .b(new_Jinkela_wire_8586),
        .c(_0245_)
    );

    spl2 new_Jinkela_splitter_322 (
        .a(_0265_),
        .b(new_Jinkela_wire_3118),
        .c(new_Jinkela_wire_3119)
    );

    bfr new_Jinkela_buffer_12437 (
        .din(new_Jinkela_wire_14938),
        .dout(new_Jinkela_wire_14939)
    );

    and_ii _2997_ (
        .a(new_Jinkela_wire_2659),
        .b(new_Jinkela_wire_5443),
        .c(_0246_)
    );

    bfr new_Jinkela_buffer_1928 (
        .din(new_Jinkela_wire_2849),
        .dout(new_Jinkela_wire_2850)
    );

    bfr new_Jinkela_buffer_12373 (
        .din(new_Jinkela_wire_14872),
        .dout(new_Jinkela_wire_14873)
    );

    and_bb _2998_ (
        .a(new_Jinkela_wire_2660),
        .b(new_Jinkela_wire_5444),
        .c(_0247_)
    );

    spl2 new_Jinkela_splitter_323 (
        .a(_0885_),
        .b(new_Jinkela_wire_3120),
        .c(new_Jinkela_wire_3121)
    );

    bfr new_Jinkela_buffer_2028 (
        .din(new_Jinkela_wire_2969),
        .dout(new_Jinkela_wire_2970)
    );

    bfr new_Jinkela_buffer_12510 (
        .din(new_Jinkela_wire_15013),
        .dout(new_Jinkela_wire_15014)
    );

    or_bb _2999_ (
        .a(new_Jinkela_wire_16873),
        .b(new_Jinkela_wire_2935),
        .c(_0248_)
    );

    bfr new_Jinkela_buffer_1929 (
        .din(new_Jinkela_wire_2850),
        .dout(new_Jinkela_wire_2851)
    );

    bfr new_Jinkela_buffer_12374 (
        .din(new_Jinkela_wire_14873),
        .dout(new_Jinkela_wire_14874)
    );

    and_ii _3000_ (
        .a(new_Jinkela_wire_1256),
        .b(new_Jinkela_wire_13045),
        .c(_0249_)
    );

    bfr new_Jinkela_buffer_15831 (
        .din(new_Jinkela_wire_18863),
        .dout(new_Jinkela_wire_18864)
    );

    bfr new_Jinkela_buffer_15923 (
        .din(new_Jinkela_wire_18975),
        .dout(new_Jinkela_wire_18976)
    );

    bfr new_Jinkela_buffer_15832 (
        .din(new_Jinkela_wire_18864),
        .dout(new_Jinkela_wire_18865)
    );

    bfr new_Jinkela_buffer_15925 (
        .din(new_Jinkela_wire_18981),
        .dout(new_Jinkela_wire_18982)
    );

    bfr new_Jinkela_buffer_15833 (
        .din(new_Jinkela_wire_18865),
        .dout(new_Jinkela_wire_18866)
    );

    spl2 new_Jinkela_splitter_1375 (
        .a(new_Jinkela_wire_18976),
        .b(new_Jinkela_wire_18977),
        .c(new_Jinkela_wire_18978)
    );

    bfr new_Jinkela_buffer_15834 (
        .din(new_Jinkela_wire_18866),
        .dout(new_Jinkela_wire_18867)
    );

    bfr new_Jinkela_buffer_15926 (
        .din(new_Jinkela_wire_18982),
        .dout(new_Jinkela_wire_18983)
    );

    bfr new_Jinkela_buffer_15835 (
        .din(new_Jinkela_wire_18867),
        .dout(new_Jinkela_wire_18868)
    );

    spl2 new_Jinkela_splitter_1380 (
        .a(_0231_),
        .b(new_Jinkela_wire_19050),
        .c(new_Jinkela_wire_19051)
    );

    bfr new_Jinkela_buffer_15836 (
        .din(new_Jinkela_wire_18868),
        .dout(new_Jinkela_wire_18869)
    );

    spl2 new_Jinkela_splitter_1379 (
        .a(_0924_),
        .b(new_Jinkela_wire_19048),
        .c(new_Jinkela_wire_19049)
    );

    bfr new_Jinkela_buffer_15837 (
        .din(new_Jinkela_wire_18869),
        .dout(new_Jinkela_wire_18870)
    );

    bfr new_Jinkela_buffer_15927 (
        .din(new_Jinkela_wire_18983),
        .dout(new_Jinkela_wire_18984)
    );

    bfr new_Jinkela_buffer_15838 (
        .din(new_Jinkela_wire_18870),
        .dout(new_Jinkela_wire_18871)
    );

    bfr new_Jinkela_buffer_15839 (
        .din(new_Jinkela_wire_18871),
        .dout(new_Jinkela_wire_18872)
    );

    bfr new_Jinkela_buffer_15928 (
        .din(new_Jinkela_wire_18984),
        .dout(new_Jinkela_wire_18985)
    );

    bfr new_Jinkela_buffer_15840 (
        .din(new_Jinkela_wire_18872),
        .dout(new_Jinkela_wire_18873)
    );

    spl2 new_Jinkela_splitter_1381 (
        .a(_1810_),
        .b(new_Jinkela_wire_19052),
        .c(new_Jinkela_wire_19053)
    );

    bfr new_Jinkela_buffer_15841 (
        .din(new_Jinkela_wire_18873),
        .dout(new_Jinkela_wire_18874)
    );

    bfr new_Jinkela_buffer_15929 (
        .din(new_Jinkela_wire_18985),
        .dout(new_Jinkela_wire_18986)
    );

    bfr new_Jinkela_buffer_15842 (
        .din(new_Jinkela_wire_18874),
        .dout(new_Jinkela_wire_18875)
    );

    bfr new_Jinkela_buffer_15987 (
        .din(_0386_),
        .dout(new_Jinkela_wire_19054)
    );

    bfr new_Jinkela_buffer_15843 (
        .din(new_Jinkela_wire_18875),
        .dout(new_Jinkela_wire_18876)
    );

    bfr new_Jinkela_buffer_15930 (
        .din(new_Jinkela_wire_18986),
        .dout(new_Jinkela_wire_18987)
    );

    bfr new_Jinkela_buffer_15844 (
        .din(new_Jinkela_wire_18876),
        .dout(new_Jinkela_wire_18877)
    );

    bfr new_Jinkela_buffer_15988 (
        .din(_0725_),
        .dout(new_Jinkela_wire_19057)
    );

    spl2 new_Jinkela_splitter_1382 (
        .a(_0530_),
        .b(new_Jinkela_wire_19055),
        .c(new_Jinkela_wire_19056)
    );

    bfr new_Jinkela_buffer_15845 (
        .din(new_Jinkela_wire_18877),
        .dout(new_Jinkela_wire_18878)
    );

    bfr new_Jinkela_buffer_15931 (
        .din(new_Jinkela_wire_18987),
        .dout(new_Jinkela_wire_18988)
    );

    bfr new_Jinkela_buffer_15846 (
        .din(new_Jinkela_wire_18878),
        .dout(new_Jinkela_wire_18879)
    );

    spl2 new_Jinkela_splitter_1385 (
        .a(_0784_),
        .b(new_Jinkela_wire_19063),
        .c(new_Jinkela_wire_19064)
    );

    bfr new_Jinkela_buffer_15847 (
        .din(new_Jinkela_wire_18879),
        .dout(new_Jinkela_wire_18880)
    );

    bfr new_Jinkela_buffer_15932 (
        .din(new_Jinkela_wire_18988),
        .dout(new_Jinkela_wire_18989)
    );

    bfr new_Jinkela_buffer_15848 (
        .din(new_Jinkela_wire_18880),
        .dout(new_Jinkela_wire_18881)
    );

    spl2 new_Jinkela_splitter_1384 (
        .a(_0661_),
        .b(new_Jinkela_wire_19061),
        .c(new_Jinkela_wire_19062)
    );

    bfr new_Jinkela_buffer_15849 (
        .din(new_Jinkela_wire_18881),
        .dout(new_Jinkela_wire_18882)
    );

    bfr new_Jinkela_buffer_15933 (
        .din(new_Jinkela_wire_18989),
        .dout(new_Jinkela_wire_18990)
    );

    bfr new_Jinkela_buffer_15850 (
        .din(new_Jinkela_wire_18882),
        .dout(new_Jinkela_wire_18883)
    );

    bfr new_Jinkela_buffer_15989 (
        .din(new_Jinkela_wire_19057),
        .dout(new_Jinkela_wire_19058)
    );

    bfr new_Jinkela_buffer_15851 (
        .din(new_Jinkela_wire_18883),
        .dout(new_Jinkela_wire_18884)
    );

    bfr new_Jinkela_buffer_15934 (
        .din(new_Jinkela_wire_18990),
        .dout(new_Jinkela_wire_18991)
    );

    bfr new_Jinkela_buffer_8916 (
        .din(new_Jinkela_wire_10907),
        .dout(new_Jinkela_wire_10908)
    );

    bfr new_Jinkela_buffer_9210 (
        .din(_0884_),
        .dout(new_Jinkela_wire_11234)
    );

    bfr new_Jinkela_buffer_8917 (
        .din(new_Jinkela_wire_10908),
        .dout(new_Jinkela_wire_10909)
    );

    bfr new_Jinkela_buffer_8996 (
        .din(new_Jinkela_wire_11001),
        .dout(new_Jinkela_wire_11002)
    );

    bfr new_Jinkela_buffer_8918 (
        .din(new_Jinkela_wire_10909),
        .dout(new_Jinkela_wire_10910)
    );

    bfr new_Jinkela_buffer_9024 (
        .din(new_Jinkela_wire_11033),
        .dout(new_Jinkela_wire_11034)
    );

    bfr new_Jinkela_buffer_8919 (
        .din(new_Jinkela_wire_10910),
        .dout(new_Jinkela_wire_10911)
    );

    bfr new_Jinkela_buffer_8997 (
        .din(new_Jinkela_wire_11002),
        .dout(new_Jinkela_wire_11003)
    );

    bfr new_Jinkela_buffer_8920 (
        .din(new_Jinkela_wire_10911),
        .dout(new_Jinkela_wire_10912)
    );

    bfr new_Jinkela_buffer_9035 (
        .din(new_Jinkela_wire_11050),
        .dout(new_Jinkela_wire_11051)
    );

    bfr new_Jinkela_buffer_8921 (
        .din(new_Jinkela_wire_10912),
        .dout(new_Jinkela_wire_10913)
    );

    bfr new_Jinkela_buffer_8998 (
        .din(new_Jinkela_wire_11003),
        .dout(new_Jinkela_wire_11004)
    );

    bfr new_Jinkela_buffer_8922 (
        .din(new_Jinkela_wire_10913),
        .dout(new_Jinkela_wire_10914)
    );

    bfr new_Jinkela_buffer_9025 (
        .din(new_Jinkela_wire_11034),
        .dout(new_Jinkela_wire_11035)
    );

    bfr new_Jinkela_buffer_8923 (
        .din(new_Jinkela_wire_10914),
        .dout(new_Jinkela_wire_10915)
    );

    bfr new_Jinkela_buffer_8999 (
        .din(new_Jinkela_wire_11004),
        .dout(new_Jinkela_wire_11005)
    );

    bfr new_Jinkela_buffer_8924 (
        .din(new_Jinkela_wire_10915),
        .dout(new_Jinkela_wire_10916)
    );

    bfr new_Jinkela_buffer_9119 (
        .din(new_Jinkela_wire_11138),
        .dout(new_Jinkela_wire_11139)
    );

    bfr new_Jinkela_buffer_8925 (
        .din(new_Jinkela_wire_10916),
        .dout(new_Jinkela_wire_10917)
    );

    bfr new_Jinkela_buffer_9000 (
        .din(new_Jinkela_wire_11005),
        .dout(new_Jinkela_wire_11006)
    );

    bfr new_Jinkela_buffer_8926 (
        .din(new_Jinkela_wire_10917),
        .dout(new_Jinkela_wire_10918)
    );

    bfr new_Jinkela_buffer_9026 (
        .din(new_Jinkela_wire_11035),
        .dout(new_Jinkela_wire_11036)
    );

    bfr new_Jinkela_buffer_8927 (
        .din(new_Jinkela_wire_10918),
        .dout(new_Jinkela_wire_10919)
    );

    bfr new_Jinkela_buffer_9001 (
        .din(new_Jinkela_wire_11006),
        .dout(new_Jinkela_wire_11007)
    );

    bfr new_Jinkela_buffer_8928 (
        .din(new_Jinkela_wire_10919),
        .dout(new_Jinkela_wire_10920)
    );

    bfr new_Jinkela_buffer_9036 (
        .din(new_Jinkela_wire_11051),
        .dout(new_Jinkela_wire_11052)
    );

    bfr new_Jinkela_buffer_8929 (
        .din(new_Jinkela_wire_10920),
        .dout(new_Jinkela_wire_10921)
    );

    bfr new_Jinkela_buffer_9002 (
        .din(new_Jinkela_wire_11007),
        .dout(new_Jinkela_wire_11008)
    );

    bfr new_Jinkela_buffer_8930 (
        .din(new_Jinkela_wire_10921),
        .dout(new_Jinkela_wire_10922)
    );

    bfr new_Jinkela_buffer_9027 (
        .din(new_Jinkela_wire_11036),
        .dout(new_Jinkela_wire_11037)
    );

    bfr new_Jinkela_buffer_8931 (
        .din(new_Jinkela_wire_10922),
        .dout(new_Jinkela_wire_10923)
    );

    bfr new_Jinkela_buffer_9003 (
        .din(new_Jinkela_wire_11008),
        .dout(new_Jinkela_wire_11009)
    );

    bfr new_Jinkela_buffer_8932 (
        .din(new_Jinkela_wire_10923),
        .dout(new_Jinkela_wire_10924)
    );

    bfr new_Jinkela_buffer_9206 (
        .din(new_Jinkela_wire_11229),
        .dout(new_Jinkela_wire_11230)
    );

    bfr new_Jinkela_buffer_8933 (
        .din(new_Jinkela_wire_10924),
        .dout(new_Jinkela_wire_10925)
    );

    bfr new_Jinkela_buffer_9004 (
        .din(new_Jinkela_wire_11009),
        .dout(new_Jinkela_wire_11010)
    );

    bfr new_Jinkela_buffer_8934 (
        .din(new_Jinkela_wire_10925),
        .dout(new_Jinkela_wire_10926)
    );

    spl2 new_Jinkela_splitter_854 (
        .a(new_Jinkela_wire_11037),
        .b(new_Jinkela_wire_11038),
        .c(new_Jinkela_wire_11039)
    );

    bfr new_Jinkela_buffer_8935 (
        .din(new_Jinkela_wire_10926),
        .dout(new_Jinkela_wire_10927)
    );

    bfr new_Jinkela_buffer_9005 (
        .din(new_Jinkela_wire_11010),
        .dout(new_Jinkela_wire_11011)
    );

    bfr new_Jinkela_buffer_8936 (
        .din(new_Jinkela_wire_10927),
        .dout(new_Jinkela_wire_10928)
    );

    bfr new_Jinkela_buffer_9037 (
        .din(new_Jinkela_wire_11052),
        .dout(new_Jinkela_wire_11053)
    );

    bfr new_Jinkela_buffer_5428 (
        .din(new_Jinkela_wire_6955),
        .dout(new_Jinkela_wire_6956)
    );

    or_bb _2077_ (
        .a(new_Jinkela_wire_2123),
        .b(new_Jinkela_wire_7691),
        .c(_1123_)
    );

    bfr new_Jinkela_buffer_5490 (
        .din(new_Jinkela_wire_7025),
        .dout(new_Jinkela_wire_7026)
    );

    or_bb _2078_ (
        .a(new_Jinkela_wire_10678),
        .b(new_Jinkela_wire_4238),
        .c(_1124_)
    );

    spl2 new_Jinkela_splitter_613 (
        .a(new_Jinkela_wire_6956),
        .b(new_Jinkela_wire_6957),
        .c(new_Jinkela_wire_6958)
    );

    and_bb _2079_ (
        .a(new_Jinkela_wire_451),
        .b(new_Jinkela_wire_343),
        .c(_1125_)
    );

    bfr new_Jinkela_buffer_5491 (
        .din(new_Jinkela_wire_7026),
        .dout(new_Jinkela_wire_7027)
    );

    and_bb _2080_ (
        .a(new_Jinkela_wire_10679),
        .b(new_Jinkela_wire_4239),
        .c(_1126_)
    );

    bfr new_Jinkela_buffer_5531 (
        .din(new_Jinkela_wire_7068),
        .dout(new_Jinkela_wire_7069)
    );

    or_bi _2081_ (
        .a(new_Jinkela_wire_13719),
        .b(new_Jinkela_wire_13316),
        .c(_1127_)
    );

    bfr new_Jinkela_buffer_5598 (
        .din(new_Jinkela_wire_7143),
        .dout(new_Jinkela_wire_7144)
    );

    and_ii _2082_ (
        .a(new_Jinkela_wire_16111),
        .b(new_Jinkela_wire_10672),
        .c(_1128_)
    );

    bfr new_Jinkela_buffer_5492 (
        .din(new_Jinkela_wire_7027),
        .dout(new_Jinkela_wire_7028)
    );

    and_bi _2083_ (
        .a(new_Jinkela_wire_13321),
        .b(new_Jinkela_wire_13955),
        .c(_1129_)
    );

    bfr new_Jinkela_buffer_5532 (
        .din(new_Jinkela_wire_7069),
        .dout(new_Jinkela_wire_7070)
    );

    and_bb _2084_ (
        .a(new_Jinkela_wire_104),
        .b(new_Jinkela_wire_463),
        .c(_1130_)
    );

    bfr new_Jinkela_buffer_5493 (
        .din(new_Jinkela_wire_7028),
        .dout(new_Jinkela_wire_7029)
    );

    and_bi _2085_ (
        .a(new_Jinkela_wire_11453),
        .b(new_Jinkela_wire_7692),
        .c(_1131_)
    );

    and_bb _2086_ (
        .a(new_Jinkela_wire_251),
        .b(new_Jinkela_wire_571),
        .c(_1132_)
    );

    spl2 new_Jinkela_splitter_625 (
        .a(_0334_),
        .b(new_Jinkela_wire_7184),
        .c(new_Jinkela_wire_7185)
    );

    bfr new_Jinkela_buffer_5494 (
        .din(new_Jinkela_wire_7029),
        .dout(new_Jinkela_wire_7030)
    );

    and_bi _2087_ (
        .a(new_Jinkela_wire_9555),
        .b(new_Jinkela_wire_7585),
        .c(_1133_)
    );

    bfr new_Jinkela_buffer_5533 (
        .din(new_Jinkela_wire_7070),
        .dout(new_Jinkela_wire_7071)
    );

    and_bb _2088_ (
        .a(new_Jinkela_wire_272),
        .b(new_Jinkela_wire_291),
        .c(_1134_)
    );

    bfr new_Jinkela_buffer_5495 (
        .din(new_Jinkela_wire_7030),
        .dout(new_Jinkela_wire_7031)
    );

    and_bi _2089_ (
        .a(new_Jinkela_wire_18790),
        .b(new_Jinkela_wire_3272),
        .c(_1135_)
    );

    bfr new_Jinkela_buffer_5599 (
        .din(new_Jinkela_wire_7144),
        .dout(new_Jinkela_wire_7145)
    );

    and_bb _2090_ (
        .a(new_Jinkela_wire_72),
        .b(new_Jinkela_wire_45),
        .c(_1136_)
    );

    bfr new_Jinkela_buffer_5496 (
        .din(new_Jinkela_wire_7031),
        .dout(new_Jinkela_wire_7032)
    );

    and_bi _2091_ (
        .a(new_Jinkela_wire_20338),
        .b(new_Jinkela_wire_15663),
        .c(_1137_)
    );

    bfr new_Jinkela_buffer_5534 (
        .din(new_Jinkela_wire_7071),
        .dout(new_Jinkela_wire_7072)
    );

    and_bb _2092_ (
        .a(new_Jinkela_wire_477),
        .b(new_Jinkela_wire_656),
        .c(_1138_)
    );

    bfr new_Jinkela_buffer_5497 (
        .din(new_Jinkela_wire_7032),
        .dout(new_Jinkela_wire_7033)
    );

    and_bi _2093_ (
        .a(new_Jinkela_wire_5103),
        .b(new_Jinkela_wire_20143),
        .c(_1139_)
    );

    and_bb _2094_ (
        .a(new_Jinkela_wire_363),
        .b(new_Jinkela_wire_633),
        .c(_1140_)
    );

    bfr new_Jinkela_buffer_5498 (
        .din(new_Jinkela_wire_7033),
        .dout(new_Jinkela_wire_7034)
    );

    and_bi _2095_ (
        .a(new_Jinkela_wire_8287),
        .b(new_Jinkela_wire_3891),
        .c(_1141_)
    );

    bfr new_Jinkela_buffer_5535 (
        .din(new_Jinkela_wire_7072),
        .dout(new_Jinkela_wire_7073)
    );

    and_bb _2096_ (
        .a(new_Jinkela_wire_691),
        .b(new_Jinkela_wire_537),
        .c(_1142_)
    );

    bfr new_Jinkela_buffer_5499 (
        .din(new_Jinkela_wire_7034),
        .dout(new_Jinkela_wire_7035)
    );

    or_ii _2097_ (
        .a(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_23),
        .c(_1143_)
    );

    bfr new_Jinkela_buffer_5600 (
        .din(new_Jinkela_wire_7145),
        .dout(new_Jinkela_wire_7146)
    );

    and_bi _2098_ (
        .a(new_Jinkela_wire_17068),
        .b(new_Jinkela_wire_1568),
        .c(_1144_)
    );

    bfr new_Jinkela_buffer_5500 (
        .din(new_Jinkela_wire_7035),
        .dout(new_Jinkela_wire_7036)
    );

    and_bb _2099_ (
        .a(new_Jinkela_wire_238),
        .b(new_Jinkela_wire_43),
        .c(_1145_)
    );

    bfr new_Jinkela_buffer_5536 (
        .din(new_Jinkela_wire_7073),
        .dout(new_Jinkela_wire_7074)
    );

    and_bi _2100_ (
        .a(new_Jinkela_wire_5433),
        .b(new_Jinkela_wire_17049),
        .c(_1146_)
    );

    bfr new_Jinkela_buffer_5501 (
        .din(new_Jinkela_wire_7036),
        .dout(new_Jinkela_wire_7037)
    );

    and_ii _2101_ (
        .a(new_Jinkela_wire_5720),
        .b(new_Jinkela_wire_3958),
        .c(_1147_)
    );

    bfr new_Jinkela_buffer_5629 (
        .din(new_Jinkela_wire_7178),
        .dout(new_Jinkela_wire_7179)
    );

    or_bb _2102_ (
        .a(new_Jinkela_wire_15754),
        .b(new_Jinkela_wire_4302),
        .c(_1148_)
    );

    bfr new_Jinkela_buffer_5502 (
        .din(new_Jinkela_wire_7037),
        .dout(new_Jinkela_wire_7038)
    );

    or_ii _2103_ (
        .a(new_Jinkela_wire_15755),
        .b(new_Jinkela_wire_4301),
        .c(_1149_)
    );

    bfr new_Jinkela_buffer_5537 (
        .din(new_Jinkela_wire_7074),
        .dout(new_Jinkela_wire_7075)
    );

    or_ii _2104_ (
        .a(new_Jinkela_wire_21123),
        .b(new_Jinkela_wire_3703),
        .c(_1150_)
    );

    bfr new_Jinkela_buffer_5503 (
        .din(new_Jinkela_wire_7038),
        .dout(new_Jinkela_wire_7039)
    );

    and_ii _2105_ (
        .a(new_Jinkela_wire_9094),
        .b(new_Jinkela_wire_16378),
        .c(_1151_)
    );

    bfr new_Jinkela_buffer_5601 (
        .din(new_Jinkela_wire_7146),
        .dout(new_Jinkela_wire_7147)
    );

    and_bb _2106_ (
        .a(new_Jinkela_wire_9095),
        .b(new_Jinkela_wire_16379),
        .c(_1152_)
    );

    bfr new_Jinkela_buffer_5504 (
        .din(new_Jinkela_wire_7039),
        .dout(new_Jinkela_wire_7040)
    );

    or_bb _2107_ (
        .a(new_Jinkela_wire_18121),
        .b(new_Jinkela_wire_18761),
        .c(_1153_)
    );

    bfr new_Jinkela_buffer_5538 (
        .din(new_Jinkela_wire_7075),
        .dout(new_Jinkela_wire_7076)
    );

    or_bb _2108_ (
        .a(new_Jinkela_wire_17079),
        .b(new_Jinkela_wire_14307),
        .c(_1154_)
    );

    bfr new_Jinkela_buffer_5505 (
        .din(new_Jinkela_wire_7040),
        .dout(new_Jinkela_wire_7041)
    );

    or_ii _2109_ (
        .a(new_Jinkela_wire_17080),
        .b(new_Jinkela_wire_14308),
        .c(_1155_)
    );

    bfr new_Jinkela_buffer_5633 (
        .din(_1689_),
        .dout(new_Jinkela_wire_7187)
    );

    or_ii _2110_ (
        .a(new_Jinkela_wire_17994),
        .b(new_Jinkela_wire_12615),
        .c(_1156_)
    );

    bfr new_Jinkela_buffer_5632 (
        .din(_1607_),
        .dout(new_Jinkela_wire_7186)
    );

    bfr new_Jinkela_buffer_5506 (
        .din(new_Jinkela_wire_7041),
        .dout(new_Jinkela_wire_7042)
    );

    and_ii _2111_ (
        .a(new_Jinkela_wire_3439),
        .b(new_Jinkela_wire_1001),
        .c(_1157_)
    );

    bfr new_Jinkela_buffer_5539 (
        .din(new_Jinkela_wire_7076),
        .dout(new_Jinkela_wire_7077)
    );

    and_bb _2112_ (
        .a(new_Jinkela_wire_3440),
        .b(new_Jinkela_wire_1002),
        .c(_1158_)
    );

    bfr new_Jinkela_buffer_5507 (
        .din(new_Jinkela_wire_7042),
        .dout(new_Jinkela_wire_7043)
    );

    or_bb _2113_ (
        .a(new_Jinkela_wire_18103),
        .b(new_Jinkela_wire_5995),
        .c(_1159_)
    );

    bfr new_Jinkela_buffer_5602 (
        .din(new_Jinkela_wire_7147),
        .dout(new_Jinkela_wire_7148)
    );

    or_bb _2114_ (
        .a(new_Jinkela_wire_4829),
        .b(new_Jinkela_wire_6238),
        .c(_1160_)
    );

    bfr new_Jinkela_buffer_5508 (
        .din(new_Jinkela_wire_7043),
        .dout(new_Jinkela_wire_7044)
    );

    or_ii _2115_ (
        .a(new_Jinkela_wire_4830),
        .b(new_Jinkela_wire_6239),
        .c(_1161_)
    );

    bfr new_Jinkela_buffer_5540 (
        .din(new_Jinkela_wire_7077),
        .dout(new_Jinkela_wire_7078)
    );

    or_ii _2116_ (
        .a(new_Jinkela_wire_12737),
        .b(new_Jinkela_wire_17031),
        .c(_1162_)
    );

    bfr new_Jinkela_buffer_5509 (
        .din(new_Jinkela_wire_7044),
        .dout(new_Jinkela_wire_7045)
    );

    and_ii _2117_ (
        .a(new_Jinkela_wire_14325),
        .b(new_Jinkela_wire_16939),
        .c(_1163_)
    );

    bfr new_Jinkela_buffer_5630 (
        .din(new_Jinkela_wire_7179),
        .dout(new_Jinkela_wire_7180)
    );

    and_bb _2118_ (
        .a(new_Jinkela_wire_14326),
        .b(new_Jinkela_wire_16940),
        .c(_1164_)
    );

    bfr new_Jinkela_buffer_12438 (
        .din(new_Jinkela_wire_14939),
        .dout(new_Jinkela_wire_14940)
    );

    bfr new_Jinkela_buffer_12375 (
        .din(new_Jinkela_wire_14874),
        .dout(new_Jinkela_wire_14875)
    );

    bfr new_Jinkela_buffer_12531 (
        .din(new_Jinkela_wire_15038),
        .dout(new_Jinkela_wire_15039)
    );

    bfr new_Jinkela_buffer_12376 (
        .din(new_Jinkela_wire_14875),
        .dout(new_Jinkela_wire_14876)
    );

    bfr new_Jinkela_buffer_12439 (
        .din(new_Jinkela_wire_14940),
        .dout(new_Jinkela_wire_14941)
    );

    bfr new_Jinkela_buffer_12377 (
        .din(new_Jinkela_wire_14876),
        .dout(new_Jinkela_wire_14877)
    );

    bfr new_Jinkela_buffer_12511 (
        .din(new_Jinkela_wire_15014),
        .dout(new_Jinkela_wire_15015)
    );

    bfr new_Jinkela_buffer_12378 (
        .din(new_Jinkela_wire_14877),
        .dout(new_Jinkela_wire_14878)
    );

    bfr new_Jinkela_buffer_12440 (
        .din(new_Jinkela_wire_14941),
        .dout(new_Jinkela_wire_14942)
    );

    bfr new_Jinkela_buffer_12379 (
        .din(new_Jinkela_wire_14878),
        .dout(new_Jinkela_wire_14879)
    );

    bfr new_Jinkela_buffer_12613 (
        .din(new_Jinkela_wire_15128),
        .dout(new_Jinkela_wire_15129)
    );

    bfr new_Jinkela_buffer_12380 (
        .din(new_Jinkela_wire_14879),
        .dout(new_Jinkela_wire_14880)
    );

    bfr new_Jinkela_buffer_12441 (
        .din(new_Jinkela_wire_14942),
        .dout(new_Jinkela_wire_14943)
    );

    bfr new_Jinkela_buffer_12381 (
        .din(new_Jinkela_wire_14880),
        .dout(new_Jinkela_wire_14881)
    );

    bfr new_Jinkela_buffer_12512 (
        .din(new_Jinkela_wire_15015),
        .dout(new_Jinkela_wire_15016)
    );

    bfr new_Jinkela_buffer_12382 (
        .din(new_Jinkela_wire_14881),
        .dout(new_Jinkela_wire_14882)
    );

    bfr new_Jinkela_buffer_12442 (
        .din(new_Jinkela_wire_14943),
        .dout(new_Jinkela_wire_14944)
    );

    bfr new_Jinkela_buffer_12383 (
        .din(new_Jinkela_wire_14882),
        .dout(new_Jinkela_wire_14883)
    );

    bfr new_Jinkela_buffer_12532 (
        .din(new_Jinkela_wire_15039),
        .dout(new_Jinkela_wire_15040)
    );

    bfr new_Jinkela_buffer_12384 (
        .din(new_Jinkela_wire_14883),
        .dout(new_Jinkela_wire_14884)
    );

    bfr new_Jinkela_buffer_12443 (
        .din(new_Jinkela_wire_14944),
        .dout(new_Jinkela_wire_14945)
    );

    bfr new_Jinkela_buffer_12385 (
        .din(new_Jinkela_wire_14884),
        .dout(new_Jinkela_wire_14885)
    );

    bfr new_Jinkela_buffer_12513 (
        .din(new_Jinkela_wire_15016),
        .dout(new_Jinkela_wire_15017)
    );

    bfr new_Jinkela_buffer_12386 (
        .din(new_Jinkela_wire_14885),
        .dout(new_Jinkela_wire_14886)
    );

    bfr new_Jinkela_buffer_12444 (
        .din(new_Jinkela_wire_14945),
        .dout(new_Jinkela_wire_14946)
    );

    bfr new_Jinkela_buffer_12387 (
        .din(new_Jinkela_wire_14886),
        .dout(new_Jinkela_wire_14887)
    );

    bfr new_Jinkela_buffer_12684 (
        .din(_0747_),
        .dout(new_Jinkela_wire_15206)
    );

    bfr new_Jinkela_buffer_12388 (
        .din(new_Jinkela_wire_14887),
        .dout(new_Jinkela_wire_14888)
    );

    bfr new_Jinkela_buffer_12445 (
        .din(new_Jinkela_wire_14946),
        .dout(new_Jinkela_wire_14947)
    );

    bfr new_Jinkela_buffer_12389 (
        .din(new_Jinkela_wire_14888),
        .dout(new_Jinkela_wire_14889)
    );

    bfr new_Jinkela_buffer_12514 (
        .din(new_Jinkela_wire_15017),
        .dout(new_Jinkela_wire_15018)
    );

    spl2 new_Jinkela_splitter_1099 (
        .a(new_Jinkela_wire_14889),
        .b(new_Jinkela_wire_14890),
        .c(new_Jinkela_wire_14891)
    );

    bfr new_Jinkela_buffer_12533 (
        .din(new_Jinkela_wire_15040),
        .dout(new_Jinkela_wire_15041)
    );

    bfr new_Jinkela_buffer_12446 (
        .din(new_Jinkela_wire_14947),
        .dout(new_Jinkela_wire_14948)
    );

    bfr new_Jinkela_buffer_12447 (
        .din(new_Jinkela_wire_14948),
        .dout(new_Jinkela_wire_14949)
    );

    bfr new_Jinkela_buffer_12515 (
        .din(new_Jinkela_wire_15018),
        .dout(new_Jinkela_wire_15019)
    );

    bfr new_Jinkela_buffer_12448 (
        .din(new_Jinkela_wire_14949),
        .dout(new_Jinkela_wire_14950)
    );

    bfr new_Jinkela_buffer_12614 (
        .din(new_Jinkela_wire_15129),
        .dout(new_Jinkela_wire_15130)
    );

    bfr new_Jinkela_buffer_12449 (
        .din(new_Jinkela_wire_14950),
        .dout(new_Jinkela_wire_14951)
    );

    bfr new_Jinkela_buffer_12516 (
        .din(new_Jinkela_wire_15019),
        .dout(new_Jinkela_wire_15020)
    );

    bfr new_Jinkela_buffer_12450 (
        .din(new_Jinkela_wire_14951),
        .dout(new_Jinkela_wire_14952)
    );

    bfr new_Jinkela_buffer_12534 (
        .din(new_Jinkela_wire_15041),
        .dout(new_Jinkela_wire_15042)
    );

    bfr new_Jinkela_buffer_15852 (
        .din(new_Jinkela_wire_18884),
        .dout(new_Jinkela_wire_18885)
    );

    bfr new_Jinkela_buffer_15853 (
        .din(new_Jinkela_wire_18885),
        .dout(new_Jinkela_wire_18886)
    );

    bfr new_Jinkela_buffer_15935 (
        .din(new_Jinkela_wire_18991),
        .dout(new_Jinkela_wire_18992)
    );

    bfr new_Jinkela_buffer_15854 (
        .din(new_Jinkela_wire_18886),
        .dout(new_Jinkela_wire_18887)
    );

    spl2 new_Jinkela_splitter_1383 (
        .a(new_Jinkela_wire_19058),
        .b(new_Jinkela_wire_19059),
        .c(new_Jinkela_wire_19060)
    );

    bfr new_Jinkela_buffer_15855 (
        .din(new_Jinkela_wire_18887),
        .dout(new_Jinkela_wire_18888)
    );

    bfr new_Jinkela_buffer_15936 (
        .din(new_Jinkela_wire_18992),
        .dout(new_Jinkela_wire_18993)
    );

    bfr new_Jinkela_buffer_15856 (
        .din(new_Jinkela_wire_18888),
        .dout(new_Jinkela_wire_18889)
    );

    bfr new_Jinkela_buffer_15998 (
        .din(_1514_),
        .dout(new_Jinkela_wire_19079)
    );

    bfr new_Jinkela_buffer_15990 (
        .din(_1219_),
        .dout(new_Jinkela_wire_19067)
    );

    bfr new_Jinkela_buffer_15857 (
        .din(new_Jinkela_wire_18889),
        .dout(new_Jinkela_wire_18890)
    );

    bfr new_Jinkela_buffer_15937 (
        .din(new_Jinkela_wire_18993),
        .dout(new_Jinkela_wire_18994)
    );

    bfr new_Jinkela_buffer_15858 (
        .din(new_Jinkela_wire_18890),
        .dout(new_Jinkela_wire_18891)
    );

    spl2 new_Jinkela_splitter_1386 (
        .a(_1722_),
        .b(new_Jinkela_wire_19065),
        .c(new_Jinkela_wire_19066)
    );

    bfr new_Jinkela_buffer_15859 (
        .din(new_Jinkela_wire_18891),
        .dout(new_Jinkela_wire_18892)
    );

    bfr new_Jinkela_buffer_15938 (
        .din(new_Jinkela_wire_18994),
        .dout(new_Jinkela_wire_18995)
    );

    bfr new_Jinkela_buffer_15860 (
        .din(new_Jinkela_wire_18892),
        .dout(new_Jinkela_wire_18893)
    );

    bfr new_Jinkela_buffer_15999 (
        .din(_1647_),
        .dout(new_Jinkela_wire_19080)
    );

    spl2 new_Jinkela_splitter_1388 (
        .a(_1275_),
        .b(new_Jinkela_wire_19077),
        .c(new_Jinkela_wire_19078)
    );

    bfr new_Jinkela_buffer_15861 (
        .din(new_Jinkela_wire_18893),
        .dout(new_Jinkela_wire_18894)
    );

    bfr new_Jinkela_buffer_15939 (
        .din(new_Jinkela_wire_18995),
        .dout(new_Jinkela_wire_18996)
    );

    bfr new_Jinkela_buffer_15862 (
        .din(new_Jinkela_wire_18894),
        .dout(new_Jinkela_wire_18895)
    );

    bfr new_Jinkela_buffer_15991 (
        .din(new_Jinkela_wire_19067),
        .dout(new_Jinkela_wire_19068)
    );

    bfr new_Jinkela_buffer_15863 (
        .din(new_Jinkela_wire_18895),
        .dout(new_Jinkela_wire_18896)
    );

    bfr new_Jinkela_buffer_15940 (
        .din(new_Jinkela_wire_18996),
        .dout(new_Jinkela_wire_18997)
    );

    bfr new_Jinkela_buffer_15864 (
        .din(new_Jinkela_wire_18896),
        .dout(new_Jinkela_wire_18897)
    );

    bfr new_Jinkela_buffer_16000 (
        .din(_1026_),
        .dout(new_Jinkela_wire_19081)
    );

    bfr new_Jinkela_buffer_15865 (
        .din(new_Jinkela_wire_18897),
        .dout(new_Jinkela_wire_18898)
    );

    bfr new_Jinkela_buffer_15941 (
        .din(new_Jinkela_wire_18997),
        .dout(new_Jinkela_wire_18998)
    );

    bfr new_Jinkela_buffer_15866 (
        .din(new_Jinkela_wire_18898),
        .dout(new_Jinkela_wire_18899)
    );

    bfr new_Jinkela_buffer_15992 (
        .din(new_Jinkela_wire_19068),
        .dout(new_Jinkela_wire_19069)
    );

    bfr new_Jinkela_buffer_15867 (
        .din(new_Jinkela_wire_18899),
        .dout(new_Jinkela_wire_18900)
    );

    bfr new_Jinkela_buffer_15942 (
        .din(new_Jinkela_wire_18998),
        .dout(new_Jinkela_wire_18999)
    );

    bfr new_Jinkela_buffer_15868 (
        .din(new_Jinkela_wire_18900),
        .dout(new_Jinkela_wire_18901)
    );

    bfr new_Jinkela_buffer_15993 (
        .din(new_Jinkela_wire_19069),
        .dout(new_Jinkela_wire_19070)
    );

    bfr new_Jinkela_buffer_15869 (
        .din(new_Jinkela_wire_18901),
        .dout(new_Jinkela_wire_18902)
    );

    bfr new_Jinkela_buffer_15943 (
        .din(new_Jinkela_wire_18999),
        .dout(new_Jinkela_wire_19000)
    );

    bfr new_Jinkela_buffer_15870 (
        .din(new_Jinkela_wire_18902),
        .dout(new_Jinkela_wire_18903)
    );

    bfr new_Jinkela_buffer_15871 (
        .din(new_Jinkela_wire_18903),
        .dout(new_Jinkela_wire_18904)
    );

    bfr new_Jinkela_buffer_15944 (
        .din(new_Jinkela_wire_19000),
        .dout(new_Jinkela_wire_19001)
    );

    bfr new_Jinkela_buffer_15872 (
        .din(new_Jinkela_wire_18904),
        .dout(new_Jinkela_wire_18905)
    );

    spl2 new_Jinkela_splitter_1390 (
        .a(_1193_),
        .b(new_Jinkela_wire_19107),
        .c(new_Jinkela_wire_19108)
    );

    bfr new_Jinkela_buffer_8937 (
        .din(new_Jinkela_wire_10928),
        .dout(new_Jinkela_wire_10929)
    );

    and_bb _3001_ (
        .a(new_Jinkela_wire_1257),
        .b(new_Jinkela_wire_13046),
        .c(_0250_)
    );

    bfr new_Jinkela_buffer_9006 (
        .din(new_Jinkela_wire_11011),
        .dout(new_Jinkela_wire_11012)
    );

    or_bb _3002_ (
        .a(new_Jinkela_wire_6737),
        .b(new_Jinkela_wire_19118),
        .c(_0251_)
    );

    bfr new_Jinkela_buffer_8938 (
        .din(new_Jinkela_wire_10929),
        .dout(new_Jinkela_wire_10930)
    );

    and_ii _3003_ (
        .a(new_Jinkela_wire_9181),
        .b(new_Jinkela_wire_2941),
        .c(_0253_)
    );

    bfr new_Jinkela_buffer_9120 (
        .din(new_Jinkela_wire_11139),
        .dout(new_Jinkela_wire_11140)
    );

    and_bb _3004_ (
        .a(new_Jinkela_wire_9182),
        .b(new_Jinkela_wire_2942),
        .c(_0254_)
    );

    bfr new_Jinkela_buffer_8939 (
        .din(new_Jinkela_wire_10930),
        .dout(new_Jinkela_wire_10931)
    );

    or_bb _3005_ (
        .a(new_Jinkela_wire_14213),
        .b(new_Jinkela_wire_16694),
        .c(_0255_)
    );

    bfr new_Jinkela_buffer_9007 (
        .din(new_Jinkela_wire_11012),
        .dout(new_Jinkela_wire_11013)
    );

    and_ii _3006_ (
        .a(new_Jinkela_wire_3193),
        .b(new_Jinkela_wire_10202),
        .c(_0256_)
    );

    bfr new_Jinkela_buffer_8940 (
        .din(new_Jinkela_wire_10931),
        .dout(new_Jinkela_wire_10932)
    );

    and_bb _3007_ (
        .a(new_Jinkela_wire_3194),
        .b(new_Jinkela_wire_10203),
        .c(_0257_)
    );

    bfr new_Jinkela_buffer_9038 (
        .din(new_Jinkela_wire_11053),
        .dout(new_Jinkela_wire_11054)
    );

    or_bb _3008_ (
        .a(new_Jinkela_wire_7737),
        .b(new_Jinkela_wire_2653),
        .c(_0258_)
    );

    bfr new_Jinkela_buffer_8941 (
        .din(new_Jinkela_wire_10932),
        .dout(new_Jinkela_wire_10933)
    );

    and_ii _3009_ (
        .a(new_Jinkela_wire_5282),
        .b(new_Jinkela_wire_19050),
        .c(_0259_)
    );

    bfr new_Jinkela_buffer_9008 (
        .din(new_Jinkela_wire_11013),
        .dout(new_Jinkela_wire_11014)
    );

    and_bb _3010_ (
        .a(new_Jinkela_wire_5283),
        .b(new_Jinkela_wire_19051),
        .c(_0260_)
    );

    bfr new_Jinkela_buffer_8942 (
        .din(new_Jinkela_wire_10933),
        .dout(new_Jinkela_wire_10934)
    );

    or_bb _3011_ (
        .a(new_Jinkela_wire_10674),
        .b(new_Jinkela_wire_2137),
        .c(_0261_)
    );

    and_ii _3012_ (
        .a(new_Jinkela_wire_16114),
        .b(new_Jinkela_wire_18443),
        .c(_0262_)
    );

    bfr new_Jinkela_buffer_9314 (
        .din(_0277_),
        .dout(new_Jinkela_wire_11340)
    );

    bfr new_Jinkela_buffer_8943 (
        .din(new_Jinkela_wire_10934),
        .dout(new_Jinkela_wire_10935)
    );

    and_bb _3013_ (
        .a(new_Jinkela_wire_16115),
        .b(new_Jinkela_wire_18444),
        .c(_0264_)
    );

    bfr new_Jinkela_buffer_9009 (
        .din(new_Jinkela_wire_11014),
        .dout(new_Jinkela_wire_11015)
    );

    or_bb _3014_ (
        .a(new_Jinkela_wire_18380),
        .b(new_Jinkela_wire_2135),
        .c(_0265_)
    );

    bfr new_Jinkela_buffer_8944 (
        .din(new_Jinkela_wire_10935),
        .dout(new_Jinkela_wire_10936)
    );

    and_ii _3015_ (
        .a(new_Jinkela_wire_3118),
        .b(new_Jinkela_wire_8691),
        .c(_0266_)
    );

    bfr new_Jinkela_buffer_9039 (
        .din(new_Jinkela_wire_11054),
        .dout(new_Jinkela_wire_11055)
    );

    and_bb _3016_ (
        .a(new_Jinkela_wire_3119),
        .b(new_Jinkela_wire_8692),
        .c(_0267_)
    );

    bfr new_Jinkela_buffer_8945 (
        .din(new_Jinkela_wire_10936),
        .dout(new_Jinkela_wire_10937)
    );

    or_bb _3017_ (
        .a(new_Jinkela_wire_2945),
        .b(new_Jinkela_wire_11422),
        .c(_0268_)
    );

    spl2 new_Jinkela_splitter_852 (
        .a(new_Jinkela_wire_11015),
        .b(new_Jinkela_wire_11016),
        .c(new_Jinkela_wire_11017)
    );

    and_ii _3018_ (
        .a(new_Jinkela_wire_13464),
        .b(new_Jinkela_wire_17856),
        .c(_0269_)
    );

    bfr new_Jinkela_buffer_8946 (
        .din(new_Jinkela_wire_10937),
        .dout(new_Jinkela_wire_10938)
    );

    and_bb _3019_ (
        .a(new_Jinkela_wire_13465),
        .b(new_Jinkela_wire_17857),
        .c(_0270_)
    );

    bfr new_Jinkela_buffer_9040 (
        .din(new_Jinkela_wire_11055),
        .dout(new_Jinkela_wire_11056)
    );

    or_bb _3020_ (
        .a(new_Jinkela_wire_14100),
        .b(new_Jinkela_wire_10261),
        .c(_0271_)
    );

    bfr new_Jinkela_buffer_8947 (
        .din(new_Jinkela_wire_10938),
        .dout(new_Jinkela_wire_10939)
    );

    and_ii _3021_ (
        .a(new_Jinkela_wire_1009),
        .b(new_Jinkela_wire_5437),
        .c(_0272_)
    );

    bfr new_Jinkela_buffer_9121 (
        .din(new_Jinkela_wire_11140),
        .dout(new_Jinkela_wire_11141)
    );

    and_bb _3022_ (
        .a(new_Jinkela_wire_1010),
        .b(new_Jinkela_wire_5438),
        .c(_0273_)
    );

    bfr new_Jinkela_buffer_8948 (
        .din(new_Jinkela_wire_10939),
        .dout(new_Jinkela_wire_10940)
    );

    or_bb _3023_ (
        .a(new_Jinkela_wire_15752),
        .b(new_Jinkela_wire_4696),
        .c(_0275_)
    );

    and_ii _3024_ (
        .a(new_Jinkela_wire_5129),
        .b(new_Jinkela_wire_20208),
        .c(_0276_)
    );

    bfr new_Jinkela_buffer_9315 (
        .din(_1637_),
        .dout(new_Jinkela_wire_11341)
    );

    bfr new_Jinkela_buffer_8949 (
        .din(new_Jinkela_wire_10940),
        .dout(new_Jinkela_wire_10941)
    );

    and_bb _3025_ (
        .a(new_Jinkela_wire_5130),
        .b(new_Jinkela_wire_20209),
        .c(_0277_)
    );

    bfr new_Jinkela_buffer_9041 (
        .din(new_Jinkela_wire_11056),
        .dout(new_Jinkela_wire_11057)
    );

    or_bb _3026_ (
        .a(new_Jinkela_wire_11340),
        .b(new_Jinkela_wire_21164),
        .c(_0278_)
    );

    bfr new_Jinkela_buffer_8950 (
        .din(new_Jinkela_wire_10941),
        .dout(new_Jinkela_wire_10942)
    );

    and_ii _3027_ (
        .a(new_Jinkela_wire_4569),
        .b(new_Jinkela_wire_13392),
        .c(_0279_)
    );

    bfr new_Jinkela_buffer_9122 (
        .din(new_Jinkela_wire_11141),
        .dout(new_Jinkela_wire_11142)
    );

    and_bb _3028_ (
        .a(new_Jinkela_wire_4570),
        .b(new_Jinkela_wire_13393),
        .c(_0280_)
    );

    bfr new_Jinkela_buffer_8951 (
        .din(new_Jinkela_wire_10942),
        .dout(new_Jinkela_wire_10943)
    );

    or_bb _3029_ (
        .a(new_Jinkela_wire_5739),
        .b(new_Jinkela_wire_15996),
        .c(_0281_)
    );

    bfr new_Jinkela_buffer_9042 (
        .din(new_Jinkela_wire_11057),
        .dout(new_Jinkela_wire_11058)
    );

    and_ii _3030_ (
        .a(new_Jinkela_wire_5445),
        .b(new_Jinkela_wire_15467),
        .c(_0282_)
    );

    bfr new_Jinkela_buffer_8952 (
        .din(new_Jinkela_wire_10943),
        .dout(new_Jinkela_wire_10944)
    );

    and_bb _3031_ (
        .a(new_Jinkela_wire_5446),
        .b(new_Jinkela_wire_15468),
        .c(_0283_)
    );

    bfr new_Jinkela_buffer_9207 (
        .din(new_Jinkela_wire_11230),
        .dout(new_Jinkela_wire_11231)
    );

    or_bb _3032_ (
        .a(new_Jinkela_wire_6678),
        .b(new_Jinkela_wire_13149),
        .c(_0284_)
    );

    bfr new_Jinkela_buffer_8953 (
        .din(new_Jinkela_wire_10944),
        .dout(new_Jinkela_wire_10945)
    );

    and_ii _3033_ (
        .a(new_Jinkela_wire_11404),
        .b(new_Jinkela_wire_12065),
        .c(_0286_)
    );

    bfr new_Jinkela_buffer_9043 (
        .din(new_Jinkela_wire_11058),
        .dout(new_Jinkela_wire_11059)
    );

    and_bb _3034_ (
        .a(new_Jinkela_wire_11405),
        .b(new_Jinkela_wire_12066),
        .c(_0287_)
    );

    bfr new_Jinkela_buffer_8954 (
        .din(new_Jinkela_wire_10945),
        .dout(new_Jinkela_wire_10946)
    );

    or_bb _3035_ (
        .a(new_Jinkela_wire_14198),
        .b(new_Jinkela_wire_14266),
        .c(_0288_)
    );

    bfr new_Jinkela_buffer_9123 (
        .din(new_Jinkela_wire_11142),
        .dout(new_Jinkela_wire_11143)
    );

    and_ii _3036_ (
        .a(new_Jinkela_wire_17668),
        .b(new_Jinkela_wire_9444),
        .c(_0289_)
    );

    bfr new_Jinkela_buffer_8955 (
        .din(new_Jinkela_wire_10946),
        .dout(new_Jinkela_wire_10947)
    );

    and_bb _3037_ (
        .a(new_Jinkela_wire_17669),
        .b(new_Jinkela_wire_9445),
        .c(_0290_)
    );

    bfr new_Jinkela_buffer_9044 (
        .din(new_Jinkela_wire_11059),
        .dout(new_Jinkela_wire_11060)
    );

    or_bb _3038_ (
        .a(new_Jinkela_wire_5703),
        .b(new_Jinkela_wire_17547),
        .c(_0291_)
    );

    bfr new_Jinkela_buffer_8956 (
        .din(new_Jinkela_wire_10947),
        .dout(new_Jinkela_wire_10948)
    );

    and_ii _3039_ (
        .a(new_Jinkela_wire_17798),
        .b(new_Jinkela_wire_18961),
        .c(_0292_)
    );

    bfr new_Jinkela_buffer_9211 (
        .din(new_Jinkela_wire_11234),
        .dout(new_Jinkela_wire_11235)
    );

    and_bb _3040_ (
        .a(new_Jinkela_wire_17799),
        .b(new_Jinkela_wire_18962),
        .c(_0293_)
    );

    spl2 new_Jinkela_splitter_845 (
        .a(new_Jinkela_wire_10948),
        .b(new_Jinkela_wire_10949),
        .c(new_Jinkela_wire_10950)
    );

    or_bb _3041_ (
        .a(new_Jinkela_wire_9746),
        .b(new_Jinkela_wire_13724),
        .c(_0294_)
    );

    bfr new_Jinkela_buffer_9045 (
        .din(new_Jinkela_wire_11060),
        .dout(new_Jinkela_wire_11061)
    );

    and_ii _3042_ (
        .a(new_Jinkela_wire_10112),
        .b(new_Jinkela_wire_6510),
        .c(_0295_)
    );

    bfr new_Jinkela_buffer_1930 (
        .din(new_Jinkela_wire_2851),
        .dout(new_Jinkela_wire_2852)
    );

    bfr new_Jinkela_buffer_2172 (
        .din(_1573_),
        .dout(new_Jinkela_wire_3122)
    );

    bfr new_Jinkela_buffer_2029 (
        .din(new_Jinkela_wire_2970),
        .dout(new_Jinkela_wire_2971)
    );

    bfr new_Jinkela_buffer_1931 (
        .din(new_Jinkela_wire_2852),
        .dout(new_Jinkela_wire_2853)
    );

    spl2 new_Jinkela_splitter_326 (
        .a(_0943_),
        .b(new_Jinkela_wire_3182),
        .c(new_Jinkela_wire_3183)
    );

    bfr new_Jinkela_buffer_1932 (
        .din(new_Jinkela_wire_2853),
        .dout(new_Jinkela_wire_2854)
    );

    bfr new_Jinkela_buffer_2030 (
        .din(new_Jinkela_wire_2971),
        .dout(new_Jinkela_wire_2972)
    );

    bfr new_Jinkela_buffer_1933 (
        .din(new_Jinkela_wire_2854),
        .dout(new_Jinkela_wire_2855)
    );

    spl2 new_Jinkela_splitter_325 (
        .a(_1163_),
        .b(new_Jinkela_wire_3180),
        .c(new_Jinkela_wire_3181)
    );

    bfr new_Jinkela_buffer_1934 (
        .din(new_Jinkela_wire_2855),
        .dout(new_Jinkela_wire_2856)
    );

    bfr new_Jinkela_buffer_2173 (
        .din(new_Jinkela_wire_3122),
        .dout(new_Jinkela_wire_3123)
    );

    bfr new_Jinkela_buffer_2031 (
        .din(new_Jinkela_wire_2972),
        .dout(new_Jinkela_wire_2973)
    );

    bfr new_Jinkela_buffer_1935 (
        .din(new_Jinkela_wire_2856),
        .dout(new_Jinkela_wire_2857)
    );

    bfr new_Jinkela_buffer_1936 (
        .din(new_Jinkela_wire_2857),
        .dout(new_Jinkela_wire_2858)
    );

    bfr new_Jinkela_buffer_2032 (
        .din(new_Jinkela_wire_2973),
        .dout(new_Jinkela_wire_2974)
    );

    bfr new_Jinkela_buffer_1937 (
        .din(new_Jinkela_wire_2858),
        .dout(new_Jinkela_wire_2859)
    );

    bfr new_Jinkela_buffer_1938 (
        .din(new_Jinkela_wire_2859),
        .dout(new_Jinkela_wire_2860)
    );

    bfr new_Jinkela_buffer_2174 (
        .din(new_Jinkela_wire_3123),
        .dout(new_Jinkela_wire_3124)
    );

    bfr new_Jinkela_buffer_2033 (
        .din(new_Jinkela_wire_2974),
        .dout(new_Jinkela_wire_2975)
    );

    bfr new_Jinkela_buffer_1939 (
        .din(new_Jinkela_wire_2860),
        .dout(new_Jinkela_wire_2861)
    );

    bfr new_Jinkela_buffer_1940 (
        .din(new_Jinkela_wire_2861),
        .dout(new_Jinkela_wire_2862)
    );

    bfr new_Jinkela_buffer_2034 (
        .din(new_Jinkela_wire_2975),
        .dout(new_Jinkela_wire_2976)
    );

    bfr new_Jinkela_buffer_1941 (
        .din(new_Jinkela_wire_2862),
        .dout(new_Jinkela_wire_2863)
    );

    spl2 new_Jinkela_splitter_327 (
        .a(_1574_),
        .b(new_Jinkela_wire_3184),
        .c(new_Jinkela_wire_3185)
    );

    bfr new_Jinkela_buffer_1942 (
        .din(new_Jinkela_wire_2863),
        .dout(new_Jinkela_wire_2864)
    );

    bfr new_Jinkela_buffer_2175 (
        .din(new_Jinkela_wire_3124),
        .dout(new_Jinkela_wire_3125)
    );

    bfr new_Jinkela_buffer_2035 (
        .din(new_Jinkela_wire_2976),
        .dout(new_Jinkela_wire_2977)
    );

    bfr new_Jinkela_buffer_1943 (
        .din(new_Jinkela_wire_2864),
        .dout(new_Jinkela_wire_2865)
    );

    bfr new_Jinkela_buffer_1944 (
        .din(new_Jinkela_wire_2865),
        .dout(new_Jinkela_wire_2866)
    );

    bfr new_Jinkela_buffer_2036 (
        .din(new_Jinkela_wire_2977),
        .dout(new_Jinkela_wire_2978)
    );

    bfr new_Jinkela_buffer_1945 (
        .din(new_Jinkela_wire_2866),
        .dout(new_Jinkela_wire_2867)
    );

    bfr new_Jinkela_buffer_2228 (
        .din(_1043_),
        .dout(new_Jinkela_wire_3186)
    );

    bfr new_Jinkela_buffer_1946 (
        .din(new_Jinkela_wire_2867),
        .dout(new_Jinkela_wire_2868)
    );

    bfr new_Jinkela_buffer_2176 (
        .din(new_Jinkela_wire_3125),
        .dout(new_Jinkela_wire_3126)
    );

    bfr new_Jinkela_buffer_2037 (
        .din(new_Jinkela_wire_2978),
        .dout(new_Jinkela_wire_2979)
    );

    bfr new_Jinkela_buffer_1947 (
        .din(new_Jinkela_wire_2868),
        .dout(new_Jinkela_wire_2869)
    );

    bfr new_Jinkela_buffer_1948 (
        .din(new_Jinkela_wire_2869),
        .dout(new_Jinkela_wire_2870)
    );

    bfr new_Jinkela_buffer_2229 (
        .din(_0138_),
        .dout(new_Jinkela_wire_3189)
    );

    bfr new_Jinkela_buffer_2038 (
        .din(new_Jinkela_wire_2979),
        .dout(new_Jinkela_wire_2980)
    );

    bfr new_Jinkela_buffer_1949 (
        .din(new_Jinkela_wire_2870),
        .dout(new_Jinkela_wire_2871)
    );

    spl2 new_Jinkela_splitter_328 (
        .a(_0132_),
        .b(new_Jinkela_wire_3187),
        .c(new_Jinkela_wire_3188)
    );

    bfr new_Jinkela_buffer_1950 (
        .din(new_Jinkela_wire_2871),
        .dout(new_Jinkela_wire_2872)
    );

    bfr new_Jinkela_buffer_2177 (
        .din(new_Jinkela_wire_3126),
        .dout(new_Jinkela_wire_3127)
    );

    bfr new_Jinkela_buffer_15873 (
        .din(new_Jinkela_wire_18905),
        .dout(new_Jinkela_wire_18906)
    );

    or_bb _2119_ (
        .a(new_Jinkela_wire_6193),
        .b(new_Jinkela_wire_3180),
        .c(_1165_)
    );

    bfr new_Jinkela_buffer_15945 (
        .din(new_Jinkela_wire_19001),
        .dout(new_Jinkela_wire_19002)
    );

    or_bb _2120_ (
        .a(new_Jinkela_wire_8276),
        .b(new_Jinkela_wire_16971),
        .c(_1166_)
    );

    bfr new_Jinkela_buffer_15874 (
        .din(new_Jinkela_wire_18906),
        .dout(new_Jinkela_wire_18907)
    );

    or_ii _2121_ (
        .a(new_Jinkela_wire_8277),
        .b(new_Jinkela_wire_16972),
        .c(_1167_)
    );

    bfr new_Jinkela_buffer_15994 (
        .din(new_Jinkela_wire_19070),
        .dout(new_Jinkela_wire_19071)
    );

    or_ii _2122_ (
        .a(new_Jinkela_wire_6421),
        .b(new_Jinkela_wire_1003),
        .c(_1168_)
    );

    bfr new_Jinkela_buffer_15875 (
        .din(new_Jinkela_wire_18907),
        .dout(new_Jinkela_wire_18908)
    );

    and_ii _2123_ (
        .a(new_Jinkela_wire_15203),
        .b(new_Jinkela_wire_8016),
        .c(_1169_)
    );

    bfr new_Jinkela_buffer_15946 (
        .din(new_Jinkela_wire_19002),
        .dout(new_Jinkela_wire_19003)
    );

    and_bb _2124_ (
        .a(new_Jinkela_wire_15204),
        .b(new_Jinkela_wire_8017),
        .c(_1170_)
    );

    bfr new_Jinkela_buffer_15876 (
        .din(new_Jinkela_wire_18908),
        .dout(new_Jinkela_wire_18909)
    );

    or_bb _2125_ (
        .a(new_Jinkela_wire_14327),
        .b(new_Jinkela_wire_10835),
        .c(_1171_)
    );

    or_bb _2126_ (
        .a(new_Jinkela_wire_15200),
        .b(new_Jinkela_wire_19739),
        .c(_1172_)
    );

    bfr new_Jinkela_buffer_16024 (
        .din(_0306_),
        .dout(new_Jinkela_wire_19109)
    );

    bfr new_Jinkela_buffer_15877 (
        .din(new_Jinkela_wire_18909),
        .dout(new_Jinkela_wire_18910)
    );

    or_ii _2127_ (
        .a(new_Jinkela_wire_15201),
        .b(new_Jinkela_wire_19740),
        .c(_1173_)
    );

    bfr new_Jinkela_buffer_15947 (
        .din(new_Jinkela_wire_19003),
        .dout(new_Jinkela_wire_19004)
    );

    or_ii _2128_ (
        .a(new_Jinkela_wire_4082),
        .b(new_Jinkela_wire_8843),
        .c(_1174_)
    );

    bfr new_Jinkela_buffer_15878 (
        .din(new_Jinkela_wire_18910),
        .dout(new_Jinkela_wire_18911)
    );

    and_ii _2129_ (
        .a(new_Jinkela_wire_18535),
        .b(new_Jinkela_wire_6732),
        .c(_1175_)
    );

    bfr new_Jinkela_buffer_15995 (
        .din(new_Jinkela_wire_19071),
        .dout(new_Jinkela_wire_19072)
    );

    and_bb _2130_ (
        .a(new_Jinkela_wire_18536),
        .b(new_Jinkela_wire_6733),
        .c(_1176_)
    );

    bfr new_Jinkela_buffer_15879 (
        .din(new_Jinkela_wire_18911),
        .dout(new_Jinkela_wire_18912)
    );

    or_bb _2131_ (
        .a(new_Jinkela_wire_832),
        .b(new_Jinkela_wire_2458),
        .c(_1177_)
    );

    bfr new_Jinkela_buffer_15948 (
        .din(new_Jinkela_wire_19004),
        .dout(new_Jinkela_wire_19005)
    );

    or_bb _2132_ (
        .a(new_Jinkela_wire_5439),
        .b(new_Jinkela_wire_19274),
        .c(_1178_)
    );

    bfr new_Jinkela_buffer_15880 (
        .din(new_Jinkela_wire_18912),
        .dout(new_Jinkela_wire_18913)
    );

    or_ii _2133_ (
        .a(new_Jinkela_wire_5440),
        .b(new_Jinkela_wire_19275),
        .c(_1179_)
    );

    bfr new_Jinkela_buffer_16001 (
        .din(new_Jinkela_wire_19081),
        .dout(new_Jinkela_wire_19082)
    );

    or_ii _2134_ (
        .a(new_Jinkela_wire_4988),
        .b(new_Jinkela_wire_13574),
        .c(_1180_)
    );

    bfr new_Jinkela_buffer_15881 (
        .din(new_Jinkela_wire_18913),
        .dout(new_Jinkela_wire_18914)
    );

    and_ii _2135_ (
        .a(new_Jinkela_wire_14010),
        .b(new_Jinkela_wire_2651),
        .c(_1181_)
    );

    bfr new_Jinkela_buffer_15949 (
        .din(new_Jinkela_wire_19005),
        .dout(new_Jinkela_wire_19006)
    );

    and_bb _2136_ (
        .a(new_Jinkela_wire_14011),
        .b(new_Jinkela_wire_2652),
        .c(_1182_)
    );

    bfr new_Jinkela_buffer_15882 (
        .din(new_Jinkela_wire_18914),
        .dout(new_Jinkela_wire_18915)
    );

    or_bb _2137_ (
        .a(new_Jinkela_wire_14310),
        .b(new_Jinkela_wire_11395),
        .c(_1183_)
    );

    bfr new_Jinkela_buffer_15996 (
        .din(new_Jinkela_wire_19072),
        .dout(new_Jinkela_wire_19073)
    );

    or_bb _2138_ (
        .a(new_Jinkela_wire_19908),
        .b(new_Jinkela_wire_20265),
        .c(_1184_)
    );

    bfr new_Jinkela_buffer_15883 (
        .din(new_Jinkela_wire_18915),
        .dout(new_Jinkela_wire_18916)
    );

    or_ii _2139_ (
        .a(new_Jinkela_wire_19909),
        .b(new_Jinkela_wire_20266),
        .c(_1185_)
    );

    bfr new_Jinkela_buffer_15950 (
        .din(new_Jinkela_wire_19006),
        .dout(new_Jinkela_wire_19007)
    );

    or_ii _2140_ (
        .a(new_Jinkela_wire_15836),
        .b(new_Jinkela_wire_10951),
        .c(_1186_)
    );

    bfr new_Jinkela_buffer_15884 (
        .din(new_Jinkela_wire_18916),
        .dout(new_Jinkela_wire_18917)
    );

    and_ii _2141_ (
        .a(new_Jinkela_wire_13195),
        .b(new_Jinkela_wire_3950),
        .c(_1187_)
    );

    and_bb _2142_ (
        .a(new_Jinkela_wire_13196),
        .b(new_Jinkela_wire_3951),
        .c(_1188_)
    );

    bfr new_Jinkela_buffer_15885 (
        .din(new_Jinkela_wire_18917),
        .dout(new_Jinkela_wire_18918)
    );

    or_bb _2143_ (
        .a(new_Jinkela_wire_16120),
        .b(new_Jinkela_wire_7273),
        .c(_1189_)
    );

    bfr new_Jinkela_buffer_15951 (
        .din(new_Jinkela_wire_19007),
        .dout(new_Jinkela_wire_19008)
    );

    or_bb _2144_ (
        .a(new_Jinkela_wire_11616),
        .b(new_Jinkela_wire_20396),
        .c(_1190_)
    );

    bfr new_Jinkela_buffer_15886 (
        .din(new_Jinkela_wire_18918),
        .dout(new_Jinkela_wire_18919)
    );

    and_bb _2145_ (
        .a(new_Jinkela_wire_11617),
        .b(new_Jinkela_wire_20397),
        .c(_1191_)
    );

    bfr new_Jinkela_buffer_15997 (
        .din(new_Jinkela_wire_19073),
        .dout(new_Jinkela_wire_19074)
    );

    or_bi _2146_ (
        .a(new_Jinkela_wire_13389),
        .b(new_Jinkela_wire_6242),
        .c(_1192_)
    );

    bfr new_Jinkela_buffer_15887 (
        .din(new_Jinkela_wire_18919),
        .dout(new_Jinkela_wire_18920)
    );

    and_ii _2147_ (
        .a(new_Jinkela_wire_19791),
        .b(new_Jinkela_wire_19538),
        .c(_1193_)
    );

    bfr new_Jinkela_buffer_15952 (
        .din(new_Jinkela_wire_19008),
        .dout(new_Jinkela_wire_19009)
    );

    and_bb _2148_ (
        .a(new_Jinkela_wire_19792),
        .b(new_Jinkela_wire_19539),
        .c(_1194_)
    );

    bfr new_Jinkela_buffer_15888 (
        .din(new_Jinkela_wire_18920),
        .dout(new_Jinkela_wire_18921)
    );

    or_bb _2149_ (
        .a(new_Jinkela_wire_5126),
        .b(new_Jinkela_wire_19107),
        .c(new_net_3956)
    );

    bfr new_Jinkela_buffer_16002 (
        .din(new_Jinkela_wire_19082),
        .dout(new_Jinkela_wire_19083)
    );

    or_ii _2150_ (
        .a(new_Jinkela_wire_308),
        .b(new_Jinkela_wire_330),
        .c(_1195_)
    );

    bfr new_Jinkela_buffer_15889 (
        .din(new_Jinkela_wire_18921),
        .dout(new_Jinkela_wire_18922)
    );

    and_bi _2151_ (
        .a(new_Jinkela_wire_5132),
        .b(new_Jinkela_wire_5429),
        .c(_1196_)
    );

    bfr new_Jinkela_buffer_15953 (
        .din(new_Jinkela_wire_19009),
        .dout(new_Jinkela_wire_19010)
    );

    and_bi _2152_ (
        .a(new_Jinkela_wire_16106),
        .b(new_Jinkela_wire_1572),
        .c(new_net_3958)
    );

    bfr new_Jinkela_buffer_15890 (
        .din(new_Jinkela_wire_18922),
        .dout(new_Jinkela_wire_18923)
    );

    and_bb _2153_ (
        .a(new_Jinkela_wire_4906),
        .b(new_Jinkela_wire_18308),
        .c(_1197_)
    );

    spl2 new_Jinkela_splitter_1387 (
        .a(new_Jinkela_wire_19074),
        .b(new_Jinkela_wire_19075),
        .c(new_Jinkela_wire_19076)
    );

    or_bb _2154_ (
        .a(new_Jinkela_wire_18106),
        .b(new_Jinkela_wire_5543),
        .c(new_net_3930)
    );

    bfr new_Jinkela_buffer_15891 (
        .din(new_Jinkela_wire_18923),
        .dout(new_Jinkela_wire_18924)
    );

    and_bb _2155_ (
        .a(new_Jinkela_wire_17859),
        .b(new_Jinkela_wire_5042),
        .c(_1198_)
    );

    bfr new_Jinkela_buffer_15954 (
        .din(new_Jinkela_wire_19010),
        .dout(new_Jinkela_wire_19011)
    );

    or_bb _2156_ (
        .a(new_Jinkela_wire_21197),
        .b(new_Jinkela_wire_6860),
        .c(new_net_3950)
    );

    bfr new_Jinkela_buffer_15892 (
        .din(new_Jinkela_wire_18924),
        .dout(new_Jinkela_wire_18925)
    );

    and_bb _2157_ (
        .a(new_Jinkela_wire_16112),
        .b(new_Jinkela_wire_10673),
        .c(_1199_)
    );

    spl2 new_Jinkela_splitter_1392 (
        .a(_0870_),
        .b(new_Jinkela_wire_19112),
        .c(new_Jinkela_wire_19113)
    );

    or_bb _2158_ (
        .a(new_Jinkela_wire_984),
        .b(new_Jinkela_wire_13956),
        .c(new_net_3928)
    );

    spl2 new_Jinkela_splitter_1391 (
        .a(_0474_),
        .b(new_Jinkela_wire_19110),
        .c(new_Jinkela_wire_19111)
    );

    bfr new_Jinkela_buffer_15893 (
        .din(new_Jinkela_wire_18925),
        .dout(new_Jinkela_wire_18926)
    );

    and_bb _2159_ (
        .a(new_Jinkela_wire_13054),
        .b(new_Jinkela_wire_7501),
        .c(_1200_)
    );

    bfr new_Jinkela_buffer_15955 (
        .din(new_Jinkela_wire_19011),
        .dout(new_Jinkela_wire_19012)
    );

    or_bb _2160_ (
        .a(new_Jinkela_wire_6691),
        .b(new_Jinkela_wire_19327),
        .c(new_net_3932)
    );

    bfr new_Jinkela_buffer_5510 (
        .din(new_Jinkela_wire_7045),
        .dout(new_Jinkela_wire_7046)
    );

    bfr new_Jinkela_buffer_5541 (
        .din(new_Jinkela_wire_7078),
        .dout(new_Jinkela_wire_7079)
    );

    bfr new_Jinkela_buffer_5511 (
        .din(new_Jinkela_wire_7046),
        .dout(new_Jinkela_wire_7047)
    );

    bfr new_Jinkela_buffer_5603 (
        .din(new_Jinkela_wire_7148),
        .dout(new_Jinkela_wire_7149)
    );

    bfr new_Jinkela_buffer_5512 (
        .din(new_Jinkela_wire_7047),
        .dout(new_Jinkela_wire_7048)
    );

    bfr new_Jinkela_buffer_5542 (
        .din(new_Jinkela_wire_7079),
        .dout(new_Jinkela_wire_7080)
    );

    bfr new_Jinkela_buffer_5513 (
        .din(new_Jinkela_wire_7048),
        .dout(new_Jinkela_wire_7049)
    );

    bfr new_Jinkela_buffer_5705 (
        .din(_1014_),
        .dout(new_Jinkela_wire_7261)
    );

    bfr new_Jinkela_buffer_5514 (
        .din(new_Jinkela_wire_7049),
        .dout(new_Jinkela_wire_7050)
    );

    bfr new_Jinkela_buffer_5543 (
        .din(new_Jinkela_wire_7080),
        .dout(new_Jinkela_wire_7081)
    );

    spl2 new_Jinkela_splitter_617 (
        .a(new_Jinkela_wire_7050),
        .b(new_Jinkela_wire_7051),
        .c(new_Jinkela_wire_7052)
    );

    bfr new_Jinkela_buffer_5544 (
        .din(new_Jinkela_wire_7081),
        .dout(new_Jinkela_wire_7082)
    );

    bfr new_Jinkela_buffer_5604 (
        .din(new_Jinkela_wire_7149),
        .dout(new_Jinkela_wire_7150)
    );

    bfr new_Jinkela_buffer_5631 (
        .din(new_Jinkela_wire_7180),
        .dout(new_Jinkela_wire_7181)
    );

    bfr new_Jinkela_buffer_5545 (
        .din(new_Jinkela_wire_7082),
        .dout(new_Jinkela_wire_7083)
    );

    bfr new_Jinkela_buffer_5605 (
        .din(new_Jinkela_wire_7150),
        .dout(new_Jinkela_wire_7151)
    );

    bfr new_Jinkela_buffer_5546 (
        .din(new_Jinkela_wire_7083),
        .dout(new_Jinkela_wire_7084)
    );

    bfr new_Jinkela_buffer_5706 (
        .din(_0204_),
        .dout(new_Jinkela_wire_7262)
    );

    bfr new_Jinkela_buffer_5547 (
        .din(new_Jinkela_wire_7084),
        .dout(new_Jinkela_wire_7085)
    );

    bfr new_Jinkela_buffer_5606 (
        .din(new_Jinkela_wire_7151),
        .dout(new_Jinkela_wire_7152)
    );

    bfr new_Jinkela_buffer_5548 (
        .din(new_Jinkela_wire_7085),
        .dout(new_Jinkela_wire_7086)
    );

    bfr new_Jinkela_buffer_5634 (
        .din(new_Jinkela_wire_7187),
        .dout(new_Jinkela_wire_7188)
    );

    bfr new_Jinkela_buffer_5549 (
        .din(new_Jinkela_wire_7086),
        .dout(new_Jinkela_wire_7087)
    );

    bfr new_Jinkela_buffer_5607 (
        .din(new_Jinkela_wire_7152),
        .dout(new_Jinkela_wire_7153)
    );

    bfr new_Jinkela_buffer_5550 (
        .din(new_Jinkela_wire_7087),
        .dout(new_Jinkela_wire_7088)
    );

    spl2 new_Jinkela_splitter_627 (
        .a(_0669_),
        .b(new_Jinkela_wire_7263),
        .c(new_Jinkela_wire_7264)
    );

    bfr new_Jinkela_buffer_5551 (
        .din(new_Jinkela_wire_7088),
        .dout(new_Jinkela_wire_7089)
    );

    bfr new_Jinkela_buffer_5608 (
        .din(new_Jinkela_wire_7153),
        .dout(new_Jinkela_wire_7154)
    );

    bfr new_Jinkela_buffer_5552 (
        .din(new_Jinkela_wire_7089),
        .dout(new_Jinkela_wire_7090)
    );

    bfr new_Jinkela_buffer_5635 (
        .din(new_Jinkela_wire_7188),
        .dout(new_Jinkela_wire_7189)
    );

    bfr new_Jinkela_buffer_5553 (
        .din(new_Jinkela_wire_7090),
        .dout(new_Jinkela_wire_7091)
    );

    bfr new_Jinkela_buffer_5609 (
        .din(new_Jinkela_wire_7154),
        .dout(new_Jinkela_wire_7155)
    );

    bfr new_Jinkela_buffer_5554 (
        .din(new_Jinkela_wire_7091),
        .dout(new_Jinkela_wire_7092)
    );

    bfr new_Jinkela_buffer_5711 (
        .din(_1439_),
        .dout(new_Jinkela_wire_7269)
    );

    bfr new_Jinkela_buffer_5707 (
        .din(new_Jinkela_wire_7264),
        .dout(new_Jinkela_wire_7265)
    );

    bfr new_Jinkela_buffer_5555 (
        .din(new_Jinkela_wire_7092),
        .dout(new_Jinkela_wire_7093)
    );

    bfr new_Jinkela_buffer_5610 (
        .din(new_Jinkela_wire_7155),
        .dout(new_Jinkela_wire_7156)
    );

    bfr new_Jinkela_buffer_5556 (
        .din(new_Jinkela_wire_7093),
        .dout(new_Jinkela_wire_7094)
    );

    bfr new_Jinkela_buffer_5636 (
        .din(new_Jinkela_wire_7189),
        .dout(new_Jinkela_wire_7190)
    );

    bfr new_Jinkela_buffer_5557 (
        .din(new_Jinkela_wire_7094),
        .dout(new_Jinkela_wire_7095)
    );

    bfr new_Jinkela_buffer_5611 (
        .din(new_Jinkela_wire_7156),
        .dout(new_Jinkela_wire_7157)
    );

    bfr new_Jinkela_buffer_5558 (
        .din(new_Jinkela_wire_7095),
        .dout(new_Jinkela_wire_7096)
    );

    bfr new_Jinkela_buffer_2039 (
        .din(new_Jinkela_wire_2980),
        .dout(new_Jinkela_wire_2981)
    );

    bfr new_Jinkela_buffer_12451 (
        .din(new_Jinkela_wire_14952),
        .dout(new_Jinkela_wire_14953)
    );

    bfr new_Jinkela_buffer_15894 (
        .din(new_Jinkela_wire_18926),
        .dout(new_Jinkela_wire_18927)
    );

    bfr new_Jinkela_buffer_1951 (
        .din(new_Jinkela_wire_2872),
        .dout(new_Jinkela_wire_2873)
    );

    bfr new_Jinkela_buffer_12517 (
        .din(new_Jinkela_wire_15020),
        .dout(new_Jinkela_wire_15021)
    );

    bfr new_Jinkela_buffer_16003 (
        .din(new_Jinkela_wire_19083),
        .dout(new_Jinkela_wire_19084)
    );

    bfr new_Jinkela_buffer_12452 (
        .din(new_Jinkela_wire_14953),
        .dout(new_Jinkela_wire_14954)
    );

    bfr new_Jinkela_buffer_15895 (
        .din(new_Jinkela_wire_18927),
        .dout(new_Jinkela_wire_18928)
    );

    bfr new_Jinkela_buffer_1952 (
        .din(new_Jinkela_wire_2873),
        .dout(new_Jinkela_wire_2874)
    );

    bfr new_Jinkela_buffer_15956 (
        .din(new_Jinkela_wire_19012),
        .dout(new_Jinkela_wire_19013)
    );

    bfr new_Jinkela_buffer_12685 (
        .din(new_net_3958),
        .dout(new_Jinkela_wire_15207)
    );

    bfr new_Jinkela_buffer_2040 (
        .din(new_Jinkela_wire_2981),
        .dout(new_Jinkela_wire_2982)
    );

    bfr new_Jinkela_buffer_12453 (
        .din(new_Jinkela_wire_14954),
        .dout(new_Jinkela_wire_14955)
    );

    bfr new_Jinkela_buffer_15896 (
        .din(new_Jinkela_wire_18928),
        .dout(new_Jinkela_wire_18929)
    );

    bfr new_Jinkela_buffer_1953 (
        .din(new_Jinkela_wire_2874),
        .dout(new_Jinkela_wire_2875)
    );

    bfr new_Jinkela_buffer_12518 (
        .din(new_Jinkela_wire_15021),
        .dout(new_Jinkela_wire_15022)
    );

    spl2 new_Jinkela_splitter_329 (
        .a(_1572_),
        .b(new_Jinkela_wire_3191),
        .c(new_Jinkela_wire_3192)
    );

    bfr new_Jinkela_buffer_12454 (
        .din(new_Jinkela_wire_14955),
        .dout(new_Jinkela_wire_14956)
    );

    bfr new_Jinkela_buffer_15897 (
        .din(new_Jinkela_wire_18929),
        .dout(new_Jinkela_wire_18930)
    );

    bfr new_Jinkela_buffer_1954 (
        .din(new_Jinkela_wire_2875),
        .dout(new_Jinkela_wire_2876)
    );

    bfr new_Jinkela_buffer_12535 (
        .din(new_Jinkela_wire_15042),
        .dout(new_Jinkela_wire_15043)
    );

    bfr new_Jinkela_buffer_15957 (
        .din(new_Jinkela_wire_19013),
        .dout(new_Jinkela_wire_19014)
    );

    bfr new_Jinkela_buffer_2178 (
        .din(new_Jinkela_wire_3127),
        .dout(new_Jinkela_wire_3128)
    );

    bfr new_Jinkela_buffer_2041 (
        .din(new_Jinkela_wire_2982),
        .dout(new_Jinkela_wire_2983)
    );

    bfr new_Jinkela_buffer_12455 (
        .din(new_Jinkela_wire_14956),
        .dout(new_Jinkela_wire_14957)
    );

    bfr new_Jinkela_buffer_15898 (
        .din(new_Jinkela_wire_18930),
        .dout(new_Jinkela_wire_18931)
    );

    bfr new_Jinkela_buffer_1955 (
        .din(new_Jinkela_wire_2876),
        .dout(new_Jinkela_wire_2877)
    );

    spl2 new_Jinkela_splitter_1101 (
        .a(new_Jinkela_wire_15022),
        .b(new_Jinkela_wire_15023),
        .c(new_Jinkela_wire_15024)
    );

    bfr new_Jinkela_buffer_16004 (
        .din(new_Jinkela_wire_19084),
        .dout(new_Jinkela_wire_19085)
    );

    bfr new_Jinkela_buffer_12456 (
        .din(new_Jinkela_wire_14957),
        .dout(new_Jinkela_wire_14958)
    );

    bfr new_Jinkela_buffer_15899 (
        .din(new_Jinkela_wire_18931),
        .dout(new_Jinkela_wire_18932)
    );

    bfr new_Jinkela_buffer_1956 (
        .din(new_Jinkela_wire_2877),
        .dout(new_Jinkela_wire_2878)
    );

    bfr new_Jinkela_buffer_12536 (
        .din(new_Jinkela_wire_15043),
        .dout(new_Jinkela_wire_15044)
    );

    bfr new_Jinkela_buffer_15958 (
        .din(new_Jinkela_wire_19014),
        .dout(new_Jinkela_wire_19015)
    );

    bfr new_Jinkela_buffer_2042 (
        .din(new_Jinkela_wire_2983),
        .dout(new_Jinkela_wire_2984)
    );

    bfr new_Jinkela_buffer_12457 (
        .din(new_Jinkela_wire_14958),
        .dout(new_Jinkela_wire_14959)
    );

    bfr new_Jinkela_buffer_15900 (
        .din(new_Jinkela_wire_18932),
        .dout(new_Jinkela_wire_18933)
    );

    bfr new_Jinkela_buffer_1957 (
        .din(new_Jinkela_wire_2878),
        .dout(new_Jinkela_wire_2879)
    );

    bfr new_Jinkela_buffer_12615 (
        .din(new_Jinkela_wire_15130),
        .dout(new_Jinkela_wire_15131)
    );

    spl2 new_Jinkela_splitter_1393 (
        .a(_1715_),
        .b(new_Jinkela_wire_19114),
        .c(new_Jinkela_wire_19115)
    );

    bfr new_Jinkela_buffer_2230 (
        .din(_1710_),
        .dout(new_Jinkela_wire_3190)
    );

    bfr new_Jinkela_buffer_12458 (
        .din(new_Jinkela_wire_14959),
        .dout(new_Jinkela_wire_14960)
    );

    bfr new_Jinkela_buffer_15901 (
        .din(new_Jinkela_wire_18933),
        .dout(new_Jinkela_wire_18934)
    );

    bfr new_Jinkela_buffer_1958 (
        .din(new_Jinkela_wire_2879),
        .dout(new_Jinkela_wire_2880)
    );

    bfr new_Jinkela_buffer_15959 (
        .din(new_Jinkela_wire_19015),
        .dout(new_Jinkela_wire_19016)
    );

    bfr new_Jinkela_buffer_2179 (
        .din(new_Jinkela_wire_3128),
        .dout(new_Jinkela_wire_3129)
    );

    bfr new_Jinkela_buffer_12857 (
        .din(new_net_3924),
        .dout(new_Jinkela_wire_15379)
    );

    bfr new_Jinkela_buffer_2043 (
        .din(new_Jinkela_wire_2984),
        .dout(new_Jinkela_wire_2985)
    );

    bfr new_Jinkela_buffer_12459 (
        .din(new_Jinkela_wire_14960),
        .dout(new_Jinkela_wire_14961)
    );

    bfr new_Jinkela_buffer_15902 (
        .din(new_Jinkela_wire_18934),
        .dout(new_Jinkela_wire_18935)
    );

    bfr new_Jinkela_buffer_1959 (
        .din(new_Jinkela_wire_2880),
        .dout(new_Jinkela_wire_2881)
    );

    bfr new_Jinkela_buffer_12537 (
        .din(new_Jinkela_wire_15044),
        .dout(new_Jinkela_wire_15045)
    );

    bfr new_Jinkela_buffer_16005 (
        .din(new_Jinkela_wire_19085),
        .dout(new_Jinkela_wire_19086)
    );

    bfr new_Jinkela_buffer_12460 (
        .din(new_Jinkela_wire_14961),
        .dout(new_Jinkela_wire_14962)
    );

    bfr new_Jinkela_buffer_15903 (
        .din(new_Jinkela_wire_18935),
        .dout(new_Jinkela_wire_18936)
    );

    bfr new_Jinkela_buffer_1960 (
        .din(new_Jinkela_wire_2881),
        .dout(new_Jinkela_wire_2882)
    );

    bfr new_Jinkela_buffer_12616 (
        .din(new_Jinkela_wire_15131),
        .dout(new_Jinkela_wire_15132)
    );

    bfr new_Jinkela_buffer_15960 (
        .din(new_Jinkela_wire_19016),
        .dout(new_Jinkela_wire_19017)
    );

    spl2 new_Jinkela_splitter_330 (
        .a(_0255_),
        .b(new_Jinkela_wire_3193),
        .c(new_Jinkela_wire_3194)
    );

    bfr new_Jinkela_buffer_2044 (
        .din(new_Jinkela_wire_2985),
        .dout(new_Jinkela_wire_2986)
    );

    bfr new_Jinkela_buffer_12461 (
        .din(new_Jinkela_wire_14962),
        .dout(new_Jinkela_wire_14963)
    );

    bfr new_Jinkela_buffer_15904 (
        .din(new_Jinkela_wire_18936),
        .dout(new_Jinkela_wire_18937)
    );

    bfr new_Jinkela_buffer_1961 (
        .din(new_Jinkela_wire_2882),
        .dout(new_Jinkela_wire_2883)
    );

    bfr new_Jinkela_buffer_12538 (
        .din(new_Jinkela_wire_15045),
        .dout(new_Jinkela_wire_15046)
    );

    spl2 new_Jinkela_splitter_1394 (
        .a(_0644_),
        .b(new_Jinkela_wire_19116),
        .c(new_Jinkela_wire_19117)
    );

    bfr new_Jinkela_buffer_2231 (
        .din(_1578_),
        .dout(new_Jinkela_wire_3197)
    );

    bfr new_Jinkela_buffer_12462 (
        .din(new_Jinkela_wire_14963),
        .dout(new_Jinkela_wire_14964)
    );

    bfr new_Jinkela_buffer_15905 (
        .din(new_Jinkela_wire_18937),
        .dout(new_Jinkela_wire_18938)
    );

    bfr new_Jinkela_buffer_1962 (
        .din(new_Jinkela_wire_2883),
        .dout(new_Jinkela_wire_2884)
    );

    bfr new_Jinkela_buffer_15961 (
        .din(new_Jinkela_wire_19017),
        .dout(new_Jinkela_wire_19018)
    );

    bfr new_Jinkela_buffer_2180 (
        .din(new_Jinkela_wire_3129),
        .dout(new_Jinkela_wire_3130)
    );

    bfr new_Jinkela_buffer_12686 (
        .din(new_Jinkela_wire_15207),
        .dout(new_Jinkela_wire_15208)
    );

    bfr new_Jinkela_buffer_2045 (
        .din(new_Jinkela_wire_2986),
        .dout(new_Jinkela_wire_2987)
    );

    bfr new_Jinkela_buffer_12463 (
        .din(new_Jinkela_wire_14964),
        .dout(new_Jinkela_wire_14965)
    );

    bfr new_Jinkela_buffer_15906 (
        .din(new_Jinkela_wire_18938),
        .dout(new_Jinkela_wire_18939)
    );

    bfr new_Jinkela_buffer_1963 (
        .din(new_Jinkela_wire_2884),
        .dout(new_Jinkela_wire_2885)
    );

    bfr new_Jinkela_buffer_12539 (
        .din(new_Jinkela_wire_15046),
        .dout(new_Jinkela_wire_15047)
    );

    bfr new_Jinkela_buffer_16006 (
        .din(new_Jinkela_wire_19086),
        .dout(new_Jinkela_wire_19087)
    );

    bfr new_Jinkela_buffer_12464 (
        .din(new_Jinkela_wire_14965),
        .dout(new_Jinkela_wire_14966)
    );

    spl2 new_Jinkela_splitter_1365 (
        .a(new_Jinkela_wire_18939),
        .b(new_Jinkela_wire_18940),
        .c(new_Jinkela_wire_18941)
    );

    bfr new_Jinkela_buffer_1964 (
        .din(new_Jinkela_wire_2885),
        .dout(new_Jinkela_wire_2886)
    );

    bfr new_Jinkela_buffer_12617 (
        .din(new_Jinkela_wire_15132),
        .dout(new_Jinkela_wire_15133)
    );

    spl2 new_Jinkela_splitter_1395 (
        .a(_0249_),
        .b(new_Jinkela_wire_19118),
        .c(new_Jinkela_wire_19119)
    );

    bfr new_Jinkela_buffer_2046 (
        .din(new_Jinkela_wire_2987),
        .dout(new_Jinkela_wire_2988)
    );

    bfr new_Jinkela_buffer_12465 (
        .din(new_Jinkela_wire_14966),
        .dout(new_Jinkela_wire_14967)
    );

    bfr new_Jinkela_buffer_15962 (
        .din(new_Jinkela_wire_19018),
        .dout(new_Jinkela_wire_19019)
    );

    bfr new_Jinkela_buffer_1965 (
        .din(new_Jinkela_wire_2886),
        .dout(new_Jinkela_wire_2887)
    );

    bfr new_Jinkela_buffer_12540 (
        .din(new_Jinkela_wire_15047),
        .dout(new_Jinkela_wire_15048)
    );

    bfr new_Jinkela_buffer_15963 (
        .din(new_Jinkela_wire_19019),
        .dout(new_Jinkela_wire_19020)
    );

    bfr new_Jinkela_buffer_12466 (
        .din(new_Jinkela_wire_14967),
        .dout(new_Jinkela_wire_14968)
    );

    bfr new_Jinkela_buffer_16007 (
        .din(new_Jinkela_wire_19087),
        .dout(new_Jinkela_wire_19088)
    );

    bfr new_Jinkela_buffer_1966 (
        .din(new_Jinkela_wire_2887),
        .dout(new_Jinkela_wire_2888)
    );

    bfr new_Jinkela_buffer_15964 (
        .din(new_Jinkela_wire_19020),
        .dout(new_Jinkela_wire_19021)
    );

    bfr new_Jinkela_buffer_2181 (
        .din(new_Jinkela_wire_3130),
        .dout(new_Jinkela_wire_3131)
    );

    bfr new_Jinkela_buffer_12873 (
        .din(_0223_),
        .dout(new_Jinkela_wire_15395)
    );

    bfr new_Jinkela_buffer_2047 (
        .din(new_Jinkela_wire_2988),
        .dout(new_Jinkela_wire_2989)
    );

    bfr new_Jinkela_buffer_12467 (
        .din(new_Jinkela_wire_14968),
        .dout(new_Jinkela_wire_14969)
    );

    bfr new_Jinkela_buffer_1967 (
        .din(new_Jinkela_wire_2888),
        .dout(new_Jinkela_wire_2889)
    );

    spl2 new_Jinkela_splitter_1396 (
        .a(_0694_),
        .b(new_Jinkela_wire_19120),
        .c(new_Jinkela_wire_19121)
    );

    bfr new_Jinkela_buffer_12541 (
        .din(new_Jinkela_wire_15048),
        .dout(new_Jinkela_wire_15049)
    );

    bfr new_Jinkela_buffer_15965 (
        .din(new_Jinkela_wire_19021),
        .dout(new_Jinkela_wire_19022)
    );

    bfr new_Jinkela_buffer_12468 (
        .din(new_Jinkela_wire_14969),
        .dout(new_Jinkela_wire_14970)
    );

    bfr new_Jinkela_buffer_16008 (
        .din(new_Jinkela_wire_19088),
        .dout(new_Jinkela_wire_19089)
    );

    bfr new_Jinkela_buffer_1968 (
        .din(new_Jinkela_wire_2889),
        .dout(new_Jinkela_wire_2890)
    );

    bfr new_Jinkela_buffer_12618 (
        .din(new_Jinkela_wire_15133),
        .dout(new_Jinkela_wire_15134)
    );

    bfr new_Jinkela_buffer_15966 (
        .din(new_Jinkela_wire_19022),
        .dout(new_Jinkela_wire_19023)
    );

    bfr new_Jinkela_buffer_2048 (
        .din(new_Jinkela_wire_2989),
        .dout(new_Jinkela_wire_2990)
    );

    bfr new_Jinkela_buffer_12469 (
        .din(new_Jinkela_wire_14970),
        .dout(new_Jinkela_wire_14971)
    );

    spl2 new_Jinkela_splitter_1399 (
        .a(_0911_),
        .b(new_Jinkela_wire_19128),
        .c(new_Jinkela_wire_19129)
    );

    bfr new_Jinkela_buffer_1969 (
        .din(new_Jinkela_wire_2890),
        .dout(new_Jinkela_wire_2891)
    );

    bfr new_Jinkela_buffer_16025 (
        .din(_0978_),
        .dout(new_Jinkela_wire_19122)
    );

    bfr new_Jinkela_buffer_12542 (
        .din(new_Jinkela_wire_15049),
        .dout(new_Jinkela_wire_15050)
    );

    bfr new_Jinkela_buffer_15967 (
        .din(new_Jinkela_wire_19023),
        .dout(new_Jinkela_wire_19024)
    );

    spl2 new_Jinkela_splitter_331 (
        .a(_1322_),
        .b(new_Jinkela_wire_3195),
        .c(new_Jinkela_wire_3196)
    );

    bfr new_Jinkela_buffer_12470 (
        .din(new_Jinkela_wire_14971),
        .dout(new_Jinkela_wire_14972)
    );

    bfr new_Jinkela_buffer_16009 (
        .din(new_Jinkela_wire_19089),
        .dout(new_Jinkela_wire_19090)
    );

    bfr new_Jinkela_buffer_1970 (
        .din(new_Jinkela_wire_2891),
        .dout(new_Jinkela_wire_2892)
    );

    bfr new_Jinkela_buffer_12945 (
        .din(new_net_3960),
        .dout(new_Jinkela_wire_15469)
    );

    bfr new_Jinkela_buffer_15968 (
        .din(new_Jinkela_wire_19024),
        .dout(new_Jinkela_wire_19025)
    );

    bfr new_Jinkela_buffer_2182 (
        .din(new_Jinkela_wire_3131),
        .dout(new_Jinkela_wire_3132)
    );

    bfr new_Jinkela_buffer_12687 (
        .din(new_Jinkela_wire_15208),
        .dout(new_Jinkela_wire_15209)
    );

    bfr new_Jinkela_buffer_2049 (
        .din(new_Jinkela_wire_2990),
        .dout(new_Jinkela_wire_2991)
    );

    bfr new_Jinkela_buffer_12471 (
        .din(new_Jinkela_wire_14972),
        .dout(new_Jinkela_wire_14973)
    );

    bfr new_Jinkela_buffer_1971 (
        .din(new_Jinkela_wire_2892),
        .dout(new_Jinkela_wire_2893)
    );

    spl2 new_Jinkela_splitter_1398 (
        .a(_1818_),
        .b(new_Jinkela_wire_19126),
        .c(new_Jinkela_wire_19127)
    );

    bfr new_Jinkela_buffer_12543 (
        .din(new_Jinkela_wire_15050),
        .dout(new_Jinkela_wire_15051)
    );

    bfr new_Jinkela_buffer_15969 (
        .din(new_Jinkela_wire_19025),
        .dout(new_Jinkela_wire_19026)
    );

    and_bb _3043_ (
        .a(new_Jinkela_wire_10113),
        .b(new_Jinkela_wire_6511),
        .c(_0297_)
    );

    and_ii _1885_ (
        .a(new_Jinkela_wire_9607),
        .b(new_Jinkela_wire_10449),
        .c(_0132_)
    );

    or_bb _3044_ (
        .a(new_Jinkela_wire_11411),
        .b(new_Jinkela_wire_13394),
        .c(_0298_)
    );

    and_ii _3045_ (
        .a(new_Jinkela_wire_8361),
        .b(new_Jinkela_wire_7589),
        .c(_0299_)
    );

    and_bb _3046_ (
        .a(new_Jinkela_wire_8362),
        .b(new_Jinkela_wire_7590),
        .c(_0300_)
    );

    or_bb _3047_ (
        .a(new_Jinkela_wire_21203),
        .b(new_Jinkela_wire_1898),
        .c(_0301_)
    );

    and_ii _3048_ (
        .a(new_Jinkela_wire_17983),
        .b(new_Jinkela_wire_6191),
        .c(_0302_)
    );

    and_bb _3049_ (
        .a(new_Jinkela_wire_17984),
        .b(new_Jinkela_wire_6192),
        .c(_0303_)
    );

    or_bb _3050_ (
        .a(new_Jinkela_wire_7442),
        .b(new_Jinkela_wire_6808),
        .c(_0304_)
    );

    and_ii _3051_ (
        .a(new_Jinkela_wire_14196),
        .b(new_Jinkela_wire_4826),
        .c(_0305_)
    );

    or_bb _3056_ (
        .a(new_Jinkela_wire_3551),
        .b(new_Jinkela_wire_14012),
        .c(_0311_)
    );

    and_ii _3057_ (
        .a(new_Jinkela_wire_17995),
        .b(new_Jinkela_wire_5884),
        .c(_0312_)
    );

    and_bb _3058_ (
        .a(new_Jinkela_wire_17996),
        .b(new_Jinkela_wire_5885),
        .c(_0313_)
    );

    or_bb _3059_ (
        .a(new_Jinkela_wire_18290),
        .b(new_Jinkela_wire_8964),
        .c(_0314_)
    );

    and_ii _3060_ (
        .a(new_Jinkela_wire_4680),
        .b(new_Jinkela_wire_5662),
        .c(_0315_)
    );

    and_bb _3061_ (
        .a(new_Jinkela_wire_4681),
        .b(new_Jinkela_wire_5663),
        .c(_0316_)
    );

    or_bb _3062_ (
        .a(new_Jinkela_wire_21332),
        .b(new_Jinkela_wire_19972),
        .c(_0317_)
    );

    and_ii _3063_ (
        .a(new_Jinkela_wire_2343),
        .b(new_Jinkela_wire_7842),
        .c(_0319_)
    );

    and_bb _3064_ (
        .a(new_Jinkela_wire_2344),
        .b(new_Jinkela_wire_7843),
        .c(_0320_)
    );

    or_bb _3065_ (
        .a(new_Jinkela_wire_21168),
        .b(new_Jinkela_wire_19134),
        .c(_0321_)
    );

    and_bi _3066_ (
        .a(new_Jinkela_wire_9609),
        .b(new_Jinkela_wire_21160),
        .c(_0322_)
    );

    and_bi _3067_ (
        .a(new_Jinkela_wire_21161),
        .b(new_Jinkela_wire_9610),
        .c(_0323_)
    );

    or_bb _3068_ (
        .a(new_Jinkela_wire_15202),
        .b(new_Jinkela_wire_17361),
        .c(new_net_3960)
    );

    or_bb _3069_ (
        .a(new_Jinkela_wire_17362),
        .b(new_Jinkela_wire_19143),
        .c(_0324_)
    );

    and_ii _3070_ (
        .a(new_Jinkela_wire_19973),
        .b(new_Jinkela_wire_8969),
        .c(_0325_)
    );

    and_bb _3071_ (
        .a(new_Jinkela_wire_67),
        .b(new_Jinkela_wire_660),
        .c(_0326_)
    );

    and_ii _3072_ (
        .a(new_Jinkela_wire_14013),
        .b(new_Jinkela_wire_8024),
        .c(_0327_)
    );

    and_bb _3073_ (
        .a(new_Jinkela_wire_483),
        .b(new_Jinkela_wire_526),
        .c(_0329_)
    );

    and_ii _3074_ (
        .a(new_Jinkela_wire_6809),
        .b(new_Jinkela_wire_1903),
        .c(_0330_)
    );

    and_bb _3075_ (
        .a(new_Jinkela_wire_361),
        .b(new_Jinkela_wire_135),
        .c(_0331_)
    );

    and_ii _3076_ (
        .a(new_Jinkela_wire_13395),
        .b(new_Jinkela_wire_13729),
        .c(_0332_)
    );

    and_bb _3077_ (
        .a(new_Jinkela_wire_684),
        .b(new_Jinkela_wire_204),
        .c(_0333_)
    );

    and_ii _3078_ (
        .a(new_Jinkela_wire_17548),
        .b(new_Jinkela_wire_14271),
        .c(_0334_)
    );

    and_bb _3079_ (
        .a(new_Jinkela_wire_577),
        .b(new_Jinkela_wire_500),
        .c(_0335_)
    );

    and_ii _3080_ (
        .a(new_Jinkela_wire_13150),
        .b(new_Jinkela_wire_16001),
        .c(_0336_)
    );

    and_bb _3081_ (
        .a(new_Jinkela_wire_122),
        .b(new_Jinkela_wire_33),
        .c(_0337_)
    );

    and_ii _3082_ (
        .a(new_Jinkela_wire_21165),
        .b(new_Jinkela_wire_4701),
        .c(_0338_)
    );

    and_bb _3083_ (
        .a(new_Jinkela_wire_180),
        .b(new_Jinkela_wire_6),
        .c(_0340_)
    );

    and_ii _3084_ (
        .a(new_Jinkela_wire_10262),
        .b(new_Jinkela_wire_11427),
        .c(_0341_)
    );

    and_bb _3085_ (
        .a(new_Jinkela_wire_377),
        .b(new_Jinkela_wire_462),
        .c(_0342_)
    );

    and_ii _3086_ (
        .a(new_Jinkela_wire_2136),
        .b(new_Jinkela_wire_2142),
        .c(_0343_)
    );

    and_bb _3087_ (
        .a(new_Jinkela_wire_397),
        .b(new_Jinkela_wire_250),
        .c(_0344_)
    );

    bfr new_Jinkela_buffer_12472 (
        .din(new_Jinkela_wire_14973),
        .dout(new_Jinkela_wire_14974)
    );

    bfr new_Jinkela_buffer_12619 (
        .din(new_Jinkela_wire_15134),
        .dout(new_Jinkela_wire_15135)
    );

    bfr new_Jinkela_buffer_12473 (
        .din(new_Jinkela_wire_14974),
        .dout(new_Jinkela_wire_14975)
    );

    bfr new_Jinkela_buffer_12544 (
        .din(new_Jinkela_wire_15051),
        .dout(new_Jinkela_wire_15052)
    );

    bfr new_Jinkela_buffer_12474 (
        .din(new_Jinkela_wire_14975),
        .dout(new_Jinkela_wire_14976)
    );

    bfr new_Jinkela_buffer_12858 (
        .din(new_Jinkela_wire_15379),
        .dout(new_Jinkela_wire_15380)
    );

    bfr new_Jinkela_buffer_12475 (
        .din(new_Jinkela_wire_14976),
        .dout(new_Jinkela_wire_14977)
    );

    bfr new_Jinkela_buffer_12545 (
        .din(new_Jinkela_wire_15052),
        .dout(new_Jinkela_wire_15053)
    );

    bfr new_Jinkela_buffer_12476 (
        .din(new_Jinkela_wire_14977),
        .dout(new_Jinkela_wire_14978)
    );

    bfr new_Jinkela_buffer_12620 (
        .din(new_Jinkela_wire_15135),
        .dout(new_Jinkela_wire_15136)
    );

    bfr new_Jinkela_buffer_12477 (
        .din(new_Jinkela_wire_14978),
        .dout(new_Jinkela_wire_14979)
    );

    bfr new_Jinkela_buffer_12546 (
        .din(new_Jinkela_wire_15053),
        .dout(new_Jinkela_wire_15054)
    );

    bfr new_Jinkela_buffer_12478 (
        .din(new_Jinkela_wire_14979),
        .dout(new_Jinkela_wire_14980)
    );

    bfr new_Jinkela_buffer_12688 (
        .din(new_Jinkela_wire_15209),
        .dout(new_Jinkela_wire_15210)
    );

    bfr new_Jinkela_buffer_12479 (
        .din(new_Jinkela_wire_14980),
        .dout(new_Jinkela_wire_14981)
    );

    bfr new_Jinkela_buffer_12547 (
        .din(new_Jinkela_wire_15054),
        .dout(new_Jinkela_wire_15055)
    );

    bfr new_Jinkela_buffer_12480 (
        .din(new_Jinkela_wire_14981),
        .dout(new_Jinkela_wire_14982)
    );

    bfr new_Jinkela_buffer_12621 (
        .din(new_Jinkela_wire_15136),
        .dout(new_Jinkela_wire_15137)
    );

    bfr new_Jinkela_buffer_12481 (
        .din(new_Jinkela_wire_14982),
        .dout(new_Jinkela_wire_14983)
    );

    bfr new_Jinkela_buffer_12548 (
        .din(new_Jinkela_wire_15055),
        .dout(new_Jinkela_wire_15056)
    );

    bfr new_Jinkela_buffer_12482 (
        .din(new_Jinkela_wire_14983),
        .dout(new_Jinkela_wire_14984)
    );

    bfr new_Jinkela_buffer_12483 (
        .din(new_Jinkela_wire_14984),
        .dout(new_Jinkela_wire_14985)
    );

    bfr new_Jinkela_buffer_12549 (
        .din(new_Jinkela_wire_15056),
        .dout(new_Jinkela_wire_15057)
    );

    bfr new_Jinkela_buffer_12484 (
        .din(new_Jinkela_wire_14985),
        .dout(new_Jinkela_wire_14986)
    );

    bfr new_Jinkela_buffer_12622 (
        .din(new_Jinkela_wire_15137),
        .dout(new_Jinkela_wire_15138)
    );

    bfr new_Jinkela_buffer_12485 (
        .din(new_Jinkela_wire_14986),
        .dout(new_Jinkela_wire_14987)
    );

    bfr new_Jinkela_buffer_12550 (
        .din(new_Jinkela_wire_15057),
        .dout(new_Jinkela_wire_15058)
    );

    spl2 new_Jinkela_splitter_1100 (
        .a(new_Jinkela_wire_14987),
        .b(new_Jinkela_wire_14988),
        .c(new_Jinkela_wire_14989)
    );

    bfr new_Jinkela_buffer_12551 (
        .din(new_Jinkela_wire_15058),
        .dout(new_Jinkela_wire_15059)
    );

    bfr new_Jinkela_buffer_12689 (
        .din(new_Jinkela_wire_15210),
        .dout(new_Jinkela_wire_15211)
    );

    bfr new_Jinkela_buffer_12623 (
        .din(new_Jinkela_wire_15138),
        .dout(new_Jinkela_wire_15139)
    );

    bfr new_Jinkela_buffer_12552 (
        .din(new_Jinkela_wire_15059),
        .dout(new_Jinkela_wire_15060)
    );

    bfr new_Jinkela_buffer_12859 (
        .din(new_Jinkela_wire_15380),
        .dout(new_Jinkela_wire_15381)
    );

    bfr new_Jinkela_buffer_12553 (
        .din(new_Jinkela_wire_15060),
        .dout(new_Jinkela_wire_15061)
    );

    bfr new_Jinkela_buffer_12624 (
        .din(new_Jinkela_wire_15139),
        .dout(new_Jinkela_wire_15140)
    );

    bfr new_Jinkela_buffer_12554 (
        .din(new_Jinkela_wire_15061),
        .dout(new_Jinkela_wire_15062)
    );

    bfr new_Jinkela_buffer_12690 (
        .din(new_Jinkela_wire_15211),
        .dout(new_Jinkela_wire_15212)
    );

    bfr new_Jinkela_buffer_12555 (
        .din(new_Jinkela_wire_15062),
        .dout(new_Jinkela_wire_15063)
    );

    bfr new_Jinkela_buffer_12625 (
        .din(new_Jinkela_wire_15140),
        .dout(new_Jinkela_wire_15141)
    );

    bfr new_Jinkela_buffer_12556 (
        .din(new_Jinkela_wire_15063),
        .dout(new_Jinkela_wire_15064)
    );

    spl2 new_Jinkela_splitter_1111 (
        .a(_0553_),
        .b(new_Jinkela_wire_15517),
        .c(new_Jinkela_wire_15518)
    );

    bfr new_Jinkela_buffer_5559 (
        .din(new_Jinkela_wire_7096),
        .dout(new_Jinkela_wire_7097)
    );

    bfr new_Jinkela_buffer_1972 (
        .din(new_Jinkela_wire_2893),
        .dout(new_Jinkela_wire_2894)
    );

    bfr new_Jinkela_buffer_5612 (
        .din(new_Jinkela_wire_7157),
        .dout(new_Jinkela_wire_7158)
    );

    bfr new_Jinkela_buffer_2277 (
        .din(_1634_),
        .dout(new_Jinkela_wire_3257)
    );

    bfr new_Jinkela_buffer_2050 (
        .din(new_Jinkela_wire_2991),
        .dout(new_Jinkela_wire_2992)
    );

    bfr new_Jinkela_buffer_5560 (
        .din(new_Jinkela_wire_7097),
        .dout(new_Jinkela_wire_7098)
    );

    bfr new_Jinkela_buffer_1973 (
        .din(new_Jinkela_wire_2894),
        .dout(new_Jinkela_wire_2895)
    );

    bfr new_Jinkela_buffer_5637 (
        .din(new_Jinkela_wire_7190),
        .dout(new_Jinkela_wire_7191)
    );

    bfr new_Jinkela_buffer_5561 (
        .din(new_Jinkela_wire_7098),
        .dout(new_Jinkela_wire_7099)
    );

    bfr new_Jinkela_buffer_1974 (
        .din(new_Jinkela_wire_2895),
        .dout(new_Jinkela_wire_2896)
    );

    bfr new_Jinkela_buffer_5613 (
        .din(new_Jinkela_wire_7158),
        .dout(new_Jinkela_wire_7159)
    );

    bfr new_Jinkela_buffer_2183 (
        .din(new_Jinkela_wire_3132),
        .dout(new_Jinkela_wire_3133)
    );

    bfr new_Jinkela_buffer_2051 (
        .din(new_Jinkela_wire_2992),
        .dout(new_Jinkela_wire_2993)
    );

    bfr new_Jinkela_buffer_5562 (
        .din(new_Jinkela_wire_7099),
        .dout(new_Jinkela_wire_7100)
    );

    bfr new_Jinkela_buffer_1975 (
        .din(new_Jinkela_wire_2896),
        .dout(new_Jinkela_wire_2897)
    );

    spl2 new_Jinkela_splitter_628 (
        .a(_0150_),
        .b(new_Jinkela_wire_7270),
        .c(new_Jinkela_wire_7271)
    );

    bfr new_Jinkela_buffer_5563 (
        .din(new_Jinkela_wire_7100),
        .dout(new_Jinkela_wire_7101)
    );

    bfr new_Jinkela_buffer_1976 (
        .din(new_Jinkela_wire_2897),
        .dout(new_Jinkela_wire_2898)
    );

    bfr new_Jinkela_buffer_5614 (
        .din(new_Jinkela_wire_7159),
        .dout(new_Jinkela_wire_7160)
    );

    bfr new_Jinkela_buffer_2052 (
        .din(new_Jinkela_wire_2993),
        .dout(new_Jinkela_wire_2994)
    );

    bfr new_Jinkela_buffer_5564 (
        .din(new_Jinkela_wire_7101),
        .dout(new_Jinkela_wire_7102)
    );

    bfr new_Jinkela_buffer_1977 (
        .din(new_Jinkela_wire_2898),
        .dout(new_Jinkela_wire_2899)
    );

    bfr new_Jinkela_buffer_5638 (
        .din(new_Jinkela_wire_7191),
        .dout(new_Jinkela_wire_7192)
    );

    spl2 new_Jinkela_splitter_339 (
        .a(_0472_),
        .b(new_Jinkela_wire_3258),
        .c(new_Jinkela_wire_3259)
    );

    bfr new_Jinkela_buffer_5565 (
        .din(new_Jinkela_wire_7102),
        .dout(new_Jinkela_wire_7103)
    );

    bfr new_Jinkela_buffer_1978 (
        .din(new_Jinkela_wire_2899),
        .dout(new_Jinkela_wire_2900)
    );

    bfr new_Jinkela_buffer_5615 (
        .din(new_Jinkela_wire_7160),
        .dout(new_Jinkela_wire_7161)
    );

    bfr new_Jinkela_buffer_2184 (
        .din(new_Jinkela_wire_3133),
        .dout(new_Jinkela_wire_3134)
    );

    bfr new_Jinkela_buffer_2053 (
        .din(new_Jinkela_wire_2994),
        .dout(new_Jinkela_wire_2995)
    );

    bfr new_Jinkela_buffer_5566 (
        .din(new_Jinkela_wire_7103),
        .dout(new_Jinkela_wire_7104)
    );

    bfr new_Jinkela_buffer_1979 (
        .din(new_Jinkela_wire_2900),
        .dout(new_Jinkela_wire_2901)
    );

    bfr new_Jinkela_buffer_5712 (
        .din(_1795_),
        .dout(new_Jinkela_wire_7272)
    );

    bfr new_Jinkela_buffer_5567 (
        .din(new_Jinkela_wire_7104),
        .dout(new_Jinkela_wire_7105)
    );

    bfr new_Jinkela_buffer_1980 (
        .din(new_Jinkela_wire_2901),
        .dout(new_Jinkela_wire_2902)
    );

    bfr new_Jinkela_buffer_5616 (
        .din(new_Jinkela_wire_7161),
        .dout(new_Jinkela_wire_7162)
    );

    bfr new_Jinkela_buffer_2240 (
        .din(new_Jinkela_wire_3205),
        .dout(new_Jinkela_wire_3206)
    );

    bfr new_Jinkela_buffer_2054 (
        .din(new_Jinkela_wire_2995),
        .dout(new_Jinkela_wire_2996)
    );

    bfr new_Jinkela_buffer_5568 (
        .din(new_Jinkela_wire_7105),
        .dout(new_Jinkela_wire_7106)
    );

    bfr new_Jinkela_buffer_1981 (
        .din(new_Jinkela_wire_2902),
        .dout(new_Jinkela_wire_2903)
    );

    bfr new_Jinkela_buffer_5639 (
        .din(new_Jinkela_wire_7192),
        .dout(new_Jinkela_wire_7193)
    );

    bfr new_Jinkela_buffer_5569 (
        .din(new_Jinkela_wire_7106),
        .dout(new_Jinkela_wire_7107)
    );

    bfr new_Jinkela_buffer_1982 (
        .din(new_Jinkela_wire_2903),
        .dout(new_Jinkela_wire_2904)
    );

    bfr new_Jinkela_buffer_5617 (
        .din(new_Jinkela_wire_7162),
        .dout(new_Jinkela_wire_7163)
    );

    bfr new_Jinkela_buffer_2185 (
        .din(new_Jinkela_wire_3134),
        .dout(new_Jinkela_wire_3135)
    );

    bfr new_Jinkela_buffer_2055 (
        .din(new_Jinkela_wire_2996),
        .dout(new_Jinkela_wire_2997)
    );

    bfr new_Jinkela_buffer_5570 (
        .din(new_Jinkela_wire_7107),
        .dout(new_Jinkela_wire_7108)
    );

    bfr new_Jinkela_buffer_1983 (
        .din(new_Jinkela_wire_2904),
        .dout(new_Jinkela_wire_2905)
    );

    bfr new_Jinkela_buffer_5708 (
        .din(new_Jinkela_wire_7265),
        .dout(new_Jinkela_wire_7266)
    );

    bfr new_Jinkela_buffer_5571 (
        .din(new_Jinkela_wire_7108),
        .dout(new_Jinkela_wire_7109)
    );

    bfr new_Jinkela_buffer_1984 (
        .din(new_Jinkela_wire_2905),
        .dout(new_Jinkela_wire_2906)
    );

    bfr new_Jinkela_buffer_5618 (
        .din(new_Jinkela_wire_7163),
        .dout(new_Jinkela_wire_7164)
    );

    bfr new_Jinkela_buffer_2274 (
        .din(new_Jinkela_wire_3249),
        .dout(new_Jinkela_wire_3250)
    );

    bfr new_Jinkela_buffer_2056 (
        .din(new_Jinkela_wire_2997),
        .dout(new_Jinkela_wire_2998)
    );

    bfr new_Jinkela_buffer_5572 (
        .din(new_Jinkela_wire_7109),
        .dout(new_Jinkela_wire_7110)
    );

    bfr new_Jinkela_buffer_1985 (
        .din(new_Jinkela_wire_2906),
        .dout(new_Jinkela_wire_2907)
    );

    bfr new_Jinkela_buffer_5640 (
        .din(new_Jinkela_wire_7193),
        .dout(new_Jinkela_wire_7194)
    );

    bfr new_Jinkela_buffer_5573 (
        .din(new_Jinkela_wire_7110),
        .dout(new_Jinkela_wire_7111)
    );

    bfr new_Jinkela_buffer_1986 (
        .din(new_Jinkela_wire_2907),
        .dout(new_Jinkela_wire_2908)
    );

    bfr new_Jinkela_buffer_5619 (
        .din(new_Jinkela_wire_7164),
        .dout(new_Jinkela_wire_7165)
    );

    bfr new_Jinkela_buffer_2186 (
        .din(new_Jinkela_wire_3135),
        .dout(new_Jinkela_wire_3136)
    );

    bfr new_Jinkela_buffer_2057 (
        .din(new_Jinkela_wire_2998),
        .dout(new_Jinkela_wire_2999)
    );

    bfr new_Jinkela_buffer_5574 (
        .din(new_Jinkela_wire_7111),
        .dout(new_Jinkela_wire_7112)
    );

    bfr new_Jinkela_buffer_1987 (
        .din(new_Jinkela_wire_2908),
        .dout(new_Jinkela_wire_2909)
    );

    spl2 new_Jinkela_splitter_629 (
        .a(_1187_),
        .b(new_Jinkela_wire_7273),
        .c(new_Jinkela_wire_7274)
    );

    bfr new_Jinkela_buffer_5575 (
        .din(new_Jinkela_wire_7112),
        .dout(new_Jinkela_wire_7113)
    );

    bfr new_Jinkela_buffer_1988 (
        .din(new_Jinkela_wire_2909),
        .dout(new_Jinkela_wire_2910)
    );

    bfr new_Jinkela_buffer_5620 (
        .din(new_Jinkela_wire_7165),
        .dout(new_Jinkela_wire_7166)
    );

    bfr new_Jinkela_buffer_2241 (
        .din(new_Jinkela_wire_3206),
        .dout(new_Jinkela_wire_3207)
    );

    bfr new_Jinkela_buffer_2058 (
        .din(new_Jinkela_wire_2999),
        .dout(new_Jinkela_wire_3000)
    );

    bfr new_Jinkela_buffer_5576 (
        .din(new_Jinkela_wire_7113),
        .dout(new_Jinkela_wire_7114)
    );

    bfr new_Jinkela_buffer_1989 (
        .din(new_Jinkela_wire_2910),
        .dout(new_Jinkela_wire_2911)
    );

    bfr new_Jinkela_buffer_5641 (
        .din(new_Jinkela_wire_7194),
        .dout(new_Jinkela_wire_7195)
    );

    bfr new_Jinkela_buffer_5577 (
        .din(new_Jinkela_wire_7114),
        .dout(new_Jinkela_wire_7115)
    );

    bfr new_Jinkela_buffer_1990 (
        .din(new_Jinkela_wire_2911),
        .dout(new_Jinkela_wire_2912)
    );

    bfr new_Jinkela_buffer_5621 (
        .din(new_Jinkela_wire_7166),
        .dout(new_Jinkela_wire_7167)
    );

    bfr new_Jinkela_buffer_2187 (
        .din(new_Jinkela_wire_3136),
        .dout(new_Jinkela_wire_3137)
    );

    bfr new_Jinkela_buffer_2059 (
        .din(new_Jinkela_wire_3000),
        .dout(new_Jinkela_wire_3001)
    );

    bfr new_Jinkela_buffer_5578 (
        .din(new_Jinkela_wire_7115),
        .dout(new_Jinkela_wire_7116)
    );

    bfr new_Jinkela_buffer_1991 (
        .din(new_Jinkela_wire_2912),
        .dout(new_Jinkela_wire_2913)
    );

    bfr new_Jinkela_buffer_5709 (
        .din(new_Jinkela_wire_7266),
        .dout(new_Jinkela_wire_7267)
    );

    bfr new_Jinkela_buffer_5579 (
        .din(new_Jinkela_wire_7116),
        .dout(new_Jinkela_wire_7117)
    );

    bfr new_Jinkela_buffer_1992 (
        .din(new_Jinkela_wire_2913),
        .dout(new_Jinkela_wire_2914)
    );

    bfr new_Jinkela_buffer_5622 (
        .din(new_Jinkela_wire_7167),
        .dout(new_Jinkela_wire_7168)
    );

    bfr new_Jinkela_buffer_9124 (
        .din(new_Jinkela_wire_11143),
        .dout(new_Jinkela_wire_11144)
    );

    bfr new_Jinkela_buffer_9046 (
        .din(new_Jinkela_wire_11061),
        .dout(new_Jinkela_wire_11062)
    );

    bfr new_Jinkela_buffer_9208 (
        .din(new_Jinkela_wire_11231),
        .dout(new_Jinkela_wire_11232)
    );

    bfr new_Jinkela_buffer_9047 (
        .din(new_Jinkela_wire_11062),
        .dout(new_Jinkela_wire_11063)
    );

    bfr new_Jinkela_buffer_9125 (
        .din(new_Jinkela_wire_11144),
        .dout(new_Jinkela_wire_11145)
    );

    bfr new_Jinkela_buffer_9048 (
        .din(new_Jinkela_wire_11063),
        .dout(new_Jinkela_wire_11064)
    );

    spl2 new_Jinkela_splitter_862 (
        .a(_1248_),
        .b(new_Jinkela_wire_11342),
        .c(new_Jinkela_wire_11343)
    );

    bfr new_Jinkela_buffer_9049 (
        .din(new_Jinkela_wire_11064),
        .dout(new_Jinkela_wire_11065)
    );

    bfr new_Jinkela_buffer_9126 (
        .din(new_Jinkela_wire_11145),
        .dout(new_Jinkela_wire_11146)
    );

    bfr new_Jinkela_buffer_9050 (
        .din(new_Jinkela_wire_11065),
        .dout(new_Jinkela_wire_11066)
    );

    bfr new_Jinkela_buffer_9209 (
        .din(new_Jinkela_wire_11232),
        .dout(new_Jinkela_wire_11233)
    );

    bfr new_Jinkela_buffer_9051 (
        .din(new_Jinkela_wire_11066),
        .dout(new_Jinkela_wire_11067)
    );

    bfr new_Jinkela_buffer_9127 (
        .din(new_Jinkela_wire_11146),
        .dout(new_Jinkela_wire_11147)
    );

    bfr new_Jinkela_buffer_9052 (
        .din(new_Jinkela_wire_11067),
        .dout(new_Jinkela_wire_11068)
    );

    bfr new_Jinkela_buffer_9212 (
        .din(new_Jinkela_wire_11235),
        .dout(new_Jinkela_wire_11236)
    );

    bfr new_Jinkela_buffer_9053 (
        .din(new_Jinkela_wire_11068),
        .dout(new_Jinkela_wire_11069)
    );

    bfr new_Jinkela_buffer_9128 (
        .din(new_Jinkela_wire_11147),
        .dout(new_Jinkela_wire_11148)
    );

    bfr new_Jinkela_buffer_9054 (
        .din(new_Jinkela_wire_11069),
        .dout(new_Jinkela_wire_11070)
    );

    spl2 new_Jinkela_splitter_863 (
        .a(_0468_),
        .b(new_Jinkela_wire_11344),
        .c(new_Jinkela_wire_11345)
    );

    bfr new_Jinkela_buffer_9055 (
        .din(new_Jinkela_wire_11070),
        .dout(new_Jinkela_wire_11071)
    );

    bfr new_Jinkela_buffer_9129 (
        .din(new_Jinkela_wire_11148),
        .dout(new_Jinkela_wire_11149)
    );

    bfr new_Jinkela_buffer_9056 (
        .din(new_Jinkela_wire_11071),
        .dout(new_Jinkela_wire_11072)
    );

    bfr new_Jinkela_buffer_9213 (
        .din(new_Jinkela_wire_11236),
        .dout(new_Jinkela_wire_11237)
    );

    bfr new_Jinkela_buffer_9057 (
        .din(new_Jinkela_wire_11072),
        .dout(new_Jinkela_wire_11073)
    );

    bfr new_Jinkela_buffer_9130 (
        .din(new_Jinkela_wire_11149),
        .dout(new_Jinkela_wire_11150)
    );

    bfr new_Jinkela_buffer_9058 (
        .din(new_Jinkela_wire_11073),
        .dout(new_Jinkela_wire_11074)
    );

    bfr new_Jinkela_buffer_9316 (
        .din(new_Jinkela_wire_11345),
        .dout(new_Jinkela_wire_11346)
    );

    bfr new_Jinkela_buffer_9059 (
        .din(new_Jinkela_wire_11074),
        .dout(new_Jinkela_wire_11075)
    );

    bfr new_Jinkela_buffer_9131 (
        .din(new_Jinkela_wire_11150),
        .dout(new_Jinkela_wire_11151)
    );

    bfr new_Jinkela_buffer_9060 (
        .din(new_Jinkela_wire_11075),
        .dout(new_Jinkela_wire_11076)
    );

    bfr new_Jinkela_buffer_9214 (
        .din(new_Jinkela_wire_11237),
        .dout(new_Jinkela_wire_11238)
    );

    bfr new_Jinkela_buffer_9061 (
        .din(new_Jinkela_wire_11076),
        .dout(new_Jinkela_wire_11077)
    );

    bfr new_Jinkela_buffer_9132 (
        .din(new_Jinkela_wire_11151),
        .dout(new_Jinkela_wire_11152)
    );

    bfr new_Jinkela_buffer_9062 (
        .din(new_Jinkela_wire_11077),
        .dout(new_Jinkela_wire_11078)
    );

    bfr new_Jinkela_buffer_9320 (
        .din(_0452_),
        .dout(new_Jinkela_wire_11350)
    );

    bfr new_Jinkela_buffer_9063 (
        .din(new_Jinkela_wire_11078),
        .dout(new_Jinkela_wire_11079)
    );

    bfr new_Jinkela_buffer_9133 (
        .din(new_Jinkela_wire_11152),
        .dout(new_Jinkela_wire_11153)
    );

    bfr new_Jinkela_buffer_9064 (
        .din(new_Jinkela_wire_11079),
        .dout(new_Jinkela_wire_11080)
    );

    bfr new_Jinkela_buffer_9215 (
        .din(new_Jinkela_wire_11238),
        .dout(new_Jinkela_wire_11239)
    );

    bfr new_Jinkela_buffer_9065 (
        .din(new_Jinkela_wire_11080),
        .dout(new_Jinkela_wire_11081)
    );

    bfr new_Jinkela_buffer_9134 (
        .din(new_Jinkela_wire_11153),
        .dout(new_Jinkela_wire_11154)
    );

    bfr new_Jinkela_buffer_9066 (
        .din(new_Jinkela_wire_11081),
        .dout(new_Jinkela_wire_11082)
    );

    bfr new_Jinkela_buffer_2060 (
        .din(new_Jinkela_wire_3001),
        .dout(new_Jinkela_wire_3002)
    );

    bfr new_Jinkela_buffer_1993 (
        .din(new_Jinkela_wire_2914),
        .dout(new_Jinkela_wire_2915)
    );

    bfr new_Jinkela_buffer_1994 (
        .din(new_Jinkela_wire_2915),
        .dout(new_Jinkela_wire_2916)
    );

    bfr new_Jinkela_buffer_2188 (
        .din(new_Jinkela_wire_3137),
        .dout(new_Jinkela_wire_3138)
    );

    bfr new_Jinkela_buffer_2061 (
        .din(new_Jinkela_wire_3002),
        .dout(new_Jinkela_wire_3003)
    );

    bfr new_Jinkela_buffer_1995 (
        .din(new_Jinkela_wire_2916),
        .dout(new_Jinkela_wire_2917)
    );

    bfr new_Jinkela_buffer_1996 (
        .din(new_Jinkela_wire_2917),
        .dout(new_Jinkela_wire_2918)
    );

    bfr new_Jinkela_buffer_2062 (
        .din(new_Jinkela_wire_3003),
        .dout(new_Jinkela_wire_3004)
    );

    bfr new_Jinkela_buffer_1997 (
        .din(new_Jinkela_wire_2918),
        .dout(new_Jinkela_wire_2919)
    );

    spl2 new_Jinkela_splitter_334 (
        .a(_0103_),
        .b(new_Jinkela_wire_3243),
        .c(new_Jinkela_wire_3244)
    );

    bfr new_Jinkela_buffer_1998 (
        .din(new_Jinkela_wire_2919),
        .dout(new_Jinkela_wire_2920)
    );

    bfr new_Jinkela_buffer_2189 (
        .din(new_Jinkela_wire_3138),
        .dout(new_Jinkela_wire_3139)
    );

    bfr new_Jinkela_buffer_2063 (
        .din(new_Jinkela_wire_3004),
        .dout(new_Jinkela_wire_3005)
    );

    bfr new_Jinkela_buffer_1999 (
        .din(new_Jinkela_wire_2920),
        .dout(new_Jinkela_wire_2921)
    );

    bfr new_Jinkela_buffer_2000 (
        .din(new_Jinkela_wire_2921),
        .dout(new_Jinkela_wire_2922)
    );

    bfr new_Jinkela_buffer_2232 (
        .din(new_Jinkela_wire_3197),
        .dout(new_Jinkela_wire_3198)
    );

    bfr new_Jinkela_buffer_2064 (
        .din(new_Jinkela_wire_3005),
        .dout(new_Jinkela_wire_3006)
    );

    bfr new_Jinkela_buffer_2001 (
        .din(new_Jinkela_wire_2922),
        .dout(new_Jinkela_wire_2923)
    );

    bfr new_Jinkela_buffer_2002 (
        .din(new_Jinkela_wire_2923),
        .dout(new_Jinkela_wire_2924)
    );

    bfr new_Jinkela_buffer_2190 (
        .din(new_Jinkela_wire_3139),
        .dout(new_Jinkela_wire_3140)
    );

    bfr new_Jinkela_buffer_2065 (
        .din(new_Jinkela_wire_3006),
        .dout(new_Jinkela_wire_3007)
    );

    bfr new_Jinkela_buffer_2003 (
        .din(new_Jinkela_wire_2924),
        .dout(new_Jinkela_wire_2925)
    );

    bfr new_Jinkela_buffer_2004 (
        .din(new_Jinkela_wire_2925),
        .dout(new_Jinkela_wire_2926)
    );

    bfr new_Jinkela_buffer_2066 (
        .din(new_Jinkela_wire_3007),
        .dout(new_Jinkela_wire_3008)
    );

    bfr new_Jinkela_buffer_2005 (
        .din(new_Jinkela_wire_2926),
        .dout(new_Jinkela_wire_2927)
    );

    spl2 new_Jinkela_splitter_335 (
        .a(_0950_),
        .b(new_Jinkela_wire_3245),
        .c(new_Jinkela_wire_3246)
    );

    bfr new_Jinkela_buffer_2006 (
        .din(new_Jinkela_wire_2927),
        .dout(new_Jinkela_wire_2928)
    );

    bfr new_Jinkela_buffer_2191 (
        .din(new_Jinkela_wire_3140),
        .dout(new_Jinkela_wire_3141)
    );

    bfr new_Jinkela_buffer_2067 (
        .din(new_Jinkela_wire_3008),
        .dout(new_Jinkela_wire_3009)
    );

    bfr new_Jinkela_buffer_2007 (
        .din(new_Jinkela_wire_2928),
        .dout(new_Jinkela_wire_2929)
    );

    bfr new_Jinkela_buffer_2008 (
        .din(new_Jinkela_wire_2929),
        .dout(new_Jinkela_wire_2930)
    );

    bfr new_Jinkela_buffer_2233 (
        .din(new_Jinkela_wire_3198),
        .dout(new_Jinkela_wire_3199)
    );

    bfr new_Jinkela_buffer_2068 (
        .din(new_Jinkela_wire_3009),
        .dout(new_Jinkela_wire_3010)
    );

    bfr new_Jinkela_buffer_2009 (
        .din(new_Jinkela_wire_2930),
        .dout(new_Jinkela_wire_2931)
    );

    spl2 new_Jinkela_splitter_310 (
        .a(new_Jinkela_wire_2931),
        .b(new_Jinkela_wire_2932),
        .c(new_Jinkela_wire_2933)
    );

    bfr new_Jinkela_buffer_2192 (
        .din(new_Jinkela_wire_3141),
        .dout(new_Jinkela_wire_3142)
    );

    bfr new_Jinkela_buffer_2069 (
        .din(new_Jinkela_wire_3010),
        .dout(new_Jinkela_wire_3011)
    );

    bfr new_Jinkela_buffer_2272 (
        .din(new_Jinkela_wire_3239),
        .dout(new_Jinkela_wire_3240)
    );

    bfr new_Jinkela_buffer_2070 (
        .din(new_Jinkela_wire_3011),
        .dout(new_Jinkela_wire_3012)
    );

    bfr new_Jinkela_buffer_2193 (
        .din(new_Jinkela_wire_3142),
        .dout(new_Jinkela_wire_3143)
    );

    bfr new_Jinkela_buffer_2071 (
        .din(new_Jinkela_wire_3012),
        .dout(new_Jinkela_wire_3013)
    );

    bfr new_Jinkela_buffer_2271 (
        .din(_1832_),
        .dout(new_Jinkela_wire_3239)
    );

    and_ii _3088_ (
        .a(new_Jinkela_wire_2654),
        .b(new_Jinkela_wire_16699),
        .c(_0345_)
    );

    bfr new_Jinkela_buffer_5580 (
        .din(new_Jinkela_wire_7117),
        .dout(new_Jinkela_wire_7118)
    );

    bfr new_Jinkela_buffer_16010 (
        .din(new_Jinkela_wire_19090),
        .dout(new_Jinkela_wire_19091)
    );

    and_bb _3089_ (
        .a(new_Jinkela_wire_161),
        .b(new_Jinkela_wire_298),
        .c(_0346_)
    );

    bfr new_Jinkela_buffer_5642 (
        .din(new_Jinkela_wire_7195),
        .dout(new_Jinkela_wire_7196)
    );

    bfr new_Jinkela_buffer_15970 (
        .din(new_Jinkela_wire_19026),
        .dout(new_Jinkela_wire_19027)
    );

    and_ii _3090_ (
        .a(new_Jinkela_wire_19119),
        .b(new_Jinkela_wire_2940),
        .c(_0347_)
    );

    bfr new_Jinkela_buffer_5581 (
        .din(new_Jinkela_wire_7118),
        .dout(new_Jinkela_wire_7119)
    );

    bfr new_Jinkela_buffer_16026 (
        .din(new_Jinkela_wire_19122),
        .dout(new_Jinkela_wire_19123)
    );

    and_bb _3091_ (
        .a(new_Jinkela_wire_608),
        .b(new_Jinkela_wire_48),
        .c(_0348_)
    );

    bfr new_Jinkela_buffer_5623 (
        .din(new_Jinkela_wire_7168),
        .dout(new_Jinkela_wire_7169)
    );

    bfr new_Jinkela_buffer_15971 (
        .din(new_Jinkela_wire_19027),
        .dout(new_Jinkela_wire_19028)
    );

    and_bb _3092_ (
        .a(new_Jinkela_wire_427),
        .b(new_Jinkela_wire_641),
        .c(_0349_)
    );

    bfr new_Jinkela_buffer_5582 (
        .din(new_Jinkela_wire_7119),
        .dout(new_Jinkela_wire_7120)
    );

    bfr new_Jinkela_buffer_16011 (
        .din(new_Jinkela_wire_19091),
        .dout(new_Jinkela_wire_19092)
    );

    and_ii _3093_ (
        .a(new_Jinkela_wire_8587),
        .b(new_Jinkela_wire_10750),
        .c(_0351_)
    );

    spl2 new_Jinkela_splitter_630 (
        .a(_0230_),
        .b(new_Jinkela_wire_7275),
        .c(new_Jinkela_wire_7276)
    );

    bfr new_Jinkela_buffer_15972 (
        .din(new_Jinkela_wire_19028),
        .dout(new_Jinkela_wire_19029)
    );

    and_ii _3094_ (
        .a(new_Jinkela_wire_20355),
        .b(new_Jinkela_wire_18831),
        .c(_0352_)
    );

    bfr new_Jinkela_buffer_5583 (
        .din(new_Jinkela_wire_7120),
        .dout(new_Jinkela_wire_7121)
    );

    and_bb _3095_ (
        .a(new_Jinkela_wire_20356),
        .b(new_Jinkela_wire_18832),
        .c(_0353_)
    );

    bfr new_Jinkela_buffer_5624 (
        .din(new_Jinkela_wire_7169),
        .dout(new_Jinkela_wire_7170)
    );

    bfr new_Jinkela_buffer_15973 (
        .din(new_Jinkela_wire_19029),
        .dout(new_Jinkela_wire_19030)
    );

    or_bb _3096_ (
        .a(new_Jinkela_wire_6734),
        .b(new_Jinkela_wire_5806),
        .c(_0354_)
    );

    bfr new_Jinkela_buffer_5584 (
        .din(new_Jinkela_wire_7121),
        .dout(new_Jinkela_wire_7122)
    );

    bfr new_Jinkela_buffer_16012 (
        .din(new_Jinkela_wire_19092),
        .dout(new_Jinkela_wire_19093)
    );

    and_ii _3097_ (
        .a(new_Jinkela_wire_18446),
        .b(new_Jinkela_wire_20574),
        .c(_0355_)
    );

    bfr new_Jinkela_buffer_5643 (
        .din(new_Jinkela_wire_7196),
        .dout(new_Jinkela_wire_7197)
    );

    bfr new_Jinkela_buffer_15974 (
        .din(new_Jinkela_wire_19030),
        .dout(new_Jinkela_wire_19031)
    );

    and_bb _3098_ (
        .a(new_Jinkela_wire_18447),
        .b(new_Jinkela_wire_20575),
        .c(_0356_)
    );

    bfr new_Jinkela_buffer_5585 (
        .din(new_Jinkela_wire_7122),
        .dout(new_Jinkela_wire_7123)
    );

    spl2 new_Jinkela_splitter_1397 (
        .a(new_Jinkela_wire_19123),
        .b(new_Jinkela_wire_19124),
        .c(new_Jinkela_wire_19125)
    );

    or_bb _3099_ (
        .a(new_Jinkela_wire_12621),
        .b(new_Jinkela_wire_12522),
        .c(_0357_)
    );

    bfr new_Jinkela_buffer_5625 (
        .din(new_Jinkela_wire_7170),
        .dout(new_Jinkela_wire_7171)
    );

    bfr new_Jinkela_buffer_15975 (
        .din(new_Jinkela_wire_19031),
        .dout(new_Jinkela_wire_19032)
    );

    and_ii _3100_ (
        .a(new_Jinkela_wire_21173),
        .b(new_Jinkela_wire_17357),
        .c(_0358_)
    );

    bfr new_Jinkela_buffer_5586 (
        .din(new_Jinkela_wire_7123),
        .dout(new_Jinkela_wire_7124)
    );

    bfr new_Jinkela_buffer_16013 (
        .din(new_Jinkela_wire_19093),
        .dout(new_Jinkela_wire_19094)
    );

    and_bb _3101_ (
        .a(new_Jinkela_wire_21174),
        .b(new_Jinkela_wire_17358),
        .c(_0359_)
    );

    bfr new_Jinkela_buffer_5710 (
        .din(new_Jinkela_wire_7267),
        .dout(new_Jinkela_wire_7268)
    );

    bfr new_Jinkela_buffer_15976 (
        .din(new_Jinkela_wire_19032),
        .dout(new_Jinkela_wire_19033)
    );

    or_bb _3102_ (
        .a(new_Jinkela_wire_14428),
        .b(new_Jinkela_wire_5136),
        .c(_0360_)
    );

    bfr new_Jinkela_buffer_5587 (
        .din(new_Jinkela_wire_7124),
        .dout(new_Jinkela_wire_7125)
    );

    bfr new_Jinkela_buffer_16027 (
        .din(new_Jinkela_wire_19129),
        .dout(new_Jinkela_wire_19130)
    );

    spl2 new_Jinkela_splitter_1401 (
        .a(_1338_),
        .b(new_Jinkela_wire_19144),
        .c(new_Jinkela_wire_19145)
    );

    and_ii _3103_ (
        .a(new_Jinkela_wire_2601),
        .b(new_Jinkela_wire_19391),
        .c(_0362_)
    );

    bfr new_Jinkela_buffer_5626 (
        .din(new_Jinkela_wire_7171),
        .dout(new_Jinkela_wire_7172)
    );

    bfr new_Jinkela_buffer_15977 (
        .din(new_Jinkela_wire_19033),
        .dout(new_Jinkela_wire_19034)
    );

    and_bb _3104_ (
        .a(new_Jinkela_wire_2602),
        .b(new_Jinkela_wire_19392),
        .c(_0363_)
    );

    spl2 new_Jinkela_splitter_618 (
        .a(new_Jinkela_wire_7125),
        .b(new_Jinkela_wire_7126),
        .c(new_Jinkela_wire_7127)
    );

    bfr new_Jinkela_buffer_16014 (
        .din(new_Jinkela_wire_19094),
        .dout(new_Jinkela_wire_19095)
    );

    or_bb _3105_ (
        .a(new_Jinkela_wire_4670),
        .b(new_Jinkela_wire_3709),
        .c(_0364_)
    );

    bfr new_Jinkela_buffer_5627 (
        .din(new_Jinkela_wire_7172),
        .dout(new_Jinkela_wire_7173)
    );

    bfr new_Jinkela_buffer_15978 (
        .din(new_Jinkela_wire_19034),
        .dout(new_Jinkela_wire_19035)
    );

    and_ii _3106_ (
        .a(new_Jinkela_wire_7314),
        .b(new_Jinkela_wire_11412),
        .c(_0365_)
    );

    bfr new_Jinkela_buffer_5644 (
        .din(new_Jinkela_wire_7197),
        .dout(new_Jinkela_wire_7198)
    );

    spl2 new_Jinkela_splitter_1400 (
        .a(_0319_),
        .b(new_Jinkela_wire_19134),
        .c(new_Jinkela_wire_19135)
    );

    and_bb _3107_ (
        .a(new_Jinkela_wire_7315),
        .b(new_Jinkela_wire_11413),
        .c(_0366_)
    );

    bfr new_Jinkela_buffer_15979 (
        .din(new_Jinkela_wire_19035),
        .dout(new_Jinkela_wire_19036)
    );

    or_bb _3108_ (
        .a(new_Jinkela_wire_17670),
        .b(new_Jinkela_wire_1596),
        .c(_0367_)
    );

    spl2 new_Jinkela_splitter_622 (
        .a(new_Jinkela_wire_7173),
        .b(new_Jinkela_wire_7174),
        .c(new_Jinkela_wire_7175)
    );

    bfr new_Jinkela_buffer_16015 (
        .din(new_Jinkela_wire_19095),
        .dout(new_Jinkela_wire_19096)
    );

    and_ii _3109_ (
        .a(new_Jinkela_wire_5284),
        .b(new_Jinkela_wire_18275),
        .c(_0368_)
    );

    bfr new_Jinkela_buffer_15980 (
        .din(new_Jinkela_wire_19036),
        .dout(new_Jinkela_wire_19037)
    );

    spl2 new_Jinkela_splitter_631 (
        .a(_1054_),
        .b(new_Jinkela_wire_7281),
        .c(new_Jinkela_wire_7282)
    );

    and_bb _3110_ (
        .a(new_Jinkela_wire_5285),
        .b(new_Jinkela_wire_18276),
        .c(_0369_)
    );

    bfr new_Jinkela_buffer_5645 (
        .din(new_Jinkela_wire_7198),
        .dout(new_Jinkela_wire_7199)
    );

    or_bb _3111_ (
        .a(new_Jinkela_wire_18699),
        .b(new_Jinkela_wire_14685),
        .c(_0370_)
    );

    bfr new_Jinkela_buffer_5646 (
        .din(new_Jinkela_wire_7199),
        .dout(new_Jinkela_wire_7200)
    );

    bfr new_Jinkela_buffer_15981 (
        .din(new_Jinkela_wire_19037),
        .dout(new_Jinkela_wire_19038)
    );

    and_ii _3112_ (
        .a(new_Jinkela_wire_5882),
        .b(new_Jinkela_wire_13572),
        .c(_0371_)
    );

    bfr new_Jinkela_buffer_5713 (
        .din(new_Jinkela_wire_7276),
        .dout(new_Jinkela_wire_7277)
    );

    bfr new_Jinkela_buffer_16016 (
        .din(new_Jinkela_wire_19096),
        .dout(new_Jinkela_wire_19097)
    );

    bfr new_Jinkela_buffer_5721 (
        .din(_0522_),
        .dout(new_Jinkela_wire_7287)
    );

    and_bb _3113_ (
        .a(new_Jinkela_wire_5883),
        .b(new_Jinkela_wire_13573),
        .c(_0373_)
    );

    bfr new_Jinkela_buffer_5647 (
        .din(new_Jinkela_wire_7200),
        .dout(new_Jinkela_wire_7201)
    );

    bfr new_Jinkela_buffer_15982 (
        .din(new_Jinkela_wire_19038),
        .dout(new_Jinkela_wire_19039)
    );

    or_bb _3114_ (
        .a(new_Jinkela_wire_1017),
        .b(new_Jinkela_wire_19964),
        .c(_0374_)
    );

    bfr new_Jinkela_buffer_16028 (
        .din(new_Jinkela_wire_19130),
        .dout(new_Jinkela_wire_19131)
    );

    and_ii _3115_ (
        .a(new_Jinkela_wire_10969),
        .b(new_Jinkela_wire_9805),
        .c(_0375_)
    );

    bfr new_Jinkela_buffer_5648 (
        .din(new_Jinkela_wire_7201),
        .dout(new_Jinkela_wire_7202)
    );

    bfr new_Jinkela_buffer_15983 (
        .din(new_Jinkela_wire_19039),
        .dout(new_Jinkela_wire_19040)
    );

    and_bb _3116_ (
        .a(new_Jinkela_wire_10970),
        .b(new_Jinkela_wire_9806),
        .c(_0376_)
    );

    bfr new_Jinkela_buffer_5714 (
        .din(new_Jinkela_wire_7277),
        .dout(new_Jinkela_wire_7278)
    );

    bfr new_Jinkela_buffer_16017 (
        .din(new_Jinkela_wire_19097),
        .dout(new_Jinkela_wire_19098)
    );

    or_bb _3117_ (
        .a(new_Jinkela_wire_20135),
        .b(new_Jinkela_wire_2711),
        .c(_0377_)
    );

    bfr new_Jinkela_buffer_5649 (
        .din(new_Jinkela_wire_7202),
        .dout(new_Jinkela_wire_7203)
    );

    bfr new_Jinkela_buffer_15984 (
        .din(new_Jinkela_wire_19040),
        .dout(new_Jinkela_wire_19041)
    );

    and_ii _3118_ (
        .a(new_Jinkela_wire_16904),
        .b(new_Jinkela_wire_12052),
        .c(_0378_)
    );

    bfr new_Jinkela_buffer_5717 (
        .din(new_Jinkela_wire_7282),
        .dout(new_Jinkela_wire_7283)
    );

    bfr new_Jinkela_buffer_16031 (
        .din(new_Jinkela_wire_19135),
        .dout(new_Jinkela_wire_19136)
    );

    bfr new_Jinkela_buffer_5722 (
        .din(_0131_),
        .dout(new_Jinkela_wire_7288)
    );

    spl2 new_Jinkela_splitter_1402 (
        .a(_1758_),
        .b(new_Jinkela_wire_19150),
        .c(new_Jinkela_wire_19151)
    );

    and_bb _3119_ (
        .a(new_Jinkela_wire_16905),
        .b(new_Jinkela_wire_12053),
        .c(_0379_)
    );

    bfr new_Jinkela_buffer_5650 (
        .din(new_Jinkela_wire_7203),
        .dout(new_Jinkela_wire_7204)
    );

    bfr new_Jinkela_buffer_15985 (
        .din(new_Jinkela_wire_19041),
        .dout(new_Jinkela_wire_19042)
    );

    or_bb _3120_ (
        .a(new_Jinkela_wire_13198),
        .b(new_Jinkela_wire_2129),
        .c(_0380_)
    );

    bfr new_Jinkela_buffer_5715 (
        .din(new_Jinkela_wire_7278),
        .dout(new_Jinkela_wire_7279)
    );

    bfr new_Jinkela_buffer_16018 (
        .din(new_Jinkela_wire_19098),
        .dout(new_Jinkela_wire_19099)
    );

    and_ii _3121_ (
        .a(new_Jinkela_wire_10395),
        .b(new_Jinkela_wire_3549),
        .c(_0381_)
    );

    bfr new_Jinkela_buffer_5651 (
        .din(new_Jinkela_wire_7204),
        .dout(new_Jinkela_wire_7205)
    );

    spl2 new_Jinkela_splitter_1377 (
        .a(new_Jinkela_wire_19042),
        .b(new_Jinkela_wire_19043),
        .c(new_Jinkela_wire_19044)
    );

    and_bb _3122_ (
        .a(new_Jinkela_wire_10396),
        .b(new_Jinkela_wire_3550),
        .c(_0382_)
    );

    bfr new_Jinkela_buffer_16019 (
        .din(new_Jinkela_wire_19099),
        .dout(new_Jinkela_wire_19100)
    );

    spl2 new_Jinkela_splitter_632 (
        .a(_1257_),
        .b(new_Jinkela_wire_7289),
        .c(new_Jinkela_wire_7290)
    );

    or_bb _3123_ (
        .a(new_Jinkela_wire_18687),
        .b(new_Jinkela_wire_2595),
        .c(_0384_)
    );

    bfr new_Jinkela_buffer_5652 (
        .din(new_Jinkela_wire_7205),
        .dout(new_Jinkela_wire_7206)
    );

    bfr new_Jinkela_buffer_16029 (
        .din(new_Jinkela_wire_19131),
        .dout(new_Jinkela_wire_19132)
    );

    and_ii _3124_ (
        .a(new_Jinkela_wire_17026),
        .b(new_Jinkela_wire_3817),
        .c(_0385_)
    );

    bfr new_Jinkela_buffer_5716 (
        .din(new_Jinkela_wire_7279),
        .dout(new_Jinkela_wire_7280)
    );

    bfr new_Jinkela_buffer_16039 (
        .din(new_Jinkela_wire_19145),
        .dout(new_Jinkela_wire_19146)
    );

    and_bb _3125_ (
        .a(new_Jinkela_wire_17027),
        .b(new_Jinkela_wire_3818),
        .c(_0386_)
    );

    bfr new_Jinkela_buffer_5653 (
        .din(new_Jinkela_wire_7206),
        .dout(new_Jinkela_wire_7207)
    );

    bfr new_Jinkela_buffer_16020 (
        .din(new_Jinkela_wire_19100),
        .dout(new_Jinkela_wire_19101)
    );

    or_bb _3126_ (
        .a(new_Jinkela_wire_19054),
        .b(new_Jinkela_wire_14311),
        .c(_0387_)
    );

    bfr new_Jinkela_buffer_5718 (
        .din(new_Jinkela_wire_7283),
        .dout(new_Jinkela_wire_7284)
    );

    bfr new_Jinkela_buffer_16030 (
        .din(new_Jinkela_wire_19132),
        .dout(new_Jinkela_wire_19133)
    );

    and_ii _3127_ (
        .a(new_Jinkela_wire_6804),
        .b(new_Jinkela_wire_2417),
        .c(_0388_)
    );

    bfr new_Jinkela_buffer_5654 (
        .din(new_Jinkela_wire_7207),
        .dout(new_Jinkela_wire_7208)
    );

    bfr new_Jinkela_buffer_16021 (
        .din(new_Jinkela_wire_19101),
        .dout(new_Jinkela_wire_19102)
    );

    and_bb _3128_ (
        .a(new_Jinkela_wire_6805),
        .b(new_Jinkela_wire_2418),
        .c(_0389_)
    );

    bfr new_Jinkela_buffer_5723 (
        .din(_0730_),
        .dout(new_Jinkela_wire_7291)
    );

    bfr new_Jinkela_buffer_16032 (
        .din(new_Jinkela_wire_19136),
        .dout(new_Jinkela_wire_19137)
    );

    or_bb _3129_ (
        .a(new_Jinkela_wire_15666),
        .b(new_Jinkela_wire_2787),
        .c(_0390_)
    );

    bfr new_Jinkela_buffer_5655 (
        .din(new_Jinkela_wire_7208),
        .dout(new_Jinkela_wire_7209)
    );

    bfr new_Jinkela_buffer_16022 (
        .din(new_Jinkela_wire_19102),
        .dout(new_Jinkela_wire_19103)
    );

    spl2 new_Jinkela_splitter_865 (
        .a(_1039_),
        .b(new_Jinkela_wire_11386),
        .c(new_Jinkela_wire_11387)
    );

    bfr new_Jinkela_buffer_9067 (
        .din(new_Jinkela_wire_11082),
        .dout(new_Jinkela_wire_11083)
    );

    bfr new_Jinkela_buffer_9135 (
        .din(new_Jinkela_wire_11154),
        .dout(new_Jinkela_wire_11155)
    );

    bfr new_Jinkela_buffer_9068 (
        .din(new_Jinkela_wire_11083),
        .dout(new_Jinkela_wire_11084)
    );

    bfr new_Jinkela_buffer_9216 (
        .din(new_Jinkela_wire_11239),
        .dout(new_Jinkela_wire_11240)
    );

    bfr new_Jinkela_buffer_9069 (
        .din(new_Jinkela_wire_11084),
        .dout(new_Jinkela_wire_11085)
    );

    bfr new_Jinkela_buffer_9136 (
        .din(new_Jinkela_wire_11155),
        .dout(new_Jinkela_wire_11156)
    );

    bfr new_Jinkela_buffer_9070 (
        .din(new_Jinkela_wire_11085),
        .dout(new_Jinkela_wire_11086)
    );

    spl2 new_Jinkela_splitter_866 (
        .a(_1093_),
        .b(new_Jinkela_wire_11388),
        .c(new_Jinkela_wire_11389)
    );

    bfr new_Jinkela_buffer_9071 (
        .din(new_Jinkela_wire_11086),
        .dout(new_Jinkela_wire_11087)
    );

    bfr new_Jinkela_buffer_9137 (
        .din(new_Jinkela_wire_11156),
        .dout(new_Jinkela_wire_11157)
    );

    bfr new_Jinkela_buffer_9072 (
        .din(new_Jinkela_wire_11087),
        .dout(new_Jinkela_wire_11088)
    );

    bfr new_Jinkela_buffer_9217 (
        .din(new_Jinkela_wire_11240),
        .dout(new_Jinkela_wire_11241)
    );

    bfr new_Jinkela_buffer_9073 (
        .din(new_Jinkela_wire_11088),
        .dout(new_Jinkela_wire_11089)
    );

    bfr new_Jinkela_buffer_9138 (
        .din(new_Jinkela_wire_11157),
        .dout(new_Jinkela_wire_11158)
    );

    bfr new_Jinkela_buffer_9074 (
        .din(new_Jinkela_wire_11089),
        .dout(new_Jinkela_wire_11090)
    );

    bfr new_Jinkela_buffer_9317 (
        .din(new_Jinkela_wire_11346),
        .dout(new_Jinkela_wire_11347)
    );

    bfr new_Jinkela_buffer_9075 (
        .din(new_Jinkela_wire_11090),
        .dout(new_Jinkela_wire_11091)
    );

    bfr new_Jinkela_buffer_9139 (
        .din(new_Jinkela_wire_11158),
        .dout(new_Jinkela_wire_11159)
    );

    bfr new_Jinkela_buffer_9076 (
        .din(new_Jinkela_wire_11091),
        .dout(new_Jinkela_wire_11092)
    );

    bfr new_Jinkela_buffer_9218 (
        .din(new_Jinkela_wire_11241),
        .dout(new_Jinkela_wire_11242)
    );

    bfr new_Jinkela_buffer_9077 (
        .din(new_Jinkela_wire_11092),
        .dout(new_Jinkela_wire_11093)
    );

    bfr new_Jinkela_buffer_9140 (
        .din(new_Jinkela_wire_11159),
        .dout(new_Jinkela_wire_11160)
    );

    bfr new_Jinkela_buffer_9078 (
        .din(new_Jinkela_wire_11093),
        .dout(new_Jinkela_wire_11094)
    );

    bfr new_Jinkela_buffer_9321 (
        .din(new_Jinkela_wire_11350),
        .dout(new_Jinkela_wire_11351)
    );

    bfr new_Jinkela_buffer_9079 (
        .din(new_Jinkela_wire_11094),
        .dout(new_Jinkela_wire_11095)
    );

    bfr new_Jinkela_buffer_9141 (
        .din(new_Jinkela_wire_11160),
        .dout(new_Jinkela_wire_11161)
    );

    bfr new_Jinkela_buffer_9080 (
        .din(new_Jinkela_wire_11095),
        .dout(new_Jinkela_wire_11096)
    );

    bfr new_Jinkela_buffer_9219 (
        .din(new_Jinkela_wire_11242),
        .dout(new_Jinkela_wire_11243)
    );

    bfr new_Jinkela_buffer_9081 (
        .din(new_Jinkela_wire_11096),
        .dout(new_Jinkela_wire_11097)
    );

    bfr new_Jinkela_buffer_9142 (
        .din(new_Jinkela_wire_11161),
        .dout(new_Jinkela_wire_11162)
    );

    bfr new_Jinkela_buffer_9082 (
        .din(new_Jinkela_wire_11097),
        .dout(new_Jinkela_wire_11098)
    );

    bfr new_Jinkela_buffer_9318 (
        .din(new_Jinkela_wire_11347),
        .dout(new_Jinkela_wire_11348)
    );

    bfr new_Jinkela_buffer_9083 (
        .din(new_Jinkela_wire_11098),
        .dout(new_Jinkela_wire_11099)
    );

    bfr new_Jinkela_buffer_9143 (
        .din(new_Jinkela_wire_11162),
        .dout(new_Jinkela_wire_11163)
    );

    bfr new_Jinkela_buffer_9084 (
        .din(new_Jinkela_wire_11099),
        .dout(new_Jinkela_wire_11100)
    );

    bfr new_Jinkela_buffer_9220 (
        .din(new_Jinkela_wire_11243),
        .dout(new_Jinkela_wire_11244)
    );

    bfr new_Jinkela_buffer_9085 (
        .din(new_Jinkela_wire_11100),
        .dout(new_Jinkela_wire_11101)
    );

    bfr new_Jinkela_buffer_9144 (
        .din(new_Jinkela_wire_11163),
        .dout(new_Jinkela_wire_11164)
    );

    bfr new_Jinkela_buffer_9086 (
        .din(new_Jinkela_wire_11101),
        .dout(new_Jinkela_wire_11102)
    );

    bfr new_Jinkela_buffer_9354 (
        .din(_1238_),
        .dout(new_Jinkela_wire_11390)
    );

    bfr new_Jinkela_buffer_9087 (
        .din(new_Jinkela_wire_11102),
        .dout(new_Jinkela_wire_11103)
    );

    bfr new_Jinkela_buffer_12557 (
        .din(new_Jinkela_wire_15064),
        .dout(new_Jinkela_wire_15065)
    );

    bfr new_Jinkela_buffer_12626 (
        .din(new_Jinkela_wire_15141),
        .dout(new_Jinkela_wire_15142)
    );

    bfr new_Jinkela_buffer_12558 (
        .din(new_Jinkela_wire_15065),
        .dout(new_Jinkela_wire_15066)
    );

    bfr new_Jinkela_buffer_12874 (
        .din(new_Jinkela_wire_15395),
        .dout(new_Jinkela_wire_15396)
    );

    bfr new_Jinkela_buffer_12691 (
        .din(new_Jinkela_wire_15212),
        .dout(new_Jinkela_wire_15213)
    );

    bfr new_Jinkela_buffer_12559 (
        .din(new_Jinkela_wire_15066),
        .dout(new_Jinkela_wire_15067)
    );

    bfr new_Jinkela_buffer_12627 (
        .din(new_Jinkela_wire_15142),
        .dout(new_Jinkela_wire_15143)
    );

    bfr new_Jinkela_buffer_12560 (
        .din(new_Jinkela_wire_15067),
        .dout(new_Jinkela_wire_15068)
    );

    bfr new_Jinkela_buffer_12860 (
        .din(new_Jinkela_wire_15381),
        .dout(new_Jinkela_wire_15382)
    );

    bfr new_Jinkela_buffer_12561 (
        .din(new_Jinkela_wire_15068),
        .dout(new_Jinkela_wire_15069)
    );

    bfr new_Jinkela_buffer_12628 (
        .din(new_Jinkela_wire_15143),
        .dout(new_Jinkela_wire_15144)
    );

    bfr new_Jinkela_buffer_12562 (
        .din(new_Jinkela_wire_15069),
        .dout(new_Jinkela_wire_15070)
    );

    bfr new_Jinkela_buffer_12692 (
        .din(new_Jinkela_wire_15213),
        .dout(new_Jinkela_wire_15214)
    );

    bfr new_Jinkela_buffer_12563 (
        .din(new_Jinkela_wire_15070),
        .dout(new_Jinkela_wire_15071)
    );

    bfr new_Jinkela_buffer_12629 (
        .din(new_Jinkela_wire_15144),
        .dout(new_Jinkela_wire_15145)
    );

    bfr new_Jinkela_buffer_12564 (
        .din(new_Jinkela_wire_15071),
        .dout(new_Jinkela_wire_15072)
    );

    bfr new_Jinkela_buffer_12565 (
        .din(new_Jinkela_wire_15072),
        .dout(new_Jinkela_wire_15073)
    );

    bfr new_Jinkela_buffer_12630 (
        .din(new_Jinkela_wire_15145),
        .dout(new_Jinkela_wire_15146)
    );

    bfr new_Jinkela_buffer_12566 (
        .din(new_Jinkela_wire_15073),
        .dout(new_Jinkela_wire_15074)
    );

    bfr new_Jinkela_buffer_12693 (
        .din(new_Jinkela_wire_15214),
        .dout(new_Jinkela_wire_15215)
    );

    bfr new_Jinkela_buffer_12567 (
        .din(new_Jinkela_wire_15074),
        .dout(new_Jinkela_wire_15075)
    );

    bfr new_Jinkela_buffer_12631 (
        .din(new_Jinkela_wire_15146),
        .dout(new_Jinkela_wire_15147)
    );

    bfr new_Jinkela_buffer_12568 (
        .din(new_Jinkela_wire_15075),
        .dout(new_Jinkela_wire_15076)
    );

    bfr new_Jinkela_buffer_12861 (
        .din(new_Jinkela_wire_15382),
        .dout(new_Jinkela_wire_15383)
    );

    bfr new_Jinkela_buffer_12569 (
        .din(new_Jinkela_wire_15076),
        .dout(new_Jinkela_wire_15077)
    );

    bfr new_Jinkela_buffer_12632 (
        .din(new_Jinkela_wire_15147),
        .dout(new_Jinkela_wire_15148)
    );

    bfr new_Jinkela_buffer_12570 (
        .din(new_Jinkela_wire_15077),
        .dout(new_Jinkela_wire_15078)
    );

    bfr new_Jinkela_buffer_12694 (
        .din(new_Jinkela_wire_15215),
        .dout(new_Jinkela_wire_15216)
    );

    bfr new_Jinkela_buffer_12571 (
        .din(new_Jinkela_wire_15078),
        .dout(new_Jinkela_wire_15079)
    );

    bfr new_Jinkela_buffer_12633 (
        .din(new_Jinkela_wire_15148),
        .dout(new_Jinkela_wire_15149)
    );

    bfr new_Jinkela_buffer_12572 (
        .din(new_Jinkela_wire_15079),
        .dout(new_Jinkela_wire_15080)
    );

    bfr new_Jinkela_buffer_12946 (
        .din(new_Jinkela_wire_15469),
        .dout(new_Jinkela_wire_15470)
    );

    bfr new_Jinkela_buffer_12573 (
        .din(new_Jinkela_wire_15080),
        .dout(new_Jinkela_wire_15081)
    );

    bfr new_Jinkela_buffer_12634 (
        .din(new_Jinkela_wire_15149),
        .dout(new_Jinkela_wire_15150)
    );

    bfr new_Jinkela_buffer_12574 (
        .din(new_Jinkela_wire_15081),
        .dout(new_Jinkela_wire_15082)
    );

    bfr new_Jinkela_buffer_12875 (
        .din(new_Jinkela_wire_15396),
        .dout(new_Jinkela_wire_15397)
    );

    bfr new_Jinkela_buffer_12695 (
        .din(new_Jinkela_wire_15216),
        .dout(new_Jinkela_wire_15217)
    );

    bfr new_Jinkela_buffer_12575 (
        .din(new_Jinkela_wire_15082),
        .dout(new_Jinkela_wire_15083)
    );

    bfr new_Jinkela_buffer_12635 (
        .din(new_Jinkela_wire_15150),
        .dout(new_Jinkela_wire_15151)
    );

    bfr new_Jinkela_buffer_12576 (
        .din(new_Jinkela_wire_15083),
        .dout(new_Jinkela_wire_15084)
    );

    bfr new_Jinkela_buffer_12862 (
        .din(new_Jinkela_wire_15383),
        .dout(new_Jinkela_wire_15384)
    );

    bfr new_Jinkela_buffer_12577 (
        .din(new_Jinkela_wire_15084),
        .dout(new_Jinkela_wire_15085)
    );

    bfr new_Jinkela_buffer_12636 (
        .din(new_Jinkela_wire_15151),
        .dout(new_Jinkela_wire_15152)
    );

    bfr new_Jinkela_buffer_9145 (
        .din(new_Jinkela_wire_11164),
        .dout(new_Jinkela_wire_11165)
    );

    bfr new_Jinkela_buffer_9088 (
        .din(new_Jinkela_wire_11103),
        .dout(new_Jinkela_wire_11104)
    );

    bfr new_Jinkela_buffer_9221 (
        .din(new_Jinkela_wire_11244),
        .dout(new_Jinkela_wire_11245)
    );

    bfr new_Jinkela_buffer_9089 (
        .din(new_Jinkela_wire_11104),
        .dout(new_Jinkela_wire_11105)
    );

    bfr new_Jinkela_buffer_9146 (
        .din(new_Jinkela_wire_11165),
        .dout(new_Jinkela_wire_11166)
    );

    bfr new_Jinkela_buffer_9090 (
        .din(new_Jinkela_wire_11105),
        .dout(new_Jinkela_wire_11106)
    );

    bfr new_Jinkela_buffer_9319 (
        .din(new_Jinkela_wire_11348),
        .dout(new_Jinkela_wire_11349)
    );

    bfr new_Jinkela_buffer_9091 (
        .din(new_Jinkela_wire_11106),
        .dout(new_Jinkela_wire_11107)
    );

    bfr new_Jinkela_buffer_9147 (
        .din(new_Jinkela_wire_11166),
        .dout(new_Jinkela_wire_11167)
    );

    bfr new_Jinkela_buffer_9092 (
        .din(new_Jinkela_wire_11107),
        .dout(new_Jinkela_wire_11108)
    );

    bfr new_Jinkela_buffer_9222 (
        .din(new_Jinkela_wire_11245),
        .dout(new_Jinkela_wire_11246)
    );

    bfr new_Jinkela_buffer_9093 (
        .din(new_Jinkela_wire_11108),
        .dout(new_Jinkela_wire_11109)
    );

    bfr new_Jinkela_buffer_9148 (
        .din(new_Jinkela_wire_11167),
        .dout(new_Jinkela_wire_11168)
    );

    bfr new_Jinkela_buffer_9094 (
        .din(new_Jinkela_wire_11109),
        .dout(new_Jinkela_wire_11110)
    );

    bfr new_Jinkela_buffer_9322 (
        .din(new_Jinkela_wire_11351),
        .dout(new_Jinkela_wire_11352)
    );

    bfr new_Jinkela_buffer_9095 (
        .din(new_Jinkela_wire_11110),
        .dout(new_Jinkela_wire_11111)
    );

    bfr new_Jinkela_buffer_9149 (
        .din(new_Jinkela_wire_11168),
        .dout(new_Jinkela_wire_11169)
    );

    bfr new_Jinkela_buffer_9096 (
        .din(new_Jinkela_wire_11111),
        .dout(new_Jinkela_wire_11112)
    );

    bfr new_Jinkela_buffer_9223 (
        .din(new_Jinkela_wire_11246),
        .dout(new_Jinkela_wire_11247)
    );

    bfr new_Jinkela_buffer_9097 (
        .din(new_Jinkela_wire_11112),
        .dout(new_Jinkela_wire_11113)
    );

    bfr new_Jinkela_buffer_9150 (
        .din(new_Jinkela_wire_11169),
        .dout(new_Jinkela_wire_11170)
    );

    bfr new_Jinkela_buffer_9098 (
        .din(new_Jinkela_wire_11113),
        .dout(new_Jinkela_wire_11114)
    );

    spl2 new_Jinkela_splitter_868 (
        .a(_0565_),
        .b(new_Jinkela_wire_11393),
        .c(new_Jinkela_wire_11394)
    );

    bfr new_Jinkela_buffer_9099 (
        .din(new_Jinkela_wire_11114),
        .dout(new_Jinkela_wire_11115)
    );

    bfr new_Jinkela_buffer_9151 (
        .din(new_Jinkela_wire_11170),
        .dout(new_Jinkela_wire_11171)
    );

    bfr new_Jinkela_buffer_9100 (
        .din(new_Jinkela_wire_11115),
        .dout(new_Jinkela_wire_11116)
    );

    bfr new_Jinkela_buffer_9224 (
        .din(new_Jinkela_wire_11247),
        .dout(new_Jinkela_wire_11248)
    );

    bfr new_Jinkela_buffer_9101 (
        .din(new_Jinkela_wire_11116),
        .dout(new_Jinkela_wire_11117)
    );

    bfr new_Jinkela_buffer_9152 (
        .din(new_Jinkela_wire_11171),
        .dout(new_Jinkela_wire_11172)
    );

    bfr new_Jinkela_buffer_9102 (
        .din(new_Jinkela_wire_11117),
        .dout(new_Jinkela_wire_11118)
    );

    bfr new_Jinkela_buffer_9323 (
        .din(new_Jinkela_wire_11352),
        .dout(new_Jinkela_wire_11353)
    );

    bfr new_Jinkela_buffer_9103 (
        .din(new_Jinkela_wire_11118),
        .dout(new_Jinkela_wire_11119)
    );

    bfr new_Jinkela_buffer_9153 (
        .din(new_Jinkela_wire_11172),
        .dout(new_Jinkela_wire_11173)
    );

    bfr new_Jinkela_buffer_9104 (
        .din(new_Jinkela_wire_11119),
        .dout(new_Jinkela_wire_11120)
    );

    bfr new_Jinkela_buffer_9225 (
        .din(new_Jinkela_wire_11248),
        .dout(new_Jinkela_wire_11249)
    );

    bfr new_Jinkela_buffer_9105 (
        .din(new_Jinkela_wire_11120),
        .dout(new_Jinkela_wire_11121)
    );

    bfr new_Jinkela_buffer_9154 (
        .din(new_Jinkela_wire_11173),
        .dout(new_Jinkela_wire_11174)
    );

    bfr new_Jinkela_buffer_9106 (
        .din(new_Jinkela_wire_11121),
        .dout(new_Jinkela_wire_11122)
    );

    spl2 new_Jinkela_splitter_867 (
        .a(_0457_),
        .b(new_Jinkela_wire_11391),
        .c(new_Jinkela_wire_11392)
    );

    bfr new_Jinkela_buffer_9107 (
        .din(new_Jinkela_wire_11122),
        .dout(new_Jinkela_wire_11123)
    );

    bfr new_Jinkela_buffer_9155 (
        .din(new_Jinkela_wire_11174),
        .dout(new_Jinkela_wire_11175)
    );

    bfr new_Jinkela_buffer_9108 (
        .din(new_Jinkela_wire_11123),
        .dout(new_Jinkela_wire_11124)
    );

    bfr new_Jinkela_buffer_5719 (
        .din(new_Jinkela_wire_7284),
        .dout(new_Jinkela_wire_7285)
    );

    bfr new_Jinkela_buffer_9226 (
        .din(new_Jinkela_wire_11249),
        .dout(new_Jinkela_wire_11250)
    );

    bfr new_Jinkela_buffer_12578 (
        .din(new_Jinkela_wire_15085),
        .dout(new_Jinkela_wire_15086)
    );

    spl2 new_Jinkela_splitter_1403 (
        .a(_1486_),
        .b(new_Jinkela_wire_19156),
        .c(new_Jinkela_wire_19157)
    );

    bfr new_Jinkela_buffer_5656 (
        .din(new_Jinkela_wire_7209),
        .dout(new_Jinkela_wire_7210)
    );

    bfr new_Jinkela_buffer_9109 (
        .din(new_Jinkela_wire_11124),
        .dout(new_Jinkela_wire_11125)
    );

    bfr new_Jinkela_buffer_16023 (
        .din(new_Jinkela_wire_19103),
        .dout(new_Jinkela_wire_19104)
    );

    bfr new_Jinkela_buffer_12696 (
        .din(new_Jinkela_wire_15217),
        .dout(new_Jinkela_wire_15218)
    );

    spl2 new_Jinkela_splitter_634 (
        .a(_0557_),
        .b(new_Jinkela_wire_7294),
        .c(new_Jinkela_wire_7295)
    );

    bfr new_Jinkela_buffer_9156 (
        .din(new_Jinkela_wire_11175),
        .dout(new_Jinkela_wire_11176)
    );

    bfr new_Jinkela_buffer_12579 (
        .din(new_Jinkela_wire_15086),
        .dout(new_Jinkela_wire_15087)
    );

    bfr new_Jinkela_buffer_16033 (
        .din(new_Jinkela_wire_19137),
        .dout(new_Jinkela_wire_19138)
    );

    bfr new_Jinkela_buffer_5657 (
        .din(new_Jinkela_wire_7210),
        .dout(new_Jinkela_wire_7211)
    );

    bfr new_Jinkela_buffer_9110 (
        .din(new_Jinkela_wire_11125),
        .dout(new_Jinkela_wire_11126)
    );

    bfr new_Jinkela_buffer_12637 (
        .din(new_Jinkela_wire_15152),
        .dout(new_Jinkela_wire_15153)
    );

    spl2 new_Jinkela_splitter_1389 (
        .a(new_Jinkela_wire_19104),
        .b(new_Jinkela_wire_19105),
        .c(new_Jinkela_wire_19106)
    );

    bfr new_Jinkela_buffer_5720 (
        .din(new_Jinkela_wire_7285),
        .dout(new_Jinkela_wire_7286)
    );

    bfr new_Jinkela_buffer_9324 (
        .din(new_Jinkela_wire_11353),
        .dout(new_Jinkela_wire_11354)
    );

    bfr new_Jinkela_buffer_12580 (
        .din(new_Jinkela_wire_15087),
        .dout(new_Jinkela_wire_15088)
    );

    bfr new_Jinkela_buffer_16034 (
        .din(new_Jinkela_wire_19138),
        .dout(new_Jinkela_wire_19139)
    );

    bfr new_Jinkela_buffer_5658 (
        .din(new_Jinkela_wire_7211),
        .dout(new_Jinkela_wire_7212)
    );

    bfr new_Jinkela_buffer_9111 (
        .din(new_Jinkela_wire_11126),
        .dout(new_Jinkela_wire_11127)
    );

    bfr new_Jinkela_buffer_9157 (
        .din(new_Jinkela_wire_11176),
        .dout(new_Jinkela_wire_11177)
    );

    bfr new_Jinkela_buffer_12581 (
        .din(new_Jinkela_wire_15088),
        .dout(new_Jinkela_wire_15089)
    );

    bfr new_Jinkela_buffer_16040 (
        .din(new_Jinkela_wire_19146),
        .dout(new_Jinkela_wire_19147)
    );

    spl2 new_Jinkela_splitter_633 (
        .a(_1234_),
        .b(new_Jinkela_wire_7292),
        .c(new_Jinkela_wire_7293)
    );

    bfr new_Jinkela_buffer_5659 (
        .din(new_Jinkela_wire_7212),
        .dout(new_Jinkela_wire_7213)
    );

    bfr new_Jinkela_buffer_9112 (
        .din(new_Jinkela_wire_11127),
        .dout(new_Jinkela_wire_11128)
    );

    bfr new_Jinkela_buffer_12638 (
        .din(new_Jinkela_wire_15153),
        .dout(new_Jinkela_wire_15154)
    );

    bfr new_Jinkela_buffer_16035 (
        .din(new_Jinkela_wire_19139),
        .dout(new_Jinkela_wire_19140)
    );

    bfr new_Jinkela_buffer_9227 (
        .din(new_Jinkela_wire_11250),
        .dout(new_Jinkela_wire_11251)
    );

    bfr new_Jinkela_buffer_12582 (
        .din(new_Jinkela_wire_15089),
        .dout(new_Jinkela_wire_15090)
    );

    bfr new_Jinkela_buffer_16043 (
        .din(new_Jinkela_wire_19151),
        .dout(new_Jinkela_wire_19152)
    );

    bfr new_Jinkela_buffer_16047 (
        .din(_0974_),
        .dout(new_Jinkela_wire_19158)
    );

    bfr new_Jinkela_buffer_5660 (
        .din(new_Jinkela_wire_7213),
        .dout(new_Jinkela_wire_7214)
    );

    bfr new_Jinkela_buffer_9113 (
        .din(new_Jinkela_wire_11128),
        .dout(new_Jinkela_wire_11129)
    );

    bfr new_Jinkela_buffer_16036 (
        .din(new_Jinkela_wire_19140),
        .dout(new_Jinkela_wire_19141)
    );

    bfr new_Jinkela_buffer_12697 (
        .din(new_Jinkela_wire_15218),
        .dout(new_Jinkela_wire_15219)
    );

    bfr new_Jinkela_buffer_9158 (
        .din(new_Jinkela_wire_11177),
        .dout(new_Jinkela_wire_11178)
    );

    bfr new_Jinkela_buffer_12583 (
        .din(new_Jinkela_wire_15090),
        .dout(new_Jinkela_wire_15091)
    );

    bfr new_Jinkela_buffer_16041 (
        .din(new_Jinkela_wire_19147),
        .dout(new_Jinkela_wire_19148)
    );

    spl2 new_Jinkela_splitter_635 (
        .a(_0552_),
        .b(new_Jinkela_wire_7296),
        .c(new_Jinkela_wire_7297)
    );

    bfr new_Jinkela_buffer_5661 (
        .din(new_Jinkela_wire_7214),
        .dout(new_Jinkela_wire_7215)
    );

    bfr new_Jinkela_buffer_9114 (
        .din(new_Jinkela_wire_11129),
        .dout(new_Jinkela_wire_11130)
    );

    bfr new_Jinkela_buffer_12639 (
        .din(new_Jinkela_wire_15154),
        .dout(new_Jinkela_wire_15155)
    );

    bfr new_Jinkela_buffer_16037 (
        .din(new_Jinkela_wire_19141),
        .dout(new_Jinkela_wire_19142)
    );

    bfr new_Jinkela_buffer_12584 (
        .din(new_Jinkela_wire_15091),
        .dout(new_Jinkela_wire_15092)
    );

    spl2 new_Jinkela_splitter_636 (
        .a(_1276_),
        .b(new_Jinkela_wire_7298),
        .c(new_Jinkela_wire_7299)
    );

    bfr new_Jinkela_buffer_5662 (
        .din(new_Jinkela_wire_7215),
        .dout(new_Jinkela_wire_7216)
    );

    bfr new_Jinkela_buffer_9115 (
        .din(new_Jinkela_wire_11130),
        .dout(new_Jinkela_wire_11131)
    );

    bfr new_Jinkela_buffer_16038 (
        .din(new_Jinkela_wire_19142),
        .dout(new_Jinkela_wire_19143)
    );

    bfr new_Jinkela_buffer_12863 (
        .din(new_Jinkela_wire_15384),
        .dout(new_Jinkela_wire_15385)
    );

    bfr new_Jinkela_buffer_5725 (
        .din(new_Jinkela_wire_7302),
        .dout(new_Jinkela_wire_7303)
    );

    bfr new_Jinkela_buffer_9159 (
        .din(new_Jinkela_wire_11178),
        .dout(new_Jinkela_wire_11179)
    );

    bfr new_Jinkela_buffer_12585 (
        .din(new_Jinkela_wire_15092),
        .dout(new_Jinkela_wire_15093)
    );

    bfr new_Jinkela_buffer_5724 (
        .din(_1049_),
        .dout(new_Jinkela_wire_7300)
    );

    bfr new_Jinkela_buffer_16042 (
        .din(new_Jinkela_wire_19148),
        .dout(new_Jinkela_wire_19149)
    );

    bfr new_Jinkela_buffer_5663 (
        .din(new_Jinkela_wire_7216),
        .dout(new_Jinkela_wire_7217)
    );

    bfr new_Jinkela_buffer_9116 (
        .din(new_Jinkela_wire_11131),
        .dout(new_Jinkela_wire_11132)
    );

    bfr new_Jinkela_buffer_12640 (
        .din(new_Jinkela_wire_15155),
        .dout(new_Jinkela_wire_15156)
    );

    bfr new_Jinkela_buffer_16044 (
        .din(new_Jinkela_wire_19152),
        .dout(new_Jinkela_wire_19153)
    );

    spl2 new_Jinkela_splitter_638 (
        .a(_0082_),
        .b(new_Jinkela_wire_7307),
        .c(new_Jinkela_wire_7308)
    );

    bfr new_Jinkela_buffer_9228 (
        .din(new_Jinkela_wire_11251),
        .dout(new_Jinkela_wire_11252)
    );

    bfr new_Jinkela_buffer_12586 (
        .din(new_Jinkela_wire_15093),
        .dout(new_Jinkela_wire_15094)
    );

    spl2 new_Jinkela_splitter_637 (
        .a(_0752_),
        .b(new_Jinkela_wire_7301),
        .c(new_Jinkela_wire_7302)
    );

    spl2 new_Jinkela_splitter_1404 (
        .a(_1096_),
        .b(new_Jinkela_wire_19159),
        .c(new_Jinkela_wire_19160)
    );

    spl2 new_Jinkela_splitter_1405 (
        .a(_0109_),
        .b(new_Jinkela_wire_19161),
        .c(new_Jinkela_wire_19162)
    );

    bfr new_Jinkela_buffer_5664 (
        .din(new_Jinkela_wire_7217),
        .dout(new_Jinkela_wire_7218)
    );

    bfr new_Jinkela_buffer_9117 (
        .din(new_Jinkela_wire_11132),
        .dout(new_Jinkela_wire_11133)
    );

    bfr new_Jinkela_buffer_16045 (
        .din(new_Jinkela_wire_19153),
        .dout(new_Jinkela_wire_19154)
    );

    bfr new_Jinkela_buffer_12698 (
        .din(new_Jinkela_wire_15219),
        .dout(new_Jinkela_wire_15220)
    );

    bfr new_Jinkela_buffer_9160 (
        .din(new_Jinkela_wire_11179),
        .dout(new_Jinkela_wire_11180)
    );

    bfr new_Jinkela_buffer_12587 (
        .din(new_Jinkela_wire_15094),
        .dout(new_Jinkela_wire_15095)
    );

    bfr new_Jinkela_buffer_5665 (
        .din(new_Jinkela_wire_7218),
        .dout(new_Jinkela_wire_7219)
    );

    spl2 new_Jinkela_splitter_857 (
        .a(new_Jinkela_wire_11133),
        .b(new_Jinkela_wire_11134),
        .c(new_Jinkela_wire_11135)
    );

    bfr new_Jinkela_buffer_12641 (
        .din(new_Jinkela_wire_15156),
        .dout(new_Jinkela_wire_15157)
    );

    bfr new_Jinkela_buffer_16046 (
        .din(new_Jinkela_wire_19154),
        .dout(new_Jinkela_wire_19155)
    );

    bfr new_Jinkela_buffer_9161 (
        .din(new_Jinkela_wire_11180),
        .dout(new_Jinkela_wire_11181)
    );

    bfr new_Jinkela_buffer_12588 (
        .din(new_Jinkela_wire_15095),
        .dout(new_Jinkela_wire_15096)
    );

    spl2 new_Jinkela_splitter_639 (
        .a(_1709_),
        .b(new_Jinkela_wire_7309),
        .c(new_Jinkela_wire_7310)
    );

    bfr new_Jinkela_buffer_16048 (
        .din(_0579_),
        .dout(new_Jinkela_wire_19163)
    );

    bfr new_Jinkela_buffer_5666 (
        .din(new_Jinkela_wire_7219),
        .dout(new_Jinkela_wire_7220)
    );

    bfr new_Jinkela_buffer_9325 (
        .din(new_Jinkela_wire_11354),
        .dout(new_Jinkela_wire_11355)
    );

    spl2 new_Jinkela_splitter_1407 (
        .a(_0800_),
        .b(new_Jinkela_wire_19182),
        .c(new_Jinkela_wire_19183)
    );

    bfr new_Jinkela_buffer_16049 (
        .din(_0318_),
        .dout(new_Jinkela_wire_19164)
    );

    bfr new_Jinkela_buffer_9229 (
        .din(new_Jinkela_wire_11252),
        .dout(new_Jinkela_wire_11253)
    );

    bfr new_Jinkela_buffer_12589 (
        .din(new_Jinkela_wire_15096),
        .dout(new_Jinkela_wire_15097)
    );

    bfr new_Jinkela_buffer_16065 (
        .din(_0412_),
        .dout(new_Jinkela_wire_19184)
    );

    bfr new_Jinkela_buffer_5667 (
        .din(new_Jinkela_wire_7220),
        .dout(new_Jinkela_wire_7221)
    );

    bfr new_Jinkela_buffer_9162 (
        .din(new_Jinkela_wire_11181),
        .dout(new_Jinkela_wire_11182)
    );

    bfr new_Jinkela_buffer_12642 (
        .din(new_Jinkela_wire_15157),
        .dout(new_Jinkela_wire_15158)
    );

    bfr new_Jinkela_buffer_16050 (
        .din(new_Jinkela_wire_19164),
        .dout(new_Jinkela_wire_19165)
    );

    bfr new_Jinkela_buffer_5726 (
        .din(new_Jinkela_wire_7303),
        .dout(new_Jinkela_wire_7304)
    );

    bfr new_Jinkela_buffer_12590 (
        .din(new_Jinkela_wire_15097),
        .dout(new_Jinkela_wire_15098)
    );

    spl2 new_Jinkela_splitter_869 (
        .a(_1181_),
        .b(new_Jinkela_wire_11395),
        .c(new_Jinkela_wire_11396)
    );

    bfr new_Jinkela_buffer_5668 (
        .din(new_Jinkela_wire_7221),
        .dout(new_Jinkela_wire_7222)
    );

    bfr new_Jinkela_buffer_9163 (
        .din(new_Jinkela_wire_11182),
        .dout(new_Jinkela_wire_11183)
    );

    bfr new_Jinkela_buffer_12876 (
        .din(new_Jinkela_wire_15397),
        .dout(new_Jinkela_wire_15398)
    );

    bfr new_Jinkela_buffer_12699 (
        .din(new_Jinkela_wire_15220),
        .dout(new_Jinkela_wire_15221)
    );

    bfr new_Jinkela_buffer_16051 (
        .din(new_Jinkela_wire_19165),
        .dout(new_Jinkela_wire_19166)
    );

    bfr new_Jinkela_buffer_9230 (
        .din(new_Jinkela_wire_11253),
        .dout(new_Jinkela_wire_11254)
    );

    bfr new_Jinkela_buffer_12591 (
        .din(new_Jinkela_wire_15098),
        .dout(new_Jinkela_wire_15099)
    );

    spl2 new_Jinkela_splitter_1409 (
        .a(_0390_),
        .b(new_Jinkela_wire_19187),
        .c(new_Jinkela_wire_19188)
    );

    bfr new_Jinkela_buffer_5730 (
        .din(_0364_),
        .dout(new_Jinkela_wire_7312)
    );

    spl2 new_Jinkela_splitter_1408 (
        .a(_0851_),
        .b(new_Jinkela_wire_19185),
        .c(new_Jinkela_wire_19186)
    );

    bfr new_Jinkela_buffer_5669 (
        .din(new_Jinkela_wire_7222),
        .dout(new_Jinkela_wire_7223)
    );

    bfr new_Jinkela_buffer_9164 (
        .din(new_Jinkela_wire_11183),
        .dout(new_Jinkela_wire_11184)
    );

    bfr new_Jinkela_buffer_12643 (
        .din(new_Jinkela_wire_15158),
        .dout(new_Jinkela_wire_15159)
    );

    bfr new_Jinkela_buffer_16052 (
        .din(new_Jinkela_wire_19166),
        .dout(new_Jinkela_wire_19167)
    );

    bfr new_Jinkela_buffer_5727 (
        .din(new_Jinkela_wire_7304),
        .dout(new_Jinkela_wire_7305)
    );

    bfr new_Jinkela_buffer_9326 (
        .din(new_Jinkela_wire_11355),
        .dout(new_Jinkela_wire_11356)
    );

    bfr new_Jinkela_buffer_12592 (
        .din(new_Jinkela_wire_15099),
        .dout(new_Jinkela_wire_15100)
    );

    bfr new_Jinkela_buffer_5670 (
        .din(new_Jinkela_wire_7223),
        .dout(new_Jinkela_wire_7224)
    );

    bfr new_Jinkela_buffer_9165 (
        .din(new_Jinkela_wire_11184),
        .dout(new_Jinkela_wire_11185)
    );

    bfr new_Jinkela_buffer_16053 (
        .din(new_Jinkela_wire_19167),
        .dout(new_Jinkela_wire_19168)
    );

    bfr new_Jinkela_buffer_12864 (
        .din(new_Jinkela_wire_15385),
        .dout(new_Jinkela_wire_15386)
    );

    bfr new_Jinkela_buffer_5729 (
        .din(new_Jinkela_wire_7310),
        .dout(new_Jinkela_wire_7311)
    );

    bfr new_Jinkela_buffer_9231 (
        .din(new_Jinkela_wire_11254),
        .dout(new_Jinkela_wire_11255)
    );

    bfr new_Jinkela_buffer_12593 (
        .din(new_Jinkela_wire_15100),
        .dout(new_Jinkela_wire_15101)
    );

    spl2 new_Jinkela_splitter_641 (
        .a(_1311_),
        .b(new_Jinkela_wire_7316),
        .c(new_Jinkela_wire_7317)
    );

    bfr new_Jinkela_buffer_16066 (
        .din(_0805_),
        .dout(new_Jinkela_wire_19189)
    );

    bfr new_Jinkela_buffer_5671 (
        .din(new_Jinkela_wire_7224),
        .dout(new_Jinkela_wire_7225)
    );

    bfr new_Jinkela_buffer_9166 (
        .din(new_Jinkela_wire_11185),
        .dout(new_Jinkela_wire_11186)
    );

    bfr new_Jinkela_buffer_12644 (
        .din(new_Jinkela_wire_15159),
        .dout(new_Jinkela_wire_15160)
    );

    bfr new_Jinkela_buffer_16054 (
        .din(new_Jinkela_wire_19168),
        .dout(new_Jinkela_wire_19169)
    );

    bfr new_Jinkela_buffer_5728 (
        .din(new_Jinkela_wire_7305),
        .dout(new_Jinkela_wire_7306)
    );

    bfr new_Jinkela_buffer_12594 (
        .din(new_Jinkela_wire_15101),
        .dout(new_Jinkela_wire_15102)
    );

    bfr new_Jinkela_buffer_16067 (
        .din(_0335_),
        .dout(new_Jinkela_wire_19192)
    );

    spl2 new_Jinkela_splitter_870 (
        .a(_0877_),
        .b(new_Jinkela_wire_11397),
        .c(new_Jinkela_wire_11398)
    );

    spl2 new_Jinkela_splitter_1410 (
        .a(_0192_),
        .b(new_Jinkela_wire_19190),
        .c(new_Jinkela_wire_19191)
    );

    bfr new_Jinkela_buffer_5672 (
        .din(new_Jinkela_wire_7225),
        .dout(new_Jinkela_wire_7226)
    );

    bfr new_Jinkela_buffer_9167 (
        .din(new_Jinkela_wire_11186),
        .dout(new_Jinkela_wire_11187)
    );

    bfr new_Jinkela_buffer_16055 (
        .din(new_Jinkela_wire_19169),
        .dout(new_Jinkela_wire_19170)
    );

    bfr new_Jinkela_buffer_12700 (
        .din(new_Jinkela_wire_15221),
        .dout(new_Jinkela_wire_15222)
    );

    bfr new_Jinkela_buffer_9232 (
        .din(new_Jinkela_wire_11255),
        .dout(new_Jinkela_wire_11256)
    );

    bfr new_Jinkela_buffer_12595 (
        .din(new_Jinkela_wire_15102),
        .dout(new_Jinkela_wire_15103)
    );

    spl2 new_Jinkela_splitter_1413 (
        .a(_1738_),
        .b(new_Jinkela_wire_19276),
        .c(new_Jinkela_wire_19277)
    );

    spl2 new_Jinkela_splitter_642 (
        .a(_1495_),
        .b(new_Jinkela_wire_7318),
        .c(new_Jinkela_wire_7319)
    );

    bfr new_Jinkela_buffer_5673 (
        .din(new_Jinkela_wire_7226),
        .dout(new_Jinkela_wire_7227)
    );

    bfr new_Jinkela_buffer_9168 (
        .din(new_Jinkela_wire_11187),
        .dout(new_Jinkela_wire_11188)
    );

    bfr new_Jinkela_buffer_12645 (
        .din(new_Jinkela_wire_15160),
        .dout(new_Jinkela_wire_15161)
    );

    bfr new_Jinkela_buffer_16056 (
        .din(new_Jinkela_wire_19170),
        .dout(new_Jinkela_wire_19171)
    );

    bfr new_Jinkela_buffer_5731 (
        .din(new_Jinkela_wire_7312),
        .dout(new_Jinkela_wire_7313)
    );

    bfr new_Jinkela_buffer_9327 (
        .din(new_Jinkela_wire_11356),
        .dout(new_Jinkela_wire_11357)
    );

    bfr new_Jinkela_buffer_12596 (
        .din(new_Jinkela_wire_15103),
        .dout(new_Jinkela_wire_15104)
    );

    spl2 new_Jinkela_splitter_643 (
        .a(_0808_),
        .b(new_Jinkela_wire_7320),
        .c(new_Jinkela_wire_7321)
    );

    spl2 new_Jinkela_splitter_1412 (
        .a(_1133_),
        .b(new_Jinkela_wire_19274),
        .c(new_Jinkela_wire_19275)
    );

    bfr new_Jinkela_buffer_5674 (
        .din(new_Jinkela_wire_7227),
        .dout(new_Jinkela_wire_7228)
    );

    bfr new_Jinkela_buffer_9169 (
        .din(new_Jinkela_wire_11188),
        .dout(new_Jinkela_wire_11189)
    );

    bfr new_Jinkela_buffer_16057 (
        .din(new_Jinkela_wire_19171),
        .dout(new_Jinkela_wire_19172)
    );

    bfr new_Jinkela_buffer_9233 (
        .din(new_Jinkela_wire_11256),
        .dout(new_Jinkela_wire_11257)
    );

    bfr new_Jinkela_buffer_12597 (
        .din(new_Jinkela_wire_15104),
        .dout(new_Jinkela_wire_15105)
    );

    bfr new_Jinkela_buffer_16068 (
        .din(new_Jinkela_wire_19192),
        .dout(new_Jinkela_wire_19193)
    );

    bfr new_Jinkela_buffer_5675 (
        .din(new_Jinkela_wire_7228),
        .dout(new_Jinkela_wire_7229)
    );

    bfr new_Jinkela_buffer_9170 (
        .din(new_Jinkela_wire_11189),
        .dout(new_Jinkela_wire_11190)
    );

    bfr new_Jinkela_buffer_12646 (
        .din(new_Jinkela_wire_15161),
        .dout(new_Jinkela_wire_15162)
    );

    bfr new_Jinkela_buffer_16058 (
        .din(new_Jinkela_wire_19172),
        .dout(new_Jinkela_wire_19173)
    );

    spl2 new_Jinkela_splitter_640 (
        .a(new_Jinkela_wire_7313),
        .b(new_Jinkela_wire_7314),
        .c(new_Jinkela_wire_7315)
    );

    bfr new_Jinkela_buffer_9356 (
        .din(_1002_),
        .dout(new_Jinkela_wire_11400)
    );

    bfr new_Jinkela_buffer_12598 (
        .din(new_Jinkela_wire_15105),
        .dout(new_Jinkela_wire_15106)
    );

    bfr new_Jinkela_buffer_9355 (
        .din(_0977_),
        .dout(new_Jinkela_wire_11399)
    );

    spl2 new_Jinkela_splitter_1414 (
        .a(_1413_),
        .b(new_Jinkela_wire_19282),
        .c(new_Jinkela_wire_19283)
    );

    bfr new_Jinkela_buffer_5676 (
        .din(new_Jinkela_wire_7229),
        .dout(new_Jinkela_wire_7230)
    );

    bfr new_Jinkela_buffer_9171 (
        .din(new_Jinkela_wire_11190),
        .dout(new_Jinkela_wire_11191)
    );

    spl2 new_Jinkela_splitter_1113 (
        .a(_1399_),
        .b(new_Jinkela_wire_15521),
        .c(new_Jinkela_wire_15522)
    );

    bfr new_Jinkela_buffer_12701 (
        .din(new_Jinkela_wire_15222),
        .dout(new_Jinkela_wire_15223)
    );

    bfr new_Jinkela_buffer_16059 (
        .din(new_Jinkela_wire_19173),
        .dout(new_Jinkela_wire_19174)
    );

    and_ii _3130_ (
        .a(new_Jinkela_wire_19187),
        .b(new_Jinkela_wire_21181),
        .c(_0391_)
    );

    and_bb _3131_ (
        .a(new_Jinkela_wire_19188),
        .b(new_Jinkela_wire_21182),
        .c(_0392_)
    );

    or_bb _3132_ (
        .a(new_Jinkela_wire_20366),
        .b(new_Jinkela_wire_8095),
        .c(_0393_)
    );

    and_ii _3133_ (
        .a(new_Jinkela_wire_11827),
        .b(new_Jinkela_wire_19272),
        .c(_0395_)
    );

    and_bb _3134_ (
        .a(new_Jinkela_wire_11828),
        .b(new_Jinkela_wire_19273),
        .c(_0396_)
    );

    or_bb _3135_ (
        .a(new_Jinkela_wire_21202),
        .b(new_Jinkela_wire_15781),
        .c(_0397_)
    );

    and_ii _3136_ (
        .a(new_Jinkela_wire_14286),
        .b(new_Jinkela_wire_7184),
        .c(_0398_)
    );

    and_bb _3137_ (
        .a(new_Jinkela_wire_14287),
        .b(new_Jinkela_wire_7185),
        .c(_0399_)
    );

    or_bb _3138_ (
        .a(new_Jinkela_wire_13197),
        .b(new_Jinkela_wire_17005),
        .c(_0400_)
    );

    and_ii _3139_ (
        .a(new_Jinkela_wire_14660),
        .b(new_Jinkela_wire_16100),
        .c(_0401_)
    );

    and_bb _3140_ (
        .a(new_Jinkela_wire_14661),
        .b(new_Jinkela_wire_16101),
        .c(_0402_)
    );

    or_bb _3141_ (
        .a(new_Jinkela_wire_9859),
        .b(new_Jinkela_wire_1259),
        .c(_0403_)
    );

    and_ii _3142_ (
        .a(new_Jinkela_wire_11955),
        .b(new_Jinkela_wire_14034),
        .c(_0404_)
    );

    and_bb _3143_ (
        .a(new_Jinkela_wire_11956),
        .b(new_Jinkela_wire_14035),
        .c(_0406_)
    );

    or_bb _3144_ (
        .a(new_Jinkela_wire_833),
        .b(new_Jinkela_wire_20375),
        .c(_0407_)
    );

    and_ii _3145_ (
        .a(new_Jinkela_wire_6240),
        .b(new_Jinkela_wire_4824),
        .c(_0408_)
    );

    and_bb _3146_ (
        .a(new_Jinkela_wire_6241),
        .b(new_Jinkela_wire_4825),
        .c(_0409_)
    );

    or_bb _3147_ (
        .a(new_Jinkela_wire_13307),
        .b(new_Jinkela_wire_13582),
        .c(_0410_)
    );

    and_ii _3148_ (
        .a(new_Jinkela_wire_5441),
        .b(new_Jinkela_wire_11531),
        .c(_0411_)
    );

    and_bb _3149_ (
        .a(new_Jinkela_wire_5442),
        .b(new_Jinkela_wire_11532),
        .c(_0412_)
    );

    or_bb _3150_ (
        .a(new_Jinkela_wire_19184),
        .b(new_Jinkela_wire_16436),
        .c(_0413_)
    );

    and_ii _3151_ (
        .a(new_Jinkela_wire_11414),
        .b(new_Jinkela_wire_15660),
        .c(_0414_)
    );

    and_bb _3152_ (
        .a(new_Jinkela_wire_11415),
        .b(new_Jinkela_wire_15661),
        .c(_0415_)
    );

    or_bb _3153_ (
        .a(new_Jinkela_wire_7982),
        .b(new_Jinkela_wire_4673),
        .c(_0417_)
    );

    and_ii _3154_ (
        .a(new_Jinkela_wire_12054),
        .b(new_Jinkela_wire_16943),
        .c(_0418_)
    );

    and_bb _3155_ (
        .a(new_Jinkela_wire_12055),
        .b(new_Jinkela_wire_16944),
        .c(_0419_)
    );

    or_bb _3156_ (
        .a(new_Jinkela_wire_16508),
        .b(new_Jinkela_wire_18516),
        .c(_0420_)
    );

    and_ii _3157_ (
        .a(new_Jinkela_wire_13722),
        .b(new_Jinkela_wire_16330),
        .c(_0421_)
    );

    and_bb _3158_ (
        .a(new_Jinkela_wire_13723),
        .b(new_Jinkela_wire_16331),
        .c(_0422_)
    );

    or_bb _3159_ (
        .a(new_Jinkela_wire_3816),
        .b(new_Jinkela_wire_14683),
        .c(_0423_)
    );

    and_ii _3160_ (
        .a(new_Jinkela_wire_7746),
        .b(new_Jinkela_wire_1619),
        .c(_0424_)
    );

    and_bb _3161_ (
        .a(new_Jinkela_wire_7747),
        .b(new_Jinkela_wire_1620),
        .c(_0425_)
    );

    or_bb _3162_ (
        .a(new_Jinkela_wire_9096),
        .b(new_Jinkela_wire_5667),
        .c(_0426_)
    );

    and_bi _3163_ (
        .a(new_Jinkela_wire_20283),
        .b(new_Jinkela_wire_10273),
        .c(_0428_)
    );

    and_bi _3164_ (
        .a(new_Jinkela_wire_10274),
        .b(new_Jinkela_wire_20284),
        .c(_0429_)
    );

    or_bb _3165_ (
        .a(new_Jinkela_wire_18807),
        .b(new_Jinkela_wire_4283),
        .c(new_net_3934)
    );

    or_bb _3166_ (
        .a(new_Jinkela_wire_4284),
        .b(new_Jinkela_wire_5680),
        .c(_0430_)
    );

    and_ii _3167_ (
        .a(new_Jinkela_wire_14684),
        .b(new_Jinkela_wire_18521),
        .c(_0431_)
    );

    and_bb _3168_ (
        .a(new_Jinkela_wire_475),
        .b(new_Jinkela_wire_675),
        .c(_0432_)
    );

    and_ii _3169_ (
        .a(new_Jinkela_wire_4674),
        .b(new_Jinkela_wire_16441),
        .c(_0433_)
    );

    and_bb _3170_ (
        .a(new_Jinkela_wire_354),
        .b(new_Jinkela_wire_515),
        .c(_0434_)
    );

    and_ii _3171_ (
        .a(new_Jinkela_wire_13583),
        .b(new_Jinkela_wire_20380),
        .c(_0435_)
    );

    bfr new_Jinkela_buffer_2072 (
        .din(new_Jinkela_wire_3013),
        .dout(new_Jinkela_wire_3014)
    );

    bfr new_Jinkela_buffer_2194 (
        .din(new_Jinkela_wire_3143),
        .dout(new_Jinkela_wire_3144)
    );

    bfr new_Jinkela_buffer_2073 (
        .din(new_Jinkela_wire_3014),
        .dout(new_Jinkela_wire_3015)
    );

    bfr new_Jinkela_buffer_2074 (
        .din(new_Jinkela_wire_3015),
        .dout(new_Jinkela_wire_3016)
    );

    bfr new_Jinkela_buffer_2195 (
        .din(new_Jinkela_wire_3144),
        .dout(new_Jinkela_wire_3145)
    );

    bfr new_Jinkela_buffer_2075 (
        .din(new_Jinkela_wire_3016),
        .dout(new_Jinkela_wire_3017)
    );

    bfr new_Jinkela_buffer_2235 (
        .din(new_Jinkela_wire_3200),
        .dout(new_Jinkela_wire_3201)
    );

    bfr new_Jinkela_buffer_2076 (
        .din(new_Jinkela_wire_3017),
        .dout(new_Jinkela_wire_3018)
    );

    bfr new_Jinkela_buffer_2196 (
        .din(new_Jinkela_wire_3145),
        .dout(new_Jinkela_wire_3146)
    );

    bfr new_Jinkela_buffer_2077 (
        .din(new_Jinkela_wire_3018),
        .dout(new_Jinkela_wire_3019)
    );

    spl2 new_Jinkela_splitter_333 (
        .a(new_Jinkela_wire_3240),
        .b(new_Jinkela_wire_3241),
        .c(new_Jinkela_wire_3242)
    );

    bfr new_Jinkela_buffer_2078 (
        .din(new_Jinkela_wire_3019),
        .dout(new_Jinkela_wire_3020)
    );

    bfr new_Jinkela_buffer_2197 (
        .din(new_Jinkela_wire_3146),
        .dout(new_Jinkela_wire_3147)
    );

    bfr new_Jinkela_buffer_2079 (
        .din(new_Jinkela_wire_3020),
        .dout(new_Jinkela_wire_3021)
    );

    bfr new_Jinkela_buffer_2236 (
        .din(new_Jinkela_wire_3201),
        .dout(new_Jinkela_wire_3202)
    );

    bfr new_Jinkela_buffer_2080 (
        .din(new_Jinkela_wire_3021),
        .dout(new_Jinkela_wire_3022)
    );

    bfr new_Jinkela_buffer_2198 (
        .din(new_Jinkela_wire_3147),
        .dout(new_Jinkela_wire_3148)
    );

    bfr new_Jinkela_buffer_2081 (
        .din(new_Jinkela_wire_3022),
        .dout(new_Jinkela_wire_3023)
    );

    bfr new_Jinkela_buffer_2082 (
        .din(new_Jinkela_wire_3023),
        .dout(new_Jinkela_wire_3024)
    );

    spl2 new_Jinkela_splitter_337 (
        .a(_0021_),
        .b(new_Jinkela_wire_3253),
        .c(new_Jinkela_wire_3254)
    );

    bfr new_Jinkela_buffer_2199 (
        .din(new_Jinkela_wire_3148),
        .dout(new_Jinkela_wire_3149)
    );

    bfr new_Jinkela_buffer_2083 (
        .din(new_Jinkela_wire_3024),
        .dout(new_Jinkela_wire_3025)
    );

    bfr new_Jinkela_buffer_2237 (
        .din(new_Jinkela_wire_3202),
        .dout(new_Jinkela_wire_3203)
    );

    bfr new_Jinkela_buffer_2084 (
        .din(new_Jinkela_wire_3025),
        .dout(new_Jinkela_wire_3026)
    );

    bfr new_Jinkela_buffer_2200 (
        .din(new_Jinkela_wire_3149),
        .dout(new_Jinkela_wire_3150)
    );

    bfr new_Jinkela_buffer_2085 (
        .din(new_Jinkela_wire_3026),
        .dout(new_Jinkela_wire_3027)
    );

    bfr new_Jinkela_buffer_2086 (
        .din(new_Jinkela_wire_3027),
        .dout(new_Jinkela_wire_3028)
    );

    spl2 new_Jinkela_splitter_336 (
        .a(_0180_),
        .b(new_Jinkela_wire_3247),
        .c(new_Jinkela_wire_3248)
    );

    bfr new_Jinkela_buffer_2201 (
        .din(new_Jinkela_wire_3150),
        .dout(new_Jinkela_wire_3151)
    );

    bfr new_Jinkela_buffer_2087 (
        .din(new_Jinkela_wire_3028),
        .dout(new_Jinkela_wire_3029)
    );

    bfr new_Jinkela_buffer_2238 (
        .din(new_Jinkela_wire_3203),
        .dout(new_Jinkela_wire_3204)
    );

    bfr new_Jinkela_buffer_2088 (
        .din(new_Jinkela_wire_3029),
        .dout(new_Jinkela_wire_3030)
    );

    bfr new_Jinkela_buffer_2202 (
        .din(new_Jinkela_wire_3151),
        .dout(new_Jinkela_wire_3152)
    );

    bfr new_Jinkela_buffer_2089 (
        .din(new_Jinkela_wire_3030),
        .dout(new_Jinkela_wire_3031)
    );

    bfr new_Jinkela_buffer_2273 (
        .din(new_Jinkela_wire_3248),
        .dout(new_Jinkela_wire_3249)
    );

    bfr new_Jinkela_buffer_2090 (
        .din(new_Jinkela_wire_3031),
        .dout(new_Jinkela_wire_3032)
    );

    spl2 new_Jinkela_splitter_338 (
        .a(_1254_),
        .b(new_Jinkela_wire_3255),
        .c(new_Jinkela_wire_3256)
    );

    bfr new_Jinkela_buffer_2203 (
        .din(new_Jinkela_wire_3152),
        .dout(new_Jinkela_wire_3153)
    );

    bfr new_Jinkela_buffer_2091 (
        .din(new_Jinkela_wire_3032),
        .dout(new_Jinkela_wire_3033)
    );

    bfr new_Jinkela_buffer_2239 (
        .din(new_Jinkela_wire_3204),
        .dout(new_Jinkela_wire_3205)
    );

    bfr new_Jinkela_buffer_2092 (
        .din(new_Jinkela_wire_3033),
        .dout(new_Jinkela_wire_3034)
    );

    bfr new_Jinkela_buffer_2234 (
        .din(new_Jinkela_wire_3199),
        .dout(new_Jinkela_wire_3200)
    );

    bfr new_Jinkela_buffer_2204 (
        .din(new_Jinkela_wire_3153),
        .dout(new_Jinkela_wire_3154)
    );

    bfr new_Jinkela_buffer_12599 (
        .din(new_Jinkela_wire_15106),
        .dout(new_Jinkela_wire_15107)
    );

    bfr new_Jinkela_buffer_5736 (
        .din(_0084_),
        .dout(new_Jinkela_wire_7326)
    );

    bfr new_Jinkela_buffer_5677 (
        .din(new_Jinkela_wire_7230),
        .dout(new_Jinkela_wire_7231)
    );

    bfr new_Jinkela_buffer_12647 (
        .din(new_Jinkela_wire_15162),
        .dout(new_Jinkela_wire_15163)
    );

    bfr new_Jinkela_buffer_12600 (
        .din(new_Jinkela_wire_15107),
        .dout(new_Jinkela_wire_15108)
    );

    bfr new_Jinkela_buffer_5678 (
        .din(new_Jinkela_wire_7231),
        .dout(new_Jinkela_wire_7232)
    );

    bfr new_Jinkela_buffer_12865 (
        .din(new_Jinkela_wire_15386),
        .dout(new_Jinkela_wire_15387)
    );

    bfr new_Jinkela_buffer_5732 (
        .din(new_Jinkela_wire_7321),
        .dout(new_Jinkela_wire_7322)
    );

    bfr new_Jinkela_buffer_12601 (
        .din(new_Jinkela_wire_15108),
        .dout(new_Jinkela_wire_15109)
    );

    spl2 new_Jinkela_splitter_645 (
        .a(_1724_),
        .b(new_Jinkela_wire_7440),
        .c(new_Jinkela_wire_7441)
    );

    bfr new_Jinkela_buffer_5679 (
        .din(new_Jinkela_wire_7232),
        .dout(new_Jinkela_wire_7233)
    );

    bfr new_Jinkela_buffer_12648 (
        .din(new_Jinkela_wire_15163),
        .dout(new_Jinkela_wire_15164)
    );

    bfr new_Jinkela_buffer_12602 (
        .din(new_Jinkela_wire_15109),
        .dout(new_Jinkela_wire_15110)
    );

    bfr new_Jinkela_buffer_5848 (
        .din(_0303_),
        .dout(new_Jinkela_wire_7442)
    );

    bfr new_Jinkela_buffer_5680 (
        .din(new_Jinkela_wire_7233),
        .dout(new_Jinkela_wire_7234)
    );

    bfr new_Jinkela_buffer_12702 (
        .din(new_Jinkela_wire_15223),
        .dout(new_Jinkela_wire_15224)
    );

    bfr new_Jinkela_buffer_5733 (
        .din(new_Jinkela_wire_7322),
        .dout(new_Jinkela_wire_7323)
    );

    bfr new_Jinkela_buffer_12603 (
        .din(new_Jinkela_wire_15110),
        .dout(new_Jinkela_wire_15111)
    );

    bfr new_Jinkela_buffer_5681 (
        .din(new_Jinkela_wire_7234),
        .dout(new_Jinkela_wire_7235)
    );

    bfr new_Jinkela_buffer_12649 (
        .din(new_Jinkela_wire_15164),
        .dout(new_Jinkela_wire_15165)
    );

    bfr new_Jinkela_buffer_5737 (
        .din(new_Jinkela_wire_7326),
        .dout(new_Jinkela_wire_7327)
    );

    bfr new_Jinkela_buffer_12604 (
        .din(new_Jinkela_wire_15111),
        .dout(new_Jinkela_wire_15112)
    );

    bfr new_Jinkela_buffer_5682 (
        .din(new_Jinkela_wire_7235),
        .dout(new_Jinkela_wire_7236)
    );

    bfr new_Jinkela_buffer_12947 (
        .din(new_Jinkela_wire_15470),
        .dout(new_Jinkela_wire_15471)
    );

    bfr new_Jinkela_buffer_5734 (
        .din(new_Jinkela_wire_7323),
        .dout(new_Jinkela_wire_7324)
    );

    bfr new_Jinkela_buffer_12605 (
        .din(new_Jinkela_wire_15112),
        .dout(new_Jinkela_wire_15113)
    );

    bfr new_Jinkela_buffer_5683 (
        .din(new_Jinkela_wire_7236),
        .dout(new_Jinkela_wire_7237)
    );

    bfr new_Jinkela_buffer_12650 (
        .din(new_Jinkela_wire_15165),
        .dout(new_Jinkela_wire_15166)
    );

    bfr new_Jinkela_buffer_12606 (
        .din(new_Jinkela_wire_15113),
        .dout(new_Jinkela_wire_15114)
    );

    bfr new_Jinkela_buffer_5684 (
        .din(new_Jinkela_wire_7237),
        .dout(new_Jinkela_wire_7238)
    );

    bfr new_Jinkela_buffer_12877 (
        .din(new_Jinkela_wire_15398),
        .dout(new_Jinkela_wire_15399)
    );

    bfr new_Jinkela_buffer_12703 (
        .din(new_Jinkela_wire_15224),
        .dout(new_Jinkela_wire_15225)
    );

    bfr new_Jinkela_buffer_5735 (
        .din(new_Jinkela_wire_7324),
        .dout(new_Jinkela_wire_7325)
    );

    bfr new_Jinkela_buffer_12607 (
        .din(new_Jinkela_wire_15114),
        .dout(new_Jinkela_wire_15115)
    );

    bfr new_Jinkela_buffer_5685 (
        .din(new_Jinkela_wire_7238),
        .dout(new_Jinkela_wire_7239)
    );

    bfr new_Jinkela_buffer_12651 (
        .din(new_Jinkela_wire_15166),
        .dout(new_Jinkela_wire_15167)
    );

    bfr new_Jinkela_buffer_5738 (
        .din(new_Jinkela_wire_7327),
        .dout(new_Jinkela_wire_7328)
    );

    bfr new_Jinkela_buffer_12608 (
        .din(new_Jinkela_wire_15115),
        .dout(new_Jinkela_wire_15116)
    );

    bfr new_Jinkela_buffer_5686 (
        .din(new_Jinkela_wire_7239),
        .dout(new_Jinkela_wire_7240)
    );

    bfr new_Jinkela_buffer_12866 (
        .din(new_Jinkela_wire_15387),
        .dout(new_Jinkela_wire_15388)
    );

    spl2 new_Jinkela_splitter_647 (
        .a(_0031_),
        .b(new_Jinkela_wire_7445),
        .c(new_Jinkela_wire_7446)
    );

    spl2 new_Jinkela_splitter_1103 (
        .a(new_Jinkela_wire_15116),
        .b(new_Jinkela_wire_15117),
        .c(new_Jinkela_wire_15118)
    );

    spl2 new_Jinkela_splitter_646 (
        .a(_1416_),
        .b(new_Jinkela_wire_7443),
        .c(new_Jinkela_wire_7444)
    );

    bfr new_Jinkela_buffer_5687 (
        .din(new_Jinkela_wire_7240),
        .dout(new_Jinkela_wire_7241)
    );

    bfr new_Jinkela_buffer_12704 (
        .din(new_Jinkela_wire_15225),
        .dout(new_Jinkela_wire_15226)
    );

    bfr new_Jinkela_buffer_5739 (
        .din(new_Jinkela_wire_7328),
        .dout(new_Jinkela_wire_7329)
    );

    bfr new_Jinkela_buffer_12652 (
        .din(new_Jinkela_wire_15167),
        .dout(new_Jinkela_wire_15168)
    );

    bfr new_Jinkela_buffer_5688 (
        .din(new_Jinkela_wire_7241),
        .dout(new_Jinkela_wire_7242)
    );

    bfr new_Jinkela_buffer_12653 (
        .din(new_Jinkela_wire_15168),
        .dout(new_Jinkela_wire_15169)
    );

    bfr new_Jinkela_buffer_5689 (
        .din(new_Jinkela_wire_7242),
        .dout(new_Jinkela_wire_7243)
    );

    bfr new_Jinkela_buffer_12654 (
        .din(new_Jinkela_wire_15169),
        .dout(new_Jinkela_wire_15170)
    );

    bfr new_Jinkela_buffer_5740 (
        .din(new_Jinkela_wire_7329),
        .dout(new_Jinkela_wire_7330)
    );

    bfr new_Jinkela_buffer_12705 (
        .din(new_Jinkela_wire_15226),
        .dout(new_Jinkela_wire_15227)
    );

    bfr new_Jinkela_buffer_5690 (
        .din(new_Jinkela_wire_7243),
        .dout(new_Jinkela_wire_7244)
    );

    bfr new_Jinkela_buffer_12655 (
        .din(new_Jinkela_wire_15170),
        .dout(new_Jinkela_wire_15171)
    );

    bfr new_Jinkela_buffer_5853 (
        .din(_1095_),
        .dout(new_Jinkela_wire_7451)
    );

    bfr new_Jinkela_buffer_12867 (
        .din(new_Jinkela_wire_15388),
        .dout(new_Jinkela_wire_15389)
    );

    bfr new_Jinkela_buffer_5691 (
        .din(new_Jinkela_wire_7244),
        .dout(new_Jinkela_wire_7245)
    );

    bfr new_Jinkela_buffer_12656 (
        .din(new_Jinkela_wire_15171),
        .dout(new_Jinkela_wire_15172)
    );

    bfr new_Jinkela_buffer_5741 (
        .din(new_Jinkela_wire_7330),
        .dout(new_Jinkela_wire_7331)
    );

    bfr new_Jinkela_buffer_12706 (
        .din(new_Jinkela_wire_15227),
        .dout(new_Jinkela_wire_15228)
    );

    bfr new_Jinkela_buffer_5692 (
        .din(new_Jinkela_wire_7245),
        .dout(new_Jinkela_wire_7246)
    );

    bfr new_Jinkela_buffer_12657 (
        .din(new_Jinkela_wire_15172),
        .dout(new_Jinkela_wire_15173)
    );

    bfr new_Jinkela_buffer_5849 (
        .din(new_Jinkela_wire_7446),
        .dout(new_Jinkela_wire_7447)
    );

    bfr new_Jinkela_buffer_5854 (
        .din(_1067_),
        .dout(new_Jinkela_wire_7452)
    );

    spl2 new_Jinkela_splitter_1112 (
        .a(_1408_),
        .b(new_Jinkela_wire_15519),
        .c(new_Jinkela_wire_15520)
    );

    bfr new_Jinkela_buffer_5693 (
        .din(new_Jinkela_wire_7246),
        .dout(new_Jinkela_wire_7247)
    );

    bfr new_Jinkela_buffer_12658 (
        .din(new_Jinkela_wire_15173),
        .dout(new_Jinkela_wire_15174)
    );

    bfr new_Jinkela_buffer_5742 (
        .din(new_Jinkela_wire_7331),
        .dout(new_Jinkela_wire_7332)
    );

    bfr new_Jinkela_buffer_12878 (
        .din(new_Jinkela_wire_15399),
        .dout(new_Jinkela_wire_15400)
    );

    bfr new_Jinkela_buffer_12707 (
        .din(new_Jinkela_wire_15228),
        .dout(new_Jinkela_wire_15229)
    );

    bfr new_Jinkela_buffer_5694 (
        .din(new_Jinkela_wire_7247),
        .dout(new_Jinkela_wire_7248)
    );

    bfr new_Jinkela_buffer_12659 (
        .din(new_Jinkela_wire_15174),
        .dout(new_Jinkela_wire_15175)
    );

    spl2 new_Jinkela_splitter_649 (
        .a(_0827_),
        .b(new_Jinkela_wire_7502),
        .c(new_Jinkela_wire_7503)
    );

    bfr new_Jinkela_buffer_12868 (
        .din(new_Jinkela_wire_15389),
        .dout(new_Jinkela_wire_15390)
    );

    bfr new_Jinkela_buffer_5695 (
        .din(new_Jinkela_wire_7248),
        .dout(new_Jinkela_wire_7249)
    );

    bfr new_Jinkela_buffer_12660 (
        .din(new_Jinkela_wire_15175),
        .dout(new_Jinkela_wire_15176)
    );

    bfr new_Jinkela_buffer_5743 (
        .din(new_Jinkela_wire_7332),
        .dout(new_Jinkela_wire_7333)
    );

    bfr new_Jinkela_buffer_12708 (
        .din(new_Jinkela_wire_15229),
        .dout(new_Jinkela_wire_15230)
    );

    bfr new_Jinkela_buffer_5696 (
        .din(new_Jinkela_wire_7249),
        .dout(new_Jinkela_wire_7250)
    );

    bfr new_Jinkela_buffer_12661 (
        .din(new_Jinkela_wire_15176),
        .dout(new_Jinkela_wire_15177)
    );

    bfr new_Jinkela_buffer_5850 (
        .din(new_Jinkela_wire_7447),
        .dout(new_Jinkela_wire_7448)
    );

    bfr new_Jinkela_buffer_5697 (
        .din(new_Jinkela_wire_7250),
        .dout(new_Jinkela_wire_7251)
    );

    bfr new_Jinkela_buffer_12662 (
        .din(new_Jinkela_wire_15177),
        .dout(new_Jinkela_wire_15178)
    );

    bfr new_Jinkela_buffer_2093 (
        .din(new_Jinkela_wire_3034),
        .dout(new_Jinkela_wire_3035)
    );

    bfr new_Jinkela_buffer_16069 (
        .din(new_Jinkela_wire_19193),
        .dout(new_Jinkela_wire_19194)
    );

    bfr new_Jinkela_buffer_16060 (
        .din(new_Jinkela_wire_19174),
        .dout(new_Jinkela_wire_19175)
    );

    bfr new_Jinkela_buffer_2242 (
        .din(new_Jinkela_wire_3207),
        .dout(new_Jinkela_wire_3208)
    );

    bfr new_Jinkela_buffer_2094 (
        .din(new_Jinkela_wire_3035),
        .dout(new_Jinkela_wire_3036)
    );

    bfr new_Jinkela_buffer_16147 (
        .din(new_Jinkela_wire_19277),
        .dout(new_Jinkela_wire_19278)
    );

    bfr new_Jinkela_buffer_16061 (
        .din(new_Jinkela_wire_19175),
        .dout(new_Jinkela_wire_19176)
    );

    bfr new_Jinkela_buffer_2205 (
        .din(new_Jinkela_wire_3154),
        .dout(new_Jinkela_wire_3155)
    );

    bfr new_Jinkela_buffer_2095 (
        .din(new_Jinkela_wire_3036),
        .dout(new_Jinkela_wire_3037)
    );

    bfr new_Jinkela_buffer_16070 (
        .din(new_Jinkela_wire_19194),
        .dout(new_Jinkela_wire_19195)
    );

    bfr new_Jinkela_buffer_16062 (
        .din(new_Jinkela_wire_19176),
        .dout(new_Jinkela_wire_19177)
    );

    bfr new_Jinkela_buffer_2275 (
        .din(new_Jinkela_wire_3250),
        .dout(new_Jinkela_wire_3251)
    );

    bfr new_Jinkela_buffer_2096 (
        .din(new_Jinkela_wire_3037),
        .dout(new_Jinkela_wire_3038)
    );

    spl2 new_Jinkela_splitter_1415 (
        .a(_1593_),
        .b(new_Jinkela_wire_19284),
        .c(new_Jinkela_wire_19285)
    );

    bfr new_Jinkela_buffer_16063 (
        .din(new_Jinkela_wire_19177),
        .dout(new_Jinkela_wire_19178)
    );

    bfr new_Jinkela_buffer_2206 (
        .din(new_Jinkela_wire_3155),
        .dout(new_Jinkela_wire_3156)
    );

    bfr new_Jinkela_buffer_2097 (
        .din(new_Jinkela_wire_3038),
        .dout(new_Jinkela_wire_3039)
    );

    bfr new_Jinkela_buffer_16071 (
        .din(new_Jinkela_wire_19195),
        .dout(new_Jinkela_wire_19196)
    );

    bfr new_Jinkela_buffer_16064 (
        .din(new_Jinkela_wire_19178),
        .dout(new_Jinkela_wire_19179)
    );

    bfr new_Jinkela_buffer_2243 (
        .din(new_Jinkela_wire_3208),
        .dout(new_Jinkela_wire_3209)
    );

    bfr new_Jinkela_buffer_2098 (
        .din(new_Jinkela_wire_3039),
        .dout(new_Jinkela_wire_3040)
    );

    spl2 new_Jinkela_splitter_1406 (
        .a(new_Jinkela_wire_19179),
        .b(new_Jinkela_wire_19180),
        .c(new_Jinkela_wire_19181)
    );

    bfr new_Jinkela_buffer_2207 (
        .din(new_Jinkela_wire_3156),
        .dout(new_Jinkela_wire_3157)
    );

    bfr new_Jinkela_buffer_2099 (
        .din(new_Jinkela_wire_3040),
        .dout(new_Jinkela_wire_3041)
    );

    bfr new_Jinkela_buffer_16148 (
        .din(new_Jinkela_wire_19278),
        .dout(new_Jinkela_wire_19279)
    );

    bfr new_Jinkela_buffer_16072 (
        .din(new_Jinkela_wire_19196),
        .dout(new_Jinkela_wire_19197)
    );

    bfr new_Jinkela_buffer_2278 (
        .din(_0610_),
        .dout(new_Jinkela_wire_3260)
    );

    bfr new_Jinkela_buffer_2100 (
        .din(new_Jinkela_wire_3041),
        .dout(new_Jinkela_wire_3042)
    );

    bfr new_Jinkela_buffer_16073 (
        .din(new_Jinkela_wire_19197),
        .dout(new_Jinkela_wire_19198)
    );

    spl2 new_Jinkela_splitter_341 (
        .a(_1281_),
        .b(new_Jinkela_wire_3269),
        .c(new_Jinkela_wire_3270)
    );

    bfr new_Jinkela_buffer_2208 (
        .din(new_Jinkela_wire_3157),
        .dout(new_Jinkela_wire_3158)
    );

    spl2 new_Jinkela_splitter_1416 (
        .a(_0905_),
        .b(new_Jinkela_wire_19290),
        .c(new_Jinkela_wire_19291)
    );

    bfr new_Jinkela_buffer_2101 (
        .din(new_Jinkela_wire_3042),
        .dout(new_Jinkela_wire_3043)
    );

    bfr new_Jinkela_buffer_16074 (
        .din(new_Jinkela_wire_19198),
        .dout(new_Jinkela_wire_19199)
    );

    bfr new_Jinkela_buffer_16149 (
        .din(new_Jinkela_wire_19279),
        .dout(new_Jinkela_wire_19280)
    );

    bfr new_Jinkela_buffer_2244 (
        .din(new_Jinkela_wire_3209),
        .dout(new_Jinkela_wire_3210)
    );

    bfr new_Jinkela_buffer_2102 (
        .din(new_Jinkela_wire_3043),
        .dout(new_Jinkela_wire_3044)
    );

    bfr new_Jinkela_buffer_16075 (
        .din(new_Jinkela_wire_19199),
        .dout(new_Jinkela_wire_19200)
    );

    bfr new_Jinkela_buffer_16151 (
        .din(new_Jinkela_wire_19285),
        .dout(new_Jinkela_wire_19286)
    );

    bfr new_Jinkela_buffer_2209 (
        .din(new_Jinkela_wire_3158),
        .dout(new_Jinkela_wire_3159)
    );

    spl2 new_Jinkela_splitter_1417 (
        .a(_1519_),
        .b(new_Jinkela_wire_19296),
        .c(new_Jinkela_wire_19297)
    );

    bfr new_Jinkela_buffer_2103 (
        .din(new_Jinkela_wire_3044),
        .dout(new_Jinkela_wire_3045)
    );

    bfr new_Jinkela_buffer_16076 (
        .din(new_Jinkela_wire_19200),
        .dout(new_Jinkela_wire_19201)
    );

    bfr new_Jinkela_buffer_16150 (
        .din(new_Jinkela_wire_19280),
        .dout(new_Jinkela_wire_19281)
    );

    bfr new_Jinkela_buffer_2276 (
        .din(new_Jinkela_wire_3251),
        .dout(new_Jinkela_wire_3252)
    );

    bfr new_Jinkela_buffer_2104 (
        .din(new_Jinkela_wire_3045),
        .dout(new_Jinkela_wire_3046)
    );

    bfr new_Jinkela_buffer_16077 (
        .din(new_Jinkela_wire_19201),
        .dout(new_Jinkela_wire_19202)
    );

    bfr new_Jinkela_buffer_2210 (
        .din(new_Jinkela_wire_3159),
        .dout(new_Jinkela_wire_3160)
    );

    bfr new_Jinkela_buffer_2105 (
        .din(new_Jinkela_wire_3046),
        .dout(new_Jinkela_wire_3047)
    );

    bfr new_Jinkela_buffer_16078 (
        .din(new_Jinkela_wire_19202),
        .dout(new_Jinkela_wire_19203)
    );

    bfr new_Jinkela_buffer_16152 (
        .din(new_Jinkela_wire_19286),
        .dout(new_Jinkela_wire_19287)
    );

    bfr new_Jinkela_buffer_2245 (
        .din(new_Jinkela_wire_3210),
        .dout(new_Jinkela_wire_3211)
    );

    bfr new_Jinkela_buffer_2106 (
        .din(new_Jinkela_wire_3047),
        .dout(new_Jinkela_wire_3048)
    );

    bfr new_Jinkela_buffer_16079 (
        .din(new_Jinkela_wire_19203),
        .dout(new_Jinkela_wire_19204)
    );

    bfr new_Jinkela_buffer_16155 (
        .din(new_Jinkela_wire_19291),
        .dout(new_Jinkela_wire_19292)
    );

    bfr new_Jinkela_buffer_2211 (
        .din(new_Jinkela_wire_3160),
        .dout(new_Jinkela_wire_3161)
    );

    bfr new_Jinkela_buffer_16159 (
        .din(_0236_),
        .dout(new_Jinkela_wire_19298)
    );

    bfr new_Jinkela_buffer_2107 (
        .din(new_Jinkela_wire_3048),
        .dout(new_Jinkela_wire_3049)
    );

    bfr new_Jinkela_buffer_16080 (
        .din(new_Jinkela_wire_19204),
        .dout(new_Jinkela_wire_19205)
    );

    bfr new_Jinkela_buffer_16153 (
        .din(new_Jinkela_wire_19287),
        .dout(new_Jinkela_wire_19288)
    );

    bfr new_Jinkela_buffer_2108 (
        .din(new_Jinkela_wire_3049),
        .dout(new_Jinkela_wire_3050)
    );

    bfr new_Jinkela_buffer_16081 (
        .din(new_Jinkela_wire_19205),
        .dout(new_Jinkela_wire_19206)
    );

    spl2 new_Jinkela_splitter_1420 (
        .a(_0535_),
        .b(new_Jinkela_wire_19320),
        .c(new_Jinkela_wire_19321)
    );

    bfr new_Jinkela_buffer_2212 (
        .din(new_Jinkela_wire_3161),
        .dout(new_Jinkela_wire_3162)
    );

    bfr new_Jinkela_buffer_2109 (
        .din(new_Jinkela_wire_3050),
        .dout(new_Jinkela_wire_3051)
    );

    bfr new_Jinkela_buffer_16082 (
        .din(new_Jinkela_wire_19206),
        .dout(new_Jinkela_wire_19207)
    );

    bfr new_Jinkela_buffer_16154 (
        .din(new_Jinkela_wire_19288),
        .dout(new_Jinkela_wire_19289)
    );

    bfr new_Jinkela_buffer_2246 (
        .din(new_Jinkela_wire_3211),
        .dout(new_Jinkela_wire_3212)
    );

    bfr new_Jinkela_buffer_2110 (
        .din(new_Jinkela_wire_3051),
        .dout(new_Jinkela_wire_3052)
    );

    bfr new_Jinkela_buffer_16083 (
        .din(new_Jinkela_wire_19207),
        .dout(new_Jinkela_wire_19208)
    );

    bfr new_Jinkela_buffer_16156 (
        .din(new_Jinkela_wire_19292),
        .dout(new_Jinkela_wire_19293)
    );

    bfr new_Jinkela_buffer_2213 (
        .din(new_Jinkela_wire_3162),
        .dout(new_Jinkela_wire_3163)
    );

    bfr new_Jinkela_buffer_2111 (
        .din(new_Jinkela_wire_3052),
        .dout(new_Jinkela_wire_3053)
    );

    bfr new_Jinkela_buffer_16084 (
        .din(new_Jinkela_wire_19208),
        .dout(new_Jinkela_wire_19209)
    );

    spl2 new_Jinkela_splitter_1419 (
        .a(_0712_),
        .b(new_Jinkela_wire_19318),
        .c(new_Jinkela_wire_19319)
    );

    bfr new_Jinkela_buffer_2112 (
        .din(new_Jinkela_wire_3053),
        .dout(new_Jinkela_wire_3054)
    );

    bfr new_Jinkela_buffer_16085 (
        .din(new_Jinkela_wire_19209),
        .dout(new_Jinkela_wire_19210)
    );

    bfr new_Jinkela_buffer_2279 (
        .din(_1706_),
        .dout(new_Jinkela_wire_3261)
    );

    bfr new_Jinkela_buffer_16157 (
        .din(new_Jinkela_wire_19293),
        .dout(new_Jinkela_wire_19294)
    );

    bfr new_Jinkela_buffer_2214 (
        .din(new_Jinkela_wire_3163),
        .dout(new_Jinkela_wire_3164)
    );

    bfr new_Jinkela_buffer_2113 (
        .din(new_Jinkela_wire_3054),
        .dout(new_Jinkela_wire_3055)
    );

    bfr new_Jinkela_buffer_16086 (
        .din(new_Jinkela_wire_19210),
        .dout(new_Jinkela_wire_19211)
    );

    bfr new_Jinkela_buffer_16160 (
        .din(new_Jinkela_wire_19298),
        .dout(new_Jinkela_wire_19299)
    );

    bfr new_Jinkela_buffer_2247 (
        .din(new_Jinkela_wire_3212),
        .dout(new_Jinkela_wire_3213)
    );

    and_bb _3172_ (
        .a(new_Jinkela_wire_699),
        .b(new_Jinkela_wire_134),
        .c(_0436_)
    );

    and_ii _3173_ (
        .a(new_Jinkela_wire_1260),
        .b(new_Jinkela_wire_17010),
        .c(_0438_)
    );

    and_bb _3174_ (
        .a(new_Jinkela_wire_207),
        .b(new_Jinkela_wire_495),
        .c(_0439_)
    );

    and_ii _3175_ (
        .a(new_Jinkela_wire_15782),
        .b(new_Jinkela_wire_8100),
        .c(_0440_)
    );

    and_bb _3176_ (
        .a(new_Jinkela_wire_582),
        .b(new_Jinkela_wire_40),
        .c(_0441_)
    );

    and_ii _3177_ (
        .a(new_Jinkela_wire_2788),
        .b(new_Jinkela_wire_14316),
        .c(_0442_)
    );

    and_bb _3178_ (
        .a(new_Jinkela_wire_181),
        .b(new_Jinkela_wire_112),
        .c(_0443_)
    );

    and_ii _3179_ (
        .a(new_Jinkela_wire_2596),
        .b(new_Jinkela_wire_2134),
        .c(_0444_)
    );

    and_bb _3180_ (
        .a(new_Jinkela_wire_387),
        .b(new_Jinkela_wire_9),
        .c(_0445_)
    );

    and_ii _3181_ (
        .a(new_Jinkela_wire_2712),
        .b(new_Jinkela_wire_19969),
        .c(_0446_)
    );

    and_bb _3182_ (
        .a(new_Jinkela_wire_408),
        .b(new_Jinkela_wire_452),
        .c(_0447_)
    );

    and_ii _3183_ (
        .a(new_Jinkela_wire_14686),
        .b(new_Jinkela_wire_1601),
        .c(_0449_)
    );

    and_bb _3184_ (
        .a(new_Jinkela_wire_153),
        .b(new_Jinkela_wire_256),
        .c(_0450_)
    );

    and_ii _3185_ (
        .a(new_Jinkela_wire_3710),
        .b(new_Jinkela_wire_5141),
        .c(_0451_)
    );

    and_bb _3186_ (
        .a(new_Jinkela_wire_599),
        .b(new_Jinkela_wire_299),
        .c(_0452_)
    );

    and_bb _3187_ (
        .a(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_55),
        .c(_0453_)
    );

    and_ii _3188_ (
        .a(new_Jinkela_wire_12523),
        .b(new_Jinkela_wire_5811),
        .c(_0454_)
    );

    and_ii _3189_ (
        .a(new_Jinkela_wire_8582),
        .b(new_Jinkela_wire_3699),
        .c(_0455_)
    );

    and_bb _3190_ (
        .a(new_Jinkela_wire_8583),
        .b(new_Jinkela_wire_3700),
        .c(_0456_)
    );

    or_bb _3191_ (
        .a(new_Jinkela_wire_14694),
        .b(new_Jinkela_wire_1797),
        .c(_0457_)
    );

    and_ii _3192_ (
        .a(new_Jinkela_wire_11391),
        .b(new_Jinkela_wire_11384),
        .c(_0458_)
    );

    and_bb _3193_ (
        .a(new_Jinkela_wire_11392),
        .b(new_Jinkela_wire_11385),
        .c(_0460_)
    );

    or_bb _3194_ (
        .a(new_Jinkela_wire_7970),
        .b(new_Jinkela_wire_20357),
        .c(_0461_)
    );

    and_ii _3195_ (
        .a(new_Jinkela_wire_14083),
        .b(new_Jinkela_wire_10064),
        .c(_0462_)
    );

    and_bb _3196_ (
        .a(new_Jinkela_wire_14084),
        .b(new_Jinkela_wire_10065),
        .c(_0463_)
    );

    or_bb _3197_ (
        .a(new_Jinkela_wire_845),
        .b(new_Jinkela_wire_17317),
        .c(_0464_)
    );

    and_ii _3198_ (
        .a(new_Jinkela_wire_19349),
        .b(new_Jinkela_wire_9345),
        .c(_0465_)
    );

    and_bb _3199_ (
        .a(new_Jinkela_wire_19350),
        .b(new_Jinkela_wire_9346),
        .c(_0466_)
    );

    or_bb _3200_ (
        .a(new_Jinkela_wire_5160),
        .b(new_Jinkela_wire_14687),
        .c(_0467_)
    );

    and_ii _3201_ (
        .a(new_Jinkela_wire_12727),
        .b(new_Jinkela_wire_14096),
        .c(_0468_)
    );

    and_bb _3202_ (
        .a(new_Jinkela_wire_12728),
        .b(new_Jinkela_wire_14097),
        .c(_0469_)
    );

    or_bb _3203_ (
        .a(new_Jinkela_wire_16332),
        .b(new_Jinkela_wire_11344),
        .c(_0471_)
    );

    and_ii _3204_ (
        .a(new_Jinkela_wire_6757),
        .b(new_Jinkela_wire_3877),
        .c(_0472_)
    );

    and_bb _3205_ (
        .a(new_Jinkela_wire_6758),
        .b(new_Jinkela_wire_3878),
        .c(_0473_)
    );

    or_bb _3206_ (
        .a(new_Jinkela_wire_10275),
        .b(new_Jinkela_wire_3258),
        .c(_0474_)
    );

    and_ii _3207_ (
        .a(new_Jinkela_wire_19110),
        .b(new_Jinkela_wire_13459),
        .c(_0475_)
    );

    and_bb _3208_ (
        .a(new_Jinkela_wire_19111),
        .b(new_Jinkela_wire_13460),
        .c(_0476_)
    );

    or_bb _3209_ (
        .a(new_Jinkela_wire_19790),
        .b(new_Jinkela_wire_20962),
        .c(_0477_)
    );

    and_ii _3210_ (
        .a(new_Jinkela_wire_14194),
        .b(new_Jinkela_wire_16506),
        .c(_0478_)
    );

    and_bb _3211_ (
        .a(new_Jinkela_wire_14195),
        .b(new_Jinkela_wire_16507),
        .c(_0479_)
    );

    or_bb _3212_ (
        .a(new_Jinkela_wire_19346),
        .b(new_Jinkela_wire_20269),
        .c(_0480_)
    );

    and_ii _3213_ (
        .a(new_Jinkela_wire_13308),
        .b(new_Jinkela_wire_1896),
        .c(_0482_)
    );

    bfr new_Jinkela_buffer_9234 (
        .din(new_Jinkela_wire_11257),
        .dout(new_Jinkela_wire_11258)
    );

    bfr new_Jinkela_buffer_9172 (
        .din(new_Jinkela_wire_11191),
        .dout(new_Jinkela_wire_11192)
    );

    bfr new_Jinkela_buffer_9328 (
        .din(new_Jinkela_wire_11357),
        .dout(new_Jinkela_wire_11358)
    );

    bfr new_Jinkela_buffer_9173 (
        .din(new_Jinkela_wire_11192),
        .dout(new_Jinkela_wire_11193)
    );

    bfr new_Jinkela_buffer_9235 (
        .din(new_Jinkela_wire_11258),
        .dout(new_Jinkela_wire_11259)
    );

    bfr new_Jinkela_buffer_9174 (
        .din(new_Jinkela_wire_11193),
        .dout(new_Jinkela_wire_11194)
    );

    spl2 new_Jinkela_splitter_871 (
        .a(_1777_),
        .b(new_Jinkela_wire_11401),
        .c(new_Jinkela_wire_11402)
    );

    bfr new_Jinkela_buffer_9175 (
        .din(new_Jinkela_wire_11194),
        .dout(new_Jinkela_wire_11195)
    );

    bfr new_Jinkela_buffer_9236 (
        .din(new_Jinkela_wire_11259),
        .dout(new_Jinkela_wire_11260)
    );

    bfr new_Jinkela_buffer_9176 (
        .din(new_Jinkela_wire_11195),
        .dout(new_Jinkela_wire_11196)
    );

    bfr new_Jinkela_buffer_9329 (
        .din(new_Jinkela_wire_11358),
        .dout(new_Jinkela_wire_11359)
    );

    bfr new_Jinkela_buffer_9177 (
        .din(new_Jinkela_wire_11196),
        .dout(new_Jinkela_wire_11197)
    );

    bfr new_Jinkela_buffer_9237 (
        .din(new_Jinkela_wire_11260),
        .dout(new_Jinkela_wire_11261)
    );

    bfr new_Jinkela_buffer_9178 (
        .din(new_Jinkela_wire_11197),
        .dout(new_Jinkela_wire_11198)
    );

    bfr new_Jinkela_buffer_9357 (
        .din(_0009_),
        .dout(new_Jinkela_wire_11403)
    );

    bfr new_Jinkela_buffer_9358 (
        .din(_1333_),
        .dout(new_Jinkela_wire_11406)
    );

    bfr new_Jinkela_buffer_9179 (
        .din(new_Jinkela_wire_11198),
        .dout(new_Jinkela_wire_11199)
    );

    bfr new_Jinkela_buffer_9238 (
        .din(new_Jinkela_wire_11261),
        .dout(new_Jinkela_wire_11262)
    );

    bfr new_Jinkela_buffer_9180 (
        .din(new_Jinkela_wire_11199),
        .dout(new_Jinkela_wire_11200)
    );

    bfr new_Jinkela_buffer_9330 (
        .din(new_Jinkela_wire_11359),
        .dout(new_Jinkela_wire_11360)
    );

    bfr new_Jinkela_buffer_9181 (
        .din(new_Jinkela_wire_11200),
        .dout(new_Jinkela_wire_11201)
    );

    bfr new_Jinkela_buffer_9239 (
        .din(new_Jinkela_wire_11262),
        .dout(new_Jinkela_wire_11263)
    );

    bfr new_Jinkela_buffer_9182 (
        .din(new_Jinkela_wire_11201),
        .dout(new_Jinkela_wire_11202)
    );

    bfr new_Jinkela_buffer_9183 (
        .din(new_Jinkela_wire_11202),
        .dout(new_Jinkela_wire_11203)
    );

    bfr new_Jinkela_buffer_9240 (
        .din(new_Jinkela_wire_11263),
        .dout(new_Jinkela_wire_11264)
    );

    bfr new_Jinkela_buffer_9184 (
        .din(new_Jinkela_wire_11203),
        .dout(new_Jinkela_wire_11204)
    );

    bfr new_Jinkela_buffer_9331 (
        .din(new_Jinkela_wire_11360),
        .dout(new_Jinkela_wire_11361)
    );

    bfr new_Jinkela_buffer_9185 (
        .din(new_Jinkela_wire_11204),
        .dout(new_Jinkela_wire_11205)
    );

    bfr new_Jinkela_buffer_9241 (
        .din(new_Jinkela_wire_11264),
        .dout(new_Jinkela_wire_11265)
    );

    bfr new_Jinkela_buffer_9186 (
        .din(new_Jinkela_wire_11205),
        .dout(new_Jinkela_wire_11206)
    );

    spl2 new_Jinkela_splitter_872 (
        .a(_0284_),
        .b(new_Jinkela_wire_11404),
        .c(new_Jinkela_wire_11405)
    );

    bfr new_Jinkela_buffer_9187 (
        .din(new_Jinkela_wire_11206),
        .dout(new_Jinkela_wire_11207)
    );

    bfr new_Jinkela_buffer_9242 (
        .din(new_Jinkela_wire_11265),
        .dout(new_Jinkela_wire_11266)
    );

    bfr new_Jinkela_buffer_9188 (
        .din(new_Jinkela_wire_11207),
        .dout(new_Jinkela_wire_11208)
    );

    bfr new_Jinkela_buffer_9332 (
        .din(new_Jinkela_wire_11361),
        .dout(new_Jinkela_wire_11362)
    );

    bfr new_Jinkela_buffer_9189 (
        .din(new_Jinkela_wire_11208),
        .dout(new_Jinkela_wire_11209)
    );

    bfr new_Jinkela_buffer_9243 (
        .din(new_Jinkela_wire_11266),
        .dout(new_Jinkela_wire_11267)
    );

    bfr new_Jinkela_buffer_9190 (
        .din(new_Jinkela_wire_11209),
        .dout(new_Jinkela_wire_11210)
    );

    spl2 new_Jinkela_splitter_873 (
        .a(_1111_),
        .b(new_Jinkela_wire_11407),
        .c(new_Jinkela_wire_11408)
    );

    bfr new_Jinkela_buffer_9191 (
        .din(new_Jinkela_wire_11210),
        .dout(new_Jinkela_wire_11211)
    );

    bfr new_Jinkela_buffer_9244 (
        .din(new_Jinkela_wire_11267),
        .dout(new_Jinkela_wire_11268)
    );

    bfr new_Jinkela_buffer_9192 (
        .din(new_Jinkela_wire_11211),
        .dout(new_Jinkela_wire_11212)
    );

    bfr new_Jinkela_buffer_5744 (
        .din(new_Jinkela_wire_7333),
        .dout(new_Jinkela_wire_7334)
    );

    bfr new_Jinkela_buffer_5698 (
        .din(new_Jinkela_wire_7251),
        .dout(new_Jinkela_wire_7252)
    );

    bfr new_Jinkela_buffer_5902 (
        .din(_1520_),
        .dout(new_Jinkela_wire_7504)
    );

    bfr new_Jinkela_buffer_5699 (
        .din(new_Jinkela_wire_7252),
        .dout(new_Jinkela_wire_7253)
    );

    bfr new_Jinkela_buffer_5745 (
        .din(new_Jinkela_wire_7334),
        .dout(new_Jinkela_wire_7335)
    );

    bfr new_Jinkela_buffer_5700 (
        .din(new_Jinkela_wire_7253),
        .dout(new_Jinkela_wire_7254)
    );

    bfr new_Jinkela_buffer_5851 (
        .din(new_Jinkela_wire_7448),
        .dout(new_Jinkela_wire_7449)
    );

    bfr new_Jinkela_buffer_5701 (
        .din(new_Jinkela_wire_7254),
        .dout(new_Jinkela_wire_7255)
    );

    bfr new_Jinkela_buffer_5746 (
        .din(new_Jinkela_wire_7335),
        .dout(new_Jinkela_wire_7336)
    );

    bfr new_Jinkela_buffer_5702 (
        .din(new_Jinkela_wire_7255),
        .dout(new_Jinkela_wire_7256)
    );

    bfr new_Jinkela_buffer_5855 (
        .din(new_Jinkela_wire_7452),
        .dout(new_Jinkela_wire_7453)
    );

    bfr new_Jinkela_buffer_5703 (
        .din(new_Jinkela_wire_7256),
        .dout(new_Jinkela_wire_7257)
    );

    bfr new_Jinkela_buffer_5747 (
        .din(new_Jinkela_wire_7336),
        .dout(new_Jinkela_wire_7337)
    );

    bfr new_Jinkela_buffer_5704 (
        .din(new_Jinkela_wire_7257),
        .dout(new_Jinkela_wire_7258)
    );

    bfr new_Jinkela_buffer_5852 (
        .din(new_Jinkela_wire_7449),
        .dout(new_Jinkela_wire_7450)
    );

    spl2 new_Jinkela_splitter_626 (
        .a(new_Jinkela_wire_7258),
        .b(new_Jinkela_wire_7259),
        .c(new_Jinkela_wire_7260)
    );

    spl2 new_Jinkela_splitter_650 (
        .a(_1745_),
        .b(new_Jinkela_wire_7506),
        .c(new_Jinkela_wire_7507)
    );

    bfr new_Jinkela_buffer_5748 (
        .din(new_Jinkela_wire_7337),
        .dout(new_Jinkela_wire_7338)
    );

    bfr new_Jinkela_buffer_5749 (
        .din(new_Jinkela_wire_7338),
        .dout(new_Jinkela_wire_7339)
    );

    bfr new_Jinkela_buffer_5856 (
        .din(new_Jinkela_wire_7453),
        .dout(new_Jinkela_wire_7454)
    );

    bfr new_Jinkela_buffer_5750 (
        .din(new_Jinkela_wire_7339),
        .dout(new_Jinkela_wire_7340)
    );

    bfr new_Jinkela_buffer_5903 (
        .din(_1670_),
        .dout(new_Jinkela_wire_7505)
    );

    bfr new_Jinkela_buffer_5751 (
        .din(new_Jinkela_wire_7340),
        .dout(new_Jinkela_wire_7341)
    );

    bfr new_Jinkela_buffer_5857 (
        .din(new_Jinkela_wire_7454),
        .dout(new_Jinkela_wire_7455)
    );

    bfr new_Jinkela_buffer_5752 (
        .din(new_Jinkela_wire_7341),
        .dout(new_Jinkela_wire_7342)
    );

    spl2 new_Jinkela_splitter_651 (
        .a(_1805_),
        .b(new_Jinkela_wire_7512),
        .c(new_Jinkela_wire_7513)
    );

    bfr new_Jinkela_buffer_5904 (
        .din(new_Jinkela_wire_7507),
        .dout(new_Jinkela_wire_7508)
    );

    bfr new_Jinkela_buffer_5753 (
        .din(new_Jinkela_wire_7342),
        .dout(new_Jinkela_wire_7343)
    );

    bfr new_Jinkela_buffer_5858 (
        .din(new_Jinkela_wire_7455),
        .dout(new_Jinkela_wire_7456)
    );

    bfr new_Jinkela_buffer_5754 (
        .din(new_Jinkela_wire_7343),
        .dout(new_Jinkela_wire_7344)
    );

    bfr new_Jinkela_buffer_5755 (
        .din(new_Jinkela_wire_7344),
        .dout(new_Jinkela_wire_7345)
    );

    bfr new_Jinkela_buffer_5859 (
        .din(new_Jinkela_wire_7456),
        .dout(new_Jinkela_wire_7457)
    );

    bfr new_Jinkela_buffer_5756 (
        .din(new_Jinkela_wire_7345),
        .dout(new_Jinkela_wire_7346)
    );

    spl2 new_Jinkela_splitter_652 (
        .a(_0768_),
        .b(new_Jinkela_wire_7514),
        .c(new_Jinkela_wire_7515)
    );

    bfr new_Jinkela_buffer_5757 (
        .din(new_Jinkela_wire_7346),
        .dout(new_Jinkela_wire_7347)
    );

    bfr new_Jinkela_buffer_5860 (
        .din(new_Jinkela_wire_7457),
        .dout(new_Jinkela_wire_7458)
    );

    bfr new_Jinkela_buffer_5758 (
        .din(new_Jinkela_wire_7347),
        .dout(new_Jinkela_wire_7348)
    );

    bfr new_Jinkela_buffer_5908 (
        .din(_1815_),
        .dout(new_Jinkela_wire_7516)
    );

    bfr new_Jinkela_buffer_5759 (
        .din(new_Jinkela_wire_7348),
        .dout(new_Jinkela_wire_7349)
    );

    bfr new_Jinkela_buffer_5861 (
        .din(new_Jinkela_wire_7458),
        .dout(new_Jinkela_wire_7459)
    );

    bfr new_Jinkela_buffer_5760 (
        .din(new_Jinkela_wire_7349),
        .dout(new_Jinkela_wire_7350)
    );

    bfr new_Jinkela_buffer_5905 (
        .din(new_Jinkela_wire_7508),
        .dout(new_Jinkela_wire_7509)
    );

    bfr new_Jinkela_buffer_2114 (
        .din(new_Jinkela_wire_3055),
        .dout(new_Jinkela_wire_3056)
    );

    bfr new_Jinkela_buffer_2215 (
        .din(new_Jinkela_wire_3164),
        .dout(new_Jinkela_wire_3165)
    );

    bfr new_Jinkela_buffer_2115 (
        .din(new_Jinkela_wire_3056),
        .dout(new_Jinkela_wire_3057)
    );

    bfr new_Jinkela_buffer_2116 (
        .din(new_Jinkela_wire_3057),
        .dout(new_Jinkela_wire_3058)
    );

    spl2 new_Jinkela_splitter_342 (
        .a(_1109_),
        .b(new_Jinkela_wire_3271),
        .c(new_Jinkela_wire_3272)
    );

    bfr new_Jinkela_buffer_2216 (
        .din(new_Jinkela_wire_3165),
        .dout(new_Jinkela_wire_3166)
    );

    bfr new_Jinkela_buffer_2117 (
        .din(new_Jinkela_wire_3058),
        .dout(new_Jinkela_wire_3059)
    );

    bfr new_Jinkela_buffer_2248 (
        .din(new_Jinkela_wire_3213),
        .dout(new_Jinkela_wire_3214)
    );

    bfr new_Jinkela_buffer_2118 (
        .din(new_Jinkela_wire_3059),
        .dout(new_Jinkela_wire_3060)
    );

    bfr new_Jinkela_buffer_2217 (
        .din(new_Jinkela_wire_3166),
        .dout(new_Jinkela_wire_3167)
    );

    bfr new_Jinkela_buffer_2119 (
        .din(new_Jinkela_wire_3060),
        .dout(new_Jinkela_wire_3061)
    );

    bfr new_Jinkela_buffer_2280 (
        .din(new_Jinkela_wire_3261),
        .dout(new_Jinkela_wire_3262)
    );

    bfr new_Jinkela_buffer_2120 (
        .din(new_Jinkela_wire_3061),
        .dout(new_Jinkela_wire_3062)
    );

    bfr new_Jinkela_buffer_2218 (
        .din(new_Jinkela_wire_3167),
        .dout(new_Jinkela_wire_3168)
    );

    bfr new_Jinkela_buffer_2121 (
        .din(new_Jinkela_wire_3062),
        .dout(new_Jinkela_wire_3063)
    );

    bfr new_Jinkela_buffer_2249 (
        .din(new_Jinkela_wire_3214),
        .dout(new_Jinkela_wire_3215)
    );

    bfr new_Jinkela_buffer_2122 (
        .din(new_Jinkela_wire_3063),
        .dout(new_Jinkela_wire_3064)
    );

    bfr new_Jinkela_buffer_2219 (
        .din(new_Jinkela_wire_3168),
        .dout(new_Jinkela_wire_3169)
    );

    bfr new_Jinkela_buffer_2123 (
        .din(new_Jinkela_wire_3064),
        .dout(new_Jinkela_wire_3065)
    );

    bfr new_Jinkela_buffer_2124 (
        .din(new_Jinkela_wire_3065),
        .dout(new_Jinkela_wire_3066)
    );

    bfr new_Jinkela_buffer_2220 (
        .din(new_Jinkela_wire_3169),
        .dout(new_Jinkela_wire_3170)
    );

    bfr new_Jinkela_buffer_2125 (
        .din(new_Jinkela_wire_3066),
        .dout(new_Jinkela_wire_3067)
    );

    bfr new_Jinkela_buffer_2250 (
        .din(new_Jinkela_wire_3215),
        .dout(new_Jinkela_wire_3216)
    );

    bfr new_Jinkela_buffer_2126 (
        .din(new_Jinkela_wire_3067),
        .dout(new_Jinkela_wire_3068)
    );

    bfr new_Jinkela_buffer_2221 (
        .din(new_Jinkela_wire_3170),
        .dout(new_Jinkela_wire_3171)
    );

    bfr new_Jinkela_buffer_2127 (
        .din(new_Jinkela_wire_3068),
        .dout(new_Jinkela_wire_3069)
    );

    bfr new_Jinkela_buffer_2281 (
        .din(new_Jinkela_wire_3262),
        .dout(new_Jinkela_wire_3263)
    );

    bfr new_Jinkela_buffer_2128 (
        .din(new_Jinkela_wire_3069),
        .dout(new_Jinkela_wire_3070)
    );

    bfr new_Jinkela_buffer_2222 (
        .din(new_Jinkela_wire_3171),
        .dout(new_Jinkela_wire_3172)
    );

    bfr new_Jinkela_buffer_2129 (
        .din(new_Jinkela_wire_3070),
        .dout(new_Jinkela_wire_3071)
    );

    bfr new_Jinkela_buffer_2251 (
        .din(new_Jinkela_wire_3216),
        .dout(new_Jinkela_wire_3217)
    );

    bfr new_Jinkela_buffer_2130 (
        .din(new_Jinkela_wire_3071),
        .dout(new_Jinkela_wire_3072)
    );

    bfr new_Jinkela_buffer_2223 (
        .din(new_Jinkela_wire_3172),
        .dout(new_Jinkela_wire_3173)
    );

    bfr new_Jinkela_buffer_2131 (
        .din(new_Jinkela_wire_3072),
        .dout(new_Jinkela_wire_3073)
    );

    spl2 new_Jinkela_splitter_344 (
        .a(_1228_),
        .b(new_Jinkela_wire_3361),
        .c(new_Jinkela_wire_3362)
    );

    bfr new_Jinkela_buffer_2132 (
        .din(new_Jinkela_wire_3073),
        .dout(new_Jinkela_wire_3074)
    );

    bfr new_Jinkela_buffer_2285 (
        .din(_0835_),
        .dout(new_Jinkela_wire_3273)
    );

    bfr new_Jinkela_buffer_2224 (
        .din(new_Jinkela_wire_3173),
        .dout(new_Jinkela_wire_3174)
    );

    bfr new_Jinkela_buffer_2133 (
        .din(new_Jinkela_wire_3074),
        .dout(new_Jinkela_wire_3075)
    );

    bfr new_Jinkela_buffer_2252 (
        .din(new_Jinkela_wire_3217),
        .dout(new_Jinkela_wire_3218)
    );

    bfr new_Jinkela_buffer_2134 (
        .din(new_Jinkela_wire_3075),
        .dout(new_Jinkela_wire_3076)
    );

    bfr new_Jinkela_buffer_2225 (
        .din(new_Jinkela_wire_3174),
        .dout(new_Jinkela_wire_3175)
    );

    bfr new_Jinkela_buffer_2135 (
        .din(new_Jinkela_wire_3076),
        .dout(new_Jinkela_wire_3077)
    );

    bfr new_Jinkela_buffer_16087 (
        .din(new_Jinkela_wire_19211),
        .dout(new_Jinkela_wire_19212)
    );

    bfr new_Jinkela_buffer_16158 (
        .din(new_Jinkela_wire_19294),
        .dout(new_Jinkela_wire_19295)
    );

    bfr new_Jinkela_buffer_16088 (
        .din(new_Jinkela_wire_19212),
        .dout(new_Jinkela_wire_19213)
    );

    bfr new_Jinkela_buffer_16089 (
        .din(new_Jinkela_wire_19213),
        .dout(new_Jinkela_wire_19214)
    );

    bfr new_Jinkela_buffer_16161 (
        .din(new_Jinkela_wire_19299),
        .dout(new_Jinkela_wire_19300)
    );

    bfr new_Jinkela_buffer_16090 (
        .din(new_Jinkela_wire_19214),
        .dout(new_Jinkela_wire_19215)
    );

    spl2 new_Jinkela_splitter_1421 (
        .a(_1070_),
        .b(new_Jinkela_wire_19326),
        .c(new_Jinkela_wire_19327)
    );

    bfr new_Jinkela_buffer_16091 (
        .din(new_Jinkela_wire_19215),
        .dout(new_Jinkela_wire_19216)
    );

    bfr new_Jinkela_buffer_16162 (
        .din(new_Jinkela_wire_19300),
        .dout(new_Jinkela_wire_19301)
    );

    bfr new_Jinkela_buffer_16092 (
        .din(new_Jinkela_wire_19216),
        .dout(new_Jinkela_wire_19217)
    );

    bfr new_Jinkela_buffer_16177 (
        .din(new_Jinkela_wire_19321),
        .dout(new_Jinkela_wire_19322)
    );

    spl2 new_Jinkela_splitter_1422 (
        .a(_0051_),
        .b(new_Jinkela_wire_19328),
        .c(new_Jinkela_wire_19329)
    );

    bfr new_Jinkela_buffer_16093 (
        .din(new_Jinkela_wire_19217),
        .dout(new_Jinkela_wire_19218)
    );

    bfr new_Jinkela_buffer_16163 (
        .din(new_Jinkela_wire_19301),
        .dout(new_Jinkela_wire_19302)
    );

    bfr new_Jinkela_buffer_16094 (
        .din(new_Jinkela_wire_19218),
        .dout(new_Jinkela_wire_19219)
    );

    bfr new_Jinkela_buffer_16095 (
        .din(new_Jinkela_wire_19219),
        .dout(new_Jinkela_wire_19220)
    );

    bfr new_Jinkela_buffer_16164 (
        .din(new_Jinkela_wire_19302),
        .dout(new_Jinkela_wire_19303)
    );

    bfr new_Jinkela_buffer_16096 (
        .din(new_Jinkela_wire_19220),
        .dout(new_Jinkela_wire_19221)
    );

    bfr new_Jinkela_buffer_16178 (
        .din(new_Jinkela_wire_19322),
        .dout(new_Jinkela_wire_19323)
    );

    bfr new_Jinkela_buffer_16097 (
        .din(new_Jinkela_wire_19221),
        .dout(new_Jinkela_wire_19222)
    );

    bfr new_Jinkela_buffer_16165 (
        .din(new_Jinkela_wire_19303),
        .dout(new_Jinkela_wire_19304)
    );

    bfr new_Jinkela_buffer_16098 (
        .din(new_Jinkela_wire_19222),
        .dout(new_Jinkela_wire_19223)
    );

    bfr new_Jinkela_buffer_16185 (
        .din(_0016_),
        .dout(new_Jinkela_wire_19334)
    );

    bfr new_Jinkela_buffer_16099 (
        .din(new_Jinkela_wire_19223),
        .dout(new_Jinkela_wire_19224)
    );

    bfr new_Jinkela_buffer_16166 (
        .din(new_Jinkela_wire_19304),
        .dout(new_Jinkela_wire_19305)
    );

    bfr new_Jinkela_buffer_16100 (
        .din(new_Jinkela_wire_19224),
        .dout(new_Jinkela_wire_19225)
    );

    bfr new_Jinkela_buffer_16179 (
        .din(new_Jinkela_wire_19323),
        .dout(new_Jinkela_wire_19324)
    );

    bfr new_Jinkela_buffer_16101 (
        .din(new_Jinkela_wire_19225),
        .dout(new_Jinkela_wire_19226)
    );

    bfr new_Jinkela_buffer_16167 (
        .din(new_Jinkela_wire_19305),
        .dout(new_Jinkela_wire_19306)
    );

    bfr new_Jinkela_buffer_16102 (
        .din(new_Jinkela_wire_19226),
        .dout(new_Jinkela_wire_19227)
    );

    bfr new_Jinkela_buffer_16181 (
        .din(new_Jinkela_wire_19329),
        .dout(new_Jinkela_wire_19330)
    );

    spl2 new_Jinkela_splitter_1423 (
        .a(_0739_),
        .b(new_Jinkela_wire_19335),
        .c(new_Jinkela_wire_19336)
    );

    bfr new_Jinkela_buffer_16103 (
        .din(new_Jinkela_wire_19227),
        .dout(new_Jinkela_wire_19228)
    );

    bfr new_Jinkela_buffer_16168 (
        .din(new_Jinkela_wire_19306),
        .dout(new_Jinkela_wire_19307)
    );

    bfr new_Jinkela_buffer_16104 (
        .din(new_Jinkela_wire_19228),
        .dout(new_Jinkela_wire_19229)
    );

    bfr new_Jinkela_buffer_16180 (
        .din(new_Jinkela_wire_19324),
        .dout(new_Jinkela_wire_19325)
    );

    bfr new_Jinkela_buffer_16105 (
        .din(new_Jinkela_wire_19229),
        .dout(new_Jinkela_wire_19230)
    );

    bfr new_Jinkela_buffer_16169 (
        .din(new_Jinkela_wire_19307),
        .dout(new_Jinkela_wire_19308)
    );

    bfr new_Jinkela_buffer_16106 (
        .din(new_Jinkela_wire_19230),
        .dout(new_Jinkela_wire_19231)
    );

    bfr new_Jinkela_buffer_16190 (
        .din(_1104_),
        .dout(new_Jinkela_wire_19341)
    );

    bfr new_Jinkela_buffer_16107 (
        .din(new_Jinkela_wire_19231),
        .dout(new_Jinkela_wire_19232)
    );

    bfr new_Jinkela_buffer_16170 (
        .din(new_Jinkela_wire_19308),
        .dout(new_Jinkela_wire_19309)
    );

    and_bb _2497_ (
        .a(new_Jinkela_wire_13200),
        .b(new_Jinkela_wire_12904),
        .c(_1540_)
    );

    or_bb _2498_ (
        .a(new_Jinkela_wire_16333),
        .b(new_Jinkela_wire_14017),
        .c(_1541_)
    );

    or_bb _2499_ (
        .a(new_Jinkela_wire_8292),
        .b(new_Jinkela_wire_17424),
        .c(_1542_)
    );

    or_ii _2500_ (
        .a(new_Jinkela_wire_8293),
        .b(new_Jinkela_wire_17425),
        .c(_1543_)
    );

    or_ii _2501_ (
        .a(new_Jinkela_wire_15733),
        .b(new_Jinkela_wire_3429),
        .c(_1544_)
    );

    and_ii _2502_ (
        .a(new_Jinkela_wire_830),
        .b(new_Jinkela_wire_6615),
        .c(_1545_)
    );

    and_bb _2503_ (
        .a(new_Jinkela_wire_831),
        .b(new_Jinkela_wire_6616),
        .c(_1546_)
    );

    or_bb _2504_ (
        .a(new_Jinkela_wire_14258),
        .b(new_Jinkela_wire_2419),
        .c(_1547_)
    );

    or_bb _2505_ (
        .a(new_Jinkela_wire_5740),
        .b(new_Jinkela_wire_7710),
        .c(_1548_)
    );

    or_ii _2506_ (
        .a(new_Jinkela_wire_5741),
        .b(new_Jinkela_wire_7711),
        .c(_1549_)
    );

    or_ii _2507_ (
        .a(new_Jinkela_wire_2421),
        .b(new_Jinkela_wire_16516),
        .c(_1550_)
    );

    and_ii _2508_ (
        .a(new_Jinkela_wire_13970),
        .b(new_Jinkela_wire_12613),
        .c(_1551_)
    );

    and_bb _2509_ (
        .a(new_Jinkela_wire_13971),
        .b(new_Jinkela_wire_12614),
        .c(_1552_)
    );

    or_bb _2510_ (
        .a(new_Jinkela_wire_7588),
        .b(new_Jinkela_wire_9185),
        .c(_1553_)
    );

    or_bb _2511_ (
        .a(new_Jinkela_wire_9864),
        .b(new_Jinkela_wire_13205),
        .c(_1554_)
    );

    and_bb _2512_ (
        .a(new_Jinkela_wire_9865),
        .b(new_Jinkela_wire_13206),
        .c(_1555_)
    );

    or_bi _2513_ (
        .a(new_Jinkela_wire_7728),
        .b(new_Jinkela_wire_13342),
        .c(_1557_)
    );

    and_ii _2514_ (
        .a(new_Jinkela_wire_2315),
        .b(new_Jinkela_wire_6957),
        .c(_1558_)
    );

    and_bb _2515_ (
        .a(new_Jinkela_wire_2316),
        .b(new_Jinkela_wire_6958),
        .c(_1559_)
    );

    or_bb _2516_ (
        .a(new_Jinkela_wire_18108),
        .b(new_Jinkela_wire_20903),
        .c(new_net_3962)
    );

    and_bb _2517_ (
        .a(new_Jinkela_wire_335),
        .b(new_Jinkela_wire_512),
        .c(_1560_)
    );

    and_bi _2518_ (
        .a(new_Jinkela_wire_13347),
        .b(new_Jinkela_wire_20904),
        .c(_1561_)
    );

    and_bb _2519_ (
        .a(new_Jinkela_wire_94),
        .b(new_Jinkela_wire_149),
        .c(_1562_)
    );

    and_bi _2520_ (
        .a(new_Jinkela_wire_16521),
        .b(new_Jinkela_wire_9186),
        .c(_1563_)
    );

    and_bb _2521_ (
        .a(new_Jinkela_wire_214),
        .b(new_Jinkela_wire_564),
        .c(_1564_)
    );

    and_bi _2522_ (
        .a(new_Jinkela_wire_3434),
        .b(new_Jinkela_wire_2420),
        .c(_1565_)
    );

    and_bb _2523_ (
        .a(new_Jinkela_wire_269),
        .b(new_Jinkela_wire_591),
        .c(_1567_)
    );

    and_bi _2524_ (
        .a(new_Jinkela_wire_13690),
        .b(new_Jinkela_wire_14018),
        .c(_1568_)
    );

    and_bb _2525_ (
        .a(new_Jinkela_wire_84),
        .b(new_Jinkela_wire_108),
        .c(_1569_)
    );

    and_bi _2526_ (
        .a(new_Jinkela_wire_8872),
        .b(new_Jinkela_wire_4689),
        .c(_1570_)
    );

    and_bb _2527_ (
        .a(new_Jinkela_wire_485),
        .b(new_Jinkela_wire_10),
        .c(_1571_)
    );

    and_bi _2528_ (
        .a(new_Jinkela_wire_17004),
        .b(new_Jinkela_wire_9522),
        .c(_1572_)
    );

    and_bb _2529_ (
        .a(new_Jinkela_wire_355),
        .b(new_Jinkela_wire_459),
        .c(_1573_)
    );

    and_bi _2530_ (
        .a(new_Jinkela_wire_4079),
        .b(new_Jinkela_wire_19297),
        .c(_1574_)
    );

    and_bb _2531_ (
        .a(new_Jinkela_wire_696),
        .b(new_Jinkela_wire_257),
        .c(_1575_)
    );

    and_bi _2532_ (
        .a(new_Jinkela_wire_1582),
        .b(new_Jinkela_wire_13215),
        .c(_1576_)
    );

    and_bb _2533_ (
        .a(new_Jinkela_wire_293),
        .b(new_Jinkela_wire_494),
        .c(_1578_)
    );

    and_bi _2534_ (
        .a(new_Jinkela_wire_13995),
        .b(new_Jinkela_wire_6736),
        .c(_1579_)
    );

    and_bb _2535_ (
        .a(new_Jinkela_wire_30),
        .b(new_Jinkela_wire_52),
        .c(_1580_)
    );

    and_bi _2536_ (
        .a(new_Jinkela_wire_11233),
        .b(new_Jinkela_wire_6364),
        .c(_1581_)
    );

    and_bb _2537_ (
        .a(new_Jinkela_wire_186),
        .b(new_Jinkela_wire_642),
        .c(_1582_)
    );

    and_bi _2538_ (
        .a(new_Jinkela_wire_18796),
        .b(new_Jinkela_wire_17980),
        .c(_1583_)
    );

    bfr new_Jinkela_buffer_15317 (
        .din(new_Jinkela_wire_18257),
        .dout(new_Jinkela_wire_18258)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_2112),
        .dout(new_Jinkela_wire_2113)
    );

    bfr new_Jinkela_buffer_15255 (
        .din(new_Jinkela_wire_18189),
        .dout(new_Jinkela_wire_18190)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_2186),
        .dout(new_Jinkela_wire_2187)
    );

    bfr new_Jinkela_buffer_15358 (
        .din(new_Jinkela_wire_18312),
        .dout(new_Jinkela_wire_18313)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(new_Jinkela_wire_2113),
        .dout(new_Jinkela_wire_2114)
    );

    bfr new_Jinkela_buffer_15256 (
        .din(new_Jinkela_wire_18190),
        .dout(new_Jinkela_wire_18191)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(new_Jinkela_wire_2328),
        .dout(new_Jinkela_wire_2329)
    );

    bfr new_Jinkela_buffer_15318 (
        .din(new_Jinkela_wire_18258),
        .dout(new_Jinkela_wire_18259)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(new_Jinkela_wire_2114),
        .b(new_Jinkela_wire_2115),
        .c(new_Jinkela_wire_2116)
    );

    bfr new_Jinkela_buffer_15257 (
        .din(new_Jinkela_wire_18191),
        .dout(new_Jinkela_wire_18192)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_2275),
        .dout(new_Jinkela_wire_2276)
    );

    bfr new_Jinkela_buffer_15355 (
        .din(new_Jinkela_wire_18305),
        .dout(new_Jinkela_wire_18306)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_2187),
        .dout(new_Jinkela_wire_2188)
    );

    bfr new_Jinkela_buffer_15258 (
        .din(new_Jinkela_wire_18192),
        .dout(new_Jinkela_wire_18193)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_2188),
        .dout(new_Jinkela_wire_2189)
    );

    bfr new_Jinkela_buffer_15319 (
        .din(new_Jinkela_wire_18259),
        .dout(new_Jinkela_wire_18260)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_Jinkela_wire_2332),
        .dout(new_Jinkela_wire_2333)
    );

    bfr new_Jinkela_buffer_15259 (
        .din(new_Jinkela_wire_18193),
        .dout(new_Jinkela_wire_18194)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_2189),
        .dout(new_Jinkela_wire_2190)
    );

    spl2 new_Jinkela_splitter_1329 (
        .a(_1320_),
        .b(new_Jinkela_wire_18381),
        .c(new_Jinkela_wire_18382)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(new_Jinkela_wire_2276),
        .dout(new_Jinkela_wire_2277)
    );

    bfr new_Jinkela_buffer_15260 (
        .din(new_Jinkela_wire_18194),
        .dout(new_Jinkela_wire_18195)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_2190),
        .dout(new_Jinkela_wire_2191)
    );

    bfr new_Jinkela_buffer_15320 (
        .din(new_Jinkela_wire_18260),
        .dout(new_Jinkela_wire_18261)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_2329),
        .dout(new_Jinkela_wire_2330)
    );

    bfr new_Jinkela_buffer_15261 (
        .din(new_Jinkela_wire_18195),
        .dout(new_Jinkela_wire_18196)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_Jinkela_wire_2191),
        .dout(new_Jinkela_wire_2192)
    );

    spl2 new_Jinkela_splitter_1324 (
        .a(new_Jinkela_wire_18306),
        .b(new_Jinkela_wire_18307),
        .c(new_Jinkela_wire_18308)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(new_Jinkela_wire_2277),
        .dout(new_Jinkela_wire_2278)
    );

    bfr new_Jinkela_buffer_15262 (
        .din(new_Jinkela_wire_18196),
        .dout(new_Jinkela_wire_18197)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_2192),
        .dout(new_Jinkela_wire_2193)
    );

    bfr new_Jinkela_buffer_15321 (
        .din(new_Jinkela_wire_18261),
        .dout(new_Jinkela_wire_18262)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(_0337_),
        .dout(new_Jinkela_wire_2345)
    );

    bfr new_Jinkela_buffer_15263 (
        .din(new_Jinkela_wire_18197),
        .dout(new_Jinkela_wire_18198)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_2193),
        .dout(new_Jinkela_wire_2194)
    );

    bfr new_Jinkela_buffer_15362 (
        .din(new_Jinkela_wire_18316),
        .dout(new_Jinkela_wire_18317)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_2278),
        .dout(new_Jinkela_wire_2279)
    );

    bfr new_Jinkela_buffer_15264 (
        .din(new_Jinkela_wire_18198),
        .dout(new_Jinkela_wire_18199)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_2194),
        .dout(new_Jinkela_wire_2195)
    );

    bfr new_Jinkela_buffer_15322 (
        .din(new_Jinkela_wire_18262),
        .dout(new_Jinkela_wire_18263)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_2330),
        .dout(new_Jinkela_wire_2331)
    );

    bfr new_Jinkela_buffer_15265 (
        .din(new_Jinkela_wire_18199),
        .dout(new_Jinkela_wire_18200)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_2195),
        .dout(new_Jinkela_wire_2196)
    );

    bfr new_Jinkela_buffer_15359 (
        .din(new_Jinkela_wire_18313),
        .dout(new_Jinkela_wire_18314)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_2279),
        .dout(new_Jinkela_wire_2280)
    );

    bfr new_Jinkela_buffer_15266 (
        .din(new_Jinkela_wire_18200),
        .dout(new_Jinkela_wire_18201)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(new_Jinkela_wire_2196),
        .dout(new_Jinkela_wire_2197)
    );

    bfr new_Jinkela_buffer_15323 (
        .din(new_Jinkela_wire_18263),
        .dout(new_Jinkela_wire_18264)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(new_Jinkela_wire_2333),
        .dout(new_Jinkela_wire_2334)
    );

    bfr new_Jinkela_buffer_15267 (
        .din(new_Jinkela_wire_18201),
        .dout(new_Jinkela_wire_18202)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(new_Jinkela_wire_2197),
        .dout(new_Jinkela_wire_2198)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_2280),
        .dout(new_Jinkela_wire_2281)
    );

    bfr new_Jinkela_buffer_15418 (
        .din(_1339_),
        .dout(new_Jinkela_wire_18379)
    );

    bfr new_Jinkela_buffer_15268 (
        .din(new_Jinkela_wire_18202),
        .dout(new_Jinkela_wire_18203)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(new_Jinkela_wire_2198),
        .dout(new_Jinkela_wire_2199)
    );

    bfr new_Jinkela_buffer_15324 (
        .din(new_Jinkela_wire_18264),
        .dout(new_Jinkela_wire_18265)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(_1549_),
        .dout(new_Jinkela_wire_2421)
    );

    bfr new_Jinkela_buffer_15269 (
        .din(new_Jinkela_wire_18203),
        .dout(new_Jinkela_wire_18204)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_2199),
        .dout(new_Jinkela_wire_2200)
    );

    bfr new_Jinkela_buffer_15363 (
        .din(new_Jinkela_wire_18317),
        .dout(new_Jinkela_wire_18318)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(new_Jinkela_wire_2281),
        .dout(new_Jinkela_wire_2282)
    );

    bfr new_Jinkela_buffer_15270 (
        .din(new_Jinkela_wire_18204),
        .dout(new_Jinkela_wire_18205)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_2200),
        .dout(new_Jinkela_wire_2201)
    );

    bfr new_Jinkela_buffer_15325 (
        .din(new_Jinkela_wire_18265),
        .dout(new_Jinkela_wire_18266)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_2334),
        .dout(new_Jinkela_wire_2335)
    );

    bfr new_Jinkela_buffer_15271 (
        .din(new_Jinkela_wire_18205),
        .dout(new_Jinkela_wire_18206)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(new_Jinkela_wire_2201),
        .dout(new_Jinkela_wire_2202)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(new_Jinkela_wire_2282),
        .dout(new_Jinkela_wire_2283)
    );

    bfr new_Jinkela_buffer_15419 (
        .din(_0264_),
        .dout(new_Jinkela_wire_18380)
    );

    bfr new_Jinkela_buffer_15272 (
        .din(new_Jinkela_wire_18206),
        .dout(new_Jinkela_wire_18207)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_2202),
        .dout(new_Jinkela_wire_2203)
    );

    bfr new_Jinkela_buffer_15326 (
        .din(new_Jinkela_wire_18266),
        .dout(new_Jinkela_wire_18267)
    );

    spl2 new_Jinkela_splitter_289 (
        .a(_1545_),
        .b(new_Jinkela_wire_2419),
        .c(new_Jinkela_wire_2420)
    );

    bfr new_Jinkela_buffer_15273 (
        .din(new_Jinkela_wire_18207),
        .dout(new_Jinkela_wire_18208)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_2203),
        .dout(new_Jinkela_wire_2204)
    );

    bfr new_Jinkela_buffer_15364 (
        .din(new_Jinkela_wire_18318),
        .dout(new_Jinkela_wire_18319)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(new_Jinkela_wire_2283),
        .dout(new_Jinkela_wire_2284)
    );

    bfr new_Jinkela_buffer_15274 (
        .din(new_Jinkela_wire_18208),
        .dout(new_Jinkela_wire_18209)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_2204),
        .dout(new_Jinkela_wire_2205)
    );

    bfr new_Jinkela_buffer_15327 (
        .din(new_Jinkela_wire_18267),
        .dout(new_Jinkela_wire_18268)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(new_Jinkela_wire_2335),
        .dout(new_Jinkela_wire_2336)
    );

    bfr new_Jinkela_buffer_15275 (
        .din(new_Jinkela_wire_18209),
        .dout(new_Jinkela_wire_18210)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_2205),
        .dout(new_Jinkela_wire_2206)
    );

    bfr new_Jinkela_buffer_4969 (
        .din(new_Jinkela_wire_6428),
        .dout(new_Jinkela_wire_6429)
    );

    bfr new_Jinkela_buffer_8360 (
        .din(new_Jinkela_wire_10301),
        .dout(new_Jinkela_wire_10302)
    );

    bfr new_Jinkela_buffer_4882 (
        .din(new_Jinkela_wire_6313),
        .dout(new_Jinkela_wire_6314)
    );

    bfr new_Jinkela_buffer_5061 (
        .din(_1456_),
        .dout(new_Jinkela_wire_6535)
    );

    bfr new_Jinkela_buffer_8361 (
        .din(new_Jinkela_wire_10302),
        .dout(new_Jinkela_wire_10303)
    );

    bfr new_Jinkela_buffer_4883 (
        .din(new_Jinkela_wire_6314),
        .dout(new_Jinkela_wire_6315)
    );

    bfr new_Jinkela_buffer_8460 (
        .din(new_Jinkela_wire_10409),
        .dout(new_Jinkela_wire_10410)
    );

    bfr new_Jinkela_buffer_8362 (
        .din(new_Jinkela_wire_10303),
        .dout(new_Jinkela_wire_10304)
    );

    bfr new_Jinkela_buffer_4884 (
        .din(new_Jinkela_wire_6315),
        .dout(new_Jinkela_wire_6316)
    );

    bfr new_Jinkela_buffer_8496 (
        .din(new_Jinkela_wire_10445),
        .dout(new_Jinkela_wire_10446)
    );

    bfr new_Jinkela_buffer_5052 (
        .din(_0731_),
        .dout(new_Jinkela_wire_6524)
    );

    bfr new_Jinkela_buffer_4970 (
        .din(new_Jinkela_wire_6429),
        .dout(new_Jinkela_wire_6430)
    );

    bfr new_Jinkela_buffer_8363 (
        .din(new_Jinkela_wire_10304),
        .dout(new_Jinkela_wire_10305)
    );

    bfr new_Jinkela_buffer_4885 (
        .din(new_Jinkela_wire_6316),
        .dout(new_Jinkela_wire_6317)
    );

    bfr new_Jinkela_buffer_8461 (
        .din(new_Jinkela_wire_10410),
        .dout(new_Jinkela_wire_10411)
    );

    bfr new_Jinkela_buffer_8364 (
        .din(new_Jinkela_wire_10305),
        .dout(new_Jinkela_wire_10306)
    );

    bfr new_Jinkela_buffer_4886 (
        .din(new_Jinkela_wire_6317),
        .dout(new_Jinkela_wire_6318)
    );

    bfr new_Jinkela_buffer_8502 (
        .din(new_Jinkela_wire_10453),
        .dout(new_Jinkela_wire_10454)
    );

    bfr new_Jinkela_buffer_5141 (
        .din(_0721_),
        .dout(new_Jinkela_wire_6617)
    );

    bfr new_Jinkela_buffer_4971 (
        .din(new_Jinkela_wire_6430),
        .dout(new_Jinkela_wire_6431)
    );

    bfr new_Jinkela_buffer_8365 (
        .din(new_Jinkela_wire_10306),
        .dout(new_Jinkela_wire_10307)
    );

    bfr new_Jinkela_buffer_4887 (
        .din(new_Jinkela_wire_6318),
        .dout(new_Jinkela_wire_6319)
    );

    bfr new_Jinkela_buffer_8462 (
        .din(new_Jinkela_wire_10411),
        .dout(new_Jinkela_wire_10412)
    );

    bfr new_Jinkela_buffer_5053 (
        .din(new_Jinkela_wire_6524),
        .dout(new_Jinkela_wire_6525)
    );

    bfr new_Jinkela_buffer_8366 (
        .din(new_Jinkela_wire_10307),
        .dout(new_Jinkela_wire_10308)
    );

    bfr new_Jinkela_buffer_4888 (
        .din(new_Jinkela_wire_6319),
        .dout(new_Jinkela_wire_6320)
    );

    bfr new_Jinkela_buffer_8497 (
        .din(new_Jinkela_wire_10446),
        .dout(new_Jinkela_wire_10447)
    );

    bfr new_Jinkela_buffer_4972 (
        .din(new_Jinkela_wire_6431),
        .dout(new_Jinkela_wire_6432)
    );

    bfr new_Jinkela_buffer_8367 (
        .din(new_Jinkela_wire_10308),
        .dout(new_Jinkela_wire_10309)
    );

    bfr new_Jinkela_buffer_4889 (
        .din(new_Jinkela_wire_6320),
        .dout(new_Jinkela_wire_6321)
    );

    bfr new_Jinkela_buffer_8463 (
        .din(new_Jinkela_wire_10412),
        .dout(new_Jinkela_wire_10413)
    );

    bfr new_Jinkela_buffer_8368 (
        .din(new_Jinkela_wire_10309),
        .dout(new_Jinkela_wire_10310)
    );

    bfr new_Jinkela_buffer_4890 (
        .din(new_Jinkela_wire_6321),
        .dout(new_Jinkela_wire_6322)
    );

    spl2 new_Jinkela_splitter_587 (
        .a(_1730_),
        .b(new_Jinkela_wire_6618),
        .c(new_Jinkela_wire_6619)
    );

    spl2 new_Jinkela_splitter_828 (
        .a(_0160_),
        .b(new_Jinkela_wire_10562),
        .c(new_Jinkela_wire_10563)
    );

    bfr new_Jinkela_buffer_4973 (
        .din(new_Jinkela_wire_6432),
        .dout(new_Jinkela_wire_6433)
    );

    bfr new_Jinkela_buffer_8369 (
        .din(new_Jinkela_wire_10310),
        .dout(new_Jinkela_wire_10311)
    );

    bfr new_Jinkela_buffer_4891 (
        .din(new_Jinkela_wire_6322),
        .dout(new_Jinkela_wire_6323)
    );

    bfr new_Jinkela_buffer_8464 (
        .din(new_Jinkela_wire_10413),
        .dout(new_Jinkela_wire_10414)
    );

    bfr new_Jinkela_buffer_5054 (
        .din(new_Jinkela_wire_6525),
        .dout(new_Jinkela_wire_6526)
    );

    bfr new_Jinkela_buffer_8370 (
        .din(new_Jinkela_wire_10311),
        .dout(new_Jinkela_wire_10312)
    );

    bfr new_Jinkela_buffer_4892 (
        .din(new_Jinkela_wire_6323),
        .dout(new_Jinkela_wire_6324)
    );

    bfr new_Jinkela_buffer_8498 (
        .din(new_Jinkela_wire_10447),
        .dout(new_Jinkela_wire_10448)
    );

    bfr new_Jinkela_buffer_4974 (
        .din(new_Jinkela_wire_6433),
        .dout(new_Jinkela_wire_6434)
    );

    bfr new_Jinkela_buffer_8371 (
        .din(new_Jinkela_wire_10312),
        .dout(new_Jinkela_wire_10313)
    );

    bfr new_Jinkela_buffer_4893 (
        .din(new_Jinkela_wire_6324),
        .dout(new_Jinkela_wire_6325)
    );

    bfr new_Jinkela_buffer_8465 (
        .din(new_Jinkela_wire_10414),
        .dout(new_Jinkela_wire_10415)
    );

    bfr new_Jinkela_buffer_5062 (
        .din(new_Jinkela_wire_6535),
        .dout(new_Jinkela_wire_6536)
    );

    bfr new_Jinkela_buffer_8372 (
        .din(new_Jinkela_wire_10313),
        .dout(new_Jinkela_wire_10314)
    );

    bfr new_Jinkela_buffer_4894 (
        .din(new_Jinkela_wire_6325),
        .dout(new_Jinkela_wire_6326)
    );

    bfr new_Jinkela_buffer_8503 (
        .din(new_Jinkela_wire_10454),
        .dout(new_Jinkela_wire_10455)
    );

    bfr new_Jinkela_buffer_5055 (
        .din(new_Jinkela_wire_6526),
        .dout(new_Jinkela_wire_6527)
    );

    bfr new_Jinkela_buffer_4975 (
        .din(new_Jinkela_wire_6434),
        .dout(new_Jinkela_wire_6435)
    );

    bfr new_Jinkela_buffer_8373 (
        .din(new_Jinkela_wire_10314),
        .dout(new_Jinkela_wire_10315)
    );

    bfr new_Jinkela_buffer_4895 (
        .din(new_Jinkela_wire_6326),
        .dout(new_Jinkela_wire_6327)
    );

    bfr new_Jinkela_buffer_8466 (
        .din(new_Jinkela_wire_10415),
        .dout(new_Jinkela_wire_10416)
    );

    bfr new_Jinkela_buffer_8374 (
        .din(new_Jinkela_wire_10315),
        .dout(new_Jinkela_wire_10316)
    );

    bfr new_Jinkela_buffer_4896 (
        .din(new_Jinkela_wire_6327),
        .dout(new_Jinkela_wire_6328)
    );

    spl2 new_Jinkela_splitter_824 (
        .a(new_Jinkela_wire_10448),
        .b(new_Jinkela_wire_10449),
        .c(new_Jinkela_wire_10450)
    );

    bfr new_Jinkela_buffer_4976 (
        .din(new_Jinkela_wire_6435),
        .dout(new_Jinkela_wire_6436)
    );

    bfr new_Jinkela_buffer_8375 (
        .din(new_Jinkela_wire_10316),
        .dout(new_Jinkela_wire_10317)
    );

    bfr new_Jinkela_buffer_4897 (
        .din(new_Jinkela_wire_6328),
        .dout(new_Jinkela_wire_6329)
    );

    bfr new_Jinkela_buffer_8467 (
        .din(new_Jinkela_wire_10416),
        .dout(new_Jinkela_wire_10417)
    );

    bfr new_Jinkela_buffer_5142 (
        .din(_0711_),
        .dout(new_Jinkela_wire_6620)
    );

    bfr new_Jinkela_buffer_8376 (
        .din(new_Jinkela_wire_10317),
        .dout(new_Jinkela_wire_10318)
    );

    bfr new_Jinkela_buffer_4898 (
        .din(new_Jinkela_wire_6329),
        .dout(new_Jinkela_wire_6330)
    );

    bfr new_Jinkela_buffer_8504 (
        .din(new_Jinkela_wire_10455),
        .dout(new_Jinkela_wire_10456)
    );

    bfr new_Jinkela_buffer_4977 (
        .din(new_Jinkela_wire_6436),
        .dout(new_Jinkela_wire_6437)
    );

    bfr new_Jinkela_buffer_8377 (
        .din(new_Jinkela_wire_10318),
        .dout(new_Jinkela_wire_10319)
    );

    bfr new_Jinkela_buffer_4899 (
        .din(new_Jinkela_wire_6330),
        .dout(new_Jinkela_wire_6331)
    );

    bfr new_Jinkela_buffer_8468 (
        .din(new_Jinkela_wire_10417),
        .dout(new_Jinkela_wire_10418)
    );

    bfr new_Jinkela_buffer_5056 (
        .din(new_Jinkela_wire_6527),
        .dout(new_Jinkela_wire_6528)
    );

    bfr new_Jinkela_buffer_8378 (
        .din(new_Jinkela_wire_10319),
        .dout(new_Jinkela_wire_10320)
    );

    bfr new_Jinkela_buffer_4900 (
        .din(new_Jinkela_wire_6331),
        .dout(new_Jinkela_wire_6332)
    );

    spl2 new_Jinkela_splitter_829 (
        .a(_1036_),
        .b(new_Jinkela_wire_10568),
        .c(new_Jinkela_wire_10569)
    );

    bfr new_Jinkela_buffer_4978 (
        .din(new_Jinkela_wire_6437),
        .dout(new_Jinkela_wire_6438)
    );

    bfr new_Jinkela_buffer_8379 (
        .din(new_Jinkela_wire_10320),
        .dout(new_Jinkela_wire_10321)
    );

    bfr new_Jinkela_buffer_4901 (
        .din(new_Jinkela_wire_6332),
        .dout(new_Jinkela_wire_6333)
    );

    bfr new_Jinkela_buffer_8469 (
        .din(new_Jinkela_wire_10418),
        .dout(new_Jinkela_wire_10419)
    );

    bfr new_Jinkela_buffer_5063 (
        .din(new_Jinkela_wire_6536),
        .dout(new_Jinkela_wire_6537)
    );

    bfr new_Jinkela_buffer_8380 (
        .din(new_Jinkela_wire_10321),
        .dout(new_Jinkela_wire_10322)
    );

    bfr new_Jinkela_buffer_4902 (
        .din(new_Jinkela_wire_6333),
        .dout(new_Jinkela_wire_6334)
    );

    bfr new_Jinkela_buffer_8604 (
        .din(new_Jinkela_wire_10563),
        .dout(new_Jinkela_wire_10564)
    );

    spl2 new_Jinkela_splitter_830 (
        .a(_0589_),
        .b(new_Jinkela_wire_10574),
        .c(new_Jinkela_wire_10575)
    );

    spl2 new_Jinkela_splitter_1330 (
        .a(_0405_),
        .b(new_Jinkela_wire_18387),
        .c(new_Jinkela_wire_18388)
    );

    bfr new_Jinkela_buffer_15420 (
        .din(new_Jinkela_wire_18382),
        .dout(new_Jinkela_wire_18383)
    );

    bfr new_Jinkela_buffer_15276 (
        .din(new_Jinkela_wire_18210),
        .dout(new_Jinkela_wire_18211)
    );

    bfr new_Jinkela_buffer_15328 (
        .din(new_Jinkela_wire_18268),
        .dout(new_Jinkela_wire_18269)
    );

    bfr new_Jinkela_buffer_15277 (
        .din(new_Jinkela_wire_18211),
        .dout(new_Jinkela_wire_18212)
    );

    bfr new_Jinkela_buffer_15365 (
        .din(new_Jinkela_wire_18319),
        .dout(new_Jinkela_wire_18320)
    );

    bfr new_Jinkela_buffer_15278 (
        .din(new_Jinkela_wire_18212),
        .dout(new_Jinkela_wire_18213)
    );

    bfr new_Jinkela_buffer_15329 (
        .din(new_Jinkela_wire_18269),
        .dout(new_Jinkela_wire_18270)
    );

    bfr new_Jinkela_buffer_15279 (
        .din(new_Jinkela_wire_18213),
        .dout(new_Jinkela_wire_18214)
    );

    bfr new_Jinkela_buffer_15280 (
        .din(new_Jinkela_wire_18214),
        .dout(new_Jinkela_wire_18215)
    );

    bfr new_Jinkela_buffer_15330 (
        .din(new_Jinkela_wire_18270),
        .dout(new_Jinkela_wire_18271)
    );

    bfr new_Jinkela_buffer_15281 (
        .din(new_Jinkela_wire_18215),
        .dout(new_Jinkela_wire_18216)
    );

    bfr new_Jinkela_buffer_15366 (
        .din(new_Jinkela_wire_18320),
        .dout(new_Jinkela_wire_18321)
    );

    bfr new_Jinkela_buffer_15282 (
        .din(new_Jinkela_wire_18216),
        .dout(new_Jinkela_wire_18217)
    );

    bfr new_Jinkela_buffer_15331 (
        .din(new_Jinkela_wire_18271),
        .dout(new_Jinkela_wire_18272)
    );

    bfr new_Jinkela_buffer_15283 (
        .din(new_Jinkela_wire_18217),
        .dout(new_Jinkela_wire_18218)
    );

    spl2 new_Jinkela_splitter_1331 (
        .a(_1352_),
        .b(new_Jinkela_wire_18393),
        .c(new_Jinkela_wire_18394)
    );

    bfr new_Jinkela_buffer_15284 (
        .din(new_Jinkela_wire_18218),
        .dout(new_Jinkela_wire_18219)
    );

    bfr new_Jinkela_buffer_15332 (
        .din(new_Jinkela_wire_18272),
        .dout(new_Jinkela_wire_18273)
    );

    spl2 new_Jinkela_splitter_1316 (
        .a(new_Jinkela_wire_18219),
        .b(new_Jinkela_wire_18220),
        .c(new_Jinkela_wire_18221)
    );

    bfr new_Jinkela_buffer_15333 (
        .din(new_Jinkela_wire_18273),
        .dout(new_Jinkela_wire_18274)
    );

    bfr new_Jinkela_buffer_15367 (
        .din(new_Jinkela_wire_18321),
        .dout(new_Jinkela_wire_18322)
    );

    spl2 new_Jinkela_splitter_1319 (
        .a(new_Jinkela_wire_18274),
        .b(new_Jinkela_wire_18275),
        .c(new_Jinkela_wire_18276)
    );

    bfr new_Jinkela_buffer_15421 (
        .din(new_Jinkela_wire_18383),
        .dout(new_Jinkela_wire_18384)
    );

    bfr new_Jinkela_buffer_15368 (
        .din(new_Jinkela_wire_18322),
        .dout(new_Jinkela_wire_18323)
    );

    bfr new_Jinkela_buffer_15369 (
        .din(new_Jinkela_wire_18323),
        .dout(new_Jinkela_wire_18324)
    );

    bfr new_Jinkela_buffer_15424 (
        .din(new_Jinkela_wire_18388),
        .dout(new_Jinkela_wire_18389)
    );

    bfr new_Jinkela_buffer_15428 (
        .din(_0229_),
        .dout(new_Jinkela_wire_18395)
    );

    bfr new_Jinkela_buffer_15370 (
        .din(new_Jinkela_wire_18324),
        .dout(new_Jinkela_wire_18325)
    );

    bfr new_Jinkela_buffer_15422 (
        .din(new_Jinkela_wire_18384),
        .dout(new_Jinkela_wire_18385)
    );

    bfr new_Jinkela_buffer_15371 (
        .din(new_Jinkela_wire_18325),
        .dout(new_Jinkela_wire_18326)
    );

    spl2 new_Jinkela_splitter_1333 (
        .a(_0354_),
        .b(new_Jinkela_wire_18446),
        .c(new_Jinkela_wire_18447)
    );

    bfr new_Jinkela_buffer_15372 (
        .din(new_Jinkela_wire_18326),
        .dout(new_Jinkela_wire_18327)
    );

    bfr new_Jinkela_buffer_15423 (
        .din(new_Jinkela_wire_18385),
        .dout(new_Jinkela_wire_18386)
    );

    bfr new_Jinkela_buffer_15373 (
        .din(new_Jinkela_wire_18327),
        .dout(new_Jinkela_wire_18328)
    );

    bfr new_Jinkela_buffer_15425 (
        .din(new_Jinkela_wire_18389),
        .dout(new_Jinkela_wire_18390)
    );

    bfr new_Jinkela_buffer_15374 (
        .din(new_Jinkela_wire_18328),
        .dout(new_Jinkela_wire_18329)
    );

    bfr new_Jinkela_buffer_15476 (
        .din(_1708_),
        .dout(new_Jinkela_wire_18445)
    );

    bfr new_Jinkela_buffer_15375 (
        .din(new_Jinkela_wire_18329),
        .dout(new_Jinkela_wire_18330)
    );

    bfr new_Jinkela_buffer_15426 (
        .din(new_Jinkela_wire_18390),
        .dout(new_Jinkela_wire_18391)
    );

    bfr new_Jinkela_buffer_15376 (
        .din(new_Jinkela_wire_18330),
        .dout(new_Jinkela_wire_18331)
    );

    bfr new_Jinkela_buffer_15429 (
        .din(new_Jinkela_wire_18395),
        .dout(new_Jinkela_wire_18396)
    );

    bfr new_Jinkela_buffer_8381 (
        .din(new_Jinkela_wire_10322),
        .dout(new_Jinkela_wire_10323)
    );

    bfr new_Jinkela_buffer_8470 (
        .din(new_Jinkela_wire_10419),
        .dout(new_Jinkela_wire_10420)
    );

    bfr new_Jinkela_buffer_8382 (
        .din(new_Jinkela_wire_10323),
        .dout(new_Jinkela_wire_10324)
    );

    bfr new_Jinkela_buffer_8505 (
        .din(new_Jinkela_wire_10456),
        .dout(new_Jinkela_wire_10457)
    );

    bfr new_Jinkela_buffer_8383 (
        .din(new_Jinkela_wire_10324),
        .dout(new_Jinkela_wire_10325)
    );

    bfr new_Jinkela_buffer_8471 (
        .din(new_Jinkela_wire_10420),
        .dout(new_Jinkela_wire_10421)
    );

    bfr new_Jinkela_buffer_8384 (
        .din(new_Jinkela_wire_10325),
        .dout(new_Jinkela_wire_10326)
    );

    bfr new_Jinkela_buffer_8608 (
        .din(new_Jinkela_wire_10569),
        .dout(new_Jinkela_wire_10570)
    );

    bfr new_Jinkela_buffer_8385 (
        .din(new_Jinkela_wire_10326),
        .dout(new_Jinkela_wire_10327)
    );

    bfr new_Jinkela_buffer_8472 (
        .din(new_Jinkela_wire_10421),
        .dout(new_Jinkela_wire_10422)
    );

    bfr new_Jinkela_buffer_8386 (
        .din(new_Jinkela_wire_10327),
        .dout(new_Jinkela_wire_10328)
    );

    bfr new_Jinkela_buffer_8506 (
        .din(new_Jinkela_wire_10457),
        .dout(new_Jinkela_wire_10458)
    );

    bfr new_Jinkela_buffer_8387 (
        .din(new_Jinkela_wire_10328),
        .dout(new_Jinkela_wire_10329)
    );

    bfr new_Jinkela_buffer_8473 (
        .din(new_Jinkela_wire_10422),
        .dout(new_Jinkela_wire_10423)
    );

    bfr new_Jinkela_buffer_8388 (
        .din(new_Jinkela_wire_10329),
        .dout(new_Jinkela_wire_10330)
    );

    bfr new_Jinkela_buffer_8605 (
        .din(new_Jinkela_wire_10564),
        .dout(new_Jinkela_wire_10565)
    );

    bfr new_Jinkela_buffer_8389 (
        .din(new_Jinkela_wire_10330),
        .dout(new_Jinkela_wire_10331)
    );

    bfr new_Jinkela_buffer_8474 (
        .din(new_Jinkela_wire_10423),
        .dout(new_Jinkela_wire_10424)
    );

    bfr new_Jinkela_buffer_8390 (
        .din(new_Jinkela_wire_10331),
        .dout(new_Jinkela_wire_10332)
    );

    bfr new_Jinkela_buffer_8507 (
        .din(new_Jinkela_wire_10458),
        .dout(new_Jinkela_wire_10459)
    );

    bfr new_Jinkela_buffer_8391 (
        .din(new_Jinkela_wire_10332),
        .dout(new_Jinkela_wire_10333)
    );

    bfr new_Jinkela_buffer_8475 (
        .din(new_Jinkela_wire_10424),
        .dout(new_Jinkela_wire_10425)
    );

    bfr new_Jinkela_buffer_8392 (
        .din(new_Jinkela_wire_10333),
        .dout(new_Jinkela_wire_10334)
    );

    bfr new_Jinkela_buffer_8616 (
        .din(_1290_),
        .dout(new_Jinkela_wire_10580)
    );

    bfr new_Jinkela_buffer_8393 (
        .din(new_Jinkela_wire_10334),
        .dout(new_Jinkela_wire_10335)
    );

    bfr new_Jinkela_buffer_8476 (
        .din(new_Jinkela_wire_10425),
        .dout(new_Jinkela_wire_10426)
    );

    bfr new_Jinkela_buffer_8394 (
        .din(new_Jinkela_wire_10335),
        .dout(new_Jinkela_wire_10336)
    );

    bfr new_Jinkela_buffer_8508 (
        .din(new_Jinkela_wire_10459),
        .dout(new_Jinkela_wire_10460)
    );

    bfr new_Jinkela_buffer_8395 (
        .din(new_Jinkela_wire_10336),
        .dout(new_Jinkela_wire_10337)
    );

    bfr new_Jinkela_buffer_8477 (
        .din(new_Jinkela_wire_10426),
        .dout(new_Jinkela_wire_10427)
    );

    bfr new_Jinkela_buffer_8396 (
        .din(new_Jinkela_wire_10337),
        .dout(new_Jinkela_wire_10338)
    );

    bfr new_Jinkela_buffer_8606 (
        .din(new_Jinkela_wire_10565),
        .dout(new_Jinkela_wire_10566)
    );

    bfr new_Jinkela_buffer_8397 (
        .din(new_Jinkela_wire_10338),
        .dout(new_Jinkela_wire_10339)
    );

    bfr new_Jinkela_buffer_8478 (
        .din(new_Jinkela_wire_10427),
        .dout(new_Jinkela_wire_10428)
    );

    bfr new_Jinkela_buffer_8398 (
        .din(new_Jinkela_wire_10339),
        .dout(new_Jinkela_wire_10340)
    );

    bfr new_Jinkela_buffer_8509 (
        .din(new_Jinkela_wire_10460),
        .dout(new_Jinkela_wire_10461)
    );

    bfr new_Jinkela_buffer_8399 (
        .din(new_Jinkela_wire_10340),
        .dout(new_Jinkela_wire_10341)
    );

    bfr new_Jinkela_buffer_8479 (
        .din(new_Jinkela_wire_10428),
        .dout(new_Jinkela_wire_10429)
    );

    bfr new_Jinkela_buffer_8400 (
        .din(new_Jinkela_wire_10341),
        .dout(new_Jinkela_wire_10342)
    );

    bfr new_Jinkela_buffer_8612 (
        .din(new_Jinkela_wire_10575),
        .dout(new_Jinkela_wire_10576)
    );

    bfr new_Jinkela_buffer_8401 (
        .din(new_Jinkela_wire_10342),
        .dout(new_Jinkela_wire_10343)
    );

    bfr new_Jinkela_buffer_8480 (
        .din(new_Jinkela_wire_10429),
        .dout(new_Jinkela_wire_10430)
    );

    bfr new_Jinkela_buffer_4979 (
        .din(new_Jinkela_wire_6438),
        .dout(new_Jinkela_wire_6439)
    );

    bfr new_Jinkela_buffer_4903 (
        .din(new_Jinkela_wire_6334),
        .dout(new_Jinkela_wire_6335)
    );

    bfr new_Jinkela_buffer_5057 (
        .din(new_Jinkela_wire_6528),
        .dout(new_Jinkela_wire_6529)
    );

    bfr new_Jinkela_buffer_4904 (
        .din(new_Jinkela_wire_6335),
        .dout(new_Jinkela_wire_6336)
    );

    bfr new_Jinkela_buffer_4980 (
        .din(new_Jinkela_wire_6439),
        .dout(new_Jinkela_wire_6440)
    );

    bfr new_Jinkela_buffer_4905 (
        .din(new_Jinkela_wire_6336),
        .dout(new_Jinkela_wire_6337)
    );

    bfr new_Jinkela_buffer_4906 (
        .din(new_Jinkela_wire_6337),
        .dout(new_Jinkela_wire_6338)
    );

    bfr new_Jinkela_buffer_5196 (
        .din(_0283_),
        .dout(new_Jinkela_wire_6678)
    );

    bfr new_Jinkela_buffer_4981 (
        .din(new_Jinkela_wire_6440),
        .dout(new_Jinkela_wire_6441)
    );

    bfr new_Jinkela_buffer_4907 (
        .din(new_Jinkela_wire_6338),
        .dout(new_Jinkela_wire_6339)
    );

    bfr new_Jinkela_buffer_5058 (
        .din(new_Jinkela_wire_6529),
        .dout(new_Jinkela_wire_6530)
    );

    bfr new_Jinkela_buffer_4908 (
        .din(new_Jinkela_wire_6339),
        .dout(new_Jinkela_wire_6340)
    );

    bfr new_Jinkela_buffer_4982 (
        .din(new_Jinkela_wire_6441),
        .dout(new_Jinkela_wire_6442)
    );

    bfr new_Jinkela_buffer_4909 (
        .din(new_Jinkela_wire_6340),
        .dout(new_Jinkela_wire_6341)
    );

    bfr new_Jinkela_buffer_5064 (
        .din(new_Jinkela_wire_6537),
        .dout(new_Jinkela_wire_6538)
    );

    bfr new_Jinkela_buffer_4910 (
        .din(new_Jinkela_wire_6341),
        .dout(new_Jinkela_wire_6342)
    );

    bfr new_Jinkela_buffer_4983 (
        .din(new_Jinkela_wire_6442),
        .dout(new_Jinkela_wire_6443)
    );

    bfr new_Jinkela_buffer_4911 (
        .din(new_Jinkela_wire_6342),
        .dout(new_Jinkela_wire_6343)
    );

    bfr new_Jinkela_buffer_5059 (
        .din(new_Jinkela_wire_6530),
        .dout(new_Jinkela_wire_6531)
    );

    bfr new_Jinkela_buffer_4912 (
        .din(new_Jinkela_wire_6343),
        .dout(new_Jinkela_wire_6344)
    );

    bfr new_Jinkela_buffer_4984 (
        .din(new_Jinkela_wire_6443),
        .dout(new_Jinkela_wire_6444)
    );

    bfr new_Jinkela_buffer_4913 (
        .din(new_Jinkela_wire_6344),
        .dout(new_Jinkela_wire_6345)
    );

    bfr new_Jinkela_buffer_4914 (
        .din(new_Jinkela_wire_6345),
        .dout(new_Jinkela_wire_6346)
    );

    spl2 new_Jinkela_splitter_589 (
        .a(_1645_),
        .b(new_Jinkela_wire_6676),
        .c(new_Jinkela_wire_6677)
    );

    bfr new_Jinkela_buffer_4985 (
        .din(new_Jinkela_wire_6444),
        .dout(new_Jinkela_wire_6445)
    );

    bfr new_Jinkela_buffer_4915 (
        .din(new_Jinkela_wire_6346),
        .dout(new_Jinkela_wire_6347)
    );

    bfr new_Jinkela_buffer_5060 (
        .din(new_Jinkela_wire_6531),
        .dout(new_Jinkela_wire_6532)
    );

    bfr new_Jinkela_buffer_4916 (
        .din(new_Jinkela_wire_6347),
        .dout(new_Jinkela_wire_6348)
    );

    bfr new_Jinkela_buffer_4986 (
        .din(new_Jinkela_wire_6445),
        .dout(new_Jinkela_wire_6446)
    );

    bfr new_Jinkela_buffer_4917 (
        .din(new_Jinkela_wire_6348),
        .dout(new_Jinkela_wire_6349)
    );

    bfr new_Jinkela_buffer_5065 (
        .din(new_Jinkela_wire_6538),
        .dout(new_Jinkela_wire_6539)
    );

    bfr new_Jinkela_buffer_4918 (
        .din(new_Jinkela_wire_6349),
        .dout(new_Jinkela_wire_6350)
    );

    bfr new_Jinkela_buffer_4987 (
        .din(new_Jinkela_wire_6446),
        .dout(new_Jinkela_wire_6447)
    );

    bfr new_Jinkela_buffer_4919 (
        .din(new_Jinkela_wire_6350),
        .dout(new_Jinkela_wire_6351)
    );

    spl2 new_Jinkela_splitter_585 (
        .a(new_Jinkela_wire_6532),
        .b(new_Jinkela_wire_6533),
        .c(new_Jinkela_wire_6534)
    );

    bfr new_Jinkela_buffer_4920 (
        .din(new_Jinkela_wire_6351),
        .dout(new_Jinkela_wire_6352)
    );

    bfr new_Jinkela_buffer_4988 (
        .din(new_Jinkela_wire_6447),
        .dout(new_Jinkela_wire_6448)
    );

    bfr new_Jinkela_buffer_4921 (
        .din(new_Jinkela_wire_6352),
        .dout(new_Jinkela_wire_6353)
    );

    bfr new_Jinkela_buffer_5143 (
        .din(new_Jinkela_wire_6620),
        .dout(new_Jinkela_wire_6621)
    );

    bfr new_Jinkela_buffer_4922 (
        .din(new_Jinkela_wire_6353),
        .dout(new_Jinkela_wire_6354)
    );

    bfr new_Jinkela_buffer_4989 (
        .din(new_Jinkela_wire_6448),
        .dout(new_Jinkela_wire_6449)
    );

    bfr new_Jinkela_buffer_4923 (
        .din(new_Jinkela_wire_6354),
        .dout(new_Jinkela_wire_6355)
    );

    bfr new_Jinkela_buffer_11858 (
        .din(_1807_),
        .dout(new_Jinkela_wire_14330)
    );

    and_bb _2539_ (
        .a(new_Jinkela_wire_384),
        .b(new_Jinkela_wire_619),
        .c(_1584_)
    );

    bfr new_Jinkela_buffer_11855 (
        .din(new_Jinkela_wire_14322),
        .dout(new_Jinkela_wire_14323)
    );

    and_bi _2540_ (
        .a(new_Jinkela_wire_18768),
        .b(new_Jinkela_wire_19157),
        .c(_1585_)
    );

    bfr new_Jinkela_buffer_11955 (
        .din(_0077_),
        .dout(new_Jinkela_wire_14429)
    );

    and_bb _2541_ (
        .a(new_Jinkela_wire_403),
        .b(new_Jinkela_wire_547),
        .c(_1586_)
    );

    bfr new_Jinkela_buffer_11856 (
        .din(new_Jinkela_wire_14323),
        .dout(new_Jinkela_wire_14324)
    );

    or_ii _2542_ (
        .a(new_Jinkela_wire_598),
        .b(new_Jinkela_wire_325),
        .c(_1587_)
    );

    or_bb _2543_ (
        .a(new_Jinkela_wire_17109),
        .b(new_Jinkela_wire_19541),
        .c(_1589_)
    );

    bfr new_Jinkela_buffer_11954 (
        .din(_0359_),
        .dout(new_Jinkela_wire_14428)
    );

    bfr new_Jinkela_buffer_11859 (
        .din(new_Jinkela_wire_14330),
        .dout(new_Jinkela_wire_14331)
    );

    and_bb _2544_ (
        .a(new_Jinkela_wire_607),
        .b(new_Jinkela_wire_231),
        .c(_1590_)
    );

    and_bi _2545_ (
        .a(new_Jinkela_wire_17088),
        .b(new_Jinkela_wire_18971),
        .c(_1591_)
    );

    bfr new_Jinkela_buffer_11956 (
        .din(_0987_),
        .dout(new_Jinkela_wire_14430)
    );

    bfr new_Jinkela_buffer_11860 (
        .din(new_Jinkela_wire_14331),
        .dout(new_Jinkela_wire_14332)
    );

    and_bi _2546_ (
        .a(new_Jinkela_wire_11456),
        .b(new_Jinkela_wire_18522),
        .c(_1592_)
    );

    spl2 new_Jinkela_splitter_1087 (
        .a(_0713_),
        .b(new_Jinkela_wire_14538),
        .c(new_Jinkela_wire_14539)
    );

    or_bb _2547_ (
        .a(new_Jinkela_wire_1594),
        .b(new_Jinkela_wire_19929),
        .c(_1593_)
    );

    bfr new_Jinkela_buffer_11861 (
        .din(new_Jinkela_wire_14332),
        .dout(new_Jinkela_wire_14333)
    );

    or_ii _2548_ (
        .a(new_Jinkela_wire_1595),
        .b(new_Jinkela_wire_19928),
        .c(_1594_)
    );

    or_ii _2549_ (
        .a(new_Jinkela_wire_5157),
        .b(new_Jinkela_wire_19284),
        .c(_1595_)
    );

    bfr new_Jinkela_buffer_12066 (
        .din(new_net_3966),
        .dout(new_Jinkela_wire_14544)
    );

    bfr new_Jinkela_buffer_11862 (
        .din(new_Jinkela_wire_14333),
        .dout(new_Jinkela_wire_14334)
    );

    and_ii _2550_ (
        .a(new_Jinkela_wire_16955),
        .b(new_Jinkela_wire_9518),
        .c(_1596_)
    );

    bfr new_Jinkela_buffer_11957 (
        .din(new_Jinkela_wire_14430),
        .dout(new_Jinkela_wire_14431)
    );

    and_bb _2551_ (
        .a(new_Jinkela_wire_16956),
        .b(new_Jinkela_wire_9519),
        .c(_1597_)
    );

    bfr new_Jinkela_buffer_11863 (
        .din(new_Jinkela_wire_14334),
        .dout(new_Jinkela_wire_14335)
    );

    or_bb _2552_ (
        .a(new_Jinkela_wire_8207),
        .b(new_Jinkela_wire_14019),
        .c(_1598_)
    );

    or_bb _2553_ (
        .a(new_Jinkela_wire_1391),
        .b(new_Jinkela_wire_11442),
        .c(_1600_)
    );

    bfr new_Jinkela_buffer_11864 (
        .din(new_Jinkela_wire_14335),
        .dout(new_Jinkela_wire_14336)
    );

    or_ii _2554_ (
        .a(new_Jinkela_wire_1392),
        .b(new_Jinkela_wire_11443),
        .c(_1601_)
    );

    bfr new_Jinkela_buffer_11958 (
        .din(new_Jinkela_wire_14431),
        .dout(new_Jinkela_wire_14432)
    );

    or_ii _2555_ (
        .a(new_Jinkela_wire_13057),
        .b(new_Jinkela_wire_16125),
        .c(_1602_)
    );

    bfr new_Jinkela_buffer_11865 (
        .din(new_Jinkela_wire_14336),
        .dout(new_Jinkela_wire_14337)
    );

    and_ii _2556_ (
        .a(new_Jinkela_wire_5812),
        .b(new_Jinkela_wire_6755),
        .c(_1603_)
    );

    bfr new_Jinkela_buffer_12062 (
        .din(new_Jinkela_wire_14539),
        .dout(new_Jinkela_wire_14540)
    );

    and_bb _2557_ (
        .a(new_Jinkela_wire_5813),
        .b(new_Jinkela_wire_6756),
        .c(_1604_)
    );

    bfr new_Jinkela_buffer_12102 (
        .din(new_net_3962),
        .dout(new_Jinkela_wire_14580)
    );

    bfr new_Jinkela_buffer_11866 (
        .din(new_Jinkela_wire_14337),
        .dout(new_Jinkela_wire_14338)
    );

    or_bb _2558_ (
        .a(new_Jinkela_wire_2149),
        .b(new_Jinkela_wire_4986),
        .c(_1605_)
    );

    bfr new_Jinkela_buffer_11959 (
        .din(new_Jinkela_wire_14432),
        .dout(new_Jinkela_wire_14433)
    );

    or_bb _2559_ (
        .a(new_Jinkela_wire_20381),
        .b(new_Jinkela_wire_6512),
        .c(_1606_)
    );

    bfr new_Jinkela_buffer_11867 (
        .din(new_Jinkela_wire_14338),
        .dout(new_Jinkela_wire_14339)
    );

    or_ii _2560_ (
        .a(new_Jinkela_wire_20382),
        .b(new_Jinkela_wire_6513),
        .c(_1607_)
    );

    or_ii _2561_ (
        .a(new_Jinkela_wire_7186),
        .b(new_Jinkela_wire_12105),
        .c(_1608_)
    );

    bfr new_Jinkela_buffer_12067 (
        .din(new_Jinkela_wire_14544),
        .dout(new_Jinkela_wire_14545)
    );

    bfr new_Jinkela_buffer_11868 (
        .din(new_Jinkela_wire_14339),
        .dout(new_Jinkela_wire_14340)
    );

    and_ii _2562_ (
        .a(new_Jinkela_wire_18122),
        .b(new_Jinkela_wire_16997),
        .c(_1609_)
    );

    bfr new_Jinkela_buffer_11960 (
        .din(new_Jinkela_wire_14433),
        .dout(new_Jinkela_wire_14434)
    );

    and_bb _2563_ (
        .a(new_Jinkela_wire_18123),
        .b(new_Jinkela_wire_16998),
        .c(_1611_)
    );

    bfr new_Jinkela_buffer_11869 (
        .din(new_Jinkela_wire_14340),
        .dout(new_Jinkela_wire_14341)
    );

    or_bb _2564_ (
        .a(new_Jinkela_wire_13999),
        .b(new_Jinkela_wire_4717),
        .c(_1612_)
    );

    bfr new_Jinkela_buffer_12063 (
        .din(new_Jinkela_wire_14540),
        .dout(new_Jinkela_wire_14541)
    );

    or_bb _2565_ (
        .a(new_Jinkela_wire_18942),
        .b(new_Jinkela_wire_17085),
        .c(_1613_)
    );

    bfr new_Jinkela_buffer_11870 (
        .din(new_Jinkela_wire_14341),
        .dout(new_Jinkela_wire_14342)
    );

    or_ii _2566_ (
        .a(new_Jinkela_wire_18943),
        .b(new_Jinkela_wire_17086),
        .c(_1614_)
    );

    bfr new_Jinkela_buffer_11961 (
        .din(new_Jinkela_wire_14434),
        .dout(new_Jinkela_wire_14435)
    );

    or_ii _2567_ (
        .a(new_Jinkela_wire_19910),
        .b(new_Jinkela_wire_10957),
        .c(_1615_)
    );

    bfr new_Jinkela_buffer_11871 (
        .din(new_Jinkela_wire_14342),
        .dout(new_Jinkela_wire_14343)
    );

    and_ii _2568_ (
        .a(new_Jinkela_wire_20960),
        .b(new_Jinkela_wire_12101),
        .c(_1616_)
    );

    and_bb _2569_ (
        .a(new_Jinkela_wire_20961),
        .b(new_Jinkela_wire_12102),
        .c(_1617_)
    );

    spl2 new_Jinkela_splitter_1088 (
        .a(_1757_),
        .b(new_Jinkela_wire_14656),
        .c(new_Jinkela_wire_14657)
    );

    bfr new_Jinkela_buffer_11872 (
        .din(new_Jinkela_wire_14343),
        .dout(new_Jinkela_wire_14344)
    );

    or_bb _2570_ (
        .a(new_Jinkela_wire_8682),
        .b(new_Jinkela_wire_16102),
        .c(_1618_)
    );

    bfr new_Jinkela_buffer_11962 (
        .din(new_Jinkela_wire_14435),
        .dout(new_Jinkela_wire_14436)
    );

    or_bb _2571_ (
        .a(new_Jinkela_wire_10081),
        .b(new_Jinkela_wire_4243),
        .c(_1619_)
    );

    bfr new_Jinkela_buffer_11873 (
        .din(new_Jinkela_wire_14344),
        .dout(new_Jinkela_wire_14345)
    );

    or_ii _2572_ (
        .a(new_Jinkela_wire_10082),
        .b(new_Jinkela_wire_4244),
        .c(_1620_)
    );

    bfr new_Jinkela_buffer_12064 (
        .din(new_Jinkela_wire_14541),
        .dout(new_Jinkela_wire_14542)
    );

    or_ii _2573_ (
        .a(new_Jinkela_wire_17542),
        .b(new_Jinkela_wire_4682),
        .c(_1622_)
    );

    bfr new_Jinkela_buffer_11874 (
        .din(new_Jinkela_wire_14345),
        .dout(new_Jinkela_wire_14346)
    );

    and_ii _2574_ (
        .a(new_Jinkela_wire_1573),
        .b(new_Jinkela_wire_3237),
        .c(_1623_)
    );

    bfr new_Jinkela_buffer_11963 (
        .din(new_Jinkela_wire_14436),
        .dout(new_Jinkela_wire_14437)
    );

    and_bb _2575_ (
        .a(new_Jinkela_wire_1574),
        .b(new_Jinkela_wire_3238),
        .c(_1624_)
    );

    bfr new_Jinkela_buffer_11875 (
        .din(new_Jinkela_wire_14346),
        .dout(new_Jinkela_wire_14347)
    );

    or_bb _2576_ (
        .a(new_Jinkela_wire_4677),
        .b(new_Jinkela_wire_12711),
        .c(_1625_)
    );

    spl2 new_Jinkela_splitter_1089 (
        .a(_0758_),
        .b(new_Jinkela_wire_14658),
        .c(new_Jinkela_wire_14659)
    );

    or_bb _2577_ (
        .a(new_Jinkela_wire_15554),
        .b(new_Jinkela_wire_16951),
        .c(_1626_)
    );

    bfr new_Jinkela_buffer_12068 (
        .din(new_Jinkela_wire_14545),
        .dout(new_Jinkela_wire_14546)
    );

    bfr new_Jinkela_buffer_11876 (
        .din(new_Jinkela_wire_14347),
        .dout(new_Jinkela_wire_14348)
    );

    or_ii _2578_ (
        .a(new_Jinkela_wire_15555),
        .b(new_Jinkela_wire_16952),
        .c(_1627_)
    );

    bfr new_Jinkela_buffer_11964 (
        .din(new_Jinkela_wire_14437),
        .dout(new_Jinkela_wire_14438)
    );

    or_ii _2579_ (
        .a(new_Jinkela_wire_2952),
        .b(new_Jinkela_wire_12331),
        .c(_1628_)
    );

    bfr new_Jinkela_buffer_11877 (
        .din(new_Jinkela_wire_14348),
        .dout(new_Jinkela_wire_14349)
    );

    and_ii _2580_ (
        .a(new_Jinkela_wire_11454),
        .b(new_Jinkela_wire_12219),
        .c(_1629_)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(new_Jinkela_wire_2284),
        .dout(new_Jinkela_wire_2285)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_2206),
        .dout(new_Jinkela_wire_2207)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_2345),
        .dout(new_Jinkela_wire_2346)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_2207),
        .dout(new_Jinkela_wire_2208)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(new_Jinkela_wire_2285),
        .dout(new_Jinkela_wire_2286)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(new_Jinkela_wire_2208),
        .dout(new_Jinkela_wire_2209)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(new_Jinkela_wire_2336),
        .dout(new_Jinkela_wire_2337)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_2209),
        .dout(new_Jinkela_wire_2210)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(new_Jinkela_wire_2286),
        .dout(new_Jinkela_wire_2287)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_2210),
        .dout(new_Jinkela_wire_2211)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(_1076_),
        .dout(new_Jinkela_wire_2423)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(new_Jinkela_wire_2211),
        .dout(new_Jinkela_wire_2212)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(new_Jinkela_wire_2287),
        .dout(new_Jinkela_wire_2288)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(new_Jinkela_wire_2212),
        .dout(new_Jinkela_wire_2213)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(new_Jinkela_wire_2337),
        .dout(new_Jinkela_wire_2338)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_2213),
        .dout(new_Jinkela_wire_2214)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(new_Jinkela_wire_2288),
        .dout(new_Jinkela_wire_2289)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_2214),
        .dout(new_Jinkela_wire_2215)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(new_Jinkela_wire_2346),
        .dout(new_Jinkela_wire_2347)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_2215),
        .dout(new_Jinkela_wire_2216)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_2289),
        .dout(new_Jinkela_wire_2290)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(new_Jinkela_wire_2216),
        .dout(new_Jinkela_wire_2217)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_Jinkela_wire_2338),
        .dout(new_Jinkela_wire_2339)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(new_Jinkela_wire_2217),
        .dout(new_Jinkela_wire_2218)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(new_Jinkela_wire_2290),
        .dout(new_Jinkela_wire_2291)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_2218),
        .dout(new_Jinkela_wire_2219)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(_1533_),
        .dout(new_Jinkela_wire_2422)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(new_Jinkela_wire_2219),
        .dout(new_Jinkela_wire_2220)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_2291),
        .dout(new_Jinkela_wire_2292)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(new_Jinkela_wire_2220),
        .dout(new_Jinkela_wire_2221)
    );

    spl2 new_Jinkela_splitter_286 (
        .a(new_Jinkela_wire_2339),
        .b(new_Jinkela_wire_2340),
        .c(new_Jinkela_wire_2341)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(new_Jinkela_wire_2221),
        .dout(new_Jinkela_wire_2222)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_2292),
        .dout(new_Jinkela_wire_2293)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_2222),
        .dout(new_Jinkela_wire_2223)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(_0760_),
        .dout(new_Jinkela_wire_2457)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(new_Jinkela_wire_2223),
        .dout(new_Jinkela_wire_2224)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_2293),
        .dout(new_Jinkela_wire_2294)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(new_Jinkela_wire_2224),
        .dout(new_Jinkela_wire_2225)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(new_Jinkela_wire_2347),
        .dout(new_Jinkela_wire_2348)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(new_Jinkela_wire_2225),
        .dout(new_Jinkela_wire_2226)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_2294),
        .dout(new_Jinkela_wire_2295)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_Jinkela_wire_2226),
        .dout(new_Jinkela_wire_2227)
    );

    bfr new_Jinkela_buffer_5066 (
        .din(new_Jinkela_wire_6539),
        .dout(new_Jinkela_wire_6540)
    );

    bfr new_Jinkela_buffer_4924 (
        .din(new_Jinkela_wire_6355),
        .dout(new_Jinkela_wire_6356)
    );

    bfr new_Jinkela_buffer_4990 (
        .din(new_Jinkela_wire_6449),
        .dout(new_Jinkela_wire_6450)
    );

    bfr new_Jinkela_buffer_4925 (
        .din(new_Jinkela_wire_6356),
        .dout(new_Jinkela_wire_6357)
    );

    bfr new_Jinkela_buffer_4926 (
        .din(new_Jinkela_wire_6357),
        .dout(new_Jinkela_wire_6358)
    );

    spl2 new_Jinkela_splitter_590 (
        .a(_0169_),
        .b(new_Jinkela_wire_6680),
        .c(new_Jinkela_wire_6681)
    );

    bfr new_Jinkela_buffer_4991 (
        .din(new_Jinkela_wire_6450),
        .dout(new_Jinkela_wire_6451)
    );

    bfr new_Jinkela_buffer_4927 (
        .din(new_Jinkela_wire_6358),
        .dout(new_Jinkela_wire_6359)
    );

    bfr new_Jinkela_buffer_5067 (
        .din(new_Jinkela_wire_6540),
        .dout(new_Jinkela_wire_6541)
    );

    bfr new_Jinkela_buffer_4928 (
        .din(new_Jinkela_wire_6359),
        .dout(new_Jinkela_wire_6360)
    );

    bfr new_Jinkela_buffer_4992 (
        .din(new_Jinkela_wire_6451),
        .dout(new_Jinkela_wire_6452)
    );

    bfr new_Jinkela_buffer_4929 (
        .din(new_Jinkela_wire_6360),
        .dout(new_Jinkela_wire_6361)
    );

    bfr new_Jinkela_buffer_5144 (
        .din(new_Jinkela_wire_6621),
        .dout(new_Jinkela_wire_6622)
    );

    bfr new_Jinkela_buffer_4993 (
        .din(new_Jinkela_wire_6452),
        .dout(new_Jinkela_wire_6453)
    );

    bfr new_Jinkela_buffer_5068 (
        .din(new_Jinkela_wire_6541),
        .dout(new_Jinkela_wire_6542)
    );

    bfr new_Jinkela_buffer_4994 (
        .din(new_Jinkela_wire_6453),
        .dout(new_Jinkela_wire_6454)
    );

    bfr new_Jinkela_buffer_5197 (
        .din(_1782_),
        .dout(new_Jinkela_wire_6679)
    );

    bfr new_Jinkela_buffer_4995 (
        .din(new_Jinkela_wire_6454),
        .dout(new_Jinkela_wire_6455)
    );

    bfr new_Jinkela_buffer_5069 (
        .din(new_Jinkela_wire_6542),
        .dout(new_Jinkela_wire_6543)
    );

    bfr new_Jinkela_buffer_4996 (
        .din(new_Jinkela_wire_6455),
        .dout(new_Jinkela_wire_6456)
    );

    bfr new_Jinkela_buffer_5145 (
        .din(new_Jinkela_wire_6622),
        .dout(new_Jinkela_wire_6623)
    );

    bfr new_Jinkela_buffer_4997 (
        .din(new_Jinkela_wire_6456),
        .dout(new_Jinkela_wire_6457)
    );

    bfr new_Jinkela_buffer_5070 (
        .din(new_Jinkela_wire_6543),
        .dout(new_Jinkela_wire_6544)
    );

    bfr new_Jinkela_buffer_4998 (
        .din(new_Jinkela_wire_6457),
        .dout(new_Jinkela_wire_6458)
    );

    spl2 new_Jinkela_splitter_591 (
        .a(_0646_),
        .b(new_Jinkela_wire_6682),
        .c(new_Jinkela_wire_6683)
    );

    spl2 new_Jinkela_splitter_592 (
        .a(_0570_),
        .b(new_Jinkela_wire_6685),
        .c(new_Jinkela_wire_6686)
    );

    bfr new_Jinkela_buffer_4999 (
        .din(new_Jinkela_wire_6458),
        .dout(new_Jinkela_wire_6459)
    );

    bfr new_Jinkela_buffer_5071 (
        .din(new_Jinkela_wire_6544),
        .dout(new_Jinkela_wire_6545)
    );

    bfr new_Jinkela_buffer_5000 (
        .din(new_Jinkela_wire_6459),
        .dout(new_Jinkela_wire_6460)
    );

    bfr new_Jinkela_buffer_5146 (
        .din(new_Jinkela_wire_6623),
        .dout(new_Jinkela_wire_6624)
    );

    bfr new_Jinkela_buffer_5001 (
        .din(new_Jinkela_wire_6460),
        .dout(new_Jinkela_wire_6461)
    );

    bfr new_Jinkela_buffer_5072 (
        .din(new_Jinkela_wire_6545),
        .dout(new_Jinkela_wire_6546)
    );

    bfr new_Jinkela_buffer_5002 (
        .din(new_Jinkela_wire_6461),
        .dout(new_Jinkela_wire_6462)
    );

    bfr new_Jinkela_buffer_5003 (
        .din(new_Jinkela_wire_6462),
        .dout(new_Jinkela_wire_6463)
    );

    bfr new_Jinkela_buffer_5073 (
        .din(new_Jinkela_wire_6546),
        .dout(new_Jinkela_wire_6547)
    );

    bfr new_Jinkela_buffer_5004 (
        .din(new_Jinkela_wire_6463),
        .dout(new_Jinkela_wire_6464)
    );

    bfr new_Jinkela_buffer_5147 (
        .din(new_Jinkela_wire_6624),
        .dout(new_Jinkela_wire_6625)
    );

    bfr new_Jinkela_buffer_5005 (
        .din(new_Jinkela_wire_6464),
        .dout(new_Jinkela_wire_6465)
    );

    bfr new_Jinkela_buffer_5074 (
        .din(new_Jinkela_wire_6547),
        .dout(new_Jinkela_wire_6548)
    );

    bfr new_Jinkela_buffer_5006 (
        .din(new_Jinkela_wire_6465),
        .dout(new_Jinkela_wire_6466)
    );

    bfr new_Jinkela_buffer_5198 (
        .din(_0151_),
        .dout(new_Jinkela_wire_6684)
    );

    bfr new_Jinkela_buffer_5007 (
        .din(new_Jinkela_wire_6466),
        .dout(new_Jinkela_wire_6467)
    );

    bfr new_Jinkela_buffer_8402 (
        .din(new_Jinkela_wire_10343),
        .dout(new_Jinkela_wire_10344)
    );

    bfr new_Jinkela_buffer_12065 (
        .din(new_Jinkela_wire_14542),
        .dout(new_Jinkela_wire_14543)
    );

    bfr new_Jinkela_buffer_8510 (
        .din(new_Jinkela_wire_10461),
        .dout(new_Jinkela_wire_10462)
    );

    bfr new_Jinkela_buffer_11878 (
        .din(new_Jinkela_wire_14349),
        .dout(new_Jinkela_wire_14350)
    );

    bfr new_Jinkela_buffer_8403 (
        .din(new_Jinkela_wire_10344),
        .dout(new_Jinkela_wire_10345)
    );

    bfr new_Jinkela_buffer_11965 (
        .din(new_Jinkela_wire_14438),
        .dout(new_Jinkela_wire_14439)
    );

    bfr new_Jinkela_buffer_8481 (
        .din(new_Jinkela_wire_10430),
        .dout(new_Jinkela_wire_10431)
    );

    bfr new_Jinkela_buffer_11879 (
        .din(new_Jinkela_wire_14350),
        .dout(new_Jinkela_wire_14351)
    );

    bfr new_Jinkela_buffer_8404 (
        .din(new_Jinkela_wire_10345),
        .dout(new_Jinkela_wire_10346)
    );

    bfr new_Jinkela_buffer_12103 (
        .din(new_Jinkela_wire_14580),
        .dout(new_Jinkela_wire_14581)
    );

    bfr new_Jinkela_buffer_8607 (
        .din(new_Jinkela_wire_10566),
        .dout(new_Jinkela_wire_10567)
    );

    bfr new_Jinkela_buffer_11880 (
        .din(new_Jinkela_wire_14351),
        .dout(new_Jinkela_wire_14352)
    );

    bfr new_Jinkela_buffer_8405 (
        .din(new_Jinkela_wire_10346),
        .dout(new_Jinkela_wire_10347)
    );

    bfr new_Jinkela_buffer_11966 (
        .din(new_Jinkela_wire_14439),
        .dout(new_Jinkela_wire_14440)
    );

    bfr new_Jinkela_buffer_8482 (
        .din(new_Jinkela_wire_10431),
        .dout(new_Jinkela_wire_10432)
    );

    bfr new_Jinkela_buffer_11881 (
        .din(new_Jinkela_wire_14352),
        .dout(new_Jinkela_wire_14353)
    );

    bfr new_Jinkela_buffer_8406 (
        .din(new_Jinkela_wire_10347),
        .dout(new_Jinkela_wire_10348)
    );

    bfr new_Jinkela_buffer_12069 (
        .din(new_Jinkela_wire_14546),
        .dout(new_Jinkela_wire_14547)
    );

    bfr new_Jinkela_buffer_8511 (
        .din(new_Jinkela_wire_10462),
        .dout(new_Jinkela_wire_10463)
    );

    bfr new_Jinkela_buffer_11882 (
        .din(new_Jinkela_wire_14353),
        .dout(new_Jinkela_wire_14354)
    );

    bfr new_Jinkela_buffer_8407 (
        .din(new_Jinkela_wire_10348),
        .dout(new_Jinkela_wire_10349)
    );

    bfr new_Jinkela_buffer_11967 (
        .din(new_Jinkela_wire_14440),
        .dout(new_Jinkela_wire_14441)
    );

    bfr new_Jinkela_buffer_8483 (
        .din(new_Jinkela_wire_10432),
        .dout(new_Jinkela_wire_10433)
    );

    bfr new_Jinkela_buffer_11883 (
        .din(new_Jinkela_wire_14354),
        .dout(new_Jinkela_wire_14355)
    );

    bfr new_Jinkela_buffer_8408 (
        .din(new_Jinkela_wire_10349),
        .dout(new_Jinkela_wire_10350)
    );

    bfr new_Jinkela_buffer_8609 (
        .din(new_Jinkela_wire_10570),
        .dout(new_Jinkela_wire_10571)
    );

    bfr new_Jinkela_buffer_11884 (
        .din(new_Jinkela_wire_14355),
        .dout(new_Jinkela_wire_14356)
    );

    bfr new_Jinkela_buffer_8409 (
        .din(new_Jinkela_wire_10350),
        .dout(new_Jinkela_wire_10351)
    );

    bfr new_Jinkela_buffer_11968 (
        .din(new_Jinkela_wire_14441),
        .dout(new_Jinkela_wire_14442)
    );

    bfr new_Jinkela_buffer_8484 (
        .din(new_Jinkela_wire_10433),
        .dout(new_Jinkela_wire_10434)
    );

    bfr new_Jinkela_buffer_11885 (
        .din(new_Jinkela_wire_14356),
        .dout(new_Jinkela_wire_14357)
    );

    bfr new_Jinkela_buffer_8410 (
        .din(new_Jinkela_wire_10351),
        .dout(new_Jinkela_wire_10352)
    );

    spl2 new_Jinkela_splitter_1090 (
        .a(_0400_),
        .b(new_Jinkela_wire_14660),
        .c(new_Jinkela_wire_14661)
    );

    bfr new_Jinkela_buffer_12070 (
        .din(new_Jinkela_wire_14547),
        .dout(new_Jinkela_wire_14548)
    );

    bfr new_Jinkela_buffer_8512 (
        .din(new_Jinkela_wire_10463),
        .dout(new_Jinkela_wire_10464)
    );

    bfr new_Jinkela_buffer_11886 (
        .din(new_Jinkela_wire_14357),
        .dout(new_Jinkela_wire_14358)
    );

    bfr new_Jinkela_buffer_8411 (
        .din(new_Jinkela_wire_10352),
        .dout(new_Jinkela_wire_10353)
    );

    bfr new_Jinkela_buffer_11969 (
        .din(new_Jinkela_wire_14442),
        .dout(new_Jinkela_wire_14443)
    );

    bfr new_Jinkela_buffer_8485 (
        .din(new_Jinkela_wire_10434),
        .dout(new_Jinkela_wire_10435)
    );

    bfr new_Jinkela_buffer_11887 (
        .din(new_Jinkela_wire_14358),
        .dout(new_Jinkela_wire_14359)
    );

    bfr new_Jinkela_buffer_8412 (
        .din(new_Jinkela_wire_10353),
        .dout(new_Jinkela_wire_10354)
    );

    bfr new_Jinkela_buffer_12104 (
        .din(new_Jinkela_wire_14581),
        .dout(new_Jinkela_wire_14582)
    );

    bfr new_Jinkela_buffer_11888 (
        .din(new_Jinkela_wire_14359),
        .dout(new_Jinkela_wire_14360)
    );

    spl2 new_Jinkela_splitter_832 (
        .a(_0608_),
        .b(new_Jinkela_wire_10614),
        .c(new_Jinkela_wire_10615)
    );

    bfr new_Jinkela_buffer_8413 (
        .din(new_Jinkela_wire_10354),
        .dout(new_Jinkela_wire_10355)
    );

    bfr new_Jinkela_buffer_11970 (
        .din(new_Jinkela_wire_14443),
        .dout(new_Jinkela_wire_14444)
    );

    bfr new_Jinkela_buffer_8486 (
        .din(new_Jinkela_wire_10435),
        .dout(new_Jinkela_wire_10436)
    );

    bfr new_Jinkela_buffer_11889 (
        .din(new_Jinkela_wire_14360),
        .dout(new_Jinkela_wire_14361)
    );

    bfr new_Jinkela_buffer_8414 (
        .din(new_Jinkela_wire_10355),
        .dout(new_Jinkela_wire_10356)
    );

    bfr new_Jinkela_buffer_12071 (
        .din(new_Jinkela_wire_14548),
        .dout(new_Jinkela_wire_14549)
    );

    bfr new_Jinkela_buffer_8513 (
        .din(new_Jinkela_wire_10464),
        .dout(new_Jinkela_wire_10465)
    );

    bfr new_Jinkela_buffer_11890 (
        .din(new_Jinkela_wire_14361),
        .dout(new_Jinkela_wire_14362)
    );

    bfr new_Jinkela_buffer_8415 (
        .din(new_Jinkela_wire_10356),
        .dout(new_Jinkela_wire_10357)
    );

    bfr new_Jinkela_buffer_11971 (
        .din(new_Jinkela_wire_14444),
        .dout(new_Jinkela_wire_14445)
    );

    bfr new_Jinkela_buffer_8487 (
        .din(new_Jinkela_wire_10436),
        .dout(new_Jinkela_wire_10437)
    );

    bfr new_Jinkela_buffer_11891 (
        .din(new_Jinkela_wire_14362),
        .dout(new_Jinkela_wire_14363)
    );

    bfr new_Jinkela_buffer_8416 (
        .din(new_Jinkela_wire_10357),
        .dout(new_Jinkela_wire_10358)
    );

    bfr new_Jinkela_buffer_8610 (
        .din(new_Jinkela_wire_10571),
        .dout(new_Jinkela_wire_10572)
    );

    bfr new_Jinkela_buffer_11892 (
        .din(new_Jinkela_wire_14363),
        .dout(new_Jinkela_wire_14364)
    );

    bfr new_Jinkela_buffer_8417 (
        .din(new_Jinkela_wire_10358),
        .dout(new_Jinkela_wire_10359)
    );

    bfr new_Jinkela_buffer_11972 (
        .din(new_Jinkela_wire_14445),
        .dout(new_Jinkela_wire_14446)
    );

    bfr new_Jinkela_buffer_8488 (
        .din(new_Jinkela_wire_10437),
        .dout(new_Jinkela_wire_10438)
    );

    bfr new_Jinkela_buffer_11893 (
        .din(new_Jinkela_wire_14364),
        .dout(new_Jinkela_wire_14365)
    );

    bfr new_Jinkela_buffer_8418 (
        .din(new_Jinkela_wire_10359),
        .dout(new_Jinkela_wire_10360)
    );

    bfr new_Jinkela_buffer_12072 (
        .din(new_Jinkela_wire_14549),
        .dout(new_Jinkela_wire_14550)
    );

    bfr new_Jinkela_buffer_8514 (
        .din(new_Jinkela_wire_10465),
        .dout(new_Jinkela_wire_10466)
    );

    bfr new_Jinkela_buffer_11894 (
        .din(new_Jinkela_wire_14365),
        .dout(new_Jinkela_wire_14366)
    );

    bfr new_Jinkela_buffer_8419 (
        .din(new_Jinkela_wire_10360),
        .dout(new_Jinkela_wire_10361)
    );

    bfr new_Jinkela_buffer_11973 (
        .din(new_Jinkela_wire_14446),
        .dout(new_Jinkela_wire_14447)
    );

    bfr new_Jinkela_buffer_8489 (
        .din(new_Jinkela_wire_10438),
        .dout(new_Jinkela_wire_10439)
    );

    bfr new_Jinkela_buffer_11895 (
        .din(new_Jinkela_wire_14366),
        .dout(new_Jinkela_wire_14367)
    );

    bfr new_Jinkela_buffer_8420 (
        .din(new_Jinkela_wire_10361),
        .dout(new_Jinkela_wire_10362)
    );

    bfr new_Jinkela_buffer_12105 (
        .din(new_Jinkela_wire_14582),
        .dout(new_Jinkela_wire_14583)
    );

    bfr new_Jinkela_buffer_11896 (
        .din(new_Jinkela_wire_14367),
        .dout(new_Jinkela_wire_14368)
    );

    bfr new_Jinkela_buffer_8648 (
        .din(_1125_),
        .dout(new_Jinkela_wire_10616)
    );

    bfr new_Jinkela_buffer_8421 (
        .din(new_Jinkela_wire_10362),
        .dout(new_Jinkela_wire_10363)
    );

    bfr new_Jinkela_buffer_11974 (
        .din(new_Jinkela_wire_14447),
        .dout(new_Jinkela_wire_14448)
    );

    bfr new_Jinkela_buffer_8490 (
        .din(new_Jinkela_wire_10439),
        .dout(new_Jinkela_wire_10440)
    );

    bfr new_Jinkela_buffer_11897 (
        .din(new_Jinkela_wire_14368),
        .dout(new_Jinkela_wire_14369)
    );

    bfr new_Jinkela_buffer_8422 (
        .din(new_Jinkela_wire_10363),
        .dout(new_Jinkela_wire_10364)
    );

    bfr new_Jinkela_buffer_12073 (
        .din(new_Jinkela_wire_14550),
        .dout(new_Jinkela_wire_14551)
    );

    bfr new_Jinkela_buffer_8515 (
        .din(new_Jinkela_wire_10466),
        .dout(new_Jinkela_wire_10467)
    );

    bfr new_Jinkela_buffer_11898 (
        .din(new_Jinkela_wire_14369),
        .dout(new_Jinkela_wire_14370)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_2348),
        .dout(new_Jinkela_wire_2349)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_2227),
        .dout(new_Jinkela_wire_2228)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_2295),
        .dout(new_Jinkela_wire_2296)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_2228),
        .dout(new_Jinkela_wire_2229)
    );

    spl2 new_Jinkela_splitter_291 (
        .a(_1175_),
        .b(new_Jinkela_wire_2458),
        .c(new_Jinkela_wire_2459)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(new_Jinkela_wire_2229),
        .dout(new_Jinkela_wire_2230)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_2296),
        .dout(new_Jinkela_wire_2297)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_2230),
        .dout(new_Jinkela_wire_2231)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(new_Jinkela_wire_2349),
        .dout(new_Jinkela_wire_2350)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_2231),
        .dout(new_Jinkela_wire_2232)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(new_Jinkela_wire_2297),
        .dout(new_Jinkela_wire_2298)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_2232),
        .dout(new_Jinkela_wire_2233)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(new_Jinkela_wire_2423),
        .dout(new_Jinkela_wire_2424)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_2233),
        .dout(new_Jinkela_wire_2234)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_2298),
        .dout(new_Jinkela_wire_2299)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_2234),
        .dout(new_Jinkela_wire_2235)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(new_Jinkela_wire_2350),
        .dout(new_Jinkela_wire_2351)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_2235),
        .dout(new_Jinkela_wire_2236)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_2299),
        .dout(new_Jinkela_wire_2300)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_2236),
        .dout(new_Jinkela_wire_2237)
    );

    spl2 new_Jinkela_splitter_292 (
        .a(_0575_),
        .b(new_Jinkela_wire_2460),
        .c(new_Jinkela_wire_2461)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_2237),
        .dout(new_Jinkela_wire_2238)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(new_Jinkela_wire_2300),
        .dout(new_Jinkela_wire_2301)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_2238),
        .dout(new_Jinkela_wire_2239)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(new_Jinkela_wire_2351),
        .dout(new_Jinkela_wire_2352)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_2239),
        .dout(new_Jinkela_wire_2240)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(new_Jinkela_wire_2301),
        .dout(new_Jinkela_wire_2302)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_2240),
        .dout(new_Jinkela_wire_2241)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_2424),
        .dout(new_Jinkela_wire_2425)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_2241),
        .dout(new_Jinkela_wire_2242)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(new_Jinkela_wire_2302),
        .dout(new_Jinkela_wire_2303)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(new_Jinkela_wire_2242),
        .dout(new_Jinkela_wire_2243)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_2352),
        .dout(new_Jinkela_wire_2353)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_2243),
        .dout(new_Jinkela_wire_2244)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(new_Jinkela_wire_2303),
        .dout(new_Jinkela_wire_2304)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_2244),
        .dout(new_Jinkela_wire_2245)
    );

    spl2 new_Jinkela_splitter_293 (
        .a(_1341_),
        .b(new_Jinkela_wire_2462),
        .c(new_Jinkela_wire_2463)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_2245),
        .dout(new_Jinkela_wire_2246)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_2304),
        .dout(new_Jinkela_wire_2305)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_2246),
        .dout(new_Jinkela_wire_2247)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_2353),
        .dout(new_Jinkela_wire_2354)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_2247),
        .dout(new_Jinkela_wire_2248)
    );

    bfr new_Jinkela_buffer_15377 (
        .din(new_Jinkela_wire_18331),
        .dout(new_Jinkela_wire_18332)
    );

    bfr new_Jinkela_buffer_8423 (
        .din(new_Jinkela_wire_10364),
        .dout(new_Jinkela_wire_10365)
    );

    bfr new_Jinkela_buffer_15427 (
        .din(new_Jinkela_wire_18391),
        .dout(new_Jinkela_wire_18392)
    );

    bfr new_Jinkela_buffer_8611 (
        .din(new_Jinkela_wire_10572),
        .dout(new_Jinkela_wire_10573)
    );

    bfr new_Jinkela_buffer_15378 (
        .din(new_Jinkela_wire_18332),
        .dout(new_Jinkela_wire_18333)
    );

    bfr new_Jinkela_buffer_8424 (
        .din(new_Jinkela_wire_10365),
        .dout(new_Jinkela_wire_10366)
    );

    spl2 new_Jinkela_splitter_1334 (
        .a(_0592_),
        .b(new_Jinkela_wire_18448),
        .c(new_Jinkela_wire_18449)
    );

    bfr new_Jinkela_buffer_8516 (
        .din(new_Jinkela_wire_10467),
        .dout(new_Jinkela_wire_10468)
    );

    spl2 new_Jinkela_splitter_1337 (
        .a(_0418_),
        .b(new_Jinkela_wire_18516),
        .c(new_Jinkela_wire_18517)
    );

    bfr new_Jinkela_buffer_15379 (
        .din(new_Jinkela_wire_18333),
        .dout(new_Jinkela_wire_18334)
    );

    bfr new_Jinkela_buffer_8425 (
        .din(new_Jinkela_wire_10366),
        .dout(new_Jinkela_wire_10367)
    );

    bfr new_Jinkela_buffer_15430 (
        .din(new_Jinkela_wire_18396),
        .dout(new_Jinkela_wire_18397)
    );

    bfr new_Jinkela_buffer_8613 (
        .din(new_Jinkela_wire_10576),
        .dout(new_Jinkela_wire_10577)
    );

    bfr new_Jinkela_buffer_15380 (
        .din(new_Jinkela_wire_18334),
        .dout(new_Jinkela_wire_18335)
    );

    bfr new_Jinkela_buffer_8426 (
        .din(new_Jinkela_wire_10367),
        .dout(new_Jinkela_wire_10368)
    );

    bfr new_Jinkela_buffer_8517 (
        .din(new_Jinkela_wire_10468),
        .dout(new_Jinkela_wire_10469)
    );

    bfr new_Jinkela_buffer_15381 (
        .din(new_Jinkela_wire_18335),
        .dout(new_Jinkela_wire_18336)
    );

    bfr new_Jinkela_buffer_8427 (
        .din(new_Jinkela_wire_10368),
        .dout(new_Jinkela_wire_10369)
    );

    bfr new_Jinkela_buffer_15431 (
        .din(new_Jinkela_wire_18397),
        .dout(new_Jinkela_wire_18398)
    );

    bfr new_Jinkela_buffer_8617 (
        .din(new_Jinkela_wire_10580),
        .dout(new_Jinkela_wire_10581)
    );

    bfr new_Jinkela_buffer_15382 (
        .din(new_Jinkela_wire_18336),
        .dout(new_Jinkela_wire_18337)
    );

    bfr new_Jinkela_buffer_8428 (
        .din(new_Jinkela_wire_10369),
        .dout(new_Jinkela_wire_10370)
    );

    bfr new_Jinkela_buffer_8518 (
        .din(new_Jinkela_wire_10469),
        .dout(new_Jinkela_wire_10470)
    );

    bfr new_Jinkela_buffer_15477 (
        .din(_0547_),
        .dout(new_Jinkela_wire_18450)
    );

    bfr new_Jinkela_buffer_15383 (
        .din(new_Jinkela_wire_18337),
        .dout(new_Jinkela_wire_18338)
    );

    bfr new_Jinkela_buffer_8429 (
        .din(new_Jinkela_wire_10370),
        .dout(new_Jinkela_wire_10371)
    );

    bfr new_Jinkela_buffer_15432 (
        .din(new_Jinkela_wire_18398),
        .dout(new_Jinkela_wire_18399)
    );

    bfr new_Jinkela_buffer_8614 (
        .din(new_Jinkela_wire_10577),
        .dout(new_Jinkela_wire_10578)
    );

    bfr new_Jinkela_buffer_15384 (
        .din(new_Jinkela_wire_18338),
        .dout(new_Jinkela_wire_18339)
    );

    bfr new_Jinkela_buffer_8430 (
        .din(new_Jinkela_wire_10371),
        .dout(new_Jinkela_wire_10372)
    );

    bfr new_Jinkela_buffer_8519 (
        .din(new_Jinkela_wire_10470),
        .dout(new_Jinkela_wire_10471)
    );

    bfr new_Jinkela_buffer_15519 (
        .din(_0691_),
        .dout(new_Jinkela_wire_18494)
    );

    bfr new_Jinkela_buffer_15385 (
        .din(new_Jinkela_wire_18339),
        .dout(new_Jinkela_wire_18340)
    );

    bfr new_Jinkela_buffer_8431 (
        .din(new_Jinkela_wire_10372),
        .dout(new_Jinkela_wire_10373)
    );

    bfr new_Jinkela_buffer_15433 (
        .din(new_Jinkela_wire_18399),
        .dout(new_Jinkela_wire_18400)
    );

    spl2 new_Jinkela_splitter_834 (
        .a(_0459_),
        .b(new_Jinkela_wire_10675),
        .c(new_Jinkela_wire_10676)
    );

    bfr new_Jinkela_buffer_15386 (
        .din(new_Jinkela_wire_18340),
        .dout(new_Jinkela_wire_18341)
    );

    bfr new_Jinkela_buffer_8432 (
        .din(new_Jinkela_wire_10373),
        .dout(new_Jinkela_wire_10374)
    );

    bfr new_Jinkela_buffer_15478 (
        .din(new_Jinkela_wire_18450),
        .dout(new_Jinkela_wire_18451)
    );

    bfr new_Jinkela_buffer_8520 (
        .din(new_Jinkela_wire_10471),
        .dout(new_Jinkela_wire_10472)
    );

    bfr new_Jinkela_buffer_15387 (
        .din(new_Jinkela_wire_18341),
        .dout(new_Jinkela_wire_18342)
    );

    bfr new_Jinkela_buffer_8433 (
        .din(new_Jinkela_wire_10374),
        .dout(new_Jinkela_wire_10375)
    );

    bfr new_Jinkela_buffer_15434 (
        .din(new_Jinkela_wire_18400),
        .dout(new_Jinkela_wire_18401)
    );

    bfr new_Jinkela_buffer_8615 (
        .din(new_Jinkela_wire_10578),
        .dout(new_Jinkela_wire_10579)
    );

    bfr new_Jinkela_buffer_15388 (
        .din(new_Jinkela_wire_18342),
        .dout(new_Jinkela_wire_18343)
    );

    bfr new_Jinkela_buffer_8434 (
        .din(new_Jinkela_wire_10375),
        .dout(new_Jinkela_wire_10376)
    );

    bfr new_Jinkela_buffer_8521 (
        .din(new_Jinkela_wire_10472),
        .dout(new_Jinkela_wire_10473)
    );

    bfr new_Jinkela_buffer_15543 (
        .din(_1591_),
        .dout(new_Jinkela_wire_18522)
    );

    bfr new_Jinkela_buffer_15389 (
        .din(new_Jinkela_wire_18343),
        .dout(new_Jinkela_wire_18344)
    );

    bfr new_Jinkela_buffer_8435 (
        .din(new_Jinkela_wire_10376),
        .dout(new_Jinkela_wire_10377)
    );

    bfr new_Jinkela_buffer_15435 (
        .din(new_Jinkela_wire_18401),
        .dout(new_Jinkela_wire_18402)
    );

    bfr new_Jinkela_buffer_8618 (
        .din(new_Jinkela_wire_10581),
        .dout(new_Jinkela_wire_10582)
    );

    bfr new_Jinkela_buffer_15390 (
        .din(new_Jinkela_wire_18344),
        .dout(new_Jinkela_wire_18345)
    );

    bfr new_Jinkela_buffer_8436 (
        .din(new_Jinkela_wire_10377),
        .dout(new_Jinkela_wire_10378)
    );

    bfr new_Jinkela_buffer_15479 (
        .din(new_Jinkela_wire_18451),
        .dout(new_Jinkela_wire_18452)
    );

    bfr new_Jinkela_buffer_8522 (
        .din(new_Jinkela_wire_10473),
        .dout(new_Jinkela_wire_10474)
    );

    bfr new_Jinkela_buffer_15391 (
        .din(new_Jinkela_wire_18345),
        .dout(new_Jinkela_wire_18346)
    );

    bfr new_Jinkela_buffer_8437 (
        .din(new_Jinkela_wire_10378),
        .dout(new_Jinkela_wire_10379)
    );

    bfr new_Jinkela_buffer_15436 (
        .din(new_Jinkela_wire_18402),
        .dout(new_Jinkela_wire_18403)
    );

    bfr new_Jinkela_buffer_8704 (
        .din(_0260_),
        .dout(new_Jinkela_wire_10674)
    );

    bfr new_Jinkela_buffer_15392 (
        .din(new_Jinkela_wire_18346),
        .dout(new_Jinkela_wire_18347)
    );

    bfr new_Jinkela_buffer_8438 (
        .din(new_Jinkela_wire_10379),
        .dout(new_Jinkela_wire_10380)
    );

    bfr new_Jinkela_buffer_15520 (
        .din(new_Jinkela_wire_18494),
        .dout(new_Jinkela_wire_18495)
    );

    bfr new_Jinkela_buffer_8523 (
        .din(new_Jinkela_wire_10474),
        .dout(new_Jinkela_wire_10475)
    );

    bfr new_Jinkela_buffer_15393 (
        .din(new_Jinkela_wire_18347),
        .dout(new_Jinkela_wire_18348)
    );

    bfr new_Jinkela_buffer_8439 (
        .din(new_Jinkela_wire_10380),
        .dout(new_Jinkela_wire_10381)
    );

    bfr new_Jinkela_buffer_15437 (
        .din(new_Jinkela_wire_18403),
        .dout(new_Jinkela_wire_18404)
    );

    bfr new_Jinkela_buffer_8619 (
        .din(new_Jinkela_wire_10582),
        .dout(new_Jinkela_wire_10583)
    );

    bfr new_Jinkela_buffer_15394 (
        .din(new_Jinkela_wire_18348),
        .dout(new_Jinkela_wire_18349)
    );

    bfr new_Jinkela_buffer_8440 (
        .din(new_Jinkela_wire_10381),
        .dout(new_Jinkela_wire_10382)
    );

    bfr new_Jinkela_buffer_15480 (
        .din(new_Jinkela_wire_18452),
        .dout(new_Jinkela_wire_18453)
    );

    bfr new_Jinkela_buffer_8524 (
        .din(new_Jinkela_wire_10475),
        .dout(new_Jinkela_wire_10476)
    );

    bfr new_Jinkela_buffer_15395 (
        .din(new_Jinkela_wire_18349),
        .dout(new_Jinkela_wire_18350)
    );

    bfr new_Jinkela_buffer_8441 (
        .din(new_Jinkela_wire_10382),
        .dout(new_Jinkela_wire_10383)
    );

    bfr new_Jinkela_buffer_15438 (
        .din(new_Jinkela_wire_18404),
        .dout(new_Jinkela_wire_18405)
    );

    bfr new_Jinkela_buffer_8649 (
        .din(new_Jinkela_wire_10616),
        .dout(new_Jinkela_wire_10617)
    );

    bfr new_Jinkela_buffer_15396 (
        .din(new_Jinkela_wire_18350),
        .dout(new_Jinkela_wire_18351)
    );

    bfr new_Jinkela_buffer_8442 (
        .din(new_Jinkela_wire_10383),
        .dout(new_Jinkela_wire_10384)
    );

    bfr new_Jinkela_buffer_8525 (
        .din(new_Jinkela_wire_10476),
        .dout(new_Jinkela_wire_10477)
    );

    bfr new_Jinkela_buffer_15539 (
        .din(new_Jinkela_wire_18517),
        .dout(new_Jinkela_wire_18518)
    );

    bfr new_Jinkela_buffer_15397 (
        .din(new_Jinkela_wire_18351),
        .dout(new_Jinkela_wire_18352)
    );

    bfr new_Jinkela_buffer_8443 (
        .din(new_Jinkela_wire_10384),
        .dout(new_Jinkela_wire_10385)
    );

    bfr new_Jinkela_buffer_15439 (
        .din(new_Jinkela_wire_18405),
        .dout(new_Jinkela_wire_18406)
    );

    bfr new_Jinkela_buffer_8620 (
        .din(new_Jinkela_wire_10583),
        .dout(new_Jinkela_wire_10584)
    );

    bfr new_Jinkela_buffer_11975 (
        .din(new_Jinkela_wire_14448),
        .dout(new_Jinkela_wire_14449)
    );

    and_bb _2581_ (
        .a(new_Jinkela_wire_11455),
        .b(new_Jinkela_wire_12220),
        .c(_1630_)
    );

    bfr new_Jinkela_buffer_11899 (
        .din(new_Jinkela_wire_14370),
        .dout(new_Jinkela_wire_14371)
    );

    or_bb _2582_ (
        .a(new_Jinkela_wire_7741),
        .b(new_Jinkela_wire_11724),
        .c(_1631_)
    );

    or_bb _2583_ (
        .a(new_Jinkela_wire_21192),
        .b(new_Jinkela_wire_3184),
        .c(_1633_)
    );

    bfr new_Jinkela_buffer_11900 (
        .din(new_Jinkela_wire_14371),
        .dout(new_Jinkela_wire_14372)
    );

    or_ii _2584_ (
        .a(new_Jinkela_wire_21193),
        .b(new_Jinkela_wire_3185),
        .c(_1634_)
    );

    bfr new_Jinkela_buffer_11976 (
        .din(new_Jinkela_wire_14449),
        .dout(new_Jinkela_wire_14450)
    );

    or_ii _2585_ (
        .a(new_Jinkela_wire_3257),
        .b(new_Jinkela_wire_17662),
        .c(_1635_)
    );

    bfr new_Jinkela_buffer_11901 (
        .din(new_Jinkela_wire_14372),
        .dout(new_Jinkela_wire_14373)
    );

    and_ii _2586_ (
        .a(new_Jinkela_wire_18950),
        .b(new_Jinkela_wire_3178),
        .c(_1636_)
    );

    bfr new_Jinkela_buffer_12178 (
        .din(_1497_),
        .dout(new_Jinkela_wire_14662)
    );

    and_bb _2587_ (
        .a(new_Jinkela_wire_18951),
        .b(new_Jinkela_wire_3179),
        .c(_1637_)
    );

    bfr new_Jinkela_buffer_12074 (
        .din(new_Jinkela_wire_14551),
        .dout(new_Jinkela_wire_14552)
    );

    bfr new_Jinkela_buffer_11902 (
        .din(new_Jinkela_wire_14373),
        .dout(new_Jinkela_wire_14374)
    );

    or_bb _2588_ (
        .a(new_Jinkela_wire_11341),
        .b(new_Jinkela_wire_1138),
        .c(_1638_)
    );

    bfr new_Jinkela_buffer_11977 (
        .din(new_Jinkela_wire_14450),
        .dout(new_Jinkela_wire_14451)
    );

    or_bb _2589_ (
        .a(new_Jinkela_wire_17977),
        .b(new_Jinkela_wire_3191),
        .c(_1639_)
    );

    bfr new_Jinkela_buffer_11903 (
        .din(new_Jinkela_wire_14374),
        .dout(new_Jinkela_wire_14375)
    );

    or_ii _2590_ (
        .a(new_Jinkela_wire_17978),
        .b(new_Jinkela_wire_3192),
        .c(_1640_)
    );

    or_ii _2591_ (
        .a(new_Jinkela_wire_2957),
        .b(new_Jinkela_wire_13207),
        .c(_1641_)
    );

    bfr new_Jinkela_buffer_12106 (
        .din(new_Jinkela_wire_14583),
        .dout(new_Jinkela_wire_14584)
    );

    bfr new_Jinkela_buffer_11904 (
        .din(new_Jinkela_wire_14375),
        .dout(new_Jinkela_wire_14376)
    );

    and_ii _2592_ (
        .a(new_Jinkela_wire_16777),
        .b(new_Jinkela_wire_16864),
        .c(_1642_)
    );

    bfr new_Jinkela_buffer_11978 (
        .din(new_Jinkela_wire_14451),
        .dout(new_Jinkela_wire_14452)
    );

    and_bb _2593_ (
        .a(new_Jinkela_wire_16778),
        .b(new_Jinkela_wire_16865),
        .c(_1644_)
    );

    bfr new_Jinkela_buffer_11905 (
        .din(new_Jinkela_wire_14376),
        .dout(new_Jinkela_wire_14377)
    );

    or_bb _2594_ (
        .a(new_Jinkela_wire_6959),
        .b(new_Jinkela_wire_13967),
        .c(_1645_)
    );

    or_bb _2595_ (
        .a(new_Jinkela_wire_6676),
        .b(new_Jinkela_wire_1584),
        .c(_1646_)
    );

    bfr new_Jinkela_buffer_12075 (
        .din(new_Jinkela_wire_14552),
        .dout(new_Jinkela_wire_14553)
    );

    bfr new_Jinkela_buffer_11906 (
        .din(new_Jinkela_wire_14377),
        .dout(new_Jinkela_wire_14378)
    );

    or_ii _2596_ (
        .a(new_Jinkela_wire_6677),
        .b(new_Jinkela_wire_1585),
        .c(_1647_)
    );

    bfr new_Jinkela_buffer_11979 (
        .din(new_Jinkela_wire_14452),
        .dout(new_Jinkela_wire_14453)
    );

    or_ii _2597_ (
        .a(new_Jinkela_wire_19080),
        .b(new_Jinkela_wire_13381),
        .c(_1648_)
    );

    bfr new_Jinkela_buffer_11907 (
        .din(new_Jinkela_wire_14378),
        .dout(new_Jinkela_wire_14379)
    );

    and_ii _2598_ (
        .a(new_Jinkela_wire_5418),
        .b(new_Jinkela_wire_19466),
        .c(_1649_)
    );

    and_bb _2599_ (
        .a(new_Jinkela_wire_5419),
        .b(new_Jinkela_wire_19467),
        .c(_1650_)
    );

    bfr new_Jinkela_buffer_11908 (
        .din(new_Jinkela_wire_14379),
        .dout(new_Jinkela_wire_14380)
    );

    or_bb _2600_ (
        .a(new_Jinkela_wire_11954),
        .b(new_Jinkela_wire_2598),
        .c(_1651_)
    );

    bfr new_Jinkela_buffer_11980 (
        .din(new_Jinkela_wire_14453),
        .dout(new_Jinkela_wire_14454)
    );

    or_bb _2601_ (
        .a(new_Jinkela_wire_20039),
        .b(new_Jinkela_wire_3713),
        .c(_1652_)
    );

    bfr new_Jinkela_buffer_11909 (
        .din(new_Jinkela_wire_14380),
        .dout(new_Jinkela_wire_14381)
    );

    or_ii _2602_ (
        .a(new_Jinkela_wire_20040),
        .b(new_Jinkela_wire_3714),
        .c(_1653_)
    );

    bfr new_Jinkela_buffer_12179 (
        .din(_1217_),
        .dout(new_Jinkela_wire_14665)
    );

    or_ii _2603_ (
        .a(new_Jinkela_wire_7835),
        .b(new_Jinkela_wire_16909),
        .c(_1655_)
    );

    bfr new_Jinkela_buffer_12076 (
        .din(new_Jinkela_wire_14553),
        .dout(new_Jinkela_wire_14554)
    );

    bfr new_Jinkela_buffer_11910 (
        .din(new_Jinkela_wire_14381),
        .dout(new_Jinkela_wire_14382)
    );

    and_ii _2604_ (
        .a(new_Jinkela_wire_14098),
        .b(new_Jinkela_wire_10833),
        .c(_1656_)
    );

    bfr new_Jinkela_buffer_11981 (
        .din(new_Jinkela_wire_14454),
        .dout(new_Jinkela_wire_14455)
    );

    and_bb _2605_ (
        .a(new_Jinkela_wire_14099),
        .b(new_Jinkela_wire_10834),
        .c(_1657_)
    );

    bfr new_Jinkela_buffer_11911 (
        .din(new_Jinkela_wire_14382),
        .dout(new_Jinkela_wire_14383)
    );

    or_bb _2606_ (
        .a(new_Jinkela_wire_10101),
        .b(new_Jinkela_wire_12341),
        .c(_1658_)
    );

    or_bb _2607_ (
        .a(new_Jinkela_wire_11957),
        .b(new_Jinkela_wire_17011),
        .c(_1659_)
    );

    bfr new_Jinkela_buffer_12107 (
        .din(new_Jinkela_wire_14584),
        .dout(new_Jinkela_wire_14585)
    );

    bfr new_Jinkela_buffer_11912 (
        .din(new_Jinkela_wire_14383),
        .dout(new_Jinkela_wire_14384)
    );

    or_ii _2608_ (
        .a(new_Jinkela_wire_11958),
        .b(new_Jinkela_wire_17012),
        .c(_1660_)
    );

    bfr new_Jinkela_buffer_11982 (
        .din(new_Jinkela_wire_14455),
        .dout(new_Jinkela_wire_14456)
    );

    or_ii _2609_ (
        .a(new_Jinkela_wire_20348),
        .b(new_Jinkela_wire_12045),
        .c(_1661_)
    );

    bfr new_Jinkela_buffer_11913 (
        .din(new_Jinkela_wire_14384),
        .dout(new_Jinkela_wire_14385)
    );

    and_ii _2610_ (
        .a(new_Jinkela_wire_5540),
        .b(new_Jinkela_wire_11226),
        .c(_1662_)
    );

    and_bb _2611_ (
        .a(new_Jinkela_wire_5541),
        .b(new_Jinkela_wire_11227),
        .c(_1663_)
    );

    bfr new_Jinkela_buffer_12077 (
        .din(new_Jinkela_wire_14554),
        .dout(new_Jinkela_wire_14555)
    );

    bfr new_Jinkela_buffer_11914 (
        .din(new_Jinkela_wire_14385),
        .dout(new_Jinkela_wire_14386)
    );

    or_bb _2612_ (
        .a(new_Jinkela_wire_13348),
        .b(new_Jinkela_wire_2143),
        .c(_1664_)
    );

    bfr new_Jinkela_buffer_11983 (
        .din(new_Jinkela_wire_14456),
        .dout(new_Jinkela_wire_14457)
    );

    or_bb _2613_ (
        .a(new_Jinkela_wire_1389),
        .b(new_Jinkela_wire_17053),
        .c(_1666_)
    );

    bfr new_Jinkela_buffer_11915 (
        .din(new_Jinkela_wire_14386),
        .dout(new_Jinkela_wire_14387)
    );

    or_ii _2614_ (
        .a(new_Jinkela_wire_1390),
        .b(new_Jinkela_wire_17054),
        .c(_1667_)
    );

    or_ii _2615_ (
        .a(new_Jinkela_wire_16369),
        .b(new_Jinkela_wire_708),
        .c(_1668_)
    );

    spl2 new_Jinkela_splitter_1091 (
        .a(_1214_),
        .b(new_Jinkela_wire_14663),
        .c(new_Jinkela_wire_14664)
    );

    bfr new_Jinkela_buffer_11916 (
        .din(new_Jinkela_wire_14387),
        .dout(new_Jinkela_wire_14388)
    );

    and_ii _2616_ (
        .a(new_Jinkela_wire_1912),
        .b(new_Jinkela_wire_13003),
        .c(_1669_)
    );

    bfr new_Jinkela_buffer_11984 (
        .din(new_Jinkela_wire_14457),
        .dout(new_Jinkela_wire_14458)
    );

    and_bb _2617_ (
        .a(new_Jinkela_wire_1913),
        .b(new_Jinkela_wire_13004),
        .c(_1670_)
    );

    bfr new_Jinkela_buffer_11917 (
        .din(new_Jinkela_wire_14388),
        .dout(new_Jinkela_wire_14389)
    );

    or_bb _2618_ (
        .a(new_Jinkela_wire_7505),
        .b(new_Jinkela_wire_17359),
        .c(_1671_)
    );

    or_bb _2619_ (
        .a(new_Jinkela_wire_6419),
        .b(new_Jinkela_wire_17795),
        .c(_1672_)
    );

    bfr new_Jinkela_buffer_12078 (
        .din(new_Jinkela_wire_14555),
        .dout(new_Jinkela_wire_14556)
    );

    bfr new_Jinkela_buffer_11918 (
        .din(new_Jinkela_wire_14389),
        .dout(new_Jinkela_wire_14390)
    );

    and_bb _2620_ (
        .a(new_Jinkela_wire_6420),
        .b(new_Jinkela_wire_17796),
        .c(_1673_)
    );

    bfr new_Jinkela_buffer_11985 (
        .din(new_Jinkela_wire_14458),
        .dout(new_Jinkela_wire_14459)
    );

    or_bi _2621_ (
        .a(new_Jinkela_wire_4997),
        .b(new_Jinkela_wire_5092),
        .c(_1674_)
    );

    bfr new_Jinkela_buffer_11919 (
        .din(new_Jinkela_wire_14390),
        .dout(new_Jinkela_wire_14391)
    );

    and_ii _2622_ (
        .a(new_Jinkela_wire_10973),
        .b(new_Jinkela_wire_3661),
        .c(_1675_)
    );

    bfr new_Jinkela_buffer_15398 (
        .din(new_Jinkela_wire_18352),
        .dout(new_Jinkela_wire_18353)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(new_Jinkela_wire_2305),
        .dout(new_Jinkela_wire_2306)
    );

    bfr new_Jinkela_buffer_15481 (
        .din(new_Jinkela_wire_18453),
        .dout(new_Jinkela_wire_18454)
    );

    spl2 new_Jinkela_splitter_275 (
        .a(new_Jinkela_wire_2248),
        .b(new_Jinkela_wire_2249),
        .c(new_Jinkela_wire_2250)
    );

    bfr new_Jinkela_buffer_15399 (
        .din(new_Jinkela_wire_18353),
        .dout(new_Jinkela_wire_18354)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_2306),
        .dout(new_Jinkela_wire_2307)
    );

    bfr new_Jinkela_buffer_15440 (
        .din(new_Jinkela_wire_18406),
        .dout(new_Jinkela_wire_18407)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_Jinkela_wire_2425),
        .dout(new_Jinkela_wire_2426)
    );

    bfr new_Jinkela_buffer_15400 (
        .din(new_Jinkela_wire_18354),
        .dout(new_Jinkela_wire_18355)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_2354),
        .dout(new_Jinkela_wire_2355)
    );

    bfr new_Jinkela_buffer_15521 (
        .din(new_Jinkela_wire_18495),
        .dout(new_Jinkela_wire_18496)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_Jinkela_wire_2307),
        .dout(new_Jinkela_wire_2308)
    );

    bfr new_Jinkela_buffer_15401 (
        .din(new_Jinkela_wire_18355),
        .dout(new_Jinkela_wire_18356)
    );

    bfr new_Jinkela_buffer_15441 (
        .din(new_Jinkela_wire_18407),
        .dout(new_Jinkela_wire_18408)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_2308),
        .dout(new_Jinkela_wire_2309)
    );

    bfr new_Jinkela_buffer_15402 (
        .din(new_Jinkela_wire_18356),
        .dout(new_Jinkela_wire_18357)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(new_Jinkela_wire_2355),
        .dout(new_Jinkela_wire_2356)
    );

    bfr new_Jinkela_buffer_15482 (
        .din(new_Jinkela_wire_18454),
        .dout(new_Jinkela_wire_18455)
    );

    spl2 new_Jinkela_splitter_279 (
        .a(new_Jinkela_wire_2309),
        .b(new_Jinkela_wire_2310),
        .c(new_Jinkela_wire_2311)
    );

    bfr new_Jinkela_buffer_15403 (
        .din(new_Jinkela_wire_18357),
        .dout(new_Jinkela_wire_18358)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(new_Jinkela_wire_2356),
        .dout(new_Jinkela_wire_2357)
    );

    bfr new_Jinkela_buffer_15442 (
        .din(new_Jinkela_wire_18408),
        .dout(new_Jinkela_wire_18409)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(new_Jinkela_wire_2426),
        .dout(new_Jinkela_wire_2427)
    );

    bfr new_Jinkela_buffer_15404 (
        .din(new_Jinkela_wire_18358),
        .dout(new_Jinkela_wire_18359)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(_0604_),
        .dout(new_Jinkela_wire_2464)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_2357),
        .dout(new_Jinkela_wire_2358)
    );

    spl2 new_Jinkela_splitter_1338 (
        .a(_1297_),
        .b(new_Jinkela_wire_18523),
        .c(new_Jinkela_wire_18524)
    );

    bfr new_Jinkela_buffer_15405 (
        .din(new_Jinkela_wire_18359),
        .dout(new_Jinkela_wire_18360)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_2427),
        .dout(new_Jinkela_wire_2428)
    );

    bfr new_Jinkela_buffer_15443 (
        .din(new_Jinkela_wire_18409),
        .dout(new_Jinkela_wire_18410)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(new_Jinkela_wire_2358),
        .dout(new_Jinkela_wire_2359)
    );

    bfr new_Jinkela_buffer_15406 (
        .din(new_Jinkela_wire_18360),
        .dout(new_Jinkela_wire_18361)
    );

    spl2 new_Jinkela_splitter_295 (
        .a(_0527_),
        .b(new_Jinkela_wire_2481),
        .c(new_Jinkela_wire_2482)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(_0237_),
        .dout(new_Jinkela_wire_2465)
    );

    bfr new_Jinkela_buffer_15483 (
        .din(new_Jinkela_wire_18455),
        .dout(new_Jinkela_wire_18456)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(new_Jinkela_wire_2359),
        .dout(new_Jinkela_wire_2360)
    );

    bfr new_Jinkela_buffer_15407 (
        .din(new_Jinkela_wire_18361),
        .dout(new_Jinkela_wire_18362)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_2428),
        .dout(new_Jinkela_wire_2429)
    );

    bfr new_Jinkela_buffer_15444 (
        .din(new_Jinkela_wire_18410),
        .dout(new_Jinkela_wire_18411)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(new_Jinkela_wire_2360),
        .dout(new_Jinkela_wire_2361)
    );

    bfr new_Jinkela_buffer_15408 (
        .din(new_Jinkela_wire_18362),
        .dout(new_Jinkela_wire_18363)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(_1336_),
        .dout(new_Jinkela_wire_2483)
    );

    bfr new_Jinkela_buffer_15522 (
        .din(new_Jinkela_wire_18496),
        .dout(new_Jinkela_wire_18497)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_2361),
        .dout(new_Jinkela_wire_2362)
    );

    bfr new_Jinkela_buffer_15409 (
        .din(new_Jinkela_wire_18363),
        .dout(new_Jinkela_wire_18364)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_2429),
        .dout(new_Jinkela_wire_2430)
    );

    bfr new_Jinkela_buffer_15445 (
        .din(new_Jinkela_wire_18411),
        .dout(new_Jinkela_wire_18412)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(new_Jinkela_wire_2362),
        .dout(new_Jinkela_wire_2363)
    );

    bfr new_Jinkela_buffer_15410 (
        .din(new_Jinkela_wire_18364),
        .dout(new_Jinkela_wire_18365)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(new_Jinkela_wire_2465),
        .dout(new_Jinkela_wire_2466)
    );

    bfr new_Jinkela_buffer_15484 (
        .din(new_Jinkela_wire_18456),
        .dout(new_Jinkela_wire_18457)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(new_Jinkela_wire_2363),
        .dout(new_Jinkela_wire_2364)
    );

    bfr new_Jinkela_buffer_15411 (
        .din(new_Jinkela_wire_18365),
        .dout(new_Jinkela_wire_18366)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_2430),
        .dout(new_Jinkela_wire_2431)
    );

    bfr new_Jinkela_buffer_15446 (
        .din(new_Jinkela_wire_18412),
        .dout(new_Jinkela_wire_18413)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(new_Jinkela_wire_2364),
        .dout(new_Jinkela_wire_2365)
    );

    bfr new_Jinkela_buffer_15412 (
        .din(new_Jinkela_wire_18366),
        .dout(new_Jinkela_wire_18367)
    );

    spl2 new_Jinkela_splitter_296 (
        .a(_1681_),
        .b(new_Jinkela_wire_2485),
        .c(new_Jinkela_wire_2486)
    );

    bfr new_Jinkela_buffer_15544 (
        .din(_0845_),
        .dout(new_Jinkela_wire_18525)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(new_Jinkela_wire_2365),
        .dout(new_Jinkela_wire_2366)
    );

    bfr new_Jinkela_buffer_15413 (
        .din(new_Jinkela_wire_18367),
        .dout(new_Jinkela_wire_18368)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_2431),
        .dout(new_Jinkela_wire_2432)
    );

    bfr new_Jinkela_buffer_15447 (
        .din(new_Jinkela_wire_18413),
        .dout(new_Jinkela_wire_18414)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_2366),
        .dout(new_Jinkela_wire_2367)
    );

    bfr new_Jinkela_buffer_15414 (
        .din(new_Jinkela_wire_18368),
        .dout(new_Jinkela_wire_18369)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(new_Jinkela_wire_2466),
        .dout(new_Jinkela_wire_2467)
    );

    bfr new_Jinkela_buffer_15485 (
        .din(new_Jinkela_wire_18457),
        .dout(new_Jinkela_wire_18458)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(new_Jinkela_wire_2367),
        .dout(new_Jinkela_wire_2368)
    );

    bfr new_Jinkela_buffer_15415 (
        .din(new_Jinkela_wire_18369),
        .dout(new_Jinkela_wire_18370)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_2432),
        .dout(new_Jinkela_wire_2433)
    );

    bfr new_Jinkela_buffer_15448 (
        .din(new_Jinkela_wire_18414),
        .dout(new_Jinkela_wire_18415)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_2368),
        .dout(new_Jinkela_wire_2369)
    );

    bfr new_Jinkela_buffer_15416 (
        .din(new_Jinkela_wire_18370),
        .dout(new_Jinkela_wire_18371)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(_0875_),
        .dout(new_Jinkela_wire_2484)
    );

    bfr new_Jinkela_buffer_15523 (
        .din(new_Jinkela_wire_18497),
        .dout(new_Jinkela_wire_18498)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_2369),
        .dout(new_Jinkela_wire_2370)
    );

    bfr new_Jinkela_buffer_15417 (
        .din(new_Jinkela_wire_18371),
        .dout(new_Jinkela_wire_18372)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_2433),
        .dout(new_Jinkela_wire_2434)
    );

    bfr new_Jinkela_buffer_15449 (
        .din(new_Jinkela_wire_18415),
        .dout(new_Jinkela_wire_18416)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(new_Jinkela_wire_2370),
        .dout(new_Jinkela_wire_2371)
    );

    spl2 new_Jinkela_splitter_1326 (
        .a(new_Jinkela_wire_18372),
        .b(new_Jinkela_wire_18373),
        .c(new_Jinkela_wire_18374)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(new_Jinkela_wire_2467),
        .dout(new_Jinkela_wire_2468)
    );

    bfr new_Jinkela_buffer_15486 (
        .din(new_Jinkela_wire_18458),
        .dout(new_Jinkela_wire_18459)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(new_Jinkela_wire_2371),
        .dout(new_Jinkela_wire_2372)
    );

    bfr new_Jinkela_buffer_12108 (
        .din(new_Jinkela_wire_14585),
        .dout(new_Jinkela_wire_14586)
    );

    bfr new_Jinkela_buffer_11920 (
        .din(new_Jinkela_wire_14391),
        .dout(new_Jinkela_wire_14392)
    );

    bfr new_Jinkela_buffer_11986 (
        .din(new_Jinkela_wire_14459),
        .dout(new_Jinkela_wire_14460)
    );

    bfr new_Jinkela_buffer_11921 (
        .din(new_Jinkela_wire_14392),
        .dout(new_Jinkela_wire_14393)
    );

    bfr new_Jinkela_buffer_12079 (
        .din(new_Jinkela_wire_14556),
        .dout(new_Jinkela_wire_14557)
    );

    bfr new_Jinkela_buffer_11922 (
        .din(new_Jinkela_wire_14393),
        .dout(new_Jinkela_wire_14394)
    );

    bfr new_Jinkela_buffer_11987 (
        .din(new_Jinkela_wire_14460),
        .dout(new_Jinkela_wire_14461)
    );

    bfr new_Jinkela_buffer_11923 (
        .din(new_Jinkela_wire_14394),
        .dout(new_Jinkela_wire_14395)
    );

    spl2 new_Jinkela_splitter_1094 (
        .a(_0368_),
        .b(new_Jinkela_wire_14685),
        .c(new_Jinkela_wire_14686)
    );

    bfr new_Jinkela_buffer_11924 (
        .din(new_Jinkela_wire_14395),
        .dout(new_Jinkela_wire_14396)
    );

    bfr new_Jinkela_buffer_11988 (
        .din(new_Jinkela_wire_14461),
        .dout(new_Jinkela_wire_14462)
    );

    bfr new_Jinkela_buffer_11925 (
        .din(new_Jinkela_wire_14396),
        .dout(new_Jinkela_wire_14397)
    );

    spl2 new_Jinkela_splitter_1093 (
        .a(_0421_),
        .b(new_Jinkela_wire_14683),
        .c(new_Jinkela_wire_14684)
    );

    bfr new_Jinkela_buffer_12080 (
        .din(new_Jinkela_wire_14557),
        .dout(new_Jinkela_wire_14558)
    );

    bfr new_Jinkela_buffer_11926 (
        .din(new_Jinkela_wire_14397),
        .dout(new_Jinkela_wire_14398)
    );

    bfr new_Jinkela_buffer_11989 (
        .din(new_Jinkela_wire_14462),
        .dout(new_Jinkela_wire_14463)
    );

    bfr new_Jinkela_buffer_11927 (
        .din(new_Jinkela_wire_14398),
        .dout(new_Jinkela_wire_14399)
    );

    bfr new_Jinkela_buffer_12109 (
        .din(new_Jinkela_wire_14586),
        .dout(new_Jinkela_wire_14587)
    );

    bfr new_Jinkela_buffer_11928 (
        .din(new_Jinkela_wire_14399),
        .dout(new_Jinkela_wire_14400)
    );

    bfr new_Jinkela_buffer_11990 (
        .din(new_Jinkela_wire_14463),
        .dout(new_Jinkela_wire_14464)
    );

    bfr new_Jinkela_buffer_11929 (
        .din(new_Jinkela_wire_14400),
        .dout(new_Jinkela_wire_14401)
    );

    bfr new_Jinkela_buffer_12081 (
        .din(new_Jinkela_wire_14558),
        .dout(new_Jinkela_wire_14559)
    );

    bfr new_Jinkela_buffer_11930 (
        .din(new_Jinkela_wire_14401),
        .dout(new_Jinkela_wire_14402)
    );

    bfr new_Jinkela_buffer_11991 (
        .din(new_Jinkela_wire_14464),
        .dout(new_Jinkela_wire_14465)
    );

    bfr new_Jinkela_buffer_11931 (
        .din(new_Jinkela_wire_14402),
        .dout(new_Jinkela_wire_14403)
    );

    bfr new_Jinkela_buffer_11932 (
        .din(new_Jinkela_wire_14403),
        .dout(new_Jinkela_wire_14404)
    );

    bfr new_Jinkela_buffer_11992 (
        .din(new_Jinkela_wire_14465),
        .dout(new_Jinkela_wire_14466)
    );

    bfr new_Jinkela_buffer_11933 (
        .din(new_Jinkela_wire_14404),
        .dout(new_Jinkela_wire_14405)
    );

    bfr new_Jinkela_buffer_12180 (
        .din(new_Jinkela_wire_14665),
        .dout(new_Jinkela_wire_14666)
    );

    bfr new_Jinkela_buffer_12082 (
        .din(new_Jinkela_wire_14559),
        .dout(new_Jinkela_wire_14560)
    );

    bfr new_Jinkela_buffer_11934 (
        .din(new_Jinkela_wire_14405),
        .dout(new_Jinkela_wire_14406)
    );

    bfr new_Jinkela_buffer_11993 (
        .din(new_Jinkela_wire_14466),
        .dout(new_Jinkela_wire_14467)
    );

    bfr new_Jinkela_buffer_11935 (
        .din(new_Jinkela_wire_14406),
        .dout(new_Jinkela_wire_14407)
    );

    bfr new_Jinkela_buffer_12110 (
        .din(new_Jinkela_wire_14587),
        .dout(new_Jinkela_wire_14588)
    );

    bfr new_Jinkela_buffer_11936 (
        .din(new_Jinkela_wire_14407),
        .dout(new_Jinkela_wire_14408)
    );

    bfr new_Jinkela_buffer_11994 (
        .din(new_Jinkela_wire_14467),
        .dout(new_Jinkela_wire_14468)
    );

    bfr new_Jinkela_buffer_11937 (
        .din(new_Jinkela_wire_14408),
        .dout(new_Jinkela_wire_14409)
    );

    bfr new_Jinkela_buffer_12083 (
        .din(new_Jinkela_wire_14560),
        .dout(new_Jinkela_wire_14561)
    );

    bfr new_Jinkela_buffer_11938 (
        .din(new_Jinkela_wire_14409),
        .dout(new_Jinkela_wire_14410)
    );

    bfr new_Jinkela_buffer_11995 (
        .din(new_Jinkela_wire_14468),
        .dout(new_Jinkela_wire_14469)
    );

    bfr new_Jinkela_buffer_11939 (
        .din(new_Jinkela_wire_14410),
        .dout(new_Jinkela_wire_14411)
    );

    bfr new_Jinkela_buffer_11940 (
        .din(new_Jinkela_wire_14411),
        .dout(new_Jinkela_wire_14412)
    );

    bfr new_Jinkela_buffer_8444 (
        .din(new_Jinkela_wire_10385),
        .dout(new_Jinkela_wire_10386)
    );

    bfr new_Jinkela_buffer_8526 (
        .din(new_Jinkela_wire_10477),
        .dout(new_Jinkela_wire_10478)
    );

    bfr new_Jinkela_buffer_8445 (
        .din(new_Jinkela_wire_10386),
        .dout(new_Jinkela_wire_10387)
    );

    bfr new_Jinkela_buffer_8705 (
        .din(_0252_),
        .dout(new_Jinkela_wire_10677)
    );

    bfr new_Jinkela_buffer_8706 (
        .din(_0110_),
        .dout(new_Jinkela_wire_10680)
    );

    bfr new_Jinkela_buffer_8446 (
        .din(new_Jinkela_wire_10387),
        .dout(new_Jinkela_wire_10388)
    );

    bfr new_Jinkela_buffer_8527 (
        .din(new_Jinkela_wire_10478),
        .dout(new_Jinkela_wire_10479)
    );

    bfr new_Jinkela_buffer_8447 (
        .din(new_Jinkela_wire_10388),
        .dout(new_Jinkela_wire_10389)
    );

    bfr new_Jinkela_buffer_8621 (
        .din(new_Jinkela_wire_10584),
        .dout(new_Jinkela_wire_10585)
    );

    bfr new_Jinkela_buffer_8448 (
        .din(new_Jinkela_wire_10389),
        .dout(new_Jinkela_wire_10390)
    );

    bfr new_Jinkela_buffer_8528 (
        .din(new_Jinkela_wire_10479),
        .dout(new_Jinkela_wire_10480)
    );

    bfr new_Jinkela_buffer_8449 (
        .din(new_Jinkela_wire_10390),
        .dout(new_Jinkela_wire_10391)
    );

    bfr new_Jinkela_buffer_8650 (
        .din(new_Jinkela_wire_10617),
        .dout(new_Jinkela_wire_10618)
    );

    spl2 new_Jinkela_splitter_820 (
        .a(new_Jinkela_wire_10391),
        .b(new_Jinkela_wire_10392),
        .c(new_Jinkela_wire_10393)
    );

    bfr new_Jinkela_buffer_8622 (
        .din(new_Jinkela_wire_10585),
        .dout(new_Jinkela_wire_10586)
    );

    bfr new_Jinkela_buffer_8529 (
        .din(new_Jinkela_wire_10480),
        .dout(new_Jinkela_wire_10481)
    );

    bfr new_Jinkela_buffer_8530 (
        .din(new_Jinkela_wire_10481),
        .dout(new_Jinkela_wire_10482)
    );

    bfr new_Jinkela_buffer_8531 (
        .din(new_Jinkela_wire_10482),
        .dout(new_Jinkela_wire_10483)
    );

    bfr new_Jinkela_buffer_8623 (
        .din(new_Jinkela_wire_10586),
        .dout(new_Jinkela_wire_10587)
    );

    bfr new_Jinkela_buffer_8532 (
        .din(new_Jinkela_wire_10483),
        .dout(new_Jinkela_wire_10484)
    );

    bfr new_Jinkela_buffer_8651 (
        .din(new_Jinkela_wire_10618),
        .dout(new_Jinkela_wire_10619)
    );

    bfr new_Jinkela_buffer_8533 (
        .din(new_Jinkela_wire_10484),
        .dout(new_Jinkela_wire_10485)
    );

    bfr new_Jinkela_buffer_8624 (
        .din(new_Jinkela_wire_10587),
        .dout(new_Jinkela_wire_10588)
    );

    bfr new_Jinkela_buffer_8534 (
        .din(new_Jinkela_wire_10485),
        .dout(new_Jinkela_wire_10486)
    );

    spl2 new_Jinkela_splitter_835 (
        .a(_1123_),
        .b(new_Jinkela_wire_10678),
        .c(new_Jinkela_wire_10679)
    );

    bfr new_Jinkela_buffer_8535 (
        .din(new_Jinkela_wire_10486),
        .dout(new_Jinkela_wire_10487)
    );

    bfr new_Jinkela_buffer_8625 (
        .din(new_Jinkela_wire_10588),
        .dout(new_Jinkela_wire_10589)
    );

    bfr new_Jinkela_buffer_8536 (
        .din(new_Jinkela_wire_10487),
        .dout(new_Jinkela_wire_10488)
    );

    bfr new_Jinkela_buffer_8652 (
        .din(new_Jinkela_wire_10619),
        .dout(new_Jinkela_wire_10620)
    );

    bfr new_Jinkela_buffer_8537 (
        .din(new_Jinkela_wire_10488),
        .dout(new_Jinkela_wire_10489)
    );

    bfr new_Jinkela_buffer_8626 (
        .din(new_Jinkela_wire_10589),
        .dout(new_Jinkela_wire_10590)
    );

    bfr new_Jinkela_buffer_8538 (
        .din(new_Jinkela_wire_10489),
        .dout(new_Jinkela_wire_10490)
    );

    spl2 new_Jinkela_splitter_836 (
        .a(_0983_),
        .b(new_Jinkela_wire_10682),
        .c(new_Jinkela_wire_10683)
    );

    bfr new_Jinkela_buffer_8539 (
        .din(new_Jinkela_wire_10490),
        .dout(new_Jinkela_wire_10491)
    );

    bfr new_Jinkela_buffer_8627 (
        .din(new_Jinkela_wire_10590),
        .dout(new_Jinkela_wire_10591)
    );

    bfr new_Jinkela_buffer_8540 (
        .din(new_Jinkela_wire_10491),
        .dout(new_Jinkela_wire_10492)
    );

    bfr new_Jinkela_buffer_8653 (
        .din(new_Jinkela_wire_10620),
        .dout(new_Jinkela_wire_10621)
    );

    bfr new_Jinkela_buffer_8541 (
        .din(new_Jinkela_wire_10492),
        .dout(new_Jinkela_wire_10493)
    );

    bfr new_Jinkela_buffer_8628 (
        .din(new_Jinkela_wire_10591),
        .dout(new_Jinkela_wire_10592)
    );

    bfr new_Jinkela_buffer_8542 (
        .din(new_Jinkela_wire_10493),
        .dout(new_Jinkela_wire_10494)
    );

    bfr new_Jinkela_buffer_8707 (
        .din(_1253_),
        .dout(new_Jinkela_wire_10681)
    );

    bfr new_Jinkela_buffer_8543 (
        .din(new_Jinkela_wire_10494),
        .dout(new_Jinkela_wire_10495)
    );

    bfr new_Jinkela_buffer_5075 (
        .din(new_Jinkela_wire_6548),
        .dout(new_Jinkela_wire_6549)
    );

    bfr new_Jinkela_buffer_5008 (
        .din(new_Jinkela_wire_6467),
        .dout(new_Jinkela_wire_6468)
    );

    bfr new_Jinkela_buffer_5148 (
        .din(new_Jinkela_wire_6625),
        .dout(new_Jinkela_wire_6626)
    );

    bfr new_Jinkela_buffer_5009 (
        .din(new_Jinkela_wire_6468),
        .dout(new_Jinkela_wire_6469)
    );

    bfr new_Jinkela_buffer_5076 (
        .din(new_Jinkela_wire_6549),
        .dout(new_Jinkela_wire_6550)
    );

    bfr new_Jinkela_buffer_5010 (
        .din(new_Jinkela_wire_6469),
        .dout(new_Jinkela_wire_6470)
    );

    bfr new_Jinkela_buffer_5203 (
        .din(_1200_),
        .dout(new_Jinkela_wire_6691)
    );

    bfr new_Jinkela_buffer_5199 (
        .din(new_Jinkela_wire_6686),
        .dout(new_Jinkela_wire_6687)
    );

    bfr new_Jinkela_buffer_5011 (
        .din(new_Jinkela_wire_6470),
        .dout(new_Jinkela_wire_6471)
    );

    bfr new_Jinkela_buffer_5077 (
        .din(new_Jinkela_wire_6550),
        .dout(new_Jinkela_wire_6551)
    );

    bfr new_Jinkela_buffer_5012 (
        .din(new_Jinkela_wire_6471),
        .dout(new_Jinkela_wire_6472)
    );

    bfr new_Jinkela_buffer_5149 (
        .din(new_Jinkela_wire_6626),
        .dout(new_Jinkela_wire_6627)
    );

    bfr new_Jinkela_buffer_5013 (
        .din(new_Jinkela_wire_6472),
        .dout(new_Jinkela_wire_6473)
    );

    bfr new_Jinkela_buffer_5078 (
        .din(new_Jinkela_wire_6551),
        .dout(new_Jinkela_wire_6552)
    );

    bfr new_Jinkela_buffer_5014 (
        .din(new_Jinkela_wire_6473),
        .dout(new_Jinkela_wire_6474)
    );

    bfr new_Jinkela_buffer_5015 (
        .din(new_Jinkela_wire_6474),
        .dout(new_Jinkela_wire_6475)
    );

    bfr new_Jinkela_buffer_5079 (
        .din(new_Jinkela_wire_6552),
        .dout(new_Jinkela_wire_6553)
    );

    bfr new_Jinkela_buffer_5016 (
        .din(new_Jinkela_wire_6475),
        .dout(new_Jinkela_wire_6476)
    );

    bfr new_Jinkela_buffer_5150 (
        .din(new_Jinkela_wire_6627),
        .dout(new_Jinkela_wire_6628)
    );

    bfr new_Jinkela_buffer_5017 (
        .din(new_Jinkela_wire_6476),
        .dout(new_Jinkela_wire_6477)
    );

    bfr new_Jinkela_buffer_5080 (
        .din(new_Jinkela_wire_6553),
        .dout(new_Jinkela_wire_6554)
    );

    bfr new_Jinkela_buffer_5018 (
        .din(new_Jinkela_wire_6477),
        .dout(new_Jinkela_wire_6478)
    );

    bfr new_Jinkela_buffer_5204 (
        .din(_1134_),
        .dout(new_Jinkela_wire_6692)
    );

    bfr new_Jinkela_buffer_5019 (
        .din(new_Jinkela_wire_6478),
        .dout(new_Jinkela_wire_6479)
    );

    bfr new_Jinkela_buffer_5081 (
        .din(new_Jinkela_wire_6554),
        .dout(new_Jinkela_wire_6555)
    );

    bfr new_Jinkela_buffer_5020 (
        .din(new_Jinkela_wire_6479),
        .dout(new_Jinkela_wire_6480)
    );

    bfr new_Jinkela_buffer_5151 (
        .din(new_Jinkela_wire_6628),
        .dout(new_Jinkela_wire_6629)
    );

    bfr new_Jinkela_buffer_5021 (
        .din(new_Jinkela_wire_6480),
        .dout(new_Jinkela_wire_6481)
    );

    bfr new_Jinkela_buffer_5082 (
        .din(new_Jinkela_wire_6555),
        .dout(new_Jinkela_wire_6556)
    );

    bfr new_Jinkela_buffer_5022 (
        .din(new_Jinkela_wire_6481),
        .dout(new_Jinkela_wire_6482)
    );

    bfr new_Jinkela_buffer_5244 (
        .din(_0353_),
        .dout(new_Jinkela_wire_6734)
    );

    bfr new_Jinkela_buffer_5023 (
        .din(new_Jinkela_wire_6482),
        .dout(new_Jinkela_wire_6483)
    );

    bfr new_Jinkela_buffer_5083 (
        .din(new_Jinkela_wire_6556),
        .dout(new_Jinkela_wire_6557)
    );

    bfr new_Jinkela_buffer_5024 (
        .din(new_Jinkela_wire_6483),
        .dout(new_Jinkela_wire_6484)
    );

    bfr new_Jinkela_buffer_5152 (
        .din(new_Jinkela_wire_6629),
        .dout(new_Jinkela_wire_6630)
    );

    bfr new_Jinkela_buffer_5025 (
        .din(new_Jinkela_wire_6484),
        .dout(new_Jinkela_wire_6485)
    );

    bfr new_Jinkela_buffer_5084 (
        .din(new_Jinkela_wire_6557),
        .dout(new_Jinkela_wire_6558)
    );

    bfr new_Jinkela_buffer_5026 (
        .din(new_Jinkela_wire_6485),
        .dout(new_Jinkela_wire_6486)
    );

    bfr new_Jinkela_buffer_5200 (
        .din(new_Jinkela_wire_6687),
        .dout(new_Jinkela_wire_6688)
    );

    bfr new_Jinkela_buffer_5027 (
        .din(new_Jinkela_wire_6486),
        .dout(new_Jinkela_wire_6487)
    );

    bfr new_Jinkela_buffer_5085 (
        .din(new_Jinkela_wire_6558),
        .dout(new_Jinkela_wire_6559)
    );

    bfr new_Jinkela_buffer_5028 (
        .din(new_Jinkela_wire_6487),
        .dout(new_Jinkela_wire_6488)
    );

    bfr new_Jinkela_buffer_11996 (
        .din(new_Jinkela_wire_14469),
        .dout(new_Jinkela_wire_14470)
    );

    and_bb _2623_ (
        .a(new_Jinkela_wire_10974),
        .b(new_Jinkela_wire_3662),
        .c(_1677_)
    );

    bfr new_Jinkela_buffer_11941 (
        .din(new_Jinkela_wire_14412),
        .dout(new_Jinkela_wire_14413)
    );

    or_bb _2624_ (
        .a(new_Jinkela_wire_16969),
        .b(new_Jinkela_wire_2120),
        .c(new_net_3942)
    );

    bfr new_Jinkela_buffer_12195 (
        .din(_0967_),
        .dout(new_Jinkela_wire_14689)
    );

    and_bb _2625_ (
        .a(new_Jinkela_wire_667),
        .b(new_Jinkela_wire_348),
        .c(_1678_)
    );

    bfr new_Jinkela_buffer_12084 (
        .din(new_Jinkela_wire_14561),
        .dout(new_Jinkela_wire_14562)
    );

    bfr new_Jinkela_buffer_11942 (
        .din(new_Jinkela_wire_14413),
        .dout(new_Jinkela_wire_14414)
    );

    and_bi _2626_ (
        .a(new_Jinkela_wire_5097),
        .b(new_Jinkela_wire_2121),
        .c(_1679_)
    );

    bfr new_Jinkela_buffer_11997 (
        .din(new_Jinkela_wire_14470),
        .dout(new_Jinkela_wire_14471)
    );

    and_bb _2627_ (
        .a(new_Jinkela_wire_91),
        .b(new_Jinkela_wire_527),
        .c(_1680_)
    );

    bfr new_Jinkela_buffer_11943 (
        .din(new_Jinkela_wire_14414),
        .dout(new_Jinkela_wire_14415)
    );

    and_bi _2628_ (
        .a(new_Jinkela_wire_713),
        .b(new_Jinkela_wire_17360),
        .c(_1681_)
    );

    and_bb _2629_ (
        .a(new_Jinkela_wire_148),
        .b(new_Jinkela_wire_556),
        .c(_1682_)
    );

    bfr new_Jinkela_buffer_12111 (
        .din(new_Jinkela_wire_14588),
        .dout(new_Jinkela_wire_14589)
    );

    bfr new_Jinkela_buffer_11944 (
        .din(new_Jinkela_wire_14415),
        .dout(new_Jinkela_wire_14416)
    );

    and_bi _2630_ (
        .a(new_Jinkela_wire_12050),
        .b(new_Jinkela_wire_2144),
        .c(_1683_)
    );

    bfr new_Jinkela_buffer_11998 (
        .din(new_Jinkela_wire_14471),
        .dout(new_Jinkela_wire_14472)
    );

    and_bb _2631_ (
        .a(new_Jinkela_wire_278),
        .b(new_Jinkela_wire_209),
        .c(_1684_)
    );

    bfr new_Jinkela_buffer_11945 (
        .din(new_Jinkela_wire_14416),
        .dout(new_Jinkela_wire_14417)
    );

    and_bi _2632_ (
        .a(new_Jinkela_wire_16914),
        .b(new_Jinkela_wire_12342),
        .c(_1685_)
    );

    and_bb _2633_ (
        .a(new_Jinkela_wire_77),
        .b(new_Jinkela_wire_573),
        .c(_1687_)
    );

    bfr new_Jinkela_buffer_12085 (
        .din(new_Jinkela_wire_14562),
        .dout(new_Jinkela_wire_14563)
    );

    bfr new_Jinkela_buffer_11946 (
        .din(new_Jinkela_wire_14417),
        .dout(new_Jinkela_wire_14418)
    );

    and_bi _2634_ (
        .a(new_Jinkela_wire_13386),
        .b(new_Jinkela_wire_2599),
        .c(_1688_)
    );

    bfr new_Jinkela_buffer_11999 (
        .din(new_Jinkela_wire_14472),
        .dout(new_Jinkela_wire_14473)
    );

    and_bb _2635_ (
        .a(new_Jinkela_wire_472),
        .b(new_Jinkela_wire_125),
        .c(_1689_)
    );

    bfr new_Jinkela_buffer_11947 (
        .din(new_Jinkela_wire_14418),
        .dout(new_Jinkela_wire_14419)
    );

    and_bi _2636_ (
        .a(new_Jinkela_wire_13212),
        .b(new_Jinkela_wire_13968),
        .c(_1690_)
    );

    and_bb _2637_ (
        .a(new_Jinkela_wire_353),
        .b(new_Jinkela_wire_18),
        .c(_1691_)
    );

    bfr new_Jinkela_buffer_11948 (
        .din(new_Jinkela_wire_14419),
        .dout(new_Jinkela_wire_14420)
    );

    and_bi _2638_ (
        .a(new_Jinkela_wire_17667),
        .b(new_Jinkela_wire_1139),
        .c(_1692_)
    );

    bfr new_Jinkela_buffer_12000 (
        .din(new_Jinkela_wire_14473),
        .dout(new_Jinkela_wire_14474)
    );

    and_bb _2639_ (
        .a(new_Jinkela_wire_688),
        .b(new_Jinkela_wire_454),
        .c(_1693_)
    );

    bfr new_Jinkela_buffer_11949 (
        .din(new_Jinkela_wire_14420),
        .dout(new_Jinkela_wire_14421)
    );

    and_bi _2640_ (
        .a(new_Jinkela_wire_12336),
        .b(new_Jinkela_wire_11725),
        .c(_1694_)
    );

    bfr new_Jinkela_buffer_12181 (
        .din(new_Jinkela_wire_14666),
        .dout(new_Jinkela_wire_14667)
    );

    and_bb _2641_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_505),
        .c(_1695_)
    );

    bfr new_Jinkela_buffer_12086 (
        .din(new_Jinkela_wire_14563),
        .dout(new_Jinkela_wire_14564)
    );

    bfr new_Jinkela_buffer_11950 (
        .din(new_Jinkela_wire_14421),
        .dout(new_Jinkela_wire_14422)
    );

    and_bi _2642_ (
        .a(new_Jinkela_wire_4687),
        .b(new_Jinkela_wire_12712),
        .c(_1696_)
    );

    bfr new_Jinkela_buffer_12001 (
        .din(new_Jinkela_wire_14474),
        .dout(new_Jinkela_wire_14475)
    );

    and_bb _2643_ (
        .a(new_Jinkela_wire_31),
        .b(new_Jinkela_wire_301),
        .c(_1698_)
    );

    bfr new_Jinkela_buffer_11951 (
        .din(new_Jinkela_wire_14422),
        .dout(new_Jinkela_wire_14423)
    );

    and_bi _2644_ (
        .a(new_Jinkela_wire_10962),
        .b(new_Jinkela_wire_16103),
        .c(_1699_)
    );

    and_bb _2645_ (
        .a(new_Jinkela_wire_194),
        .b(new_Jinkela_wire_63),
        .c(_1700_)
    );

    bfr new_Jinkela_buffer_12112 (
        .din(new_Jinkela_wire_14589),
        .dout(new_Jinkela_wire_14590)
    );

    bfr new_Jinkela_buffer_11952 (
        .din(new_Jinkela_wire_14423),
        .dout(new_Jinkela_wire_14424)
    );

    and_bi _2646_ (
        .a(new_Jinkela_wire_12110),
        .b(new_Jinkela_wire_4718),
        .c(_1701_)
    );

    bfr new_Jinkela_buffer_12002 (
        .din(new_Jinkela_wire_14475),
        .dout(new_Jinkela_wire_14476)
    );

    and_bb _2647_ (
        .a(new_Jinkela_wire_375),
        .b(new_Jinkela_wire_650),
        .c(_1702_)
    );

    bfr new_Jinkela_buffer_11953 (
        .din(new_Jinkela_wire_14424),
        .dout(new_Jinkela_wire_14425)
    );

    and_bi _2648_ (
        .a(new_Jinkela_wire_16130),
        .b(new_Jinkela_wire_4987),
        .c(_1703_)
    );

    and_bb _2649_ (
        .a(new_Jinkela_wire_402),
        .b(new_Jinkela_wire_624),
        .c(_1704_)
    );

    bfr new_Jinkela_buffer_12087 (
        .din(new_Jinkela_wire_14564),
        .dout(new_Jinkela_wire_14565)
    );

    spl2 new_Jinkela_splitter_1085 (
        .a(new_Jinkela_wire_14425),
        .b(new_Jinkela_wire_14426),
        .c(new_Jinkela_wire_14427)
    );

    and_bi _2650_ (
        .a(new_Jinkela_wire_19289),
        .b(new_Jinkela_wire_14020),
        .c(_1705_)
    );

    and_bb _2651_ (
        .a(new_Jinkela_wire_171),
        .b(new_Jinkela_wire_543),
        .c(_1706_)
    );

    bfr new_Jinkela_buffer_12003 (
        .din(new_Jinkela_wire_14476),
        .dout(new_Jinkela_wire_14477)
    );

    and_ii _2652_ (
        .a(new_Jinkela_wire_11458),
        .b(new_Jinkela_wire_442),
        .c(_1707_)
    );

    bfr new_Jinkela_buffer_12004 (
        .din(new_Jinkela_wire_14477),
        .dout(new_Jinkela_wire_14478)
    );

    and_bb _2653_ (
        .a(new_Jinkela_wire_432),
        .b(new_Jinkela_wire_230),
        .c(_1709_)
    );

    and_bi _2654_ (
        .a(new_Jinkela_wire_17108),
        .b(new_Jinkela_wire_7309),
        .c(_1710_)
    );

    bfr new_Jinkela_buffer_12088 (
        .din(new_Jinkela_wire_14565),
        .dout(new_Jinkela_wire_14566)
    );

    bfr new_Jinkela_buffer_12005 (
        .din(new_Jinkela_wire_14478),
        .dout(new_Jinkela_wire_14479)
    );

    or_bb _2655_ (
        .a(new_Jinkela_wire_17110),
        .b(new_Jinkela_wire_176),
        .c(_1711_)
    );

    and_bi _2656_ (
        .a(new_Jinkela_wire_7311),
        .b(_1711_),
        .c(_1712_)
    );

    bfr new_Jinkela_buffer_12113 (
        .din(new_Jinkela_wire_14590),
        .dout(new_Jinkela_wire_14591)
    );

    bfr new_Jinkela_buffer_12006 (
        .din(new_Jinkela_wire_14479),
        .dout(new_Jinkela_wire_14480)
    );

    or_bb _2657_ (
        .a(_1712_),
        .b(new_Jinkela_wire_3190),
        .c(_1713_)
    );

    or_bb _2658_ (
        .a(new_Jinkela_wire_15689),
        .b(_1707_),
        .c(_1714_)
    );

    bfr new_Jinkela_buffer_12089 (
        .din(new_Jinkela_wire_14566),
        .dout(new_Jinkela_wire_14567)
    );

    bfr new_Jinkela_buffer_12007 (
        .din(new_Jinkela_wire_14480),
        .dout(new_Jinkela_wire_14481)
    );

    and_ii _2659_ (
        .a(new_Jinkela_wire_8683),
        .b(new_Jinkela_wire_3267),
        .c(_1715_)
    );

    and_bb _2660_ (
        .a(new_Jinkela_wire_8684),
        .b(new_Jinkela_wire_3268),
        .c(_1716_)
    );

    spl2 new_Jinkela_splitter_1095 (
        .a(_0465_),
        .b(new_Jinkela_wire_14687),
        .c(new_Jinkela_wire_14688)
    );

    bfr new_Jinkela_buffer_12008 (
        .din(new_Jinkela_wire_14481),
        .dout(new_Jinkela_wire_14482)
    );

    or_bb _2661_ (
        .a(new_Jinkela_wire_18952),
        .b(new_Jinkela_wire_19114),
        .c(_1717_)
    );

    bfr new_Jinkela_buffer_12182 (
        .din(new_Jinkela_wire_14667),
        .dout(new_Jinkela_wire_14668)
    );

    or_bb _2662_ (
        .a(new_Jinkela_wire_17786),
        .b(new_Jinkela_wire_5800),
        .c(_1718_)
    );

    bfr new_Jinkela_buffer_12090 (
        .din(new_Jinkela_wire_14567),
        .dout(new_Jinkela_wire_14568)
    );

    bfr new_Jinkela_buffer_12009 (
        .din(new_Jinkela_wire_14482),
        .dout(new_Jinkela_wire_14483)
    );

    or_ii _2663_ (
        .a(new_Jinkela_wire_17787),
        .b(new_Jinkela_wire_5801),
        .c(_1720_)
    );

    or_ii _2664_ (
        .a(new_Jinkela_wire_12723),
        .b(new_Jinkela_wire_21099),
        .c(_1721_)
    );

    bfr new_Jinkela_buffer_12114 (
        .din(new_Jinkela_wire_14591),
        .dout(new_Jinkela_wire_14592)
    );

    bfr new_Jinkela_buffer_5153 (
        .din(new_Jinkela_wire_6630),
        .dout(new_Jinkela_wire_6631)
    );

    bfr new_Jinkela_buffer_5029 (
        .din(new_Jinkela_wire_6488),
        .dout(new_Jinkela_wire_6489)
    );

    bfr new_Jinkela_buffer_5086 (
        .din(new_Jinkela_wire_6559),
        .dout(new_Jinkela_wire_6560)
    );

    bfr new_Jinkela_buffer_5030 (
        .din(new_Jinkela_wire_6489),
        .dout(new_Jinkela_wire_6490)
    );

    spl2 new_Jinkela_splitter_594 (
        .a(_1506_),
        .b(new_Jinkela_wire_6735),
        .c(new_Jinkela_wire_6736)
    );

    bfr new_Jinkela_buffer_5031 (
        .din(new_Jinkela_wire_6490),
        .dout(new_Jinkela_wire_6491)
    );

    bfr new_Jinkela_buffer_5087 (
        .din(new_Jinkela_wire_6560),
        .dout(new_Jinkela_wire_6561)
    );

    bfr new_Jinkela_buffer_5032 (
        .din(new_Jinkela_wire_6491),
        .dout(new_Jinkela_wire_6492)
    );

    bfr new_Jinkela_buffer_5154 (
        .din(new_Jinkela_wire_6631),
        .dout(new_Jinkela_wire_6632)
    );

    bfr new_Jinkela_buffer_5033 (
        .din(new_Jinkela_wire_6492),
        .dout(new_Jinkela_wire_6493)
    );

    bfr new_Jinkela_buffer_5088 (
        .din(new_Jinkela_wire_6561),
        .dout(new_Jinkela_wire_6562)
    );

    bfr new_Jinkela_buffer_5034 (
        .din(new_Jinkela_wire_6493),
        .dout(new_Jinkela_wire_6494)
    );

    bfr new_Jinkela_buffer_5201 (
        .din(new_Jinkela_wire_6688),
        .dout(new_Jinkela_wire_6689)
    );

    bfr new_Jinkela_buffer_5035 (
        .din(new_Jinkela_wire_6494),
        .dout(new_Jinkela_wire_6495)
    );

    bfr new_Jinkela_buffer_5089 (
        .din(new_Jinkela_wire_6562),
        .dout(new_Jinkela_wire_6563)
    );

    bfr new_Jinkela_buffer_5036 (
        .din(new_Jinkela_wire_6495),
        .dout(new_Jinkela_wire_6496)
    );

    bfr new_Jinkela_buffer_5155 (
        .din(new_Jinkela_wire_6632),
        .dout(new_Jinkela_wire_6633)
    );

    bfr new_Jinkela_buffer_5037 (
        .din(new_Jinkela_wire_6496),
        .dout(new_Jinkela_wire_6497)
    );

    bfr new_Jinkela_buffer_5090 (
        .din(new_Jinkela_wire_6563),
        .dout(new_Jinkela_wire_6564)
    );

    bfr new_Jinkela_buffer_5038 (
        .din(new_Jinkela_wire_6497),
        .dout(new_Jinkela_wire_6498)
    );

    bfr new_Jinkela_buffer_5205 (
        .din(new_Jinkela_wire_6692),
        .dout(new_Jinkela_wire_6693)
    );

    bfr new_Jinkela_buffer_5039 (
        .din(new_Jinkela_wire_6498),
        .dout(new_Jinkela_wire_6499)
    );

    bfr new_Jinkela_buffer_5091 (
        .din(new_Jinkela_wire_6564),
        .dout(new_Jinkela_wire_6565)
    );

    bfr new_Jinkela_buffer_5040 (
        .din(new_Jinkela_wire_6499),
        .dout(new_Jinkela_wire_6500)
    );

    bfr new_Jinkela_buffer_5156 (
        .din(new_Jinkela_wire_6633),
        .dout(new_Jinkela_wire_6634)
    );

    bfr new_Jinkela_buffer_5041 (
        .din(new_Jinkela_wire_6500),
        .dout(new_Jinkela_wire_6501)
    );

    bfr new_Jinkela_buffer_5092 (
        .din(new_Jinkela_wire_6565),
        .dout(new_Jinkela_wire_6566)
    );

    bfr new_Jinkela_buffer_5042 (
        .din(new_Jinkela_wire_6501),
        .dout(new_Jinkela_wire_6502)
    );

    bfr new_Jinkela_buffer_5202 (
        .din(new_Jinkela_wire_6689),
        .dout(new_Jinkela_wire_6690)
    );

    bfr new_Jinkela_buffer_5043 (
        .din(new_Jinkela_wire_6502),
        .dout(new_Jinkela_wire_6503)
    );

    bfr new_Jinkela_buffer_5093 (
        .din(new_Jinkela_wire_6566),
        .dout(new_Jinkela_wire_6567)
    );

    bfr new_Jinkela_buffer_5044 (
        .din(new_Jinkela_wire_6503),
        .dout(new_Jinkela_wire_6504)
    );

    bfr new_Jinkela_buffer_5157 (
        .din(new_Jinkela_wire_6634),
        .dout(new_Jinkela_wire_6635)
    );

    bfr new_Jinkela_buffer_5045 (
        .din(new_Jinkela_wire_6504),
        .dout(new_Jinkela_wire_6505)
    );

    bfr new_Jinkela_buffer_5094 (
        .din(new_Jinkela_wire_6567),
        .dout(new_Jinkela_wire_6568)
    );

    bfr new_Jinkela_buffer_5046 (
        .din(new_Jinkela_wire_6505),
        .dout(new_Jinkela_wire_6506)
    );

    bfr new_Jinkela_buffer_5245 (
        .din(_0250_),
        .dout(new_Jinkela_wire_6737)
    );

    bfr new_Jinkela_buffer_5047 (
        .din(new_Jinkela_wire_6506),
        .dout(new_Jinkela_wire_6507)
    );

    bfr new_Jinkela_buffer_5095 (
        .din(new_Jinkela_wire_6568),
        .dout(new_Jinkela_wire_6569)
    );

    bfr new_Jinkela_buffer_5048 (
        .din(new_Jinkela_wire_6507),
        .dout(new_Jinkela_wire_6508)
    );

    bfr new_Jinkela_buffer_5158 (
        .din(new_Jinkela_wire_6635),
        .dout(new_Jinkela_wire_6636)
    );

    bfr new_Jinkela_buffer_5049 (
        .din(new_Jinkela_wire_6508),
        .dout(new_Jinkela_wire_6509)
    );

    bfr new_Jinkela_buffer_15450 (
        .din(new_Jinkela_wire_18416),
        .dout(new_Jinkela_wire_18417)
    );

    bfr new_Jinkela_buffer_15540 (
        .din(new_Jinkela_wire_18518),
        .dout(new_Jinkela_wire_18519)
    );

    bfr new_Jinkela_buffer_15451 (
        .din(new_Jinkela_wire_18417),
        .dout(new_Jinkela_wire_18418)
    );

    bfr new_Jinkela_buffer_15487 (
        .din(new_Jinkela_wire_18459),
        .dout(new_Jinkela_wire_18460)
    );

    bfr new_Jinkela_buffer_15452 (
        .din(new_Jinkela_wire_18418),
        .dout(new_Jinkela_wire_18419)
    );

    bfr new_Jinkela_buffer_15524 (
        .din(new_Jinkela_wire_18498),
        .dout(new_Jinkela_wire_18499)
    );

    bfr new_Jinkela_buffer_15453 (
        .din(new_Jinkela_wire_18419),
        .dout(new_Jinkela_wire_18420)
    );

    bfr new_Jinkela_buffer_15488 (
        .din(new_Jinkela_wire_18460),
        .dout(new_Jinkela_wire_18461)
    );

    bfr new_Jinkela_buffer_15454 (
        .din(new_Jinkela_wire_18420),
        .dout(new_Jinkela_wire_18421)
    );

    spl2 new_Jinkela_splitter_1340 (
        .a(_1374_),
        .b(new_Jinkela_wire_18528),
        .c(new_Jinkela_wire_18529)
    );

    bfr new_Jinkela_buffer_15455 (
        .din(new_Jinkela_wire_18421),
        .dout(new_Jinkela_wire_18422)
    );

    bfr new_Jinkela_buffer_15489 (
        .din(new_Jinkela_wire_18461),
        .dout(new_Jinkela_wire_18462)
    );

    bfr new_Jinkela_buffer_15456 (
        .din(new_Jinkela_wire_18422),
        .dout(new_Jinkela_wire_18423)
    );

    bfr new_Jinkela_buffer_15525 (
        .din(new_Jinkela_wire_18499),
        .dout(new_Jinkela_wire_18500)
    );

    bfr new_Jinkela_buffer_15457 (
        .din(new_Jinkela_wire_18423),
        .dout(new_Jinkela_wire_18424)
    );

    bfr new_Jinkela_buffer_15490 (
        .din(new_Jinkela_wire_18462),
        .dout(new_Jinkela_wire_18463)
    );

    bfr new_Jinkela_buffer_15458 (
        .din(new_Jinkela_wire_18424),
        .dout(new_Jinkela_wire_18425)
    );

    bfr new_Jinkela_buffer_15541 (
        .din(new_Jinkela_wire_18519),
        .dout(new_Jinkela_wire_18520)
    );

    bfr new_Jinkela_buffer_15459 (
        .din(new_Jinkela_wire_18425),
        .dout(new_Jinkela_wire_18426)
    );

    bfr new_Jinkela_buffer_15491 (
        .din(new_Jinkela_wire_18463),
        .dout(new_Jinkela_wire_18464)
    );

    bfr new_Jinkela_buffer_15460 (
        .din(new_Jinkela_wire_18426),
        .dout(new_Jinkela_wire_18427)
    );

    bfr new_Jinkela_buffer_15526 (
        .din(new_Jinkela_wire_18500),
        .dout(new_Jinkela_wire_18501)
    );

    bfr new_Jinkela_buffer_15461 (
        .din(new_Jinkela_wire_18427),
        .dout(new_Jinkela_wire_18428)
    );

    bfr new_Jinkela_buffer_15492 (
        .din(new_Jinkela_wire_18464),
        .dout(new_Jinkela_wire_18465)
    );

    bfr new_Jinkela_buffer_15462 (
        .din(new_Jinkela_wire_18428),
        .dout(new_Jinkela_wire_18429)
    );

    spl2 new_Jinkela_splitter_1339 (
        .a(_1230_),
        .b(new_Jinkela_wire_18526),
        .c(new_Jinkela_wire_18527)
    );

    bfr new_Jinkela_buffer_15463 (
        .din(new_Jinkela_wire_18429),
        .dout(new_Jinkela_wire_18430)
    );

    bfr new_Jinkela_buffer_15493 (
        .din(new_Jinkela_wire_18465),
        .dout(new_Jinkela_wire_18466)
    );

    bfr new_Jinkela_buffer_15464 (
        .din(new_Jinkela_wire_18430),
        .dout(new_Jinkela_wire_18431)
    );

    bfr new_Jinkela_buffer_15527 (
        .din(new_Jinkela_wire_18501),
        .dout(new_Jinkela_wire_18502)
    );

    bfr new_Jinkela_buffer_15465 (
        .din(new_Jinkela_wire_18431),
        .dout(new_Jinkela_wire_18432)
    );

    bfr new_Jinkela_buffer_15494 (
        .din(new_Jinkela_wire_18466),
        .dout(new_Jinkela_wire_18467)
    );

    bfr new_Jinkela_buffer_15466 (
        .din(new_Jinkela_wire_18432),
        .dout(new_Jinkela_wire_18433)
    );

    bfr new_Jinkela_buffer_15542 (
        .din(new_Jinkela_wire_18520),
        .dout(new_Jinkela_wire_18521)
    );

    bfr new_Jinkela_buffer_15467 (
        .din(new_Jinkela_wire_18433),
        .dout(new_Jinkela_wire_18434)
    );

    bfr new_Jinkela_buffer_15495 (
        .din(new_Jinkela_wire_18467),
        .dout(new_Jinkela_wire_18468)
    );

    bfr new_Jinkela_buffer_15468 (
        .din(new_Jinkela_wire_18434),
        .dout(new_Jinkela_wire_18435)
    );

    bfr new_Jinkela_buffer_15528 (
        .din(new_Jinkela_wire_18502),
        .dout(new_Jinkela_wire_18503)
    );

    bfr new_Jinkela_buffer_15469 (
        .din(new_Jinkela_wire_18435),
        .dout(new_Jinkela_wire_18436)
    );

    bfr new_Jinkela_buffer_15496 (
        .din(new_Jinkela_wire_18468),
        .dout(new_Jinkela_wire_18469)
    );

    bfr new_Jinkela_buffer_15470 (
        .din(new_Jinkela_wire_18436),
        .dout(new_Jinkela_wire_18437)
    );

    spl2 new_Jinkela_splitter_1341 (
        .a(_0655_),
        .b(new_Jinkela_wire_18530),
        .c(new_Jinkela_wire_18531)
    );

    bfr new_Jinkela_buffer_5096 (
        .din(new_Jinkela_wire_6569),
        .dout(new_Jinkela_wire_6570)
    );

    spl2 new_Jinkela_splitter_579 (
        .a(new_Jinkela_wire_6509),
        .b(new_Jinkela_wire_6510),
        .c(new_Jinkela_wire_6511)
    );

    bfr new_Jinkela_buffer_5097 (
        .din(new_Jinkela_wire_6570),
        .dout(new_Jinkela_wire_6571)
    );

    bfr new_Jinkela_buffer_5206 (
        .din(new_Jinkela_wire_6693),
        .dout(new_Jinkela_wire_6694)
    );

    bfr new_Jinkela_buffer_5159 (
        .din(new_Jinkela_wire_6636),
        .dout(new_Jinkela_wire_6637)
    );

    bfr new_Jinkela_buffer_5098 (
        .din(new_Jinkela_wire_6571),
        .dout(new_Jinkela_wire_6572)
    );

    bfr new_Jinkela_buffer_5247 (
        .din(_1584_),
        .dout(new_Jinkela_wire_6739)
    );

    bfr new_Jinkela_buffer_5099 (
        .din(new_Jinkela_wire_6572),
        .dout(new_Jinkela_wire_6573)
    );

    bfr new_Jinkela_buffer_5160 (
        .din(new_Jinkela_wire_6637),
        .dout(new_Jinkela_wire_6638)
    );

    bfr new_Jinkela_buffer_5100 (
        .din(new_Jinkela_wire_6573),
        .dout(new_Jinkela_wire_6574)
    );

    bfr new_Jinkela_buffer_5207 (
        .din(new_Jinkela_wire_6694),
        .dout(new_Jinkela_wire_6695)
    );

    bfr new_Jinkela_buffer_5101 (
        .din(new_Jinkela_wire_6574),
        .dout(new_Jinkela_wire_6575)
    );

    bfr new_Jinkela_buffer_5161 (
        .din(new_Jinkela_wire_6638),
        .dout(new_Jinkela_wire_6639)
    );

    bfr new_Jinkela_buffer_5102 (
        .din(new_Jinkela_wire_6575),
        .dout(new_Jinkela_wire_6576)
    );

    bfr new_Jinkela_buffer_5246 (
        .din(_1442_),
        .dout(new_Jinkela_wire_6738)
    );

    bfr new_Jinkela_buffer_5103 (
        .din(new_Jinkela_wire_6576),
        .dout(new_Jinkela_wire_6577)
    );

    bfr new_Jinkela_buffer_5162 (
        .din(new_Jinkela_wire_6639),
        .dout(new_Jinkela_wire_6640)
    );

    bfr new_Jinkela_buffer_5104 (
        .din(new_Jinkela_wire_6577),
        .dout(new_Jinkela_wire_6578)
    );

    bfr new_Jinkela_buffer_5208 (
        .din(new_Jinkela_wire_6695),
        .dout(new_Jinkela_wire_6696)
    );

    bfr new_Jinkela_buffer_5105 (
        .din(new_Jinkela_wire_6578),
        .dout(new_Jinkela_wire_6579)
    );

    bfr new_Jinkela_buffer_5163 (
        .din(new_Jinkela_wire_6640),
        .dout(new_Jinkela_wire_6641)
    );

    bfr new_Jinkela_buffer_5106 (
        .din(new_Jinkela_wire_6579),
        .dout(new_Jinkela_wire_6580)
    );

    spl2 new_Jinkela_splitter_596 (
        .a(_0471_),
        .b(new_Jinkela_wire_6757),
        .c(new_Jinkela_wire_6758)
    );

    bfr new_Jinkela_buffer_5107 (
        .din(new_Jinkela_wire_6580),
        .dout(new_Jinkela_wire_6581)
    );

    bfr new_Jinkela_buffer_5164 (
        .din(new_Jinkela_wire_6641),
        .dout(new_Jinkela_wire_6642)
    );

    bfr new_Jinkela_buffer_5108 (
        .din(new_Jinkela_wire_6581),
        .dout(new_Jinkela_wire_6582)
    );

    bfr new_Jinkela_buffer_5209 (
        .din(new_Jinkela_wire_6696),
        .dout(new_Jinkela_wire_6697)
    );

    bfr new_Jinkela_buffer_5109 (
        .din(new_Jinkela_wire_6582),
        .dout(new_Jinkela_wire_6583)
    );

    bfr new_Jinkela_buffer_5165 (
        .din(new_Jinkela_wire_6642),
        .dout(new_Jinkela_wire_6643)
    );

    bfr new_Jinkela_buffer_5110 (
        .din(new_Jinkela_wire_6583),
        .dout(new_Jinkela_wire_6584)
    );

    spl2 new_Jinkela_splitter_597 (
        .a(_0620_),
        .b(new_Jinkela_wire_6759),
        .c(new_Jinkela_wire_6760)
    );

    bfr new_Jinkela_buffer_5111 (
        .din(new_Jinkela_wire_6584),
        .dout(new_Jinkela_wire_6585)
    );

    bfr new_Jinkela_buffer_5166 (
        .din(new_Jinkela_wire_6643),
        .dout(new_Jinkela_wire_6644)
    );

    bfr new_Jinkela_buffer_5112 (
        .din(new_Jinkela_wire_6585),
        .dout(new_Jinkela_wire_6586)
    );

    bfr new_Jinkela_buffer_5210 (
        .din(new_Jinkela_wire_6697),
        .dout(new_Jinkela_wire_6698)
    );

    bfr new_Jinkela_buffer_5113 (
        .din(new_Jinkela_wire_6586),
        .dout(new_Jinkela_wire_6587)
    );

    bfr new_Jinkela_buffer_5167 (
        .din(new_Jinkela_wire_6644),
        .dout(new_Jinkela_wire_6645)
    );

    bfr new_Jinkela_buffer_5114 (
        .din(new_Jinkela_wire_6587),
        .dout(new_Jinkela_wire_6588)
    );

    bfr new_Jinkela_buffer_5248 (
        .din(new_Jinkela_wire_6739),
        .dout(new_Jinkela_wire_6740)
    );

    bfr new_Jinkela_buffer_5115 (
        .din(new_Jinkela_wire_6588),
        .dout(new_Jinkela_wire_6589)
    );

    bfr new_Jinkela_buffer_5168 (
        .din(new_Jinkela_wire_6645),
        .dout(new_Jinkela_wire_6646)
    );

    bfr new_Jinkela_buffer_5116 (
        .din(new_Jinkela_wire_6589),
        .dout(new_Jinkela_wire_6590)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_2434),
        .dout(new_Jinkela_wire_2435)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(new_Jinkela_wire_2372),
        .dout(new_Jinkela_wire_2373)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(_0928_),
        .dout(new_Jinkela_wire_2487)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_2373),
        .dout(new_Jinkela_wire_2374)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_2435),
        .dout(new_Jinkela_wire_2436)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_2374),
        .dout(new_Jinkela_wire_2375)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_2468),
        .dout(new_Jinkela_wire_2469)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(new_Jinkela_wire_2375),
        .dout(new_Jinkela_wire_2376)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_2436),
        .dout(new_Jinkela_wire_2437)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(new_Jinkela_wire_2376),
        .dout(new_Jinkela_wire_2377)
    );

    spl2 new_Jinkela_splitter_298 (
        .a(_1820_),
        .b(new_Jinkela_wire_2592),
        .c(new_Jinkela_wire_2593)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(new_Jinkela_wire_2377),
        .dout(new_Jinkela_wire_2378)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_2437),
        .dout(new_Jinkela_wire_2438)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_Jinkela_wire_2378),
        .dout(new_Jinkela_wire_2379)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(new_Jinkela_wire_2469),
        .dout(new_Jinkela_wire_2470)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_2379),
        .dout(new_Jinkela_wire_2380)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_2438),
        .dout(new_Jinkela_wire_2439)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_2380),
        .dout(new_Jinkela_wire_2381)
    );

    bfr new_Jinkela_buffer_1693 (
        .din(_0667_),
        .dout(new_Jinkela_wire_2591)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_2381),
        .dout(new_Jinkela_wire_2382)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_2439),
        .dout(new_Jinkela_wire_2440)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(new_Jinkela_wire_2382),
        .dout(new_Jinkela_wire_2383)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_2470),
        .dout(new_Jinkela_wire_2471)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(new_Jinkela_wire_2383),
        .dout(new_Jinkela_wire_2384)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_2440),
        .dout(new_Jinkela_wire_2441)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_2384),
        .dout(new_Jinkela_wire_2385)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_2487),
        .dout(new_Jinkela_wire_2488)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_2385),
        .dout(new_Jinkela_wire_2386)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_2441),
        .dout(new_Jinkela_wire_2442)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_2386),
        .dout(new_Jinkela_wire_2387)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_2471),
        .dout(new_Jinkela_wire_2472)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_2387),
        .dout(new_Jinkela_wire_2388)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(new_Jinkela_wire_2442),
        .dout(new_Jinkela_wire_2443)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_2388),
        .dout(new_Jinkela_wire_2389)
    );

    bfr new_Jinkela_buffer_1694 (
        .din(_1762_),
        .dout(new_Jinkela_wire_2594)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_2389),
        .dout(new_Jinkela_wire_2390)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(new_Jinkela_wire_2443),
        .dout(new_Jinkela_wire_2444)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_2390),
        .dout(new_Jinkela_wire_2391)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(new_Jinkela_wire_2472),
        .dout(new_Jinkela_wire_2473)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_2391),
        .dout(new_Jinkela_wire_2392)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_2444),
        .dout(new_Jinkela_wire_2445)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_2392),
        .dout(new_Jinkela_wire_2393)
    );

    bfr new_Jinkela_buffer_8629 (
        .din(new_Jinkela_wire_10592),
        .dout(new_Jinkela_wire_10593)
    );

    bfr new_Jinkela_buffer_8544 (
        .din(new_Jinkela_wire_10495),
        .dout(new_Jinkela_wire_10496)
    );

    bfr new_Jinkela_buffer_8654 (
        .din(new_Jinkela_wire_10621),
        .dout(new_Jinkela_wire_10622)
    );

    bfr new_Jinkela_buffer_8545 (
        .din(new_Jinkela_wire_10496),
        .dout(new_Jinkela_wire_10497)
    );

    bfr new_Jinkela_buffer_8630 (
        .din(new_Jinkela_wire_10593),
        .dout(new_Jinkela_wire_10594)
    );

    bfr new_Jinkela_buffer_8546 (
        .din(new_Jinkela_wire_10497),
        .dout(new_Jinkela_wire_10498)
    );

    spl2 new_Jinkela_splitter_837 (
        .a(_0960_),
        .b(new_Jinkela_wire_10684),
        .c(new_Jinkela_wire_10685)
    );

    bfr new_Jinkela_buffer_8547 (
        .din(new_Jinkela_wire_10498),
        .dout(new_Jinkela_wire_10499)
    );

    bfr new_Jinkela_buffer_8631 (
        .din(new_Jinkela_wire_10594),
        .dout(new_Jinkela_wire_10595)
    );

    bfr new_Jinkela_buffer_8548 (
        .din(new_Jinkela_wire_10499),
        .dout(new_Jinkela_wire_10500)
    );

    bfr new_Jinkela_buffer_8655 (
        .din(new_Jinkela_wire_10622),
        .dout(new_Jinkela_wire_10623)
    );

    bfr new_Jinkela_buffer_8549 (
        .din(new_Jinkela_wire_10500),
        .dout(new_Jinkela_wire_10501)
    );

    bfr new_Jinkela_buffer_8632 (
        .din(new_Jinkela_wire_10595),
        .dout(new_Jinkela_wire_10596)
    );

    bfr new_Jinkela_buffer_8550 (
        .din(new_Jinkela_wire_10501),
        .dout(new_Jinkela_wire_10502)
    );

    bfr new_Jinkela_buffer_8551 (
        .din(new_Jinkela_wire_10502),
        .dout(new_Jinkela_wire_10503)
    );

    bfr new_Jinkela_buffer_8633 (
        .din(new_Jinkela_wire_10596),
        .dout(new_Jinkela_wire_10597)
    );

    bfr new_Jinkela_buffer_8552 (
        .din(new_Jinkela_wire_10503),
        .dout(new_Jinkela_wire_10504)
    );

    bfr new_Jinkela_buffer_8656 (
        .din(new_Jinkela_wire_10623),
        .dout(new_Jinkela_wire_10624)
    );

    bfr new_Jinkela_buffer_8553 (
        .din(new_Jinkela_wire_10504),
        .dout(new_Jinkela_wire_10505)
    );

    bfr new_Jinkela_buffer_8634 (
        .din(new_Jinkela_wire_10597),
        .dout(new_Jinkela_wire_10598)
    );

    bfr new_Jinkela_buffer_8554 (
        .din(new_Jinkela_wire_10505),
        .dout(new_Jinkela_wire_10506)
    );

    spl2 new_Jinkela_splitter_838 (
        .a(_0788_),
        .b(new_Jinkela_wire_10686),
        .c(new_Jinkela_wire_10687)
    );

    bfr new_Jinkela_buffer_8555 (
        .din(new_Jinkela_wire_10506),
        .dout(new_Jinkela_wire_10507)
    );

    bfr new_Jinkela_buffer_8635 (
        .din(new_Jinkela_wire_10598),
        .dout(new_Jinkela_wire_10599)
    );

    bfr new_Jinkela_buffer_8556 (
        .din(new_Jinkela_wire_10507),
        .dout(new_Jinkela_wire_10508)
    );

    bfr new_Jinkela_buffer_8657 (
        .din(new_Jinkela_wire_10624),
        .dout(new_Jinkela_wire_10625)
    );

    bfr new_Jinkela_buffer_8557 (
        .din(new_Jinkela_wire_10508),
        .dout(new_Jinkela_wire_10509)
    );

    bfr new_Jinkela_buffer_8636 (
        .din(new_Jinkela_wire_10599),
        .dout(new_Jinkela_wire_10600)
    );

    bfr new_Jinkela_buffer_8558 (
        .din(new_Jinkela_wire_10509),
        .dout(new_Jinkela_wire_10510)
    );

    spl2 new_Jinkela_splitter_839 (
        .a(_0722_),
        .b(new_Jinkela_wire_10692),
        .c(new_Jinkela_wire_10693)
    );

    bfr new_Jinkela_buffer_8559 (
        .din(new_Jinkela_wire_10510),
        .dout(new_Jinkela_wire_10511)
    );

    bfr new_Jinkela_buffer_8637 (
        .din(new_Jinkela_wire_10600),
        .dout(new_Jinkela_wire_10601)
    );

    bfr new_Jinkela_buffer_8560 (
        .din(new_Jinkela_wire_10511),
        .dout(new_Jinkela_wire_10512)
    );

    bfr new_Jinkela_buffer_8658 (
        .din(new_Jinkela_wire_10625),
        .dout(new_Jinkela_wire_10626)
    );

    bfr new_Jinkela_buffer_8561 (
        .din(new_Jinkela_wire_10512),
        .dout(new_Jinkela_wire_10513)
    );

    bfr new_Jinkela_buffer_8638 (
        .din(new_Jinkela_wire_10601),
        .dout(new_Jinkela_wire_10602)
    );

    bfr new_Jinkela_buffer_8562 (
        .din(new_Jinkela_wire_10513),
        .dout(new_Jinkela_wire_10514)
    );

    bfr new_Jinkela_buffer_8708 (
        .din(new_Jinkela_wire_10687),
        .dout(new_Jinkela_wire_10688)
    );

    bfr new_Jinkela_buffer_8712 (
        .din(_0574_),
        .dout(new_Jinkela_wire_10694)
    );

    bfr new_Jinkela_buffer_8563 (
        .din(new_Jinkela_wire_10514),
        .dout(new_Jinkela_wire_10515)
    );

    bfr new_Jinkela_buffer_8639 (
        .din(new_Jinkela_wire_10602),
        .dout(new_Jinkela_wire_10603)
    );

    bfr new_Jinkela_buffer_8564 (
        .din(new_Jinkela_wire_10515),
        .dout(new_Jinkela_wire_10516)
    );

    bfr new_Jinkela_buffer_15471 (
        .din(new_Jinkela_wire_18437),
        .dout(new_Jinkela_wire_18438)
    );

    and_ii _2665_ (
        .a(new_Jinkela_wire_2117),
        .b(new_Jinkela_wire_17654),
        .c(_1722_)
    );

    bfr new_Jinkela_buffer_15497 (
        .din(new_Jinkela_wire_18469),
        .dout(new_Jinkela_wire_18470)
    );

    and_bb _2666_ (
        .a(new_Jinkela_wire_2118),
        .b(new_Jinkela_wire_17655),
        .c(_1723_)
    );

    bfr new_Jinkela_buffer_15472 (
        .din(new_Jinkela_wire_18438),
        .dout(new_Jinkela_wire_18439)
    );

    or_bb _2667_ (
        .a(new_Jinkela_wire_7583),
        .b(new_Jinkela_wire_19065),
        .c(_1724_)
    );

    bfr new_Jinkela_buffer_15529 (
        .din(new_Jinkela_wire_18503),
        .dout(new_Jinkela_wire_18504)
    );

    or_bb _2668_ (
        .a(new_Jinkela_wire_7440),
        .b(new_Jinkela_wire_20287),
        .c(_1725_)
    );

    bfr new_Jinkela_buffer_15473 (
        .din(new_Jinkela_wire_18439),
        .dout(new_Jinkela_wire_18440)
    );

    or_ii _2669_ (
        .a(new_Jinkela_wire_7441),
        .b(new_Jinkela_wire_20288),
        .c(_1726_)
    );

    bfr new_Jinkela_buffer_15498 (
        .din(new_Jinkela_wire_18470),
        .dout(new_Jinkela_wire_18471)
    );

    or_ii _2670_ (
        .a(new_Jinkela_wire_16368),
        .b(new_Jinkela_wire_17056),
        .c(_1727_)
    );

    bfr new_Jinkela_buffer_15474 (
        .din(new_Jinkela_wire_18440),
        .dout(new_Jinkela_wire_18441)
    );

    and_ii _2671_ (
        .a(new_Jinkela_wire_12339),
        .b(new_Jinkela_wire_4567),
        .c(_1728_)
    );

    bfr new_Jinkela_buffer_15547 (
        .din(_0516_),
        .dout(new_Jinkela_wire_18534)
    );

    and_bb _2672_ (
        .a(new_Jinkela_wire_12340),
        .b(new_Jinkela_wire_4568),
        .c(_1729_)
    );

    bfr new_Jinkela_buffer_15475 (
        .din(new_Jinkela_wire_18441),
        .dout(new_Jinkela_wire_18442)
    );

    or_bb _2673_ (
        .a(new_Jinkela_wire_13410),
        .b(new_Jinkela_wire_16779),
        .c(_1731_)
    );

    bfr new_Jinkela_buffer_15499 (
        .din(new_Jinkela_wire_18471),
        .dout(new_Jinkela_wire_18472)
    );

    or_bb _2674_ (
        .a(new_Jinkela_wire_6202),
        .b(new_Jinkela_wire_16947),
        .c(_1732_)
    );

    spl2 new_Jinkela_splitter_1332 (
        .a(new_Jinkela_wire_18442),
        .b(new_Jinkela_wire_18443),
        .c(new_Jinkela_wire_18444)
    );

    or_ii _2675_ (
        .a(new_Jinkela_wire_6203),
        .b(new_Jinkela_wire_16948),
        .c(_1733_)
    );

    bfr new_Jinkela_buffer_15500 (
        .din(new_Jinkela_wire_18472),
        .dout(new_Jinkela_wire_18473)
    );

    or_ii _2676_ (
        .a(new_Jinkela_wire_20047),
        .b(new_Jinkela_wire_20349),
        .c(_1734_)
    );

    bfr new_Jinkela_buffer_15530 (
        .din(new_Jinkela_wire_18504),
        .dout(new_Jinkela_wire_18505)
    );

    and_ii _2677_ (
        .a(new_Jinkela_wire_4834),
        .b(new_Jinkela_wire_17355),
        .c(_1735_)
    );

    and_bb _2678_ (
        .a(new_Jinkela_wire_4835),
        .b(new_Jinkela_wire_17356),
        .c(_1736_)
    );

    bfr new_Jinkela_buffer_15545 (
        .din(_0561_),
        .dout(new_Jinkela_wire_18532)
    );

    bfr new_Jinkela_buffer_15501 (
        .din(new_Jinkela_wire_18473),
        .dout(new_Jinkela_wire_18474)
    );

    or_bb _2679_ (
        .a(new_Jinkela_wire_16776),
        .b(new_Jinkela_wire_11529),
        .c(_1737_)
    );

    bfr new_Jinkela_buffer_15531 (
        .din(new_Jinkela_wire_18505),
        .dout(new_Jinkela_wire_18506)
    );

    or_bb _2680_ (
        .a(new_Jinkela_wire_13012),
        .b(new_Jinkela_wire_17071),
        .c(_1738_)
    );

    bfr new_Jinkela_buffer_15502 (
        .din(new_Jinkela_wire_18474),
        .dout(new_Jinkela_wire_18475)
    );

    or_ii _2681_ (
        .a(new_Jinkela_wire_13013),
        .b(new_Jinkela_wire_17072),
        .c(_1739_)
    );

    or_ii _2682_ (
        .a(new_Jinkela_wire_9520),
        .b(new_Jinkela_wire_19276),
        .c(_1740_)
    );

    bfr new_Jinkela_buffer_15546 (
        .din(_0782_),
        .dout(new_Jinkela_wire_18533)
    );

    bfr new_Jinkela_buffer_15503 (
        .din(new_Jinkela_wire_18475),
        .dout(new_Jinkela_wire_18476)
    );

    and_ii _2683_ (
        .a(new_Jinkela_wire_14692),
        .b(new_Jinkela_wire_19781),
        .c(_1742_)
    );

    bfr new_Jinkela_buffer_15532 (
        .din(new_Jinkela_wire_18506),
        .dout(new_Jinkela_wire_18507)
    );

    and_bb _2684_ (
        .a(new_Jinkela_wire_14693),
        .b(new_Jinkela_wire_19782),
        .c(_1743_)
    );

    bfr new_Jinkela_buffer_15504 (
        .din(new_Jinkela_wire_18476),
        .dout(new_Jinkela_wire_18477)
    );

    or_bb _2685_ (
        .a(new_Jinkela_wire_16205),
        .b(new_Jinkela_wire_21097),
        .c(_1744_)
    );

    or_bb _2686_ (
        .a(new_Jinkela_wire_4903),
        .b(new_Jinkela_wire_5993),
        .c(_1745_)
    );

    spl2 new_Jinkela_splitter_1342 (
        .a(_1174_),
        .b(new_Jinkela_wire_18535),
        .c(new_Jinkela_wire_18536)
    );

    bfr new_Jinkela_buffer_15505 (
        .din(new_Jinkela_wire_18477),
        .dout(new_Jinkela_wire_18478)
    );

    or_ii _2687_ (
        .a(new_Jinkela_wire_4904),
        .b(new_Jinkela_wire_5994),
        .c(_1746_)
    );

    bfr new_Jinkela_buffer_15533 (
        .din(new_Jinkela_wire_18507),
        .dout(new_Jinkela_wire_18508)
    );

    or_ii _2688_ (
        .a(new_Jinkela_wire_4247),
        .b(new_Jinkela_wire_7506),
        .c(_1747_)
    );

    bfr new_Jinkela_buffer_15506 (
        .din(new_Jinkela_wire_18478),
        .dout(new_Jinkela_wire_18479)
    );

    and_ii _2689_ (
        .a(new_Jinkela_wire_1134),
        .b(new_Jinkela_wire_10255),
        .c(_1748_)
    );

    spl2 new_Jinkela_splitter_1343 (
        .a(_0689_),
        .b(new_Jinkela_wire_18537),
        .c(new_Jinkela_wire_18538)
    );

    and_bb _2690_ (
        .a(new_Jinkela_wire_1135),
        .b(new_Jinkela_wire_10256),
        .c(_1749_)
    );

    bfr new_Jinkela_buffer_15507 (
        .din(new_Jinkela_wire_18479),
        .dout(new_Jinkela_wire_18480)
    );

    or_bb _2691_ (
        .a(new_Jinkela_wire_1626),
        .b(new_Jinkela_wire_1267),
        .c(_1750_)
    );

    bfr new_Jinkela_buffer_15534 (
        .din(new_Jinkela_wire_18508),
        .dout(new_Jinkela_wire_18509)
    );

    or_bb _2692_ (
        .a(new_Jinkela_wire_16700),
        .b(new_Jinkela_wire_4083),
        .c(_1751_)
    );

    bfr new_Jinkela_buffer_15508 (
        .din(new_Jinkela_wire_18480),
        .dout(new_Jinkela_wire_18481)
    );

    or_ii _2693_ (
        .a(new_Jinkela_wire_16701),
        .b(new_Jinkela_wire_4084),
        .c(_1753_)
    );

    or_ii _2694_ (
        .a(new_Jinkela_wire_6854),
        .b(new_Jinkela_wire_11830),
        .c(_1754_)
    );

    bfr new_Jinkela_buffer_15509 (
        .din(new_Jinkela_wire_18481),
        .dout(new_Jinkela_wire_18482)
    );

    and_ii _2695_ (
        .a(new_Jinkela_wire_19788),
        .b(new_Jinkela_wire_17973),
        .c(_1755_)
    );

    bfr new_Jinkela_buffer_15535 (
        .din(new_Jinkela_wire_18509),
        .dout(new_Jinkela_wire_18510)
    );

    and_bb _2696_ (
        .a(new_Jinkela_wire_19789),
        .b(new_Jinkela_wire_17974),
        .c(_1756_)
    );

    bfr new_Jinkela_buffer_15510 (
        .din(new_Jinkela_wire_18482),
        .dout(new_Jinkela_wire_18483)
    );

    or_bb _2697_ (
        .a(new_Jinkela_wire_4913),
        .b(new_Jinkela_wire_12739),
        .c(_1757_)
    );

    or_bb _2698_ (
        .a(new_Jinkela_wire_14656),
        .b(new_Jinkela_wire_8295),
        .c(_1758_)
    );

    bfr new_Jinkela_buffer_15572 (
        .din(_1412_),
        .dout(new_Jinkela_wire_18563)
    );

    bfr new_Jinkela_buffer_15511 (
        .din(new_Jinkela_wire_18483),
        .dout(new_Jinkela_wire_18484)
    );

    or_ii _2699_ (
        .a(new_Jinkela_wire_14657),
        .b(new_Jinkela_wire_8296),
        .c(_1759_)
    );

    bfr new_Jinkela_buffer_15536 (
        .din(new_Jinkela_wire_18510),
        .dout(new_Jinkela_wire_18511)
    );

    or_ii _2700_ (
        .a(new_Jinkela_wire_19918),
        .b(new_Jinkela_wire_19150),
        .c(_1760_)
    );

    bfr new_Jinkela_buffer_15512 (
        .din(new_Jinkela_wire_18484),
        .dout(new_Jinkela_wire_18485)
    );

    and_ii _2701_ (
        .a(new_Jinkela_wire_6846),
        .b(new_Jinkela_wire_9171),
        .c(_1761_)
    );

    bfr new_Jinkela_buffer_15548 (
        .din(new_Jinkela_wire_18538),
        .dout(new_Jinkela_wire_18539)
    );

    and_bb _2702_ (
        .a(new_Jinkela_wire_6847),
        .b(new_Jinkela_wire_9172),
        .c(_1762_)
    );

    spl2 new_Jinkela_splitter_1344 (
        .a(_1679_),
        .b(new_Jinkela_wire_18564),
        .c(new_Jinkela_wire_18565)
    );

    bfr new_Jinkela_buffer_15513 (
        .din(new_Jinkela_wire_18485),
        .dout(new_Jinkela_wire_18486)
    );

    or_bb _2703_ (
        .a(new_Jinkela_wire_2594),
        .b(new_Jinkela_wire_21110),
        .c(_1764_)
    );

    bfr new_Jinkela_buffer_15537 (
        .din(new_Jinkela_wire_18511),
        .dout(new_Jinkela_wire_18512)
    );

    or_bb _2704_ (
        .a(new_Jinkela_wire_17545),
        .b(new_Jinkela_wire_3116),
        .c(_1765_)
    );

    bfr new_Jinkela_buffer_15514 (
        .din(new_Jinkela_wire_18486),
        .dout(new_Jinkela_wire_18487)
    );

    or_ii _2705_ (
        .a(new_Jinkela_wire_17546),
        .b(new_Jinkela_wire_3117),
        .c(_1766_)
    );

    spl2 new_Jinkela_splitter_1345 (
        .a(_0045_),
        .b(new_Jinkela_wire_18566),
        .c(new_Jinkela_wire_18567)
    );

    or_ii _2706_ (
        .a(new_Jinkela_wire_17015),
        .b(new_Jinkela_wire_16783),
        .c(_1767_)
    );

    bfr new_Jinkela_buffer_12010 (
        .din(new_Jinkela_wire_14483),
        .dout(new_Jinkela_wire_14484)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_2488),
        .dout(new_Jinkela_wire_2489)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_2393),
        .dout(new_Jinkela_wire_2394)
    );

    bfr new_Jinkela_buffer_12091 (
        .din(new_Jinkela_wire_14568),
        .dout(new_Jinkela_wire_14569)
    );

    bfr new_Jinkela_buffer_12011 (
        .din(new_Jinkela_wire_14484),
        .dout(new_Jinkela_wire_14485)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_2445),
        .dout(new_Jinkela_wire_2446)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_2394),
        .dout(new_Jinkela_wire_2395)
    );

    bfr new_Jinkela_buffer_12012 (
        .din(new_Jinkela_wire_14485),
        .dout(new_Jinkela_wire_14486)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_Jinkela_wire_2473),
        .dout(new_Jinkela_wire_2474)
    );

    spl2 new_Jinkela_splitter_1097 (
        .a(_1740_),
        .b(new_Jinkela_wire_14692),
        .c(new_Jinkela_wire_14693)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_2395),
        .dout(new_Jinkela_wire_2396)
    );

    bfr new_Jinkela_buffer_12092 (
        .din(new_Jinkela_wire_14569),
        .dout(new_Jinkela_wire_14570)
    );

    bfr new_Jinkela_buffer_12013 (
        .din(new_Jinkela_wire_14486),
        .dout(new_Jinkela_wire_14487)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_2446),
        .dout(new_Jinkela_wire_2447)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(new_Jinkela_wire_2396),
        .dout(new_Jinkela_wire_2397)
    );

    bfr new_Jinkela_buffer_12115 (
        .din(new_Jinkela_wire_14592),
        .dout(new_Jinkela_wire_14593)
    );

    bfr new_Jinkela_buffer_12014 (
        .din(new_Jinkela_wire_14487),
        .dout(new_Jinkela_wire_14488)
    );

    bfr new_Jinkela_buffer_1695 (
        .din(_1524_),
        .dout(new_Jinkela_wire_2597)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_2397),
        .dout(new_Jinkela_wire_2398)
    );

    bfr new_Jinkela_buffer_12093 (
        .din(new_Jinkela_wire_14570),
        .dout(new_Jinkela_wire_14571)
    );

    bfr new_Jinkela_buffer_12015 (
        .din(new_Jinkela_wire_14488),
        .dout(new_Jinkela_wire_14489)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(new_Jinkela_wire_2447),
        .dout(new_Jinkela_wire_2448)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_2398),
        .dout(new_Jinkela_wire_2399)
    );

    bfr new_Jinkela_buffer_12016 (
        .din(new_Jinkela_wire_14489),
        .dout(new_Jinkela_wire_14490)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_Jinkela_wire_2474),
        .dout(new_Jinkela_wire_2475)
    );

    bfr new_Jinkela_buffer_12183 (
        .din(new_Jinkela_wire_14668),
        .dout(new_Jinkela_wire_14669)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_2399),
        .dout(new_Jinkela_wire_2400)
    );

    bfr new_Jinkela_buffer_12094 (
        .din(new_Jinkela_wire_14571),
        .dout(new_Jinkela_wire_14572)
    );

    bfr new_Jinkela_buffer_12017 (
        .din(new_Jinkela_wire_14490),
        .dout(new_Jinkela_wire_14491)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_2448),
        .dout(new_Jinkela_wire_2449)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_2400),
        .dout(new_Jinkela_wire_2401)
    );

    bfr new_Jinkela_buffer_12116 (
        .din(new_Jinkela_wire_14593),
        .dout(new_Jinkela_wire_14594)
    );

    bfr new_Jinkela_buffer_12018 (
        .din(new_Jinkela_wire_14491),
        .dout(new_Jinkela_wire_14492)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_2489),
        .dout(new_Jinkela_wire_2490)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_2401),
        .dout(new_Jinkela_wire_2402)
    );

    bfr new_Jinkela_buffer_12095 (
        .din(new_Jinkela_wire_14572),
        .dout(new_Jinkela_wire_14573)
    );

    bfr new_Jinkela_buffer_12019 (
        .din(new_Jinkela_wire_14492),
        .dout(new_Jinkela_wire_14493)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(new_Jinkela_wire_2449),
        .dout(new_Jinkela_wire_2450)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_2402),
        .dout(new_Jinkela_wire_2403)
    );

    bfr new_Jinkela_buffer_12020 (
        .din(new_Jinkela_wire_14493),
        .dout(new_Jinkela_wire_14494)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_2475),
        .dout(new_Jinkela_wire_2476)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_2403),
        .dout(new_Jinkela_wire_2404)
    );

    bfr new_Jinkela_buffer_12096 (
        .din(new_Jinkela_wire_14573),
        .dout(new_Jinkela_wire_14574)
    );

    bfr new_Jinkela_buffer_12021 (
        .din(new_Jinkela_wire_14494),
        .dout(new_Jinkela_wire_14495)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_2450),
        .dout(new_Jinkela_wire_2451)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(new_Jinkela_wire_2404),
        .dout(new_Jinkela_wire_2405)
    );

    bfr new_Jinkela_buffer_12117 (
        .din(new_Jinkela_wire_14594),
        .dout(new_Jinkela_wire_14595)
    );

    bfr new_Jinkela_buffer_12022 (
        .din(new_Jinkela_wire_14495),
        .dout(new_Jinkela_wire_14496)
    );

    spl2 new_Jinkela_splitter_299 (
        .a(_0381_),
        .b(new_Jinkela_wire_2595),
        .c(new_Jinkela_wire_2596)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(new_Jinkela_wire_2405),
        .dout(new_Jinkela_wire_2406)
    );

    bfr new_Jinkela_buffer_12097 (
        .din(new_Jinkela_wire_14574),
        .dout(new_Jinkela_wire_14575)
    );

    bfr new_Jinkela_buffer_12023 (
        .din(new_Jinkela_wire_14496),
        .dout(new_Jinkela_wire_14497)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(new_Jinkela_wire_2451),
        .dout(new_Jinkela_wire_2452)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(new_Jinkela_wire_2406),
        .dout(new_Jinkela_wire_2407)
    );

    spl2 new_Jinkela_splitter_1096 (
        .a(_1291_),
        .b(new_Jinkela_wire_14690),
        .c(new_Jinkela_wire_14691)
    );

    bfr new_Jinkela_buffer_12024 (
        .din(new_Jinkela_wire_14497),
        .dout(new_Jinkela_wire_14498)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_2476),
        .dout(new_Jinkela_wire_2477)
    );

    bfr new_Jinkela_buffer_12184 (
        .din(new_Jinkela_wire_14669),
        .dout(new_Jinkela_wire_14670)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(new_Jinkela_wire_2407),
        .dout(new_Jinkela_wire_2408)
    );

    bfr new_Jinkela_buffer_12098 (
        .din(new_Jinkela_wire_14575),
        .dout(new_Jinkela_wire_14576)
    );

    bfr new_Jinkela_buffer_12025 (
        .din(new_Jinkela_wire_14498),
        .dout(new_Jinkela_wire_14499)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(new_Jinkela_wire_2452),
        .dout(new_Jinkela_wire_2453)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(new_Jinkela_wire_2408),
        .dout(new_Jinkela_wire_2409)
    );

    bfr new_Jinkela_buffer_12118 (
        .din(new_Jinkela_wire_14595),
        .dout(new_Jinkela_wire_14596)
    );

    bfr new_Jinkela_buffer_12026 (
        .din(new_Jinkela_wire_14499),
        .dout(new_Jinkela_wire_14500)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_2490),
        .dout(new_Jinkela_wire_2491)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(new_Jinkela_wire_2409),
        .dout(new_Jinkela_wire_2410)
    );

    bfr new_Jinkela_buffer_12099 (
        .din(new_Jinkela_wire_14576),
        .dout(new_Jinkela_wire_14577)
    );

    bfr new_Jinkela_buffer_12027 (
        .din(new_Jinkela_wire_14500),
        .dout(new_Jinkela_wire_14501)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_Jinkela_wire_2453),
        .dout(new_Jinkela_wire_2454)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_2410),
        .dout(new_Jinkela_wire_2411)
    );

    bfr new_Jinkela_buffer_12028 (
        .din(new_Jinkela_wire_14501),
        .dout(new_Jinkela_wire_14502)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_2477),
        .dout(new_Jinkela_wire_2478)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_2411),
        .dout(new_Jinkela_wire_2412)
    );

    bfr new_Jinkela_buffer_12100 (
        .din(new_Jinkela_wire_14577),
        .dout(new_Jinkela_wire_14578)
    );

    bfr new_Jinkela_buffer_12029 (
        .din(new_Jinkela_wire_14502),
        .dout(new_Jinkela_wire_14503)
    );

    spl2 new_Jinkela_splitter_290 (
        .a(new_Jinkela_wire_2454),
        .b(new_Jinkela_wire_2455),
        .c(new_Jinkela_wire_2456)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_2412),
        .dout(new_Jinkela_wire_2413)
    );

    bfr new_Jinkela_buffer_12119 (
        .din(new_Jinkela_wire_14596),
        .dout(new_Jinkela_wire_14597)
    );

    bfr new_Jinkela_buffer_12030 (
        .din(new_Jinkela_wire_14503),
        .dout(new_Jinkela_wire_14504)
    );

    spl2 new_Jinkela_splitter_300 (
        .a(_1649_),
        .b(new_Jinkela_wire_2598),
        .c(new_Jinkela_wire_2599)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(new_Jinkela_wire_2413),
        .dout(new_Jinkela_wire_2414)
    );

    bfr new_Jinkela_buffer_12101 (
        .din(new_Jinkela_wire_14578),
        .dout(new_Jinkela_wire_14579)
    );

    bfr new_Jinkela_buffer_8659 (
        .din(new_Jinkela_wire_10626),
        .dout(new_Jinkela_wire_10627)
    );

    bfr new_Jinkela_buffer_8565 (
        .din(new_Jinkela_wire_10516),
        .dout(new_Jinkela_wire_10517)
    );

    bfr new_Jinkela_buffer_8640 (
        .din(new_Jinkela_wire_10603),
        .dout(new_Jinkela_wire_10604)
    );

    bfr new_Jinkela_buffer_8566 (
        .din(new_Jinkela_wire_10517),
        .dout(new_Jinkela_wire_10518)
    );

    spl2 new_Jinkela_splitter_841 (
        .a(_0239_),
        .b(new_Jinkela_wire_10745),
        .c(new_Jinkela_wire_10746)
    );

    bfr new_Jinkela_buffer_8567 (
        .din(new_Jinkela_wire_10518),
        .dout(new_Jinkela_wire_10519)
    );

    bfr new_Jinkela_buffer_8641 (
        .din(new_Jinkela_wire_10604),
        .dout(new_Jinkela_wire_10605)
    );

    bfr new_Jinkela_buffer_8568 (
        .din(new_Jinkela_wire_10519),
        .dout(new_Jinkela_wire_10520)
    );

    bfr new_Jinkela_buffer_8660 (
        .din(new_Jinkela_wire_10627),
        .dout(new_Jinkela_wire_10628)
    );

    bfr new_Jinkela_buffer_8569 (
        .din(new_Jinkela_wire_10520),
        .dout(new_Jinkela_wire_10521)
    );

    bfr new_Jinkela_buffer_8642 (
        .din(new_Jinkela_wire_10605),
        .dout(new_Jinkela_wire_10606)
    );

    bfr new_Jinkela_buffer_8570 (
        .din(new_Jinkela_wire_10521),
        .dout(new_Jinkela_wire_10522)
    );

    bfr new_Jinkela_buffer_8709 (
        .din(new_Jinkela_wire_10688),
        .dout(new_Jinkela_wire_10689)
    );

    bfr new_Jinkela_buffer_8571 (
        .din(new_Jinkela_wire_10522),
        .dout(new_Jinkela_wire_10523)
    );

    bfr new_Jinkela_buffer_8643 (
        .din(new_Jinkela_wire_10606),
        .dout(new_Jinkela_wire_10607)
    );

    bfr new_Jinkela_buffer_8572 (
        .din(new_Jinkela_wire_10523),
        .dout(new_Jinkela_wire_10524)
    );

    bfr new_Jinkela_buffer_8661 (
        .din(new_Jinkela_wire_10628),
        .dout(new_Jinkela_wire_10629)
    );

    bfr new_Jinkela_buffer_8573 (
        .din(new_Jinkela_wire_10524),
        .dout(new_Jinkela_wire_10525)
    );

    bfr new_Jinkela_buffer_8644 (
        .din(new_Jinkela_wire_10607),
        .dout(new_Jinkela_wire_10608)
    );

    bfr new_Jinkela_buffer_8574 (
        .din(new_Jinkela_wire_10525),
        .dout(new_Jinkela_wire_10526)
    );

    bfr new_Jinkela_buffer_8713 (
        .din(_0102_),
        .dout(new_Jinkela_wire_10695)
    );

    bfr new_Jinkela_buffer_8575 (
        .din(new_Jinkela_wire_10526),
        .dout(new_Jinkela_wire_10527)
    );

    bfr new_Jinkela_buffer_8645 (
        .din(new_Jinkela_wire_10608),
        .dout(new_Jinkela_wire_10609)
    );

    bfr new_Jinkela_buffer_8576 (
        .din(new_Jinkela_wire_10527),
        .dout(new_Jinkela_wire_10528)
    );

    bfr new_Jinkela_buffer_8662 (
        .din(new_Jinkela_wire_10629),
        .dout(new_Jinkela_wire_10630)
    );

    bfr new_Jinkela_buffer_8577 (
        .din(new_Jinkela_wire_10528),
        .dout(new_Jinkela_wire_10529)
    );

    bfr new_Jinkela_buffer_8646 (
        .din(new_Jinkela_wire_10609),
        .dout(new_Jinkela_wire_10610)
    );

    bfr new_Jinkela_buffer_8578 (
        .din(new_Jinkela_wire_10529),
        .dout(new_Jinkela_wire_10530)
    );

    bfr new_Jinkela_buffer_8710 (
        .din(new_Jinkela_wire_10689),
        .dout(new_Jinkela_wire_10690)
    );

    bfr new_Jinkela_buffer_8579 (
        .din(new_Jinkela_wire_10530),
        .dout(new_Jinkela_wire_10531)
    );

    bfr new_Jinkela_buffer_8647 (
        .din(new_Jinkela_wire_10610),
        .dout(new_Jinkela_wire_10611)
    );

    bfr new_Jinkela_buffer_8580 (
        .din(new_Jinkela_wire_10531),
        .dout(new_Jinkela_wire_10532)
    );

    bfr new_Jinkela_buffer_8663 (
        .din(new_Jinkela_wire_10630),
        .dout(new_Jinkela_wire_10631)
    );

    bfr new_Jinkela_buffer_8581 (
        .din(new_Jinkela_wire_10532),
        .dout(new_Jinkela_wire_10533)
    );

    spl2 new_Jinkela_splitter_831 (
        .a(new_Jinkela_wire_10611),
        .b(new_Jinkela_wire_10612),
        .c(new_Jinkela_wire_10613)
    );

    bfr new_Jinkela_buffer_8582 (
        .din(new_Jinkela_wire_10533),
        .dout(new_Jinkela_wire_10534)
    );

    bfr new_Jinkela_buffer_8664 (
        .din(new_Jinkela_wire_10631),
        .dout(new_Jinkela_wire_10632)
    );

    bfr new_Jinkela_buffer_8583 (
        .din(new_Jinkela_wire_10534),
        .dout(new_Jinkela_wire_10535)
    );

    spl2 new_Jinkela_splitter_842 (
        .a(_0993_),
        .b(new_Jinkela_wire_10751),
        .c(new_Jinkela_wire_10752)
    );

    bfr new_Jinkela_buffer_8584 (
        .din(new_Jinkela_wire_10535),
        .dout(new_Jinkela_wire_10536)
    );

    bfr new_Jinkela_buffer_8711 (
        .din(new_Jinkela_wire_10690),
        .dout(new_Jinkela_wire_10691)
    );

    bfr new_Jinkela_buffer_8585 (
        .din(new_Jinkela_wire_10536),
        .dout(new_Jinkela_wire_10537)
    );

    bfr new_Jinkela_buffer_12031 (
        .din(new_Jinkela_wire_14504),
        .dout(new_Jinkela_wire_14505)
    );

    bfr new_Jinkela_buffer_5211 (
        .din(new_Jinkela_wire_6698),
        .dout(new_Jinkela_wire_6699)
    );

    bfr new_Jinkela_buffer_15515 (
        .din(new_Jinkela_wire_18487),
        .dout(new_Jinkela_wire_18488)
    );

    spl2 new_Jinkela_splitter_294 (
        .a(new_Jinkela_wire_2478),
        .b(new_Jinkela_wire_2479),
        .c(new_Jinkela_wire_2480)
    );

    bfr new_Jinkela_buffer_15538 (
        .din(new_Jinkela_wire_18512),
        .dout(new_Jinkela_wire_18513)
    );

    bfr new_Jinkela_buffer_5117 (
        .din(new_Jinkela_wire_6590),
        .dout(new_Jinkela_wire_6591)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_2414),
        .dout(new_Jinkela_wire_2415)
    );

    bfr new_Jinkela_buffer_12032 (
        .din(new_Jinkela_wire_14505),
        .dout(new_Jinkela_wire_14506)
    );

    bfr new_Jinkela_buffer_5169 (
        .din(new_Jinkela_wire_6646),
        .dout(new_Jinkela_wire_6647)
    );

    bfr new_Jinkela_buffer_15516 (
        .din(new_Jinkela_wire_18488),
        .dout(new_Jinkela_wire_18489)
    );

    bfr new_Jinkela_buffer_1696 (
        .din(_0125_),
        .dout(new_Jinkela_wire_2600)
    );

    bfr new_Jinkela_buffer_5118 (
        .din(new_Jinkela_wire_6591),
        .dout(new_Jinkela_wire_6592)
    );

    bfr new_Jinkela_buffer_1697 (
        .din(_1132_),
        .dout(new_Jinkela_wire_2603)
    );

    bfr new_Jinkela_buffer_12185 (
        .din(new_Jinkela_wire_14670),
        .dout(new_Jinkela_wire_14671)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_2415),
        .dout(new_Jinkela_wire_2416)
    );

    bfr new_Jinkela_buffer_12120 (
        .din(new_Jinkela_wire_14597),
        .dout(new_Jinkela_wire_14598)
    );

    bfr new_Jinkela_buffer_15549 (
        .din(new_Jinkela_wire_18539),
        .dout(new_Jinkela_wire_18540)
    );

    bfr new_Jinkela_buffer_15517 (
        .din(new_Jinkela_wire_18489),
        .dout(new_Jinkela_wire_18490)
    );

    bfr new_Jinkela_buffer_12033 (
        .din(new_Jinkela_wire_14506),
        .dout(new_Jinkela_wire_14507)
    );

    bfr new_Jinkela_buffer_1596 (
        .din(new_Jinkela_wire_2491),
        .dout(new_Jinkela_wire_2492)
    );

    spl2 new_Jinkela_splitter_1336 (
        .a(new_Jinkela_wire_18513),
        .b(new_Jinkela_wire_18514),
        .c(new_Jinkela_wire_18515)
    );

    bfr new_Jinkela_buffer_5119 (
        .din(new_Jinkela_wire_6592),
        .dout(new_Jinkela_wire_6593)
    );

    spl2 new_Jinkela_splitter_288 (
        .a(new_Jinkela_wire_2416),
        .b(new_Jinkela_wire_2417),
        .c(new_Jinkela_wire_2418)
    );

    bfr new_Jinkela_buffer_12034 (
        .din(new_Jinkela_wire_14507),
        .dout(new_Jinkela_wire_14508)
    );

    bfr new_Jinkela_buffer_5170 (
        .din(new_Jinkela_wire_6647),
        .dout(new_Jinkela_wire_6648)
    );

    bfr new_Jinkela_buffer_15518 (
        .din(new_Jinkela_wire_18490),
        .dout(new_Jinkela_wire_18491)
    );

    bfr new_Jinkela_buffer_12196 (
        .din(_0456_),
        .dout(new_Jinkela_wire_14694)
    );

    bfr new_Jinkela_buffer_5120 (
        .din(new_Jinkela_wire_6593),
        .dout(new_Jinkela_wire_6594)
    );

    bfr new_Jinkela_buffer_15550 (
        .din(new_Jinkela_wire_18540),
        .dout(new_Jinkela_wire_18541)
    );

    bfr new_Jinkela_buffer_1597 (
        .din(new_Jinkela_wire_2492),
        .dout(new_Jinkela_wire_2493)
    );

    bfr new_Jinkela_buffer_12121 (
        .din(new_Jinkela_wire_14598),
        .dout(new_Jinkela_wire_14599)
    );

    bfr new_Jinkela_buffer_12035 (
        .din(new_Jinkela_wire_14508),
        .dout(new_Jinkela_wire_14509)
    );

    bfr new_Jinkela_buffer_5212 (
        .din(new_Jinkela_wire_6699),
        .dout(new_Jinkela_wire_6700)
    );

    spl2 new_Jinkela_splitter_1335 (
        .a(new_Jinkela_wire_18491),
        .b(new_Jinkela_wire_18492),
        .c(new_Jinkela_wire_18493)
    );

    bfr new_Jinkela_buffer_1598 (
        .din(new_Jinkela_wire_2493),
        .dout(new_Jinkela_wire_2494)
    );

    bfr new_Jinkela_buffer_5121 (
        .din(new_Jinkela_wire_6594),
        .dout(new_Jinkela_wire_6595)
    );

    bfr new_Jinkela_buffer_12198 (
        .din(_1278_),
        .dout(new_Jinkela_wire_14696)
    );

    bfr new_Jinkela_buffer_15577 (
        .din(_0971_),
        .dout(new_Jinkela_wire_18572)
    );

    bfr new_Jinkela_buffer_5171 (
        .din(new_Jinkela_wire_6648),
        .dout(new_Jinkela_wire_6649)
    );

    spl2 new_Jinkela_splitter_301 (
        .a(_0360_),
        .b(new_Jinkela_wire_2601),
        .c(new_Jinkela_wire_2602)
    );

    bfr new_Jinkela_buffer_12036 (
        .din(new_Jinkela_wire_14509),
        .dout(new_Jinkela_wire_14510)
    );

    bfr new_Jinkela_buffer_1599 (
        .din(new_Jinkela_wire_2494),
        .dout(new_Jinkela_wire_2495)
    );

    bfr new_Jinkela_buffer_12186 (
        .din(new_Jinkela_wire_14671),
        .dout(new_Jinkela_wire_14672)
    );

    bfr new_Jinkela_buffer_5122 (
        .din(new_Jinkela_wire_6595),
        .dout(new_Jinkela_wire_6596)
    );

    bfr new_Jinkela_buffer_15551 (
        .din(new_Jinkela_wire_18541),
        .dout(new_Jinkela_wire_18542)
    );

    bfr new_Jinkela_buffer_1745 (
        .din(_0245_),
        .dout(new_Jinkela_wire_2655)
    );

    bfr new_Jinkela_buffer_12122 (
        .din(new_Jinkela_wire_14599),
        .dout(new_Jinkela_wire_14600)
    );

    bfr new_Jinkela_buffer_12037 (
        .din(new_Jinkela_wire_14510),
        .dout(new_Jinkela_wire_14511)
    );

    bfr new_Jinkela_buffer_5249 (
        .din(new_Jinkela_wire_6740),
        .dout(new_Jinkela_wire_6741)
    );

    bfr new_Jinkela_buffer_15573 (
        .din(new_Jinkela_wire_18567),
        .dout(new_Jinkela_wire_18568)
    );

    bfr new_Jinkela_buffer_1600 (
        .din(new_Jinkela_wire_2495),
        .dout(new_Jinkela_wire_2496)
    );

    spl2 new_Jinkela_splitter_1346 (
        .a(_0515_),
        .b(new_Jinkela_wire_18573),
        .c(new_Jinkela_wire_18574)
    );

    bfr new_Jinkela_buffer_15552 (
        .din(new_Jinkela_wire_18542),
        .dout(new_Jinkela_wire_18543)
    );

    bfr new_Jinkela_buffer_5123 (
        .din(new_Jinkela_wire_6596),
        .dout(new_Jinkela_wire_6597)
    );

    bfr new_Jinkela_buffer_5172 (
        .din(new_Jinkela_wire_6649),
        .dout(new_Jinkela_wire_6650)
    );

    spl2 new_Jinkela_splitter_303 (
        .a(_0256_),
        .b(new_Jinkela_wire_2653),
        .c(new_Jinkela_wire_2654)
    );

    bfr new_Jinkela_buffer_12038 (
        .din(new_Jinkela_wire_14511),
        .dout(new_Jinkela_wire_14512)
    );

    bfr new_Jinkela_buffer_1601 (
        .din(new_Jinkela_wire_2496),
        .dout(new_Jinkela_wire_2497)
    );

    bfr new_Jinkela_buffer_15578 (
        .din(new_Jinkela_wire_18574),
        .dout(new_Jinkela_wire_18575)
    );

    bfr new_Jinkela_buffer_15582 (
        .din(_0846_),
        .dout(new_Jinkela_wire_18579)
    );

    bfr new_Jinkela_buffer_15553 (
        .din(new_Jinkela_wire_18543),
        .dout(new_Jinkela_wire_18544)
    );

    bfr new_Jinkela_buffer_5124 (
        .din(new_Jinkela_wire_6597),
        .dout(new_Jinkela_wire_6598)
    );

    bfr new_Jinkela_buffer_1698 (
        .din(new_Jinkela_wire_2603),
        .dout(new_Jinkela_wire_2604)
    );

    bfr new_Jinkela_buffer_12123 (
        .din(new_Jinkela_wire_14600),
        .dout(new_Jinkela_wire_14601)
    );

    bfr new_Jinkela_buffer_12039 (
        .din(new_Jinkela_wire_14512),
        .dout(new_Jinkela_wire_14513)
    );

    bfr new_Jinkela_buffer_5213 (
        .din(new_Jinkela_wire_6700),
        .dout(new_Jinkela_wire_6701)
    );

    bfr new_Jinkela_buffer_15574 (
        .din(new_Jinkela_wire_18568),
        .dout(new_Jinkela_wire_18569)
    );

    bfr new_Jinkela_buffer_1602 (
        .din(new_Jinkela_wire_2497),
        .dout(new_Jinkela_wire_2498)
    );

    bfr new_Jinkela_buffer_15554 (
        .din(new_Jinkela_wire_18544),
        .dout(new_Jinkela_wire_18545)
    );

    bfr new_Jinkela_buffer_5125 (
        .din(new_Jinkela_wire_6598),
        .dout(new_Jinkela_wire_6599)
    );

    spl2 new_Jinkela_splitter_306 (
        .a(_0375_),
        .b(new_Jinkela_wire_2711),
        .c(new_Jinkela_wire_2712)
    );

    bfr new_Jinkela_buffer_12197 (
        .din(_1494_),
        .dout(new_Jinkela_wire_14695)
    );

    bfr new_Jinkela_buffer_12040 (
        .din(new_Jinkela_wire_14513),
        .dout(new_Jinkela_wire_14514)
    );

    bfr new_Jinkela_buffer_5173 (
        .din(new_Jinkela_wire_6650),
        .dout(new_Jinkela_wire_6651)
    );

    bfr new_Jinkela_buffer_1603 (
        .din(new_Jinkela_wire_2498),
        .dout(new_Jinkela_wire_2499)
    );

    bfr new_Jinkela_buffer_12187 (
        .din(new_Jinkela_wire_14672),
        .dout(new_Jinkela_wire_14673)
    );

    bfr new_Jinkela_buffer_5126 (
        .din(new_Jinkela_wire_6599),
        .dout(new_Jinkela_wire_6600)
    );

    bfr new_Jinkela_buffer_15555 (
        .din(new_Jinkela_wire_18545),
        .dout(new_Jinkela_wire_18546)
    );

    bfr new_Jinkela_buffer_1699 (
        .din(new_Jinkela_wire_2604),
        .dout(new_Jinkela_wire_2605)
    );

    bfr new_Jinkela_buffer_12124 (
        .din(new_Jinkela_wire_14601),
        .dout(new_Jinkela_wire_14602)
    );

    bfr new_Jinkela_buffer_15575 (
        .din(new_Jinkela_wire_18569),
        .dout(new_Jinkela_wire_18570)
    );

    bfr new_Jinkela_buffer_12041 (
        .din(new_Jinkela_wire_14514),
        .dout(new_Jinkela_wire_14515)
    );

    bfr new_Jinkela_buffer_1604 (
        .din(new_Jinkela_wire_2499),
        .dout(new_Jinkela_wire_2500)
    );

    spl2 new_Jinkela_splitter_598 (
        .a(_1781_),
        .b(new_Jinkela_wire_6761),
        .c(new_Jinkela_wire_6762)
    );

    bfr new_Jinkela_buffer_15556 (
        .din(new_Jinkela_wire_18546),
        .dout(new_Jinkela_wire_18547)
    );

    bfr new_Jinkela_buffer_5127 (
        .din(new_Jinkela_wire_6600),
        .dout(new_Jinkela_wire_6601)
    );

    bfr new_Jinkela_buffer_1797 (
        .din(_1203_),
        .dout(new_Jinkela_wire_2713)
    );

    bfr new_Jinkela_buffer_5174 (
        .din(new_Jinkela_wire_6651),
        .dout(new_Jinkela_wire_6652)
    );

    bfr new_Jinkela_buffer_1749 (
        .din(_1819_),
        .dout(new_Jinkela_wire_2661)
    );

    bfr new_Jinkela_buffer_12042 (
        .din(new_Jinkela_wire_14515),
        .dout(new_Jinkela_wire_14516)
    );

    bfr new_Jinkela_buffer_1605 (
        .din(new_Jinkela_wire_2500),
        .dout(new_Jinkela_wire_2501)
    );

    bfr new_Jinkela_buffer_15586 (
        .din(new_net_3922),
        .dout(new_Jinkela_wire_18585)
    );

    bfr new_Jinkela_buffer_12278 (
        .din(_0617_),
        .dout(new_Jinkela_wire_14778)
    );

    bfr new_Jinkela_buffer_5128 (
        .din(new_Jinkela_wire_6601),
        .dout(new_Jinkela_wire_6602)
    );

    bfr new_Jinkela_buffer_15557 (
        .din(new_Jinkela_wire_18547),
        .dout(new_Jinkela_wire_18548)
    );

    bfr new_Jinkela_buffer_1700 (
        .din(new_Jinkela_wire_2605),
        .dout(new_Jinkela_wire_2606)
    );

    bfr new_Jinkela_buffer_12125 (
        .din(new_Jinkela_wire_14602),
        .dout(new_Jinkela_wire_14603)
    );

    bfr new_Jinkela_buffer_12043 (
        .din(new_Jinkela_wire_14516),
        .dout(new_Jinkela_wire_14517)
    );

    bfr new_Jinkela_buffer_5214 (
        .din(new_Jinkela_wire_6701),
        .dout(new_Jinkela_wire_6702)
    );

    bfr new_Jinkela_buffer_15576 (
        .din(new_Jinkela_wire_18570),
        .dout(new_Jinkela_wire_18571)
    );

    bfr new_Jinkela_buffer_1606 (
        .din(new_Jinkela_wire_2501),
        .dout(new_Jinkela_wire_2502)
    );

    bfr new_Jinkela_buffer_15558 (
        .din(new_Jinkela_wire_18548),
        .dout(new_Jinkela_wire_18549)
    );

    bfr new_Jinkela_buffer_5129 (
        .din(new_Jinkela_wire_6602),
        .dout(new_Jinkela_wire_6603)
    );

    bfr new_Jinkela_buffer_1746 (
        .din(new_Jinkela_wire_2655),
        .dout(new_Jinkela_wire_2656)
    );

    bfr new_Jinkela_buffer_12044 (
        .din(new_Jinkela_wire_14517),
        .dout(new_Jinkela_wire_14518)
    );

    bfr new_Jinkela_buffer_5175 (
        .din(new_Jinkela_wire_6652),
        .dout(new_Jinkela_wire_6653)
    );

    bfr new_Jinkela_buffer_15587 (
        .din(new_Jinkela_wire_18585),
        .dout(new_Jinkela_wire_18586)
    );

    bfr new_Jinkela_buffer_1607 (
        .din(new_Jinkela_wire_2502),
        .dout(new_Jinkela_wire_2503)
    );

    spl2 new_Jinkela_splitter_1348 (
        .a(_0749_),
        .b(new_Jinkela_wire_18685),
        .c(new_Jinkela_wire_18686)
    );

    bfr new_Jinkela_buffer_12188 (
        .din(new_Jinkela_wire_14673),
        .dout(new_Jinkela_wire_14674)
    );

    bfr new_Jinkela_buffer_5130 (
        .din(new_Jinkela_wire_6603),
        .dout(new_Jinkela_wire_6604)
    );

    bfr new_Jinkela_buffer_15559 (
        .din(new_Jinkela_wire_18549),
        .dout(new_Jinkela_wire_18550)
    );

    bfr new_Jinkela_buffer_1701 (
        .din(new_Jinkela_wire_2606),
        .dout(new_Jinkela_wire_2607)
    );

    bfr new_Jinkela_buffer_12126 (
        .din(new_Jinkela_wire_14603),
        .dout(new_Jinkela_wire_14604)
    );

    bfr new_Jinkela_buffer_12045 (
        .din(new_Jinkela_wire_14518),
        .dout(new_Jinkela_wire_14519)
    );

    bfr new_Jinkela_buffer_5250 (
        .din(new_Jinkela_wire_6741),
        .dout(new_Jinkela_wire_6742)
    );

    bfr new_Jinkela_buffer_15579 (
        .din(new_Jinkela_wire_18575),
        .dout(new_Jinkela_wire_18576)
    );

    bfr new_Jinkela_buffer_1608 (
        .din(new_Jinkela_wire_2503),
        .dout(new_Jinkela_wire_2504)
    );

    bfr new_Jinkela_buffer_15560 (
        .din(new_Jinkela_wire_18550),
        .dout(new_Jinkela_wire_18551)
    );

    bfr new_Jinkela_buffer_5131 (
        .din(new_Jinkela_wire_6604),
        .dout(new_Jinkela_wire_6605)
    );

    bfr new_Jinkela_buffer_5176 (
        .din(new_Jinkela_wire_6653),
        .dout(new_Jinkela_wire_6654)
    );

    bfr new_Jinkela_buffer_1747 (
        .din(new_Jinkela_wire_2656),
        .dout(new_Jinkela_wire_2657)
    );

    bfr new_Jinkela_buffer_12046 (
        .din(new_Jinkela_wire_14519),
        .dout(new_Jinkela_wire_14520)
    );

    bfr new_Jinkela_buffer_1609 (
        .din(new_Jinkela_wire_2504),
        .dout(new_Jinkela_wire_2505)
    );

    bfr new_Jinkela_buffer_15583 (
        .din(new_Jinkela_wire_18579),
        .dout(new_Jinkela_wire_18580)
    );

    bfr new_Jinkela_buffer_15561 (
        .din(new_Jinkela_wire_18551),
        .dout(new_Jinkela_wire_18552)
    );

    bfr new_Jinkela_buffer_5132 (
        .din(new_Jinkela_wire_6605),
        .dout(new_Jinkela_wire_6606)
    );

    bfr new_Jinkela_buffer_1702 (
        .din(new_Jinkela_wire_2607),
        .dout(new_Jinkela_wire_2608)
    );

    bfr new_Jinkela_buffer_12127 (
        .din(new_Jinkela_wire_14604),
        .dout(new_Jinkela_wire_14605)
    );

    bfr new_Jinkela_buffer_12047 (
        .din(new_Jinkela_wire_14520),
        .dout(new_Jinkela_wire_14521)
    );

    bfr new_Jinkela_buffer_5215 (
        .din(new_Jinkela_wire_6702),
        .dout(new_Jinkela_wire_6703)
    );

    bfr new_Jinkela_buffer_15580 (
        .din(new_Jinkela_wire_18576),
        .dout(new_Jinkela_wire_18577)
    );

    bfr new_Jinkela_buffer_1610 (
        .din(new_Jinkela_wire_2505),
        .dout(new_Jinkela_wire_2506)
    );

    bfr new_Jinkela_buffer_15562 (
        .din(new_Jinkela_wire_18552),
        .dout(new_Jinkela_wire_18553)
    );

    bfr new_Jinkela_buffer_5133 (
        .din(new_Jinkela_wire_6606),
        .dout(new_Jinkela_wire_6607)
    );

    bfr new_Jinkela_buffer_12390 (
        .din(_1682_),
        .dout(new_Jinkela_wire_14892)
    );

    bfr new_Jinkela_buffer_12048 (
        .din(new_Jinkela_wire_14521),
        .dout(new_Jinkela_wire_14522)
    );

    bfr new_Jinkela_buffer_5177 (
        .din(new_Jinkela_wire_6654),
        .dout(new_Jinkela_wire_6655)
    );

    bfr new_Jinkela_buffer_15686 (
        .din(_0382_),
        .dout(new_Jinkela_wire_18687)
    );

    bfr new_Jinkela_buffer_1611 (
        .din(new_Jinkela_wire_2506),
        .dout(new_Jinkela_wire_2507)
    );

    bfr new_Jinkela_buffer_15584 (
        .din(new_Jinkela_wire_18580),
        .dout(new_Jinkela_wire_18581)
    );

    bfr new_Jinkela_buffer_12189 (
        .din(new_Jinkela_wire_14674),
        .dout(new_Jinkela_wire_14675)
    );

    bfr new_Jinkela_buffer_5134 (
        .din(new_Jinkela_wire_6607),
        .dout(new_Jinkela_wire_6608)
    );

    bfr new_Jinkela_buffer_15563 (
        .din(new_Jinkela_wire_18553),
        .dout(new_Jinkela_wire_18554)
    );

    bfr new_Jinkela_buffer_1703 (
        .din(new_Jinkela_wire_2608),
        .dout(new_Jinkela_wire_2609)
    );

    bfr new_Jinkela_buffer_12128 (
        .din(new_Jinkela_wire_14605),
        .dout(new_Jinkela_wire_14606)
    );

    bfr new_Jinkela_buffer_12049 (
        .din(new_Jinkela_wire_14522),
        .dout(new_Jinkela_wire_14523)
    );

    spl2 new_Jinkela_splitter_601 (
        .a(_1511_),
        .b(new_Jinkela_wire_6768),
        .c(new_Jinkela_wire_6769)
    );

    bfr new_Jinkela_buffer_15581 (
        .din(new_Jinkela_wire_18577),
        .dout(new_Jinkela_wire_18578)
    );

    bfr new_Jinkela_buffer_1612 (
        .din(new_Jinkela_wire_2507),
        .dout(new_Jinkela_wire_2508)
    );

    spl2 new_Jinkela_splitter_599 (
        .a(_1654_),
        .b(new_Jinkela_wire_6763),
        .c(new_Jinkela_wire_6764)
    );

    bfr new_Jinkela_buffer_15564 (
        .din(new_Jinkela_wire_18554),
        .dout(new_Jinkela_wire_18555)
    );

    bfr new_Jinkela_buffer_5135 (
        .din(new_Jinkela_wire_6608),
        .dout(new_Jinkela_wire_6609)
    );

    bfr new_Jinkela_buffer_1750 (
        .din(new_Jinkela_wire_2661),
        .dout(new_Jinkela_wire_2662)
    );

    bfr new_Jinkela_buffer_12050 (
        .din(new_Jinkela_wire_14523),
        .dout(new_Jinkela_wire_14524)
    );

    bfr new_Jinkela_buffer_5178 (
        .din(new_Jinkela_wire_6655),
        .dout(new_Jinkela_wire_6656)
    );

    bfr new_Jinkela_buffer_1613 (
        .din(new_Jinkela_wire_2508),
        .dout(new_Jinkela_wire_2509)
    );

    bfr new_Jinkela_buffer_12199 (
        .din(new_Jinkela_wire_14696),
        .dout(new_Jinkela_wire_14697)
    );

    bfr new_Jinkela_buffer_5136 (
        .din(new_Jinkela_wire_6609),
        .dout(new_Jinkela_wire_6610)
    );

    bfr new_Jinkela_buffer_15565 (
        .din(new_Jinkela_wire_18555),
        .dout(new_Jinkela_wire_18556)
    );

    bfr new_Jinkela_buffer_1704 (
        .din(new_Jinkela_wire_2609),
        .dout(new_Jinkela_wire_2610)
    );

    bfr new_Jinkela_buffer_12129 (
        .din(new_Jinkela_wire_14606),
        .dout(new_Jinkela_wire_14607)
    );

    bfr new_Jinkela_buffer_12051 (
        .din(new_Jinkela_wire_14524),
        .dout(new_Jinkela_wire_14525)
    );

    bfr new_Jinkela_buffer_5216 (
        .din(new_Jinkela_wire_6703),
        .dout(new_Jinkela_wire_6704)
    );

    bfr new_Jinkela_buffer_1614 (
        .din(new_Jinkela_wire_2509),
        .dout(new_Jinkela_wire_2510)
    );

    bfr new_Jinkela_buffer_15566 (
        .din(new_Jinkela_wire_18556),
        .dout(new_Jinkela_wire_18557)
    );

    bfr new_Jinkela_buffer_5137 (
        .din(new_Jinkela_wire_6610),
        .dout(new_Jinkela_wire_6611)
    );

    bfr new_Jinkela_buffer_1748 (
        .din(new_Jinkela_wire_2657),
        .dout(new_Jinkela_wire_2658)
    );

    bfr new_Jinkela_buffer_8665 (
        .din(new_Jinkela_wire_10632),
        .dout(new_Jinkela_wire_10633)
    );

    and_ii _2707_ (
        .a(new_Jinkela_wire_4251),
        .b(new_Jinkela_wire_7259),
        .c(_1768_)
    );

    bfr new_Jinkela_buffer_8586 (
        .din(new_Jinkela_wire_10537),
        .dout(new_Jinkela_wire_10538)
    );

    and_bb _2708_ (
        .a(new_Jinkela_wire_4252),
        .b(new_Jinkela_wire_7260),
        .c(_1769_)
    );

    bfr new_Jinkela_buffer_8714 (
        .din(new_Jinkela_wire_10695),
        .dout(new_Jinkela_wire_10696)
    );

    or_bb _2709_ (
        .a(new_Jinkela_wire_3815),
        .b(new_Jinkela_wire_5463),
        .c(_1770_)
    );

    bfr new_Jinkela_buffer_8587 (
        .din(new_Jinkela_wire_10538),
        .dout(new_Jinkela_wire_10539)
    );

    or_bb _2710_ (
        .a(new_Jinkela_wire_13846),
        .b(new_Jinkela_wire_18953),
        .c(_1771_)
    );

    bfr new_Jinkela_buffer_8666 (
        .din(new_Jinkela_wire_10633),
        .dout(new_Jinkela_wire_10634)
    );

    or_ii _2711_ (
        .a(new_Jinkela_wire_13847),
        .b(new_Jinkela_wire_18954),
        .c(_1772_)
    );

    bfr new_Jinkela_buffer_8588 (
        .din(new_Jinkela_wire_10539),
        .dout(new_Jinkela_wire_10540)
    );

    or_ii _2712_ (
        .a(new_Jinkela_wire_7971),
        .b(new_Jinkela_wire_17675),
        .c(_1773_)
    );

    bfr new_Jinkela_buffer_8761 (
        .din(new_Jinkela_wire_10746),
        .dout(new_Jinkela_wire_10747)
    );

    and_ii _2713_ (
        .a(new_Jinkela_wire_13151),
        .b(new_Jinkela_wire_6093),
        .c(_1775_)
    );

    bfr new_Jinkela_buffer_8589 (
        .din(new_Jinkela_wire_10540),
        .dout(new_Jinkela_wire_10541)
    );

    and_bb _2714_ (
        .a(new_Jinkela_wire_13152),
        .b(new_Jinkela_wire_6094),
        .c(_1776_)
    );

    bfr new_Jinkela_buffer_8667 (
        .din(new_Jinkela_wire_10634),
        .dout(new_Jinkela_wire_10635)
    );

    or_bb _2715_ (
        .a(new_Jinkela_wire_21155),
        .b(new_Jinkela_wire_1387),
        .c(_1777_)
    );

    bfr new_Jinkela_buffer_8590 (
        .din(new_Jinkela_wire_10541),
        .dout(new_Jinkela_wire_10542)
    );

    or_bb _2716_ (
        .a(new_Jinkela_wire_11401),
        .b(new_Jinkela_wire_18979),
        .c(_1778_)
    );

    bfr new_Jinkela_buffer_8715 (
        .din(new_Jinkela_wire_10696),
        .dout(new_Jinkela_wire_10697)
    );

    or_ii _2717_ (
        .a(new_Jinkela_wire_11402),
        .b(new_Jinkela_wire_18980),
        .c(_1779_)
    );

    bfr new_Jinkela_buffer_8591 (
        .din(new_Jinkela_wire_10542),
        .dout(new_Jinkela_wire_10543)
    );

    or_ii _2718_ (
        .a(new_Jinkela_wire_19566),
        .b(new_Jinkela_wire_14090),
        .c(_1780_)
    );

    bfr new_Jinkela_buffer_8668 (
        .din(new_Jinkela_wire_10635),
        .dout(new_Jinkela_wire_10636)
    );

    and_ii _2719_ (
        .a(new_Jinkela_wire_18375),
        .b(new_Jinkela_wire_8961),
        .c(_1781_)
    );

    bfr new_Jinkela_buffer_8592 (
        .din(new_Jinkela_wire_10543),
        .dout(new_Jinkela_wire_10544)
    );

    and_bb _2720_ (
        .a(new_Jinkela_wire_18376),
        .b(new_Jinkela_wire_8962),
        .c(_1782_)
    );

    or_bb _2721_ (
        .a(new_Jinkela_wire_6679),
        .b(new_Jinkela_wire_6761),
        .c(_1783_)
    );

    bfr new_Jinkela_buffer_8765 (
        .din(_1567_),
        .dout(new_Jinkela_wire_10753)
    );

    bfr new_Jinkela_buffer_8593 (
        .din(new_Jinkela_wire_10544),
        .dout(new_Jinkela_wire_10545)
    );

    or_bb _2722_ (
        .a(new_Jinkela_wire_1283),
        .b(new_Jinkela_wire_11961),
        .c(_1784_)
    );

    bfr new_Jinkela_buffer_8669 (
        .din(new_Jinkela_wire_10636),
        .dout(new_Jinkela_wire_10637)
    );

    or_ii _2723_ (
        .a(new_Jinkela_wire_1284),
        .b(new_Jinkela_wire_11962),
        .c(_1786_)
    );

    bfr new_Jinkela_buffer_8594 (
        .din(new_Jinkela_wire_10545),
        .dout(new_Jinkela_wire_10546)
    );

    or_ii _2724_ (
        .a(new_Jinkela_wire_20385),
        .b(new_Jinkela_wire_7868),
        .c(_1787_)
    );

    bfr new_Jinkela_buffer_8716 (
        .din(new_Jinkela_wire_10697),
        .dout(new_Jinkela_wire_10698)
    );

    and_ii _2725_ (
        .a(new_Jinkela_wire_19960),
        .b(new_Jinkela_wire_14988),
        .c(_1788_)
    );

    bfr new_Jinkela_buffer_8595 (
        .din(new_Jinkela_wire_10546),
        .dout(new_Jinkela_wire_10547)
    );

    and_bb _2726_ (
        .a(new_Jinkela_wire_19961),
        .b(new_Jinkela_wire_14989),
        .c(_1789_)
    );

    bfr new_Jinkela_buffer_8670 (
        .din(new_Jinkela_wire_10637),
        .dout(new_Jinkela_wire_10638)
    );

    or_bb _2727_ (
        .a(new_Jinkela_wire_11838),
        .b(new_Jinkela_wire_7847),
        .c(_1790_)
    );

    bfr new_Jinkela_buffer_8596 (
        .din(new_Jinkela_wire_10547),
        .dout(new_Jinkela_wire_10548)
    );

    or_bb _2728_ (
        .a(new_Jinkela_wire_13154),
        .b(new_Jinkela_wire_2485),
        .c(_1791_)
    );

    bfr new_Jinkela_buffer_8845 (
        .din(_0696_),
        .dout(new_Jinkela_wire_10837)
    );

    or_ii _2729_ (
        .a(new_Jinkela_wire_13155),
        .b(new_Jinkela_wire_2486),
        .c(_1792_)
    );

    bfr new_Jinkela_buffer_8597 (
        .din(new_Jinkela_wire_10548),
        .dout(new_Jinkela_wire_10549)
    );

    or_ii _2730_ (
        .a(new_Jinkela_wire_2934),
        .b(new_Jinkela_wire_20388),
        .c(_1793_)
    );

    bfr new_Jinkela_buffer_8671 (
        .din(new_Jinkela_wire_10638),
        .dout(new_Jinkela_wire_10639)
    );

    and_ii _2731_ (
        .a(new_Jinkela_wire_6405),
        .b(new_Jinkela_wire_17530),
        .c(_1794_)
    );

    bfr new_Jinkela_buffer_8598 (
        .din(new_Jinkela_wire_10549),
        .dout(new_Jinkela_wire_10550)
    );

    and_bb _2732_ (
        .a(new_Jinkela_wire_6406),
        .b(new_Jinkela_wire_17531),
        .c(_1795_)
    );

    bfr new_Jinkela_buffer_8717 (
        .din(new_Jinkela_wire_10698),
        .dout(new_Jinkela_wire_10699)
    );

    or_bb _2733_ (
        .a(new_Jinkela_wire_7272),
        .b(new_Jinkela_wire_7734),
        .c(_1797_)
    );

    bfr new_Jinkela_buffer_8599 (
        .din(new_Jinkela_wire_10550),
        .dout(new_Jinkela_wire_10551)
    );

    and_ii _2734_ (
        .a(new_Jinkela_wire_15664),
        .b(new_Jinkela_wire_18564),
        .c(_1798_)
    );

    bfr new_Jinkela_buffer_8672 (
        .din(new_Jinkela_wire_10639),
        .dout(new_Jinkela_wire_10640)
    );

    and_bb _2735_ (
        .a(new_Jinkela_wire_15665),
        .b(new_Jinkela_wire_18565),
        .c(_1799_)
    );

    bfr new_Jinkela_buffer_8600 (
        .din(new_Jinkela_wire_10551),
        .dout(new_Jinkela_wire_10552)
    );

    or_bb _2736_ (
        .a(new_Jinkela_wire_16510),
        .b(new_Jinkela_wire_3952),
        .c(_1800_)
    );

    bfr new_Jinkela_buffer_8762 (
        .din(new_Jinkela_wire_10747),
        .dout(new_Jinkela_wire_10748)
    );

    and_ii _2737_ (
        .a(new_Jinkela_wire_17987),
        .b(new_Jinkela_wire_1252),
        .c(_1801_)
    );

    bfr new_Jinkela_buffer_8601 (
        .din(new_Jinkela_wire_10552),
        .dout(new_Jinkela_wire_10553)
    );

    and_bb _2738_ (
        .a(new_Jinkela_wire_17988),
        .b(new_Jinkela_wire_1253),
        .c(_1802_)
    );

    bfr new_Jinkela_buffer_8673 (
        .din(new_Jinkela_wire_10640),
        .dout(new_Jinkela_wire_10641)
    );

    or_bb _2739_ (
        .a(new_Jinkela_wire_13978),
        .b(new_Jinkela_wire_2145),
        .c(new_net_3920)
    );

    bfr new_Jinkela_buffer_8602 (
        .din(new_Jinkela_wire_10553),
        .dout(new_Jinkela_wire_10554)
    );

    and_bi _2740_ (
        .a(new_Jinkela_wire_20393),
        .b(new_Jinkela_wire_7735),
        .c(_1803_)
    );

    bfr new_Jinkela_buffer_8718 (
        .din(new_Jinkela_wire_10699),
        .dout(new_Jinkela_wire_10700)
    );

    and_bb _2741_ (
        .a(new_Jinkela_wire_523),
        .b(new_Jinkela_wire_559),
        .c(_1804_)
    );

    bfr new_Jinkela_buffer_8603 (
        .din(new_Jinkela_wire_10554),
        .dout(new_Jinkela_wire_10555)
    );

    and_bi _2742_ (
        .a(new_Jinkela_wire_7873),
        .b(new_Jinkela_wire_7848),
        .c(_1805_)
    );

    bfr new_Jinkela_buffer_8674 (
        .din(new_Jinkela_wire_10641),
        .dout(new_Jinkela_wire_10642)
    );

    and_bb _2743_ (
        .a(new_Jinkela_wire_271),
        .b(new_Jinkela_wire_138),
        .c(_1807_)
    );

    spl2 new_Jinkela_splitter_825 (
        .a(new_Jinkela_wire_10555),
        .b(new_Jinkela_wire_10556),
        .c(new_Jinkela_wire_10557)
    );

    and_bi _2744_ (
        .a(new_Jinkela_wire_14095),
        .b(new_Jinkela_wire_6762),
        .c(_1808_)
    );

    bfr new_Jinkela_buffer_8675 (
        .din(new_Jinkela_wire_10642),
        .dout(new_Jinkela_wire_10643)
    );

    and_bb _2745_ (
        .a(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_199),
        .c(_1809_)
    );

    and_bi _2746_ (
        .a(new_Jinkela_wire_17680),
        .b(new_Jinkela_wire_1388),
        .c(_1810_)
    );

    spl2 new_Jinkela_splitter_844 (
        .a(_1169_),
        .b(new_Jinkela_wire_10835),
        .c(new_Jinkela_wire_10836)
    );

    bfr new_Jinkela_buffer_8719 (
        .din(new_Jinkela_wire_10700),
        .dout(new_Jinkela_wire_10701)
    );

    and_bb _2747_ (
        .a(new_Jinkela_wire_479),
        .b(new_Jinkela_wire_576),
        .c(_1811_)
    );

    bfr new_Jinkela_buffer_8676 (
        .din(new_Jinkela_wire_10643),
        .dout(new_Jinkela_wire_10644)
    );

    and_bi _2748_ (
        .a(new_Jinkela_wire_16788),
        .b(new_Jinkela_wire_5464),
        .c(_1812_)
    );

    bfr new_Jinkela_buffer_5179 (
        .din(new_Jinkela_wire_6656),
        .dout(new_Jinkela_wire_6657)
    );

    bfr new_Jinkela_buffer_5138 (
        .din(new_Jinkela_wire_6611),
        .dout(new_Jinkela_wire_6612)
    );

    bfr new_Jinkela_buffer_5251 (
        .din(new_Jinkela_wire_6742),
        .dout(new_Jinkela_wire_6743)
    );

    bfr new_Jinkela_buffer_5139 (
        .din(new_Jinkela_wire_6612),
        .dout(new_Jinkela_wire_6613)
    );

    bfr new_Jinkela_buffer_5180 (
        .din(new_Jinkela_wire_6657),
        .dout(new_Jinkela_wire_6658)
    );

    bfr new_Jinkela_buffer_5140 (
        .din(new_Jinkela_wire_6613),
        .dout(new_Jinkela_wire_6614)
    );

    bfr new_Jinkela_buffer_5217 (
        .din(new_Jinkela_wire_6704),
        .dout(new_Jinkela_wire_6705)
    );

    spl2 new_Jinkela_splitter_586 (
        .a(new_Jinkela_wire_6614),
        .b(new_Jinkela_wire_6615),
        .c(new_Jinkela_wire_6616)
    );

    bfr new_Jinkela_buffer_5181 (
        .din(new_Jinkela_wire_6658),
        .dout(new_Jinkela_wire_6659)
    );

    bfr new_Jinkela_buffer_5182 (
        .din(new_Jinkela_wire_6659),
        .dout(new_Jinkela_wire_6660)
    );

    bfr new_Jinkela_buffer_5218 (
        .din(new_Jinkela_wire_6705),
        .dout(new_Jinkela_wire_6706)
    );

    bfr new_Jinkela_buffer_5183 (
        .din(new_Jinkela_wire_6660),
        .dout(new_Jinkela_wire_6661)
    );

    bfr new_Jinkela_buffer_5252 (
        .din(new_Jinkela_wire_6743),
        .dout(new_Jinkela_wire_6744)
    );

    bfr new_Jinkela_buffer_5184 (
        .din(new_Jinkela_wire_6661),
        .dout(new_Jinkela_wire_6662)
    );

    bfr new_Jinkela_buffer_5219 (
        .din(new_Jinkela_wire_6706),
        .dout(new_Jinkela_wire_6707)
    );

    bfr new_Jinkela_buffer_5185 (
        .din(new_Jinkela_wire_6662),
        .dout(new_Jinkela_wire_6663)
    );

    bfr new_Jinkela_buffer_5272 (
        .din(new_Jinkela_wire_6777),
        .dout(new_Jinkela_wire_6778)
    );

    spl2 new_Jinkela_splitter_609 (
        .a(_0966_),
        .b(new_Jinkela_wire_6848),
        .c(new_Jinkela_wire_6849)
    );

    bfr new_Jinkela_buffer_5186 (
        .din(new_Jinkela_wire_6663),
        .dout(new_Jinkela_wire_6664)
    );

    bfr new_Jinkela_buffer_5220 (
        .din(new_Jinkela_wire_6707),
        .dout(new_Jinkela_wire_6708)
    );

    bfr new_Jinkela_buffer_5187 (
        .din(new_Jinkela_wire_6664),
        .dout(new_Jinkela_wire_6665)
    );

    bfr new_Jinkela_buffer_5253 (
        .din(new_Jinkela_wire_6744),
        .dout(new_Jinkela_wire_6745)
    );

    bfr new_Jinkela_buffer_5188 (
        .din(new_Jinkela_wire_6665),
        .dout(new_Jinkela_wire_6666)
    );

    bfr new_Jinkela_buffer_5221 (
        .din(new_Jinkela_wire_6708),
        .dout(new_Jinkela_wire_6709)
    );

    bfr new_Jinkela_buffer_5189 (
        .din(new_Jinkela_wire_6666),
        .dout(new_Jinkela_wire_6667)
    );

    bfr new_Jinkela_buffer_5263 (
        .din(new_Jinkela_wire_6764),
        .dout(new_Jinkela_wire_6765)
    );

    bfr new_Jinkela_buffer_5190 (
        .din(new_Jinkela_wire_6667),
        .dout(new_Jinkela_wire_6668)
    );

    bfr new_Jinkela_buffer_5222 (
        .din(new_Jinkela_wire_6709),
        .dout(new_Jinkela_wire_6710)
    );

    bfr new_Jinkela_buffer_5191 (
        .din(new_Jinkela_wire_6668),
        .dout(new_Jinkela_wire_6669)
    );

    bfr new_Jinkela_buffer_5254 (
        .din(new_Jinkela_wire_6745),
        .dout(new_Jinkela_wire_6746)
    );

    bfr new_Jinkela_buffer_5192 (
        .din(new_Jinkela_wire_6669),
        .dout(new_Jinkela_wire_6670)
    );

    bfr new_Jinkela_buffer_5223 (
        .din(new_Jinkela_wire_6710),
        .dout(new_Jinkela_wire_6711)
    );

    bfr new_Jinkela_buffer_5193 (
        .din(new_Jinkela_wire_6670),
        .dout(new_Jinkela_wire_6671)
    );

    spl2 new_Jinkela_splitter_600 (
        .a(new_Jinkela_wire_6765),
        .b(new_Jinkela_wire_6766),
        .c(new_Jinkela_wire_6767)
    );

    bfr new_Jinkela_buffer_5194 (
        .din(new_Jinkela_wire_6671),
        .dout(new_Jinkela_wire_6672)
    );

    bfr new_Jinkela_buffer_5224 (
        .din(new_Jinkela_wire_6711),
        .dout(new_Jinkela_wire_6712)
    );

    bfr new_Jinkela_buffer_5195 (
        .din(new_Jinkela_wire_6672),
        .dout(new_Jinkela_wire_6673)
    );

    bfr new_Jinkela_buffer_5255 (
        .din(new_Jinkela_wire_6746),
        .dout(new_Jinkela_wire_6747)
    );

    spl2 new_Jinkela_splitter_588 (
        .a(new_Jinkela_wire_6673),
        .b(new_Jinkela_wire_6674),
        .c(new_Jinkela_wire_6675)
    );

    bfr new_Jinkela_buffer_5298 (
        .din(new_Jinkela_wire_6813),
        .dout(new_Jinkela_wire_6814)
    );

    bfr new_Jinkela_buffer_5225 (
        .din(new_Jinkela_wire_6712),
        .dout(new_Jinkela_wire_6713)
    );

    bfr new_Jinkela_buffer_5226 (
        .din(new_Jinkela_wire_6713),
        .dout(new_Jinkela_wire_6714)
    );

    bfr new_Jinkela_buffer_12052 (
        .din(new_Jinkela_wire_14525),
        .dout(new_Jinkela_wire_14526)
    );

    bfr new_Jinkela_buffer_12190 (
        .din(new_Jinkela_wire_14675),
        .dout(new_Jinkela_wire_14676)
    );

    bfr new_Jinkela_buffer_12130 (
        .din(new_Jinkela_wire_14607),
        .dout(new_Jinkela_wire_14608)
    );

    bfr new_Jinkela_buffer_12053 (
        .din(new_Jinkela_wire_14526),
        .dout(new_Jinkela_wire_14527)
    );

    bfr new_Jinkela_buffer_12054 (
        .din(new_Jinkela_wire_14527),
        .dout(new_Jinkela_wire_14528)
    );

    bfr new_Jinkela_buffer_12131 (
        .din(new_Jinkela_wire_14608),
        .dout(new_Jinkela_wire_14609)
    );

    bfr new_Jinkela_buffer_12055 (
        .din(new_Jinkela_wire_14528),
        .dout(new_Jinkela_wire_14529)
    );

    bfr new_Jinkela_buffer_12486 (
        .din(_1406_),
        .dout(new_Jinkela_wire_14990)
    );

    bfr new_Jinkela_buffer_12056 (
        .din(new_Jinkela_wire_14529),
        .dout(new_Jinkela_wire_14530)
    );

    bfr new_Jinkela_buffer_12191 (
        .din(new_Jinkela_wire_14676),
        .dout(new_Jinkela_wire_14677)
    );

    bfr new_Jinkela_buffer_12132 (
        .din(new_Jinkela_wire_14609),
        .dout(new_Jinkela_wire_14610)
    );

    bfr new_Jinkela_buffer_12057 (
        .din(new_Jinkela_wire_14530),
        .dout(new_Jinkela_wire_14531)
    );

    bfr new_Jinkela_buffer_12058 (
        .din(new_Jinkela_wire_14531),
        .dout(new_Jinkela_wire_14532)
    );

    bfr new_Jinkela_buffer_12200 (
        .din(new_Jinkela_wire_14697),
        .dout(new_Jinkela_wire_14698)
    );

    bfr new_Jinkela_buffer_12133 (
        .din(new_Jinkela_wire_14610),
        .dout(new_Jinkela_wire_14611)
    );

    bfr new_Jinkela_buffer_12059 (
        .din(new_Jinkela_wire_14532),
        .dout(new_Jinkela_wire_14533)
    );

    bfr new_Jinkela_buffer_12060 (
        .din(new_Jinkela_wire_14533),
        .dout(new_Jinkela_wire_14534)
    );

    bfr new_Jinkela_buffer_12192 (
        .din(new_Jinkela_wire_14677),
        .dout(new_Jinkela_wire_14678)
    );

    bfr new_Jinkela_buffer_12134 (
        .din(new_Jinkela_wire_14611),
        .dout(new_Jinkela_wire_14612)
    );

    bfr new_Jinkela_buffer_12061 (
        .din(new_Jinkela_wire_14534),
        .dout(new_Jinkela_wire_14535)
    );

    spl2 new_Jinkela_splitter_1086 (
        .a(new_Jinkela_wire_14535),
        .b(new_Jinkela_wire_14536),
        .c(new_Jinkela_wire_14537)
    );

    bfr new_Jinkela_buffer_12279 (
        .din(new_Jinkela_wire_14778),
        .dout(new_Jinkela_wire_14779)
    );

    bfr new_Jinkela_buffer_12135 (
        .din(new_Jinkela_wire_14612),
        .dout(new_Jinkela_wire_14613)
    );

    bfr new_Jinkela_buffer_12193 (
        .din(new_Jinkela_wire_14678),
        .dout(new_Jinkela_wire_14679)
    );

    bfr new_Jinkela_buffer_12136 (
        .din(new_Jinkela_wire_14613),
        .dout(new_Jinkela_wire_14614)
    );

    bfr new_Jinkela_buffer_12201 (
        .din(new_Jinkela_wire_14698),
        .dout(new_Jinkela_wire_14699)
    );

    bfr new_Jinkela_buffer_12137 (
        .din(new_Jinkela_wire_14614),
        .dout(new_Jinkela_wire_14615)
    );

    bfr new_Jinkela_buffer_12194 (
        .din(new_Jinkela_wire_14679),
        .dout(new_Jinkela_wire_14680)
    );

    bfr new_Jinkela_buffer_12138 (
        .din(new_Jinkela_wire_14615),
        .dout(new_Jinkela_wire_14616)
    );

    bfr new_Jinkela_buffer_12139 (
        .din(new_Jinkela_wire_14616),
        .dout(new_Jinkela_wire_14617)
    );

    bfr new_Jinkela_buffer_12487 (
        .din(_1470_),
        .dout(new_Jinkela_wire_14991)
    );

    spl2 new_Jinkela_splitter_1092 (
        .a(new_Jinkela_wire_14680),
        .b(new_Jinkela_wire_14681),
        .c(new_Jinkela_wire_14682)
    );

    bfr new_Jinkela_buffer_12140 (
        .din(new_Jinkela_wire_14617),
        .dout(new_Jinkela_wire_14618)
    );

    bfr new_Jinkela_buffer_12280 (
        .din(new_Jinkela_wire_14779),
        .dout(new_Jinkela_wire_14780)
    );

    bfr new_Jinkela_buffer_12141 (
        .din(new_Jinkela_wire_14618),
        .dout(new_Jinkela_wire_14619)
    );

    bfr new_Jinkela_buffer_12202 (
        .din(new_Jinkela_wire_14699),
        .dout(new_Jinkela_wire_14700)
    );

    bfr new_Jinkela_buffer_12142 (
        .din(new_Jinkela_wire_14619),
        .dout(new_Jinkela_wire_14620)
    );

    bfr new_Jinkela_buffer_12203 (
        .din(new_Jinkela_wire_14700),
        .dout(new_Jinkela_wire_14701)
    );

    bfr new_Jinkela_buffer_12143 (
        .din(new_Jinkela_wire_14620),
        .dout(new_Jinkela_wire_14621)
    );

    bfr new_Jinkela_buffer_12391 (
        .din(new_Jinkela_wire_14892),
        .dout(new_Jinkela_wire_14893)
    );

    bfr new_Jinkela_buffer_12144 (
        .din(new_Jinkela_wire_14621),
        .dout(new_Jinkela_wire_14622)
    );

    bfr new_Jinkela_buffer_12204 (
        .din(new_Jinkela_wire_14701),
        .dout(new_Jinkela_wire_14702)
    );

    bfr new_Jinkela_buffer_12145 (
        .din(new_Jinkela_wire_14622),
        .dout(new_Jinkela_wire_14623)
    );

    bfr new_Jinkela_buffer_15585 (
        .din(new_Jinkela_wire_18581),
        .dout(new_Jinkela_wire_18582)
    );

    bfr new_Jinkela_buffer_15567 (
        .din(new_Jinkela_wire_18557),
        .dout(new_Jinkela_wire_18558)
    );

    bfr new_Jinkela_buffer_15588 (
        .din(new_Jinkela_wire_18586),
        .dout(new_Jinkela_wire_18587)
    );

    bfr new_Jinkela_buffer_15568 (
        .din(new_Jinkela_wire_18558),
        .dout(new_Jinkela_wire_18559)
    );

    spl2 new_Jinkela_splitter_1347 (
        .a(new_Jinkela_wire_18582),
        .b(new_Jinkela_wire_18583),
        .c(new_Jinkela_wire_18584)
    );

    bfr new_Jinkela_buffer_15569 (
        .din(new_Jinkela_wire_18559),
        .dout(new_Jinkela_wire_18560)
    );

    bfr new_Jinkela_buffer_15589 (
        .din(new_Jinkela_wire_18587),
        .dout(new_Jinkela_wire_18588)
    );

    bfr new_Jinkela_buffer_15570 (
        .din(new_Jinkela_wire_18560),
        .dout(new_Jinkela_wire_18561)
    );

    spl2 new_Jinkela_splitter_1349 (
        .a(_1836_),
        .b(new_Jinkela_wire_18689),
        .c(new_Jinkela_wire_18690)
    );

    bfr new_Jinkela_buffer_15571 (
        .din(new_Jinkela_wire_18561),
        .dout(new_Jinkela_wire_18562)
    );

    bfr new_Jinkela_buffer_15687 (
        .din(_1517_),
        .dout(new_Jinkela_wire_18688)
    );

    spl2 new_Jinkela_splitter_1350 (
        .a(_0791_),
        .b(new_Jinkela_wire_18695),
        .c(new_Jinkela_wire_18696)
    );

    bfr new_Jinkela_buffer_15590 (
        .din(new_Jinkela_wire_18588),
        .dout(new_Jinkela_wire_18589)
    );

    bfr new_Jinkela_buffer_15688 (
        .din(new_Jinkela_wire_18690),
        .dout(new_Jinkela_wire_18691)
    );

    bfr new_Jinkela_buffer_15591 (
        .din(new_Jinkela_wire_18589),
        .dout(new_Jinkela_wire_18590)
    );

    bfr new_Jinkela_buffer_15592 (
        .din(new_Jinkela_wire_18590),
        .dout(new_Jinkela_wire_18591)
    );

    spl2 new_Jinkela_splitter_1351 (
        .a(_1431_),
        .b(new_Jinkela_wire_18697),
        .c(new_Jinkela_wire_18698)
    );

    bfr new_Jinkela_buffer_15593 (
        .din(new_Jinkela_wire_18591),
        .dout(new_Jinkela_wire_18592)
    );

    bfr new_Jinkela_buffer_15689 (
        .din(new_Jinkela_wire_18691),
        .dout(new_Jinkela_wire_18692)
    );

    bfr new_Jinkela_buffer_15594 (
        .din(new_Jinkela_wire_18592),
        .dout(new_Jinkela_wire_18593)
    );

    bfr new_Jinkela_buffer_15595 (
        .din(new_Jinkela_wire_18593),
        .dout(new_Jinkela_wire_18594)
    );

    bfr new_Jinkela_buffer_15692 (
        .din(_0369_),
        .dout(new_Jinkela_wire_18699)
    );

    bfr new_Jinkela_buffer_15690 (
        .din(new_Jinkela_wire_18692),
        .dout(new_Jinkela_wire_18693)
    );

    bfr new_Jinkela_buffer_15596 (
        .din(new_Jinkela_wire_18594),
        .dout(new_Jinkela_wire_18595)
    );

    spl2 new_Jinkela_splitter_1353 (
        .a(_0153_),
        .b(new_Jinkela_wire_18702),
        .c(new_Jinkela_wire_18703)
    );

    bfr new_Jinkela_buffer_15597 (
        .din(new_Jinkela_wire_18595),
        .dout(new_Jinkela_wire_18596)
    );

    spl2 new_Jinkela_splitter_1352 (
        .a(_1059_),
        .b(new_Jinkela_wire_18700),
        .c(new_Jinkela_wire_18701)
    );

    bfr new_Jinkela_buffer_15691 (
        .din(new_Jinkela_wire_18693),
        .dout(new_Jinkela_wire_18694)
    );

    bfr new_Jinkela_buffer_15598 (
        .din(new_Jinkela_wire_18596),
        .dout(new_Jinkela_wire_18597)
    );

    bfr new_Jinkela_buffer_15599 (
        .din(new_Jinkela_wire_18597),
        .dout(new_Jinkela_wire_18598)
    );

    bfr new_Jinkela_buffer_15600 (
        .din(new_Jinkela_wire_18598),
        .dout(new_Jinkela_wire_18599)
    );

    bfr new_Jinkela_buffer_15697 (
        .din(_1472_),
        .dout(new_Jinkela_wire_18708)
    );

    bfr new_Jinkela_buffer_15693 (
        .din(new_Jinkela_wire_18703),
        .dout(new_Jinkela_wire_18704)
    );

    bfr new_Jinkela_buffer_15601 (
        .din(new_Jinkela_wire_18599),
        .dout(new_Jinkela_wire_18600)
    );

    bfr new_Jinkela_buffer_15721 (
        .din(_1825_),
        .dout(new_Jinkela_wire_18734)
    );

    bfr new_Jinkela_buffer_15602 (
        .din(new_Jinkela_wire_18600),
        .dout(new_Jinkela_wire_18601)
    );

    bfr new_Jinkela_buffer_15745 (
        .din(_1837_),
        .dout(new_Jinkela_wire_18760)
    );

    bfr new_Jinkela_buffer_15694 (
        .din(new_Jinkela_wire_18704),
        .dout(new_Jinkela_wire_18705)
    );

    bfr new_Jinkela_buffer_15603 (
        .din(new_Jinkela_wire_18601),
        .dout(new_Jinkela_wire_18602)
    );

    bfr new_Jinkela_buffer_15698 (
        .din(new_Jinkela_wire_18708),
        .dout(new_Jinkela_wire_18709)
    );

    bfr new_Jinkela_buffer_15604 (
        .din(new_Jinkela_wire_18602),
        .dout(new_Jinkela_wire_18603)
    );

    bfr new_Jinkela_buffer_15695 (
        .din(new_Jinkela_wire_18705),
        .dout(new_Jinkela_wire_18706)
    );

    bfr new_Jinkela_buffer_15605 (
        .din(new_Jinkela_wire_18603),
        .dout(new_Jinkela_wire_18604)
    );

    and_bb _2749_ (
        .a(new_Jinkela_wire_369),
        .b(new_Jinkela_wire_118),
        .c(_1813_)
    );

    and_bi _2750_ (
        .a(new_Jinkela_wire_19155),
        .b(new_Jinkela_wire_21111),
        .c(_1814_)
    );

    and_bb _2751_ (
        .a(new_Jinkela_wire_689),
        .b(new_Jinkela_wire_8),
        .c(_1815_)
    );

    and_bi _2752_ (
        .a(new_Jinkela_wire_11835),
        .b(new_Jinkela_wire_12740),
        .c(_1816_)
    );

    and_bb _2753_ (
        .a(new_Jinkela_wire_461),
        .b(new_Jinkela_wire_504),
        .c(_1817_)
    );

    and_bi _2754_ (
        .a(new_Jinkela_wire_7511),
        .b(new_Jinkela_wire_1268),
        .c(_1818_)
    );

    and_bb _2755_ (
        .a(new_Jinkela_wire_253),
        .b(new_Jinkela_wire_32),
        .c(_1819_)
    );

    and_bi _2756_ (
        .a(new_Jinkela_wire_19281),
        .b(new_Jinkela_wire_21098),
        .c(_1820_)
    );

    and_bb _2757_ (
        .a(new_Jinkela_wire_192),
        .b(new_Jinkela_wire_306),
        .c(_1821_)
    );

    and_bi _2758_ (
        .a(new_Jinkela_wire_20354),
        .b(new_Jinkela_wire_11530),
        .c(_1822_)
    );

    and_bb _2759_ (
        .a(new_Jinkela_wire_385),
        .b(new_Jinkela_wire_54),
        .c(_1823_)
    );

    and_bi _2760_ (
        .a(new_Jinkela_wire_17061),
        .b(new_Jinkela_wire_16780),
        .c(_1824_)
    );

    and_bb _2761_ (
        .a(new_Jinkela_wire_411),
        .b(new_Jinkela_wire_655),
        .c(_1825_)
    );

    and_bi _2762_ (
        .a(new_Jinkela_wire_21104),
        .b(new_Jinkela_wire_19066),
        .c(_1826_)
    );

    and_bb _2763_ (
        .a(new_Jinkela_wire_167),
        .b(new_Jinkela_wire_629),
        .c(_1828_)
    );

    and_ii _2764_ (
        .a(new_Jinkela_wire_19115),
        .b(new_Jinkela_wire_15694),
        .c(_1829_)
    );

    or_ii _2765_ (
        .a(new_Jinkela_wire_431),
        .b(new_Jinkela_wire_320),
        .c(_1830_)
    );

    or_bb _2766_ (
        .a(new_Jinkela_wire_14259),
        .b(new_Jinkela_wire_18972),
        .c(_1831_)
    );

    and_bb _2767_ (
        .a(new_Jinkela_wire_611),
        .b(new_Jinkela_wire_533),
        .c(_1832_)
    );

    and_ii _2768_ (
        .a(new_Jinkela_wire_3241),
        .b(new_Jinkela_wire_4294),
        .c(_1833_)
    );

    and_bb _2769_ (
        .a(new_Jinkela_wire_3242),
        .b(new_Jinkela_wire_4295),
        .c(_1834_)
    );

    or_bb _2770_ (
        .a(new_Jinkela_wire_17553),
        .b(new_Jinkela_wire_10104),
        .c(_1835_)
    );

    or_bb _2771_ (
        .a(new_Jinkela_wire_20293),
        .b(new_Jinkela_wire_15119),
        .c(_1836_)
    );

    or_ii _2772_ (
        .a(new_Jinkela_wire_20294),
        .b(new_Jinkela_wire_15120),
        .c(_1837_)
    );

    or_ii _2773_ (
        .a(new_Jinkela_wire_18760),
        .b(new_Jinkela_wire_18689),
        .c(_0001_)
    );

    and_ii _2774_ (
        .a(new_Jinkela_wire_21177),
        .b(new_Jinkela_wire_18783),
        .c(_0002_)
    );

    and_bb _2775_ (
        .a(new_Jinkela_wire_21178),
        .b(new_Jinkela_wire_18784),
        .c(_0003_)
    );

    or_bb _2776_ (
        .a(new_Jinkela_wire_13969),
        .b(new_Jinkela_wire_4995),
        .c(_0004_)
    );

    or_bb _2777_ (
        .a(new_Jinkela_wire_20273),
        .b(new_Jinkela_wire_17862),
        .c(_0005_)
    );

    or_ii _2778_ (
        .a(new_Jinkela_wire_20274),
        .b(new_Jinkela_wire_17863),
        .c(_0006_)
    );

    or_ii _2779_ (
        .a(new_Jinkela_wire_17683),
        .b(new_Jinkela_wire_17016),
        .c(_0007_)
    );

    and_ii _2780_ (
        .a(new_Jinkela_wire_5991),
        .b(new_Jinkela_wire_18758),
        .c(_0008_)
    );

    and_bb _2781_ (
        .a(new_Jinkela_wire_5992),
        .b(new_Jinkela_wire_18759),
        .c(_0009_)
    );

    or_bb _2782_ (
        .a(new_Jinkela_wire_11403),
        .b(new_Jinkela_wire_17028),
        .c(_0010_)
    );

    or_bb _2783_ (
        .a(new_Jinkela_wire_6377),
        .b(new_Jinkela_wire_15773),
        .c(_0012_)
    );

    or_ii _2784_ (
        .a(new_Jinkela_wire_6378),
        .b(new_Jinkela_wire_15774),
        .c(_0013_)
    );

    or_ii _2785_ (
        .a(new_Jinkela_wire_12624),
        .b(new_Jinkela_wire_5457),
        .c(_0014_)
    );

    and_ii _2786_ (
        .a(new_Jinkela_wire_17660),
        .b(new_Jinkela_wire_16366),
        .c(_0015_)
    );

    and_bb _2787_ (
        .a(new_Jinkela_wire_17661),
        .b(new_Jinkela_wire_16367),
        .c(_0016_)
    );

    or_bb _2788_ (
        .a(new_Jinkela_wire_19334),
        .b(new_Jinkela_wire_11445),
        .c(_0017_)
    );

    or_bb _2789_ (
        .a(new_Jinkela_wire_12625),
        .b(new_Jinkela_wire_18834),
        .c(_0018_)
    );

    or_ii _2790_ (
        .a(new_Jinkela_wire_12626),
        .b(new_Jinkela_wire_18835),
        .c(_0019_)
    );

    bfr new_Jinkela_buffer_1615 (
        .din(new_Jinkela_wire_2510),
        .dout(new_Jinkela_wire_2511)
    );

    bfr new_Jinkela_buffer_1705 (
        .din(new_Jinkela_wire_2610),
        .dout(new_Jinkela_wire_2611)
    );

    bfr new_Jinkela_buffer_1616 (
        .din(new_Jinkela_wire_2511),
        .dout(new_Jinkela_wire_2512)
    );

    spl2 new_Jinkela_splitter_309 (
        .a(_1210_),
        .b(new_Jinkela_wire_2789),
        .c(new_Jinkela_wire_2790)
    );

    bfr new_Jinkela_buffer_1617 (
        .din(new_Jinkela_wire_2512),
        .dout(new_Jinkela_wire_2513)
    );

    bfr new_Jinkela_buffer_1706 (
        .din(new_Jinkela_wire_2611),
        .dout(new_Jinkela_wire_2612)
    );

    bfr new_Jinkela_buffer_1618 (
        .din(new_Jinkela_wire_2513),
        .dout(new_Jinkela_wire_2514)
    );

    spl2 new_Jinkela_splitter_304 (
        .a(new_Jinkela_wire_2658),
        .b(new_Jinkela_wire_2659),
        .c(new_Jinkela_wire_2660)
    );

    bfr new_Jinkela_buffer_1619 (
        .din(new_Jinkela_wire_2514),
        .dout(new_Jinkela_wire_2515)
    );

    bfr new_Jinkela_buffer_1707 (
        .din(new_Jinkela_wire_2612),
        .dout(new_Jinkela_wire_2613)
    );

    bfr new_Jinkela_buffer_1620 (
        .din(new_Jinkela_wire_2515),
        .dout(new_Jinkela_wire_2516)
    );

    spl2 new_Jinkela_splitter_308 (
        .a(_0388_),
        .b(new_Jinkela_wire_2787),
        .c(new_Jinkela_wire_2788)
    );

    bfr new_Jinkela_buffer_1621 (
        .din(new_Jinkela_wire_2516),
        .dout(new_Jinkela_wire_2517)
    );

    bfr new_Jinkela_buffer_1708 (
        .din(new_Jinkela_wire_2613),
        .dout(new_Jinkela_wire_2614)
    );

    bfr new_Jinkela_buffer_1622 (
        .din(new_Jinkela_wire_2517),
        .dout(new_Jinkela_wire_2518)
    );

    bfr new_Jinkela_buffer_1751 (
        .din(new_Jinkela_wire_2662),
        .dout(new_Jinkela_wire_2663)
    );

    bfr new_Jinkela_buffer_1623 (
        .din(new_Jinkela_wire_2518),
        .dout(new_Jinkela_wire_2519)
    );

    bfr new_Jinkela_buffer_1709 (
        .din(new_Jinkela_wire_2614),
        .dout(new_Jinkela_wire_2615)
    );

    bfr new_Jinkela_buffer_1624 (
        .din(new_Jinkela_wire_2519),
        .dout(new_Jinkela_wire_2520)
    );

    bfr new_Jinkela_buffer_1752 (
        .din(new_Jinkela_wire_2663),
        .dout(new_Jinkela_wire_2664)
    );

    bfr new_Jinkela_buffer_1625 (
        .din(new_Jinkela_wire_2520),
        .dout(new_Jinkela_wire_2521)
    );

    bfr new_Jinkela_buffer_1710 (
        .din(new_Jinkela_wire_2615),
        .dout(new_Jinkela_wire_2616)
    );

    bfr new_Jinkela_buffer_1626 (
        .din(new_Jinkela_wire_2521),
        .dout(new_Jinkela_wire_2522)
    );

    bfr new_Jinkela_buffer_1798 (
        .din(new_Jinkela_wire_2713),
        .dout(new_Jinkela_wire_2714)
    );

    bfr new_Jinkela_buffer_1627 (
        .din(new_Jinkela_wire_2522),
        .dout(new_Jinkela_wire_2523)
    );

    bfr new_Jinkela_buffer_1711 (
        .din(new_Jinkela_wire_2616),
        .dout(new_Jinkela_wire_2617)
    );

    bfr new_Jinkela_buffer_1628 (
        .din(new_Jinkela_wire_2523),
        .dout(new_Jinkela_wire_2524)
    );

    bfr new_Jinkela_buffer_1753 (
        .din(new_Jinkela_wire_2664),
        .dout(new_Jinkela_wire_2665)
    );

    bfr new_Jinkela_buffer_1629 (
        .din(new_Jinkela_wire_2524),
        .dout(new_Jinkela_wire_2525)
    );

    bfr new_Jinkela_buffer_1712 (
        .din(new_Jinkela_wire_2617),
        .dout(new_Jinkela_wire_2618)
    );

    bfr new_Jinkela_buffer_1630 (
        .din(new_Jinkela_wire_2525),
        .dout(new_Jinkela_wire_2526)
    );

    bfr new_Jinkela_buffer_1869 (
        .din(new_net_3918),
        .dout(new_Jinkela_wire_2791)
    );

    bfr new_Jinkela_buffer_1631 (
        .din(new_Jinkela_wire_2526),
        .dout(new_Jinkela_wire_2527)
    );

    bfr new_Jinkela_buffer_1713 (
        .din(new_Jinkela_wire_2618),
        .dout(new_Jinkela_wire_2619)
    );

    bfr new_Jinkela_buffer_1632 (
        .din(new_Jinkela_wire_2527),
        .dout(new_Jinkela_wire_2528)
    );

    bfr new_Jinkela_buffer_1754 (
        .din(new_Jinkela_wire_2665),
        .dout(new_Jinkela_wire_2666)
    );

    bfr new_Jinkela_buffer_1633 (
        .din(new_Jinkela_wire_2528),
        .dout(new_Jinkela_wire_2529)
    );

    bfr new_Jinkela_buffer_1714 (
        .din(new_Jinkela_wire_2619),
        .dout(new_Jinkela_wire_2620)
    );

    bfr new_Jinkela_buffer_1634 (
        .din(new_Jinkela_wire_2529),
        .dout(new_Jinkela_wire_2530)
    );

    bfr new_Jinkela_buffer_1799 (
        .din(new_Jinkela_wire_2714),
        .dout(new_Jinkela_wire_2715)
    );

    bfr new_Jinkela_buffer_1635 (
        .din(new_Jinkela_wire_2530),
        .dout(new_Jinkela_wire_2531)
    );

    bfr new_Jinkela_buffer_1715 (
        .din(new_Jinkela_wire_2620),
        .dout(new_Jinkela_wire_2621)
    );

    bfr new_Jinkela_buffer_15606 (
        .din(new_Jinkela_wire_18604),
        .dout(new_Jinkela_wire_18605)
    );

    spl2 new_Jinkela_splitter_1356 (
        .a(_1151_),
        .b(new_Jinkela_wire_18761),
        .c(new_Jinkela_wire_18762)
    );

    bfr new_Jinkela_buffer_15696 (
        .din(new_Jinkela_wire_18706),
        .dout(new_Jinkela_wire_18707)
    );

    bfr new_Jinkela_buffer_15607 (
        .din(new_Jinkela_wire_18605),
        .dout(new_Jinkela_wire_18606)
    );

    bfr new_Jinkela_buffer_15699 (
        .din(new_Jinkela_wire_18709),
        .dout(new_Jinkela_wire_18710)
    );

    bfr new_Jinkela_buffer_15608 (
        .din(new_Jinkela_wire_18606),
        .dout(new_Jinkela_wire_18607)
    );

    bfr new_Jinkela_buffer_15722 (
        .din(new_Jinkela_wire_18734),
        .dout(new_Jinkela_wire_18735)
    );

    bfr new_Jinkela_buffer_15609 (
        .din(new_Jinkela_wire_18607),
        .dout(new_Jinkela_wire_18608)
    );

    bfr new_Jinkela_buffer_15700 (
        .din(new_Jinkela_wire_18710),
        .dout(new_Jinkela_wire_18711)
    );

    bfr new_Jinkela_buffer_15610 (
        .din(new_Jinkela_wire_18608),
        .dout(new_Jinkela_wire_18609)
    );

    spl2 new_Jinkela_splitter_1357 (
        .a(_1483_),
        .b(new_Jinkela_wire_18763),
        .c(new_Jinkela_wire_18764)
    );

    bfr new_Jinkela_buffer_15611 (
        .din(new_Jinkela_wire_18609),
        .dout(new_Jinkela_wire_18610)
    );

    bfr new_Jinkela_buffer_15701 (
        .din(new_Jinkela_wire_18711),
        .dout(new_Jinkela_wire_18712)
    );

    bfr new_Jinkela_buffer_15612 (
        .din(new_Jinkela_wire_18610),
        .dout(new_Jinkela_wire_18611)
    );

    bfr new_Jinkela_buffer_15723 (
        .din(new_Jinkela_wire_18735),
        .dout(new_Jinkela_wire_18736)
    );

    bfr new_Jinkela_buffer_15613 (
        .din(new_Jinkela_wire_18611),
        .dout(new_Jinkela_wire_18612)
    );

    bfr new_Jinkela_buffer_15702 (
        .din(new_Jinkela_wire_18712),
        .dout(new_Jinkela_wire_18713)
    );

    bfr new_Jinkela_buffer_15614 (
        .din(new_Jinkela_wire_18612),
        .dout(new_Jinkela_wire_18613)
    );

    bfr new_Jinkela_buffer_15615 (
        .din(new_Jinkela_wire_18613),
        .dout(new_Jinkela_wire_18614)
    );

    bfr new_Jinkela_buffer_15703 (
        .din(new_Jinkela_wire_18713),
        .dout(new_Jinkela_wire_18714)
    );

    bfr new_Jinkela_buffer_15616 (
        .din(new_Jinkela_wire_18614),
        .dout(new_Jinkela_wire_18615)
    );

    bfr new_Jinkela_buffer_15724 (
        .din(new_Jinkela_wire_18736),
        .dout(new_Jinkela_wire_18737)
    );

    bfr new_Jinkela_buffer_15617 (
        .din(new_Jinkela_wire_18615),
        .dout(new_Jinkela_wire_18616)
    );

    bfr new_Jinkela_buffer_15704 (
        .din(new_Jinkela_wire_18714),
        .dout(new_Jinkela_wire_18715)
    );

    bfr new_Jinkela_buffer_15618 (
        .din(new_Jinkela_wire_18616),
        .dout(new_Jinkela_wire_18617)
    );

    bfr new_Jinkela_buffer_15619 (
        .din(new_Jinkela_wire_18617),
        .dout(new_Jinkela_wire_18618)
    );

    bfr new_Jinkela_buffer_15750 (
        .din(_1828_),
        .dout(new_Jinkela_wire_18769)
    );

    bfr new_Jinkela_buffer_15705 (
        .din(new_Jinkela_wire_18715),
        .dout(new_Jinkela_wire_18716)
    );

    bfr new_Jinkela_buffer_15620 (
        .din(new_Jinkela_wire_18618),
        .dout(new_Jinkela_wire_18619)
    );

    bfr new_Jinkela_buffer_15725 (
        .din(new_Jinkela_wire_18737),
        .dout(new_Jinkela_wire_18738)
    );

    bfr new_Jinkela_buffer_15621 (
        .din(new_Jinkela_wire_18619),
        .dout(new_Jinkela_wire_18620)
    );

    bfr new_Jinkela_buffer_15706 (
        .din(new_Jinkela_wire_18716),
        .dout(new_Jinkela_wire_18717)
    );

    bfr new_Jinkela_buffer_15622 (
        .din(new_Jinkela_wire_18620),
        .dout(new_Jinkela_wire_18621)
    );

    bfr new_Jinkela_buffer_15746 (
        .din(new_Jinkela_wire_18764),
        .dout(new_Jinkela_wire_18765)
    );

    bfr new_Jinkela_buffer_15623 (
        .din(new_Jinkela_wire_18621),
        .dout(new_Jinkela_wire_18622)
    );

    spl2 new_Jinkela_splitter_1359 (
        .a(_1106_),
        .b(new_Jinkela_wire_18785),
        .c(new_Jinkela_wire_18786)
    );

    bfr new_Jinkela_buffer_15707 (
        .din(new_Jinkela_wire_18717),
        .dout(new_Jinkela_wire_18718)
    );

    bfr new_Jinkela_buffer_15624 (
        .din(new_Jinkela_wire_18622),
        .dout(new_Jinkela_wire_18623)
    );

    bfr new_Jinkela_buffer_15726 (
        .din(new_Jinkela_wire_18738),
        .dout(new_Jinkela_wire_18739)
    );

    bfr new_Jinkela_buffer_15625 (
        .din(new_Jinkela_wire_18623),
        .dout(new_Jinkela_wire_18624)
    );

    bfr new_Jinkela_buffer_15708 (
        .din(new_Jinkela_wire_18718),
        .dout(new_Jinkela_wire_18719)
    );

    bfr new_Jinkela_buffer_15626 (
        .din(new_Jinkela_wire_18624),
        .dout(new_Jinkela_wire_18625)
    );

    bfr new_Jinkela_buffer_5256 (
        .din(new_Jinkela_wire_6747),
        .dout(new_Jinkela_wire_6748)
    );

    bfr new_Jinkela_buffer_8763 (
        .din(new_Jinkela_wire_10748),
        .dout(new_Jinkela_wire_10749)
    );

    bfr new_Jinkela_buffer_5227 (
        .din(new_Jinkela_wire_6714),
        .dout(new_Jinkela_wire_6715)
    );

    bfr new_Jinkela_buffer_8677 (
        .din(new_Jinkela_wire_10644),
        .dout(new_Jinkela_wire_10645)
    );

    bfr new_Jinkela_buffer_8720 (
        .din(new_Jinkela_wire_10701),
        .dout(new_Jinkela_wire_10702)
    );

    spl2 new_Jinkela_splitter_603 (
        .a(_0387_),
        .b(new_Jinkela_wire_6804),
        .c(new_Jinkela_wire_6805)
    );

    bfr new_Jinkela_buffer_5228 (
        .din(new_Jinkela_wire_6715),
        .dout(new_Jinkela_wire_6716)
    );

    bfr new_Jinkela_buffer_8678 (
        .din(new_Jinkela_wire_10645),
        .dout(new_Jinkela_wire_10646)
    );

    bfr new_Jinkela_buffer_5257 (
        .din(new_Jinkela_wire_6748),
        .dout(new_Jinkela_wire_6749)
    );

    bfr new_Jinkela_buffer_8766 (
        .din(new_Jinkela_wire_10753),
        .dout(new_Jinkela_wire_10754)
    );

    bfr new_Jinkela_buffer_5229 (
        .din(new_Jinkela_wire_6716),
        .dout(new_Jinkela_wire_6717)
    );

    bfr new_Jinkela_buffer_8679 (
        .din(new_Jinkela_wire_10646),
        .dout(new_Jinkela_wire_10647)
    );

    bfr new_Jinkela_buffer_8721 (
        .din(new_Jinkela_wire_10702),
        .dout(new_Jinkela_wire_10703)
    );

    spl2 new_Jinkela_splitter_604 (
        .a(_0857_),
        .b(new_Jinkela_wire_6806),
        .c(new_Jinkela_wire_6807)
    );

    bfr new_Jinkela_buffer_5230 (
        .din(new_Jinkela_wire_6717),
        .dout(new_Jinkela_wire_6718)
    );

    bfr new_Jinkela_buffer_8680 (
        .din(new_Jinkela_wire_10647),
        .dout(new_Jinkela_wire_10648)
    );

    bfr new_Jinkela_buffer_5258 (
        .din(new_Jinkela_wire_6749),
        .dout(new_Jinkela_wire_6750)
    );

    bfr new_Jinkela_buffer_8764 (
        .din(new_Jinkela_wire_10749),
        .dout(new_Jinkela_wire_10750)
    );

    bfr new_Jinkela_buffer_5231 (
        .din(new_Jinkela_wire_6718),
        .dout(new_Jinkela_wire_6719)
    );

    bfr new_Jinkela_buffer_8681 (
        .din(new_Jinkela_wire_10648),
        .dout(new_Jinkela_wire_10649)
    );

    bfr new_Jinkela_buffer_5265 (
        .din(new_Jinkela_wire_6770),
        .dout(new_Jinkela_wire_6771)
    );

    bfr new_Jinkela_buffer_8722 (
        .din(new_Jinkela_wire_10703),
        .dout(new_Jinkela_wire_10704)
    );

    bfr new_Jinkela_buffer_5232 (
        .din(new_Jinkela_wire_6719),
        .dout(new_Jinkela_wire_6720)
    );

    bfr new_Jinkela_buffer_8682 (
        .din(new_Jinkela_wire_10649),
        .dout(new_Jinkela_wire_10650)
    );

    bfr new_Jinkela_buffer_5259 (
        .din(new_Jinkela_wire_6750),
        .dout(new_Jinkela_wire_6751)
    );

    spl2 new_Jinkela_splitter_847 (
        .a(_1613_),
        .b(new_Jinkela_wire_10957),
        .c(new_Jinkela_wire_10958)
    );

    bfr new_Jinkela_buffer_5233 (
        .din(new_Jinkela_wire_6720),
        .dout(new_Jinkela_wire_6721)
    );

    bfr new_Jinkela_buffer_8683 (
        .din(new_Jinkela_wire_10650),
        .dout(new_Jinkela_wire_10651)
    );

    bfr new_Jinkela_buffer_8723 (
        .din(new_Jinkela_wire_10704),
        .dout(new_Jinkela_wire_10705)
    );

    bfr new_Jinkela_buffer_5234 (
        .din(new_Jinkela_wire_6721),
        .dout(new_Jinkela_wire_6722)
    );

    bfr new_Jinkela_buffer_8684 (
        .din(new_Jinkela_wire_10651),
        .dout(new_Jinkela_wire_10652)
    );

    bfr new_Jinkela_buffer_5260 (
        .din(new_Jinkela_wire_6751),
        .dout(new_Jinkela_wire_6752)
    );

    bfr new_Jinkela_buffer_8767 (
        .din(new_Jinkela_wire_10754),
        .dout(new_Jinkela_wire_10755)
    );

    bfr new_Jinkela_buffer_5235 (
        .din(new_Jinkela_wire_6722),
        .dout(new_Jinkela_wire_6723)
    );

    bfr new_Jinkela_buffer_8685 (
        .din(new_Jinkela_wire_10652),
        .dout(new_Jinkela_wire_10653)
    );

    bfr new_Jinkela_buffer_5266 (
        .din(new_Jinkela_wire_6771),
        .dout(new_Jinkela_wire_6772)
    );

    bfr new_Jinkela_buffer_8724 (
        .din(new_Jinkela_wire_10705),
        .dout(new_Jinkela_wire_10706)
    );

    bfr new_Jinkela_buffer_5236 (
        .din(new_Jinkela_wire_6723),
        .dout(new_Jinkela_wire_6724)
    );

    bfr new_Jinkela_buffer_8686 (
        .din(new_Jinkela_wire_10653),
        .dout(new_Jinkela_wire_10654)
    );

    bfr new_Jinkela_buffer_5261 (
        .din(new_Jinkela_wire_6752),
        .dout(new_Jinkela_wire_6753)
    );

    spl2 new_Jinkela_splitter_846 (
        .a(_1184_),
        .b(new_Jinkela_wire_10951),
        .c(new_Jinkela_wire_10952)
    );

    bfr new_Jinkela_buffer_5237 (
        .din(new_Jinkela_wire_6724),
        .dout(new_Jinkela_wire_6725)
    );

    bfr new_Jinkela_buffer_8687 (
        .din(new_Jinkela_wire_10654),
        .dout(new_Jinkela_wire_10655)
    );

    bfr new_Jinkela_buffer_8725 (
        .din(new_Jinkela_wire_10706),
        .dout(new_Jinkela_wire_10707)
    );

    spl2 new_Jinkela_splitter_605 (
        .a(_0302_),
        .b(new_Jinkela_wire_6808),
        .c(new_Jinkela_wire_6809)
    );

    bfr new_Jinkela_buffer_5238 (
        .din(new_Jinkela_wire_6725),
        .dout(new_Jinkela_wire_6726)
    );

    bfr new_Jinkela_buffer_8688 (
        .din(new_Jinkela_wire_10655),
        .dout(new_Jinkela_wire_10656)
    );

    bfr new_Jinkela_buffer_5262 (
        .din(new_Jinkela_wire_6753),
        .dout(new_Jinkela_wire_6754)
    );

    bfr new_Jinkela_buffer_8768 (
        .din(new_Jinkela_wire_10755),
        .dout(new_Jinkela_wire_10756)
    );

    bfr new_Jinkela_buffer_5239 (
        .din(new_Jinkela_wire_6726),
        .dout(new_Jinkela_wire_6727)
    );

    bfr new_Jinkela_buffer_8689 (
        .din(new_Jinkela_wire_10656),
        .dout(new_Jinkela_wire_10657)
    );

    bfr new_Jinkela_buffer_5267 (
        .din(new_Jinkela_wire_6772),
        .dout(new_Jinkela_wire_6773)
    );

    bfr new_Jinkela_buffer_8726 (
        .din(new_Jinkela_wire_10707),
        .dout(new_Jinkela_wire_10708)
    );

    bfr new_Jinkela_buffer_5240 (
        .din(new_Jinkela_wire_6727),
        .dout(new_Jinkela_wire_6728)
    );

    bfr new_Jinkela_buffer_8690 (
        .din(new_Jinkela_wire_10657),
        .dout(new_Jinkela_wire_10658)
    );

    spl2 new_Jinkela_splitter_595 (
        .a(new_Jinkela_wire_6754),
        .b(new_Jinkela_wire_6755),
        .c(new_Jinkela_wire_6756)
    );

    bfr new_Jinkela_buffer_8846 (
        .din(new_Jinkela_wire_10837),
        .dout(new_Jinkela_wire_10838)
    );

    bfr new_Jinkela_buffer_5241 (
        .din(new_Jinkela_wire_6728),
        .dout(new_Jinkela_wire_6729)
    );

    bfr new_Jinkela_buffer_8691 (
        .din(new_Jinkela_wire_10658),
        .dout(new_Jinkela_wire_10659)
    );

    bfr new_Jinkela_buffer_5268 (
        .din(new_Jinkela_wire_6773),
        .dout(new_Jinkela_wire_6774)
    );

    bfr new_Jinkela_buffer_8727 (
        .din(new_Jinkela_wire_10708),
        .dout(new_Jinkela_wire_10709)
    );

    bfr new_Jinkela_buffer_5242 (
        .din(new_Jinkela_wire_6729),
        .dout(new_Jinkela_wire_6730)
    );

    bfr new_Jinkela_buffer_8692 (
        .din(new_Jinkela_wire_10659),
        .dout(new_Jinkela_wire_10660)
    );

    bfr new_Jinkela_buffer_8769 (
        .din(new_Jinkela_wire_10756),
        .dout(new_Jinkela_wire_10757)
    );

    spl2 new_Jinkela_splitter_606 (
        .a(_0087_),
        .b(new_Jinkela_wire_6810),
        .c(new_Jinkela_wire_6811)
    );

    bfr new_Jinkela_buffer_5243 (
        .din(new_Jinkela_wire_6730),
        .dout(new_Jinkela_wire_6731)
    );

    bfr new_Jinkela_buffer_8693 (
        .din(new_Jinkela_wire_10660),
        .dout(new_Jinkela_wire_10661)
    );

    bfr new_Jinkela_buffer_8728 (
        .din(new_Jinkela_wire_10709),
        .dout(new_Jinkela_wire_10710)
    );

    bfr new_Jinkela_buffer_5296 (
        .din(_0612_),
        .dout(new_Jinkela_wire_6812)
    );

    spl2 new_Jinkela_splitter_593 (
        .a(new_Jinkela_wire_6731),
        .b(new_Jinkela_wire_6732),
        .c(new_Jinkela_wire_6733)
    );

    bfr new_Jinkela_buffer_8694 (
        .din(new_Jinkela_wire_10661),
        .dout(new_Jinkela_wire_10662)
    );

    spl2 new_Jinkela_splitter_608 (
        .a(_1760_),
        .b(new_Jinkela_wire_6846),
        .c(new_Jinkela_wire_6847)
    );

    bfr new_Jinkela_buffer_8957 (
        .din(new_Jinkela_wire_10952),
        .dout(new_Jinkela_wire_10953)
    );

    bfr new_Jinkela_buffer_5269 (
        .din(new_Jinkela_wire_6774),
        .dout(new_Jinkela_wire_6775)
    );

    bfr new_Jinkela_buffer_8695 (
        .din(new_Jinkela_wire_10662),
        .dout(new_Jinkela_wire_10663)
    );

    bfr new_Jinkela_buffer_5270 (
        .din(new_Jinkela_wire_6775),
        .dout(new_Jinkela_wire_6776)
    );

    bfr new_Jinkela_buffer_8729 (
        .din(new_Jinkela_wire_10710),
        .dout(new_Jinkela_wire_10711)
    );

    bfr new_Jinkela_buffer_5297 (
        .din(new_Jinkela_wire_6812),
        .dout(new_Jinkela_wire_6813)
    );

    bfr new_Jinkela_buffer_8696 (
        .din(new_Jinkela_wire_10663),
        .dout(new_Jinkela_wire_10664)
    );

    bfr new_Jinkela_buffer_5271 (
        .din(new_Jinkela_wire_6776),
        .dout(new_Jinkela_wire_6777)
    );

    bfr new_Jinkela_buffer_8770 (
        .din(new_Jinkela_wire_10757),
        .dout(new_Jinkela_wire_10758)
    );

    bfr new_Jinkela_buffer_5332 (
        .din(_1753_),
        .dout(new_Jinkela_wire_6854)
    );

    bfr new_Jinkela_buffer_8697 (
        .din(new_Jinkela_wire_10664),
        .dout(new_Jinkela_wire_10665)
    );

    bfr new_Jinkela_buffer_5264 (
        .din(_1213_),
        .dout(new_Jinkela_wire_6770)
    );

    bfr new_Jinkela_buffer_8730 (
        .din(new_Jinkela_wire_10711),
        .dout(new_Jinkela_wire_10712)
    );

    bfr new_Jinkela_buffer_1636 (
        .din(new_Jinkela_wire_2531),
        .dout(new_Jinkela_wire_2532)
    );

    bfr new_Jinkela_buffer_8698 (
        .din(new_Jinkela_wire_10665),
        .dout(new_Jinkela_wire_10666)
    );

    bfr new_Jinkela_buffer_12281 (
        .din(new_Jinkela_wire_14780),
        .dout(new_Jinkela_wire_14781)
    );

    bfr new_Jinkela_buffer_1755 (
        .din(new_Jinkela_wire_2666),
        .dout(new_Jinkela_wire_2667)
    );

    bfr new_Jinkela_buffer_12146 (
        .din(new_Jinkela_wire_14623),
        .dout(new_Jinkela_wire_14624)
    );

    bfr new_Jinkela_buffer_8847 (
        .din(new_Jinkela_wire_10838),
        .dout(new_Jinkela_wire_10839)
    );

    bfr new_Jinkela_buffer_1637 (
        .din(new_Jinkela_wire_2532),
        .dout(new_Jinkela_wire_2533)
    );

    bfr new_Jinkela_buffer_8699 (
        .din(new_Jinkela_wire_10666),
        .dout(new_Jinkela_wire_10667)
    );

    bfr new_Jinkela_buffer_12205 (
        .din(new_Jinkela_wire_14702),
        .dout(new_Jinkela_wire_14703)
    );

    bfr new_Jinkela_buffer_1716 (
        .din(new_Jinkela_wire_2621),
        .dout(new_Jinkela_wire_2622)
    );

    bfr new_Jinkela_buffer_12147 (
        .din(new_Jinkela_wire_14624),
        .dout(new_Jinkela_wire_14625)
    );

    bfr new_Jinkela_buffer_8731 (
        .din(new_Jinkela_wire_10712),
        .dout(new_Jinkela_wire_10713)
    );

    bfr new_Jinkela_buffer_1638 (
        .din(new_Jinkela_wire_2533),
        .dout(new_Jinkela_wire_2534)
    );

    bfr new_Jinkela_buffer_8700 (
        .din(new_Jinkela_wire_10667),
        .dout(new_Jinkela_wire_10668)
    );

    bfr new_Jinkela_buffer_12519 (
        .din(_0577_),
        .dout(new_Jinkela_wire_15025)
    );

    bfr new_Jinkela_buffer_12148 (
        .din(new_Jinkela_wire_14625),
        .dout(new_Jinkela_wire_14626)
    );

    bfr new_Jinkela_buffer_1870 (
        .din(new_Jinkela_wire_2791),
        .dout(new_Jinkela_wire_2792)
    );

    bfr new_Jinkela_buffer_8771 (
        .din(new_Jinkela_wire_10758),
        .dout(new_Jinkela_wire_10759)
    );

    bfr new_Jinkela_buffer_1639 (
        .din(new_Jinkela_wire_2534),
        .dout(new_Jinkela_wire_2535)
    );

    bfr new_Jinkela_buffer_8701 (
        .din(new_Jinkela_wire_10668),
        .dout(new_Jinkela_wire_10669)
    );

    bfr new_Jinkela_buffer_12206 (
        .din(new_Jinkela_wire_14703),
        .dout(new_Jinkela_wire_14704)
    );

    bfr new_Jinkela_buffer_1717 (
        .din(new_Jinkela_wire_2622),
        .dout(new_Jinkela_wire_2623)
    );

    bfr new_Jinkela_buffer_12149 (
        .din(new_Jinkela_wire_14626),
        .dout(new_Jinkela_wire_14627)
    );

    bfr new_Jinkela_buffer_8732 (
        .din(new_Jinkela_wire_10713),
        .dout(new_Jinkela_wire_10714)
    );

    bfr new_Jinkela_buffer_1640 (
        .din(new_Jinkela_wire_2535),
        .dout(new_Jinkela_wire_2536)
    );

    bfr new_Jinkela_buffer_8702 (
        .din(new_Jinkela_wire_10669),
        .dout(new_Jinkela_wire_10670)
    );

    bfr new_Jinkela_buffer_12282 (
        .din(new_Jinkela_wire_14781),
        .dout(new_Jinkela_wire_14782)
    );

    bfr new_Jinkela_buffer_1756 (
        .din(new_Jinkela_wire_2667),
        .dout(new_Jinkela_wire_2668)
    );

    bfr new_Jinkela_buffer_12150 (
        .din(new_Jinkela_wire_14627),
        .dout(new_Jinkela_wire_14628)
    );

    bfr new_Jinkela_buffer_1641 (
        .din(new_Jinkela_wire_2536),
        .dout(new_Jinkela_wire_2537)
    );

    bfr new_Jinkela_buffer_8703 (
        .din(new_Jinkela_wire_10670),
        .dout(new_Jinkela_wire_10671)
    );

    bfr new_Jinkela_buffer_12207 (
        .din(new_Jinkela_wire_14704),
        .dout(new_Jinkela_wire_14705)
    );

    bfr new_Jinkela_buffer_1718 (
        .din(new_Jinkela_wire_2623),
        .dout(new_Jinkela_wire_2624)
    );

    bfr new_Jinkela_buffer_12151 (
        .din(new_Jinkela_wire_14628),
        .dout(new_Jinkela_wire_14629)
    );

    bfr new_Jinkela_buffer_8733 (
        .din(new_Jinkela_wire_10714),
        .dout(new_Jinkela_wire_10715)
    );

    bfr new_Jinkela_buffer_1642 (
        .din(new_Jinkela_wire_2537),
        .dout(new_Jinkela_wire_2538)
    );

    spl2 new_Jinkela_splitter_833 (
        .a(new_Jinkela_wire_10671),
        .b(new_Jinkela_wire_10672),
        .c(new_Jinkela_wire_10673)
    );

    bfr new_Jinkela_buffer_12392 (
        .din(new_Jinkela_wire_14893),
        .dout(new_Jinkela_wire_14894)
    );

    bfr new_Jinkela_buffer_1800 (
        .din(new_Jinkela_wire_2715),
        .dout(new_Jinkela_wire_2716)
    );

    bfr new_Jinkela_buffer_12152 (
        .din(new_Jinkela_wire_14629),
        .dout(new_Jinkela_wire_14630)
    );

    bfr new_Jinkela_buffer_8734 (
        .din(new_Jinkela_wire_10715),
        .dout(new_Jinkela_wire_10716)
    );

    bfr new_Jinkela_buffer_1643 (
        .din(new_Jinkela_wire_2538),
        .dout(new_Jinkela_wire_2539)
    );

    bfr new_Jinkela_buffer_8772 (
        .din(new_Jinkela_wire_10759),
        .dout(new_Jinkela_wire_10760)
    );

    bfr new_Jinkela_buffer_12208 (
        .din(new_Jinkela_wire_14705),
        .dout(new_Jinkela_wire_14706)
    );

    bfr new_Jinkela_buffer_1719 (
        .din(new_Jinkela_wire_2624),
        .dout(new_Jinkela_wire_2625)
    );

    bfr new_Jinkela_buffer_12153 (
        .din(new_Jinkela_wire_14630),
        .dout(new_Jinkela_wire_14631)
    );

    bfr new_Jinkela_buffer_8848 (
        .din(new_Jinkela_wire_10839),
        .dout(new_Jinkela_wire_10840)
    );

    bfr new_Jinkela_buffer_1644 (
        .din(new_Jinkela_wire_2539),
        .dout(new_Jinkela_wire_2540)
    );

    bfr new_Jinkela_buffer_8735 (
        .din(new_Jinkela_wire_10716),
        .dout(new_Jinkela_wire_10717)
    );

    bfr new_Jinkela_buffer_12283 (
        .din(new_Jinkela_wire_14782),
        .dout(new_Jinkela_wire_14783)
    );

    bfr new_Jinkela_buffer_1757 (
        .din(new_Jinkela_wire_2668),
        .dout(new_Jinkela_wire_2669)
    );

    bfr new_Jinkela_buffer_12154 (
        .din(new_Jinkela_wire_14631),
        .dout(new_Jinkela_wire_14632)
    );

    bfr new_Jinkela_buffer_8773 (
        .din(new_Jinkela_wire_10760),
        .dout(new_Jinkela_wire_10761)
    );

    bfr new_Jinkela_buffer_1645 (
        .din(new_Jinkela_wire_2540),
        .dout(new_Jinkela_wire_2541)
    );

    bfr new_Jinkela_buffer_8736 (
        .din(new_Jinkela_wire_10717),
        .dout(new_Jinkela_wire_10718)
    );

    bfr new_Jinkela_buffer_12209 (
        .din(new_Jinkela_wire_14706),
        .dout(new_Jinkela_wire_14707)
    );

    bfr new_Jinkela_buffer_1720 (
        .din(new_Jinkela_wire_2625),
        .dout(new_Jinkela_wire_2626)
    );

    bfr new_Jinkela_buffer_12155 (
        .din(new_Jinkela_wire_14632),
        .dout(new_Jinkela_wire_14633)
    );

    bfr new_Jinkela_buffer_1646 (
        .din(new_Jinkela_wire_2541),
        .dout(new_Jinkela_wire_2542)
    );

    spl2 new_Jinkela_splitter_850 (
        .a(_0096_),
        .b(new_Jinkela_wire_10971),
        .c(new_Jinkela_wire_10972)
    );

    bfr new_Jinkela_buffer_8737 (
        .din(new_Jinkela_wire_10718),
        .dout(new_Jinkela_wire_10719)
    );

    bfr new_Jinkela_buffer_12156 (
        .din(new_Jinkela_wire_14633),
        .dout(new_Jinkela_wire_14634)
    );

    bfr new_Jinkela_buffer_1897 (
        .din(_0584_),
        .dout(new_Jinkela_wire_2819)
    );

    bfr new_Jinkela_buffer_8774 (
        .din(new_Jinkela_wire_10761),
        .dout(new_Jinkela_wire_10762)
    );

    bfr new_Jinkela_buffer_1647 (
        .din(new_Jinkela_wire_2542),
        .dout(new_Jinkela_wire_2543)
    );

    spl2 new_Jinkela_splitter_1102 (
        .a(_0849_),
        .b(new_Jinkela_wire_15026),
        .c(new_Jinkela_wire_15027)
    );

    bfr new_Jinkela_buffer_8738 (
        .din(new_Jinkela_wire_10719),
        .dout(new_Jinkela_wire_10720)
    );

    bfr new_Jinkela_buffer_12210 (
        .din(new_Jinkela_wire_14707),
        .dout(new_Jinkela_wire_14708)
    );

    bfr new_Jinkela_buffer_1721 (
        .din(new_Jinkela_wire_2626),
        .dout(new_Jinkela_wire_2627)
    );

    bfr new_Jinkela_buffer_12157 (
        .din(new_Jinkela_wire_14634),
        .dout(new_Jinkela_wire_14635)
    );

    bfr new_Jinkela_buffer_8849 (
        .din(new_Jinkela_wire_10840),
        .dout(new_Jinkela_wire_10841)
    );

    bfr new_Jinkela_buffer_1648 (
        .din(new_Jinkela_wire_2543),
        .dout(new_Jinkela_wire_2544)
    );

    bfr new_Jinkela_buffer_8739 (
        .din(new_Jinkela_wire_10720),
        .dout(new_Jinkela_wire_10721)
    );

    bfr new_Jinkela_buffer_12284 (
        .din(new_Jinkela_wire_14783),
        .dout(new_Jinkela_wire_14784)
    );

    bfr new_Jinkela_buffer_1758 (
        .din(new_Jinkela_wire_2669),
        .dout(new_Jinkela_wire_2670)
    );

    bfr new_Jinkela_buffer_12158 (
        .din(new_Jinkela_wire_14635),
        .dout(new_Jinkela_wire_14636)
    );

    bfr new_Jinkela_buffer_8775 (
        .din(new_Jinkela_wire_10762),
        .dout(new_Jinkela_wire_10763)
    );

    bfr new_Jinkela_buffer_1649 (
        .din(new_Jinkela_wire_2544),
        .dout(new_Jinkela_wire_2545)
    );

    bfr new_Jinkela_buffer_8740 (
        .din(new_Jinkela_wire_10721),
        .dout(new_Jinkela_wire_10722)
    );

    bfr new_Jinkela_buffer_12211 (
        .din(new_Jinkela_wire_14708),
        .dout(new_Jinkela_wire_14709)
    );

    bfr new_Jinkela_buffer_1722 (
        .din(new_Jinkela_wire_2627),
        .dout(new_Jinkela_wire_2628)
    );

    bfr new_Jinkela_buffer_12159 (
        .din(new_Jinkela_wire_14636),
        .dout(new_Jinkela_wire_14637)
    );

    bfr new_Jinkela_buffer_8958 (
        .din(new_Jinkela_wire_10953),
        .dout(new_Jinkela_wire_10954)
    );

    bfr new_Jinkela_buffer_1650 (
        .din(new_Jinkela_wire_2545),
        .dout(new_Jinkela_wire_2546)
    );

    bfr new_Jinkela_buffer_8741 (
        .din(new_Jinkela_wire_10722),
        .dout(new_Jinkela_wire_10723)
    );

    bfr new_Jinkela_buffer_12393 (
        .din(new_Jinkela_wire_14894),
        .dout(new_Jinkela_wire_14895)
    );

    bfr new_Jinkela_buffer_1801 (
        .din(new_Jinkela_wire_2716),
        .dout(new_Jinkela_wire_2717)
    );

    bfr new_Jinkela_buffer_12160 (
        .din(new_Jinkela_wire_14637),
        .dout(new_Jinkela_wire_14638)
    );

    bfr new_Jinkela_buffer_8776 (
        .din(new_Jinkela_wire_10763),
        .dout(new_Jinkela_wire_10764)
    );

    bfr new_Jinkela_buffer_1651 (
        .din(new_Jinkela_wire_2546),
        .dout(new_Jinkela_wire_2547)
    );

    bfr new_Jinkela_buffer_8742 (
        .din(new_Jinkela_wire_10723),
        .dout(new_Jinkela_wire_10724)
    );

    bfr new_Jinkela_buffer_12212 (
        .din(new_Jinkela_wire_14709),
        .dout(new_Jinkela_wire_14710)
    );

    bfr new_Jinkela_buffer_1723 (
        .din(new_Jinkela_wire_2628),
        .dout(new_Jinkela_wire_2629)
    );

    bfr new_Jinkela_buffer_12161 (
        .din(new_Jinkela_wire_14638),
        .dout(new_Jinkela_wire_14639)
    );

    bfr new_Jinkela_buffer_8850 (
        .din(new_Jinkela_wire_10841),
        .dout(new_Jinkela_wire_10842)
    );

    bfr new_Jinkela_buffer_1652 (
        .din(new_Jinkela_wire_2547),
        .dout(new_Jinkela_wire_2548)
    );

    bfr new_Jinkela_buffer_8743 (
        .din(new_Jinkela_wire_10724),
        .dout(new_Jinkela_wire_10725)
    );

    bfr new_Jinkela_buffer_12285 (
        .din(new_Jinkela_wire_14784),
        .dout(new_Jinkela_wire_14785)
    );

    bfr new_Jinkela_buffer_1759 (
        .din(new_Jinkela_wire_2670),
        .dout(new_Jinkela_wire_2671)
    );

    bfr new_Jinkela_buffer_12162 (
        .din(new_Jinkela_wire_14639),
        .dout(new_Jinkela_wire_14640)
    );

    bfr new_Jinkela_buffer_8777 (
        .din(new_Jinkela_wire_10764),
        .dout(new_Jinkela_wire_10765)
    );

    bfr new_Jinkela_buffer_1653 (
        .din(new_Jinkela_wire_2548),
        .dout(new_Jinkela_wire_2549)
    );

    bfr new_Jinkela_buffer_8744 (
        .din(new_Jinkela_wire_10725),
        .dout(new_Jinkela_wire_10726)
    );

    bfr new_Jinkela_buffer_12213 (
        .din(new_Jinkela_wire_14710),
        .dout(new_Jinkela_wire_14711)
    );

    bfr new_Jinkela_buffer_1724 (
        .din(new_Jinkela_wire_2629),
        .dout(new_Jinkela_wire_2630)
    );

    bfr new_Jinkela_buffer_12163 (
        .din(new_Jinkela_wire_14640),
        .dout(new_Jinkela_wire_14641)
    );

    bfr new_Jinkela_buffer_8961 (
        .din(new_Jinkela_wire_10958),
        .dout(new_Jinkela_wire_10959)
    );

    bfr new_Jinkela_buffer_1654 (
        .din(new_Jinkela_wire_2549),
        .dout(new_Jinkela_wire_2550)
    );

    spl2 new_Jinkela_splitter_849 (
        .a(_0374_),
        .b(new_Jinkela_wire_10969),
        .c(new_Jinkela_wire_10970)
    );

    bfr new_Jinkela_buffer_8745 (
        .din(new_Jinkela_wire_10726),
        .dout(new_Jinkela_wire_10727)
    );

    bfr new_Jinkela_buffer_12488 (
        .din(new_Jinkela_wire_14991),
        .dout(new_Jinkela_wire_14992)
    );

    bfr new_Jinkela_buffer_12164 (
        .din(new_Jinkela_wire_14641),
        .dout(new_Jinkela_wire_14642)
    );

    bfr new_Jinkela_buffer_1898 (
        .din(_0529_),
        .dout(new_Jinkela_wire_2820)
    );

    bfr new_Jinkela_buffer_8778 (
        .din(new_Jinkela_wire_10765),
        .dout(new_Jinkela_wire_10766)
    );

    bfr new_Jinkela_buffer_1655 (
        .din(new_Jinkela_wire_2550),
        .dout(new_Jinkela_wire_2551)
    );

    bfr new_Jinkela_buffer_8746 (
        .din(new_Jinkela_wire_10727),
        .dout(new_Jinkela_wire_10728)
    );

    bfr new_Jinkela_buffer_12214 (
        .din(new_Jinkela_wire_14711),
        .dout(new_Jinkela_wire_14712)
    );

    bfr new_Jinkela_buffer_1725 (
        .din(new_Jinkela_wire_2630),
        .dout(new_Jinkela_wire_2631)
    );

    bfr new_Jinkela_buffer_12165 (
        .din(new_Jinkela_wire_14642),
        .dout(new_Jinkela_wire_14643)
    );

    bfr new_Jinkela_buffer_8851 (
        .din(new_Jinkela_wire_10842),
        .dout(new_Jinkela_wire_10843)
    );

    bfr new_Jinkela_buffer_1656 (
        .din(new_Jinkela_wire_2551),
        .dout(new_Jinkela_wire_2552)
    );

    bfr new_Jinkela_buffer_8747 (
        .din(new_Jinkela_wire_10728),
        .dout(new_Jinkela_wire_10729)
    );

    bfr new_Jinkela_buffer_12286 (
        .din(new_Jinkela_wire_14785),
        .dout(new_Jinkela_wire_14786)
    );

    bfr new_Jinkela_buffer_1760 (
        .din(new_Jinkela_wire_2671),
        .dout(new_Jinkela_wire_2672)
    );

    bfr new_Jinkela_buffer_12166 (
        .din(new_Jinkela_wire_14643),
        .dout(new_Jinkela_wire_14644)
    );

    or_ii _2791_ (
        .a(new_Jinkela_wire_20907),
        .b(new_Jinkela_wire_1011),
        .c(_0020_)
    );

    and_ii _2792_ (
        .a(new_Jinkela_wire_17065),
        .b(new_Jinkela_wire_14256),
        .c(_0021_)
    );

    and_bb _2793_ (
        .a(new_Jinkela_wire_17066),
        .b(new_Jinkela_wire_14257),
        .c(_0023_)
    );

    or_bb _2794_ (
        .a(new_Jinkela_wire_14288),
        .b(new_Jinkela_wire_3253),
        .c(_0024_)
    );

    or_bb _2795_ (
        .a(new_Jinkela_wire_7703),
        .b(new_Jinkela_wire_2592),
        .c(_0025_)
    );

    or_ii _2796_ (
        .a(new_Jinkela_wire_7704),
        .b(new_Jinkela_wire_2593),
        .c(_0026_)
    );

    or_ii _2797_ (
        .a(new_Jinkela_wire_13455),
        .b(new_Jinkela_wire_4702),
        .c(_0027_)
    );

    and_ii _2798_ (
        .a(new_Jinkela_wire_15672),
        .b(new_Jinkela_wire_2709),
        .c(_0028_)
    );

    and_bb _2799_ (
        .a(new_Jinkela_wire_15673),
        .b(new_Jinkela_wire_2710),
        .c(_0029_)
    );

    or_bb _2800_ (
        .a(new_Jinkela_wire_17423),
        .b(new_Jinkela_wire_18119),
        .c(_0030_)
    );

    or_bb _2801_ (
        .a(new_Jinkela_wire_3892),
        .b(new_Jinkela_wire_19126),
        .c(_0031_)
    );

    or_ii _2802_ (
        .a(new_Jinkela_wire_3893),
        .b(new_Jinkela_wire_19127),
        .c(_0032_)
    );

    or_ii _2803_ (
        .a(new_Jinkela_wire_13156),
        .b(new_Jinkela_wire_7445),
        .c(_0034_)
    );

    and_ii _2804_ (
        .a(new_Jinkela_wire_16866),
        .b(new_Jinkela_wire_1075),
        .c(_0035_)
    );

    and_bb _2805_ (
        .a(new_Jinkela_wire_16867),
        .b(new_Jinkela_wire_1076),
        .c(_0036_)
    );

    or_bb _2806_ (
        .a(new_Jinkela_wire_8294),
        .b(new_Jinkela_wire_16530),
        .c(_0037_)
    );

    or_bb _2807_ (
        .a(new_Jinkela_wire_12103),
        .b(new_Jinkela_wire_19045),
        .c(_0038_)
    );

    or_ii _2808_ (
        .a(new_Jinkela_wire_12104),
        .b(new_Jinkela_wire_19046),
        .c(_0039_)
    );

    or_ii _2809_ (
        .a(new_Jinkela_wire_5146),
        .b(new_Jinkela_wire_13333),
        .c(_0040_)
    );

    and_ii _2810_ (
        .a(new_Jinkela_wire_17013),
        .b(new_Jinkela_wire_7580),
        .c(_0041_)
    );

    and_bb _2811_ (
        .a(new_Jinkela_wire_17014),
        .b(new_Jinkela_wire_7581),
        .c(_0042_)
    );

    or_bb _2812_ (
        .a(new_Jinkela_wire_15893),
        .b(new_Jinkela_wire_4909),
        .c(_0043_)
    );

    or_bb _2813_ (
        .a(new_Jinkela_wire_10118),
        .b(new_Jinkela_wire_9097),
        .c(_0045_)
    );

    or_ii _2814_ (
        .a(new_Jinkela_wire_10119),
        .b(new_Jinkela_wire_9098),
        .c(_0046_)
    );

    or_ii _2815_ (
        .a(new_Jinkela_wire_5664),
        .b(new_Jinkela_wire_18566),
        .c(_0047_)
    );

    and_ii _2816_ (
        .a(new_Jinkela_wire_9175),
        .b(new_Jinkela_wire_13139),
        .c(_0048_)
    );

    and_bb _2817_ (
        .a(new_Jinkela_wire_9176),
        .b(new_Jinkela_wire_13140),
        .c(_0049_)
    );

    or_bb _2818_ (
        .a(new_Jinkela_wire_13966),
        .b(new_Jinkela_wire_13675),
        .c(_0050_)
    );

    or_bb _2819_ (
        .a(new_Jinkela_wire_8280),
        .b(new_Jinkela_wire_8841),
        .c(_0051_)
    );

    or_ii _2820_ (
        .a(new_Jinkela_wire_8281),
        .b(new_Jinkela_wire_8842),
        .c(_0052_)
    );

    or_ii _2821_ (
        .a(new_Jinkela_wire_8838),
        .b(new_Jinkela_wire_19328),
        .c(_0053_)
    );

    and_ii _2822_ (
        .a(new_Jinkela_wire_17985),
        .b(new_Jinkela_wire_14182),
        .c(_0054_)
    );

    and_bb _2823_ (
        .a(new_Jinkela_wire_17986),
        .b(new_Jinkela_wire_14183),
        .c(_0056_)
    );

    or_bb _2824_ (
        .a(new_Jinkela_wire_4666),
        .b(new_Jinkela_wire_17865),
        .c(_0057_)
    );

    or_bb _2825_ (
        .a(new_Jinkela_wire_8482),
        .b(new_Jinkela_wire_19052),
        .c(_0058_)
    );

    or_ii _2826_ (
        .a(new_Jinkela_wire_8483),
        .b(new_Jinkela_wire_19053),
        .c(_0059_)
    );

    or_ii _2827_ (
        .a(new_Jinkela_wire_18107),
        .b(new_Jinkela_wire_1791),
        .c(_0060_)
    );

    and_ii _2828_ (
        .a(new_Jinkela_wire_11614),
        .b(new_Jinkela_wire_8680),
        .c(_0061_)
    );

    and_bb _2829_ (
        .a(new_Jinkela_wire_11615),
        .b(new_Jinkela_wire_8681),
        .c(_0062_)
    );

    or_bb _2830_ (
        .a(new_Jinkela_wire_19785),
        .b(new_Jinkela_wire_13457),
        .c(_0063_)
    );

    or_bb _2831_ (
        .a(new_Jinkela_wire_18377),
        .b(new_Jinkela_wire_9347),
        .c(_0064_)
    );

    or_ii _2832_ (
        .a(new_Jinkela_wire_18378),
        .b(new_Jinkela_wire_9348),
        .c(_0065_)
    );

    bfr new_Jinkela_buffer_12215 (
        .din(new_Jinkela_wire_14712),
        .dout(new_Jinkela_wire_14713)
    );

    bfr new_Jinkela_buffer_12167 (
        .din(new_Jinkela_wire_14644),
        .dout(new_Jinkela_wire_14645)
    );

    bfr new_Jinkela_buffer_15627 (
        .din(new_Jinkela_wire_18625),
        .dout(new_Jinkela_wire_18626)
    );

    spl2 new_Jinkela_splitter_1360 (
        .a(_1489_),
        .b(new_Jinkela_wire_18791),
        .c(new_Jinkela_wire_18792)
    );

    bfr new_Jinkela_buffer_15709 (
        .din(new_Jinkela_wire_18719),
        .dout(new_Jinkela_wire_18720)
    );

    bfr new_Jinkela_buffer_12394 (
        .din(new_Jinkela_wire_14895),
        .dout(new_Jinkela_wire_14896)
    );

    bfr new_Jinkela_buffer_12168 (
        .din(new_Jinkela_wire_14645),
        .dout(new_Jinkela_wire_14646)
    );

    bfr new_Jinkela_buffer_15628 (
        .din(new_Jinkela_wire_18626),
        .dout(new_Jinkela_wire_18627)
    );

    bfr new_Jinkela_buffer_15727 (
        .din(new_Jinkela_wire_18739),
        .dout(new_Jinkela_wire_18740)
    );

    bfr new_Jinkela_buffer_12216 (
        .din(new_Jinkela_wire_14713),
        .dout(new_Jinkela_wire_14714)
    );

    bfr new_Jinkela_buffer_12169 (
        .din(new_Jinkela_wire_14646),
        .dout(new_Jinkela_wire_14647)
    );

    bfr new_Jinkela_buffer_15629 (
        .din(new_Jinkela_wire_18627),
        .dout(new_Jinkela_wire_18628)
    );

    bfr new_Jinkela_buffer_15710 (
        .din(new_Jinkela_wire_18720),
        .dout(new_Jinkela_wire_18721)
    );

    bfr new_Jinkela_buffer_12287 (
        .din(new_Jinkela_wire_14786),
        .dout(new_Jinkela_wire_14787)
    );

    bfr new_Jinkela_buffer_12170 (
        .din(new_Jinkela_wire_14647),
        .dout(new_Jinkela_wire_14648)
    );

    bfr new_Jinkela_buffer_15630 (
        .din(new_Jinkela_wire_18628),
        .dout(new_Jinkela_wire_18629)
    );

    bfr new_Jinkela_buffer_15747 (
        .din(new_Jinkela_wire_18765),
        .dout(new_Jinkela_wire_18766)
    );

    bfr new_Jinkela_buffer_12217 (
        .din(new_Jinkela_wire_14714),
        .dout(new_Jinkela_wire_14715)
    );

    bfr new_Jinkela_buffer_12171 (
        .din(new_Jinkela_wire_14648),
        .dout(new_Jinkela_wire_14649)
    );

    bfr new_Jinkela_buffer_15631 (
        .din(new_Jinkela_wire_18629),
        .dout(new_Jinkela_wire_18630)
    );

    bfr new_Jinkela_buffer_15711 (
        .din(new_Jinkela_wire_18721),
        .dout(new_Jinkela_wire_18722)
    );

    bfr new_Jinkela_buffer_12520 (
        .din(_0143_),
        .dout(new_Jinkela_wire_15028)
    );

    bfr new_Jinkela_buffer_12172 (
        .din(new_Jinkela_wire_14649),
        .dout(new_Jinkela_wire_14650)
    );

    bfr new_Jinkela_buffer_15632 (
        .din(new_Jinkela_wire_18630),
        .dout(new_Jinkela_wire_18631)
    );

    bfr new_Jinkela_buffer_15728 (
        .din(new_Jinkela_wire_18740),
        .dout(new_Jinkela_wire_18741)
    );

    bfr new_Jinkela_buffer_12218 (
        .din(new_Jinkela_wire_14715),
        .dout(new_Jinkela_wire_14716)
    );

    bfr new_Jinkela_buffer_12173 (
        .din(new_Jinkela_wire_14650),
        .dout(new_Jinkela_wire_14651)
    );

    bfr new_Jinkela_buffer_15633 (
        .din(new_Jinkela_wire_18631),
        .dout(new_Jinkela_wire_18632)
    );

    bfr new_Jinkela_buffer_15712 (
        .din(new_Jinkela_wire_18722),
        .dout(new_Jinkela_wire_18723)
    );

    bfr new_Jinkela_buffer_12288 (
        .din(new_Jinkela_wire_14787),
        .dout(new_Jinkela_wire_14788)
    );

    bfr new_Jinkela_buffer_12174 (
        .din(new_Jinkela_wire_14651),
        .dout(new_Jinkela_wire_14652)
    );

    bfr new_Jinkela_buffer_15634 (
        .din(new_Jinkela_wire_18632),
        .dout(new_Jinkela_wire_18633)
    );

    bfr new_Jinkela_buffer_15751 (
        .din(new_Jinkela_wire_18769),
        .dout(new_Jinkela_wire_18770)
    );

    bfr new_Jinkela_buffer_12219 (
        .din(new_Jinkela_wire_14716),
        .dout(new_Jinkela_wire_14717)
    );

    bfr new_Jinkela_buffer_12175 (
        .din(new_Jinkela_wire_14652),
        .dout(new_Jinkela_wire_14653)
    );

    bfr new_Jinkela_buffer_15635 (
        .din(new_Jinkela_wire_18633),
        .dout(new_Jinkela_wire_18634)
    );

    bfr new_Jinkela_buffer_15713 (
        .din(new_Jinkela_wire_18723),
        .dout(new_Jinkela_wire_18724)
    );

    bfr new_Jinkela_buffer_12395 (
        .din(new_Jinkela_wire_14896),
        .dout(new_Jinkela_wire_14897)
    );

    bfr new_Jinkela_buffer_12176 (
        .din(new_Jinkela_wire_14653),
        .dout(new_Jinkela_wire_14654)
    );

    bfr new_Jinkela_buffer_15636 (
        .din(new_Jinkela_wire_18634),
        .dout(new_Jinkela_wire_18635)
    );

    bfr new_Jinkela_buffer_15729 (
        .din(new_Jinkela_wire_18741),
        .dout(new_Jinkela_wire_18742)
    );

    bfr new_Jinkela_buffer_12220 (
        .din(new_Jinkela_wire_14717),
        .dout(new_Jinkela_wire_14718)
    );

    bfr new_Jinkela_buffer_12177 (
        .din(new_Jinkela_wire_14654),
        .dout(new_Jinkela_wire_14655)
    );

    bfr new_Jinkela_buffer_15637 (
        .din(new_Jinkela_wire_18635),
        .dout(new_Jinkela_wire_18636)
    );

    bfr new_Jinkela_buffer_15714 (
        .din(new_Jinkela_wire_18724),
        .dout(new_Jinkela_wire_18725)
    );

    bfr new_Jinkela_buffer_12289 (
        .din(new_Jinkela_wire_14788),
        .dout(new_Jinkela_wire_14789)
    );

    bfr new_Jinkela_buffer_15638 (
        .din(new_Jinkela_wire_18636),
        .dout(new_Jinkela_wire_18637)
    );

    bfr new_Jinkela_buffer_12221 (
        .din(new_Jinkela_wire_14718),
        .dout(new_Jinkela_wire_14719)
    );

    bfr new_Jinkela_buffer_15748 (
        .din(new_Jinkela_wire_18766),
        .dout(new_Jinkela_wire_18767)
    );

    bfr new_Jinkela_buffer_12489 (
        .din(new_Jinkela_wire_14992),
        .dout(new_Jinkela_wire_14993)
    );

    bfr new_Jinkela_buffer_15639 (
        .din(new_Jinkela_wire_18637),
        .dout(new_Jinkela_wire_18638)
    );

    bfr new_Jinkela_buffer_12222 (
        .din(new_Jinkela_wire_14719),
        .dout(new_Jinkela_wire_14720)
    );

    bfr new_Jinkela_buffer_15715 (
        .din(new_Jinkela_wire_18725),
        .dout(new_Jinkela_wire_18726)
    );

    bfr new_Jinkela_buffer_12290 (
        .din(new_Jinkela_wire_14789),
        .dout(new_Jinkela_wire_14790)
    );

    bfr new_Jinkela_buffer_15640 (
        .din(new_Jinkela_wire_18638),
        .dout(new_Jinkela_wire_18639)
    );

    bfr new_Jinkela_buffer_12223 (
        .din(new_Jinkela_wire_14720),
        .dout(new_Jinkela_wire_14721)
    );

    bfr new_Jinkela_buffer_15730 (
        .din(new_Jinkela_wire_18742),
        .dout(new_Jinkela_wire_18743)
    );

    bfr new_Jinkela_buffer_12396 (
        .din(new_Jinkela_wire_14897),
        .dout(new_Jinkela_wire_14898)
    );

    bfr new_Jinkela_buffer_15641 (
        .din(new_Jinkela_wire_18639),
        .dout(new_Jinkela_wire_18640)
    );

    bfr new_Jinkela_buffer_12224 (
        .din(new_Jinkela_wire_14721),
        .dout(new_Jinkela_wire_14722)
    );

    bfr new_Jinkela_buffer_15716 (
        .din(new_Jinkela_wire_18726),
        .dout(new_Jinkela_wire_18727)
    );

    bfr new_Jinkela_buffer_12291 (
        .din(new_Jinkela_wire_14790),
        .dout(new_Jinkela_wire_14791)
    );

    bfr new_Jinkela_buffer_15642 (
        .din(new_Jinkela_wire_18640),
        .dout(new_Jinkela_wire_18641)
    );

    bfr new_Jinkela_buffer_12225 (
        .din(new_Jinkela_wire_14722),
        .dout(new_Jinkela_wire_14723)
    );

    bfr new_Jinkela_buffer_12521 (
        .din(_0536_),
        .dout(new_Jinkela_wire_15029)
    );

    bfr new_Jinkela_buffer_15643 (
        .din(new_Jinkela_wire_18641),
        .dout(new_Jinkela_wire_18642)
    );

    bfr new_Jinkela_buffer_12226 (
        .din(new_Jinkela_wire_14723),
        .dout(new_Jinkela_wire_14724)
    );

    bfr new_Jinkela_buffer_15764 (
        .din(new_Jinkela_wire_18786),
        .dout(new_Jinkela_wire_18787)
    );

    bfr new_Jinkela_buffer_15717 (
        .din(new_Jinkela_wire_18727),
        .dout(new_Jinkela_wire_18728)
    );

    bfr new_Jinkela_buffer_12292 (
        .din(new_Jinkela_wire_14791),
        .dout(new_Jinkela_wire_14792)
    );

    bfr new_Jinkela_buffer_15644 (
        .din(new_Jinkela_wire_18642),
        .dout(new_Jinkela_wire_18643)
    );

    bfr new_Jinkela_buffer_12227 (
        .din(new_Jinkela_wire_14724),
        .dout(new_Jinkela_wire_14725)
    );

    bfr new_Jinkela_buffer_15731 (
        .din(new_Jinkela_wire_18743),
        .dout(new_Jinkela_wire_18744)
    );

    bfr new_Jinkela_buffer_12397 (
        .din(new_Jinkela_wire_14898),
        .dout(new_Jinkela_wire_14899)
    );

    bfr new_Jinkela_buffer_15645 (
        .din(new_Jinkela_wire_18643),
        .dout(new_Jinkela_wire_18644)
    );

    bfr new_Jinkela_buffer_12228 (
        .din(new_Jinkela_wire_14725),
        .dout(new_Jinkela_wire_14726)
    );

    bfr new_Jinkela_buffer_15718 (
        .din(new_Jinkela_wire_18728),
        .dout(new_Jinkela_wire_18729)
    );

    bfr new_Jinkela_buffer_12293 (
        .din(new_Jinkela_wire_14792),
        .dout(new_Jinkela_wire_14793)
    );

    bfr new_Jinkela_buffer_15646 (
        .din(new_Jinkela_wire_18644),
        .dout(new_Jinkela_wire_18645)
    );

    bfr new_Jinkela_buffer_12229 (
        .din(new_Jinkela_wire_14726),
        .dout(new_Jinkela_wire_14727)
    );

    bfr new_Jinkela_buffer_15749 (
        .din(new_Jinkela_wire_18767),
        .dout(new_Jinkela_wire_18768)
    );

    bfr new_Jinkela_buffer_12490 (
        .din(new_Jinkela_wire_14993),
        .dout(new_Jinkela_wire_14994)
    );

    bfr new_Jinkela_buffer_15647 (
        .din(new_Jinkela_wire_18645),
        .dout(new_Jinkela_wire_18646)
    );

    bfr new_Jinkela_buffer_1657 (
        .din(new_Jinkela_wire_2552),
        .dout(new_Jinkela_wire_2553)
    );

    bfr new_Jinkela_buffer_1726 (
        .din(new_Jinkela_wire_2631),
        .dout(new_Jinkela_wire_2632)
    );

    bfr new_Jinkela_buffer_1658 (
        .din(new_Jinkela_wire_2553),
        .dout(new_Jinkela_wire_2554)
    );

    bfr new_Jinkela_buffer_1802 (
        .din(new_Jinkela_wire_2717),
        .dout(new_Jinkela_wire_2718)
    );

    bfr new_Jinkela_buffer_1659 (
        .din(new_Jinkela_wire_2554),
        .dout(new_Jinkela_wire_2555)
    );

    bfr new_Jinkela_buffer_1727 (
        .din(new_Jinkela_wire_2632),
        .dout(new_Jinkela_wire_2633)
    );

    bfr new_Jinkela_buffer_1660 (
        .din(new_Jinkela_wire_2555),
        .dout(new_Jinkela_wire_2556)
    );

    bfr new_Jinkela_buffer_1761 (
        .din(new_Jinkela_wire_2672),
        .dout(new_Jinkela_wire_2673)
    );

    bfr new_Jinkela_buffer_1661 (
        .din(new_Jinkela_wire_2556),
        .dout(new_Jinkela_wire_2557)
    );

    bfr new_Jinkela_buffer_1728 (
        .din(new_Jinkela_wire_2633),
        .dout(new_Jinkela_wire_2634)
    );

    bfr new_Jinkela_buffer_1662 (
        .din(new_Jinkela_wire_2557),
        .dout(new_Jinkela_wire_2558)
    );

    bfr new_Jinkela_buffer_2010 (
        .din(_1792_),
        .dout(new_Jinkela_wire_2934)
    );

    bfr new_Jinkela_buffer_1871 (
        .din(new_Jinkela_wire_2792),
        .dout(new_Jinkela_wire_2793)
    );

    bfr new_Jinkela_buffer_1663 (
        .din(new_Jinkela_wire_2558),
        .dout(new_Jinkela_wire_2559)
    );

    bfr new_Jinkela_buffer_1729 (
        .din(new_Jinkela_wire_2634),
        .dout(new_Jinkela_wire_2635)
    );

    bfr new_Jinkela_buffer_1664 (
        .din(new_Jinkela_wire_2559),
        .dout(new_Jinkela_wire_2560)
    );

    bfr new_Jinkela_buffer_1762 (
        .din(new_Jinkela_wire_2673),
        .dout(new_Jinkela_wire_2674)
    );

    bfr new_Jinkela_buffer_1665 (
        .din(new_Jinkela_wire_2560),
        .dout(new_Jinkela_wire_2561)
    );

    bfr new_Jinkela_buffer_1730 (
        .din(new_Jinkela_wire_2635),
        .dout(new_Jinkela_wire_2636)
    );

    bfr new_Jinkela_buffer_1666 (
        .din(new_Jinkela_wire_2561),
        .dout(new_Jinkela_wire_2562)
    );

    bfr new_Jinkela_buffer_1803 (
        .din(new_Jinkela_wire_2718),
        .dout(new_Jinkela_wire_2719)
    );

    bfr new_Jinkela_buffer_1667 (
        .din(new_Jinkela_wire_2562),
        .dout(new_Jinkela_wire_2563)
    );

    bfr new_Jinkela_buffer_1731 (
        .din(new_Jinkela_wire_2636),
        .dout(new_Jinkela_wire_2637)
    );

    bfr new_Jinkela_buffer_1668 (
        .din(new_Jinkela_wire_2563),
        .dout(new_Jinkela_wire_2564)
    );

    bfr new_Jinkela_buffer_1763 (
        .din(new_Jinkela_wire_2674),
        .dout(new_Jinkela_wire_2675)
    );

    bfr new_Jinkela_buffer_1669 (
        .din(new_Jinkela_wire_2564),
        .dout(new_Jinkela_wire_2565)
    );

    bfr new_Jinkela_buffer_1732 (
        .din(new_Jinkela_wire_2637),
        .dout(new_Jinkela_wire_2638)
    );

    bfr new_Jinkela_buffer_1670 (
        .din(new_Jinkela_wire_2565),
        .dout(new_Jinkela_wire_2566)
    );

    bfr new_Jinkela_buffer_1671 (
        .din(new_Jinkela_wire_2566),
        .dout(new_Jinkela_wire_2567)
    );

    bfr new_Jinkela_buffer_1733 (
        .din(new_Jinkela_wire_2638),
        .dout(new_Jinkela_wire_2639)
    );

    bfr new_Jinkela_buffer_1672 (
        .din(new_Jinkela_wire_2567),
        .dout(new_Jinkela_wire_2568)
    );

    bfr new_Jinkela_buffer_1764 (
        .din(new_Jinkela_wire_2675),
        .dout(new_Jinkela_wire_2676)
    );

    bfr new_Jinkela_buffer_1673 (
        .din(new_Jinkela_wire_2568),
        .dout(new_Jinkela_wire_2569)
    );

    bfr new_Jinkela_buffer_1734 (
        .din(new_Jinkela_wire_2639),
        .dout(new_Jinkela_wire_2640)
    );

    bfr new_Jinkela_buffer_1674 (
        .din(new_Jinkela_wire_2569),
        .dout(new_Jinkela_wire_2570)
    );

    bfr new_Jinkela_buffer_1804 (
        .din(new_Jinkela_wire_2719),
        .dout(new_Jinkela_wire_2720)
    );

    bfr new_Jinkela_buffer_1675 (
        .din(new_Jinkela_wire_2570),
        .dout(new_Jinkela_wire_2571)
    );

    bfr new_Jinkela_buffer_1735 (
        .din(new_Jinkela_wire_2640),
        .dout(new_Jinkela_wire_2641)
    );

    bfr new_Jinkela_buffer_1676 (
        .din(new_Jinkela_wire_2571),
        .dout(new_Jinkela_wire_2572)
    );

    bfr new_Jinkela_buffer_1765 (
        .din(new_Jinkela_wire_2676),
        .dout(new_Jinkela_wire_2677)
    );

    bfr new_Jinkela_buffer_1677 (
        .din(new_Jinkela_wire_2572),
        .dout(new_Jinkela_wire_2573)
    );

    bfr new_Jinkela_buffer_1736 (
        .din(new_Jinkela_wire_2641),
        .dout(new_Jinkela_wire_2642)
    );

    bfr new_Jinkela_buffer_5273 (
        .din(new_Jinkela_wire_6778),
        .dout(new_Jinkela_wire_6779)
    );

    bfr new_Jinkela_buffer_5328 (
        .din(new_Jinkela_wire_6849),
        .dout(new_Jinkela_wire_6850)
    );

    bfr new_Jinkela_buffer_5274 (
        .din(new_Jinkela_wire_6779),
        .dout(new_Jinkela_wire_6780)
    );

    bfr new_Jinkela_buffer_5299 (
        .din(new_Jinkela_wire_6814),
        .dout(new_Jinkela_wire_6815)
    );

    bfr new_Jinkela_buffer_5275 (
        .din(new_Jinkela_wire_6780),
        .dout(new_Jinkela_wire_6781)
    );

    spl2 new_Jinkela_splitter_610 (
        .a(_1346_),
        .b(new_Jinkela_wire_6855),
        .c(new_Jinkela_wire_6856)
    );

    bfr new_Jinkela_buffer_5276 (
        .din(new_Jinkela_wire_6781),
        .dout(new_Jinkela_wire_6782)
    );

    bfr new_Jinkela_buffer_5300 (
        .din(new_Jinkela_wire_6815),
        .dout(new_Jinkela_wire_6816)
    );

    bfr new_Jinkela_buffer_5277 (
        .din(new_Jinkela_wire_6782),
        .dout(new_Jinkela_wire_6783)
    );

    spl2 new_Jinkela_splitter_611 (
        .a(_1390_),
        .b(new_Jinkela_wire_6857),
        .c(new_Jinkela_wire_6858)
    );

    bfr new_Jinkela_buffer_5278 (
        .din(new_Jinkela_wire_6783),
        .dout(new_Jinkela_wire_6784)
    );

    bfr new_Jinkela_buffer_5301 (
        .din(new_Jinkela_wire_6816),
        .dout(new_Jinkela_wire_6817)
    );

    bfr new_Jinkela_buffer_5279 (
        .din(new_Jinkela_wire_6784),
        .dout(new_Jinkela_wire_6785)
    );

    bfr new_Jinkela_buffer_5329 (
        .din(new_Jinkela_wire_6850),
        .dout(new_Jinkela_wire_6851)
    );

    bfr new_Jinkela_buffer_5280 (
        .din(new_Jinkela_wire_6785),
        .dout(new_Jinkela_wire_6786)
    );

    bfr new_Jinkela_buffer_5302 (
        .din(new_Jinkela_wire_6817),
        .dout(new_Jinkela_wire_6818)
    );

    bfr new_Jinkela_buffer_5281 (
        .din(new_Jinkela_wire_6786),
        .dout(new_Jinkela_wire_6787)
    );

    bfr new_Jinkela_buffer_5282 (
        .din(new_Jinkela_wire_6787),
        .dout(new_Jinkela_wire_6788)
    );

    bfr new_Jinkela_buffer_5303 (
        .din(new_Jinkela_wire_6818),
        .dout(new_Jinkela_wire_6819)
    );

    bfr new_Jinkela_buffer_5283 (
        .din(new_Jinkela_wire_6788),
        .dout(new_Jinkela_wire_6789)
    );

    bfr new_Jinkela_buffer_5330 (
        .din(new_Jinkela_wire_6851),
        .dout(new_Jinkela_wire_6852)
    );

    bfr new_Jinkela_buffer_5284 (
        .din(new_Jinkela_wire_6789),
        .dout(new_Jinkela_wire_6790)
    );

    bfr new_Jinkela_buffer_5304 (
        .din(new_Jinkela_wire_6819),
        .dout(new_Jinkela_wire_6820)
    );

    bfr new_Jinkela_buffer_5285 (
        .din(new_Jinkela_wire_6790),
        .dout(new_Jinkela_wire_6791)
    );

    spl2 new_Jinkela_splitter_612 (
        .a(_1020_),
        .b(new_Jinkela_wire_6859),
        .c(new_Jinkela_wire_6860)
    );

    bfr new_Jinkela_buffer_5286 (
        .din(new_Jinkela_wire_6791),
        .dout(new_Jinkela_wire_6792)
    );

    bfr new_Jinkela_buffer_5305 (
        .din(new_Jinkela_wire_6820),
        .dout(new_Jinkela_wire_6821)
    );

    bfr new_Jinkela_buffer_5287 (
        .din(new_Jinkela_wire_6792),
        .dout(new_Jinkela_wire_6793)
    );

    bfr new_Jinkela_buffer_5331 (
        .din(new_Jinkela_wire_6852),
        .dout(new_Jinkela_wire_6853)
    );

    bfr new_Jinkela_buffer_5288 (
        .din(new_Jinkela_wire_6793),
        .dout(new_Jinkela_wire_6794)
    );

    bfr new_Jinkela_buffer_5306 (
        .din(new_Jinkela_wire_6821),
        .dout(new_Jinkela_wire_6822)
    );

    bfr new_Jinkela_buffer_5289 (
        .din(new_Jinkela_wire_6794),
        .dout(new_Jinkela_wire_6795)
    );

    spl2 new_Jinkela_splitter_614 (
        .a(_0940_),
        .b(new_Jinkela_wire_6960),
        .c(new_Jinkela_wire_6961)
    );

    bfr new_Jinkela_buffer_5333 (
        .din(_1452_),
        .dout(new_Jinkela_wire_6861)
    );

    bfr new_Jinkela_buffer_5290 (
        .din(new_Jinkela_wire_6795),
        .dout(new_Jinkela_wire_6796)
    );

    bfr new_Jinkela_buffer_5307 (
        .din(new_Jinkela_wire_6822),
        .dout(new_Jinkela_wire_6823)
    );

    bfr new_Jinkela_buffer_5291 (
        .din(new_Jinkela_wire_6796),
        .dout(new_Jinkela_wire_6797)
    );

    bfr new_Jinkela_buffer_5429 (
        .din(_1644_),
        .dout(new_Jinkela_wire_6959)
    );

    bfr new_Jinkela_buffer_5292 (
        .din(new_Jinkela_wire_6797),
        .dout(new_Jinkela_wire_6798)
    );

    bfr new_Jinkela_buffer_5308 (
        .din(new_Jinkela_wire_6823),
        .dout(new_Jinkela_wire_6824)
    );

    bfr new_Jinkela_buffer_5293 (
        .din(new_Jinkela_wire_6798),
        .dout(new_Jinkela_wire_6799)
    );

    bfr new_Jinkela_buffer_5334 (
        .din(new_Jinkela_wire_6861),
        .dout(new_Jinkela_wire_6862)
    );

    bfr new_Jinkela_buffer_8779 (
        .din(new_Jinkela_wire_10766),
        .dout(new_Jinkela_wire_10767)
    );

    bfr new_Jinkela_buffer_8748 (
        .din(new_Jinkela_wire_10729),
        .dout(new_Jinkela_wire_10730)
    );

    bfr new_Jinkela_buffer_8959 (
        .din(new_Jinkela_wire_10954),
        .dout(new_Jinkela_wire_10955)
    );

    bfr new_Jinkela_buffer_8749 (
        .din(new_Jinkela_wire_10730),
        .dout(new_Jinkela_wire_10731)
    );

    bfr new_Jinkela_buffer_8780 (
        .din(new_Jinkela_wire_10767),
        .dout(new_Jinkela_wire_10768)
    );

    bfr new_Jinkela_buffer_8750 (
        .din(new_Jinkela_wire_10731),
        .dout(new_Jinkela_wire_10732)
    );

    bfr new_Jinkela_buffer_8852 (
        .din(new_Jinkela_wire_10843),
        .dout(new_Jinkela_wire_10844)
    );

    bfr new_Jinkela_buffer_8751 (
        .din(new_Jinkela_wire_10732),
        .dout(new_Jinkela_wire_10733)
    );

    bfr new_Jinkela_buffer_8781 (
        .din(new_Jinkela_wire_10768),
        .dout(new_Jinkela_wire_10769)
    );

    bfr new_Jinkela_buffer_8752 (
        .din(new_Jinkela_wire_10733),
        .dout(new_Jinkela_wire_10734)
    );

    bfr new_Jinkela_buffer_8753 (
        .din(new_Jinkela_wire_10734),
        .dout(new_Jinkela_wire_10735)
    );

    bfr new_Jinkela_buffer_8782 (
        .din(new_Jinkela_wire_10769),
        .dout(new_Jinkela_wire_10770)
    );

    bfr new_Jinkela_buffer_8754 (
        .din(new_Jinkela_wire_10735),
        .dout(new_Jinkela_wire_10736)
    );

    bfr new_Jinkela_buffer_8853 (
        .din(new_Jinkela_wire_10844),
        .dout(new_Jinkela_wire_10845)
    );

    bfr new_Jinkela_buffer_8755 (
        .din(new_Jinkela_wire_10736),
        .dout(new_Jinkela_wire_10737)
    );

    bfr new_Jinkela_buffer_8783 (
        .din(new_Jinkela_wire_10770),
        .dout(new_Jinkela_wire_10771)
    );

    bfr new_Jinkela_buffer_8756 (
        .din(new_Jinkela_wire_10737),
        .dout(new_Jinkela_wire_10738)
    );

    bfr new_Jinkela_buffer_8960 (
        .din(new_Jinkela_wire_10955),
        .dout(new_Jinkela_wire_10956)
    );

    bfr new_Jinkela_buffer_8757 (
        .din(new_Jinkela_wire_10738),
        .dout(new_Jinkela_wire_10739)
    );

    bfr new_Jinkela_buffer_8784 (
        .din(new_Jinkela_wire_10771),
        .dout(new_Jinkela_wire_10772)
    );

    bfr new_Jinkela_buffer_8758 (
        .din(new_Jinkela_wire_10739),
        .dout(new_Jinkela_wire_10740)
    );

    bfr new_Jinkela_buffer_8854 (
        .din(new_Jinkela_wire_10845),
        .dout(new_Jinkela_wire_10846)
    );

    bfr new_Jinkela_buffer_8759 (
        .din(new_Jinkela_wire_10740),
        .dout(new_Jinkela_wire_10741)
    );

    bfr new_Jinkela_buffer_8785 (
        .din(new_Jinkela_wire_10772),
        .dout(new_Jinkela_wire_10773)
    );

    bfr new_Jinkela_buffer_8760 (
        .din(new_Jinkela_wire_10741),
        .dout(new_Jinkela_wire_10742)
    );

    bfr new_Jinkela_buffer_8962 (
        .din(new_Jinkela_wire_10959),
        .dout(new_Jinkela_wire_10960)
    );

    spl2 new_Jinkela_splitter_840 (
        .a(new_Jinkela_wire_10742),
        .b(new_Jinkela_wire_10743),
        .c(new_Jinkela_wire_10744)
    );

    bfr new_Jinkela_buffer_8855 (
        .din(new_Jinkela_wire_10846),
        .dout(new_Jinkela_wire_10847)
    );

    bfr new_Jinkela_buffer_8786 (
        .din(new_Jinkela_wire_10773),
        .dout(new_Jinkela_wire_10774)
    );

    bfr new_Jinkela_buffer_8787 (
        .din(new_Jinkela_wire_10774),
        .dout(new_Jinkela_wire_10775)
    );

    spl2 new_Jinkela_splitter_851 (
        .a(_1674_),
        .b(new_Jinkela_wire_10973),
        .c(new_Jinkela_wire_10974)
    );

    bfr new_Jinkela_buffer_8788 (
        .din(new_Jinkela_wire_10775),
        .dout(new_Jinkela_wire_10776)
    );

    bfr new_Jinkela_buffer_8856 (
        .din(new_Jinkela_wire_10847),
        .dout(new_Jinkela_wire_10848)
    );

    bfr new_Jinkela_buffer_8789 (
        .din(new_Jinkela_wire_10776),
        .dout(new_Jinkela_wire_10777)
    );

    bfr new_Jinkela_buffer_8963 (
        .din(new_Jinkela_wire_10960),
        .dout(new_Jinkela_wire_10961)
    );

    bfr new_Jinkela_buffer_8790 (
        .din(new_Jinkela_wire_10777),
        .dout(new_Jinkela_wire_10778)
    );

    bfr new_Jinkela_buffer_8857 (
        .din(new_Jinkela_wire_10848),
        .dout(new_Jinkela_wire_10849)
    );

    bfr new_Jinkela_buffer_8791 (
        .din(new_Jinkela_wire_10778),
        .dout(new_Jinkela_wire_10779)
    );

    bfr new_Jinkela_buffer_8966 (
        .din(new_Jinkela_wire_10963),
        .dout(new_Jinkela_wire_10964)
    );

    bfr new_Jinkela_buffer_8965 (
        .din(_0641_),
        .dout(new_Jinkela_wire_10963)
    );

    bfr new_Jinkela_buffer_8792 (
        .din(new_Jinkela_wire_10779),
        .dout(new_Jinkela_wire_10780)
    );

    bfr new_Jinkela_buffer_8858 (
        .din(new_Jinkela_wire_10849),
        .dout(new_Jinkela_wire_10850)
    );

    bfr new_Jinkela_buffer_5294 (
        .din(new_Jinkela_wire_6799),
        .dout(new_Jinkela_wire_6800)
    );

    bfr new_Jinkela_buffer_1678 (
        .din(new_Jinkela_wire_2573),
        .dout(new_Jinkela_wire_2574)
    );

    bfr new_Jinkela_buffer_5309 (
        .din(new_Jinkela_wire_6824),
        .dout(new_Jinkela_wire_6825)
    );

    bfr new_Jinkela_buffer_15719 (
        .din(new_Jinkela_wire_18729),
        .dout(new_Jinkela_wire_18730)
    );

    bfr new_Jinkela_buffer_15648 (
        .din(new_Jinkela_wire_18646),
        .dout(new_Jinkela_wire_18647)
    );

    bfr new_Jinkela_buffer_1872 (
        .din(new_Jinkela_wire_2793),
        .dout(new_Jinkela_wire_2794)
    );

    bfr new_Jinkela_buffer_5295 (
        .din(new_Jinkela_wire_6800),
        .dout(new_Jinkela_wire_6801)
    );

    bfr new_Jinkela_buffer_1679 (
        .din(new_Jinkela_wire_2574),
        .dout(new_Jinkela_wire_2575)
    );

    bfr new_Jinkela_buffer_5434 (
        .din(_0761_),
        .dout(new_Jinkela_wire_6966)
    );

    bfr new_Jinkela_buffer_15732 (
        .din(new_Jinkela_wire_18744),
        .dout(new_Jinkela_wire_18745)
    );

    bfr new_Jinkela_buffer_1737 (
        .din(new_Jinkela_wire_2642),
        .dout(new_Jinkela_wire_2643)
    );

    bfr new_Jinkela_buffer_5430 (
        .din(new_Jinkela_wire_6961),
        .dout(new_Jinkela_wire_6962)
    );

    bfr new_Jinkela_buffer_15649 (
        .din(new_Jinkela_wire_18647),
        .dout(new_Jinkela_wire_18648)
    );

    spl2 new_Jinkela_splitter_602 (
        .a(new_Jinkela_wire_6801),
        .b(new_Jinkela_wire_6802),
        .c(new_Jinkela_wire_6803)
    );

    bfr new_Jinkela_buffer_1680 (
        .din(new_Jinkela_wire_2575),
        .dout(new_Jinkela_wire_2576)
    );

    bfr new_Jinkela_buffer_5335 (
        .din(new_Jinkela_wire_6862),
        .dout(new_Jinkela_wire_6863)
    );

    bfr new_Jinkela_buffer_15720 (
        .din(new_Jinkela_wire_18730),
        .dout(new_Jinkela_wire_18731)
    );

    bfr new_Jinkela_buffer_1766 (
        .din(new_Jinkela_wire_2677),
        .dout(new_Jinkela_wire_2678)
    );

    bfr new_Jinkela_buffer_15650 (
        .din(new_Jinkela_wire_18648),
        .dout(new_Jinkela_wire_18649)
    );

    bfr new_Jinkela_buffer_5310 (
        .din(new_Jinkela_wire_6825),
        .dout(new_Jinkela_wire_6826)
    );

    bfr new_Jinkela_buffer_1681 (
        .din(new_Jinkela_wire_2576),
        .dout(new_Jinkela_wire_2577)
    );

    bfr new_Jinkela_buffer_5311 (
        .din(new_Jinkela_wire_6826),
        .dout(new_Jinkela_wire_6827)
    );

    bfr new_Jinkela_buffer_15752 (
        .din(new_Jinkela_wire_18770),
        .dout(new_Jinkela_wire_18771)
    );

    bfr new_Jinkela_buffer_1738 (
        .din(new_Jinkela_wire_2643),
        .dout(new_Jinkela_wire_2644)
    );

    bfr new_Jinkela_buffer_15651 (
        .din(new_Jinkela_wire_18649),
        .dout(new_Jinkela_wire_18650)
    );

    bfr new_Jinkela_buffer_1682 (
        .din(new_Jinkela_wire_2577),
        .dout(new_Jinkela_wire_2578)
    );

    bfr new_Jinkela_buffer_5312 (
        .din(new_Jinkela_wire_6827),
        .dout(new_Jinkela_wire_6828)
    );

    spl2 new_Jinkela_splitter_1354 (
        .a(new_Jinkela_wire_18731),
        .b(new_Jinkela_wire_18732),
        .c(new_Jinkela_wire_18733)
    );

    bfr new_Jinkela_buffer_1805 (
        .din(new_Jinkela_wire_2720),
        .dout(new_Jinkela_wire_2721)
    );

    bfr new_Jinkela_buffer_15652 (
        .din(new_Jinkela_wire_18650),
        .dout(new_Jinkela_wire_18651)
    );

    bfr new_Jinkela_buffer_5336 (
        .din(new_Jinkela_wire_6863),
        .dout(new_Jinkela_wire_6864)
    );

    bfr new_Jinkela_buffer_1683 (
        .din(new_Jinkela_wire_2578),
        .dout(new_Jinkela_wire_2579)
    );

    bfr new_Jinkela_buffer_5313 (
        .din(new_Jinkela_wire_6828),
        .dout(new_Jinkela_wire_6829)
    );

    bfr new_Jinkela_buffer_1739 (
        .din(new_Jinkela_wire_2644),
        .dout(new_Jinkela_wire_2645)
    );

    bfr new_Jinkela_buffer_15653 (
        .din(new_Jinkela_wire_18651),
        .dout(new_Jinkela_wire_18652)
    );

    bfr new_Jinkela_buffer_1684 (
        .din(new_Jinkela_wire_2579),
        .dout(new_Jinkela_wire_2580)
    );

    spl2 new_Jinkela_splitter_616 (
        .a(_0894_),
        .b(new_Jinkela_wire_6992),
        .c(new_Jinkela_wire_6993)
    );

    bfr new_Jinkela_buffer_15772 (
        .din(_0587_),
        .dout(new_Jinkela_wire_18797)
    );

    bfr new_Jinkela_buffer_5314 (
        .din(new_Jinkela_wire_6829),
        .dout(new_Jinkela_wire_6830)
    );

    bfr new_Jinkela_buffer_15733 (
        .din(new_Jinkela_wire_18745),
        .dout(new_Jinkela_wire_18746)
    );

    bfr new_Jinkela_buffer_1767 (
        .din(new_Jinkela_wire_2678),
        .dout(new_Jinkela_wire_2679)
    );

    bfr new_Jinkela_buffer_15654 (
        .din(new_Jinkela_wire_18652),
        .dout(new_Jinkela_wire_18653)
    );

    bfr new_Jinkela_buffer_5337 (
        .din(new_Jinkela_wire_6864),
        .dout(new_Jinkela_wire_6865)
    );

    bfr new_Jinkela_buffer_1685 (
        .din(new_Jinkela_wire_2580),
        .dout(new_Jinkela_wire_2581)
    );

    bfr new_Jinkela_buffer_5315 (
        .din(new_Jinkela_wire_6830),
        .dout(new_Jinkela_wire_6831)
    );

    bfr new_Jinkela_buffer_15734 (
        .din(new_Jinkela_wire_18746),
        .dout(new_Jinkela_wire_18747)
    );

    bfr new_Jinkela_buffer_1740 (
        .din(new_Jinkela_wire_2645),
        .dout(new_Jinkela_wire_2646)
    );

    bfr new_Jinkela_buffer_15655 (
        .din(new_Jinkela_wire_18653),
        .dout(new_Jinkela_wire_18654)
    );

    bfr new_Jinkela_buffer_1686 (
        .din(new_Jinkela_wire_2581),
        .dout(new_Jinkela_wire_2582)
    );

    bfr new_Jinkela_buffer_5458 (
        .din(_1034_),
        .dout(new_Jinkela_wire_6994)
    );

    bfr new_Jinkela_buffer_5316 (
        .din(new_Jinkela_wire_6831),
        .dout(new_Jinkela_wire_6832)
    );

    bfr new_Jinkela_buffer_15753 (
        .din(new_Jinkela_wire_18771),
        .dout(new_Jinkela_wire_18772)
    );

    bfr new_Jinkela_buffer_15656 (
        .din(new_Jinkela_wire_18654),
        .dout(new_Jinkela_wire_18655)
    );

    spl2 new_Jinkela_splitter_311 (
        .a(_0246_),
        .b(new_Jinkela_wire_2935),
        .c(new_Jinkela_wire_2936)
    );

    bfr new_Jinkela_buffer_5338 (
        .din(new_Jinkela_wire_6865),
        .dout(new_Jinkela_wire_6866)
    );

    bfr new_Jinkela_buffer_1687 (
        .din(new_Jinkela_wire_2582),
        .dout(new_Jinkela_wire_2583)
    );

    bfr new_Jinkela_buffer_5317 (
        .din(new_Jinkela_wire_6832),
        .dout(new_Jinkela_wire_6833)
    );

    bfr new_Jinkela_buffer_15735 (
        .din(new_Jinkela_wire_18747),
        .dout(new_Jinkela_wire_18748)
    );

    bfr new_Jinkela_buffer_1741 (
        .din(new_Jinkela_wire_2646),
        .dout(new_Jinkela_wire_2647)
    );

    bfr new_Jinkela_buffer_15657 (
        .din(new_Jinkela_wire_18655),
        .dout(new_Jinkela_wire_18656)
    );

    bfr new_Jinkela_buffer_5431 (
        .din(new_Jinkela_wire_6962),
        .dout(new_Jinkela_wire_6963)
    );

    bfr new_Jinkela_buffer_1688 (
        .din(new_Jinkela_wire_2583),
        .dout(new_Jinkela_wire_2584)
    );

    bfr new_Jinkela_buffer_5318 (
        .din(new_Jinkela_wire_6833),
        .dout(new_Jinkela_wire_6834)
    );

    bfr new_Jinkela_buffer_1768 (
        .din(new_Jinkela_wire_2679),
        .dout(new_Jinkela_wire_2680)
    );

    bfr new_Jinkela_buffer_15658 (
        .din(new_Jinkela_wire_18656),
        .dout(new_Jinkela_wire_18657)
    );

    bfr new_Jinkela_buffer_5339 (
        .din(new_Jinkela_wire_6866),
        .dout(new_Jinkela_wire_6867)
    );

    bfr new_Jinkela_buffer_1689 (
        .din(new_Jinkela_wire_2584),
        .dout(new_Jinkela_wire_2585)
    );

    bfr new_Jinkela_buffer_5319 (
        .din(new_Jinkela_wire_6834),
        .dout(new_Jinkela_wire_6835)
    );

    bfr new_Jinkela_buffer_15736 (
        .din(new_Jinkela_wire_18748),
        .dout(new_Jinkela_wire_18749)
    );

    bfr new_Jinkela_buffer_1742 (
        .din(new_Jinkela_wire_2647),
        .dout(new_Jinkela_wire_2648)
    );

    bfr new_Jinkela_buffer_15659 (
        .din(new_Jinkela_wire_18657),
        .dout(new_Jinkela_wire_18658)
    );

    bfr new_Jinkela_buffer_5435 (
        .din(new_Jinkela_wire_6966),
        .dout(new_Jinkela_wire_6967)
    );

    bfr new_Jinkela_buffer_1690 (
        .din(new_Jinkela_wire_2585),
        .dout(new_Jinkela_wire_2586)
    );

    bfr new_Jinkela_buffer_5320 (
        .din(new_Jinkela_wire_6835),
        .dout(new_Jinkela_wire_6836)
    );

    bfr new_Jinkela_buffer_15754 (
        .din(new_Jinkela_wire_18772),
        .dout(new_Jinkela_wire_18773)
    );

    bfr new_Jinkela_buffer_1806 (
        .din(new_Jinkela_wire_2721),
        .dout(new_Jinkela_wire_2722)
    );

    bfr new_Jinkela_buffer_15660 (
        .din(new_Jinkela_wire_18658),
        .dout(new_Jinkela_wire_18659)
    );

    bfr new_Jinkela_buffer_5340 (
        .din(new_Jinkela_wire_6867),
        .dout(new_Jinkela_wire_6868)
    );

    bfr new_Jinkela_buffer_1691 (
        .din(new_Jinkela_wire_2586),
        .dout(new_Jinkela_wire_2587)
    );

    bfr new_Jinkela_buffer_5321 (
        .din(new_Jinkela_wire_6836),
        .dout(new_Jinkela_wire_6837)
    );

    bfr new_Jinkela_buffer_15737 (
        .din(new_Jinkela_wire_18749),
        .dout(new_Jinkela_wire_18750)
    );

    bfr new_Jinkela_buffer_1743 (
        .din(new_Jinkela_wire_2648),
        .dout(new_Jinkela_wire_2649)
    );

    bfr new_Jinkela_buffer_15661 (
        .din(new_Jinkela_wire_18659),
        .dout(new_Jinkela_wire_18660)
    );

    bfr new_Jinkela_buffer_5432 (
        .din(new_Jinkela_wire_6963),
        .dout(new_Jinkela_wire_6964)
    );

    bfr new_Jinkela_buffer_1692 (
        .din(new_Jinkela_wire_2587),
        .dout(new_Jinkela_wire_2588)
    );

    bfr new_Jinkela_buffer_5322 (
        .din(new_Jinkela_wire_6837),
        .dout(new_Jinkela_wire_6838)
    );

    bfr new_Jinkela_buffer_15765 (
        .din(new_Jinkela_wire_18787),
        .dout(new_Jinkela_wire_18788)
    );

    bfr new_Jinkela_buffer_1769 (
        .din(new_Jinkela_wire_2680),
        .dout(new_Jinkela_wire_2681)
    );

    bfr new_Jinkela_buffer_15662 (
        .din(new_Jinkela_wire_18660),
        .dout(new_Jinkela_wire_18661)
    );

    bfr new_Jinkela_buffer_5341 (
        .din(new_Jinkela_wire_6868),
        .dout(new_Jinkela_wire_6869)
    );

    spl2 new_Jinkela_splitter_297 (
        .a(new_Jinkela_wire_2588),
        .b(new_Jinkela_wire_2589),
        .c(new_Jinkela_wire_2590)
    );

    bfr new_Jinkela_buffer_5323 (
        .din(new_Jinkela_wire_6838),
        .dout(new_Jinkela_wire_6839)
    );

    bfr new_Jinkela_buffer_15738 (
        .din(new_Jinkela_wire_18750),
        .dout(new_Jinkela_wire_18751)
    );

    bfr new_Jinkela_buffer_1899 (
        .din(new_Jinkela_wire_2820),
        .dout(new_Jinkela_wire_2821)
    );

    bfr new_Jinkela_buffer_15663 (
        .din(new_Jinkela_wire_18661),
        .dout(new_Jinkela_wire_18662)
    );

    bfr new_Jinkela_buffer_1873 (
        .din(new_Jinkela_wire_2794),
        .dout(new_Jinkela_wire_2795)
    );

    bfr new_Jinkela_buffer_5459 (
        .din(_1207_),
        .dout(new_Jinkela_wire_6995)
    );

    bfr new_Jinkela_buffer_1744 (
        .din(new_Jinkela_wire_2649),
        .dout(new_Jinkela_wire_2650)
    );

    bfr new_Jinkela_buffer_5324 (
        .din(new_Jinkela_wire_6839),
        .dout(new_Jinkela_wire_6840)
    );

    bfr new_Jinkela_buffer_15755 (
        .din(new_Jinkela_wire_18773),
        .dout(new_Jinkela_wire_18774)
    );

    spl2 new_Jinkela_splitter_302 (
        .a(new_Jinkela_wire_2650),
        .b(new_Jinkela_wire_2651),
        .c(new_Jinkela_wire_2652)
    );

    bfr new_Jinkela_buffer_15664 (
        .din(new_Jinkela_wire_18662),
        .dout(new_Jinkela_wire_18663)
    );

    bfr new_Jinkela_buffer_5342 (
        .din(new_Jinkela_wire_6869),
        .dout(new_Jinkela_wire_6870)
    );

    bfr new_Jinkela_buffer_1807 (
        .din(new_Jinkela_wire_2722),
        .dout(new_Jinkela_wire_2723)
    );

    bfr new_Jinkela_buffer_5325 (
        .din(new_Jinkela_wire_6840),
        .dout(new_Jinkela_wire_6841)
    );

    bfr new_Jinkela_buffer_15739 (
        .din(new_Jinkela_wire_18751),
        .dout(new_Jinkela_wire_18752)
    );

    bfr new_Jinkela_buffer_1770 (
        .din(new_Jinkela_wire_2681),
        .dout(new_Jinkela_wire_2682)
    );

    bfr new_Jinkela_buffer_15665 (
        .din(new_Jinkela_wire_18663),
        .dout(new_Jinkela_wire_18664)
    );

    bfr new_Jinkela_buffer_5433 (
        .din(new_Jinkela_wire_6964),
        .dout(new_Jinkela_wire_6965)
    );

    bfr new_Jinkela_buffer_1771 (
        .din(new_Jinkela_wire_2682),
        .dout(new_Jinkela_wire_2683)
    );

    bfr new_Jinkela_buffer_5326 (
        .din(new_Jinkela_wire_6841),
        .dout(new_Jinkela_wire_6842)
    );

    bfr new_Jinkela_buffer_15768 (
        .din(new_Jinkela_wire_18792),
        .dout(new_Jinkela_wire_18793)
    );

    bfr new_Jinkela_buffer_15666 (
        .din(new_Jinkela_wire_18664),
        .dout(new_Jinkela_wire_18665)
    );

    bfr new_Jinkela_buffer_5343 (
        .din(new_Jinkela_wire_6870),
        .dout(new_Jinkela_wire_6871)
    );

    bfr new_Jinkela_buffer_1772 (
        .din(new_Jinkela_wire_2683),
        .dout(new_Jinkela_wire_2684)
    );

    spl2 new_Jinkela_splitter_1361 (
        .a(_1237_),
        .b(new_Jinkela_wire_18798),
        .c(new_Jinkela_wire_18799)
    );

    bfr new_Jinkela_buffer_5327 (
        .din(new_Jinkela_wire_6842),
        .dout(new_Jinkela_wire_6843)
    );

    bfr new_Jinkela_buffer_15740 (
        .din(new_Jinkela_wire_18752),
        .dout(new_Jinkela_wire_18753)
    );

    bfr new_Jinkela_buffer_1808 (
        .din(new_Jinkela_wire_2723),
        .dout(new_Jinkela_wire_2724)
    );

    bfr new_Jinkela_buffer_15667 (
        .din(new_Jinkela_wire_18665),
        .dout(new_Jinkela_wire_18666)
    );

    bfr new_Jinkela_buffer_5436 (
        .din(new_Jinkela_wire_6967),
        .dout(new_Jinkela_wire_6968)
    );

    bfr new_Jinkela_buffer_1773 (
        .din(new_Jinkela_wire_2684),
        .dout(new_Jinkela_wire_2685)
    );

    spl2 new_Jinkela_splitter_607 (
        .a(new_Jinkela_wire_6843),
        .b(new_Jinkela_wire_6844),
        .c(new_Jinkela_wire_6845)
    );

    bfr new_Jinkela_buffer_15756 (
        .din(new_Jinkela_wire_18774),
        .dout(new_Jinkela_wire_18775)
    );

    spl2 new_Jinkela_splitter_312 (
        .a(_0233_),
        .b(new_Jinkela_wire_2941),
        .c(new_Jinkela_wire_2942)
    );

    bfr new_Jinkela_buffer_15668 (
        .din(new_Jinkela_wire_18666),
        .dout(new_Jinkela_wire_18667)
    );

    or_ii _2833_ (
        .a(new_Jinkela_wire_20332),
        .b(new_Jinkela_wire_7130),
        .c(_0067_)
    );

    and_ii _2834_ (
        .a(new_Jinkela_wire_20373),
        .b(new_Jinkela_wire_14426),
        .c(_0068_)
    );

    and_bb _2835_ (
        .a(new_Jinkela_wire_20374),
        .b(new_Jinkela_wire_14427),
        .c(_0069_)
    );

    or_bb _2836_ (
        .a(new_Jinkela_wire_10060),
        .b(new_Jinkela_wire_15756),
        .c(_0070_)
    );

    or_bb _2837_ (
        .a(new_Jinkela_wire_19567),
        .b(new_Jinkela_wire_7512),
        .c(_0071_)
    );

    or_ii _2838_ (
        .a(new_Jinkela_wire_19568),
        .b(new_Jinkela_wire_7513),
        .c(_0072_)
    );

    or_ii _2839_ (
        .a(new_Jinkela_wire_15753),
        .b(new_Jinkela_wire_13005),
        .c(_0073_)
    );

    and_ii _2840_ (
        .a(new_Jinkela_wire_15124),
        .b(new_Jinkela_wire_4070),
        .c(_0074_)
    );

    and_bb _2841_ (
        .a(new_Jinkela_wire_15125),
        .b(new_Jinkela_wire_4071),
        .c(_0075_)
    );

    or_bb _2842_ (
        .a(new_Jinkela_wire_4838),
        .b(new_Jinkela_wire_5999),
        .c(_0076_)
    );

    or_bb _2843_ (
        .a(new_Jinkela_wire_15741),
        .b(new_Jinkela_wire_7182),
        .c(_0078_)
    );

    and_bb _2844_ (
        .a(new_Jinkela_wire_100),
        .b(new_Jinkela_wire_673),
        .c(_0079_)
    );

    or_ii _2845_ (
        .a(new_Jinkela_wire_15742),
        .b(new_Jinkela_wire_7183),
        .c(_0080_)
    );

    or_ii _2846_ (
        .a(new_Jinkela_wire_7844),
        .b(new_Jinkela_wire_7973),
        .c(_0081_)
    );

    and_ii _2847_ (
        .a(new_Jinkela_wire_16781),
        .b(new_Jinkela_wire_13844),
        .c(_0082_)
    );

    and_bi _2848_ (
        .a(new_Jinkela_wire_7978),
        .b(new_Jinkela_wire_7307),
        .c(_0083_)
    );

    and_bb _2849_ (
        .a(new_Jinkela_wire_664),
        .b(new_Jinkela_wire_561),
        .c(_0084_)
    );

    and_bi _2850_ (
        .a(new_Jinkela_wire_13010),
        .b(new_Jinkela_wire_6000),
        .c(_0085_)
    );

    and_bb _2851_ (
        .a(new_Jinkela_wire_279),
        .b(new_Jinkela_wire_517),
        .c(_0086_)
    );

    and_bi _2852_ (
        .a(new_Jinkela_wire_7135),
        .b(new_Jinkela_wire_15757),
        .c(_0087_)
    );

    and_bb _2853_ (
        .a(new_Jinkela_wire_73),
        .b(new_Jinkela_wire_130),
        .c(_0089_)
    );

    and_bi _2854_ (
        .a(new_Jinkela_wire_1796),
        .b(new_Jinkela_wire_13458),
        .c(_0090_)
    );

    and_bb _2855_ (
        .a(new_Jinkela_wire_474),
        .b(new_Jinkela_wire_219),
        .c(_0091_)
    );

    and_bi _2856_ (
        .a(new_Jinkela_wire_19333),
        .b(new_Jinkela_wire_17866),
        .c(_0092_)
    );

    and_bb _2857_ (
        .a(new_Jinkela_wire_360),
        .b(new_Jinkela_wire_593),
        .c(_0093_)
    );

    and_bi _2858_ (
        .a(new_Jinkela_wire_18571),
        .b(new_Jinkela_wire_13676),
        .c(_0094_)
    );

    and_bb _2859_ (
        .a(new_Jinkela_wire_701),
        .b(new_Jinkela_wire_111),
        .c(_0095_)
    );

    and_bi _2860_ (
        .a(new_Jinkela_wire_13338),
        .b(new_Jinkela_wire_4910),
        .c(_0096_)
    );

    and_bb _2861_ (
        .a(new_Jinkela_wire_19),
        .b(new_Jinkela_wire_498),
        .c(_0097_)
    );

    and_bi _2862_ (
        .a(new_Jinkela_wire_7450),
        .b(new_Jinkela_wire_16531),
        .c(_0098_)
    );

    and_bb _2863_ (
        .a(new_Jinkela_wire_458),
        .b(new_Jinkela_wire_27),
        .c(_0100_)
    );

    and_bi _2864_ (
        .a(new_Jinkela_wire_4707),
        .b(new_Jinkela_wire_18120),
        .c(_0101_)
    );

    and_bb _2865_ (
        .a(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_261),
        .c(_0102_)
    );

    and_bi _2866_ (
        .a(new_Jinkela_wire_1016),
        .b(new_Jinkela_wire_3254),
        .c(_0103_)
    );

    and_bb _2867_ (
        .a(new_Jinkela_wire_382),
        .b(new_Jinkela_wire_290),
        .c(_0104_)
    );

    and_bi _2868_ (
        .a(new_Jinkela_wire_5462),
        .b(new_Jinkela_wire_11446),
        .c(_0105_)
    );

    and_bb _2869_ (
        .a(new_Jinkela_wire_413),
        .b(new_Jinkela_wire_59),
        .c(_0106_)
    );

    and_bi _2870_ (
        .a(new_Jinkela_wire_17021),
        .b(new_Jinkela_wire_17029),
        .c(_0107_)
    );

    and_bb _2871_ (
        .a(new_Jinkela_wire_164),
        .b(new_Jinkela_wire_646),
        .c(_0108_)
    );

    and_bi _2872_ (
        .a(new_Jinkela_wire_18694),
        .b(new_Jinkela_wire_4996),
        .c(_0109_)
    );

    and_bb _2873_ (
        .a(new_Jinkela_wire_604),
        .b(new_Jinkela_wire_634),
        .c(_0111_)
    );

    and_bb _2874_ (
        .a(new_Jinkela_wire_429),
        .b(new_Jinkela_wire_538),
        .c(_0112_)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1553),
        .dout(new_Jinkela_wire_1554)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_net_3952),
        .dout(new_Jinkela_wire_1812)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1704),
        .dout(new_Jinkela_wire_1705)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1554),
        .dout(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1555),
        .dout(new_Jinkela_wire_1556)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1705),
        .dout(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1556),
        .dout(new_Jinkela_wire_1557)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1557),
        .dout(new_Jinkela_wire_1558)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(_0444_),
        .b(new_Jinkela_wire_1896),
        .c(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_1706),
        .dout(new_Jinkela_wire_1707)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1558),
        .dout(new_Jinkela_wire_1559)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_1559),
        .dout(new_Jinkela_wire_1560)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1707),
        .dout(new_Jinkela_wire_1708)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1560),
        .dout(new_Jinkela_wire_1561)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(_0299_),
        .b(new_Jinkela_wire_1898),
        .c(new_Jinkela_wire_1899)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_1708),
        .dout(new_Jinkela_wire_1709)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1709),
        .dout(new_Jinkela_wire_1710)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1564),
        .dout(new_Jinkela_wire_1565)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1565),
        .dout(new_Jinkela_wire_1566)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1710),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1711),
        .dout(new_Jinkela_wire_1712)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1712),
        .dout(new_Jinkela_wire_1713)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1713),
        .dout(new_Jinkela_wire_1714)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1814),
        .dout(new_Jinkela_wire_1815)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1714),
        .dout(new_Jinkela_wire_1715)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(_0537_),
        .b(new_Jinkela_wire_1904),
        .c(new_Jinkela_wire_1905)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1715),
        .dout(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_1899),
        .dout(new_Jinkela_wire_1900)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1815),
        .dout(new_Jinkela_wire_1816)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1716),
        .dout(new_Jinkela_wire_1717)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(_1326_),
        .b(new_Jinkela_wire_1906),
        .c(new_Jinkela_wire_1907)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1717),
        .dout(new_Jinkela_wire_1718)
    );

    bfr new_Jinkela_buffer_7919 (
        .din(new_Jinkela_wire_9786),
        .dout(new_Jinkela_wire_9787)
    );

    bfr new_Jinkela_buffer_7993 (
        .din(new_Jinkela_wire_9872),
        .dout(new_Jinkela_wire_9873)
    );

    bfr new_Jinkela_buffer_7920 (
        .din(new_Jinkela_wire_9787),
        .dout(new_Jinkela_wire_9788)
    );

    bfr new_Jinkela_buffer_7956 (
        .din(new_Jinkela_wire_9827),
        .dout(new_Jinkela_wire_9828)
    );

    bfr new_Jinkela_buffer_7921 (
        .din(new_Jinkela_wire_9788),
        .dout(new_Jinkela_wire_9789)
    );

    bfr new_Jinkela_buffer_8030 (
        .din(new_Jinkela_wire_9911),
        .dout(new_Jinkela_wire_9912)
    );

    bfr new_Jinkela_buffer_7922 (
        .din(new_Jinkela_wire_9789),
        .dout(new_Jinkela_wire_9790)
    );

    bfr new_Jinkela_buffer_7957 (
        .din(new_Jinkela_wire_9828),
        .dout(new_Jinkela_wire_9829)
    );

    bfr new_Jinkela_buffer_7923 (
        .din(new_Jinkela_wire_9790),
        .dout(new_Jinkela_wire_9791)
    );

    bfr new_Jinkela_buffer_7994 (
        .din(new_Jinkela_wire_9873),
        .dout(new_Jinkela_wire_9874)
    );

    bfr new_Jinkela_buffer_7924 (
        .din(new_Jinkela_wire_9791),
        .dout(new_Jinkela_wire_9792)
    );

    bfr new_Jinkela_buffer_7958 (
        .din(new_Jinkela_wire_9829),
        .dout(new_Jinkela_wire_9830)
    );

    bfr new_Jinkela_buffer_7925 (
        .din(new_Jinkela_wire_9792),
        .dout(new_Jinkela_wire_9793)
    );

    spl2 new_Jinkela_splitter_791 (
        .a(_0716_),
        .b(new_Jinkela_wire_10062),
        .c(new_Jinkela_wire_10063)
    );

    bfr new_Jinkela_buffer_7926 (
        .din(new_Jinkela_wire_9793),
        .dout(new_Jinkela_wire_9794)
    );

    bfr new_Jinkela_buffer_7959 (
        .din(new_Jinkela_wire_9830),
        .dout(new_Jinkela_wire_9831)
    );

    bfr new_Jinkela_buffer_7927 (
        .din(new_Jinkela_wire_9794),
        .dout(new_Jinkela_wire_9795)
    );

    bfr new_Jinkela_buffer_7995 (
        .din(new_Jinkela_wire_9874),
        .dout(new_Jinkela_wire_9875)
    );

    bfr new_Jinkela_buffer_7928 (
        .din(new_Jinkela_wire_9795),
        .dout(new_Jinkela_wire_9796)
    );

    bfr new_Jinkela_buffer_7960 (
        .din(new_Jinkela_wire_9831),
        .dout(new_Jinkela_wire_9832)
    );

    bfr new_Jinkela_buffer_7929 (
        .din(new_Jinkela_wire_9796),
        .dout(new_Jinkela_wire_9797)
    );

    bfr new_Jinkela_buffer_8168 (
        .din(new_Jinkela_wire_10049),
        .dout(new_Jinkela_wire_10050)
    );

    bfr new_Jinkela_buffer_8031 (
        .din(new_Jinkela_wire_9912),
        .dout(new_Jinkela_wire_9913)
    );

    bfr new_Jinkela_buffer_7930 (
        .din(new_Jinkela_wire_9797),
        .dout(new_Jinkela_wire_9798)
    );

    bfr new_Jinkela_buffer_7961 (
        .din(new_Jinkela_wire_9832),
        .dout(new_Jinkela_wire_9833)
    );

    bfr new_Jinkela_buffer_7931 (
        .din(new_Jinkela_wire_9798),
        .dout(new_Jinkela_wire_9799)
    );

    bfr new_Jinkela_buffer_7996 (
        .din(new_Jinkela_wire_9875),
        .dout(new_Jinkela_wire_9876)
    );

    bfr new_Jinkela_buffer_7932 (
        .din(new_Jinkela_wire_9799),
        .dout(new_Jinkela_wire_9800)
    );

    bfr new_Jinkela_buffer_7962 (
        .din(new_Jinkela_wire_9833),
        .dout(new_Jinkela_wire_9834)
    );

    bfr new_Jinkela_buffer_7933 (
        .din(new_Jinkela_wire_9800),
        .dout(new_Jinkela_wire_9801)
    );

    bfr new_Jinkela_buffer_7934 (
        .din(new_Jinkela_wire_9801),
        .dout(new_Jinkela_wire_9802)
    );

    bfr new_Jinkela_buffer_7963 (
        .din(new_Jinkela_wire_9834),
        .dout(new_Jinkela_wire_9835)
    );

    bfr new_Jinkela_buffer_7935 (
        .din(new_Jinkela_wire_9802),
        .dout(new_Jinkela_wire_9803)
    );

    bfr new_Jinkela_buffer_7997 (
        .din(new_Jinkela_wire_9876),
        .dout(new_Jinkela_wire_9877)
    );

    bfr new_Jinkela_buffer_7936 (
        .din(new_Jinkela_wire_9803),
        .dout(new_Jinkela_wire_9804)
    );

    bfr new_Jinkela_buffer_7964 (
        .din(new_Jinkela_wire_9835),
        .dout(new_Jinkela_wire_9836)
    );

    spl2 new_Jinkela_splitter_783 (
        .a(new_Jinkela_wire_9804),
        .b(new_Jinkela_wire_9805),
        .c(new_Jinkela_wire_9806)
    );

    bfr new_Jinkela_buffer_7965 (
        .din(new_Jinkela_wire_9836),
        .dout(new_Jinkela_wire_9837)
    );

    spl2 new_Jinkela_splitter_792 (
        .a(_0451_),
        .b(new_Jinkela_wire_10064),
        .c(new_Jinkela_wire_10065)
    );

    bfr new_Jinkela_buffer_8032 (
        .din(new_Jinkela_wire_9913),
        .dout(new_Jinkela_wire_9914)
    );

    bfr new_Jinkela_buffer_7998 (
        .din(new_Jinkela_wire_9877),
        .dout(new_Jinkela_wire_9878)
    );

    bfr new_Jinkela_buffer_7966 (
        .din(new_Jinkela_wire_9837),
        .dout(new_Jinkela_wire_9838)
    );

    bfr new_Jinkela_buffer_14970 (
        .din(_1371_),
        .dout(new_Jinkela_wire_17867)
    );

    spl2 new_Jinkela_splitter_1286 (
        .a(new_Jinkela_wire_17723),
        .b(new_Jinkela_wire_17724),
        .c(new_Jinkela_wire_17725)
    );

    bfr new_Jinkela_buffer_14917 (
        .din(new_Jinkela_wire_17803),
        .dout(new_Jinkela_wire_17804)
    );

    bfr new_Jinkela_buffer_14869 (
        .din(new_Jinkela_wire_17745),
        .dout(new_Jinkela_wire_17746)
    );

    bfr new_Jinkela_buffer_14870 (
        .din(new_Jinkela_wire_17746),
        .dout(new_Jinkela_wire_17747)
    );

    spl2 new_Jinkela_splitter_1296 (
        .a(_0054_),
        .b(new_Jinkela_wire_17865),
        .c(new_Jinkela_wire_17866)
    );

    bfr new_Jinkela_buffer_14871 (
        .din(new_Jinkela_wire_17747),
        .dout(new_Jinkela_wire_17748)
    );

    bfr new_Jinkela_buffer_14918 (
        .din(new_Jinkela_wire_17804),
        .dout(new_Jinkela_wire_17805)
    );

    bfr new_Jinkela_buffer_14872 (
        .din(new_Jinkela_wire_17748),
        .dout(new_Jinkela_wire_17749)
    );

    spl2 new_Jinkela_splitter_1299 (
        .a(_1251_),
        .b(new_Jinkela_wire_17975),
        .c(new_Jinkela_wire_17976)
    );

    bfr new_Jinkela_buffer_14873 (
        .din(new_Jinkela_wire_17749),
        .dout(new_Jinkela_wire_17750)
    );

    bfr new_Jinkela_buffer_14919 (
        .din(new_Jinkela_wire_17805),
        .dout(new_Jinkela_wire_17806)
    );

    bfr new_Jinkela_buffer_14874 (
        .din(new_Jinkela_wire_17750),
        .dout(new_Jinkela_wire_17751)
    );

    bfr new_Jinkela_buffer_15018 (
        .din(_1693_),
        .dout(new_Jinkela_wire_17917)
    );

    bfr new_Jinkela_buffer_14875 (
        .din(new_Jinkela_wire_17751),
        .dout(new_Jinkela_wire_17752)
    );

    bfr new_Jinkela_buffer_14920 (
        .din(new_Jinkela_wire_17806),
        .dout(new_Jinkela_wire_17807)
    );

    bfr new_Jinkela_buffer_14876 (
        .din(new_Jinkela_wire_17752),
        .dout(new_Jinkela_wire_17753)
    );

    bfr new_Jinkela_buffer_14971 (
        .din(new_Jinkela_wire_17867),
        .dout(new_Jinkela_wire_17868)
    );

    bfr new_Jinkela_buffer_14877 (
        .din(new_Jinkela_wire_17753),
        .dout(new_Jinkela_wire_17754)
    );

    bfr new_Jinkela_buffer_14921 (
        .din(new_Jinkela_wire_17807),
        .dout(new_Jinkela_wire_17808)
    );

    bfr new_Jinkela_buffer_14878 (
        .din(new_Jinkela_wire_17754),
        .dout(new_Jinkela_wire_17755)
    );

    spl2 new_Jinkela_splitter_1300 (
        .a(_1638_),
        .b(new_Jinkela_wire_17977),
        .c(new_Jinkela_wire_17978)
    );

    bfr new_Jinkela_buffer_14879 (
        .din(new_Jinkela_wire_17755),
        .dout(new_Jinkela_wire_17756)
    );

    bfr new_Jinkela_buffer_14922 (
        .din(new_Jinkela_wire_17808),
        .dout(new_Jinkela_wire_17809)
    );

    bfr new_Jinkela_buffer_14880 (
        .din(new_Jinkela_wire_17756),
        .dout(new_Jinkela_wire_17757)
    );

    bfr new_Jinkela_buffer_14972 (
        .din(new_Jinkela_wire_17868),
        .dout(new_Jinkela_wire_17869)
    );

    bfr new_Jinkela_buffer_14881 (
        .din(new_Jinkela_wire_17757),
        .dout(new_Jinkela_wire_17758)
    );

    bfr new_Jinkela_buffer_14923 (
        .din(new_Jinkela_wire_17809),
        .dout(new_Jinkela_wire_17810)
    );

    bfr new_Jinkela_buffer_14882 (
        .din(new_Jinkela_wire_17758),
        .dout(new_Jinkela_wire_17759)
    );

    bfr new_Jinkela_buffer_15019 (
        .din(new_Jinkela_wire_17917),
        .dout(new_Jinkela_wire_17918)
    );

    bfr new_Jinkela_buffer_14883 (
        .din(new_Jinkela_wire_17759),
        .dout(new_Jinkela_wire_17760)
    );

    bfr new_Jinkela_buffer_14924 (
        .din(new_Jinkela_wire_17810),
        .dout(new_Jinkela_wire_17811)
    );

    bfr new_Jinkela_buffer_14884 (
        .din(new_Jinkela_wire_17760),
        .dout(new_Jinkela_wire_17761)
    );

    bfr new_Jinkela_buffer_14973 (
        .din(new_Jinkela_wire_17869),
        .dout(new_Jinkela_wire_17870)
    );

    bfr new_Jinkela_buffer_14885 (
        .din(new_Jinkela_wire_17761),
        .dout(new_Jinkela_wire_17762)
    );

    bfr new_Jinkela_buffer_14925 (
        .din(new_Jinkela_wire_17811),
        .dout(new_Jinkela_wire_17812)
    );

    bfr new_Jinkela_buffer_14886 (
        .din(new_Jinkela_wire_17762),
        .dout(new_Jinkela_wire_17763)
    );

    spl2 new_Jinkela_splitter_1301 (
        .a(_1493_),
        .b(new_Jinkela_wire_17979),
        .c(new_Jinkela_wire_17980)
    );

    bfr new_Jinkela_buffer_14887 (
        .din(new_Jinkela_wire_17763),
        .dout(new_Jinkela_wire_17764)
    );

    bfr new_Jinkela_buffer_14926 (
        .din(new_Jinkela_wire_17812),
        .dout(new_Jinkela_wire_17813)
    );

    bfr new_Jinkela_buffer_14888 (
        .din(new_Jinkela_wire_17764),
        .dout(new_Jinkela_wire_17765)
    );

    bfr new_Jinkela_buffer_14974 (
        .din(new_Jinkela_wire_17870),
        .dout(new_Jinkela_wire_17871)
    );

    bfr new_Jinkela_buffer_4468 (
        .din(new_Jinkela_wire_5849),
        .dout(new_Jinkela_wire_5850)
    );

    bfr new_Jinkela_buffer_4513 (
        .din(new_Jinkela_wire_5902),
        .dout(new_Jinkela_wire_5903)
    );

    bfr new_Jinkela_buffer_4469 (
        .din(new_Jinkela_wire_5850),
        .dout(new_Jinkela_wire_5851)
    );

    bfr new_Jinkela_buffer_4583 (
        .din(new_Jinkela_wire_5976),
        .dout(new_Jinkela_wire_5977)
    );

    bfr new_Jinkela_buffer_4470 (
        .din(new_Jinkela_wire_5851),
        .dout(new_Jinkela_wire_5852)
    );

    bfr new_Jinkela_buffer_4514 (
        .din(new_Jinkela_wire_5903),
        .dout(new_Jinkela_wire_5904)
    );

    bfr new_Jinkela_buffer_4471 (
        .din(new_Jinkela_wire_5852),
        .dout(new_Jinkela_wire_5853)
    );

    spl2 new_Jinkela_splitter_552 (
        .a(_0173_),
        .b(new_Jinkela_wire_6001),
        .c(new_Jinkela_wire_6002)
    );

    bfr new_Jinkela_buffer_4472 (
        .din(new_Jinkela_wire_5853),
        .dout(new_Jinkela_wire_5854)
    );

    bfr new_Jinkela_buffer_4515 (
        .din(new_Jinkela_wire_5904),
        .dout(new_Jinkela_wire_5905)
    );

    bfr new_Jinkela_buffer_4473 (
        .din(new_Jinkela_wire_5854),
        .dout(new_Jinkela_wire_5855)
    );

    bfr new_Jinkela_buffer_4584 (
        .din(new_Jinkela_wire_5977),
        .dout(new_Jinkela_wire_5978)
    );

    bfr new_Jinkela_buffer_4474 (
        .din(new_Jinkela_wire_5855),
        .dout(new_Jinkela_wire_5856)
    );

    bfr new_Jinkela_buffer_4516 (
        .din(new_Jinkela_wire_5905),
        .dout(new_Jinkela_wire_5906)
    );

    bfr new_Jinkela_buffer_4475 (
        .din(new_Jinkela_wire_5856),
        .dout(new_Jinkela_wire_5857)
    );

    bfr new_Jinkela_buffer_4476 (
        .din(new_Jinkela_wire_5857),
        .dout(new_Jinkela_wire_5858)
    );

    bfr new_Jinkela_buffer_4517 (
        .din(new_Jinkela_wire_5906),
        .dout(new_Jinkela_wire_5907)
    );

    bfr new_Jinkela_buffer_4477 (
        .din(new_Jinkela_wire_5858),
        .dout(new_Jinkela_wire_5859)
    );

    bfr new_Jinkela_buffer_4585 (
        .din(new_Jinkela_wire_5978),
        .dout(new_Jinkela_wire_5979)
    );

    bfr new_Jinkela_buffer_4478 (
        .din(new_Jinkela_wire_5859),
        .dout(new_Jinkela_wire_5860)
    );

    bfr new_Jinkela_buffer_4518 (
        .din(new_Jinkela_wire_5907),
        .dout(new_Jinkela_wire_5908)
    );

    bfr new_Jinkela_buffer_4479 (
        .din(new_Jinkela_wire_5860),
        .dout(new_Jinkela_wire_5861)
    );

    spl2 new_Jinkela_splitter_553 (
        .a(_1047_),
        .b(new_Jinkela_wire_6007),
        .c(new_Jinkela_wire_6008)
    );

    bfr new_Jinkela_buffer_4480 (
        .din(new_Jinkela_wire_5861),
        .dout(new_Jinkela_wire_5862)
    );

    bfr new_Jinkela_buffer_4519 (
        .din(new_Jinkela_wire_5908),
        .dout(new_Jinkela_wire_5909)
    );

    bfr new_Jinkela_buffer_4481 (
        .din(new_Jinkela_wire_5862),
        .dout(new_Jinkela_wire_5863)
    );

    bfr new_Jinkela_buffer_4586 (
        .din(new_Jinkela_wire_5979),
        .dout(new_Jinkela_wire_5980)
    );

    bfr new_Jinkela_buffer_4482 (
        .din(new_Jinkela_wire_5863),
        .dout(new_Jinkela_wire_5864)
    );

    bfr new_Jinkela_buffer_4520 (
        .din(new_Jinkela_wire_5909),
        .dout(new_Jinkela_wire_5910)
    );

    bfr new_Jinkela_buffer_4483 (
        .din(new_Jinkela_wire_5864),
        .dout(new_Jinkela_wire_5865)
    );

    bfr new_Jinkela_buffer_4595 (
        .din(new_Jinkela_wire_6002),
        .dout(new_Jinkela_wire_6003)
    );

    bfr new_Jinkela_buffer_4599 (
        .din(_1588_),
        .dout(new_Jinkela_wire_6009)
    );

    bfr new_Jinkela_buffer_4484 (
        .din(new_Jinkela_wire_5865),
        .dout(new_Jinkela_wire_5866)
    );

    bfr new_Jinkela_buffer_4521 (
        .din(new_Jinkela_wire_5910),
        .dout(new_Jinkela_wire_5911)
    );

    bfr new_Jinkela_buffer_4485 (
        .din(new_Jinkela_wire_5866),
        .dout(new_Jinkela_wire_5867)
    );

    bfr new_Jinkela_buffer_4587 (
        .din(new_Jinkela_wire_5980),
        .dout(new_Jinkela_wire_5981)
    );

    bfr new_Jinkela_buffer_4486 (
        .din(new_Jinkela_wire_5867),
        .dout(new_Jinkela_wire_5868)
    );

    bfr new_Jinkela_buffer_4522 (
        .din(new_Jinkela_wire_5911),
        .dout(new_Jinkela_wire_5912)
    );

    bfr new_Jinkela_buffer_4487 (
        .din(new_Jinkela_wire_5868),
        .dout(new_Jinkela_wire_5869)
    );

    spl2 new_Jinkela_splitter_554 (
        .a(_1227_),
        .b(new_Jinkela_wire_6010),
        .c(new_Jinkela_wire_6011)
    );

    bfr new_Jinkela_buffer_4488 (
        .din(new_Jinkela_wire_5869),
        .dout(new_Jinkela_wire_5870)
    );

    bfr new_Jinkela_buffer_4523 (
        .din(new_Jinkela_wire_5912),
        .dout(new_Jinkela_wire_5913)
    );

    bfr new_Jinkela_buffer_11516 (
        .din(new_Jinkela_wire_13863),
        .dout(new_Jinkela_wire_13864)
    );

    bfr new_Jinkela_buffer_11423 (
        .din(new_Jinkela_wire_13766),
        .dout(new_Jinkela_wire_13767)
    );

    bfr new_Jinkela_buffer_11618 (
        .din(_0648_),
        .dout(new_Jinkela_wire_13980)
    );

    bfr new_Jinkela_buffer_11424 (
        .din(new_Jinkela_wire_13767),
        .dout(new_Jinkela_wire_13768)
    );

    bfr new_Jinkela_buffer_11517 (
        .din(new_Jinkela_wire_13864),
        .dout(new_Jinkela_wire_13865)
    );

    bfr new_Jinkela_buffer_11425 (
        .din(new_Jinkela_wire_13768),
        .dout(new_Jinkela_wire_13769)
    );

    bfr new_Jinkela_buffer_11613 (
        .din(new_Jinkela_wire_13974),
        .dout(new_Jinkela_wire_13975)
    );

    bfr new_Jinkela_buffer_11426 (
        .din(new_Jinkela_wire_13769),
        .dout(new_Jinkela_wire_13770)
    );

    bfr new_Jinkela_buffer_11518 (
        .din(new_Jinkela_wire_13865),
        .dout(new_Jinkela_wire_13866)
    );

    bfr new_Jinkela_buffer_11427 (
        .din(new_Jinkela_wire_13770),
        .dout(new_Jinkela_wire_13771)
    );

    bfr new_Jinkela_buffer_11619 (
        .din(new_Jinkela_wire_13980),
        .dout(new_Jinkela_wire_13981)
    );

    bfr new_Jinkela_buffer_11428 (
        .din(new_Jinkela_wire_13771),
        .dout(new_Jinkela_wire_13772)
    );

    bfr new_Jinkela_buffer_11519 (
        .din(new_Jinkela_wire_13866),
        .dout(new_Jinkela_wire_13867)
    );

    bfr new_Jinkela_buffer_11429 (
        .din(new_Jinkela_wire_13772),
        .dout(new_Jinkela_wire_13773)
    );

    bfr new_Jinkela_buffer_11614 (
        .din(new_Jinkela_wire_13975),
        .dout(new_Jinkela_wire_13976)
    );

    bfr new_Jinkela_buffer_11430 (
        .din(new_Jinkela_wire_13773),
        .dout(new_Jinkela_wire_13774)
    );

    bfr new_Jinkela_buffer_11520 (
        .din(new_Jinkela_wire_13867),
        .dout(new_Jinkela_wire_13868)
    );

    bfr new_Jinkela_buffer_11431 (
        .din(new_Jinkela_wire_13774),
        .dout(new_Jinkela_wire_13775)
    );

    bfr new_Jinkela_buffer_11620 (
        .din(new_Jinkela_wire_13985),
        .dout(new_Jinkela_wire_13986)
    );

    bfr new_Jinkela_buffer_11432 (
        .din(new_Jinkela_wire_13775),
        .dout(new_Jinkela_wire_13776)
    );

    bfr new_Jinkela_buffer_11521 (
        .din(new_Jinkela_wire_13868),
        .dout(new_Jinkela_wire_13869)
    );

    bfr new_Jinkela_buffer_11433 (
        .din(new_Jinkela_wire_13776),
        .dout(new_Jinkela_wire_13777)
    );

    bfr new_Jinkela_buffer_11615 (
        .din(new_Jinkela_wire_13976),
        .dout(new_Jinkela_wire_13977)
    );

    bfr new_Jinkela_buffer_11434 (
        .din(new_Jinkela_wire_13777),
        .dout(new_Jinkela_wire_13778)
    );

    bfr new_Jinkela_buffer_11522 (
        .din(new_Jinkela_wire_13869),
        .dout(new_Jinkela_wire_13870)
    );

    bfr new_Jinkela_buffer_11435 (
        .din(new_Jinkela_wire_13778),
        .dout(new_Jinkela_wire_13779)
    );

    bfr new_Jinkela_buffer_11436 (
        .din(new_Jinkela_wire_13779),
        .dout(new_Jinkela_wire_13780)
    );

    bfr new_Jinkela_buffer_11523 (
        .din(new_Jinkela_wire_13870),
        .dout(new_Jinkela_wire_13871)
    );

    bfr new_Jinkela_buffer_11437 (
        .din(new_Jinkela_wire_13780),
        .dout(new_Jinkela_wire_13781)
    );

    bfr new_Jinkela_buffer_11628 (
        .din(_0690_),
        .dout(new_Jinkela_wire_13996)
    );

    bfr new_Jinkela_buffer_11438 (
        .din(new_Jinkela_wire_13781),
        .dout(new_Jinkela_wire_13782)
    );

    bfr new_Jinkela_buffer_11524 (
        .din(new_Jinkela_wire_13871),
        .dout(new_Jinkela_wire_13872)
    );

    bfr new_Jinkela_buffer_11439 (
        .din(new_Jinkela_wire_13782),
        .dout(new_Jinkela_wire_13783)
    );

    spl2 new_Jinkela_splitter_1030 (
        .a(new_Jinkela_wire_13981),
        .b(new_Jinkela_wire_13982),
        .c(new_Jinkela_wire_13983)
    );

    bfr new_Jinkela_buffer_11440 (
        .din(new_Jinkela_wire_13783),
        .dout(new_Jinkela_wire_13784)
    );

    bfr new_Jinkela_buffer_11525 (
        .din(new_Jinkela_wire_13872),
        .dout(new_Jinkela_wire_13873)
    );

    bfr new_Jinkela_buffer_11441 (
        .din(new_Jinkela_wire_13784),
        .dout(new_Jinkela_wire_13785)
    );

    bfr new_Jinkela_buffer_11624 (
        .din(new_Jinkela_wire_13991),
        .dout(new_Jinkela_wire_13992)
    );

    bfr new_Jinkela_buffer_11442 (
        .din(new_Jinkela_wire_13785),
        .dout(new_Jinkela_wire_13786)
    );

    bfr new_Jinkela_buffer_11526 (
        .din(new_Jinkela_wire_13873),
        .dout(new_Jinkela_wire_13874)
    );

    bfr new_Jinkela_buffer_11617 (
        .din(_1040_),
        .dout(new_Jinkela_wire_13979)
    );

    bfr new_Jinkela_buffer_11443 (
        .din(new_Jinkela_wire_13786),
        .dout(new_Jinkela_wire_13787)
    );

    bfr new_Jinkela_buffer_7967 (
        .din(new_Jinkela_wire_9838),
        .dout(new_Jinkela_wire_9839)
    );

    bfr new_Jinkela_buffer_14889 (
        .din(new_Jinkela_wire_17765),
        .dout(new_Jinkela_wire_17766)
    );

    bfr new_Jinkela_buffer_7999 (
        .din(new_Jinkela_wire_9878),
        .dout(new_Jinkela_wire_9879)
    );

    bfr new_Jinkela_buffer_14927 (
        .din(new_Jinkela_wire_17813),
        .dout(new_Jinkela_wire_17814)
    );

    bfr new_Jinkela_buffer_7968 (
        .din(new_Jinkela_wire_9839),
        .dout(new_Jinkela_wire_9840)
    );

    bfr new_Jinkela_buffer_14890 (
        .din(new_Jinkela_wire_17766),
        .dout(new_Jinkela_wire_17767)
    );

    bfr new_Jinkela_buffer_8169 (
        .din(new_Jinkela_wire_10050),
        .dout(new_Jinkela_wire_10051)
    );

    bfr new_Jinkela_buffer_15020 (
        .din(new_Jinkela_wire_17918),
        .dout(new_Jinkela_wire_17919)
    );

    bfr new_Jinkela_buffer_8033 (
        .din(new_Jinkela_wire_9914),
        .dout(new_Jinkela_wire_9915)
    );

    bfr new_Jinkela_buffer_7969 (
        .din(new_Jinkela_wire_9840),
        .dout(new_Jinkela_wire_9841)
    );

    bfr new_Jinkela_buffer_14891 (
        .din(new_Jinkela_wire_17767),
        .dout(new_Jinkela_wire_17768)
    );

    bfr new_Jinkela_buffer_8000 (
        .din(new_Jinkela_wire_9879),
        .dout(new_Jinkela_wire_9880)
    );

    bfr new_Jinkela_buffer_14928 (
        .din(new_Jinkela_wire_17814),
        .dout(new_Jinkela_wire_17815)
    );

    bfr new_Jinkela_buffer_7970 (
        .din(new_Jinkela_wire_9841),
        .dout(new_Jinkela_wire_9842)
    );

    bfr new_Jinkela_buffer_14892 (
        .din(new_Jinkela_wire_17768),
        .dout(new_Jinkela_wire_17769)
    );

    bfr new_Jinkela_buffer_14975 (
        .din(new_Jinkela_wire_17871),
        .dout(new_Jinkela_wire_17872)
    );

    bfr new_Jinkela_buffer_7971 (
        .din(new_Jinkela_wire_9842),
        .dout(new_Jinkela_wire_9843)
    );

    bfr new_Jinkela_buffer_14893 (
        .din(new_Jinkela_wire_17769),
        .dout(new_Jinkela_wire_17770)
    );

    bfr new_Jinkela_buffer_8001 (
        .din(new_Jinkela_wire_9880),
        .dout(new_Jinkela_wire_9881)
    );

    bfr new_Jinkela_buffer_14929 (
        .din(new_Jinkela_wire_17815),
        .dout(new_Jinkela_wire_17816)
    );

    bfr new_Jinkela_buffer_7972 (
        .din(new_Jinkela_wire_9843),
        .dout(new_Jinkela_wire_9844)
    );

    bfr new_Jinkela_buffer_14894 (
        .din(new_Jinkela_wire_17770),
        .dout(new_Jinkela_wire_17771)
    );

    spl2 new_Jinkela_splitter_794 (
        .a(_0895_),
        .b(new_Jinkela_wire_10073),
        .c(new_Jinkela_wire_10074)
    );

    bfr new_Jinkela_buffer_8034 (
        .din(new_Jinkela_wire_9915),
        .dout(new_Jinkela_wire_9916)
    );

    bfr new_Jinkela_buffer_7973 (
        .din(new_Jinkela_wire_9844),
        .dout(new_Jinkela_wire_9845)
    );

    bfr new_Jinkela_buffer_14895 (
        .din(new_Jinkela_wire_17771),
        .dout(new_Jinkela_wire_17772)
    );

    bfr new_Jinkela_buffer_8002 (
        .din(new_Jinkela_wire_9881),
        .dout(new_Jinkela_wire_9882)
    );

    bfr new_Jinkela_buffer_14930 (
        .din(new_Jinkela_wire_17816),
        .dout(new_Jinkela_wire_17817)
    );

    bfr new_Jinkela_buffer_7974 (
        .din(new_Jinkela_wire_9845),
        .dout(new_Jinkela_wire_9846)
    );

    bfr new_Jinkela_buffer_14896 (
        .din(new_Jinkela_wire_17772),
        .dout(new_Jinkela_wire_17773)
    );

    bfr new_Jinkela_buffer_14976 (
        .din(new_Jinkela_wire_17872),
        .dout(new_Jinkela_wire_17873)
    );

    bfr new_Jinkela_buffer_7975 (
        .din(new_Jinkela_wire_9846),
        .dout(new_Jinkela_wire_9847)
    );

    bfr new_Jinkela_buffer_14897 (
        .din(new_Jinkela_wire_17773),
        .dout(new_Jinkela_wire_17774)
    );

    bfr new_Jinkela_buffer_8003 (
        .din(new_Jinkela_wire_9882),
        .dout(new_Jinkela_wire_9883)
    );

    bfr new_Jinkela_buffer_14931 (
        .din(new_Jinkela_wire_17817),
        .dout(new_Jinkela_wire_17818)
    );

    bfr new_Jinkela_buffer_7976 (
        .din(new_Jinkela_wire_9847),
        .dout(new_Jinkela_wire_9848)
    );

    bfr new_Jinkela_buffer_14898 (
        .din(new_Jinkela_wire_17774),
        .dout(new_Jinkela_wire_17775)
    );

    bfr new_Jinkela_buffer_8170 (
        .din(new_Jinkela_wire_10051),
        .dout(new_Jinkela_wire_10052)
    );

    bfr new_Jinkela_buffer_15021 (
        .din(new_Jinkela_wire_17919),
        .dout(new_Jinkela_wire_17920)
    );

    bfr new_Jinkela_buffer_8035 (
        .din(new_Jinkela_wire_9916),
        .dout(new_Jinkela_wire_9917)
    );

    bfr new_Jinkela_buffer_7977 (
        .din(new_Jinkela_wire_9848),
        .dout(new_Jinkela_wire_9849)
    );

    bfr new_Jinkela_buffer_14899 (
        .din(new_Jinkela_wire_17775),
        .dout(new_Jinkela_wire_17776)
    );

    bfr new_Jinkela_buffer_8004 (
        .din(new_Jinkela_wire_9883),
        .dout(new_Jinkela_wire_9884)
    );

    bfr new_Jinkela_buffer_14932 (
        .din(new_Jinkela_wire_17818),
        .dout(new_Jinkela_wire_17819)
    );

    bfr new_Jinkela_buffer_7978 (
        .din(new_Jinkela_wire_9849),
        .dout(new_Jinkela_wire_9850)
    );

    bfr new_Jinkela_buffer_14900 (
        .din(new_Jinkela_wire_17776),
        .dout(new_Jinkela_wire_17777)
    );

    bfr new_Jinkela_buffer_14977 (
        .din(new_Jinkela_wire_17873),
        .dout(new_Jinkela_wire_17874)
    );

    bfr new_Jinkela_buffer_7979 (
        .din(new_Jinkela_wire_9850),
        .dout(new_Jinkela_wire_9851)
    );

    bfr new_Jinkela_buffer_14901 (
        .din(new_Jinkela_wire_17777),
        .dout(new_Jinkela_wire_17778)
    );

    bfr new_Jinkela_buffer_8005 (
        .din(new_Jinkela_wire_9884),
        .dout(new_Jinkela_wire_9885)
    );

    bfr new_Jinkela_buffer_14933 (
        .din(new_Jinkela_wire_17819),
        .dout(new_Jinkela_wire_17820)
    );

    bfr new_Jinkela_buffer_7980 (
        .din(new_Jinkela_wire_9851),
        .dout(new_Jinkela_wire_9852)
    );

    bfr new_Jinkela_buffer_14902 (
        .din(new_Jinkela_wire_17778),
        .dout(new_Jinkela_wire_17779)
    );

    bfr new_Jinkela_buffer_8036 (
        .din(new_Jinkela_wire_9917),
        .dout(new_Jinkela_wire_9918)
    );

    spl2 new_Jinkela_splitter_1302 (
        .a(_1218_),
        .b(new_Jinkela_wire_17981),
        .c(new_Jinkela_wire_17982)
    );

    bfr new_Jinkela_buffer_7981 (
        .din(new_Jinkela_wire_9852),
        .dout(new_Jinkela_wire_9853)
    );

    bfr new_Jinkela_buffer_14903 (
        .din(new_Jinkela_wire_17779),
        .dout(new_Jinkela_wire_17780)
    );

    bfr new_Jinkela_buffer_8006 (
        .din(new_Jinkela_wire_9885),
        .dout(new_Jinkela_wire_9886)
    );

    bfr new_Jinkela_buffer_14934 (
        .din(new_Jinkela_wire_17820),
        .dout(new_Jinkela_wire_17821)
    );

    bfr new_Jinkela_buffer_7982 (
        .din(new_Jinkela_wire_9853),
        .dout(new_Jinkela_wire_9854)
    );

    bfr new_Jinkela_buffer_14904 (
        .din(new_Jinkela_wire_17780),
        .dout(new_Jinkela_wire_17781)
    );

    bfr new_Jinkela_buffer_14978 (
        .din(new_Jinkela_wire_17874),
        .dout(new_Jinkela_wire_17875)
    );

    bfr new_Jinkela_buffer_8178 (
        .din(_1348_),
        .dout(new_Jinkela_wire_10066)
    );

    bfr new_Jinkela_buffer_7983 (
        .din(new_Jinkela_wire_9854),
        .dout(new_Jinkela_wire_9855)
    );

    spl2 new_Jinkela_splitter_1287 (
        .a(new_Jinkela_wire_17781),
        .b(new_Jinkela_wire_17782),
        .c(new_Jinkela_wire_17783)
    );

    bfr new_Jinkela_buffer_8007 (
        .din(new_Jinkela_wire_9886),
        .dout(new_Jinkela_wire_9887)
    );

    bfr new_Jinkela_buffer_15022 (
        .din(new_Jinkela_wire_17920),
        .dout(new_Jinkela_wire_17921)
    );

    bfr new_Jinkela_buffer_7984 (
        .din(new_Jinkela_wire_9855),
        .dout(new_Jinkela_wire_9856)
    );

    bfr new_Jinkela_buffer_14935 (
        .din(new_Jinkela_wire_17821),
        .dout(new_Jinkela_wire_17822)
    );

    bfr new_Jinkela_buffer_8171 (
        .din(new_Jinkela_wire_10052),
        .dout(new_Jinkela_wire_10053)
    );

    bfr new_Jinkela_buffer_14936 (
        .din(new_Jinkela_wire_17822),
        .dout(new_Jinkela_wire_17823)
    );

    bfr new_Jinkela_buffer_8037 (
        .din(new_Jinkela_wire_9918),
        .dout(new_Jinkela_wire_9919)
    );

    spl2 new_Jinkela_splitter_785 (
        .a(new_Jinkela_wire_9856),
        .b(new_Jinkela_wire_9857),
        .c(new_Jinkela_wire_9858)
    );

    bfr new_Jinkela_buffer_14979 (
        .din(new_Jinkela_wire_17875),
        .dout(new_Jinkela_wire_17876)
    );

    bfr new_Jinkela_buffer_14937 (
        .din(new_Jinkela_wire_17823),
        .dout(new_Jinkela_wire_17824)
    );

    bfr new_Jinkela_buffer_8008 (
        .din(new_Jinkela_wire_9887),
        .dout(new_Jinkela_wire_9888)
    );

    spl2 new_Jinkela_splitter_1304 (
        .a(_0053_),
        .b(new_Jinkela_wire_17985),
        .c(new_Jinkela_wire_17986)
    );

    spl2 new_Jinkela_splitter_1303 (
        .a(_0301_),
        .b(new_Jinkela_wire_17983),
        .c(new_Jinkela_wire_17984)
    );

    bfr new_Jinkela_buffer_8009 (
        .din(new_Jinkela_wire_9888),
        .dout(new_Jinkela_wire_9889)
    );

    bfr new_Jinkela_buffer_14938 (
        .din(new_Jinkela_wire_17824),
        .dout(new_Jinkela_wire_17825)
    );

    spl2 new_Jinkela_splitter_793 (
        .a(_1763_),
        .b(new_Jinkela_wire_10067),
        .c(new_Jinkela_wire_10068)
    );

    bfr new_Jinkela_buffer_14980 (
        .din(new_Jinkela_wire_17876),
        .dout(new_Jinkela_wire_17877)
    );

    bfr new_Jinkela_buffer_8038 (
        .din(new_Jinkela_wire_9919),
        .dout(new_Jinkela_wire_9920)
    );

    bfr new_Jinkela_buffer_8010 (
        .din(new_Jinkela_wire_9889),
        .dout(new_Jinkela_wire_9890)
    );

    bfr new_Jinkela_buffer_14939 (
        .din(new_Jinkela_wire_17825),
        .dout(new_Jinkela_wire_17826)
    );

    bfr new_Jinkela_buffer_4489 (
        .din(new_Jinkela_wire_5870),
        .dout(new_Jinkela_wire_5871)
    );

    bfr new_Jinkela_buffer_4588 (
        .din(new_Jinkela_wire_5981),
        .dout(new_Jinkela_wire_5982)
    );

    bfr new_Jinkela_buffer_4490 (
        .din(new_Jinkela_wire_5871),
        .dout(new_Jinkela_wire_5872)
    );

    bfr new_Jinkela_buffer_4524 (
        .din(new_Jinkela_wire_5913),
        .dout(new_Jinkela_wire_5914)
    );

    bfr new_Jinkela_buffer_4491 (
        .din(new_Jinkela_wire_5872),
        .dout(new_Jinkela_wire_5873)
    );

    bfr new_Jinkela_buffer_4596 (
        .din(new_Jinkela_wire_6003),
        .dout(new_Jinkela_wire_6004)
    );

    bfr new_Jinkela_buffer_4492 (
        .din(new_Jinkela_wire_5873),
        .dout(new_Jinkela_wire_5874)
    );

    bfr new_Jinkela_buffer_4525 (
        .din(new_Jinkela_wire_5914),
        .dout(new_Jinkela_wire_5915)
    );

    bfr new_Jinkela_buffer_4493 (
        .din(new_Jinkela_wire_5874),
        .dout(new_Jinkela_wire_5875)
    );

    bfr new_Jinkela_buffer_4589 (
        .din(new_Jinkela_wire_5982),
        .dout(new_Jinkela_wire_5983)
    );

    bfr new_Jinkela_buffer_4494 (
        .din(new_Jinkela_wire_5875),
        .dout(new_Jinkela_wire_5876)
    );

    bfr new_Jinkela_buffer_4526 (
        .din(new_Jinkela_wire_5915),
        .dout(new_Jinkela_wire_5916)
    );

    bfr new_Jinkela_buffer_4495 (
        .din(new_Jinkela_wire_5876),
        .dout(new_Jinkela_wire_5877)
    );

    bfr new_Jinkela_buffer_4600 (
        .din(_1687_),
        .dout(new_Jinkela_wire_6012)
    );

    spl2 new_Jinkela_splitter_540 (
        .a(new_Jinkela_wire_5877),
        .b(new_Jinkela_wire_5878),
        .c(new_Jinkela_wire_5879)
    );

    bfr new_Jinkela_buffer_4590 (
        .din(new_Jinkela_wire_5983),
        .dout(new_Jinkela_wire_5984)
    );

    bfr new_Jinkela_buffer_4527 (
        .din(new_Jinkela_wire_5916),
        .dout(new_Jinkela_wire_5917)
    );

    bfr new_Jinkela_buffer_4528 (
        .din(new_Jinkela_wire_5917),
        .dout(new_Jinkela_wire_5918)
    );

    bfr new_Jinkela_buffer_4597 (
        .din(new_Jinkela_wire_6004),
        .dout(new_Jinkela_wire_6005)
    );

    bfr new_Jinkela_buffer_4529 (
        .din(new_Jinkela_wire_5918),
        .dout(new_Jinkela_wire_5919)
    );

    bfr new_Jinkela_buffer_4591 (
        .din(new_Jinkela_wire_5984),
        .dout(new_Jinkela_wire_5985)
    );

    bfr new_Jinkela_buffer_4530 (
        .din(new_Jinkela_wire_5919),
        .dout(new_Jinkela_wire_5920)
    );

    bfr new_Jinkela_buffer_4777 (
        .din(_1164_),
        .dout(new_Jinkela_wire_6193)
    );

    bfr new_Jinkela_buffer_4531 (
        .din(new_Jinkela_wire_5920),
        .dout(new_Jinkela_wire_5921)
    );

    spl2 new_Jinkela_splitter_546 (
        .a(new_Jinkela_wire_5985),
        .b(new_Jinkela_wire_5986),
        .c(new_Jinkela_wire_5987)
    );

    bfr new_Jinkela_buffer_4532 (
        .din(new_Jinkela_wire_5921),
        .dout(new_Jinkela_wire_5922)
    );

    bfr new_Jinkela_buffer_4681 (
        .din(_0216_),
        .dout(new_Jinkela_wire_6095)
    );

    bfr new_Jinkela_buffer_4533 (
        .din(new_Jinkela_wire_5922),
        .dout(new_Jinkela_wire_5923)
    );

    bfr new_Jinkela_buffer_4598 (
        .din(new_Jinkela_wire_6005),
        .dout(new_Jinkela_wire_6006)
    );

    bfr new_Jinkela_buffer_4534 (
        .din(new_Jinkela_wire_5923),
        .dout(new_Jinkela_wire_5924)
    );

    bfr new_Jinkela_buffer_4601 (
        .din(new_Jinkela_wire_6012),
        .dout(new_Jinkela_wire_6013)
    );

    bfr new_Jinkela_buffer_4535 (
        .din(new_Jinkela_wire_5924),
        .dout(new_Jinkela_wire_5925)
    );

    spl2 new_Jinkela_splitter_557 (
        .a(_1283_),
        .b(new_Jinkela_wire_6194),
        .c(new_Jinkela_wire_6195)
    );

    bfr new_Jinkela_buffer_4536 (
        .din(new_Jinkela_wire_5925),
        .dout(new_Jinkela_wire_5926)
    );

    bfr new_Jinkela_buffer_4602 (
        .din(new_Jinkela_wire_6013),
        .dout(new_Jinkela_wire_6014)
    );

    bfr new_Jinkela_buffer_4537 (
        .din(new_Jinkela_wire_5926),
        .dout(new_Jinkela_wire_5927)
    );

    bfr new_Jinkela_buffer_4682 (
        .din(new_Jinkela_wire_6095),
        .dout(new_Jinkela_wire_6096)
    );

    bfr new_Jinkela_buffer_4538 (
        .din(new_Jinkela_wire_5927),
        .dout(new_Jinkela_wire_5928)
    );

    bfr new_Jinkela_buffer_4603 (
        .din(new_Jinkela_wire_6014),
        .dout(new_Jinkela_wire_6015)
    );

    bfr new_Jinkela_buffer_4539 (
        .din(new_Jinkela_wire_5928),
        .dout(new_Jinkela_wire_5929)
    );

    spl2 new_Jinkela_splitter_558 (
        .a(_1423_),
        .b(new_Jinkela_wire_6196),
        .c(new_Jinkela_wire_6197)
    );

    bfr new_Jinkela_buffer_4540 (
        .din(new_Jinkela_wire_5929),
        .dout(new_Jinkela_wire_5930)
    );

    bfr new_Jinkela_buffer_11527 (
        .din(new_Jinkela_wire_13874),
        .dout(new_Jinkela_wire_13875)
    );

    bfr new_Jinkela_buffer_11444 (
        .din(new_Jinkela_wire_13787),
        .dout(new_Jinkela_wire_13788)
    );

    bfr new_Jinkela_buffer_11621 (
        .din(new_Jinkela_wire_13986),
        .dout(new_Jinkela_wire_13987)
    );

    bfr new_Jinkela_buffer_11445 (
        .din(new_Jinkela_wire_13788),
        .dout(new_Jinkela_wire_13789)
    );

    bfr new_Jinkela_buffer_11528 (
        .din(new_Jinkela_wire_13875),
        .dout(new_Jinkela_wire_13876)
    );

    bfr new_Jinkela_buffer_11446 (
        .din(new_Jinkela_wire_13789),
        .dout(new_Jinkela_wire_13790)
    );

    spl2 new_Jinkela_splitter_1033 (
        .a(_1004_),
        .b(new_Jinkela_wire_13997),
        .c(new_Jinkela_wire_13998)
    );

    bfr new_Jinkela_buffer_11447 (
        .din(new_Jinkela_wire_13790),
        .dout(new_Jinkela_wire_13791)
    );

    bfr new_Jinkela_buffer_11529 (
        .din(new_Jinkela_wire_13876),
        .dout(new_Jinkela_wire_13877)
    );

    bfr new_Jinkela_buffer_11448 (
        .din(new_Jinkela_wire_13791),
        .dout(new_Jinkela_wire_13792)
    );

    bfr new_Jinkela_buffer_11622 (
        .din(new_Jinkela_wire_13987),
        .dout(new_Jinkela_wire_13988)
    );

    bfr new_Jinkela_buffer_11449 (
        .din(new_Jinkela_wire_13792),
        .dout(new_Jinkela_wire_13793)
    );

    bfr new_Jinkela_buffer_11530 (
        .din(new_Jinkela_wire_13877),
        .dout(new_Jinkela_wire_13878)
    );

    bfr new_Jinkela_buffer_11450 (
        .din(new_Jinkela_wire_13793),
        .dout(new_Jinkela_wire_13794)
    );

    bfr new_Jinkela_buffer_11629 (
        .din(_1611_),
        .dout(new_Jinkela_wire_13999)
    );

    bfr new_Jinkela_buffer_11634 (
        .din(_0676_),
        .dout(new_Jinkela_wire_14006)
    );

    bfr new_Jinkela_buffer_11451 (
        .din(new_Jinkela_wire_13794),
        .dout(new_Jinkela_wire_13795)
    );

    bfr new_Jinkela_buffer_11531 (
        .din(new_Jinkela_wire_13878),
        .dout(new_Jinkela_wire_13879)
    );

    bfr new_Jinkela_buffer_11452 (
        .din(new_Jinkela_wire_13795),
        .dout(new_Jinkela_wire_13796)
    );

    bfr new_Jinkela_buffer_11623 (
        .din(new_Jinkela_wire_13988),
        .dout(new_Jinkela_wire_13989)
    );

    bfr new_Jinkela_buffer_11453 (
        .din(new_Jinkela_wire_13796),
        .dout(new_Jinkela_wire_13797)
    );

    bfr new_Jinkela_buffer_11532 (
        .din(new_Jinkela_wire_13879),
        .dout(new_Jinkela_wire_13880)
    );

    bfr new_Jinkela_buffer_11454 (
        .din(new_Jinkela_wire_13797),
        .dout(new_Jinkela_wire_13798)
    );

    bfr new_Jinkela_buffer_11625 (
        .din(new_Jinkela_wire_13992),
        .dout(new_Jinkela_wire_13993)
    );

    bfr new_Jinkela_buffer_11455 (
        .din(new_Jinkela_wire_13798),
        .dout(new_Jinkela_wire_13799)
    );

    bfr new_Jinkela_buffer_11533 (
        .din(new_Jinkela_wire_13880),
        .dout(new_Jinkela_wire_13881)
    );

    bfr new_Jinkela_buffer_11456 (
        .din(new_Jinkela_wire_13799),
        .dout(new_Jinkela_wire_13800)
    );

    bfr new_Jinkela_buffer_11457 (
        .din(new_Jinkela_wire_13800),
        .dout(new_Jinkela_wire_13801)
    );

    bfr new_Jinkela_buffer_11534 (
        .din(new_Jinkela_wire_13881),
        .dout(new_Jinkela_wire_13882)
    );

    bfr new_Jinkela_buffer_11458 (
        .din(new_Jinkela_wire_13801),
        .dout(new_Jinkela_wire_13802)
    );

    bfr new_Jinkela_buffer_11626 (
        .din(new_Jinkela_wire_13993),
        .dout(new_Jinkela_wire_13994)
    );

    bfr new_Jinkela_buffer_11459 (
        .din(new_Jinkela_wire_13802),
        .dout(new_Jinkela_wire_13803)
    );

    bfr new_Jinkela_buffer_11535 (
        .din(new_Jinkela_wire_13882),
        .dout(new_Jinkela_wire_13883)
    );

    bfr new_Jinkela_buffer_11460 (
        .din(new_Jinkela_wire_13803),
        .dout(new_Jinkela_wire_13804)
    );

    bfr new_Jinkela_buffer_11630 (
        .din(_0996_),
        .dout(new_Jinkela_wire_14000)
    );

    bfr new_Jinkela_buffer_11461 (
        .din(new_Jinkela_wire_13804),
        .dout(new_Jinkela_wire_13805)
    );

    bfr new_Jinkela_buffer_11536 (
        .din(new_Jinkela_wire_13883),
        .dout(new_Jinkela_wire_13884)
    );

    bfr new_Jinkela_buffer_11462 (
        .din(new_Jinkela_wire_13805),
        .dout(new_Jinkela_wire_13806)
    );

    bfr new_Jinkela_buffer_11627 (
        .din(new_Jinkela_wire_13994),
        .dout(new_Jinkela_wire_13995)
    );

    bfr new_Jinkela_buffer_11463 (
        .din(new_Jinkela_wire_13806),
        .dout(new_Jinkela_wire_13807)
    );

    bfr new_Jinkela_buffer_11537 (
        .din(new_Jinkela_wire_13884),
        .dout(new_Jinkela_wire_13885)
    );

    bfr new_Jinkela_buffer_11464 (
        .din(new_Jinkela_wire_13807),
        .dout(new_Jinkela_wire_13808)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1718),
        .dout(new_Jinkela_wire_1719)
    );

    bfr new_Jinkela_buffer_8011 (
        .din(new_Jinkela_wire_9890),
        .dout(new_Jinkela_wire_9891)
    );

    bfr new_Jinkela_buffer_8172 (
        .din(new_Jinkela_wire_10053),
        .dout(new_Jinkela_wire_10054)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1719),
        .dout(new_Jinkela_wire_1720)
    );

    bfr new_Jinkela_buffer_8039 (
        .din(new_Jinkela_wire_9920),
        .dout(new_Jinkela_wire_9921)
    );

    bfr new_Jinkela_buffer_8012 (
        .din(new_Jinkela_wire_9891),
        .dout(new_Jinkela_wire_9892)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1817),
        .dout(new_Jinkela_wire_1818)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1720),
        .dout(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_8013 (
        .din(new_Jinkela_wire_9892),
        .dout(new_Jinkela_wire_9893)
    );

    bfr new_Jinkela_buffer_8179 (
        .din(new_Jinkela_wire_10068),
        .dout(new_Jinkela_wire_10069)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1721),
        .dout(new_Jinkela_wire_1722)
    );

    bfr new_Jinkela_buffer_8040 (
        .din(new_Jinkela_wire_9921),
        .dout(new_Jinkela_wire_9922)
    );

    bfr new_Jinkela_buffer_8014 (
        .din(new_Jinkela_wire_9893),
        .dout(new_Jinkela_wire_9894)
    );

    spl2 new_Jinkela_splitter_259 (
        .a(_1668_),
        .b(new_Jinkela_wire_1912),
        .c(new_Jinkela_wire_1913)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(new_Jinkela_wire_1818),
        .dout(new_Jinkela_wire_1819)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1722),
        .dout(new_Jinkela_wire_1723)
    );

    bfr new_Jinkela_buffer_8015 (
        .din(new_Jinkela_wire_9894),
        .dout(new_Jinkela_wire_9895)
    );

    bfr new_Jinkela_buffer_8173 (
        .din(new_Jinkela_wire_10054),
        .dout(new_Jinkela_wire_10055)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1723),
        .dout(new_Jinkela_wire_1724)
    );

    bfr new_Jinkela_buffer_8041 (
        .din(new_Jinkela_wire_9922),
        .dout(new_Jinkela_wire_9923)
    );

    bfr new_Jinkela_buffer_8016 (
        .din(new_Jinkela_wire_9895),
        .dout(new_Jinkela_wire_9896)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1819),
        .dout(new_Jinkela_wire_1820)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1724),
        .dout(new_Jinkela_wire_1725)
    );

    bfr new_Jinkela_buffer_8017 (
        .din(new_Jinkela_wire_9896),
        .dout(new_Jinkela_wire_9897)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1725),
        .dout(new_Jinkela_wire_1726)
    );

    bfr new_Jinkela_buffer_8042 (
        .din(new_Jinkela_wire_9923),
        .dout(new_Jinkela_wire_9924)
    );

    bfr new_Jinkela_buffer_8018 (
        .din(new_Jinkela_wire_9897),
        .dout(new_Jinkela_wire_9898)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(new_Jinkela_wire_1907),
        .dout(new_Jinkela_wire_1908)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(new_Jinkela_wire_1820),
        .dout(new_Jinkela_wire_1821)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1726),
        .dout(new_Jinkela_wire_1727)
    );

    bfr new_Jinkela_buffer_8183 (
        .din(_0812_),
        .dout(new_Jinkela_wire_10075)
    );

    bfr new_Jinkela_buffer_8019 (
        .din(new_Jinkela_wire_9898),
        .dout(new_Jinkela_wire_9899)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(_0795_),
        .dout(new_Jinkela_wire_1914)
    );

    bfr new_Jinkela_buffer_8174 (
        .din(new_Jinkela_wire_10055),
        .dout(new_Jinkela_wire_10056)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1727),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_8043 (
        .din(new_Jinkela_wire_9924),
        .dout(new_Jinkela_wire_9925)
    );

    bfr new_Jinkela_buffer_8020 (
        .din(new_Jinkela_wire_9899),
        .dout(new_Jinkela_wire_9900)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1728),
        .dout(new_Jinkela_wire_1729)
    );

    bfr new_Jinkela_buffer_8021 (
        .din(new_Jinkela_wire_9900),
        .dout(new_Jinkela_wire_9901)
    );

    spl2 new_Jinkela_splitter_797 (
        .a(_1618_),
        .b(new_Jinkela_wire_10081),
        .c(new_Jinkela_wire_10082)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1729),
        .dout(new_Jinkela_wire_1730)
    );

    bfr new_Jinkela_buffer_8044 (
        .din(new_Jinkela_wire_9925),
        .dout(new_Jinkela_wire_9926)
    );

    bfr new_Jinkela_buffer_8022 (
        .din(new_Jinkela_wire_9901),
        .dout(new_Jinkela_wire_9902)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1822),
        .dout(new_Jinkela_wire_1823)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1730),
        .dout(new_Jinkela_wire_1731)
    );

    bfr new_Jinkela_buffer_8023 (
        .din(new_Jinkela_wire_9902),
        .dout(new_Jinkela_wire_9903)
    );

    bfr new_Jinkela_buffer_8175 (
        .din(new_Jinkela_wire_10056),
        .dout(new_Jinkela_wire_10057)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1731),
        .dout(new_Jinkela_wire_1732)
    );

    bfr new_Jinkela_buffer_8045 (
        .din(new_Jinkela_wire_9926),
        .dout(new_Jinkela_wire_9927)
    );

    bfr new_Jinkela_buffer_8024 (
        .din(new_Jinkela_wire_9903),
        .dout(new_Jinkela_wire_9904)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(new_Jinkela_wire_1908),
        .dout(new_Jinkela_wire_1909)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1823),
        .dout(new_Jinkela_wire_1824)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_Jinkela_wire_1732),
        .dout(new_Jinkela_wire_1733)
    );

    bfr new_Jinkela_buffer_8025 (
        .din(new_Jinkela_wire_9904),
        .dout(new_Jinkela_wire_9905)
    );

    bfr new_Jinkela_buffer_8180 (
        .din(new_Jinkela_wire_10069),
        .dout(new_Jinkela_wire_10070)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1733),
        .dout(new_Jinkela_wire_1734)
    );

    bfr new_Jinkela_buffer_8046 (
        .din(new_Jinkela_wire_9927),
        .dout(new_Jinkela_wire_9928)
    );

    spl2 new_Jinkela_splitter_789 (
        .a(new_Jinkela_wire_9905),
        .b(new_Jinkela_wire_9906),
        .c(new_Jinkela_wire_9907)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(_0525_),
        .b(new_Jinkela_wire_2013),
        .c(new_Jinkela_wire_2014)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1824),
        .dout(new_Jinkela_wire_1825)
    );

    spl2 new_Jinkela_splitter_790 (
        .a(new_Jinkela_wire_10057),
        .b(new_Jinkela_wire_10058),
        .c(new_Jinkela_wire_10059)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1734),
        .dout(new_Jinkela_wire_1735)
    );

    bfr new_Jinkela_buffer_8047 (
        .din(new_Jinkela_wire_9928),
        .dout(new_Jinkela_wire_9929)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(_0771_),
        .dout(new_Jinkela_wire_1915)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1735),
        .dout(new_Jinkela_wire_1736)
    );

    bfr new_Jinkela_buffer_8181 (
        .din(new_Jinkela_wire_10070),
        .dout(new_Jinkela_wire_10071)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_1909),
        .dout(new_Jinkela_wire_1910)
    );

    bfr new_Jinkela_buffer_8048 (
        .din(new_Jinkela_wire_9929),
        .dout(new_Jinkela_wire_9930)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1736),
        .dout(new_Jinkela_wire_1737)
    );

    spl2 new_Jinkela_splitter_796 (
        .a(_0524_),
        .b(new_Jinkela_wire_10079),
        .c(new_Jinkela_wire_10080)
    );

    bfr new_Jinkela_buffer_8049 (
        .din(new_Jinkela_wire_9930),
        .dout(new_Jinkela_wire_9931)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1737),
        .dout(new_Jinkela_wire_1738)
    );

    bfr new_Jinkela_buffer_8184 (
        .din(_0066_),
        .dout(new_Jinkela_wire_10076)
    );

    bfr new_Jinkela_buffer_8050 (
        .din(new_Jinkela_wire_9931),
        .dout(new_Jinkela_wire_9932)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1826),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1738),
        .dout(new_Jinkela_wire_1739)
    );

    bfr new_Jinkela_buffer_8182 (
        .din(new_Jinkela_wire_10071),
        .dout(new_Jinkela_wire_10072)
    );

    bfr new_Jinkela_buffer_8051 (
        .din(new_Jinkela_wire_9932),
        .dout(new_Jinkela_wire_9933)
    );

    bfr new_Jinkela_buffer_4604 (
        .din(new_Jinkela_wire_6015),
        .dout(new_Jinkela_wire_6016)
    );

    spl2 new_Jinkela_splitter_1035 (
        .a(_0628_),
        .b(new_Jinkela_wire_14007),
        .c(new_Jinkela_wire_14008)
    );

    bfr new_Jinkela_buffer_4541 (
        .din(new_Jinkela_wire_5930),
        .dout(new_Jinkela_wire_5931)
    );

    bfr new_Jinkela_buffer_11465 (
        .din(new_Jinkela_wire_13808),
        .dout(new_Jinkela_wire_13809)
    );

    bfr new_Jinkela_buffer_4683 (
        .din(new_Jinkela_wire_6096),
        .dout(new_Jinkela_wire_6097)
    );

    bfr new_Jinkela_buffer_11538 (
        .din(new_Jinkela_wire_13885),
        .dout(new_Jinkela_wire_13886)
    );

    bfr new_Jinkela_buffer_4542 (
        .din(new_Jinkela_wire_5931),
        .dout(new_Jinkela_wire_5932)
    );

    bfr new_Jinkela_buffer_11466 (
        .din(new_Jinkela_wire_13809),
        .dout(new_Jinkela_wire_13810)
    );

    bfr new_Jinkela_buffer_4605 (
        .din(new_Jinkela_wire_6016),
        .dout(new_Jinkela_wire_6017)
    );

    bfr new_Jinkela_buffer_11631 (
        .din(new_Jinkela_wire_14000),
        .dout(new_Jinkela_wire_14001)
    );

    bfr new_Jinkela_buffer_4543 (
        .din(new_Jinkela_wire_5932),
        .dout(new_Jinkela_wire_5933)
    );

    bfr new_Jinkela_buffer_11467 (
        .din(new_Jinkela_wire_13810),
        .dout(new_Jinkela_wire_13811)
    );

    bfr new_Jinkela_buffer_11539 (
        .din(new_Jinkela_wire_13886),
        .dout(new_Jinkela_wire_13887)
    );

    bfr new_Jinkela_buffer_4544 (
        .din(new_Jinkela_wire_5933),
        .dout(new_Jinkela_wire_5934)
    );

    bfr new_Jinkela_buffer_11468 (
        .din(new_Jinkela_wire_13811),
        .dout(new_Jinkela_wire_13812)
    );

    bfr new_Jinkela_buffer_4606 (
        .din(new_Jinkela_wire_6017),
        .dout(new_Jinkela_wire_6018)
    );

    bfr new_Jinkela_buffer_11635 (
        .din(_0632_),
        .dout(new_Jinkela_wire_14009)
    );

    spl2 new_Jinkela_splitter_1037 (
        .a(_0309_),
        .b(new_Jinkela_wire_14012),
        .c(new_Jinkela_wire_14013)
    );

    bfr new_Jinkela_buffer_4545 (
        .din(new_Jinkela_wire_5934),
        .dout(new_Jinkela_wire_5935)
    );

    bfr new_Jinkela_buffer_11469 (
        .din(new_Jinkela_wire_13812),
        .dout(new_Jinkela_wire_13813)
    );

    bfr new_Jinkela_buffer_4684 (
        .din(new_Jinkela_wire_6097),
        .dout(new_Jinkela_wire_6098)
    );

    bfr new_Jinkela_buffer_11540 (
        .din(new_Jinkela_wire_13887),
        .dout(new_Jinkela_wire_13888)
    );

    bfr new_Jinkela_buffer_4546 (
        .din(new_Jinkela_wire_5935),
        .dout(new_Jinkela_wire_5936)
    );

    bfr new_Jinkela_buffer_11470 (
        .din(new_Jinkela_wire_13813),
        .dout(new_Jinkela_wire_13814)
    );

    bfr new_Jinkela_buffer_4607 (
        .din(new_Jinkela_wire_6018),
        .dout(new_Jinkela_wire_6019)
    );

    bfr new_Jinkela_buffer_11632 (
        .din(new_Jinkela_wire_14001),
        .dout(new_Jinkela_wire_14002)
    );

    bfr new_Jinkela_buffer_4547 (
        .din(new_Jinkela_wire_5936),
        .dout(new_Jinkela_wire_5937)
    );

    bfr new_Jinkela_buffer_11471 (
        .din(new_Jinkela_wire_13814),
        .dout(new_Jinkela_wire_13815)
    );

    bfr new_Jinkela_buffer_11541 (
        .din(new_Jinkela_wire_13888),
        .dout(new_Jinkela_wire_13889)
    );

    spl2 new_Jinkela_splitter_559 (
        .a(_1731_),
        .b(new_Jinkela_wire_6202),
        .c(new_Jinkela_wire_6203)
    );

    bfr new_Jinkela_buffer_4548 (
        .din(new_Jinkela_wire_5937),
        .dout(new_Jinkela_wire_5938)
    );

    bfr new_Jinkela_buffer_11472 (
        .din(new_Jinkela_wire_13815),
        .dout(new_Jinkela_wire_13816)
    );

    bfr new_Jinkela_buffer_4608 (
        .din(new_Jinkela_wire_6019),
        .dout(new_Jinkela_wire_6020)
    );

    bfr new_Jinkela_buffer_4549 (
        .din(new_Jinkela_wire_5938),
        .dout(new_Jinkela_wire_5939)
    );

    bfr new_Jinkela_buffer_11473 (
        .din(new_Jinkela_wire_13816),
        .dout(new_Jinkela_wire_13817)
    );

    bfr new_Jinkela_buffer_4685 (
        .din(new_Jinkela_wire_6098),
        .dout(new_Jinkela_wire_6099)
    );

    bfr new_Jinkela_buffer_11542 (
        .din(new_Jinkela_wire_13889),
        .dout(new_Jinkela_wire_13890)
    );

    bfr new_Jinkela_buffer_4550 (
        .din(new_Jinkela_wire_5939),
        .dout(new_Jinkela_wire_5940)
    );

    bfr new_Jinkela_buffer_11474 (
        .din(new_Jinkela_wire_13817),
        .dout(new_Jinkela_wire_13818)
    );

    bfr new_Jinkela_buffer_4609 (
        .din(new_Jinkela_wire_6020),
        .dout(new_Jinkela_wire_6021)
    );

    bfr new_Jinkela_buffer_11633 (
        .din(new_Jinkela_wire_14002),
        .dout(new_Jinkela_wire_14003)
    );

    bfr new_Jinkela_buffer_4551 (
        .din(new_Jinkela_wire_5940),
        .dout(new_Jinkela_wire_5941)
    );

    bfr new_Jinkela_buffer_11475 (
        .din(new_Jinkela_wire_13818),
        .dout(new_Jinkela_wire_13819)
    );

    bfr new_Jinkela_buffer_4778 (
        .din(new_Jinkela_wire_6197),
        .dout(new_Jinkela_wire_6198)
    );

    bfr new_Jinkela_buffer_11543 (
        .din(new_Jinkela_wire_13890),
        .dout(new_Jinkela_wire_13891)
    );

    spl2 new_Jinkela_splitter_560 (
        .a(_0821_),
        .b(new_Jinkela_wire_6204),
        .c(new_Jinkela_wire_6205)
    );

    bfr new_Jinkela_buffer_4552 (
        .din(new_Jinkela_wire_5941),
        .dout(new_Jinkela_wire_5942)
    );

    bfr new_Jinkela_buffer_11476 (
        .din(new_Jinkela_wire_13819),
        .dout(new_Jinkela_wire_13820)
    );

    bfr new_Jinkela_buffer_4610 (
        .din(new_Jinkela_wire_6021),
        .dout(new_Jinkela_wire_6022)
    );

    spl2 new_Jinkela_splitter_1036 (
        .a(_1180_),
        .b(new_Jinkela_wire_14010),
        .c(new_Jinkela_wire_14011)
    );

    bfr new_Jinkela_buffer_4553 (
        .din(new_Jinkela_wire_5942),
        .dout(new_Jinkela_wire_5943)
    );

    bfr new_Jinkela_buffer_11477 (
        .din(new_Jinkela_wire_13820),
        .dout(new_Jinkela_wire_13821)
    );

    bfr new_Jinkela_buffer_4686 (
        .din(new_Jinkela_wire_6099),
        .dout(new_Jinkela_wire_6100)
    );

    bfr new_Jinkela_buffer_11544 (
        .din(new_Jinkela_wire_13891),
        .dout(new_Jinkela_wire_13892)
    );

    bfr new_Jinkela_buffer_4554 (
        .din(new_Jinkela_wire_5943),
        .dout(new_Jinkela_wire_5944)
    );

    bfr new_Jinkela_buffer_11478 (
        .din(new_Jinkela_wire_13821),
        .dout(new_Jinkela_wire_13822)
    );

    bfr new_Jinkela_buffer_4611 (
        .din(new_Jinkela_wire_6022),
        .dout(new_Jinkela_wire_6023)
    );

    spl2 new_Jinkela_splitter_1034 (
        .a(new_Jinkela_wire_14003),
        .b(new_Jinkela_wire_14004),
        .c(new_Jinkela_wire_14005)
    );

    bfr new_Jinkela_buffer_4555 (
        .din(new_Jinkela_wire_5944),
        .dout(new_Jinkela_wire_5945)
    );

    bfr new_Jinkela_buffer_11479 (
        .din(new_Jinkela_wire_13822),
        .dout(new_Jinkela_wire_13823)
    );

    spl2 new_Jinkela_splitter_561 (
        .a(_1139_),
        .b(new_Jinkela_wire_6238),
        .c(new_Jinkela_wire_6239)
    );

    bfr new_Jinkela_buffer_11545 (
        .din(new_Jinkela_wire_13892),
        .dout(new_Jinkela_wire_13893)
    );

    bfr new_Jinkela_buffer_4556 (
        .din(new_Jinkela_wire_5945),
        .dout(new_Jinkela_wire_5946)
    );

    bfr new_Jinkela_buffer_11480 (
        .din(new_Jinkela_wire_13823),
        .dout(new_Jinkela_wire_13824)
    );

    bfr new_Jinkela_buffer_4612 (
        .din(new_Jinkela_wire_6023),
        .dout(new_Jinkela_wire_6024)
    );

    spl2 new_Jinkela_splitter_1038 (
        .a(_0568_),
        .b(new_Jinkela_wire_14014),
        .c(new_Jinkela_wire_14015)
    );

    bfr new_Jinkela_buffer_4557 (
        .din(new_Jinkela_wire_5946),
        .dout(new_Jinkela_wire_5947)
    );

    bfr new_Jinkela_buffer_11481 (
        .din(new_Jinkela_wire_13824),
        .dout(new_Jinkela_wire_13825)
    );

    bfr new_Jinkela_buffer_4687 (
        .din(new_Jinkela_wire_6100),
        .dout(new_Jinkela_wire_6101)
    );

    bfr new_Jinkela_buffer_11546 (
        .din(new_Jinkela_wire_13893),
        .dout(new_Jinkela_wire_13894)
    );

    bfr new_Jinkela_buffer_4558 (
        .din(new_Jinkela_wire_5947),
        .dout(new_Jinkela_wire_5948)
    );

    bfr new_Jinkela_buffer_11482 (
        .din(new_Jinkela_wire_13825),
        .dout(new_Jinkela_wire_13826)
    );

    bfr new_Jinkela_buffer_4613 (
        .din(new_Jinkela_wire_6024),
        .dout(new_Jinkela_wire_6025)
    );

    bfr new_Jinkela_buffer_4559 (
        .din(new_Jinkela_wire_5948),
        .dout(new_Jinkela_wire_5949)
    );

    bfr new_Jinkela_buffer_11483 (
        .din(new_Jinkela_wire_13826),
        .dout(new_Jinkela_wire_13827)
    );

    bfr new_Jinkela_buffer_4779 (
        .din(new_Jinkela_wire_6198),
        .dout(new_Jinkela_wire_6199)
    );

    bfr new_Jinkela_buffer_11547 (
        .din(new_Jinkela_wire_13894),
        .dout(new_Jinkela_wire_13895)
    );

    bfr new_Jinkela_buffer_4560 (
        .din(new_Jinkela_wire_5949),
        .dout(new_Jinkela_wire_5950)
    );

    bfr new_Jinkela_buffer_11484 (
        .din(new_Jinkela_wire_13827),
        .dout(new_Jinkela_wire_13828)
    );

    bfr new_Jinkela_buffer_4614 (
        .din(new_Jinkela_wire_6025),
        .dout(new_Jinkela_wire_6026)
    );

    spl2 new_Jinkela_splitter_1039 (
        .a(_1539_),
        .b(new_Jinkela_wire_14017),
        .c(new_Jinkela_wire_14018)
    );

    bfr new_Jinkela_buffer_11636 (
        .din(_1490_),
        .dout(new_Jinkela_wire_14016)
    );

    bfr new_Jinkela_buffer_4561 (
        .din(new_Jinkela_wire_5950),
        .dout(new_Jinkela_wire_5951)
    );

    bfr new_Jinkela_buffer_11485 (
        .din(new_Jinkela_wire_13828),
        .dout(new_Jinkela_wire_13829)
    );

    bfr new_Jinkela_buffer_15023 (
        .din(new_Jinkela_wire_17921),
        .dout(new_Jinkela_wire_17922)
    );

    bfr new_Jinkela_buffer_14940 (
        .din(new_Jinkela_wire_17826),
        .dout(new_Jinkela_wire_17827)
    );

    bfr new_Jinkela_buffer_14981 (
        .din(new_Jinkela_wire_17877),
        .dout(new_Jinkela_wire_17878)
    );

    bfr new_Jinkela_buffer_14941 (
        .din(new_Jinkela_wire_17827),
        .dout(new_Jinkela_wire_17828)
    );

    bfr new_Jinkela_buffer_14942 (
        .din(new_Jinkela_wire_17828),
        .dout(new_Jinkela_wire_17829)
    );

    bfr new_Jinkela_buffer_14982 (
        .din(new_Jinkela_wire_17878),
        .dout(new_Jinkela_wire_17879)
    );

    bfr new_Jinkela_buffer_14943 (
        .din(new_Jinkela_wire_17829),
        .dout(new_Jinkela_wire_17830)
    );

    bfr new_Jinkela_buffer_15024 (
        .din(new_Jinkela_wire_17922),
        .dout(new_Jinkela_wire_17923)
    );

    bfr new_Jinkela_buffer_14944 (
        .din(new_Jinkela_wire_17830),
        .dout(new_Jinkela_wire_17831)
    );

    bfr new_Jinkela_buffer_14983 (
        .din(new_Jinkela_wire_17879),
        .dout(new_Jinkela_wire_17880)
    );

    bfr new_Jinkela_buffer_14945 (
        .din(new_Jinkela_wire_17831),
        .dout(new_Jinkela_wire_17832)
    );

    spl2 new_Jinkela_splitter_1305 (
        .a(_1800_),
        .b(new_Jinkela_wire_17987),
        .c(new_Jinkela_wire_17988)
    );

    bfr new_Jinkela_buffer_14946 (
        .din(new_Jinkela_wire_17832),
        .dout(new_Jinkela_wire_17833)
    );

    bfr new_Jinkela_buffer_14984 (
        .din(new_Jinkela_wire_17880),
        .dout(new_Jinkela_wire_17881)
    );

    bfr new_Jinkela_buffer_14947 (
        .din(new_Jinkela_wire_17833),
        .dout(new_Jinkela_wire_17834)
    );

    bfr new_Jinkela_buffer_15025 (
        .din(new_Jinkela_wire_17923),
        .dout(new_Jinkela_wire_17924)
    );

    bfr new_Jinkela_buffer_14948 (
        .din(new_Jinkela_wire_17834),
        .dout(new_Jinkela_wire_17835)
    );

    bfr new_Jinkela_buffer_14985 (
        .din(new_Jinkela_wire_17881),
        .dout(new_Jinkela_wire_17882)
    );

    bfr new_Jinkela_buffer_14949 (
        .din(new_Jinkela_wire_17835),
        .dout(new_Jinkela_wire_17836)
    );

    spl2 new_Jinkela_splitter_1306 (
        .a(_0572_),
        .b(new_Jinkela_wire_17989),
        .c(new_Jinkela_wire_17990)
    );

    bfr new_Jinkela_buffer_14950 (
        .din(new_Jinkela_wire_17836),
        .dout(new_Jinkela_wire_17837)
    );

    bfr new_Jinkela_buffer_14986 (
        .din(new_Jinkela_wire_17882),
        .dout(new_Jinkela_wire_17883)
    );

    bfr new_Jinkela_buffer_14951 (
        .din(new_Jinkela_wire_17837),
        .dout(new_Jinkela_wire_17838)
    );

    bfr new_Jinkela_buffer_15026 (
        .din(new_Jinkela_wire_17924),
        .dout(new_Jinkela_wire_17925)
    );

    bfr new_Jinkela_buffer_14952 (
        .din(new_Jinkela_wire_17838),
        .dout(new_Jinkela_wire_17839)
    );

    bfr new_Jinkela_buffer_14987 (
        .din(new_Jinkela_wire_17883),
        .dout(new_Jinkela_wire_17884)
    );

    bfr new_Jinkela_buffer_14953 (
        .din(new_Jinkela_wire_17839),
        .dout(new_Jinkela_wire_17840)
    );

    bfr new_Jinkela_buffer_15074 (
        .din(_0941_),
        .dout(new_Jinkela_wire_17991)
    );

    bfr new_Jinkela_buffer_14954 (
        .din(new_Jinkela_wire_17840),
        .dout(new_Jinkela_wire_17841)
    );

    bfr new_Jinkela_buffer_14988 (
        .din(new_Jinkela_wire_17884),
        .dout(new_Jinkela_wire_17885)
    );

    bfr new_Jinkela_buffer_14955 (
        .din(new_Jinkela_wire_17841),
        .dout(new_Jinkela_wire_17842)
    );

    bfr new_Jinkela_buffer_15027 (
        .din(new_Jinkela_wire_17925),
        .dout(new_Jinkela_wire_17926)
    );

    bfr new_Jinkela_buffer_14956 (
        .din(new_Jinkela_wire_17842),
        .dout(new_Jinkela_wire_17843)
    );

    bfr new_Jinkela_buffer_14989 (
        .din(new_Jinkela_wire_17885),
        .dout(new_Jinkela_wire_17886)
    );

    bfr new_Jinkela_buffer_14957 (
        .din(new_Jinkela_wire_17843),
        .dout(new_Jinkela_wire_17844)
    );

    bfr new_Jinkela_buffer_15075 (
        .din(_1155_),
        .dout(new_Jinkela_wire_17994)
    );

    spl2 new_Jinkela_splitter_1307 (
        .a(_1266_),
        .b(new_Jinkela_wire_17992),
        .c(new_Jinkela_wire_17993)
    );

    bfr new_Jinkela_buffer_14958 (
        .din(new_Jinkela_wire_17844),
        .dout(new_Jinkela_wire_17845)
    );

    bfr new_Jinkela_buffer_14990 (
        .din(new_Jinkela_wire_17886),
        .dout(new_Jinkela_wire_17887)
    );

    bfr new_Jinkela_buffer_14959 (
        .din(new_Jinkela_wire_17845),
        .dout(new_Jinkela_wire_17846)
    );

    bfr new_Jinkela_buffer_15028 (
        .din(new_Jinkela_wire_17926),
        .dout(new_Jinkela_wire_17927)
    );

    bfr new_Jinkela_buffer_14960 (
        .din(new_Jinkela_wire_17846),
        .dout(new_Jinkela_wire_17847)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(_0852_),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1739),
        .dout(new_Jinkela_wire_1740)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_1910),
        .dout(new_Jinkela_wire_1911)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1740),
        .dout(new_Jinkela_wire_1741)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1741),
        .dout(new_Jinkela_wire_1742)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_1915),
        .dout(new_Jinkela_wire_1916)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1742),
        .dout(new_Jinkela_wire_1743)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1743),
        .dout(new_Jinkela_wire_1744)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(_1721_),
        .b(new_Jinkela_wire_2117),
        .c(new_Jinkela_wire_2118)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1744),
        .dout(new_Jinkela_wire_1745)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1745),
        .dout(new_Jinkela_wire_1746)
    );

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_1916),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1830),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1746),
        .dout(new_Jinkela_wire_1747)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1747),
        .dout(new_Jinkela_wire_1748)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(_1430_),
        .dout(new_Jinkela_wire_2018)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1748),
        .dout(new_Jinkela_wire_1749)
    );

    spl2 new_Jinkela_splitter_262 (
        .a(_0442_),
        .b(new_Jinkela_wire_2016),
        .c(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1749),
        .dout(new_Jinkela_wire_1750)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(new_Jinkela_wire_1917),
        .dout(new_Jinkela_wire_1918)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1832),
        .dout(new_Jinkela_wire_1833)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1750),
        .dout(new_Jinkela_wire_1751)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1751),
        .dout(new_Jinkela_wire_1752)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1833),
        .dout(new_Jinkela_wire_1834)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1752),
        .dout(new_Jinkela_wire_1753)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1753),
        .dout(new_Jinkela_wire_1754)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_1918),
        .dout(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1834),
        .dout(new_Jinkela_wire_1835)
    );

    bfr new_Jinkela_buffer_971 (
        .din(new_Jinkela_wire_1754),
        .dout(new_Jinkela_wire_1755)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1755),
        .dout(new_Jinkela_wire_1756)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(_0621_),
        .dout(new_Jinkela_wire_2019)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1757),
        .dout(new_Jinkela_wire_1758)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_1919),
        .dout(new_Jinkela_wire_1920)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1758),
        .dout(new_Jinkela_wire_1759)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1759),
        .dout(new_Jinkela_wire_1760)
    );

    bfr new_Jinkela_buffer_11548 (
        .din(new_Jinkela_wire_13895),
        .dout(new_Jinkela_wire_13896)
    );

    bfr new_Jinkela_buffer_11486 (
        .din(new_Jinkela_wire_13829),
        .dout(new_Jinkela_wire_13830)
    );

    spl2 new_Jinkela_splitter_1040 (
        .a(_1596_),
        .b(new_Jinkela_wire_14019),
        .c(new_Jinkela_wire_14020)
    );

    bfr new_Jinkela_buffer_11487 (
        .din(new_Jinkela_wire_13830),
        .dout(new_Jinkela_wire_13831)
    );

    bfr new_Jinkela_buffer_11549 (
        .din(new_Jinkela_wire_13896),
        .dout(new_Jinkela_wire_13897)
    );

    bfr new_Jinkela_buffer_11488 (
        .din(new_Jinkela_wire_13831),
        .dout(new_Jinkela_wire_13832)
    );

    bfr new_Jinkela_buffer_11489 (
        .din(new_Jinkela_wire_13832),
        .dout(new_Jinkela_wire_13833)
    );

    bfr new_Jinkela_buffer_11550 (
        .din(new_Jinkela_wire_13897),
        .dout(new_Jinkela_wire_13898)
    );

    bfr new_Jinkela_buffer_11490 (
        .din(new_Jinkela_wire_13833),
        .dout(new_Jinkela_wire_13834)
    );

    bfr new_Jinkela_buffer_11637 (
        .din(_0181_),
        .dout(new_Jinkela_wire_14021)
    );

    bfr new_Jinkela_buffer_11491 (
        .din(new_Jinkela_wire_13834),
        .dout(new_Jinkela_wire_13835)
    );

    bfr new_Jinkela_buffer_11551 (
        .din(new_Jinkela_wire_13898),
        .dout(new_Jinkela_wire_13899)
    );

    bfr new_Jinkela_buffer_11492 (
        .din(new_Jinkela_wire_13835),
        .dout(new_Jinkela_wire_13836)
    );

    spl2 new_Jinkela_splitter_1042 (
        .a(_1376_),
        .b(new_Jinkela_wire_14024),
        .c(new_Jinkela_wire_14025)
    );

    spl2 new_Jinkela_splitter_1041 (
        .a(_0307_),
        .b(new_Jinkela_wire_14022),
        .c(new_Jinkela_wire_14023)
    );

    bfr new_Jinkela_buffer_11493 (
        .din(new_Jinkela_wire_13836),
        .dout(new_Jinkela_wire_13837)
    );

    bfr new_Jinkela_buffer_11552 (
        .din(new_Jinkela_wire_13899),
        .dout(new_Jinkela_wire_13900)
    );

    bfr new_Jinkela_buffer_11494 (
        .din(new_Jinkela_wire_13837),
        .dout(new_Jinkela_wire_13838)
    );

    bfr new_Jinkela_buffer_11495 (
        .din(new_Jinkela_wire_13838),
        .dout(new_Jinkela_wire_13839)
    );

    bfr new_Jinkela_buffer_11553 (
        .din(new_Jinkela_wire_13900),
        .dout(new_Jinkela_wire_13901)
    );

    bfr new_Jinkela_buffer_11496 (
        .din(new_Jinkela_wire_13839),
        .dout(new_Jinkela_wire_13840)
    );

    spl2 new_Jinkela_splitter_1043 (
        .a(_1444_),
        .b(new_Jinkela_wire_14026),
        .c(new_Jinkela_wire_14027)
    );

    bfr new_Jinkela_buffer_11497 (
        .din(new_Jinkela_wire_13840),
        .dout(new_Jinkela_wire_13841)
    );

    bfr new_Jinkela_buffer_11554 (
        .din(new_Jinkela_wire_13901),
        .dout(new_Jinkela_wire_13902)
    );

    bfr new_Jinkela_buffer_11498 (
        .din(new_Jinkela_wire_13841),
        .dout(new_Jinkela_wire_13842)
    );

    spl2 new_Jinkela_splitter_1044 (
        .a(_0490_),
        .b(new_Jinkela_wire_14028),
        .c(new_Jinkela_wire_14029)
    );

    bfr new_Jinkela_buffer_11499 (
        .din(new_Jinkela_wire_13842),
        .dout(new_Jinkela_wire_13843)
    );

    bfr new_Jinkela_buffer_11555 (
        .din(new_Jinkela_wire_13902),
        .dout(new_Jinkela_wire_13903)
    );

    spl2 new_Jinkela_splitter_1021 (
        .a(new_Jinkela_wire_13843),
        .b(new_Jinkela_wire_13844),
        .c(new_Jinkela_wire_13845)
    );

    bfr new_Jinkela_buffer_11556 (
        .din(new_Jinkela_wire_13903),
        .dout(new_Jinkela_wire_13904)
    );

    spl2 new_Jinkela_splitter_1045 (
        .a(_0915_),
        .b(new_Jinkela_wire_14030),
        .c(new_Jinkela_wire_14031)
    );

    spl2 new_Jinkela_splitter_1046 (
        .a(_0949_),
        .b(new_Jinkela_wire_14032),
        .c(new_Jinkela_wire_14033)
    );

    bfr new_Jinkela_buffer_11557 (
        .din(new_Jinkela_wire_13904),
        .dout(new_Jinkela_wire_13905)
    );

    spl2 new_Jinkela_splitter_1047 (
        .a(_0332_),
        .b(new_Jinkela_wire_14034),
        .c(new_Jinkela_wire_14035)
    );

    bfr new_Jinkela_buffer_11558 (
        .din(new_Jinkela_wire_13905),
        .dout(new_Jinkela_wire_13906)
    );

    spl2 new_Jinkela_splitter_1048 (
        .a(_1293_),
        .b(new_Jinkela_wire_14036),
        .c(new_Jinkela_wire_14037)
    );

    bfr new_Jinkela_buffer_11559 (
        .din(new_Jinkela_wire_13906),
        .dout(new_Jinkela_wire_13907)
    );

    bfr new_Jinkela_buffer_11638 (
        .din(new_Jinkela_wire_14039),
        .dout(new_Jinkela_wire_14040)
    );

    spl2 new_Jinkela_splitter_1049 (
        .a(_0636_),
        .b(new_Jinkela_wire_14038),
        .c(new_Jinkela_wire_14039)
    );

    bfr new_Jinkela_buffer_11560 (
        .din(new_Jinkela_wire_13907),
        .dout(new_Jinkela_wire_13908)
    );

    bfr new_Jinkela_buffer_11642 (
        .din(_1375_),
        .dout(new_Jinkela_wire_14044)
    );

    bfr new_Jinkela_buffer_11561 (
        .din(new_Jinkela_wire_13908),
        .dout(new_Jinkela_wire_13909)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    bfr new_Jinkela_buffer_4688 (
        .din(new_Jinkela_wire_6101),
        .dout(new_Jinkela_wire_6102)
    );

    bfr new_Jinkela_buffer_14991 (
        .din(new_Jinkela_wire_17887),
        .dout(new_Jinkela_wire_17888)
    );

    spl2 new_Jinkela_splitter_241 (
        .a(new_Jinkela_wire_1760),
        .b(new_Jinkela_wire_1761),
        .c(new_Jinkela_wire_1762)
    );

    bfr new_Jinkela_buffer_4562 (
        .din(new_Jinkela_wire_5951),
        .dout(new_Jinkela_wire_5952)
    );

    bfr new_Jinkela_buffer_14961 (
        .din(new_Jinkela_wire_17847),
        .dout(new_Jinkela_wire_17848)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_1920),
        .dout(new_Jinkela_wire_1921)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1838),
        .dout(new_Jinkela_wire_1839)
    );

    bfr new_Jinkela_buffer_4615 (
        .din(new_Jinkela_wire_6026),
        .dout(new_Jinkela_wire_6027)
    );

    bfr new_Jinkela_buffer_15076 (
        .din(_0434_),
        .dout(new_Jinkela_wire_17997)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(_0951_),
        .dout(new_Jinkela_wire_2119)
    );

    bfr new_Jinkela_buffer_4563 (
        .din(new_Jinkela_wire_5952),
        .dout(new_Jinkela_wire_5953)
    );

    bfr new_Jinkela_buffer_14962 (
        .din(new_Jinkela_wire_17848),
        .dout(new_Jinkela_wire_17849)
    );

    bfr new_Jinkela_buffer_4782 (
        .din(new_Jinkela_wire_6205),
        .dout(new_Jinkela_wire_6206)
    );

    bfr new_Jinkela_buffer_14992 (
        .din(new_Jinkela_wire_17888),
        .dout(new_Jinkela_wire_17889)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_2019),
        .dout(new_Jinkela_wire_2020)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1839),
        .dout(new_Jinkela_wire_1840)
    );

    bfr new_Jinkela_buffer_4564 (
        .din(new_Jinkela_wire_5953),
        .dout(new_Jinkela_wire_5954)
    );

    bfr new_Jinkela_buffer_14963 (
        .din(new_Jinkela_wire_17849),
        .dout(new_Jinkela_wire_17850)
    );

    bfr new_Jinkela_buffer_4616 (
        .din(new_Jinkela_wire_6027),
        .dout(new_Jinkela_wire_6028)
    );

    bfr new_Jinkela_buffer_15029 (
        .din(new_Jinkela_wire_17927),
        .dout(new_Jinkela_wire_17928)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_1921),
        .dout(new_Jinkela_wire_1922)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1840),
        .dout(new_Jinkela_wire_1841)
    );

    bfr new_Jinkela_buffer_4565 (
        .din(new_Jinkela_wire_5954),
        .dout(new_Jinkela_wire_5955)
    );

    bfr new_Jinkela_buffer_14964 (
        .din(new_Jinkela_wire_17850),
        .dout(new_Jinkela_wire_17851)
    );

    bfr new_Jinkela_buffer_4689 (
        .din(new_Jinkela_wire_6102),
        .dout(new_Jinkela_wire_6103)
    );

    bfr new_Jinkela_buffer_14993 (
        .din(new_Jinkela_wire_17889),
        .dout(new_Jinkela_wire_17890)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1841),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_4566 (
        .din(new_Jinkela_wire_5955),
        .dout(new_Jinkela_wire_5956)
    );

    bfr new_Jinkela_buffer_14965 (
        .din(new_Jinkela_wire_17851),
        .dout(new_Jinkela_wire_17852)
    );

    bfr new_Jinkela_buffer_4617 (
        .din(new_Jinkela_wire_6028),
        .dout(new_Jinkela_wire_6029)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_1922),
        .dout(new_Jinkela_wire_1923)
    );

    spl2 new_Jinkela_splitter_1308 (
        .a(_0311_),
        .b(new_Jinkela_wire_17995),
        .c(new_Jinkela_wire_17996)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1842),
        .dout(new_Jinkela_wire_1843)
    );

    bfr new_Jinkela_buffer_4567 (
        .din(new_Jinkela_wire_5956),
        .dout(new_Jinkela_wire_5957)
    );

    bfr new_Jinkela_buffer_14966 (
        .din(new_Jinkela_wire_17852),
        .dout(new_Jinkela_wire_17853)
    );

    bfr new_Jinkela_buffer_4780 (
        .din(new_Jinkela_wire_6199),
        .dout(new_Jinkela_wire_6200)
    );

    bfr new_Jinkela_buffer_14994 (
        .din(new_Jinkela_wire_17890),
        .dout(new_Jinkela_wire_17891)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_2020),
        .dout(new_Jinkela_wire_2021)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1843),
        .dout(new_Jinkela_wire_1844)
    );

    bfr new_Jinkela_buffer_4568 (
        .din(new_Jinkela_wire_5957),
        .dout(new_Jinkela_wire_5958)
    );

    bfr new_Jinkela_buffer_14967 (
        .din(new_Jinkela_wire_17853),
        .dout(new_Jinkela_wire_17854)
    );

    bfr new_Jinkela_buffer_4618 (
        .din(new_Jinkela_wire_6029),
        .dout(new_Jinkela_wire_6030)
    );

    bfr new_Jinkela_buffer_15030 (
        .din(new_Jinkela_wire_17928),
        .dout(new_Jinkela_wire_17929)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_1923),
        .dout(new_Jinkela_wire_1924)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1844),
        .dout(new_Jinkela_wire_1845)
    );

    bfr new_Jinkela_buffer_4569 (
        .din(new_Jinkela_wire_5958),
        .dout(new_Jinkela_wire_5959)
    );

    bfr new_Jinkela_buffer_14968 (
        .din(new_Jinkela_wire_17854),
        .dout(new_Jinkela_wire_17855)
    );

    bfr new_Jinkela_buffer_4690 (
        .din(new_Jinkela_wire_6103),
        .dout(new_Jinkela_wire_6104)
    );

    bfr new_Jinkela_buffer_14995 (
        .din(new_Jinkela_wire_17891),
        .dout(new_Jinkela_wire_17892)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(_0786_),
        .dout(new_Jinkela_wire_2122)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(new_Jinkela_wire_1845),
        .dout(new_Jinkela_wire_1846)
    );

    bfr new_Jinkela_buffer_4570 (
        .din(new_Jinkela_wire_5959),
        .dout(new_Jinkela_wire_5960)
    );

    spl2 new_Jinkela_splitter_1292 (
        .a(new_Jinkela_wire_17855),
        .b(new_Jinkela_wire_17856),
        .c(new_Jinkela_wire_17857)
    );

    spl2 new_Jinkela_splitter_265 (
        .a(_1675_),
        .b(new_Jinkela_wire_2120),
        .c(new_Jinkela_wire_2121)
    );

    bfr new_Jinkela_buffer_4619 (
        .din(new_Jinkela_wire_6030),
        .dout(new_Jinkela_wire_6031)
    );

    bfr new_Jinkela_buffer_14996 (
        .din(new_Jinkela_wire_17892),
        .dout(new_Jinkela_wire_17893)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_1924),
        .dout(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1846),
        .dout(new_Jinkela_wire_1847)
    );

    bfr new_Jinkela_buffer_4571 (
        .din(new_Jinkela_wire_5960),
        .dout(new_Jinkela_wire_5961)
    );

    spl2 new_Jinkela_splitter_1310 (
        .a(_1366_),
        .b(new_Jinkela_wire_18104),
        .c(new_Jinkela_wire_18105)
    );

    bfr new_Jinkela_buffer_15031 (
        .din(new_Jinkela_wire_17929),
        .dout(new_Jinkela_wire_17930)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(new_Jinkela_wire_2021),
        .dout(new_Jinkela_wire_2022)
    );

    spl2 new_Jinkela_splitter_562 (
        .a(_0407_),
        .b(new_Jinkela_wire_6240),
        .c(new_Jinkela_wire_6241)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(new_Jinkela_wire_1847),
        .dout(new_Jinkela_wire_1848)
    );

    bfr new_Jinkela_buffer_4572 (
        .din(new_Jinkela_wire_5961),
        .dout(new_Jinkela_wire_5962)
    );

    bfr new_Jinkela_buffer_14997 (
        .din(new_Jinkela_wire_17893),
        .dout(new_Jinkela_wire_17894)
    );

    bfr new_Jinkela_buffer_4620 (
        .din(new_Jinkela_wire_6031),
        .dout(new_Jinkela_wire_6032)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_1925),
        .dout(new_Jinkela_wire_1926)
    );

    bfr new_Jinkela_buffer_15180 (
        .din(_1158_),
        .dout(new_Jinkela_wire_18103)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(new_Jinkela_wire_1848),
        .dout(new_Jinkela_wire_1849)
    );

    bfr new_Jinkela_buffer_4573 (
        .din(new_Jinkela_wire_5962),
        .dout(new_Jinkela_wire_5963)
    );

    bfr new_Jinkela_buffer_14998 (
        .din(new_Jinkela_wire_17894),
        .dout(new_Jinkela_wire_17895)
    );

    bfr new_Jinkela_buffer_4691 (
        .din(new_Jinkela_wire_6104),
        .dout(new_Jinkela_wire_6105)
    );

    bfr new_Jinkela_buffer_15032 (
        .din(new_Jinkela_wire_17930),
        .dout(new_Jinkela_wire_17931)
    );

    spl2 new_Jinkela_splitter_266 (
        .a(_1009_),
        .b(new_Jinkela_wire_2124),
        .c(new_Jinkela_wire_2125)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1849),
        .dout(new_Jinkela_wire_1850)
    );

    bfr new_Jinkela_buffer_4574 (
        .din(new_Jinkela_wire_5963),
        .dout(new_Jinkela_wire_5964)
    );

    bfr new_Jinkela_buffer_14999 (
        .din(new_Jinkela_wire_17895),
        .dout(new_Jinkela_wire_17896)
    );

    bfr new_Jinkela_buffer_4621 (
        .din(new_Jinkela_wire_6032),
        .dout(new_Jinkela_wire_6033)
    );

    bfr new_Jinkela_buffer_15077 (
        .din(new_Jinkela_wire_17997),
        .dout(new_Jinkela_wire_17998)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_1926),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1850),
        .dout(new_Jinkela_wire_1851)
    );

    spl2 new_Jinkela_splitter_544 (
        .a(new_Jinkela_wire_5964),
        .b(new_Jinkela_wire_5965),
        .c(new_Jinkela_wire_5966)
    );

    bfr new_Jinkela_buffer_15000 (
        .din(new_Jinkela_wire_17896),
        .dout(new_Jinkela_wire_17897)
    );

    bfr new_Jinkela_buffer_4622 (
        .din(new_Jinkela_wire_6033),
        .dout(new_Jinkela_wire_6034)
    );

    bfr new_Jinkela_buffer_15033 (
        .din(new_Jinkela_wire_17931),
        .dout(new_Jinkela_wire_17932)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1851),
        .dout(new_Jinkela_wire_1852)
    );

    bfr new_Jinkela_buffer_4781 (
        .din(new_Jinkela_wire_6200),
        .dout(new_Jinkela_wire_6201)
    );

    bfr new_Jinkela_buffer_15001 (
        .din(new_Jinkela_wire_17897),
        .dout(new_Jinkela_wire_17898)
    );

    bfr new_Jinkela_buffer_4692 (
        .din(new_Jinkela_wire_6105),
        .dout(new_Jinkela_wire_6106)
    );

    bfr new_Jinkela_buffer_15181 (
        .din(_1197_),
        .dout(new_Jinkela_wire_18106)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1852),
        .dout(new_Jinkela_wire_1853)
    );

    bfr new_Jinkela_buffer_4623 (
        .din(new_Jinkela_wire_6034),
        .dout(new_Jinkela_wire_6035)
    );

    bfr new_Jinkela_buffer_15002 (
        .din(new_Jinkela_wire_17898),
        .dout(new_Jinkela_wire_17899)
    );

    bfr new_Jinkela_buffer_15034 (
        .din(new_Jinkela_wire_17932),
        .dout(new_Jinkela_wire_17933)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1853),
        .dout(new_Jinkela_wire_1854)
    );

    bfr new_Jinkela_buffer_4624 (
        .din(new_Jinkela_wire_6035),
        .dout(new_Jinkela_wire_6036)
    );

    bfr new_Jinkela_buffer_15003 (
        .din(new_Jinkela_wire_17899),
        .dout(new_Jinkela_wire_17900)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(_1122_),
        .dout(new_Jinkela_wire_2123)
    );

    bfr new_Jinkela_buffer_4693 (
        .din(new_Jinkela_wire_6106),
        .dout(new_Jinkela_wire_6107)
    );

    bfr new_Jinkela_buffer_15078 (
        .din(new_Jinkela_wire_17998),
        .dout(new_Jinkela_wire_17999)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_1928),
        .dout(new_Jinkela_wire_1929)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1854),
        .dout(new_Jinkela_wire_1855)
    );

    bfr new_Jinkela_buffer_4625 (
        .din(new_Jinkela_wire_6036),
        .dout(new_Jinkela_wire_6037)
    );

    bfr new_Jinkela_buffer_15004 (
        .din(new_Jinkela_wire_17900),
        .dout(new_Jinkela_wire_17901)
    );

    bfr new_Jinkela_buffer_4783 (
        .din(new_Jinkela_wire_6206),
        .dout(new_Jinkela_wire_6207)
    );

    bfr new_Jinkela_buffer_15035 (
        .din(new_Jinkela_wire_17933),
        .dout(new_Jinkela_wire_17934)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_2023),
        .dout(new_Jinkela_wire_2024)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1855),
        .dout(new_Jinkela_wire_1856)
    );

    bfr new_Jinkela_buffer_4626 (
        .din(new_Jinkela_wire_6037),
        .dout(new_Jinkela_wire_6038)
    );

    bfr new_Jinkela_buffer_15005 (
        .din(new_Jinkela_wire_17901),
        .dout(new_Jinkela_wire_17902)
    );

    bfr new_Jinkela_buffer_4694 (
        .din(new_Jinkela_wire_6107),
        .dout(new_Jinkela_wire_6108)
    );

    bfr new_Jinkela_buffer_15182 (
        .din(_0059_),
        .dout(new_Jinkela_wire_18107)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_1929),
        .dout(new_Jinkela_wire_1930)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1856),
        .dout(new_Jinkela_wire_1857)
    );

    bfr new_Jinkela_buffer_4627 (
        .din(new_Jinkela_wire_6038),
        .dout(new_Jinkela_wire_6039)
    );

    bfr new_Jinkela_buffer_15006 (
        .din(new_Jinkela_wire_17902),
        .dout(new_Jinkela_wire_17903)
    );

    spl2 new_Jinkela_splitter_564 (
        .a(_0662_),
        .b(new_Jinkela_wire_6248),
        .c(new_Jinkela_wire_6249)
    );

    bfr new_Jinkela_buffer_15036 (
        .din(new_Jinkela_wire_17934),
        .dout(new_Jinkela_wire_17935)
    );

    spl2 new_Jinkela_splitter_267 (
        .a(_0843_),
        .b(new_Jinkela_wire_2126),
        .c(new_Jinkela_wire_2127)
    );

    spl2 new_Jinkela_splitter_563 (
        .a(_1190_),
        .b(new_Jinkela_wire_6242),
        .c(new_Jinkela_wire_6243)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1857),
        .dout(new_Jinkela_wire_1858)
    );

    bfr new_Jinkela_buffer_4628 (
        .din(new_Jinkela_wire_6039),
        .dout(new_Jinkela_wire_6040)
    );

    bfr new_Jinkela_buffer_15007 (
        .din(new_Jinkela_wire_17903),
        .dout(new_Jinkela_wire_17904)
    );

    spl2 new_Jinkela_splitter_795 (
        .a(new_Jinkela_wire_10076),
        .b(new_Jinkela_wire_10077),
        .c(new_Jinkela_wire_10078)
    );

    bfr new_Jinkela_buffer_8052 (
        .din(new_Jinkela_wire_9933),
        .dout(new_Jinkela_wire_9934)
    );

    bfr new_Jinkela_buffer_8053 (
        .din(new_Jinkela_wire_9934),
        .dout(new_Jinkela_wire_9935)
    );

    spl2 new_Jinkela_splitter_798 (
        .a(_0715_),
        .b(new_Jinkela_wire_10083),
        .c(new_Jinkela_wire_10084)
    );

    bfr new_Jinkela_buffer_8054 (
        .din(new_Jinkela_wire_9935),
        .dout(new_Jinkela_wire_9936)
    );

    bfr new_Jinkela_buffer_8055 (
        .din(new_Jinkela_wire_9936),
        .dout(new_Jinkela_wire_9937)
    );

    spl2 new_Jinkela_splitter_799 (
        .a(_1344_),
        .b(new_Jinkela_wire_10085),
        .c(new_Jinkela_wire_10086)
    );

    bfr new_Jinkela_buffer_8056 (
        .din(new_Jinkela_wire_9937),
        .dout(new_Jinkela_wire_9938)
    );

    spl2 new_Jinkela_splitter_800 (
        .a(_1417_),
        .b(new_Jinkela_wire_10091),
        .c(new_Jinkela_wire_10092)
    );

    bfr new_Jinkela_buffer_8185 (
        .din(new_Jinkela_wire_10086),
        .dout(new_Jinkela_wire_10087)
    );

    bfr new_Jinkela_buffer_8057 (
        .din(new_Jinkela_wire_9938),
        .dout(new_Jinkela_wire_9939)
    );

    spl2 new_Jinkela_splitter_801 (
        .a(_0990_),
        .b(new_Jinkela_wire_10097),
        .c(new_Jinkela_wire_10098)
    );

    bfr new_Jinkela_buffer_8058 (
        .din(new_Jinkela_wire_9939),
        .dout(new_Jinkela_wire_9940)
    );

    bfr new_Jinkela_buffer_8186 (
        .din(new_Jinkela_wire_10087),
        .dout(new_Jinkela_wire_10088)
    );

    bfr new_Jinkela_buffer_8059 (
        .din(new_Jinkela_wire_9940),
        .dout(new_Jinkela_wire_9941)
    );

    bfr new_Jinkela_buffer_8189 (
        .din(new_Jinkela_wire_10092),
        .dout(new_Jinkela_wire_10093)
    );

    bfr new_Jinkela_buffer_8060 (
        .din(new_Jinkela_wire_9941),
        .dout(new_Jinkela_wire_9942)
    );

    spl2 new_Jinkela_splitter_802 (
        .a(_0497_),
        .b(new_Jinkela_wire_10099),
        .c(new_Jinkela_wire_10100)
    );

    bfr new_Jinkela_buffer_8187 (
        .din(new_Jinkela_wire_10088),
        .dout(new_Jinkela_wire_10089)
    );

    bfr new_Jinkela_buffer_8061 (
        .din(new_Jinkela_wire_9942),
        .dout(new_Jinkela_wire_9943)
    );

    bfr new_Jinkela_buffer_8062 (
        .din(new_Jinkela_wire_9943),
        .dout(new_Jinkela_wire_9944)
    );

    bfr new_Jinkela_buffer_8188 (
        .din(new_Jinkela_wire_10089),
        .dout(new_Jinkela_wire_10090)
    );

    bfr new_Jinkela_buffer_8063 (
        .din(new_Jinkela_wire_9944),
        .dout(new_Jinkela_wire_9945)
    );

    bfr new_Jinkela_buffer_8190 (
        .din(new_Jinkela_wire_10093),
        .dout(new_Jinkela_wire_10094)
    );

    bfr new_Jinkela_buffer_8064 (
        .din(new_Jinkela_wire_9945),
        .dout(new_Jinkela_wire_9946)
    );

    bfr new_Jinkela_buffer_8065 (
        .din(new_Jinkela_wire_9946),
        .dout(new_Jinkela_wire_9947)
    );

    bfr new_Jinkela_buffer_8193 (
        .din(_1657_),
        .dout(new_Jinkela_wire_10101)
    );

    bfr new_Jinkela_buffer_8191 (
        .din(new_Jinkela_wire_10094),
        .dout(new_Jinkela_wire_10095)
    );

    bfr new_Jinkela_buffer_8066 (
        .din(new_Jinkela_wire_9947),
        .dout(new_Jinkela_wire_9948)
    );

    spl2 new_Jinkela_splitter_804 (
        .a(_1833_),
        .b(new_Jinkela_wire_10104),
        .c(new_Jinkela_wire_10105)
    );

    bfr new_Jinkela_buffer_8067 (
        .din(new_Jinkela_wire_9948),
        .dout(new_Jinkela_wire_9949)
    );

    spl2 new_Jinkela_splitter_803 (
        .a(_0866_),
        .b(new_Jinkela_wire_10102),
        .c(new_Jinkela_wire_10103)
    );

    bfr new_Jinkela_buffer_8192 (
        .din(new_Jinkela_wire_10095),
        .dout(new_Jinkela_wire_10096)
    );

    bfr new_Jinkela_buffer_8068 (
        .din(new_Jinkela_wire_9949),
        .dout(new_Jinkela_wire_9950)
    );

    bfr new_Jinkela_buffer_8069 (
        .din(new_Jinkela_wire_9950),
        .dout(new_Jinkela_wire_9951)
    );

    bfr new_Jinkela_buffer_8070 (
        .din(new_Jinkela_wire_9951),
        .dout(new_Jinkela_wire_9952)
    );

    spl2 new_Jinkela_splitter_805 (
        .a(_0746_),
        .b(new_Jinkela_wire_10106),
        .c(new_Jinkela_wire_10107)
    );

    bfr new_Jinkela_buffer_8071 (
        .din(new_Jinkela_wire_9952),
        .dout(new_Jinkela_wire_9953)
    );

    spl2 new_Jinkela_splitter_806 (
        .a(_0294_),
        .b(new_Jinkela_wire_10112),
        .c(new_Jinkela_wire_10113)
    );

    bfr new_Jinkela_buffer_8194 (
        .din(new_Jinkela_wire_10107),
        .dout(new_Jinkela_wire_10108)
    );

    bfr new_Jinkela_buffer_8072 (
        .din(new_Jinkela_wire_9953),
        .dout(new_Jinkela_wire_9954)
    );

    spl2 new_Jinkela_splitter_807 (
        .a(_0698_),
        .b(new_Jinkela_wire_10114),
        .c(new_Jinkela_wire_10115)
    );

    bfr new_Jinkela_buffer_8073 (
        .din(new_Jinkela_wire_9954),
        .dout(new_Jinkela_wire_9955)
    );

    bfr new_Jinkela_buffer_8195 (
        .din(new_Jinkela_wire_10108),
        .dout(new_Jinkela_wire_10109)
    );

    bfr new_Jinkela_buffer_8074 (
        .din(new_Jinkela_wire_9955),
        .dout(new_Jinkela_wire_9956)
    );

    bfr new_Jinkela_buffer_8075 (
        .din(new_Jinkela_wire_9956),
        .dout(new_Jinkela_wire_9957)
    );

    spl2 new_Jinkela_splitter_808 (
        .a(_0658_),
        .b(new_Jinkela_wire_10116),
        .c(new_Jinkela_wire_10117)
    );

    bfr new_Jinkela_buffer_8196 (
        .din(new_Jinkela_wire_10109),
        .dout(new_Jinkela_wire_10110)
    );

    bfr new_Jinkela_buffer_8076 (
        .din(new_Jinkela_wire_9957),
        .dout(new_Jinkela_wire_9958)
    );

    bfr new_Jinkela_buffer_8077 (
        .din(new_Jinkela_wire_9958),
        .dout(new_Jinkela_wire_9959)
    );

    spl2 new_Jinkela_splitter_809 (
        .a(_0043_),
        .b(new_Jinkela_wire_10118),
        .c(new_Jinkela_wire_10119)
    );

    bfr new_Jinkela_buffer_8197 (
        .din(new_Jinkela_wire_10110),
        .dout(new_Jinkela_wire_10111)
    );

    bfr new_Jinkela_buffer_8078 (
        .din(new_Jinkela_wire_9959),
        .dout(new_Jinkela_wire_9960)
    );

    bfr new_Jinkela_buffer_8278 (
        .din(_0554_),
        .dout(new_Jinkela_wire_10204)
    );

    bfr new_Jinkela_buffer_8079 (
        .din(new_Jinkela_wire_9960),
        .dout(new_Jinkela_wire_9961)
    );

    bfr new_Jinkela_buffer_8198 (
        .din(_1022_),
        .dout(new_Jinkela_wire_10120)
    );

    bfr new_Jinkela_buffer_8080 (
        .din(new_Jinkela_wire_9961),
        .dout(new_Jinkela_wire_9962)
    );

    bfr new_Jinkela_buffer_8238 (
        .din(_0232_),
        .dout(new_Jinkela_wire_10162)
    );

    bfr new_Jinkela_buffer_8199 (
        .din(new_Jinkela_wire_10120),
        .dout(new_Jinkela_wire_10121)
    );

    bfr new_Jinkela_buffer_8081 (
        .din(new_Jinkela_wire_9962),
        .dout(new_Jinkela_wire_9963)
    );

    bfr new_Jinkela_buffer_8082 (
        .din(new_Jinkela_wire_9963),
        .dout(new_Jinkela_wire_9964)
    );

    spl2 new_Jinkela_splitter_812 (
        .a(_1260_),
        .b(new_Jinkela_wire_10205),
        .c(new_Jinkela_wire_10206)
    );

    bfr new_Jinkela_buffer_8200 (
        .din(new_Jinkela_wire_10121),
        .dout(new_Jinkela_wire_10122)
    );

    bfr new_Jinkela_buffer_8083 (
        .din(new_Jinkela_wire_9964),
        .dout(new_Jinkela_wire_9965)
    );

    bfr new_Jinkela_buffer_8239 (
        .din(new_Jinkela_wire_10162),
        .dout(new_Jinkela_wire_10163)
    );

    bfr new_Jinkela_buffer_8084 (
        .din(new_Jinkela_wire_9965),
        .dout(new_Jinkela_wire_9966)
    );

    bfr new_Jinkela_buffer_8201 (
        .din(new_Jinkela_wire_10122),
        .dout(new_Jinkela_wire_10123)
    );

    bfr new_Jinkela_buffer_8085 (
        .din(new_Jinkela_wire_9966),
        .dout(new_Jinkela_wire_9967)
    );

    bfr new_Jinkela_buffer_8279 (
        .din(_1695_),
        .dout(new_Jinkela_wire_10207)
    );

    bfr new_Jinkela_buffer_8086 (
        .din(new_Jinkela_wire_9967),
        .dout(new_Jinkela_wire_9968)
    );

    bfr new_Jinkela_buffer_8202 (
        .din(new_Jinkela_wire_10123),
        .dout(new_Jinkela_wire_10124)
    );

    bfr new_Jinkela_buffer_8087 (
        .din(new_Jinkela_wire_9968),
        .dout(new_Jinkela_wire_9969)
    );

    bfr new_Jinkela_buffer_8240 (
        .din(new_Jinkela_wire_10163),
        .dout(new_Jinkela_wire_10164)
    );

    bfr new_Jinkela_buffer_8088 (
        .din(new_Jinkela_wire_9969),
        .dout(new_Jinkela_wire_9970)
    );

    bfr new_Jinkela_buffer_8203 (
        .din(new_Jinkela_wire_10124),
        .dout(new_Jinkela_wire_10125)
    );

    bfr new_Jinkela_buffer_8089 (
        .din(new_Jinkela_wire_9970),
        .dout(new_Jinkela_wire_9971)
    );

    spl2 new_Jinkela_splitter_814 (
        .a(_1515_),
        .b(new_Jinkela_wire_10257),
        .c(new_Jinkela_wire_10258)
    );

    bfr new_Jinkela_buffer_8090 (
        .din(new_Jinkela_wire_9971),
        .dout(new_Jinkela_wire_9972)
    );

    bfr new_Jinkela_buffer_8204 (
        .din(new_Jinkela_wire_10125),
        .dout(new_Jinkela_wire_10126)
    );

    bfr new_Jinkela_buffer_8091 (
        .din(new_Jinkela_wire_9972),
        .dout(new_Jinkela_wire_9973)
    );

    bfr new_Jinkela_buffer_8241 (
        .din(new_Jinkela_wire_10164),
        .dout(new_Jinkela_wire_10165)
    );

    bfr new_Jinkela_buffer_8092 (
        .din(new_Jinkela_wire_9973),
        .dout(new_Jinkela_wire_9974)
    );

    bfr new_Jinkela_buffer_8205 (
        .din(new_Jinkela_wire_10126),
        .dout(new_Jinkela_wire_10127)
    );

    bfr new_Jinkela_buffer_8093 (
        .din(new_Jinkela_wire_9974),
        .dout(new_Jinkela_wire_9975)
    );

    bfr new_Jinkela_buffer_15079 (
        .din(new_Jinkela_wire_17999),
        .dout(new_Jinkela_wire_18000)
    );

    bfr new_Jinkela_buffer_15008 (
        .din(new_Jinkela_wire_17904),
        .dout(new_Jinkela_wire_17905)
    );

    bfr new_Jinkela_buffer_15037 (
        .din(new_Jinkela_wire_17935),
        .dout(new_Jinkela_wire_17936)
    );

    bfr new_Jinkela_buffer_15009 (
        .din(new_Jinkela_wire_17905),
        .dout(new_Jinkela_wire_17906)
    );

    bfr new_Jinkela_buffer_15183 (
        .din(_1559_),
        .dout(new_Jinkela_wire_18108)
    );

    bfr new_Jinkela_buffer_15010 (
        .din(new_Jinkela_wire_17906),
        .dout(new_Jinkela_wire_17907)
    );

    bfr new_Jinkela_buffer_15038 (
        .din(new_Jinkela_wire_17936),
        .dout(new_Jinkela_wire_17937)
    );

    bfr new_Jinkela_buffer_15011 (
        .din(new_Jinkela_wire_17907),
        .dout(new_Jinkela_wire_17908)
    );

    bfr new_Jinkela_buffer_15080 (
        .din(new_Jinkela_wire_18000),
        .dout(new_Jinkela_wire_18001)
    );

    bfr new_Jinkela_buffer_15012 (
        .din(new_Jinkela_wire_17908),
        .dout(new_Jinkela_wire_17909)
    );

    bfr new_Jinkela_buffer_15039 (
        .din(new_Jinkela_wire_17937),
        .dout(new_Jinkela_wire_17938)
    );

    bfr new_Jinkela_buffer_15013 (
        .din(new_Jinkela_wire_17909),
        .dout(new_Jinkela_wire_17910)
    );

    spl2 new_Jinkela_splitter_1311 (
        .a(_1031_),
        .b(new_Jinkela_wire_18109),
        .c(new_Jinkela_wire_18110)
    );

    bfr new_Jinkela_buffer_15014 (
        .din(new_Jinkela_wire_17910),
        .dout(new_Jinkela_wire_17911)
    );

    bfr new_Jinkela_buffer_15040 (
        .din(new_Jinkela_wire_17938),
        .dout(new_Jinkela_wire_17939)
    );

    bfr new_Jinkela_buffer_15015 (
        .din(new_Jinkela_wire_17911),
        .dout(new_Jinkela_wire_17912)
    );

    bfr new_Jinkela_buffer_15081 (
        .din(new_Jinkela_wire_18001),
        .dout(new_Jinkela_wire_18002)
    );

    bfr new_Jinkela_buffer_15016 (
        .din(new_Jinkela_wire_17912),
        .dout(new_Jinkela_wire_17913)
    );

    bfr new_Jinkela_buffer_15041 (
        .din(new_Jinkela_wire_17939),
        .dout(new_Jinkela_wire_17940)
    );

    bfr new_Jinkela_buffer_15017 (
        .din(new_Jinkela_wire_17913),
        .dout(new_Jinkela_wire_17914)
    );

    spl2 new_Jinkela_splitter_1312 (
        .a(_0488_),
        .b(new_Jinkela_wire_18111),
        .c(new_Jinkela_wire_18112)
    );

    spl2 new_Jinkela_splitter_1297 (
        .a(new_Jinkela_wire_17914),
        .b(new_Jinkela_wire_17915),
        .c(new_Jinkela_wire_17916)
    );

    bfr new_Jinkela_buffer_15082 (
        .din(new_Jinkela_wire_18002),
        .dout(new_Jinkela_wire_18003)
    );

    bfr new_Jinkela_buffer_15042 (
        .din(new_Jinkela_wire_17940),
        .dout(new_Jinkela_wire_17941)
    );

    bfr new_Jinkela_buffer_15043 (
        .din(new_Jinkela_wire_17941),
        .dout(new_Jinkela_wire_17942)
    );

    bfr new_Jinkela_buffer_15044 (
        .din(new_Jinkela_wire_17942),
        .dout(new_Jinkela_wire_17943)
    );

    bfr new_Jinkela_buffer_15083 (
        .din(new_Jinkela_wire_18003),
        .dout(new_Jinkela_wire_18004)
    );

    bfr new_Jinkela_buffer_15045 (
        .din(new_Jinkela_wire_17943),
        .dout(new_Jinkela_wire_17944)
    );

    spl2 new_Jinkela_splitter_1313 (
        .a(_0560_),
        .b(new_Jinkela_wire_18117),
        .c(new_Jinkela_wire_18118)
    );

    bfr new_Jinkela_buffer_15046 (
        .din(new_Jinkela_wire_17944),
        .dout(new_Jinkela_wire_17945)
    );

    bfr new_Jinkela_buffer_15084 (
        .din(new_Jinkela_wire_18004),
        .dout(new_Jinkela_wire_18005)
    );

    bfr new_Jinkela_buffer_15047 (
        .din(new_Jinkela_wire_17945),
        .dout(new_Jinkela_wire_17946)
    );

    bfr new_Jinkela_buffer_15184 (
        .din(new_Jinkela_wire_18112),
        .dout(new_Jinkela_wire_18113)
    );

    spl2 new_Jinkela_splitter_1314 (
        .a(_0028_),
        .b(new_Jinkela_wire_18119),
        .c(new_Jinkela_wire_18120)
    );

    bfr new_Jinkela_buffer_15048 (
        .din(new_Jinkela_wire_17946),
        .dout(new_Jinkela_wire_17947)
    );

    bfr new_Jinkela_buffer_15085 (
        .din(new_Jinkela_wire_18005),
        .dout(new_Jinkela_wire_18006)
    );

    bfr new_Jinkela_buffer_15049 (
        .din(new_Jinkela_wire_17947),
        .dout(new_Jinkela_wire_17948)
    );

    bfr new_Jinkela_buffer_15188 (
        .din(_1152_),
        .dout(new_Jinkela_wire_18121)
    );

    bfr new_Jinkela_buffer_15050 (
        .din(new_Jinkela_wire_17948),
        .dout(new_Jinkela_wire_17949)
    );

    bfr new_Jinkela_buffer_15086 (
        .din(new_Jinkela_wire_18006),
        .dout(new_Jinkela_wire_18007)
    );

    bfr new_Jinkela_buffer_15051 (
        .din(new_Jinkela_wire_17949),
        .dout(new_Jinkela_wire_17950)
    );

    bfr new_Jinkela_buffer_15185 (
        .din(new_Jinkela_wire_18113),
        .dout(new_Jinkela_wire_18114)
    );

    bfr new_Jinkela_buffer_4695 (
        .din(new_Jinkela_wire_6108),
        .dout(new_Jinkela_wire_6109)
    );

    bfr new_Jinkela_buffer_11674 (
        .din(_0899_),
        .dout(new_Jinkela_wire_14078)
    );

    bfr new_Jinkela_buffer_4629 (
        .din(new_Jinkela_wire_6040),
        .dout(new_Jinkela_wire_6041)
    );

    bfr new_Jinkela_buffer_11562 (
        .din(new_Jinkela_wire_13909),
        .dout(new_Jinkela_wire_13910)
    );

    bfr new_Jinkela_buffer_4784 (
        .din(new_Jinkela_wire_6207),
        .dout(new_Jinkela_wire_6208)
    );

    bfr new_Jinkela_buffer_11681 (
        .din(_0839_),
        .dout(new_Jinkela_wire_14089)
    );

    bfr new_Jinkela_buffer_11675 (
        .din(_0461_),
        .dout(new_Jinkela_wire_14079)
    );

    bfr new_Jinkela_buffer_4630 (
        .din(new_Jinkela_wire_6041),
        .dout(new_Jinkela_wire_6042)
    );

    bfr new_Jinkela_buffer_11563 (
        .din(new_Jinkela_wire_13910),
        .dout(new_Jinkela_wire_13911)
    );

    bfr new_Jinkela_buffer_4696 (
        .din(new_Jinkela_wire_6109),
        .dout(new_Jinkela_wire_6110)
    );

    bfr new_Jinkela_buffer_11639 (
        .din(new_Jinkela_wire_14040),
        .dout(new_Jinkela_wire_14041)
    );

    bfr new_Jinkela_buffer_4631 (
        .din(new_Jinkela_wire_6042),
        .dout(new_Jinkela_wire_6043)
    );

    bfr new_Jinkela_buffer_11564 (
        .din(new_Jinkela_wire_13911),
        .dout(new_Jinkela_wire_13912)
    );

    bfr new_Jinkela_buffer_4814 (
        .din(new_Jinkela_wire_6243),
        .dout(new_Jinkela_wire_6244)
    );

    bfr new_Jinkela_buffer_11643 (
        .din(new_Jinkela_wire_14044),
        .dout(new_Jinkela_wire_14045)
    );

    bfr new_Jinkela_buffer_4632 (
        .din(new_Jinkela_wire_6043),
        .dout(new_Jinkela_wire_6044)
    );

    bfr new_Jinkela_buffer_11565 (
        .din(new_Jinkela_wire_13912),
        .dout(new_Jinkela_wire_13913)
    );

    bfr new_Jinkela_buffer_4697 (
        .din(new_Jinkela_wire_6110),
        .dout(new_Jinkela_wire_6111)
    );

    bfr new_Jinkela_buffer_11640 (
        .din(new_Jinkela_wire_14041),
        .dout(new_Jinkela_wire_14042)
    );

    bfr new_Jinkela_buffer_4633 (
        .din(new_Jinkela_wire_6044),
        .dout(new_Jinkela_wire_6045)
    );

    bfr new_Jinkela_buffer_11566 (
        .din(new_Jinkela_wire_13913),
        .dout(new_Jinkela_wire_13914)
    );

    bfr new_Jinkela_buffer_4785 (
        .din(new_Jinkela_wire_6208),
        .dout(new_Jinkela_wire_6209)
    );

    bfr new_Jinkela_buffer_11679 (
        .din(_1388_),
        .dout(new_Jinkela_wire_14085)
    );

    bfr new_Jinkela_buffer_11680 (
        .din(_0809_),
        .dout(new_Jinkela_wire_14088)
    );

    bfr new_Jinkela_buffer_4634 (
        .din(new_Jinkela_wire_6045),
        .dout(new_Jinkela_wire_6046)
    );

    bfr new_Jinkela_buffer_11567 (
        .din(new_Jinkela_wire_13914),
        .dout(new_Jinkela_wire_13915)
    );

    bfr new_Jinkela_buffer_4698 (
        .din(new_Jinkela_wire_6111),
        .dout(new_Jinkela_wire_6112)
    );

    bfr new_Jinkela_buffer_11641 (
        .din(new_Jinkela_wire_14042),
        .dout(new_Jinkela_wire_14043)
    );

    bfr new_Jinkela_buffer_4635 (
        .din(new_Jinkela_wire_6046),
        .dout(new_Jinkela_wire_6047)
    );

    bfr new_Jinkela_buffer_11568 (
        .din(new_Jinkela_wire_13915),
        .dout(new_Jinkela_wire_13916)
    );

    bfr new_Jinkela_buffer_11644 (
        .din(new_Jinkela_wire_14045),
        .dout(new_Jinkela_wire_14046)
    );

    bfr new_Jinkela_buffer_4822 (
        .din(new_net_3956),
        .dout(new_Jinkela_wire_6254)
    );

    bfr new_Jinkela_buffer_4636 (
        .din(new_Jinkela_wire_6047),
        .dout(new_Jinkela_wire_6048)
    );

    bfr new_Jinkela_buffer_11569 (
        .din(new_Jinkela_wire_13916),
        .dout(new_Jinkela_wire_13917)
    );

    bfr new_Jinkela_buffer_4699 (
        .din(new_Jinkela_wire_6112),
        .dout(new_Jinkela_wire_6113)
    );

    spl2 new_Jinkela_splitter_1052 (
        .a(_0606_),
        .b(new_Jinkela_wire_14086),
        .c(new_Jinkela_wire_14087)
    );

    bfr new_Jinkela_buffer_4637 (
        .din(new_Jinkela_wire_6048),
        .dout(new_Jinkela_wire_6049)
    );

    bfr new_Jinkela_buffer_11570 (
        .din(new_Jinkela_wire_13917),
        .dout(new_Jinkela_wire_13918)
    );

    bfr new_Jinkela_buffer_4786 (
        .din(new_Jinkela_wire_6209),
        .dout(new_Jinkela_wire_6210)
    );

    bfr new_Jinkela_buffer_11645 (
        .din(new_Jinkela_wire_14046),
        .dout(new_Jinkela_wire_14047)
    );

    bfr new_Jinkela_buffer_4638 (
        .din(new_Jinkela_wire_6049),
        .dout(new_Jinkela_wire_6050)
    );

    bfr new_Jinkela_buffer_11571 (
        .din(new_Jinkela_wire_13918),
        .dout(new_Jinkela_wire_13919)
    );

    bfr new_Jinkela_buffer_4700 (
        .din(new_Jinkela_wire_6113),
        .dout(new_Jinkela_wire_6114)
    );

    bfr new_Jinkela_buffer_11676 (
        .din(new_Jinkela_wire_14079),
        .dout(new_Jinkela_wire_14080)
    );

    bfr new_Jinkela_buffer_4639 (
        .din(new_Jinkela_wire_6050),
        .dout(new_Jinkela_wire_6051)
    );

    bfr new_Jinkela_buffer_11572 (
        .din(new_Jinkela_wire_13919),
        .dout(new_Jinkela_wire_13920)
    );

    bfr new_Jinkela_buffer_11646 (
        .din(new_Jinkela_wire_14047),
        .dout(new_Jinkela_wire_14048)
    );

    bfr new_Jinkela_buffer_4640 (
        .din(new_Jinkela_wire_6051),
        .dout(new_Jinkela_wire_6052)
    );

    bfr new_Jinkela_buffer_11573 (
        .din(new_Jinkela_wire_13920),
        .dout(new_Jinkela_wire_13921)
    );

    bfr new_Jinkela_buffer_4701 (
        .din(new_Jinkela_wire_6114),
        .dout(new_Jinkela_wire_6115)
    );

    bfr new_Jinkela_buffer_4641 (
        .din(new_Jinkela_wire_6052),
        .dout(new_Jinkela_wire_6053)
    );

    bfr new_Jinkela_buffer_11574 (
        .din(new_Jinkela_wire_13921),
        .dout(new_Jinkela_wire_13922)
    );

    bfr new_Jinkela_buffer_4787 (
        .din(new_Jinkela_wire_6210),
        .dout(new_Jinkela_wire_6211)
    );

    bfr new_Jinkela_buffer_11647 (
        .din(new_Jinkela_wire_14048),
        .dout(new_Jinkela_wire_14049)
    );

    bfr new_Jinkela_buffer_4642 (
        .din(new_Jinkela_wire_6053),
        .dout(new_Jinkela_wire_6054)
    );

    bfr new_Jinkela_buffer_11575 (
        .din(new_Jinkela_wire_13922),
        .dout(new_Jinkela_wire_13923)
    );

    bfr new_Jinkela_buffer_4702 (
        .din(new_Jinkela_wire_6115),
        .dout(new_Jinkela_wire_6116)
    );

    bfr new_Jinkela_buffer_11677 (
        .din(new_Jinkela_wire_14080),
        .dout(new_Jinkela_wire_14081)
    );

    bfr new_Jinkela_buffer_4643 (
        .din(new_Jinkela_wire_6054),
        .dout(new_Jinkela_wire_6055)
    );

    bfr new_Jinkela_buffer_11576 (
        .din(new_Jinkela_wire_13923),
        .dout(new_Jinkela_wire_13924)
    );

    bfr new_Jinkela_buffer_4815 (
        .din(new_Jinkela_wire_6244),
        .dout(new_Jinkela_wire_6245)
    );

    bfr new_Jinkela_buffer_11648 (
        .din(new_Jinkela_wire_14049),
        .dout(new_Jinkela_wire_14050)
    );

    bfr new_Jinkela_buffer_4644 (
        .din(new_Jinkela_wire_6055),
        .dout(new_Jinkela_wire_6056)
    );

    bfr new_Jinkela_buffer_11577 (
        .din(new_Jinkela_wire_13924),
        .dout(new_Jinkela_wire_13925)
    );

    bfr new_Jinkela_buffer_4703 (
        .din(new_Jinkela_wire_6116),
        .dout(new_Jinkela_wire_6117)
    );

    spl2 new_Jinkela_splitter_1053 (
        .a(_1778_),
        .b(new_Jinkela_wire_14090),
        .c(new_Jinkela_wire_14091)
    );

    bfr new_Jinkela_buffer_4645 (
        .din(new_Jinkela_wire_6056),
        .dout(new_Jinkela_wire_6057)
    );

    bfr new_Jinkela_buffer_11578 (
        .din(new_Jinkela_wire_13925),
        .dout(new_Jinkela_wire_13926)
    );

    bfr new_Jinkela_buffer_4788 (
        .din(new_Jinkela_wire_6211),
        .dout(new_Jinkela_wire_6212)
    );

    bfr new_Jinkela_buffer_11649 (
        .din(new_Jinkela_wire_14050),
        .dout(new_Jinkela_wire_14051)
    );

    bfr new_Jinkela_buffer_4646 (
        .din(new_Jinkela_wire_6057),
        .dout(new_Jinkela_wire_6058)
    );

    bfr new_Jinkela_buffer_11579 (
        .din(new_Jinkela_wire_13926),
        .dout(new_Jinkela_wire_13927)
    );

    bfr new_Jinkela_buffer_4704 (
        .din(new_Jinkela_wire_6117),
        .dout(new_Jinkela_wire_6118)
    );

    bfr new_Jinkela_buffer_11678 (
        .din(new_Jinkela_wire_14081),
        .dout(new_Jinkela_wire_14082)
    );

    bfr new_Jinkela_buffer_4647 (
        .din(new_Jinkela_wire_6058),
        .dout(new_Jinkela_wire_6059)
    );

    bfr new_Jinkela_buffer_11580 (
        .din(new_Jinkela_wire_13927),
        .dout(new_Jinkela_wire_13928)
    );

    bfr new_Jinkela_buffer_4818 (
        .din(new_Jinkela_wire_6249),
        .dout(new_Jinkela_wire_6250)
    );

    bfr new_Jinkela_buffer_11650 (
        .din(new_Jinkela_wire_14051),
        .dout(new_Jinkela_wire_14052)
    );

    bfr new_Jinkela_buffer_4930 (
        .din(_0209_),
        .dout(new_Jinkela_wire_6362)
    );

    bfr new_Jinkela_buffer_4648 (
        .din(new_Jinkela_wire_6059),
        .dout(new_Jinkela_wire_6060)
    );

    bfr new_Jinkela_buffer_11581 (
        .din(new_Jinkela_wire_13928),
        .dout(new_Jinkela_wire_13929)
    );

    bfr new_Jinkela_buffer_4705 (
        .din(new_Jinkela_wire_6118),
        .dout(new_Jinkela_wire_6119)
    );

    bfr new_Jinkela_buffer_4649 (
        .din(new_Jinkela_wire_6060),
        .dout(new_Jinkela_wire_6061)
    );

    bfr new_Jinkela_buffer_11582 (
        .din(new_Jinkela_wire_13929),
        .dout(new_Jinkela_wire_13930)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_1930),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1858),
        .dout(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_2024),
        .dout(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(new_Jinkela_wire_1859),
        .dout(new_Jinkela_wire_1860)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_1931),
        .dout(new_Jinkela_wire_1932)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(new_Jinkela_wire_1860),
        .dout(new_Jinkela_wire_1861)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(new_Jinkela_wire_2130),
        .dout(new_Jinkela_wire_2131)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(new_Jinkela_wire_1861),
        .dout(new_Jinkela_wire_1862)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_1932),
        .dout(new_Jinkela_wire_1933)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1862),
        .dout(new_Jinkela_wire_1863)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_2025),
        .dout(new_Jinkela_wire_2026)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(new_Jinkela_wire_1863),
        .dout(new_Jinkela_wire_1864)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(new_Jinkela_wire_1933),
        .dout(new_Jinkela_wire_1934)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1864),
        .dout(new_Jinkela_wire_1865)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(new_Jinkela_wire_1865),
        .dout(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(_0936_),
        .dout(new_Jinkela_wire_2128)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_1934),
        .dout(new_Jinkela_wire_1935)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1866),
        .dout(new_Jinkela_wire_1867)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1867),
        .dout(new_Jinkela_wire_1868)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_1935),
        .dout(new_Jinkela_wire_1936)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_Jinkela_wire_1868),
        .dout(new_Jinkela_wire_1869)
    );

    spl2 new_Jinkela_splitter_269 (
        .a(_0262_),
        .b(new_Jinkela_wire_2135),
        .c(new_Jinkela_wire_2136)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(new_Jinkela_wire_1869),
        .dout(new_Jinkela_wire_1870)
    );

    spl2 new_Jinkela_splitter_268 (
        .a(_0378_),
        .b(new_Jinkela_wire_2129),
        .c(new_Jinkela_wire_2130)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_1936),
        .dout(new_Jinkela_wire_1937)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1870),
        .dout(new_Jinkela_wire_1871)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(new_Jinkela_wire_2027),
        .dout(new_Jinkela_wire_2028)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1871),
        .dout(new_Jinkela_wire_1872)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_1937),
        .dout(new_Jinkela_wire_1938)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_Jinkela_wire_1872),
        .dout(new_Jinkela_wire_1873)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1873),
        .dout(new_Jinkela_wire_1874)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_1938),
        .dout(new_Jinkela_wire_1939)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1874),
        .dout(new_Jinkela_wire_1875)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_2028),
        .dout(new_Jinkela_wire_2029)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1875),
        .dout(new_Jinkela_wire_1876)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_1939),
        .dout(new_Jinkela_wire_1940)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1876),
        .dout(new_Jinkela_wire_1877)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1877),
        .dout(new_Jinkela_wire_1878)
    );

    spl2 new_Jinkela_splitter_270 (
        .a(_0259_),
        .b(new_Jinkela_wire_2137),
        .c(new_Jinkela_wire_2138)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_1940),
        .dout(new_Jinkela_wire_1941)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(new_Jinkela_wire_1878),
        .dout(new_Jinkela_wire_1879)
    );

    bfr new_Jinkela_buffer_8094 (
        .din(new_Jinkela_wire_9975),
        .dout(new_Jinkela_wire_9976)
    );

    spl2 new_Jinkela_splitter_815 (
        .a(_0513_),
        .b(new_Jinkela_wire_10259),
        .c(new_Jinkela_wire_10260)
    );

    bfr new_Jinkela_buffer_8206 (
        .din(new_Jinkela_wire_10127),
        .dout(new_Jinkela_wire_10128)
    );

    bfr new_Jinkela_buffer_8095 (
        .din(new_Jinkela_wire_9976),
        .dout(new_Jinkela_wire_9977)
    );

    bfr new_Jinkela_buffer_8242 (
        .din(new_Jinkela_wire_10165),
        .dout(new_Jinkela_wire_10166)
    );

    bfr new_Jinkela_buffer_8096 (
        .din(new_Jinkela_wire_9977),
        .dout(new_Jinkela_wire_9978)
    );

    bfr new_Jinkela_buffer_8207 (
        .din(new_Jinkela_wire_10128),
        .dout(new_Jinkela_wire_10129)
    );

    bfr new_Jinkela_buffer_8097 (
        .din(new_Jinkela_wire_9978),
        .dout(new_Jinkela_wire_9979)
    );

    bfr new_Jinkela_buffer_8280 (
        .din(new_Jinkela_wire_10207),
        .dout(new_Jinkela_wire_10208)
    );

    bfr new_Jinkela_buffer_8098 (
        .din(new_Jinkela_wire_9979),
        .dout(new_Jinkela_wire_9980)
    );

    bfr new_Jinkela_buffer_8208 (
        .din(new_Jinkela_wire_10129),
        .dout(new_Jinkela_wire_10130)
    );

    bfr new_Jinkela_buffer_8099 (
        .din(new_Jinkela_wire_9980),
        .dout(new_Jinkela_wire_9981)
    );

    bfr new_Jinkela_buffer_8243 (
        .din(new_Jinkela_wire_10166),
        .dout(new_Jinkela_wire_10167)
    );

    bfr new_Jinkela_buffer_8100 (
        .din(new_Jinkela_wire_9981),
        .dout(new_Jinkela_wire_9982)
    );

    bfr new_Jinkela_buffer_8209 (
        .din(new_Jinkela_wire_10130),
        .dout(new_Jinkela_wire_10131)
    );

    bfr new_Jinkela_buffer_8101 (
        .din(new_Jinkela_wire_9982),
        .dout(new_Jinkela_wire_9983)
    );

    and_ii _1863_ (
        .a(new_Jinkela_wire_5106),
        .b(new_Jinkela_wire_8863),
        .c(_1730_)
    );

    bfr new_Jinkela_buffer_8102 (
        .din(new_Jinkela_wire_9983),
        .dout(new_Jinkela_wire_9984)
    );

    and_bi _1841_ (
        .a(new_Jinkela_wire_5428),
        .b(new_Jinkela_wire_13396),
        .c(_1491_)
    );

    and_bb _1839_ (
        .a(new_Jinkela_wire_98),
        .b(new_Jinkela_wire_225),
        .c(_1469_)
    );

    bfr new_Jinkela_buffer_8210 (
        .din(new_Jinkela_wire_10131),
        .dout(new_Jinkela_wire_10132)
    );

    or_ii _1840_ (
        .a(new_Jinkela_wire_328),
        .b(new_Jinkela_wire_555),
        .c(_1480_)
    );

    bfr new_Jinkela_buffer_8103 (
        .din(new_Jinkela_wire_9984),
        .dout(new_Jinkela_wire_9985)
    );

    and_bb _1838_ (
        .a(new_Jinkela_wire_630),
        .b(new_Jinkela_wire_337),
        .c(_1458_)
    );

    and_bb _1842_ (
        .a(new_Jinkela_wire_224),
        .b(new_Jinkela_wire_568),
        .c(_1502_)
    );

    bfr new_Jinkela_buffer_8244 (
        .din(new_Jinkela_wire_10167),
        .dout(new_Jinkela_wire_10168)
    );

    bfr new_Jinkela_buffer_8104 (
        .din(new_Jinkela_wire_9985),
        .dout(new_Jinkela_wire_9986)
    );

    and_bb _1846_ (
        .a(new_Jinkela_wire_239),
        .b(new_Jinkela_wire_340),
        .c(new_net_0)
    );

    and_ii _1845_ (
        .a(new_Jinkela_wire_2597),
        .b(new_Jinkela_wire_7729),
        .c(_1535_)
    );

    bfr new_Jinkela_buffer_8211 (
        .din(new_Jinkela_wire_10132),
        .dout(new_Jinkela_wire_10133)
    );

    bfr new_Jinkela_buffer_8105 (
        .din(new_Jinkela_wire_9986),
        .dout(new_Jinkela_wire_9987)
    );

    or_ii _1843_ (
        .a(new_Jinkela_wire_89),
        .b(new_Jinkela_wire_322),
        .c(_1513_)
    );

    bfr new_Jinkela_buffer_8281 (
        .din(new_Jinkela_wire_10208),
        .dout(new_Jinkela_wire_10209)
    );

    or_ii _1855_ (
        .a(new_Jinkela_wire_267),
        .b(new_Jinkela_wire_316),
        .c(_1643_)
    );

    bfr new_Jinkela_buffer_8106 (
        .din(new_Jinkela_wire_9987),
        .dout(new_Jinkela_wire_9988)
    );

    and_bi _1844_ (
        .a(new_Jinkela_wire_20360),
        .b(new_Jinkela_wire_14284),
        .c(_1524_)
    );

    or_bi _1847_ (
        .a(new_Jinkela_wire_20361),
        .b(new_Jinkela_wire_12343),
        .c(_1556_)
    );

    bfr new_Jinkela_buffer_8212 (
        .din(new_Jinkela_wire_10133),
        .dout(new_Jinkela_wire_10134)
    );

    or_bi _1848_ (
        .a(new_Jinkela_wire_20346),
        .b(new_Jinkela_wire_16109),
        .c(_1566_)
    );

    bfr new_Jinkela_buffer_8107 (
        .din(new_Jinkela_wire_9988),
        .dout(new_Jinkela_wire_9989)
    );

    and_bb _1849_ (
        .a(new_Jinkela_wire_539),
        .b(new_Jinkela_wire_350),
        .c(_1577_)
    );

    bfr new_Jinkela_buffer_8245 (
        .din(new_Jinkela_wire_10168),
        .dout(new_Jinkela_wire_10169)
    );

    and_bi _1850_ (
        .a(new_Jinkela_wire_20347),
        .b(new_Jinkela_wire_16110),
        .c(_1588_)
    );

    bfr new_Jinkela_buffer_8108 (
        .din(new_Jinkela_wire_9989),
        .dout(new_Jinkela_wire_9990)
    );

    or_bi _1851_ (
        .a(new_Jinkela_wire_6009),
        .b(new_Jinkela_wire_21326),
        .c(_1599_)
    );

    bfr new_Jinkela_buffer_8213 (
        .din(new_Jinkela_wire_10134),
        .dout(new_Jinkela_wire_10135)
    );

    and_ii _1852_ (
        .a(new_Jinkela_wire_4905),
        .b(new_Jinkela_wire_18307),
        .c(_1610_)
    );

    bfr new_Jinkela_buffer_8109 (
        .din(new_Jinkela_wire_9990),
        .dout(new_Jinkela_wire_9991)
    );

    and_bi _1853_ (
        .a(new_Jinkela_wire_21331),
        .b(new_Jinkela_wire_5542),
        .c(_1621_)
    );

    spl2 new_Jinkela_splitter_817 (
        .a(_0729_),
        .b(new_Jinkela_wire_10263),
        .c(new_Jinkela_wire_10264)
    );

    and_bb _1854_ (
        .a(new_Jinkela_wire_106),
        .b(new_Jinkela_wire_534),
        .c(_1632_)
    );

    bfr new_Jinkela_buffer_8110 (
        .din(new_Jinkela_wire_9991),
        .dout(new_Jinkela_wire_9992)
    );

    spl2 new_Jinkela_splitter_816 (
        .a(_0269_),
        .b(new_Jinkela_wire_10261),
        .c(new_Jinkela_wire_10262)
    );

    and_bi _1856_ (
        .a(new_Jinkela_wire_14285),
        .b(new_Jinkela_wire_4713),
        .c(_1654_)
    );

    bfr new_Jinkela_buffer_8214 (
        .din(new_Jinkela_wire_10135),
        .dout(new_Jinkela_wire_10136)
    );

    bfr new_Jinkela_buffer_8111 (
        .din(new_Jinkela_wire_9992),
        .dout(new_Jinkela_wire_9993)
    );

    and_bb _1857_ (
        .a(new_Jinkela_wire_277),
        .b(new_Jinkela_wire_233),
        .c(_1665_)
    );

    and_bi _1858_ (
        .a(new_Jinkela_wire_13397),
        .b(new_Jinkela_wire_5737),
        .c(_1676_)
    );

    bfr new_Jinkela_buffer_8246 (
        .din(new_Jinkela_wire_10169),
        .dout(new_Jinkela_wire_10170)
    );

    bfr new_Jinkela_buffer_8112 (
        .din(new_Jinkela_wire_9993),
        .dout(new_Jinkela_wire_9994)
    );

    and_ii _1859_ (
        .a(new_Jinkela_wire_4240),
        .b(new_Jinkela_wire_6763),
        .c(_1686_)
    );

    or_bb _1860_ (
        .a(new_Jinkela_wire_703),
        .b(new_Jinkela_wire_7733),
        .c(_1697_)
    );

    bfr new_Jinkela_buffer_8215 (
        .din(new_Jinkela_wire_10136),
        .dout(new_Jinkela_wire_10137)
    );

    bfr new_Jinkela_buffer_8113 (
        .din(new_Jinkela_wire_9994),
        .dout(new_Jinkela_wire_9995)
    );

    or_ii _1861_ (
        .a(new_Jinkela_wire_704),
        .b(new_Jinkela_wire_7732),
        .c(_1708_)
    );

    or_ii _1862_ (
        .a(new_Jinkela_wire_18445),
        .b(new_Jinkela_wire_5151),
        .c(_1719_)
    );

    bfr new_Jinkela_buffer_8282 (
        .din(new_Jinkela_wire_10209),
        .dout(new_Jinkela_wire_10210)
    );

    bfr new_Jinkela_buffer_8114 (
        .din(new_Jinkela_wire_9995),
        .dout(new_Jinkela_wire_9996)
    );

    bfr new_Jinkela_buffer_4789 (
        .din(new_Jinkela_wire_6212),
        .dout(new_Jinkela_wire_6213)
    );

    bfr new_Jinkela_buffer_11651 (
        .din(new_Jinkela_wire_14052),
        .dout(new_Jinkela_wire_14053)
    );

    bfr new_Jinkela_buffer_15052 (
        .din(new_Jinkela_wire_17950),
        .dout(new_Jinkela_wire_17951)
    );

    bfr new_Jinkela_buffer_4650 (
        .din(new_Jinkela_wire_6061),
        .dout(new_Jinkela_wire_6062)
    );

    bfr new_Jinkela_buffer_11583 (
        .din(new_Jinkela_wire_13930),
        .dout(new_Jinkela_wire_13931)
    );

    bfr new_Jinkela_buffer_15087 (
        .din(new_Jinkela_wire_18007),
        .dout(new_Jinkela_wire_18008)
    );

    bfr new_Jinkela_buffer_4706 (
        .din(new_Jinkela_wire_6119),
        .dout(new_Jinkela_wire_6120)
    );

    spl2 new_Jinkela_splitter_1051 (
        .a(new_Jinkela_wire_14082),
        .b(new_Jinkela_wire_14083),
        .c(new_Jinkela_wire_14084)
    );

    bfr new_Jinkela_buffer_15053 (
        .din(new_Jinkela_wire_17951),
        .dout(new_Jinkela_wire_17952)
    );

    bfr new_Jinkela_buffer_4651 (
        .din(new_Jinkela_wire_6062),
        .dout(new_Jinkela_wire_6063)
    );

    bfr new_Jinkela_buffer_11584 (
        .din(new_Jinkela_wire_13931),
        .dout(new_Jinkela_wire_13932)
    );

    bfr new_Jinkela_buffer_15189 (
        .din(_0701_),
        .dout(new_Jinkela_wire_18124)
    );

    bfr new_Jinkela_buffer_4816 (
        .din(new_Jinkela_wire_6245),
        .dout(new_Jinkela_wire_6246)
    );

    bfr new_Jinkela_buffer_11652 (
        .din(new_Jinkela_wire_14053),
        .dout(new_Jinkela_wire_14054)
    );

    bfr new_Jinkela_buffer_15054 (
        .din(new_Jinkela_wire_17952),
        .dout(new_Jinkela_wire_17953)
    );

    bfr new_Jinkela_buffer_4652 (
        .din(new_Jinkela_wire_6063),
        .dout(new_Jinkela_wire_6064)
    );

    bfr new_Jinkela_buffer_11585 (
        .din(new_Jinkela_wire_13932),
        .dout(new_Jinkela_wire_13933)
    );

    bfr new_Jinkela_buffer_15088 (
        .din(new_Jinkela_wire_18008),
        .dout(new_Jinkela_wire_18009)
    );

    bfr new_Jinkela_buffer_4707 (
        .din(new_Jinkela_wire_6120),
        .dout(new_Jinkela_wire_6121)
    );

    bfr new_Jinkela_buffer_15055 (
        .din(new_Jinkela_wire_17953),
        .dout(new_Jinkela_wire_17954)
    );

    bfr new_Jinkela_buffer_4653 (
        .din(new_Jinkela_wire_6064),
        .dout(new_Jinkela_wire_6065)
    );

    bfr new_Jinkela_buffer_11586 (
        .din(new_Jinkela_wire_13933),
        .dout(new_Jinkela_wire_13934)
    );

    bfr new_Jinkela_buffer_15186 (
        .din(new_Jinkela_wire_18114),
        .dout(new_Jinkela_wire_18115)
    );

    bfr new_Jinkela_buffer_4790 (
        .din(new_Jinkela_wire_6213),
        .dout(new_Jinkela_wire_6214)
    );

    bfr new_Jinkela_buffer_11653 (
        .din(new_Jinkela_wire_14054),
        .dout(new_Jinkela_wire_14055)
    );

    bfr new_Jinkela_buffer_15056 (
        .din(new_Jinkela_wire_17954),
        .dout(new_Jinkela_wire_17955)
    );

    bfr new_Jinkela_buffer_4654 (
        .din(new_Jinkela_wire_6065),
        .dout(new_Jinkela_wire_6066)
    );

    bfr new_Jinkela_buffer_11587 (
        .din(new_Jinkela_wire_13934),
        .dout(new_Jinkela_wire_13935)
    );

    bfr new_Jinkela_buffer_15089 (
        .din(new_Jinkela_wire_18009),
        .dout(new_Jinkela_wire_18010)
    );

    bfr new_Jinkela_buffer_4708 (
        .din(new_Jinkela_wire_6121),
        .dout(new_Jinkela_wire_6122)
    );

    spl2 new_Jinkela_splitter_1054 (
        .a(_0449_),
        .b(new_Jinkela_wire_14096),
        .c(new_Jinkela_wire_14097)
    );

    bfr new_Jinkela_buffer_15057 (
        .din(new_Jinkela_wire_17955),
        .dout(new_Jinkela_wire_17956)
    );

    bfr new_Jinkela_buffer_11682 (
        .din(new_Jinkela_wire_14091),
        .dout(new_Jinkela_wire_14092)
    );

    bfr new_Jinkela_buffer_4655 (
        .din(new_Jinkela_wire_6066),
        .dout(new_Jinkela_wire_6067)
    );

    bfr new_Jinkela_buffer_11588 (
        .din(new_Jinkela_wire_13935),
        .dout(new_Jinkela_wire_13936)
    );

    spl2 new_Jinkela_splitter_1315 (
        .a(_1608_),
        .b(new_Jinkela_wire_18122),
        .c(new_Jinkela_wire_18123)
    );

    bfr new_Jinkela_buffer_11654 (
        .din(new_Jinkela_wire_14055),
        .dout(new_Jinkela_wire_14056)
    );

    bfr new_Jinkela_buffer_15058 (
        .din(new_Jinkela_wire_17956),
        .dout(new_Jinkela_wire_17957)
    );

    bfr new_Jinkela_buffer_4823 (
        .din(new_Jinkela_wire_6254),
        .dout(new_Jinkela_wire_6255)
    );

    bfr new_Jinkela_buffer_4656 (
        .din(new_Jinkela_wire_6067),
        .dout(new_Jinkela_wire_6068)
    );

    bfr new_Jinkela_buffer_11589 (
        .din(new_Jinkela_wire_13936),
        .dout(new_Jinkela_wire_13937)
    );

    bfr new_Jinkela_buffer_15090 (
        .din(new_Jinkela_wire_18010),
        .dout(new_Jinkela_wire_18011)
    );

    bfr new_Jinkela_buffer_4709 (
        .din(new_Jinkela_wire_6122),
        .dout(new_Jinkela_wire_6123)
    );

    bfr new_Jinkela_buffer_15059 (
        .din(new_Jinkela_wire_17957),
        .dout(new_Jinkela_wire_17958)
    );

    spl2 new_Jinkela_splitter_1055 (
        .a(_1655_),
        .b(new_Jinkela_wire_14098),
        .c(new_Jinkela_wire_14099)
    );

    bfr new_Jinkela_buffer_4657 (
        .din(new_Jinkela_wire_6068),
        .dout(new_Jinkela_wire_6069)
    );

    bfr new_Jinkela_buffer_11590 (
        .din(new_Jinkela_wire_13937),
        .dout(new_Jinkela_wire_13938)
    );

    bfr new_Jinkela_buffer_15187 (
        .din(new_Jinkela_wire_18115),
        .dout(new_Jinkela_wire_18116)
    );

    bfr new_Jinkela_buffer_4791 (
        .din(new_Jinkela_wire_6214),
        .dout(new_Jinkela_wire_6215)
    );

    bfr new_Jinkela_buffer_11655 (
        .din(new_Jinkela_wire_14056),
        .dout(new_Jinkela_wire_14057)
    );

    bfr new_Jinkela_buffer_15060 (
        .din(new_Jinkela_wire_17958),
        .dout(new_Jinkela_wire_17959)
    );

    bfr new_Jinkela_buffer_4658 (
        .din(new_Jinkela_wire_6069),
        .dout(new_Jinkela_wire_6070)
    );

    bfr new_Jinkela_buffer_11591 (
        .din(new_Jinkela_wire_13938),
        .dout(new_Jinkela_wire_13939)
    );

    bfr new_Jinkela_buffer_15091 (
        .din(new_Jinkela_wire_18011),
        .dout(new_Jinkela_wire_18012)
    );

    bfr new_Jinkela_buffer_4710 (
        .din(new_Jinkela_wire_6123),
        .dout(new_Jinkela_wire_6124)
    );

    bfr new_Jinkela_buffer_15061 (
        .din(new_Jinkela_wire_17959),
        .dout(new_Jinkela_wire_17960)
    );

    bfr new_Jinkela_buffer_4659 (
        .din(new_Jinkela_wire_6070),
        .dout(new_Jinkela_wire_6071)
    );

    bfr new_Jinkela_buffer_11592 (
        .din(new_Jinkela_wire_13939),
        .dout(new_Jinkela_wire_13940)
    );

    spl2 new_Jinkela_splitter_1317 (
        .a(_0741_),
        .b(new_Jinkela_wire_18223),
        .c(new_Jinkela_wire_18224)
    );

    bfr new_Jinkela_buffer_4817 (
        .din(new_Jinkela_wire_6246),
        .dout(new_Jinkela_wire_6247)
    );

    bfr new_Jinkela_buffer_11656 (
        .din(new_Jinkela_wire_14057),
        .dout(new_Jinkela_wire_14058)
    );

    bfr new_Jinkela_buffer_15062 (
        .din(new_Jinkela_wire_17960),
        .dout(new_Jinkela_wire_17961)
    );

    bfr new_Jinkela_buffer_4660 (
        .din(new_Jinkela_wire_6071),
        .dout(new_Jinkela_wire_6072)
    );

    bfr new_Jinkela_buffer_11593 (
        .din(new_Jinkela_wire_13940),
        .dout(new_Jinkela_wire_13941)
    );

    bfr new_Jinkela_buffer_15092 (
        .din(new_Jinkela_wire_18012),
        .dout(new_Jinkela_wire_18013)
    );

    bfr new_Jinkela_buffer_4711 (
        .din(new_Jinkela_wire_6124),
        .dout(new_Jinkela_wire_6125)
    );

    bfr new_Jinkela_buffer_11683 (
        .din(new_Jinkela_wire_14092),
        .dout(new_Jinkela_wire_14093)
    );

    bfr new_Jinkela_buffer_15063 (
        .din(new_Jinkela_wire_17961),
        .dout(new_Jinkela_wire_17962)
    );

    bfr new_Jinkela_buffer_4661 (
        .din(new_Jinkela_wire_6072),
        .dout(new_Jinkela_wire_6073)
    );

    bfr new_Jinkela_buffer_11594 (
        .din(new_Jinkela_wire_13941),
        .dout(new_Jinkela_wire_13942)
    );

    bfr new_Jinkela_buffer_15285 (
        .din(_0906_),
        .dout(new_Jinkela_wire_18222)
    );

    bfr new_Jinkela_buffer_4792 (
        .din(new_Jinkela_wire_6215),
        .dout(new_Jinkela_wire_6216)
    );

    bfr new_Jinkela_buffer_11657 (
        .din(new_Jinkela_wire_14058),
        .dout(new_Jinkela_wire_14059)
    );

    bfr new_Jinkela_buffer_15064 (
        .din(new_Jinkela_wire_17962),
        .dout(new_Jinkela_wire_17963)
    );

    bfr new_Jinkela_buffer_4662 (
        .din(new_Jinkela_wire_6073),
        .dout(new_Jinkela_wire_6074)
    );

    bfr new_Jinkela_buffer_11595 (
        .din(new_Jinkela_wire_13942),
        .dout(new_Jinkela_wire_13943)
    );

    bfr new_Jinkela_buffer_15093 (
        .din(new_Jinkela_wire_18013),
        .dout(new_Jinkela_wire_18014)
    );

    bfr new_Jinkela_buffer_4712 (
        .din(new_Jinkela_wire_6125),
        .dout(new_Jinkela_wire_6126)
    );

    bfr new_Jinkela_buffer_11688 (
        .din(_1811_),
        .dout(new_Jinkela_wire_14102)
    );

    bfr new_Jinkela_buffer_15065 (
        .din(new_Jinkela_wire_17963),
        .dout(new_Jinkela_wire_17964)
    );

    bfr new_Jinkela_buffer_11686 (
        .din(_0270_),
        .dout(new_Jinkela_wire_14100)
    );

    bfr new_Jinkela_buffer_4663 (
        .din(new_Jinkela_wire_6074),
        .dout(new_Jinkela_wire_6075)
    );

    bfr new_Jinkela_buffer_11596 (
        .din(new_Jinkela_wire_13943),
        .dout(new_Jinkela_wire_13944)
    );

    bfr new_Jinkela_buffer_15190 (
        .din(new_Jinkela_wire_18124),
        .dout(new_Jinkela_wire_18125)
    );

    bfr new_Jinkela_buffer_4819 (
        .din(new_Jinkela_wire_6250),
        .dout(new_Jinkela_wire_6251)
    );

    bfr new_Jinkela_buffer_11658 (
        .din(new_Jinkela_wire_14059),
        .dout(new_Jinkela_wire_14060)
    );

    bfr new_Jinkela_buffer_15066 (
        .din(new_Jinkela_wire_17964),
        .dout(new_Jinkela_wire_17965)
    );

    bfr new_Jinkela_buffer_4664 (
        .din(new_Jinkela_wire_6075),
        .dout(new_Jinkela_wire_6076)
    );

    bfr new_Jinkela_buffer_11597 (
        .din(new_Jinkela_wire_13944),
        .dout(new_Jinkela_wire_13945)
    );

    bfr new_Jinkela_buffer_15094 (
        .din(new_Jinkela_wire_18014),
        .dout(new_Jinkela_wire_18015)
    );

    bfr new_Jinkela_buffer_4713 (
        .din(new_Jinkela_wire_6126),
        .dout(new_Jinkela_wire_6127)
    );

    bfr new_Jinkela_buffer_11684 (
        .din(new_Jinkela_wire_14093),
        .dout(new_Jinkela_wire_14094)
    );

    bfr new_Jinkela_buffer_15067 (
        .din(new_Jinkela_wire_17965),
        .dout(new_Jinkela_wire_17966)
    );

    bfr new_Jinkela_buffer_4665 (
        .din(new_Jinkela_wire_6076),
        .dout(new_Jinkela_wire_6077)
    );

    bfr new_Jinkela_buffer_11598 (
        .din(new_Jinkela_wire_13945),
        .dout(new_Jinkela_wire_13946)
    );

    spl2 new_Jinkela_splitter_1318 (
        .a(_1050_),
        .b(new_Jinkela_wire_18225),
        .c(new_Jinkela_wire_18226)
    );

    bfr new_Jinkela_buffer_4793 (
        .din(new_Jinkela_wire_6216),
        .dout(new_Jinkela_wire_6217)
    );

    bfr new_Jinkela_buffer_11659 (
        .din(new_Jinkela_wire_14060),
        .dout(new_Jinkela_wire_14061)
    );

    bfr new_Jinkela_buffer_15068 (
        .din(new_Jinkela_wire_17966),
        .dout(new_Jinkela_wire_17967)
    );

    bfr new_Jinkela_buffer_4666 (
        .din(new_Jinkela_wire_6077),
        .dout(new_Jinkela_wire_6078)
    );

    bfr new_Jinkela_buffer_11599 (
        .din(new_Jinkela_wire_13946),
        .dout(new_Jinkela_wire_13947)
    );

    bfr new_Jinkela_buffer_15095 (
        .din(new_Jinkela_wire_18015),
        .dout(new_Jinkela_wire_18016)
    );

    bfr new_Jinkela_buffer_4714 (
        .din(new_Jinkela_wire_6127),
        .dout(new_Jinkela_wire_6128)
    );

    bfr new_Jinkela_buffer_15069 (
        .din(new_Jinkela_wire_17967),
        .dout(new_Jinkela_wire_17968)
    );

    bfr new_Jinkela_buffer_11687 (
        .din(_1107_),
        .dout(new_Jinkela_wire_14101)
    );

    bfr new_Jinkela_buffer_4667 (
        .din(new_Jinkela_wire_6078),
        .dout(new_Jinkela_wire_6079)
    );

    bfr new_Jinkela_buffer_11600 (
        .din(new_Jinkela_wire_13947),
        .dout(new_Jinkela_wire_13948)
    );

    bfr new_Jinkela_buffer_15191 (
        .din(new_Jinkela_wire_18125),
        .dout(new_Jinkela_wire_18126)
    );

    bfr new_Jinkela_buffer_11660 (
        .din(new_Jinkela_wire_14061),
        .dout(new_Jinkela_wire_14062)
    );

    bfr new_Jinkela_buffer_15070 (
        .din(new_Jinkela_wire_17968),
        .dout(new_Jinkela_wire_17969)
    );

    spl2 new_Jinkela_splitter_565 (
        .a(_1499_),
        .b(new_Jinkela_wire_6363),
        .c(new_Jinkela_wire_6364)
    );

    bfr new_Jinkela_buffer_4668 (
        .din(new_Jinkela_wire_6079),
        .dout(new_Jinkela_wire_6080)
    );

    bfr new_Jinkela_buffer_11601 (
        .din(new_Jinkela_wire_13948),
        .dout(new_Jinkela_wire_13949)
    );

    bfr new_Jinkela_buffer_15096 (
        .din(new_Jinkela_wire_18016),
        .dout(new_Jinkela_wire_18017)
    );

    bfr new_Jinkela_buffer_4715 (
        .din(new_Jinkela_wire_6128),
        .dout(new_Jinkela_wire_6129)
    );

    bfr new_Jinkela_buffer_11685 (
        .din(new_Jinkela_wire_14094),
        .dout(new_Jinkela_wire_14095)
    );

    bfr new_Jinkela_buffer_15071 (
        .din(new_Jinkela_wire_17969),
        .dout(new_Jinkela_wire_17970)
    );

    bfr new_Jinkela_buffer_4669 (
        .din(new_Jinkela_wire_6080),
        .dout(new_Jinkela_wire_6081)
    );

    bfr new_Jinkela_buffer_11602 (
        .din(new_Jinkela_wire_13949),
        .dout(new_Jinkela_wire_13950)
    );

    bfr new_Jinkela_buffer_15286 (
        .din(_0344_),
        .dout(new_Jinkela_wire_18227)
    );

    bfr new_Jinkela_buffer_4794 (
        .din(new_Jinkela_wire_6217),
        .dout(new_Jinkela_wire_6218)
    );

    bfr new_Jinkela_buffer_11661 (
        .din(new_Jinkela_wire_14062),
        .dout(new_Jinkela_wire_14063)
    );

    bfr new_Jinkela_buffer_15072 (
        .din(new_Jinkela_wire_17970),
        .dout(new_Jinkela_wire_17971)
    );

    bfr new_Jinkela_buffer_4670 (
        .din(new_Jinkela_wire_6081),
        .dout(new_Jinkela_wire_6082)
    );

    bfr new_Jinkela_buffer_11603 (
        .din(new_Jinkela_wire_13950),
        .dout(new_Jinkela_wire_13951)
    );

    bfr new_Jinkela_buffer_15097 (
        .din(new_Jinkela_wire_18017),
        .dout(new_Jinkela_wire_18018)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_2029),
        .dout(new_Jinkela_wire_2030)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1879),
        .dout(new_Jinkela_wire_1880)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(new_Jinkela_wire_1941),
        .dout(new_Jinkela_wire_1942)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1880),
        .dout(new_Jinkela_wire_1881)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1881),
        .dout(new_Jinkela_wire_1882)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(new_Jinkela_wire_1942),
        .dout(new_Jinkela_wire_1943)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_Jinkela_wire_1882),
        .dout(new_Jinkela_wire_1883)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(new_Jinkela_wire_2030),
        .dout(new_Jinkela_wire_2031)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1883),
        .dout(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(new_Jinkela_wire_1943),
        .dout(new_Jinkela_wire_1944)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_1884),
        .dout(new_Jinkela_wire_1885)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(new_Jinkela_wire_2131),
        .dout(new_Jinkela_wire_2132)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_1885),
        .dout(new_Jinkela_wire_1886)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_Jinkela_wire_1944),
        .dout(new_Jinkela_wire_1945)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_1886),
        .dout(new_Jinkela_wire_1887)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_2031),
        .dout(new_Jinkela_wire_2032)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(new_Jinkela_wire_1887),
        .dout(new_Jinkela_wire_1888)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_1945),
        .dout(new_Jinkela_wire_1946)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_Jinkela_wire_1888),
        .dout(new_Jinkela_wire_1889)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_1889),
        .dout(new_Jinkela_wire_1890)
    );

    spl2 new_Jinkela_splitter_271 (
        .a(_1662_),
        .b(new_Jinkela_wire_2143),
        .c(new_Jinkela_wire_2144)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_1946),
        .dout(new_Jinkela_wire_1947)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_1890),
        .dout(new_Jinkela_wire_1891)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(new_Jinkela_wire_2032),
        .dout(new_Jinkela_wire_2033)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_1891),
        .dout(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(new_Jinkela_wire_1947),
        .dout(new_Jinkela_wire_1948)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_1892),
        .dout(new_Jinkela_wire_1893)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(new_Jinkela_wire_2132),
        .dout(new_Jinkela_wire_2133)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_1893),
        .dout(new_Jinkela_wire_1894)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_1948),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_1894),
        .dout(new_Jinkela_wire_1895)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_2033),
        .dout(new_Jinkela_wire_2034)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_1949),
        .dout(new_Jinkela_wire_1950)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(new_Jinkela_wire_2138),
        .dout(new_Jinkela_wire_2139)
    );

    spl2 new_Jinkela_splitter_272 (
        .a(_1801_),
        .b(new_Jinkela_wire_2145),
        .c(new_Jinkela_wire_2146)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(new_Jinkela_wire_1950),
        .dout(new_Jinkela_wire_1951)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(new_Jinkela_wire_2034),
        .dout(new_Jinkela_wire_2035)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_1951),
        .dout(new_Jinkela_wire_1952)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_2133),
        .dout(new_Jinkela_wire_2134)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_1952),
        .dout(new_Jinkela_wire_1953)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_Jinkela_wire_2035),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_1953),
        .dout(new_Jinkela_wire_1954)
    );

    bfr new_Jinkela_buffer_8216 (
        .din(new_Jinkela_wire_10137),
        .dout(new_Jinkela_wire_10138)
    );

    bfr new_Jinkela_buffer_8115 (
        .din(new_Jinkela_wire_9996),
        .dout(new_Jinkela_wire_9997)
    );

    bfr new_Jinkela_buffer_8247 (
        .din(new_Jinkela_wire_10170),
        .dout(new_Jinkela_wire_10171)
    );

    bfr new_Jinkela_buffer_8116 (
        .din(new_Jinkela_wire_9997),
        .dout(new_Jinkela_wire_9998)
    );

    bfr new_Jinkela_buffer_8217 (
        .din(new_Jinkela_wire_10138),
        .dout(new_Jinkela_wire_10139)
    );

    bfr new_Jinkela_buffer_8117 (
        .din(new_Jinkela_wire_9998),
        .dout(new_Jinkela_wire_9999)
    );

    bfr new_Jinkela_buffer_8336 (
        .din(_1448_),
        .dout(new_Jinkela_wire_10276)
    );

    bfr new_Jinkela_buffer_8118 (
        .din(new_Jinkela_wire_9999),
        .dout(new_Jinkela_wire_10000)
    );

    bfr new_Jinkela_buffer_8218 (
        .din(new_Jinkela_wire_10139),
        .dout(new_Jinkela_wire_10140)
    );

    bfr new_Jinkela_buffer_8119 (
        .din(new_Jinkela_wire_10000),
        .dout(new_Jinkela_wire_10001)
    );

    bfr new_Jinkela_buffer_8248 (
        .din(new_Jinkela_wire_10171),
        .dout(new_Jinkela_wire_10172)
    );

    bfr new_Jinkela_buffer_8120 (
        .din(new_Jinkela_wire_10001),
        .dout(new_Jinkela_wire_10002)
    );

    bfr new_Jinkela_buffer_8219 (
        .din(new_Jinkela_wire_10140),
        .dout(new_Jinkela_wire_10141)
    );

    bfr new_Jinkela_buffer_8121 (
        .din(new_Jinkela_wire_10002),
        .dout(new_Jinkela_wire_10003)
    );

    bfr new_Jinkela_buffer_8283 (
        .din(new_Jinkela_wire_10210),
        .dout(new_Jinkela_wire_10211)
    );

    bfr new_Jinkela_buffer_8122 (
        .din(new_Jinkela_wire_10003),
        .dout(new_Jinkela_wire_10004)
    );

    bfr new_Jinkela_buffer_8220 (
        .din(new_Jinkela_wire_10141),
        .dout(new_Jinkela_wire_10142)
    );

    bfr new_Jinkela_buffer_8123 (
        .din(new_Jinkela_wire_10004),
        .dout(new_Jinkela_wire_10005)
    );

    bfr new_Jinkela_buffer_8249 (
        .din(new_Jinkela_wire_10172),
        .dout(new_Jinkela_wire_10173)
    );

    bfr new_Jinkela_buffer_8124 (
        .din(new_Jinkela_wire_10005),
        .dout(new_Jinkela_wire_10006)
    );

    bfr new_Jinkela_buffer_8221 (
        .din(new_Jinkela_wire_10142),
        .dout(new_Jinkela_wire_10143)
    );

    bfr new_Jinkela_buffer_8125 (
        .din(new_Jinkela_wire_10006),
        .dout(new_Jinkela_wire_10007)
    );

    bfr new_Jinkela_buffer_8126 (
        .din(new_Jinkela_wire_10007),
        .dout(new_Jinkela_wire_10008)
    );

    bfr new_Jinkela_buffer_8327 (
        .din(_0426_),
        .dout(new_Jinkela_wire_10265)
    );

    bfr new_Jinkela_buffer_8222 (
        .din(new_Jinkela_wire_10143),
        .dout(new_Jinkela_wire_10144)
    );

    bfr new_Jinkela_buffer_8127 (
        .din(new_Jinkela_wire_10008),
        .dout(new_Jinkela_wire_10009)
    );

    bfr new_Jinkela_buffer_8250 (
        .din(new_Jinkela_wire_10173),
        .dout(new_Jinkela_wire_10174)
    );

    bfr new_Jinkela_buffer_8128 (
        .din(new_Jinkela_wire_10009),
        .dout(new_Jinkela_wire_10010)
    );

    bfr new_Jinkela_buffer_8223 (
        .din(new_Jinkela_wire_10144),
        .dout(new_Jinkela_wire_10145)
    );

    bfr new_Jinkela_buffer_8129 (
        .din(new_Jinkela_wire_10010),
        .dout(new_Jinkela_wire_10011)
    );

    bfr new_Jinkela_buffer_8284 (
        .din(new_Jinkela_wire_10211),
        .dout(new_Jinkela_wire_10212)
    );

    bfr new_Jinkela_buffer_8130 (
        .din(new_Jinkela_wire_10011),
        .dout(new_Jinkela_wire_10012)
    );

    bfr new_Jinkela_buffer_8224 (
        .din(new_Jinkela_wire_10145),
        .dout(new_Jinkela_wire_10146)
    );

    bfr new_Jinkela_buffer_8131 (
        .din(new_Jinkela_wire_10012),
        .dout(new_Jinkela_wire_10013)
    );

    bfr new_Jinkela_buffer_8251 (
        .din(new_Jinkela_wire_10174),
        .dout(new_Jinkela_wire_10175)
    );

    bfr new_Jinkela_buffer_8132 (
        .din(new_Jinkela_wire_10013),
        .dout(new_Jinkela_wire_10014)
    );

    bfr new_Jinkela_buffer_8225 (
        .din(new_Jinkela_wire_10146),
        .dout(new_Jinkela_wire_10147)
    );

    bfr new_Jinkela_buffer_8133 (
        .din(new_Jinkela_wire_10014),
        .dout(new_Jinkela_wire_10015)
    );

    bfr new_Jinkela_buffer_8134 (
        .din(new_Jinkela_wire_10015),
        .dout(new_Jinkela_wire_10016)
    );

    bfr new_Jinkela_buffer_8335 (
        .din(_0473_),
        .dout(new_Jinkela_wire_10275)
    );

    bfr new_Jinkela_buffer_8226 (
        .din(new_Jinkela_wire_10147),
        .dout(new_Jinkela_wire_10148)
    );

    bfr new_Jinkela_buffer_8135 (
        .din(new_Jinkela_wire_10016),
        .dout(new_Jinkela_wire_10017)
    );

    bfr new_Jinkela_buffer_4716 (
        .din(new_Jinkela_wire_6129),
        .dout(new_Jinkela_wire_6130)
    );

    spl2 new_Jinkela_splitter_1057 (
        .a(_0854_),
        .b(new_Jinkela_wire_14184),
        .c(new_Jinkela_wire_14185)
    );

    bfr new_Jinkela_buffer_4671 (
        .din(new_Jinkela_wire_6082),
        .dout(new_Jinkela_wire_6083)
    );

    spl2 new_Jinkela_splitter_1023 (
        .a(new_Jinkela_wire_13951),
        .b(new_Jinkela_wire_13952),
        .c(new_Jinkela_wire_13953)
    );

    bfr new_Jinkela_buffer_4820 (
        .din(new_Jinkela_wire_6251),
        .dout(new_Jinkela_wire_6252)
    );

    spl2 new_Jinkela_splitter_1058 (
        .a(_0770_),
        .b(new_Jinkela_wire_14190),
        .c(new_Jinkela_wire_14191)
    );

    bfr new_Jinkela_buffer_4672 (
        .din(new_Jinkela_wire_6083),
        .dout(new_Jinkela_wire_6084)
    );

    bfr new_Jinkela_buffer_11662 (
        .din(new_Jinkela_wire_14063),
        .dout(new_Jinkela_wire_14064)
    );

    bfr new_Jinkela_buffer_4717 (
        .din(new_Jinkela_wire_6130),
        .dout(new_Jinkela_wire_6131)
    );

    bfr new_Jinkela_buffer_11663 (
        .din(new_Jinkela_wire_14064),
        .dout(new_Jinkela_wire_14065)
    );

    bfr new_Jinkela_buffer_4673 (
        .din(new_Jinkela_wire_6084),
        .dout(new_Jinkela_wire_6085)
    );

    bfr new_Jinkela_buffer_11689 (
        .din(new_Jinkela_wire_14102),
        .dout(new_Jinkela_wire_14103)
    );

    bfr new_Jinkela_buffer_4795 (
        .din(new_Jinkela_wire_6218),
        .dout(new_Jinkela_wire_6219)
    );

    bfr new_Jinkela_buffer_11664 (
        .din(new_Jinkela_wire_14065),
        .dout(new_Jinkela_wire_14066)
    );

    bfr new_Jinkela_buffer_4674 (
        .din(new_Jinkela_wire_6085),
        .dout(new_Jinkela_wire_6086)
    );

    bfr new_Jinkela_buffer_4718 (
        .din(new_Jinkela_wire_6131),
        .dout(new_Jinkela_wire_6132)
    );

    bfr new_Jinkela_buffer_11665 (
        .din(new_Jinkela_wire_14066),
        .dout(new_Jinkela_wire_14067)
    );

    bfr new_Jinkela_buffer_4675 (
        .din(new_Jinkela_wire_6086),
        .dout(new_Jinkela_wire_6087)
    );

    bfr new_Jinkela_buffer_11690 (
        .din(new_Jinkela_wire_14103),
        .dout(new_Jinkela_wire_14104)
    );

    spl2 new_Jinkela_splitter_566 (
        .a(_1087_),
        .b(new_Jinkela_wire_6365),
        .c(new_Jinkela_wire_6366)
    );

    bfr new_Jinkela_buffer_11666 (
        .din(new_Jinkela_wire_14067),
        .dout(new_Jinkela_wire_14068)
    );

    bfr new_Jinkela_buffer_4824 (
        .din(new_Jinkela_wire_6255),
        .dout(new_Jinkela_wire_6256)
    );

    bfr new_Jinkela_buffer_4676 (
        .din(new_Jinkela_wire_6087),
        .dout(new_Jinkela_wire_6088)
    );

    bfr new_Jinkela_buffer_11768 (
        .din(new_Jinkela_wire_14185),
        .dout(new_Jinkela_wire_14186)
    );

    spl2 new_Jinkela_splitter_1059 (
        .a(_1301_),
        .b(new_Jinkela_wire_14192),
        .c(new_Jinkela_wire_14193)
    );

    bfr new_Jinkela_buffer_4719 (
        .din(new_Jinkela_wire_6132),
        .dout(new_Jinkela_wire_6133)
    );

    bfr new_Jinkela_buffer_11667 (
        .din(new_Jinkela_wire_14068),
        .dout(new_Jinkela_wire_14069)
    );

    bfr new_Jinkela_buffer_4677 (
        .din(new_Jinkela_wire_6088),
        .dout(new_Jinkela_wire_6089)
    );

    bfr new_Jinkela_buffer_11691 (
        .din(new_Jinkela_wire_14104),
        .dout(new_Jinkela_wire_14105)
    );

    bfr new_Jinkela_buffer_4796 (
        .din(new_Jinkela_wire_6219),
        .dout(new_Jinkela_wire_6220)
    );

    bfr new_Jinkela_buffer_11668 (
        .din(new_Jinkela_wire_14069),
        .dout(new_Jinkela_wire_14070)
    );

    bfr new_Jinkela_buffer_4678 (
        .din(new_Jinkela_wire_6089),
        .dout(new_Jinkela_wire_6090)
    );

    bfr new_Jinkela_buffer_4720 (
        .din(new_Jinkela_wire_6133),
        .dout(new_Jinkela_wire_6134)
    );

    bfr new_Jinkela_buffer_11669 (
        .din(new_Jinkela_wire_14070),
        .dout(new_Jinkela_wire_14071)
    );

    bfr new_Jinkela_buffer_4679 (
        .din(new_Jinkela_wire_6090),
        .dout(new_Jinkela_wire_6091)
    );

    bfr new_Jinkela_buffer_11692 (
        .din(new_Jinkela_wire_14105),
        .dout(new_Jinkela_wire_14106)
    );

    bfr new_Jinkela_buffer_4821 (
        .din(new_Jinkela_wire_6252),
        .dout(new_Jinkela_wire_6253)
    );

    bfr new_Jinkela_buffer_11670 (
        .din(new_Jinkela_wire_14071),
        .dout(new_Jinkela_wire_14072)
    );

    bfr new_Jinkela_buffer_4680 (
        .din(new_Jinkela_wire_6091),
        .dout(new_Jinkela_wire_6092)
    );

    bfr new_Jinkela_buffer_11769 (
        .din(new_Jinkela_wire_14186),
        .dout(new_Jinkela_wire_14187)
    );

    bfr new_Jinkela_buffer_4721 (
        .din(new_Jinkela_wire_6134),
        .dout(new_Jinkela_wire_6135)
    );

    bfr new_Jinkela_buffer_11671 (
        .din(new_Jinkela_wire_14072),
        .dout(new_Jinkela_wire_14073)
    );

    spl2 new_Jinkela_splitter_555 (
        .a(new_Jinkela_wire_6092),
        .b(new_Jinkela_wire_6093),
        .c(new_Jinkela_wire_6094)
    );

    bfr new_Jinkela_buffer_11693 (
        .din(new_Jinkela_wire_14106),
        .dout(new_Jinkela_wire_14107)
    );

    bfr new_Jinkela_buffer_4722 (
        .din(new_Jinkela_wire_6135),
        .dout(new_Jinkela_wire_6136)
    );

    bfr new_Jinkela_buffer_11672 (
        .din(new_Jinkela_wire_14073),
        .dout(new_Jinkela_wire_14074)
    );

    bfr new_Jinkela_buffer_4797 (
        .din(new_Jinkela_wire_6220),
        .dout(new_Jinkela_wire_6221)
    );

    spl2 new_Jinkela_splitter_1060 (
        .a(_0477_),
        .b(new_Jinkela_wire_14194),
        .c(new_Jinkela_wire_14195)
    );

    bfr new_Jinkela_buffer_11673 (
        .din(new_Jinkela_wire_14074),
        .dout(new_Jinkela_wire_14075)
    );

    spl2 new_Jinkela_splitter_567 (
        .a(_0578_),
        .b(new_Jinkela_wire_6368),
        .c(new_Jinkela_wire_6369)
    );

    bfr new_Jinkela_buffer_4723 (
        .din(new_Jinkela_wire_6136),
        .dout(new_Jinkela_wire_6137)
    );

    bfr new_Jinkela_buffer_11694 (
        .din(new_Jinkela_wire_14107),
        .dout(new_Jinkela_wire_14108)
    );

    bfr new_Jinkela_buffer_4798 (
        .din(new_Jinkela_wire_6221),
        .dout(new_Jinkela_wire_6222)
    );

    spl2 new_Jinkela_splitter_1050 (
        .a(new_Jinkela_wire_14075),
        .b(new_Jinkela_wire_14076),
        .c(new_Jinkela_wire_14077)
    );

    bfr new_Jinkela_buffer_4724 (
        .din(new_Jinkela_wire_6137),
        .dout(new_Jinkela_wire_6138)
    );

    bfr new_Jinkela_buffer_11695 (
        .din(new_Jinkela_wire_14108),
        .dout(new_Jinkela_wire_14109)
    );

    bfr new_Jinkela_buffer_11770 (
        .din(new_Jinkela_wire_14187),
        .dout(new_Jinkela_wire_14188)
    );

    bfr new_Jinkela_buffer_4825 (
        .din(new_Jinkela_wire_6256),
        .dout(new_Jinkela_wire_6257)
    );

    bfr new_Jinkela_buffer_4725 (
        .din(new_Jinkela_wire_6138),
        .dout(new_Jinkela_wire_6139)
    );

    spl2 new_Jinkela_splitter_1061 (
        .a(_0304_),
        .b(new_Jinkela_wire_14196),
        .c(new_Jinkela_wire_14197)
    );

    bfr new_Jinkela_buffer_4799 (
        .din(new_Jinkela_wire_6222),
        .dout(new_Jinkela_wire_6223)
    );

    bfr new_Jinkela_buffer_11696 (
        .din(new_Jinkela_wire_14109),
        .dout(new_Jinkela_wire_14110)
    );

    bfr new_Jinkela_buffer_4726 (
        .din(new_Jinkela_wire_6139),
        .dout(new_Jinkela_wire_6140)
    );

    bfr new_Jinkela_buffer_11771 (
        .din(new_Jinkela_wire_14188),
        .dout(new_Jinkela_wire_14189)
    );

    bfr new_Jinkela_buffer_11697 (
        .din(new_Jinkela_wire_14110),
        .dout(new_Jinkela_wire_14111)
    );

    bfr new_Jinkela_buffer_4727 (
        .din(new_Jinkela_wire_6140),
        .dout(new_Jinkela_wire_6141)
    );

    spl2 new_Jinkela_splitter_1064 (
        .a(_0099_),
        .b(new_Jinkela_wire_14204),
        .c(new_Jinkela_wire_14205)
    );

    bfr new_Jinkela_buffer_11772 (
        .din(_0287_),
        .dout(new_Jinkela_wire_14198)
    );

    bfr new_Jinkela_buffer_4800 (
        .din(new_Jinkela_wire_6223),
        .dout(new_Jinkela_wire_6224)
    );

    bfr new_Jinkela_buffer_11698 (
        .din(new_Jinkela_wire_14111),
        .dout(new_Jinkela_wire_14112)
    );

    bfr new_Jinkela_buffer_4728 (
        .din(new_Jinkela_wire_6141),
        .dout(new_Jinkela_wire_6142)
    );

    bfr new_Jinkela_buffer_11773 (
        .din(_0191_),
        .dout(new_Jinkela_wire_14201)
    );

    spl2 new_Jinkela_splitter_1062 (
        .a(_0510_),
        .b(new_Jinkela_wire_14199),
        .c(new_Jinkela_wire_14200)
    );

    bfr new_Jinkela_buffer_11699 (
        .din(new_Jinkela_wire_14112),
        .dout(new_Jinkela_wire_14113)
    );

    bfr new_Jinkela_buffer_4826 (
        .din(new_Jinkela_wire_6257),
        .dout(new_Jinkela_wire_6258)
    );

    bfr new_Jinkela_buffer_4729 (
        .din(new_Jinkela_wire_6142),
        .dout(new_Jinkela_wire_6143)
    );

    bfr new_Jinkela_buffer_4801 (
        .din(new_Jinkela_wire_6224),
        .dout(new_Jinkela_wire_6225)
    );

    bfr new_Jinkela_buffer_11700 (
        .din(new_Jinkela_wire_14113),
        .dout(new_Jinkela_wire_14114)
    );

    bfr new_Jinkela_buffer_4730 (
        .din(new_Jinkela_wire_6143),
        .dout(new_Jinkela_wire_6144)
    );

    spl2 new_Jinkela_splitter_1063 (
        .a(_0088_),
        .b(new_Jinkela_wire_14202),
        .c(new_Jinkela_wire_14203)
    );

    bfr new_Jinkela_buffer_11701 (
        .din(new_Jinkela_wire_14114),
        .dout(new_Jinkela_wire_14115)
    );

    bfr new_Jinkela_buffer_4931 (
        .din(_0896_),
        .dout(new_Jinkela_wire_6367)
    );

    bfr new_Jinkela_buffer_4731 (
        .din(new_Jinkela_wire_6144),
        .dout(new_Jinkela_wire_6145)
    );

    spl2 new_Jinkela_splitter_1065 (
        .a(_1038_),
        .b(new_Jinkela_wire_14210),
        .c(new_Jinkela_wire_14211)
    );

    bfr new_Jinkela_buffer_15073 (
        .din(new_Jinkela_wire_17971),
        .dout(new_Jinkela_wire_17972)
    );

    bfr new_Jinkela_buffer_15192 (
        .din(new_Jinkela_wire_18126),
        .dout(new_Jinkela_wire_18127)
    );

    spl2 new_Jinkela_splitter_1298 (
        .a(new_Jinkela_wire_17972),
        .b(new_Jinkela_wire_17973),
        .c(new_Jinkela_wire_17974)
    );

    spl2 new_Jinkela_splitter_1321 (
        .a(_0719_),
        .b(new_Jinkela_wire_18283),
        .c(new_Jinkela_wire_18284)
    );

    bfr new_Jinkela_buffer_15098 (
        .din(new_Jinkela_wire_18018),
        .dout(new_Jinkela_wire_18019)
    );

    bfr new_Jinkela_buffer_15099 (
        .din(new_Jinkela_wire_18019),
        .dout(new_Jinkela_wire_18020)
    );

    bfr new_Jinkela_buffer_15193 (
        .din(new_Jinkela_wire_18127),
        .dout(new_Jinkela_wire_18128)
    );

    bfr new_Jinkela_buffer_15100 (
        .din(new_Jinkela_wire_18020),
        .dout(new_Jinkela_wire_18021)
    );

    spl2 new_Jinkela_splitter_1320 (
        .a(_0601_),
        .b(new_Jinkela_wire_18277),
        .c(new_Jinkela_wire_18278)
    );

    bfr new_Jinkela_buffer_15101 (
        .din(new_Jinkela_wire_18021),
        .dout(new_Jinkela_wire_18022)
    );

    bfr new_Jinkela_buffer_15194 (
        .din(new_Jinkela_wire_18128),
        .dout(new_Jinkela_wire_18129)
    );

    bfr new_Jinkela_buffer_15102 (
        .din(new_Jinkela_wire_18022),
        .dout(new_Jinkela_wire_18023)
    );

    bfr new_Jinkela_buffer_15287 (
        .din(new_Jinkela_wire_18227),
        .dout(new_Jinkela_wire_18228)
    );

    bfr new_Jinkela_buffer_15103 (
        .din(new_Jinkela_wire_18023),
        .dout(new_Jinkela_wire_18024)
    );

    bfr new_Jinkela_buffer_15195 (
        .din(new_Jinkela_wire_18129),
        .dout(new_Jinkela_wire_18130)
    );

    bfr new_Jinkela_buffer_15104 (
        .din(new_Jinkela_wire_18024),
        .dout(new_Jinkela_wire_18025)
    );

    bfr new_Jinkela_buffer_15105 (
        .din(new_Jinkela_wire_18025),
        .dout(new_Jinkela_wire_18026)
    );

    bfr new_Jinkela_buffer_15196 (
        .din(new_Jinkela_wire_18130),
        .dout(new_Jinkela_wire_18131)
    );

    bfr new_Jinkela_buffer_15106 (
        .din(new_Jinkela_wire_18026),
        .dout(new_Jinkela_wire_18027)
    );

    bfr new_Jinkela_buffer_15288 (
        .din(new_Jinkela_wire_18228),
        .dout(new_Jinkela_wire_18229)
    );

    bfr new_Jinkela_buffer_15107 (
        .din(new_Jinkela_wire_18027),
        .dout(new_Jinkela_wire_18028)
    );

    bfr new_Jinkela_buffer_15197 (
        .din(new_Jinkela_wire_18131),
        .dout(new_Jinkela_wire_18132)
    );

    bfr new_Jinkela_buffer_15108 (
        .din(new_Jinkela_wire_18028),
        .dout(new_Jinkela_wire_18029)
    );

    bfr new_Jinkela_buffer_15334 (
        .din(new_Jinkela_wire_18278),
        .dout(new_Jinkela_wire_18279)
    );

    bfr new_Jinkela_buffer_15342 (
        .din(_0483_),
        .dout(new_Jinkela_wire_18289)
    );

    bfr new_Jinkela_buffer_15109 (
        .din(new_Jinkela_wire_18029),
        .dout(new_Jinkela_wire_18030)
    );

    bfr new_Jinkela_buffer_15198 (
        .din(new_Jinkela_wire_18132),
        .dout(new_Jinkela_wire_18133)
    );

    bfr new_Jinkela_buffer_15110 (
        .din(new_Jinkela_wire_18030),
        .dout(new_Jinkela_wire_18031)
    );

    bfr new_Jinkela_buffer_15289 (
        .din(new_Jinkela_wire_18229),
        .dout(new_Jinkela_wire_18230)
    );

    bfr new_Jinkela_buffer_15111 (
        .din(new_Jinkela_wire_18031),
        .dout(new_Jinkela_wire_18032)
    );

    bfr new_Jinkela_buffer_15199 (
        .din(new_Jinkela_wire_18133),
        .dout(new_Jinkela_wire_18134)
    );

    bfr new_Jinkela_buffer_15112 (
        .din(new_Jinkela_wire_18032),
        .dout(new_Jinkela_wire_18033)
    );

    bfr new_Jinkela_buffer_15338 (
        .din(new_Jinkela_wire_18284),
        .dout(new_Jinkela_wire_18285)
    );

    bfr new_Jinkela_buffer_15113 (
        .din(new_Jinkela_wire_18033),
        .dout(new_Jinkela_wire_18034)
    );

    bfr new_Jinkela_buffer_15200 (
        .din(new_Jinkela_wire_18134),
        .dout(new_Jinkela_wire_18135)
    );

    bfr new_Jinkela_buffer_15114 (
        .din(new_Jinkela_wire_18034),
        .dout(new_Jinkela_wire_18035)
    );

    bfr new_Jinkela_buffer_15290 (
        .din(new_Jinkela_wire_18230),
        .dout(new_Jinkela_wire_18231)
    );

    bfr new_Jinkela_buffer_15115 (
        .din(new_Jinkela_wire_18035),
        .dout(new_Jinkela_wire_18036)
    );

    bfr new_Jinkela_buffer_15201 (
        .din(new_Jinkela_wire_18135),
        .dout(new_Jinkela_wire_18136)
    );

    bfr new_Jinkela_buffer_15116 (
        .din(new_Jinkela_wire_18036),
        .dout(new_Jinkela_wire_18037)
    );

    bfr new_Jinkela_buffer_15335 (
        .din(new_Jinkela_wire_18279),
        .dout(new_Jinkela_wire_18280)
    );

    bfr new_Jinkela_buffer_15117 (
        .din(new_Jinkela_wire_18037),
        .dout(new_Jinkela_wire_18038)
    );

    bfr new_Jinkela_buffer_8252 (
        .din(new_Jinkela_wire_10175),
        .dout(new_Jinkela_wire_10176)
    );

    bfr new_Jinkela_buffer_8136 (
        .din(new_Jinkela_wire_10017),
        .dout(new_Jinkela_wire_10018)
    );

    bfr new_Jinkela_buffer_8227 (
        .din(new_Jinkela_wire_10148),
        .dout(new_Jinkela_wire_10149)
    );

    bfr new_Jinkela_buffer_8137 (
        .din(new_Jinkela_wire_10018),
        .dout(new_Jinkela_wire_10019)
    );

    bfr new_Jinkela_buffer_8285 (
        .din(new_Jinkela_wire_10212),
        .dout(new_Jinkela_wire_10213)
    );

    bfr new_Jinkela_buffer_8138 (
        .din(new_Jinkela_wire_10019),
        .dout(new_Jinkela_wire_10020)
    );

    bfr new_Jinkela_buffer_8228 (
        .din(new_Jinkela_wire_10149),
        .dout(new_Jinkela_wire_10150)
    );

    bfr new_Jinkela_buffer_8139 (
        .din(new_Jinkela_wire_10020),
        .dout(new_Jinkela_wire_10021)
    );

    bfr new_Jinkela_buffer_8253 (
        .din(new_Jinkela_wire_10176),
        .dout(new_Jinkela_wire_10177)
    );

    bfr new_Jinkela_buffer_8140 (
        .din(new_Jinkela_wire_10021),
        .dout(new_Jinkela_wire_10022)
    );

    bfr new_Jinkela_buffer_8229 (
        .din(new_Jinkela_wire_10150),
        .dout(new_Jinkela_wire_10151)
    );

    bfr new_Jinkela_buffer_8141 (
        .din(new_Jinkela_wire_10022),
        .dout(new_Jinkela_wire_10023)
    );

    bfr new_Jinkela_buffer_8328 (
        .din(new_Jinkela_wire_10265),
        .dout(new_Jinkela_wire_10266)
    );

    bfr new_Jinkela_buffer_8142 (
        .din(new_Jinkela_wire_10023),
        .dout(new_Jinkela_wire_10024)
    );

    bfr new_Jinkela_buffer_8230 (
        .din(new_Jinkela_wire_10151),
        .dout(new_Jinkela_wire_10152)
    );

    bfr new_Jinkela_buffer_8143 (
        .din(new_Jinkela_wire_10024),
        .dout(new_Jinkela_wire_10025)
    );

    bfr new_Jinkela_buffer_8254 (
        .din(new_Jinkela_wire_10177),
        .dout(new_Jinkela_wire_10178)
    );

    bfr new_Jinkela_buffer_8144 (
        .din(new_Jinkela_wire_10025),
        .dout(new_Jinkela_wire_10026)
    );

    bfr new_Jinkela_buffer_8231 (
        .din(new_Jinkela_wire_10152),
        .dout(new_Jinkela_wire_10153)
    );

    bfr new_Jinkela_buffer_8145 (
        .din(new_Jinkela_wire_10026),
        .dout(new_Jinkela_wire_10027)
    );

    bfr new_Jinkela_buffer_8286 (
        .din(new_Jinkela_wire_10213),
        .dout(new_Jinkela_wire_10214)
    );

    bfr new_Jinkela_buffer_8146 (
        .din(new_Jinkela_wire_10027),
        .dout(new_Jinkela_wire_10028)
    );

    bfr new_Jinkela_buffer_8232 (
        .din(new_Jinkela_wire_10153),
        .dout(new_Jinkela_wire_10154)
    );

    bfr new_Jinkela_buffer_8147 (
        .din(new_Jinkela_wire_10028),
        .dout(new_Jinkela_wire_10029)
    );

    bfr new_Jinkela_buffer_8255 (
        .din(new_Jinkela_wire_10178),
        .dout(new_Jinkela_wire_10179)
    );

    bfr new_Jinkela_buffer_8148 (
        .din(new_Jinkela_wire_10029),
        .dout(new_Jinkela_wire_10030)
    );

    bfr new_Jinkela_buffer_8233 (
        .din(new_Jinkela_wire_10154),
        .dout(new_Jinkela_wire_10155)
    );

    bfr new_Jinkela_buffer_8149 (
        .din(new_Jinkela_wire_10030),
        .dout(new_Jinkela_wire_10031)
    );

    bfr new_Jinkela_buffer_8150 (
        .din(new_Jinkela_wire_10031),
        .dout(new_Jinkela_wire_10032)
    );

    bfr new_Jinkela_buffer_8337 (
        .din(_0118_),
        .dout(new_Jinkela_wire_10277)
    );

    bfr new_Jinkela_buffer_8234 (
        .din(new_Jinkela_wire_10155),
        .dout(new_Jinkela_wire_10156)
    );

    bfr new_Jinkela_buffer_8151 (
        .din(new_Jinkela_wire_10032),
        .dout(new_Jinkela_wire_10033)
    );

    bfr new_Jinkela_buffer_8256 (
        .din(new_Jinkela_wire_10179),
        .dout(new_Jinkela_wire_10180)
    );

    bfr new_Jinkela_buffer_8152 (
        .din(new_Jinkela_wire_10033),
        .dout(new_Jinkela_wire_10034)
    );

    bfr new_Jinkela_buffer_8235 (
        .din(new_Jinkela_wire_10156),
        .dout(new_Jinkela_wire_10157)
    );

    bfr new_Jinkela_buffer_8153 (
        .din(new_Jinkela_wire_10034),
        .dout(new_Jinkela_wire_10035)
    );

    bfr new_Jinkela_buffer_8287 (
        .din(new_Jinkela_wire_10214),
        .dout(new_Jinkela_wire_10215)
    );

    bfr new_Jinkela_buffer_8154 (
        .din(new_Jinkela_wire_10035),
        .dout(new_Jinkela_wire_10036)
    );

    bfr new_Jinkela_buffer_8236 (
        .din(new_Jinkela_wire_10157),
        .dout(new_Jinkela_wire_10158)
    );

    bfr new_Jinkela_buffer_8155 (
        .din(new_Jinkela_wire_10036),
        .dout(new_Jinkela_wire_10037)
    );

    bfr new_Jinkela_buffer_8257 (
        .din(new_Jinkela_wire_10180),
        .dout(new_Jinkela_wire_10181)
    );

    bfr new_Jinkela_buffer_8156 (
        .din(new_Jinkela_wire_10037),
        .dout(new_Jinkela_wire_10038)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(new_Jinkela_wire_1954),
        .dout(new_Jinkela_wire_1955)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_2036),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(new_Jinkela_wire_1955),
        .dout(new_Jinkela_wire_1956)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_2139),
        .dout(new_Jinkela_wire_2140)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(new_Jinkela_wire_1956),
        .dout(new_Jinkela_wire_1957)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    spl2 new_Jinkela_splitter_273 (
        .a(_0671_),
        .b(new_Jinkela_wire_2147),
        .c(new_Jinkela_wire_2148)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_1958),
        .dout(new_Jinkela_wire_1959)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(new_Jinkela_wire_1959),
        .dout(new_Jinkela_wire_1960)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_Jinkela_wire_2140),
        .dout(new_Jinkela_wire_2141)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_Jinkela_wire_1960),
        .dout(new_Jinkela_wire_1961)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(new_Jinkela_wire_1961),
        .dout(new_Jinkela_wire_1962)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(_1604_),
        .dout(new_Jinkela_wire_2149)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(new_Jinkela_wire_1962),
        .dout(new_Jinkela_wire_1963)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_1963),
        .dout(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_2141),
        .dout(new_Jinkela_wire_2142)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_1964),
        .dout(new_Jinkela_wire_1965)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_Jinkela_wire_2041),
        .dout(new_Jinkela_wire_2042)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(_0089_),
        .dout(new_Jinkela_wire_2152)
    );

    spl2 new_Jinkela_splitter_274 (
        .a(_0820_),
        .b(new_Jinkela_wire_2150),
        .c(new_Jinkela_wire_2151)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(new_Jinkela_wire_1966),
        .dout(new_Jinkela_wire_1967)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(new_Jinkela_wire_2042),
        .dout(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(new_Jinkela_wire_1967),
        .dout(new_Jinkela_wire_1968)
    );

    spl2 new_Jinkela_splitter_277 (
        .a(_0994_),
        .b(new_Jinkela_wire_2257),
        .c(new_Jinkela_wire_2258)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_1968),
        .dout(new_Jinkela_wire_1969)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_1969),
        .dout(new_Jinkela_wire_1970)
    );

    spl2 new_Jinkela_splitter_276 (
        .a(_0140_),
        .b(new_Jinkela_wire_2251),
        .c(new_Jinkela_wire_2252)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_1970),
        .dout(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(new_Jinkela_wire_2044),
        .dout(new_Jinkela_wire_2045)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(new_Jinkela_wire_1971),
        .dout(new_Jinkela_wire_1972)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_Jinkela_wire_2152),
        .dout(new_Jinkela_wire_2153)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_1972),
        .dout(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_1973),
        .dout(new_Jinkela_wire_1974)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_2252),
        .dout(new_Jinkela_wire_2253)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_1974),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_15202 (
        .din(new_Jinkela_wire_18136),
        .dout(new_Jinkela_wire_18137)
    );

    bfr new_Jinkela_buffer_8237 (
        .din(new_Jinkela_wire_10158),
        .dout(new_Jinkela_wire_10159)
    );

    bfr new_Jinkela_buffer_15118 (
        .din(new_Jinkela_wire_18038),
        .dout(new_Jinkela_wire_18039)
    );

    bfr new_Jinkela_buffer_8157 (
        .din(new_Jinkela_wire_10038),
        .dout(new_Jinkela_wire_10039)
    );

    bfr new_Jinkela_buffer_15291 (
        .din(new_Jinkela_wire_18231),
        .dout(new_Jinkela_wire_18232)
    );

    bfr new_Jinkela_buffer_8329 (
        .din(new_Jinkela_wire_10266),
        .dout(new_Jinkela_wire_10267)
    );

    bfr new_Jinkela_buffer_15119 (
        .din(new_Jinkela_wire_18039),
        .dout(new_Jinkela_wire_18040)
    );

    bfr new_Jinkela_buffer_8158 (
        .din(new_Jinkela_wire_10039),
        .dout(new_Jinkela_wire_10040)
    );

    bfr new_Jinkela_buffer_15203 (
        .din(new_Jinkela_wire_18137),
        .dout(new_Jinkela_wire_18138)
    );

    spl2 new_Jinkela_splitter_810 (
        .a(new_Jinkela_wire_10159),
        .b(new_Jinkela_wire_10160),
        .c(new_Jinkela_wire_10161)
    );

    bfr new_Jinkela_buffer_15120 (
        .din(new_Jinkela_wire_18040),
        .dout(new_Jinkela_wire_18041)
    );

    bfr new_Jinkela_buffer_8159 (
        .din(new_Jinkela_wire_10040),
        .dout(new_Jinkela_wire_10041)
    );

    bfr new_Jinkela_buffer_15343 (
        .din(_0313_),
        .dout(new_Jinkela_wire_18290)
    );

    bfr new_Jinkela_buffer_8288 (
        .din(new_Jinkela_wire_10215),
        .dout(new_Jinkela_wire_10216)
    );

    bfr new_Jinkela_buffer_15121 (
        .din(new_Jinkela_wire_18041),
        .dout(new_Jinkela_wire_18042)
    );

    bfr new_Jinkela_buffer_8160 (
        .din(new_Jinkela_wire_10041),
        .dout(new_Jinkela_wire_10042)
    );

    bfr new_Jinkela_buffer_15204 (
        .din(new_Jinkela_wire_18138),
        .dout(new_Jinkela_wire_18139)
    );

    bfr new_Jinkela_buffer_8258 (
        .din(new_Jinkela_wire_10181),
        .dout(new_Jinkela_wire_10182)
    );

    bfr new_Jinkela_buffer_15122 (
        .din(new_Jinkela_wire_18042),
        .dout(new_Jinkela_wire_18043)
    );

    bfr new_Jinkela_buffer_8161 (
        .din(new_Jinkela_wire_10042),
        .dout(new_Jinkela_wire_10043)
    );

    bfr new_Jinkela_buffer_15292 (
        .din(new_Jinkela_wire_18232),
        .dout(new_Jinkela_wire_18233)
    );

    bfr new_Jinkela_buffer_8259 (
        .din(new_Jinkela_wire_10182),
        .dout(new_Jinkela_wire_10183)
    );

    bfr new_Jinkela_buffer_15123 (
        .din(new_Jinkela_wire_18043),
        .dout(new_Jinkela_wire_18044)
    );

    bfr new_Jinkela_buffer_8162 (
        .din(new_Jinkela_wire_10043),
        .dout(new_Jinkela_wire_10044)
    );

    bfr new_Jinkela_buffer_15205 (
        .din(new_Jinkela_wire_18139),
        .dout(new_Jinkela_wire_18140)
    );

    bfr new_Jinkela_buffer_15124 (
        .din(new_Jinkela_wire_18044),
        .dout(new_Jinkela_wire_18045)
    );

    bfr new_Jinkela_buffer_8163 (
        .din(new_Jinkela_wire_10044),
        .dout(new_Jinkela_wire_10045)
    );

    bfr new_Jinkela_buffer_15336 (
        .din(new_Jinkela_wire_18280),
        .dout(new_Jinkela_wire_18281)
    );

    spl2 new_Jinkela_splitter_819 (
        .a(_1236_),
        .b(new_Jinkela_wire_10278),
        .c(new_Jinkela_wire_10279)
    );

    bfr new_Jinkela_buffer_8260 (
        .din(new_Jinkela_wire_10183),
        .dout(new_Jinkela_wire_10184)
    );

    bfr new_Jinkela_buffer_15125 (
        .din(new_Jinkela_wire_18045),
        .dout(new_Jinkela_wire_18046)
    );

    bfr new_Jinkela_buffer_8164 (
        .din(new_Jinkela_wire_10045),
        .dout(new_Jinkela_wire_10046)
    );

    bfr new_Jinkela_buffer_15206 (
        .din(new_Jinkela_wire_18140),
        .dout(new_Jinkela_wire_18141)
    );

    bfr new_Jinkela_buffer_8289 (
        .din(new_Jinkela_wire_10216),
        .dout(new_Jinkela_wire_10217)
    );

    bfr new_Jinkela_buffer_15126 (
        .din(new_Jinkela_wire_18046),
        .dout(new_Jinkela_wire_18047)
    );

    bfr new_Jinkela_buffer_8165 (
        .din(new_Jinkela_wire_10046),
        .dout(new_Jinkela_wire_10047)
    );

    bfr new_Jinkela_buffer_15293 (
        .din(new_Jinkela_wire_18233),
        .dout(new_Jinkela_wire_18234)
    );

    bfr new_Jinkela_buffer_8261 (
        .din(new_Jinkela_wire_10184),
        .dout(new_Jinkela_wire_10185)
    );

    bfr new_Jinkela_buffer_15127 (
        .din(new_Jinkela_wire_18047),
        .dout(new_Jinkela_wire_18048)
    );

    bfr new_Jinkela_buffer_8330 (
        .din(new_Jinkela_wire_10267),
        .dout(new_Jinkela_wire_10268)
    );

    bfr new_Jinkela_buffer_15207 (
        .din(new_Jinkela_wire_18141),
        .dout(new_Jinkela_wire_18142)
    );

    bfr new_Jinkela_buffer_8262 (
        .din(new_Jinkela_wire_10185),
        .dout(new_Jinkela_wire_10186)
    );

    bfr new_Jinkela_buffer_15128 (
        .din(new_Jinkela_wire_18048),
        .dout(new_Jinkela_wire_18049)
    );

    bfr new_Jinkela_buffer_8290 (
        .din(new_Jinkela_wire_10217),
        .dout(new_Jinkela_wire_10218)
    );

    spl2 new_Jinkela_splitter_1322 (
        .a(_0732_),
        .b(new_Jinkela_wire_18291),
        .c(new_Jinkela_wire_18292)
    );

    bfr new_Jinkela_buffer_8263 (
        .din(new_Jinkela_wire_10186),
        .dout(new_Jinkela_wire_10187)
    );

    bfr new_Jinkela_buffer_15129 (
        .din(new_Jinkela_wire_18049),
        .dout(new_Jinkela_wire_18050)
    );

    bfr new_Jinkela_buffer_8338 (
        .din(_0829_),
        .dout(new_Jinkela_wire_10280)
    );

    bfr new_Jinkela_buffer_15208 (
        .din(new_Jinkela_wire_18142),
        .dout(new_Jinkela_wire_18143)
    );

    bfr new_Jinkela_buffer_8264 (
        .din(new_Jinkela_wire_10187),
        .dout(new_Jinkela_wire_10188)
    );

    bfr new_Jinkela_buffer_15130 (
        .din(new_Jinkela_wire_18050),
        .dout(new_Jinkela_wire_18051)
    );

    bfr new_Jinkela_buffer_8291 (
        .din(new_Jinkela_wire_10218),
        .dout(new_Jinkela_wire_10219)
    );

    bfr new_Jinkela_buffer_15294 (
        .din(new_Jinkela_wire_18234),
        .dout(new_Jinkela_wire_18235)
    );

    bfr new_Jinkela_buffer_8265 (
        .din(new_Jinkela_wire_10188),
        .dout(new_Jinkela_wire_10189)
    );

    bfr new_Jinkela_buffer_15131 (
        .din(new_Jinkela_wire_18051),
        .dout(new_Jinkela_wire_18052)
    );

    bfr new_Jinkela_buffer_8331 (
        .din(new_Jinkela_wire_10268),
        .dout(new_Jinkela_wire_10269)
    );

    bfr new_Jinkela_buffer_15209 (
        .din(new_Jinkela_wire_18143),
        .dout(new_Jinkela_wire_18144)
    );

    bfr new_Jinkela_buffer_8266 (
        .din(new_Jinkela_wire_10189),
        .dout(new_Jinkela_wire_10190)
    );

    bfr new_Jinkela_buffer_15132 (
        .din(new_Jinkela_wire_18052),
        .dout(new_Jinkela_wire_18053)
    );

    bfr new_Jinkela_buffer_8292 (
        .din(new_Jinkela_wire_10219),
        .dout(new_Jinkela_wire_10220)
    );

    bfr new_Jinkela_buffer_15337 (
        .din(new_Jinkela_wire_18281),
        .dout(new_Jinkela_wire_18282)
    );

    bfr new_Jinkela_buffer_8267 (
        .din(new_Jinkela_wire_10190),
        .dout(new_Jinkela_wire_10191)
    );

    bfr new_Jinkela_buffer_15133 (
        .din(new_Jinkela_wire_18053),
        .dout(new_Jinkela_wire_18054)
    );

    spl2 new_Jinkela_splitter_821 (
        .a(_0380_),
        .b(new_Jinkela_wire_10395),
        .c(new_Jinkela_wire_10396)
    );

    bfr new_Jinkela_buffer_15210 (
        .din(new_Jinkela_wire_18144),
        .dout(new_Jinkela_wire_18145)
    );

    bfr new_Jinkela_buffer_8268 (
        .din(new_Jinkela_wire_10191),
        .dout(new_Jinkela_wire_10192)
    );

    bfr new_Jinkela_buffer_15134 (
        .din(new_Jinkela_wire_18054),
        .dout(new_Jinkela_wire_18055)
    );

    bfr new_Jinkela_buffer_8293 (
        .din(new_Jinkela_wire_10220),
        .dout(new_Jinkela_wire_10221)
    );

    bfr new_Jinkela_buffer_15295 (
        .din(new_Jinkela_wire_18235),
        .dout(new_Jinkela_wire_18236)
    );

    bfr new_Jinkela_buffer_8269 (
        .din(new_Jinkela_wire_10192),
        .dout(new_Jinkela_wire_10193)
    );

    bfr new_Jinkela_buffer_15135 (
        .din(new_Jinkela_wire_18055),
        .dout(new_Jinkela_wire_18056)
    );

    bfr new_Jinkela_buffer_8332 (
        .din(new_Jinkela_wire_10269),
        .dout(new_Jinkela_wire_10270)
    );

    bfr new_Jinkela_buffer_15211 (
        .din(new_Jinkela_wire_18145),
        .dout(new_Jinkela_wire_18146)
    );

    bfr new_Jinkela_buffer_8270 (
        .din(new_Jinkela_wire_10193),
        .dout(new_Jinkela_wire_10194)
    );

    bfr new_Jinkela_buffer_15136 (
        .din(new_Jinkela_wire_18056),
        .dout(new_Jinkela_wire_18057)
    );

    bfr new_Jinkela_buffer_8294 (
        .din(new_Jinkela_wire_10221),
        .dout(new_Jinkela_wire_10222)
    );

    bfr new_Jinkela_buffer_15339 (
        .din(new_Jinkela_wire_18285),
        .dout(new_Jinkela_wire_18286)
    );

    bfr new_Jinkela_buffer_8271 (
        .din(new_Jinkela_wire_10194),
        .dout(new_Jinkela_wire_10195)
    );

    bfr new_Jinkela_buffer_15137 (
        .din(new_Jinkela_wire_18057),
        .dout(new_Jinkela_wire_18058)
    );

    bfr new_Jinkela_buffer_15212 (
        .din(new_Jinkela_wire_18146),
        .dout(new_Jinkela_wire_18147)
    );

    bfr new_Jinkela_buffer_8450 (
        .din(_1306_),
        .dout(new_Jinkela_wire_10394)
    );

    bfr new_Jinkela_buffer_8272 (
        .din(new_Jinkela_wire_10195),
        .dout(new_Jinkela_wire_10196)
    );

    bfr new_Jinkela_buffer_15138 (
        .din(new_Jinkela_wire_18058),
        .dout(new_Jinkela_wire_18059)
    );

    bfr new_Jinkela_buffer_4802 (
        .din(new_Jinkela_wire_6225),
        .dout(new_Jinkela_wire_6226)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_2046),
        .dout(new_Jinkela_wire_2047)
    );

    bfr new_Jinkela_buffer_4732 (
        .din(new_Jinkela_wire_6145),
        .dout(new_Jinkela_wire_6146)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(new_Jinkela_wire_1975),
        .dout(new_Jinkela_wire_1976)
    );

    spl2 new_Jinkela_splitter_568 (
        .a(_0908_),
        .b(new_Jinkela_wire_6370),
        .c(new_Jinkela_wire_6371)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_2153),
        .dout(new_Jinkela_wire_2154)
    );

    bfr new_Jinkela_buffer_4827 (
        .din(new_Jinkela_wire_6258),
        .dout(new_Jinkela_wire_6259)
    );

    bfr new_Jinkela_buffer_4733 (
        .din(new_Jinkela_wire_6146),
        .dout(new_Jinkela_wire_6147)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(new_Jinkela_wire_1976),
        .dout(new_Jinkela_wire_1977)
    );

    bfr new_Jinkela_buffer_4803 (
        .din(new_Jinkela_wire_6226),
        .dout(new_Jinkela_wire_6227)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_2047),
        .dout(new_Jinkela_wire_2048)
    );

    bfr new_Jinkela_buffer_4734 (
        .din(new_Jinkela_wire_6147),
        .dout(new_Jinkela_wire_6148)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_1977),
        .dout(new_Jinkela_wire_1978)
    );

    spl2 new_Jinkela_splitter_278 (
        .a(_1420_),
        .b(new_Jinkela_wire_2259),
        .c(new_Jinkela_wire_2260)
    );

    bfr new_Jinkela_buffer_4735 (
        .din(new_Jinkela_wire_6148),
        .dout(new_Jinkela_wire_6149)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(new_Jinkela_wire_1978),
        .dout(new_Jinkela_wire_1979)
    );

    bfr new_Jinkela_buffer_4804 (
        .din(new_Jinkela_wire_6227),
        .dout(new_Jinkela_wire_6228)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_Jinkela_wire_2048),
        .dout(new_Jinkela_wire_2049)
    );

    bfr new_Jinkela_buffer_4736 (
        .din(new_Jinkela_wire_6149),
        .dout(new_Jinkela_wire_6150)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_1979),
        .dout(new_Jinkela_wire_1980)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_2154),
        .dout(new_Jinkela_wire_2155)
    );

    bfr new_Jinkela_buffer_4828 (
        .din(new_Jinkela_wire_6259),
        .dout(new_Jinkela_wire_6260)
    );

    bfr new_Jinkela_buffer_4737 (
        .din(new_Jinkela_wire_6150),
        .dout(new_Jinkela_wire_6151)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_1980),
        .dout(new_Jinkela_wire_1981)
    );

    bfr new_Jinkela_buffer_4805 (
        .din(new_Jinkela_wire_6228),
        .dout(new_Jinkela_wire_6229)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_2049),
        .dout(new_Jinkela_wire_2050)
    );

    bfr new_Jinkela_buffer_4738 (
        .din(new_Jinkela_wire_6151),
        .dout(new_Jinkela_wire_6152)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(new_Jinkela_wire_1981),
        .dout(new_Jinkela_wire_1982)
    );

    bfr new_Jinkela_buffer_4739 (
        .din(new_Jinkela_wire_6152),
        .dout(new_Jinkela_wire_6153)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_1982),
        .dout(new_Jinkela_wire_1983)
    );

    bfr new_Jinkela_buffer_4806 (
        .din(new_Jinkela_wire_6229),
        .dout(new_Jinkela_wire_6230)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_2050),
        .dout(new_Jinkela_wire_2051)
    );

    bfr new_Jinkela_buffer_4740 (
        .din(new_Jinkela_wire_6153),
        .dout(new_Jinkela_wire_6154)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(new_Jinkela_wire_1983),
        .dout(new_Jinkela_wire_1984)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_2155),
        .dout(new_Jinkela_wire_2156)
    );

    bfr new_Jinkela_buffer_4829 (
        .din(new_Jinkela_wire_6260),
        .dout(new_Jinkela_wire_6261)
    );

    bfr new_Jinkela_buffer_4741 (
        .din(new_Jinkela_wire_6154),
        .dout(new_Jinkela_wire_6155)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_1984),
        .dout(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_4807 (
        .din(new_Jinkela_wire_6230),
        .dout(new_Jinkela_wire_6231)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_2051),
        .dout(new_Jinkela_wire_2052)
    );

    bfr new_Jinkela_buffer_4742 (
        .din(new_Jinkela_wire_6155),
        .dout(new_Jinkela_wire_6156)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_1985),
        .dout(new_Jinkela_wire_1986)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_2253),
        .dout(new_Jinkela_wire_2254)
    );

    spl2 new_Jinkela_splitter_569 (
        .a(_0541_),
        .b(new_Jinkela_wire_6372),
        .c(new_Jinkela_wire_6373)
    );

    bfr new_Jinkela_buffer_4743 (
        .din(new_Jinkela_wire_6156),
        .dout(new_Jinkela_wire_6157)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_1986),
        .dout(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_4808 (
        .din(new_Jinkela_wire_6231),
        .dout(new_Jinkela_wire_6232)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_2052),
        .dout(new_Jinkela_wire_2053)
    );

    bfr new_Jinkela_buffer_4744 (
        .din(new_Jinkela_wire_6157),
        .dout(new_Jinkela_wire_6158)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_1987),
        .dout(new_Jinkela_wire_1988)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(new_Jinkela_wire_2156),
        .dout(new_Jinkela_wire_2157)
    );

    bfr new_Jinkela_buffer_4830 (
        .din(new_Jinkela_wire_6261),
        .dout(new_Jinkela_wire_6262)
    );

    bfr new_Jinkela_buffer_4745 (
        .din(new_Jinkela_wire_6158),
        .dout(new_Jinkela_wire_6159)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(new_Jinkela_wire_1988),
        .dout(new_Jinkela_wire_1989)
    );

    bfr new_Jinkela_buffer_4809 (
        .din(new_Jinkela_wire_6232),
        .dout(new_Jinkela_wire_6233)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(new_Jinkela_wire_2053),
        .dout(new_Jinkela_wire_2054)
    );

    bfr new_Jinkela_buffer_4746 (
        .din(new_Jinkela_wire_6159),
        .dout(new_Jinkela_wire_6160)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(new_Jinkela_wire_1989),
        .dout(new_Jinkela_wire_1990)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(_1465_),
        .dout(new_Jinkela_wire_2262)
    );

    spl2 new_Jinkela_splitter_570 (
        .a(_0654_),
        .b(new_Jinkela_wire_6374),
        .c(new_Jinkela_wire_6375)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(_0992_),
        .dout(new_Jinkela_wire_2261)
    );

    bfr new_Jinkela_buffer_4747 (
        .din(new_Jinkela_wire_6160),
        .dout(new_Jinkela_wire_6161)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_1990),
        .dout(new_Jinkela_wire_1991)
    );

    bfr new_Jinkela_buffer_4810 (
        .din(new_Jinkela_wire_6233),
        .dout(new_Jinkela_wire_6234)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(new_Jinkela_wire_2054),
        .dout(new_Jinkela_wire_2055)
    );

    bfr new_Jinkela_buffer_4748 (
        .din(new_Jinkela_wire_6161),
        .dout(new_Jinkela_wire_6162)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(new_Jinkela_wire_1991),
        .dout(new_Jinkela_wire_1992)
    );

    spl2 new_Jinkela_splitter_571 (
        .a(_0010_),
        .b(new_Jinkela_wire_6377),
        .c(new_Jinkela_wire_6378)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(new_Jinkela_wire_2157),
        .dout(new_Jinkela_wire_2158)
    );

    bfr new_Jinkela_buffer_4831 (
        .din(new_Jinkela_wire_6262),
        .dout(new_Jinkela_wire_6263)
    );

    bfr new_Jinkela_buffer_4749 (
        .din(new_Jinkela_wire_6162),
        .dout(new_Jinkela_wire_6163)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    bfr new_Jinkela_buffer_4811 (
        .din(new_Jinkela_wire_6234),
        .dout(new_Jinkela_wire_6235)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(new_Jinkela_wire_2055),
        .dout(new_Jinkela_wire_2056)
    );

    bfr new_Jinkela_buffer_4750 (
        .din(new_Jinkela_wire_6163),
        .dout(new_Jinkela_wire_6164)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(new_Jinkela_wire_1993),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_2254),
        .dout(new_Jinkela_wire_2255)
    );

    bfr new_Jinkela_buffer_4932 (
        .din(_1011_),
        .dout(new_Jinkela_wire_6376)
    );

    bfr new_Jinkela_buffer_4751 (
        .din(new_Jinkela_wire_6164),
        .dout(new_Jinkela_wire_6165)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_4812 (
        .din(new_Jinkela_wire_6235),
        .dout(new_Jinkela_wire_6236)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(new_Jinkela_wire_2056),
        .dout(new_Jinkela_wire_2057)
    );

    bfr new_Jinkela_buffer_4752 (
        .din(new_Jinkela_wire_6165),
        .dout(new_Jinkela_wire_6166)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    bfr new_Jinkela_buffer_15296 (
        .din(new_Jinkela_wire_18236),
        .dout(new_Jinkela_wire_18237)
    );

    bfr new_Jinkela_buffer_4933 (
        .din(_1215_),
        .dout(new_Jinkela_wire_6379)
    );

    bfr new_Jinkela_buffer_4832 (
        .din(new_Jinkela_wire_6263),
        .dout(new_Jinkela_wire_6264)
    );

    bfr new_Jinkela_buffer_15139 (
        .din(new_Jinkela_wire_18059),
        .dout(new_Jinkela_wire_18060)
    );

    bfr new_Jinkela_buffer_4753 (
        .din(new_Jinkela_wire_6166),
        .dout(new_Jinkela_wire_6167)
    );

    bfr new_Jinkela_buffer_15213 (
        .din(new_Jinkela_wire_18147),
        .dout(new_Jinkela_wire_18148)
    );

    bfr new_Jinkela_buffer_4813 (
        .din(new_Jinkela_wire_6236),
        .dout(new_Jinkela_wire_6237)
    );

    bfr new_Jinkela_buffer_15140 (
        .din(new_Jinkela_wire_18060),
        .dout(new_Jinkela_wire_18061)
    );

    bfr new_Jinkela_buffer_4754 (
        .din(new_Jinkela_wire_6167),
        .dout(new_Jinkela_wire_6168)
    );

    bfr new_Jinkela_buffer_15344 (
        .din(_1101_),
        .dout(new_Jinkela_wire_18293)
    );

    bfr new_Jinkela_buffer_15141 (
        .din(new_Jinkela_wire_18061),
        .dout(new_Jinkela_wire_18062)
    );

    bfr new_Jinkela_buffer_4755 (
        .din(new_Jinkela_wire_6168),
        .dout(new_Jinkela_wire_6169)
    );

    bfr new_Jinkela_buffer_15214 (
        .din(new_Jinkela_wire_18148),
        .dout(new_Jinkela_wire_18149)
    );

    spl2 new_Jinkela_splitter_574 (
        .a(_1401_),
        .b(new_Jinkela_wire_6407),
        .c(new_Jinkela_wire_6408)
    );

    bfr new_Jinkela_buffer_4833 (
        .din(new_Jinkela_wire_6264),
        .dout(new_Jinkela_wire_6265)
    );

    bfr new_Jinkela_buffer_15142 (
        .din(new_Jinkela_wire_18062),
        .dout(new_Jinkela_wire_18063)
    );

    bfr new_Jinkela_buffer_4756 (
        .din(new_Jinkela_wire_6169),
        .dout(new_Jinkela_wire_6170)
    );

    bfr new_Jinkela_buffer_15297 (
        .din(new_Jinkela_wire_18237),
        .dout(new_Jinkela_wire_18238)
    );

    bfr new_Jinkela_buffer_15143 (
        .din(new_Jinkela_wire_18063),
        .dout(new_Jinkela_wire_18064)
    );

    bfr new_Jinkela_buffer_4757 (
        .din(new_Jinkela_wire_6170),
        .dout(new_Jinkela_wire_6171)
    );

    bfr new_Jinkela_buffer_15215 (
        .din(new_Jinkela_wire_18149),
        .dout(new_Jinkela_wire_18150)
    );

    bfr new_Jinkela_buffer_4834 (
        .din(new_Jinkela_wire_6265),
        .dout(new_Jinkela_wire_6266)
    );

    bfr new_Jinkela_buffer_15144 (
        .din(new_Jinkela_wire_18064),
        .dout(new_Jinkela_wire_18065)
    );

    bfr new_Jinkela_buffer_4758 (
        .din(new_Jinkela_wire_6171),
        .dout(new_Jinkela_wire_6172)
    );

    bfr new_Jinkela_buffer_15340 (
        .din(new_Jinkela_wire_18286),
        .dout(new_Jinkela_wire_18287)
    );

    spl2 new_Jinkela_splitter_573 (
        .a(_1793_),
        .b(new_Jinkela_wire_6405),
        .c(new_Jinkela_wire_6406)
    );

    bfr new_Jinkela_buffer_15145 (
        .din(new_Jinkela_wire_18065),
        .dout(new_Jinkela_wire_18066)
    );

    bfr new_Jinkela_buffer_4759 (
        .din(new_Jinkela_wire_6172),
        .dout(new_Jinkela_wire_6173)
    );

    bfr new_Jinkela_buffer_15216 (
        .din(new_Jinkela_wire_18150),
        .dout(new_Jinkela_wire_18151)
    );

    bfr new_Jinkela_buffer_4934 (
        .din(new_Jinkela_wire_6379),
        .dout(new_Jinkela_wire_6380)
    );

    bfr new_Jinkela_buffer_4835 (
        .din(new_Jinkela_wire_6266),
        .dout(new_Jinkela_wire_6267)
    );

    bfr new_Jinkela_buffer_15146 (
        .din(new_Jinkela_wire_18066),
        .dout(new_Jinkela_wire_18067)
    );

    bfr new_Jinkela_buffer_4760 (
        .din(new_Jinkela_wire_6173),
        .dout(new_Jinkela_wire_6174)
    );

    bfr new_Jinkela_buffer_15298 (
        .din(new_Jinkela_wire_18238),
        .dout(new_Jinkela_wire_18239)
    );

    bfr new_Jinkela_buffer_15147 (
        .din(new_Jinkela_wire_18067),
        .dout(new_Jinkela_wire_18068)
    );

    bfr new_Jinkela_buffer_4761 (
        .din(new_Jinkela_wire_6174),
        .dout(new_Jinkela_wire_6175)
    );

    bfr new_Jinkela_buffer_15217 (
        .din(new_Jinkela_wire_18151),
        .dout(new_Jinkela_wire_18152)
    );

    bfr new_Jinkela_buffer_4836 (
        .din(new_Jinkela_wire_6267),
        .dout(new_Jinkela_wire_6268)
    );

    bfr new_Jinkela_buffer_15148 (
        .din(new_Jinkela_wire_18068),
        .dout(new_Jinkela_wire_18069)
    );

    bfr new_Jinkela_buffer_4762 (
        .din(new_Jinkela_wire_6175),
        .dout(new_Jinkela_wire_6176)
    );

    spl2 new_Jinkela_splitter_1323 (
        .a(_1117_),
        .b(new_Jinkela_wire_18295),
        .c(new_Jinkela_wire_18296)
    );

    bfr new_Jinkela_buffer_15149 (
        .din(new_Jinkela_wire_18069),
        .dout(new_Jinkela_wire_18070)
    );

    bfr new_Jinkela_buffer_4763 (
        .din(new_Jinkela_wire_6176),
        .dout(new_Jinkela_wire_6177)
    );

    bfr new_Jinkela_buffer_15218 (
        .din(new_Jinkela_wire_18152),
        .dout(new_Jinkela_wire_18153)
    );

    bfr new_Jinkela_buffer_4935 (
        .din(new_Jinkela_wire_6380),
        .dout(new_Jinkela_wire_6381)
    );

    bfr new_Jinkela_buffer_4837 (
        .din(new_Jinkela_wire_6268),
        .dout(new_Jinkela_wire_6269)
    );

    bfr new_Jinkela_buffer_15150 (
        .din(new_Jinkela_wire_18070),
        .dout(new_Jinkela_wire_18071)
    );

    bfr new_Jinkela_buffer_4764 (
        .din(new_Jinkela_wire_6177),
        .dout(new_Jinkela_wire_6178)
    );

    bfr new_Jinkela_buffer_15299 (
        .din(new_Jinkela_wire_18239),
        .dout(new_Jinkela_wire_18240)
    );

    bfr new_Jinkela_buffer_15151 (
        .din(new_Jinkela_wire_18071),
        .dout(new_Jinkela_wire_18072)
    );

    bfr new_Jinkela_buffer_4765 (
        .din(new_Jinkela_wire_6178),
        .dout(new_Jinkela_wire_6179)
    );

    bfr new_Jinkela_buffer_15219 (
        .din(new_Jinkela_wire_18153),
        .dout(new_Jinkela_wire_18154)
    );

    bfr new_Jinkela_buffer_4838 (
        .din(new_Jinkela_wire_6269),
        .dout(new_Jinkela_wire_6270)
    );

    bfr new_Jinkela_buffer_15152 (
        .din(new_Jinkela_wire_18072),
        .dout(new_Jinkela_wire_18073)
    );

    bfr new_Jinkela_buffer_4766 (
        .din(new_Jinkela_wire_6179),
        .dout(new_Jinkela_wire_6180)
    );

    bfr new_Jinkela_buffer_15341 (
        .din(new_Jinkela_wire_18287),
        .dout(new_Jinkela_wire_18288)
    );

    spl2 new_Jinkela_splitter_575 (
        .a(_0580_),
        .b(new_Jinkela_wire_6409),
        .c(new_Jinkela_wire_6410)
    );

    bfr new_Jinkela_buffer_15153 (
        .din(new_Jinkela_wire_18073),
        .dout(new_Jinkela_wire_18074)
    );

    bfr new_Jinkela_buffer_4767 (
        .din(new_Jinkela_wire_6180),
        .dout(new_Jinkela_wire_6181)
    );

    bfr new_Jinkela_buffer_15220 (
        .din(new_Jinkela_wire_18154),
        .dout(new_Jinkela_wire_18155)
    );

    bfr new_Jinkela_buffer_4936 (
        .din(new_Jinkela_wire_6381),
        .dout(new_Jinkela_wire_6382)
    );

    bfr new_Jinkela_buffer_4839 (
        .din(new_Jinkela_wire_6270),
        .dout(new_Jinkela_wire_6271)
    );

    bfr new_Jinkela_buffer_15154 (
        .din(new_Jinkela_wire_18074),
        .dout(new_Jinkela_wire_18075)
    );

    bfr new_Jinkela_buffer_4768 (
        .din(new_Jinkela_wire_6181),
        .dout(new_Jinkela_wire_6182)
    );

    bfr new_Jinkela_buffer_15300 (
        .din(new_Jinkela_wire_18240),
        .dout(new_Jinkela_wire_18241)
    );

    bfr new_Jinkela_buffer_15155 (
        .din(new_Jinkela_wire_18075),
        .dout(new_Jinkela_wire_18076)
    );

    bfr new_Jinkela_buffer_4769 (
        .din(new_Jinkela_wire_6182),
        .dout(new_Jinkela_wire_6183)
    );

    bfr new_Jinkela_buffer_15221 (
        .din(new_Jinkela_wire_18155),
        .dout(new_Jinkela_wire_18156)
    );

    spl2 new_Jinkela_splitter_577 (
        .a(_0129_),
        .b(new_Jinkela_wire_6417),
        .c(new_Jinkela_wire_6418)
    );

    bfr new_Jinkela_buffer_4840 (
        .din(new_Jinkela_wire_6271),
        .dout(new_Jinkela_wire_6272)
    );

    bfr new_Jinkela_buffer_15156 (
        .din(new_Jinkela_wire_18076),
        .dout(new_Jinkela_wire_18077)
    );

    bfr new_Jinkela_buffer_4770 (
        .din(new_Jinkela_wire_6183),
        .dout(new_Jinkela_wire_6184)
    );

    spl2 new_Jinkela_splitter_576 (
        .a(_1225_),
        .b(new_Jinkela_wire_6411),
        .c(new_Jinkela_wire_6412)
    );

    bfr new_Jinkela_buffer_15345 (
        .din(_1116_),
        .dout(new_Jinkela_wire_18294)
    );

    bfr new_Jinkela_buffer_15157 (
        .din(new_Jinkela_wire_18077),
        .dout(new_Jinkela_wire_18078)
    );

    bfr new_Jinkela_buffer_4771 (
        .din(new_Jinkela_wire_6184),
        .dout(new_Jinkela_wire_6185)
    );

    bfr new_Jinkela_buffer_15222 (
        .din(new_Jinkela_wire_18156),
        .dout(new_Jinkela_wire_18157)
    );

    bfr new_Jinkela_buffer_4937 (
        .din(new_Jinkela_wire_6382),
        .dout(new_Jinkela_wire_6383)
    );

    bfr new_Jinkela_buffer_4841 (
        .din(new_Jinkela_wire_6272),
        .dout(new_Jinkela_wire_6273)
    );

    bfr new_Jinkela_buffer_15158 (
        .din(new_Jinkela_wire_18078),
        .dout(new_Jinkela_wire_18079)
    );

    bfr new_Jinkela_buffer_4772 (
        .din(new_Jinkela_wire_6185),
        .dout(new_Jinkela_wire_6186)
    );

    bfr new_Jinkela_buffer_15301 (
        .din(new_Jinkela_wire_18241),
        .dout(new_Jinkela_wire_18242)
    );

    bfr new_Jinkela_buffer_15159 (
        .din(new_Jinkela_wire_18079),
        .dout(new_Jinkela_wire_18080)
    );

    bfr new_Jinkela_buffer_4773 (
        .din(new_Jinkela_wire_6186),
        .dout(new_Jinkela_wire_6187)
    );

    bfr new_Jinkela_buffer_11702 (
        .din(new_Jinkela_wire_14115),
        .dout(new_Jinkela_wire_14116)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_2158),
        .dout(new_Jinkela_wire_2159)
    );

    bfr new_Jinkela_buffer_11774 (
        .din(new_Jinkela_wire_14205),
        .dout(new_Jinkela_wire_14206)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_1996),
        .dout(new_Jinkela_wire_1997)
    );

    bfr new_Jinkela_buffer_11703 (
        .din(new_Jinkela_wire_14116),
        .dout(new_Jinkela_wire_14117)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(new_Jinkela_wire_2057),
        .dout(new_Jinkela_wire_2058)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_1997),
        .dout(new_Jinkela_wire_1998)
    );

    bfr new_Jinkela_buffer_11778 (
        .din(_0934_),
        .dout(new_Jinkela_wire_14212)
    );

    bfr new_Jinkela_buffer_11704 (
        .din(new_Jinkela_wire_14117),
        .dout(new_Jinkela_wire_14118)
    );

    spl2 new_Jinkela_splitter_280 (
        .a(_1446_),
        .b(new_Jinkela_wire_2312),
        .c(new_Jinkela_wire_2313)
    );

    spl2 new_Jinkela_splitter_1066 (
        .a(_0498_),
        .b(new_Jinkela_wire_14214),
        .c(new_Jinkela_wire_14215)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_1998),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_11705 (
        .din(new_Jinkela_wire_14118),
        .dout(new_Jinkela_wire_14119)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_2058),
        .dout(new_Jinkela_wire_2059)
    );

    bfr new_Jinkela_buffer_11775 (
        .din(new_Jinkela_wire_14206),
        .dout(new_Jinkela_wire_14207)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_11706 (
        .din(new_Jinkela_wire_14119),
        .dout(new_Jinkela_wire_14120)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_2159),
        .dout(new_Jinkela_wire_2160)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_2000),
        .dout(new_Jinkela_wire_2001)
    );

    bfr new_Jinkela_buffer_11779 (
        .din(_0254_),
        .dout(new_Jinkela_wire_14213)
    );

    bfr new_Jinkela_buffer_11707 (
        .din(new_Jinkela_wire_14120),
        .dout(new_Jinkela_wire_14121)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_2059),
        .dout(new_Jinkela_wire_2060)
    );

    bfr new_Jinkela_buffer_11776 (
        .din(new_Jinkela_wire_14207),
        .dout(new_Jinkela_wire_14208)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(new_Jinkela_wire_2001),
        .dout(new_Jinkela_wire_2002)
    );

    bfr new_Jinkela_buffer_11708 (
        .din(new_Jinkela_wire_14121),
        .dout(new_Jinkela_wire_14122)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_2255),
        .dout(new_Jinkela_wire_2256)
    );

    bfr new_Jinkela_buffer_11780 (
        .din(_1821_),
        .dout(new_Jinkela_wire_14216)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_2002),
        .dout(new_Jinkela_wire_2003)
    );

    bfr new_Jinkela_buffer_11709 (
        .din(new_Jinkela_wire_14122),
        .dout(new_Jinkela_wire_14123)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_2060),
        .dout(new_Jinkela_wire_2061)
    );

    bfr new_Jinkela_buffer_11777 (
        .din(new_Jinkela_wire_14208),
        .dout(new_Jinkela_wire_14209)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(new_Jinkela_wire_2003),
        .dout(new_Jinkela_wire_2004)
    );

    bfr new_Jinkela_buffer_11710 (
        .din(new_Jinkela_wire_14123),
        .dout(new_Jinkela_wire_14124)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_2160),
        .dout(new_Jinkela_wire_2161)
    );

    spl2 new_Jinkela_splitter_1068 (
        .a(_1830_),
        .b(new_Jinkela_wire_14259),
        .c(new_Jinkela_wire_14260)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_2004),
        .dout(new_Jinkela_wire_2005)
    );

    bfr new_Jinkela_buffer_11711 (
        .din(new_Jinkela_wire_14124),
        .dout(new_Jinkela_wire_14125)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(new_Jinkela_wire_2061),
        .dout(new_Jinkela_wire_2062)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_2005),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_11820 (
        .din(_1546_),
        .dout(new_Jinkela_wire_14258)
    );

    bfr new_Jinkela_buffer_11712 (
        .din(new_Jinkela_wire_14125),
        .dout(new_Jinkela_wire_14126)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(_1113_),
        .dout(new_Jinkela_wire_2314)
    );

    bfr new_Jinkela_buffer_11781 (
        .din(new_Jinkela_wire_14216),
        .dout(new_Jinkela_wire_14217)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_2006),
        .dout(new_Jinkela_wire_2007)
    );

    bfr new_Jinkela_buffer_11713 (
        .din(new_Jinkela_wire_14126),
        .dout(new_Jinkela_wire_14127)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_2062),
        .dout(new_Jinkela_wire_2063)
    );

    bfr new_Jinkela_buffer_11825 (
        .din(_0995_),
        .dout(new_Jinkela_wire_14265)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_2007),
        .dout(new_Jinkela_wire_2008)
    );

    bfr new_Jinkela_buffer_11821 (
        .din(new_Jinkela_wire_14260),
        .dout(new_Jinkela_wire_14261)
    );

    bfr new_Jinkela_buffer_11714 (
        .din(new_Jinkela_wire_14127),
        .dout(new_Jinkela_wire_14128)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(new_Jinkela_wire_2161),
        .dout(new_Jinkela_wire_2162)
    );

    bfr new_Jinkela_buffer_11782 (
        .din(new_Jinkela_wire_14217),
        .dout(new_Jinkela_wire_14218)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_2008),
        .dout(new_Jinkela_wire_2009)
    );

    bfr new_Jinkela_buffer_11715 (
        .din(new_Jinkela_wire_14128),
        .dout(new_Jinkela_wire_14129)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_2063),
        .dout(new_Jinkela_wire_2064)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_2009),
        .dout(new_Jinkela_wire_2010)
    );

    bfr new_Jinkela_buffer_11716 (
        .din(new_Jinkela_wire_14129),
        .dout(new_Jinkela_wire_14130)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_2262),
        .dout(new_Jinkela_wire_2263)
    );

    bfr new_Jinkela_buffer_11783 (
        .din(new_Jinkela_wire_14218),
        .dout(new_Jinkela_wire_14219)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(new_Jinkela_wire_2010),
        .b(new_Jinkela_wire_2011),
        .c(new_Jinkela_wire_2012)
    );

    bfr new_Jinkela_buffer_11717 (
        .din(new_Jinkela_wire_14130),
        .dout(new_Jinkela_wire_14131)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(new_Jinkela_wire_2162),
        .dout(new_Jinkela_wire_2163)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_2064),
        .dout(new_Jinkela_wire_2065)
    );

    spl2 new_Jinkela_splitter_1069 (
        .a(_0286_),
        .b(new_Jinkela_wire_14266),
        .c(new_Jinkela_wire_14267)
    );

    bfr new_Jinkela_buffer_11718 (
        .din(new_Jinkela_wire_14131),
        .dout(new_Jinkela_wire_14132)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(new_Jinkela_wire_2065),
        .dout(new_Jinkela_wire_2066)
    );

    bfr new_Jinkela_buffer_11784 (
        .din(new_Jinkela_wire_14219),
        .dout(new_Jinkela_wire_14220)
    );

    spl2 new_Jinkela_splitter_282 (
        .a(_1208_),
        .b(new_Jinkela_wire_2317),
        .c(new_Jinkela_wire_2318)
    );

    bfr new_Jinkela_buffer_11719 (
        .din(new_Jinkela_wire_14132),
        .dout(new_Jinkela_wire_14133)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_2066),
        .dout(new_Jinkela_wire_2067)
    );

    bfr new_Jinkela_buffer_11830 (
        .din(_0178_),
        .dout(new_Jinkela_wire_14272)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(new_Jinkela_wire_2163),
        .dout(new_Jinkela_wire_2164)
    );

    bfr new_Jinkela_buffer_11720 (
        .din(new_Jinkela_wire_14133),
        .dout(new_Jinkela_wire_14134)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(new_Jinkela_wire_2067),
        .dout(new_Jinkela_wire_2068)
    );

    bfr new_Jinkela_buffer_11785 (
        .din(new_Jinkela_wire_14220),
        .dout(new_Jinkela_wire_14221)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_Jinkela_wire_2263),
        .dout(new_Jinkela_wire_2264)
    );

    bfr new_Jinkela_buffer_11721 (
        .din(new_Jinkela_wire_14134),
        .dout(new_Jinkela_wire_14135)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(new_Jinkela_wire_2068),
        .dout(new_Jinkela_wire_2069)
    );

    bfr new_Jinkela_buffer_11822 (
        .din(new_Jinkela_wire_14261),
        .dout(new_Jinkela_wire_14262)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(new_Jinkela_wire_2164),
        .dout(new_Jinkela_wire_2165)
    );

    bfr new_Jinkela_buffer_11722 (
        .din(new_Jinkela_wire_14135),
        .dout(new_Jinkela_wire_14136)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(new_Jinkela_wire_2069),
        .dout(new_Jinkela_wire_2070)
    );

    bfr new_Jinkela_buffer_11786 (
        .din(new_Jinkela_wire_14221),
        .dout(new_Jinkela_wire_14222)
    );

    spl2 new_Jinkela_splitter_281 (
        .a(_1557_),
        .b(new_Jinkela_wire_2315),
        .c(new_Jinkela_wire_2316)
    );

    bfr new_Jinkela_buffer_11723 (
        .din(new_Jinkela_wire_14136),
        .dout(new_Jinkela_wire_14137)
    );

    bfr new_Jinkela_buffer_11826 (
        .din(new_Jinkela_wire_14267),
        .dout(new_Jinkela_wire_14268)
    );

    bfr new_Jinkela_buffer_11724 (
        .din(new_Jinkela_wire_14137),
        .dout(new_Jinkela_wire_14138)
    );

    bfr new_Jinkela_buffer_11787 (
        .din(new_Jinkela_wire_14222),
        .dout(new_Jinkela_wire_14223)
    );

    bfr new_Jinkela_buffer_11725 (
        .din(new_Jinkela_wire_14138),
        .dout(new_Jinkela_wire_14139)
    );

    bfr new_Jinkela_buffer_11823 (
        .din(new_Jinkela_wire_14262),
        .dout(new_Jinkela_wire_14263)
    );

    bfr new_Jinkela_buffer_11726 (
        .din(new_Jinkela_wire_14139),
        .dout(new_Jinkela_wire_14140)
    );

    bfr new_Jinkela_buffer_11788 (
        .din(new_Jinkela_wire_14223),
        .dout(new_Jinkela_wire_14224)
    );

    bfr new_Jinkela_buffer_11727 (
        .din(new_Jinkela_wire_14140),
        .dout(new_Jinkela_wire_14141)
    );

    bfr new_Jinkela_buffer_11831 (
        .din(_0740_),
        .dout(new_Jinkela_wire_14273)
    );

    bfr new_Jinkela_buffer_11728 (
        .din(new_Jinkela_wire_14141),
        .dout(new_Jinkela_wire_14142)
    );

    bfr new_Jinkela_buffer_11789 (
        .din(new_Jinkela_wire_14224),
        .dout(new_Jinkela_wire_14225)
    );

    bfr new_Jinkela_buffer_11729 (
        .din(new_Jinkela_wire_14142),
        .dout(new_Jinkela_wire_14143)
    );

    bfr new_Jinkela_buffer_11824 (
        .din(new_Jinkela_wire_14263),
        .dout(new_Jinkela_wire_14264)
    );

    bfr new_Jinkela_buffer_11730 (
        .din(new_Jinkela_wire_14143),
        .dout(new_Jinkela_wire_14144)
    );

    bfr new_Jinkela_buffer_11790 (
        .din(new_Jinkela_wire_14225),
        .dout(new_Jinkela_wire_14226)
    );

    bfr new_Jinkela_buffer_11731 (
        .din(new_Jinkela_wire_14144),
        .dout(new_Jinkela_wire_14145)
    );

    bfr new_Jinkela_buffer_11832 (
        .din(_0489_),
        .dout(new_Jinkela_wire_14274)
    );

    bfr new_Jinkela_buffer_11732 (
        .din(new_Jinkela_wire_14145),
        .dout(new_Jinkela_wire_14146)
    );

    bfr new_Jinkela_buffer_11791 (
        .din(new_Jinkela_wire_14226),
        .dout(new_Jinkela_wire_14227)
    );

    bfr new_Jinkela_buffer_11733 (
        .din(new_Jinkela_wire_14146),
        .dout(new_Jinkela_wire_14147)
    );

    bfr new_Jinkela_buffer_11827 (
        .din(new_Jinkela_wire_14268),
        .dout(new_Jinkela_wire_14269)
    );

    bfr new_Jinkela_buffer_11734 (
        .din(new_Jinkela_wire_14147),
        .dout(new_Jinkela_wire_14148)
    );

    bfr new_Jinkela_buffer_11792 (
        .din(new_Jinkela_wire_14227),
        .dout(new_Jinkela_wire_14228)
    );

    bfr new_Jinkela_buffer_11735 (
        .din(new_Jinkela_wire_14148),
        .dout(new_Jinkela_wire_14149)
    );

    spl2 new_Jinkela_splitter_1070 (
        .a(_1796_),
        .b(new_Jinkela_wire_14275),
        .c(new_Jinkela_wire_14276)
    );

    bfr new_Jinkela_buffer_11736 (
        .din(new_Jinkela_wire_14149),
        .dout(new_Jinkela_wire_14150)
    );

    bfr new_Jinkela_buffer_11793 (
        .din(new_Jinkela_wire_14228),
        .dout(new_Jinkela_wire_14229)
    );

    bfr new_Jinkela_buffer_11737 (
        .din(new_Jinkela_wire_14150),
        .dout(new_Jinkela_wire_14151)
    );

    bfr new_Jinkela_buffer_11828 (
        .din(new_Jinkela_wire_14269),
        .dout(new_Jinkela_wire_14270)
    );

    bfr new_Jinkela_buffer_11738 (
        .din(new_Jinkela_wire_14151),
        .dout(new_Jinkela_wire_14152)
    );

    bfr new_Jinkela_buffer_11794 (
        .din(new_Jinkela_wire_14229),
        .dout(new_Jinkela_wire_14230)
    );

    bfr new_Jinkela_buffer_11739 (
        .din(new_Jinkela_wire_14152),
        .dout(new_Jinkela_wire_14153)
    );

    spl2 new_Jinkela_splitter_1071 (
        .a(_0679_),
        .b(new_Jinkela_wire_14277),
        .c(new_Jinkela_wire_14278)
    );

    bfr new_Jinkela_buffer_11740 (
        .din(new_Jinkela_wire_14153),
        .dout(new_Jinkela_wire_14154)
    );

    bfr new_Jinkela_buffer_11795 (
        .din(new_Jinkela_wire_14230),
        .dout(new_Jinkela_wire_14231)
    );

    bfr new_Jinkela_buffer_11741 (
        .din(new_Jinkela_wire_14154),
        .dout(new_Jinkela_wire_14155)
    );

    bfr new_Jinkela_buffer_11829 (
        .din(new_Jinkela_wire_14270),
        .dout(new_Jinkela_wire_14271)
    );

    bfr new_Jinkela_buffer_11742 (
        .din(new_Jinkela_wire_14155),
        .dout(new_Jinkela_wire_14156)
    );

    bfr new_Jinkela_buffer_11796 (
        .din(new_Jinkela_wire_14231),
        .dout(new_Jinkela_wire_14232)
    );

    bfr new_Jinkela_buffer_11743 (
        .din(new_Jinkela_wire_14156),
        .dout(new_Jinkela_wire_14157)
    );

    spl2 new_Jinkela_splitter_1072 (
        .a(_0681_),
        .b(new_Jinkela_wire_14279),
        .c(new_Jinkela_wire_14280)
    );

    bfr new_Jinkela_buffer_4957 (
        .din(new_Jinkela_wire_6412),
        .dout(new_Jinkela_wire_6413)
    );

    bfr new_Jinkela_buffer_15223 (
        .din(new_Jinkela_wire_18157),
        .dout(new_Jinkela_wire_18158)
    );

    bfr new_Jinkela_buffer_4842 (
        .din(new_Jinkela_wire_6273),
        .dout(new_Jinkela_wire_6274)
    );

    bfr new_Jinkela_buffer_4774 (
        .din(new_Jinkela_wire_6187),
        .dout(new_Jinkela_wire_6188)
    );

    bfr new_Jinkela_buffer_15160 (
        .din(new_Jinkela_wire_18080),
        .dout(new_Jinkela_wire_18081)
    );

    bfr new_Jinkela_buffer_15346 (
        .din(_1119_),
        .dout(new_Jinkela_wire_18297)
    );

    bfr new_Jinkela_buffer_4775 (
        .din(new_Jinkela_wire_6188),
        .dout(new_Jinkela_wire_6189)
    );

    bfr new_Jinkela_buffer_15161 (
        .din(new_Jinkela_wire_18081),
        .dout(new_Jinkela_wire_18082)
    );

    bfr new_Jinkela_buffer_4938 (
        .din(new_Jinkela_wire_6383),
        .dout(new_Jinkela_wire_6384)
    );

    bfr new_Jinkela_buffer_15224 (
        .din(new_Jinkela_wire_18158),
        .dout(new_Jinkela_wire_18159)
    );

    bfr new_Jinkela_buffer_4843 (
        .din(new_Jinkela_wire_6274),
        .dout(new_Jinkela_wire_6275)
    );

    bfr new_Jinkela_buffer_4776 (
        .din(new_Jinkela_wire_6189),
        .dout(new_Jinkela_wire_6190)
    );

    bfr new_Jinkela_buffer_15162 (
        .din(new_Jinkela_wire_18082),
        .dout(new_Jinkela_wire_18083)
    );

    bfr new_Jinkela_buffer_15302 (
        .din(new_Jinkela_wire_18242),
        .dout(new_Jinkela_wire_18243)
    );

    spl2 new_Jinkela_splitter_556 (
        .a(new_Jinkela_wire_6190),
        .b(new_Jinkela_wire_6191),
        .c(new_Jinkela_wire_6192)
    );

    bfr new_Jinkela_buffer_15163 (
        .din(new_Jinkela_wire_18083),
        .dout(new_Jinkela_wire_18084)
    );

    bfr new_Jinkela_buffer_15225 (
        .din(new_Jinkela_wire_18159),
        .dout(new_Jinkela_wire_18160)
    );

    spl2 new_Jinkela_splitter_578 (
        .a(_1671_),
        .b(new_Jinkela_wire_6419),
        .c(new_Jinkela_wire_6420)
    );

    bfr new_Jinkela_buffer_15164 (
        .din(new_Jinkela_wire_18084),
        .dout(new_Jinkela_wire_18085)
    );

    bfr new_Jinkela_buffer_4844 (
        .din(new_Jinkela_wire_6275),
        .dout(new_Jinkela_wire_6276)
    );

    bfr new_Jinkela_buffer_4939 (
        .din(new_Jinkela_wire_6384),
        .dout(new_Jinkela_wire_6385)
    );

    bfr new_Jinkela_buffer_15348 (
        .din(_1577_),
        .dout(new_Jinkela_wire_18299)
    );

    bfr new_Jinkela_buffer_4845 (
        .din(new_Jinkela_wire_6276),
        .dout(new_Jinkela_wire_6277)
    );

    bfr new_Jinkela_buffer_15165 (
        .din(new_Jinkela_wire_18085),
        .dout(new_Jinkela_wire_18086)
    );

    bfr new_Jinkela_buffer_15226 (
        .din(new_Jinkela_wire_18160),
        .dout(new_Jinkela_wire_18161)
    );

    bfr new_Jinkela_buffer_4846 (
        .din(new_Jinkela_wire_6277),
        .dout(new_Jinkela_wire_6278)
    );

    bfr new_Jinkela_buffer_15166 (
        .din(new_Jinkela_wire_18086),
        .dout(new_Jinkela_wire_18087)
    );

    bfr new_Jinkela_buffer_4940 (
        .din(new_Jinkela_wire_6385),
        .dout(new_Jinkela_wire_6386)
    );

    bfr new_Jinkela_buffer_15303 (
        .din(new_Jinkela_wire_18243),
        .dout(new_Jinkela_wire_18244)
    );

    bfr new_Jinkela_buffer_4847 (
        .din(new_Jinkela_wire_6278),
        .dout(new_Jinkela_wire_6279)
    );

    bfr new_Jinkela_buffer_15167 (
        .din(new_Jinkela_wire_18087),
        .dout(new_Jinkela_wire_18088)
    );

    bfr new_Jinkela_buffer_4958 (
        .din(new_Jinkela_wire_6413),
        .dout(new_Jinkela_wire_6414)
    );

    bfr new_Jinkela_buffer_15227 (
        .din(new_Jinkela_wire_18161),
        .dout(new_Jinkela_wire_18162)
    );

    bfr new_Jinkela_buffer_4848 (
        .din(new_Jinkela_wire_6279),
        .dout(new_Jinkela_wire_6280)
    );

    bfr new_Jinkela_buffer_15168 (
        .din(new_Jinkela_wire_18088),
        .dout(new_Jinkela_wire_18089)
    );

    bfr new_Jinkela_buffer_4941 (
        .din(new_Jinkela_wire_6386),
        .dout(new_Jinkela_wire_6387)
    );

    bfr new_Jinkela_buffer_4849 (
        .din(new_Jinkela_wire_6280),
        .dout(new_Jinkela_wire_6281)
    );

    bfr new_Jinkela_buffer_15347 (
        .din(_0938_),
        .dout(new_Jinkela_wire_18298)
    );

    bfr new_Jinkela_buffer_15169 (
        .din(new_Jinkela_wire_18089),
        .dout(new_Jinkela_wire_18090)
    );

    bfr new_Jinkela_buffer_15228 (
        .din(new_Jinkela_wire_18162),
        .dout(new_Jinkela_wire_18163)
    );

    bfr new_Jinkela_buffer_4850 (
        .din(new_Jinkela_wire_6281),
        .dout(new_Jinkela_wire_6282)
    );

    bfr new_Jinkela_buffer_15170 (
        .din(new_Jinkela_wire_18090),
        .dout(new_Jinkela_wire_18091)
    );

    bfr new_Jinkela_buffer_4961 (
        .din(_1167_),
        .dout(new_Jinkela_wire_6421)
    );

    bfr new_Jinkela_buffer_4942 (
        .din(new_Jinkela_wire_6387),
        .dout(new_Jinkela_wire_6388)
    );

    bfr new_Jinkela_buffer_15304 (
        .din(new_Jinkela_wire_18244),
        .dout(new_Jinkela_wire_18245)
    );

    bfr new_Jinkela_buffer_4851 (
        .din(new_Jinkela_wire_6282),
        .dout(new_Jinkela_wire_6283)
    );

    bfr new_Jinkela_buffer_15171 (
        .din(new_Jinkela_wire_18091),
        .dout(new_Jinkela_wire_18092)
    );

    bfr new_Jinkela_buffer_4959 (
        .din(new_Jinkela_wire_6414),
        .dout(new_Jinkela_wire_6415)
    );

    bfr new_Jinkela_buffer_15229 (
        .din(new_Jinkela_wire_18163),
        .dout(new_Jinkela_wire_18164)
    );

    bfr new_Jinkela_buffer_4852 (
        .din(new_Jinkela_wire_6283),
        .dout(new_Jinkela_wire_6284)
    );

    bfr new_Jinkela_buffer_15172 (
        .din(new_Jinkela_wire_18092),
        .dout(new_Jinkela_wire_18093)
    );

    bfr new_Jinkela_buffer_4943 (
        .din(new_Jinkela_wire_6388),
        .dout(new_Jinkela_wire_6389)
    );

    spl2 new_Jinkela_splitter_1325 (
        .a(_0946_),
        .b(new_Jinkela_wire_18309),
        .c(new_Jinkela_wire_18310)
    );

    bfr new_Jinkela_buffer_4853 (
        .din(new_Jinkela_wire_6284),
        .dout(new_Jinkela_wire_6285)
    );

    bfr new_Jinkela_buffer_15173 (
        .din(new_Jinkela_wire_18093),
        .dout(new_Jinkela_wire_18094)
    );

    spl2 new_Jinkela_splitter_580 (
        .a(_1583_),
        .b(new_Jinkela_wire_6512),
        .c(new_Jinkela_wire_6513)
    );

    bfr new_Jinkela_buffer_15230 (
        .din(new_Jinkela_wire_18164),
        .dout(new_Jinkela_wire_18165)
    );

    bfr new_Jinkela_buffer_4854 (
        .din(new_Jinkela_wire_6285),
        .dout(new_Jinkela_wire_6286)
    );

    bfr new_Jinkela_buffer_15174 (
        .din(new_Jinkela_wire_18094),
        .dout(new_Jinkela_wire_18095)
    );

    bfr new_Jinkela_buffer_4962 (
        .din(_0218_),
        .dout(new_Jinkela_wire_6422)
    );

    bfr new_Jinkela_buffer_4944 (
        .din(new_Jinkela_wire_6389),
        .dout(new_Jinkela_wire_6390)
    );

    bfr new_Jinkela_buffer_15305 (
        .din(new_Jinkela_wire_18245),
        .dout(new_Jinkela_wire_18246)
    );

    bfr new_Jinkela_buffer_4855 (
        .din(new_Jinkela_wire_6286),
        .dout(new_Jinkela_wire_6287)
    );

    bfr new_Jinkela_buffer_15175 (
        .din(new_Jinkela_wire_18095),
        .dout(new_Jinkela_wire_18096)
    );

    bfr new_Jinkela_buffer_4960 (
        .din(new_Jinkela_wire_6415),
        .dout(new_Jinkela_wire_6416)
    );

    bfr new_Jinkela_buffer_15231 (
        .din(new_Jinkela_wire_18165),
        .dout(new_Jinkela_wire_18166)
    );

    bfr new_Jinkela_buffer_4856 (
        .din(new_Jinkela_wire_6287),
        .dout(new_Jinkela_wire_6288)
    );

    bfr new_Jinkela_buffer_15176 (
        .din(new_Jinkela_wire_18096),
        .dout(new_Jinkela_wire_18097)
    );

    bfr new_Jinkela_buffer_4945 (
        .din(new_Jinkela_wire_6390),
        .dout(new_Jinkela_wire_6391)
    );

    bfr new_Jinkela_buffer_4857 (
        .din(new_Jinkela_wire_6288),
        .dout(new_Jinkela_wire_6289)
    );

    bfr new_Jinkela_buffer_15360 (
        .din(_0710_),
        .dout(new_Jinkela_wire_18315)
    );

    bfr new_Jinkela_buffer_15177 (
        .din(new_Jinkela_wire_18097),
        .dout(new_Jinkela_wire_18098)
    );

    bfr new_Jinkela_buffer_15232 (
        .din(new_Jinkela_wire_18166),
        .dout(new_Jinkela_wire_18167)
    );

    bfr new_Jinkela_buffer_4858 (
        .din(new_Jinkela_wire_6289),
        .dout(new_Jinkela_wire_6290)
    );

    bfr new_Jinkela_buffer_15178 (
        .din(new_Jinkela_wire_18098),
        .dout(new_Jinkela_wire_18099)
    );

    spl2 new_Jinkela_splitter_581 (
        .a(_0893_),
        .b(new_Jinkela_wire_6514),
        .c(new_Jinkela_wire_6515)
    );

    bfr new_Jinkela_buffer_4946 (
        .din(new_Jinkela_wire_6391),
        .dout(new_Jinkela_wire_6392)
    );

    bfr new_Jinkela_buffer_15306 (
        .din(new_Jinkela_wire_18246),
        .dout(new_Jinkela_wire_18247)
    );

    bfr new_Jinkela_buffer_4859 (
        .din(new_Jinkela_wire_6290),
        .dout(new_Jinkela_wire_6291)
    );

    bfr new_Jinkela_buffer_15179 (
        .din(new_Jinkela_wire_18099),
        .dout(new_Jinkela_wire_18100)
    );

    bfr new_Jinkela_buffer_4963 (
        .din(new_Jinkela_wire_6422),
        .dout(new_Jinkela_wire_6423)
    );

    bfr new_Jinkela_buffer_15233 (
        .din(new_Jinkela_wire_18167),
        .dout(new_Jinkela_wire_18168)
    );

    bfr new_Jinkela_buffer_4860 (
        .din(new_Jinkela_wire_6291),
        .dout(new_Jinkela_wire_6292)
    );

    spl2 new_Jinkela_splitter_1309 (
        .a(new_Jinkela_wire_18100),
        .b(new_Jinkela_wire_18101),
        .c(new_Jinkela_wire_18102)
    );

    bfr new_Jinkela_buffer_8295 (
        .din(new_Jinkela_wire_10222),
        .dout(new_Jinkela_wire_10223)
    );

    bfr new_Jinkela_buffer_8273 (
        .din(new_Jinkela_wire_10196),
        .dout(new_Jinkela_wire_10197)
    );

    bfr new_Jinkela_buffer_8333 (
        .din(new_Jinkela_wire_10270),
        .dout(new_Jinkela_wire_10271)
    );

    bfr new_Jinkela_buffer_8274 (
        .din(new_Jinkela_wire_10197),
        .dout(new_Jinkela_wire_10198)
    );

    bfr new_Jinkela_buffer_8296 (
        .din(new_Jinkela_wire_10223),
        .dout(new_Jinkela_wire_10224)
    );

    bfr new_Jinkela_buffer_8275 (
        .din(new_Jinkela_wire_10198),
        .dout(new_Jinkela_wire_10199)
    );

    bfr new_Jinkela_buffer_8339 (
        .din(new_Jinkela_wire_10280),
        .dout(new_Jinkela_wire_10281)
    );

    bfr new_Jinkela_buffer_8276 (
        .din(new_Jinkela_wire_10199),
        .dout(new_Jinkela_wire_10200)
    );

    bfr new_Jinkela_buffer_8297 (
        .din(new_Jinkela_wire_10224),
        .dout(new_Jinkela_wire_10225)
    );

    bfr new_Jinkela_buffer_8277 (
        .din(new_Jinkela_wire_10200),
        .dout(new_Jinkela_wire_10201)
    );

    bfr new_Jinkela_buffer_8334 (
        .din(new_Jinkela_wire_10271),
        .dout(new_Jinkela_wire_10272)
    );

    spl2 new_Jinkela_splitter_811 (
        .a(new_Jinkela_wire_10201),
        .b(new_Jinkela_wire_10202),
        .c(new_Jinkela_wire_10203)
    );

    spl2 new_Jinkela_splitter_822 (
        .a(_0435_),
        .b(new_Jinkela_wire_10397),
        .c(new_Jinkela_wire_10398)
    );

    bfr new_Jinkela_buffer_8298 (
        .din(new_Jinkela_wire_10225),
        .dout(new_Jinkela_wire_10226)
    );

    bfr new_Jinkela_buffer_8299 (
        .din(new_Jinkela_wire_10226),
        .dout(new_Jinkela_wire_10227)
    );

    spl2 new_Jinkela_splitter_818 (
        .a(new_Jinkela_wire_10272),
        .b(new_Jinkela_wire_10273),
        .c(new_Jinkela_wire_10274)
    );

    bfr new_Jinkela_buffer_8300 (
        .din(new_Jinkela_wire_10227),
        .dout(new_Jinkela_wire_10228)
    );

    bfr new_Jinkela_buffer_8301 (
        .din(new_Jinkela_wire_10228),
        .dout(new_Jinkela_wire_10229)
    );

    bfr new_Jinkela_buffer_8340 (
        .din(new_Jinkela_wire_10281),
        .dout(new_Jinkela_wire_10282)
    );

    bfr new_Jinkela_buffer_8302 (
        .din(new_Jinkela_wire_10229),
        .dout(new_Jinkela_wire_10230)
    );

    bfr new_Jinkela_buffer_8341 (
        .din(new_Jinkela_wire_10282),
        .dout(new_Jinkela_wire_10283)
    );

    bfr new_Jinkela_buffer_8303 (
        .din(new_Jinkela_wire_10230),
        .dout(new_Jinkela_wire_10231)
    );

    spl2 new_Jinkela_splitter_823 (
        .a(_0918_),
        .b(new_Jinkela_wire_10399),
        .c(new_Jinkela_wire_10400)
    );

    bfr new_Jinkela_buffer_8304 (
        .din(new_Jinkela_wire_10231),
        .dout(new_Jinkela_wire_10232)
    );

    bfr new_Jinkela_buffer_8342 (
        .din(new_Jinkela_wire_10283),
        .dout(new_Jinkela_wire_10284)
    );

    bfr new_Jinkela_buffer_8305 (
        .din(new_Jinkela_wire_10232),
        .dout(new_Jinkela_wire_10233)
    );

    bfr new_Jinkela_buffer_8491 (
        .din(_0033_),
        .dout(new_Jinkela_wire_10441)
    );

    bfr new_Jinkela_buffer_8306 (
        .din(new_Jinkela_wire_10233),
        .dout(new_Jinkela_wire_10234)
    );

    bfr new_Jinkela_buffer_8343 (
        .din(new_Jinkela_wire_10284),
        .dout(new_Jinkela_wire_10285)
    );

    bfr new_Jinkela_buffer_8307 (
        .din(new_Jinkela_wire_10234),
        .dout(new_Jinkela_wire_10235)
    );

    bfr new_Jinkela_buffer_8451 (
        .din(new_Jinkela_wire_10400),
        .dout(new_Jinkela_wire_10401)
    );

    bfr new_Jinkela_buffer_8499 (
        .din(_0774_),
        .dout(new_Jinkela_wire_10451)
    );

    bfr new_Jinkela_buffer_8308 (
        .din(new_Jinkela_wire_10235),
        .dout(new_Jinkela_wire_10236)
    );

    bfr new_Jinkela_buffer_8344 (
        .din(new_Jinkela_wire_10285),
        .dout(new_Jinkela_wire_10286)
    );

    bfr new_Jinkela_buffer_8309 (
        .din(new_Jinkela_wire_10236),
        .dout(new_Jinkela_wire_10237)
    );

    bfr new_Jinkela_buffer_8500 (
        .din(_0619_),
        .dout(new_Jinkela_wire_10452)
    );

    bfr new_Jinkela_buffer_8310 (
        .din(new_Jinkela_wire_10237),
        .dout(new_Jinkela_wire_10238)
    );

    bfr new_Jinkela_buffer_8345 (
        .din(new_Jinkela_wire_10286),
        .dout(new_Jinkela_wire_10287)
    );

    bfr new_Jinkela_buffer_8311 (
        .din(new_Jinkela_wire_10238),
        .dout(new_Jinkela_wire_10239)
    );

    bfr new_Jinkela_buffer_8452 (
        .din(new_Jinkela_wire_10401),
        .dout(new_Jinkela_wire_10402)
    );

    bfr new_Jinkela_buffer_8312 (
        .din(new_Jinkela_wire_10239),
        .dout(new_Jinkela_wire_10240)
    );

    bfr new_Jinkela_buffer_8346 (
        .din(new_Jinkela_wire_10287),
        .dout(new_Jinkela_wire_10288)
    );

    bfr new_Jinkela_buffer_11744 (
        .din(new_Jinkela_wire_14157),
        .dout(new_Jinkela_wire_14158)
    );

    bfr new_Jinkela_buffer_11797 (
        .din(new_Jinkela_wire_14232),
        .dout(new_Jinkela_wire_14233)
    );

    bfr new_Jinkela_buffer_11745 (
        .din(new_Jinkela_wire_14158),
        .dout(new_Jinkela_wire_14159)
    );

    bfr new_Jinkela_buffer_11746 (
        .din(new_Jinkela_wire_14159),
        .dout(new_Jinkela_wire_14160)
    );

    bfr new_Jinkela_buffer_11798 (
        .din(new_Jinkela_wire_14233),
        .dout(new_Jinkela_wire_14234)
    );

    bfr new_Jinkela_buffer_11747 (
        .din(new_Jinkela_wire_14160),
        .dout(new_Jinkela_wire_14161)
    );

    spl2 new_Jinkela_splitter_1073 (
        .a(_1245_),
        .b(new_Jinkela_wire_14281),
        .c(new_Jinkela_wire_14282)
    );

    bfr new_Jinkela_buffer_11748 (
        .din(new_Jinkela_wire_14161),
        .dout(new_Jinkela_wire_14162)
    );

    bfr new_Jinkela_buffer_11799 (
        .din(new_Jinkela_wire_14234),
        .dout(new_Jinkela_wire_14235)
    );

    bfr new_Jinkela_buffer_11749 (
        .din(new_Jinkela_wire_14162),
        .dout(new_Jinkela_wire_14163)
    );

    bfr new_Jinkela_buffer_11833 (
        .din(_0614_),
        .dout(new_Jinkela_wire_14283)
    );

    bfr new_Jinkela_buffer_11750 (
        .din(new_Jinkela_wire_14163),
        .dout(new_Jinkela_wire_14164)
    );

    bfr new_Jinkela_buffer_11800 (
        .din(new_Jinkela_wire_14235),
        .dout(new_Jinkela_wire_14236)
    );

    bfr new_Jinkela_buffer_11751 (
        .din(new_Jinkela_wire_14164),
        .dout(new_Jinkela_wire_14165)
    );

    spl2 new_Jinkela_splitter_1075 (
        .a(_0397_),
        .b(new_Jinkela_wire_14286),
        .c(new_Jinkela_wire_14287)
    );

    spl2 new_Jinkela_splitter_1074 (
        .a(_1502_),
        .b(new_Jinkela_wire_14284),
        .c(new_Jinkela_wire_14285)
    );

    bfr new_Jinkela_buffer_11752 (
        .din(new_Jinkela_wire_14165),
        .dout(new_Jinkela_wire_14166)
    );

    bfr new_Jinkela_buffer_11801 (
        .din(new_Jinkela_wire_14236),
        .dout(new_Jinkela_wire_14237)
    );

    bfr new_Jinkela_buffer_11753 (
        .din(new_Jinkela_wire_14166),
        .dout(new_Jinkela_wire_14167)
    );

    bfr new_Jinkela_buffer_11754 (
        .din(new_Jinkela_wire_14167),
        .dout(new_Jinkela_wire_14168)
    );

    bfr new_Jinkela_buffer_11802 (
        .din(new_Jinkela_wire_14237),
        .dout(new_Jinkela_wire_14238)
    );

    bfr new_Jinkela_buffer_11755 (
        .din(new_Jinkela_wire_14168),
        .dout(new_Jinkela_wire_14169)
    );

    bfr new_Jinkela_buffer_11834 (
        .din(_0023_),
        .dout(new_Jinkela_wire_14288)
    );

    bfr new_Jinkela_buffer_11756 (
        .din(new_Jinkela_wire_14169),
        .dout(new_Jinkela_wire_14170)
    );

    bfr new_Jinkela_buffer_11803 (
        .din(new_Jinkela_wire_14238),
        .dout(new_Jinkela_wire_14239)
    );

    bfr new_Jinkela_buffer_11757 (
        .din(new_Jinkela_wire_14170),
        .dout(new_Jinkela_wire_14171)
    );

    spl2 new_Jinkela_splitter_1077 (
        .a(_1015_),
        .b(new_Jinkela_wire_14299),
        .c(new_Jinkela_wire_14300)
    );

    bfr new_Jinkela_buffer_11835 (
        .din(_1296_),
        .dout(new_Jinkela_wire_14289)
    );

    bfr new_Jinkela_buffer_11758 (
        .din(new_Jinkela_wire_14171),
        .dout(new_Jinkela_wire_14172)
    );

    bfr new_Jinkela_buffer_11804 (
        .din(new_Jinkela_wire_14239),
        .dout(new_Jinkela_wire_14240)
    );

    bfr new_Jinkela_buffer_11759 (
        .din(new_Jinkela_wire_14172),
        .dout(new_Jinkela_wire_14173)
    );

    spl2 new_Jinkela_splitter_1078 (
        .a(_0550_),
        .b(new_Jinkela_wire_14301),
        .c(new_Jinkela_wire_14302)
    );

    bfr new_Jinkela_buffer_11760 (
        .din(new_Jinkela_wire_14173),
        .dout(new_Jinkela_wire_14174)
    );

    bfr new_Jinkela_buffer_11805 (
        .din(new_Jinkela_wire_14240),
        .dout(new_Jinkela_wire_14241)
    );

    bfr new_Jinkela_buffer_11761 (
        .din(new_Jinkela_wire_14174),
        .dout(new_Jinkela_wire_14175)
    );

    bfr new_Jinkela_buffer_11836 (
        .din(new_Jinkela_wire_14289),
        .dout(new_Jinkela_wire_14290)
    );

    bfr new_Jinkela_buffer_11762 (
        .din(new_Jinkela_wire_14175),
        .dout(new_Jinkela_wire_14176)
    );

    bfr new_Jinkela_buffer_11806 (
        .din(new_Jinkela_wire_14241),
        .dout(new_Jinkela_wire_14242)
    );

    bfr new_Jinkela_buffer_11763 (
        .din(new_Jinkela_wire_14176),
        .dout(new_Jinkela_wire_14177)
    );

    spl2 new_Jinkela_splitter_1079 (
        .a(_1141_),
        .b(new_Jinkela_wire_14307),
        .c(new_Jinkela_wire_14308)
    );

    bfr new_Jinkela_buffer_11764 (
        .din(new_Jinkela_wire_14177),
        .dout(new_Jinkela_wire_14178)
    );

    bfr new_Jinkela_buffer_11807 (
        .din(new_Jinkela_wire_14242),
        .dout(new_Jinkela_wire_14243)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_2070),
        .dout(new_Jinkela_wire_2071)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_2165),
        .dout(new_Jinkela_wire_2166)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(new_Jinkela_wire_2071),
        .dout(new_Jinkela_wire_2072)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_2264),
        .dout(new_Jinkela_wire_2265)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_2072),
        .dout(new_Jinkela_wire_2073)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(new_Jinkela_wire_2166),
        .dout(new_Jinkela_wire_2167)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_2073),
        .dout(new_Jinkela_wire_2074)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(new_Jinkela_wire_2320),
        .dout(new_Jinkela_wire_2321)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_2074),
        .dout(new_Jinkela_wire_2075)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_2167),
        .dout(new_Jinkela_wire_2168)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(new_Jinkela_wire_2075),
        .dout(new_Jinkela_wire_2076)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_2265),
        .dout(new_Jinkela_wire_2266)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_2076),
        .dout(new_Jinkela_wire_2077)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_2168),
        .dout(new_Jinkela_wire_2169)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(new_Jinkela_wire_2077),
        .dout(new_Jinkela_wire_2078)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(_0194_),
        .dout(new_Jinkela_wire_2319)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_2078),
        .dout(new_Jinkela_wire_2079)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(new_Jinkela_wire_2169),
        .dout(new_Jinkela_wire_2170)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_2079),
        .dout(new_Jinkela_wire_2080)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_2266),
        .dout(new_Jinkela_wire_2267)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_2080),
        .dout(new_Jinkela_wire_2081)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(new_Jinkela_wire_2170),
        .dout(new_Jinkela_wire_2171)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_2081),
        .dout(new_Jinkela_wire_2082)
    );

    spl2 new_Jinkela_splitter_284 (
        .a(_0708_),
        .b(new_Jinkela_wire_2324),
        .c(new_Jinkela_wire_2325)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(_0945_),
        .dout(new_Jinkela_wire_2320)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_2082),
        .dout(new_Jinkela_wire_2083)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_2171),
        .dout(new_Jinkela_wire_2172)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(new_Jinkela_wire_2083),
        .dout(new_Jinkela_wire_2084)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_2267),
        .dout(new_Jinkela_wire_2268)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_2084),
        .dout(new_Jinkela_wire_2085)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_2172),
        .dout(new_Jinkela_wire_2173)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_2085),
        .dout(new_Jinkela_wire_2086)
    );

    spl2 new_Jinkela_splitter_285 (
        .a(_0781_),
        .b(new_Jinkela_wire_2326),
        .c(new_Jinkela_wire_2327)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(new_Jinkela_wire_2086),
        .dout(new_Jinkela_wire_2087)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(new_Jinkela_wire_2173),
        .dout(new_Jinkela_wire_2174)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_2087),
        .dout(new_Jinkela_wire_2088)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_2268),
        .dout(new_Jinkela_wire_2269)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_2088),
        .dout(new_Jinkela_wire_2089)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_2174),
        .dout(new_Jinkela_wire_2175)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(new_Jinkela_wire_2089),
        .dout(new_Jinkela_wire_2090)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(new_Jinkela_wire_2090),
        .dout(new_Jinkela_wire_2091)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(new_Jinkela_wire_2175),
        .dout(new_Jinkela_wire_2176)
    );

    bfr new_Jinkela_buffer_11765 (
        .din(new_Jinkela_wire_14178),
        .dout(new_Jinkela_wire_14179)
    );

    bfr new_Jinkela_buffer_11837 (
        .din(new_Jinkela_wire_14290),
        .dout(new_Jinkela_wire_14291)
    );

    bfr new_Jinkela_buffer_11766 (
        .din(new_Jinkela_wire_14179),
        .dout(new_Jinkela_wire_14180)
    );

    bfr new_Jinkela_buffer_11808 (
        .din(new_Jinkela_wire_14243),
        .dout(new_Jinkela_wire_14244)
    );

    bfr new_Jinkela_buffer_11767 (
        .din(new_Jinkela_wire_14180),
        .dout(new_Jinkela_wire_14181)
    );

    bfr new_Jinkela_buffer_11843 (
        .din(new_Jinkela_wire_14302),
        .dout(new_Jinkela_wire_14303)
    );

    spl2 new_Jinkela_splitter_1056 (
        .a(new_Jinkela_wire_14181),
        .b(new_Jinkela_wire_14182),
        .c(new_Jinkela_wire_14183)
    );

    bfr new_Jinkela_buffer_11838 (
        .din(new_Jinkela_wire_14291),
        .dout(new_Jinkela_wire_14292)
    );

    bfr new_Jinkela_buffer_11809 (
        .din(new_Jinkela_wire_14244),
        .dout(new_Jinkela_wire_14245)
    );

    bfr new_Jinkela_buffer_11810 (
        .din(new_Jinkela_wire_14245),
        .dout(new_Jinkela_wire_14246)
    );

    bfr new_Jinkela_buffer_11847 (
        .din(_0737_),
        .dout(new_Jinkela_wire_14309)
    );

    bfr new_Jinkela_buffer_11811 (
        .din(new_Jinkela_wire_14246),
        .dout(new_Jinkela_wire_14247)
    );

    bfr new_Jinkela_buffer_11839 (
        .din(new_Jinkela_wire_14292),
        .dout(new_Jinkela_wire_14293)
    );

    bfr new_Jinkela_buffer_11812 (
        .din(new_Jinkela_wire_14247),
        .dout(new_Jinkela_wire_14248)
    );

    spl2 new_Jinkela_splitter_1080 (
        .a(_0385_),
        .b(new_Jinkela_wire_14311),
        .c(new_Jinkela_wire_14312)
    );

    bfr new_Jinkela_buffer_11813 (
        .din(new_Jinkela_wire_14248),
        .dout(new_Jinkela_wire_14249)
    );

    bfr new_Jinkela_buffer_11840 (
        .din(new_Jinkela_wire_14293),
        .dout(new_Jinkela_wire_14294)
    );

    bfr new_Jinkela_buffer_11814 (
        .din(new_Jinkela_wire_14249),
        .dout(new_Jinkela_wire_14250)
    );

    bfr new_Jinkela_buffer_11844 (
        .din(new_Jinkela_wire_14303),
        .dout(new_Jinkela_wire_14304)
    );

    bfr new_Jinkela_buffer_11815 (
        .din(new_Jinkela_wire_14250),
        .dout(new_Jinkela_wire_14251)
    );

    bfr new_Jinkela_buffer_11841 (
        .din(new_Jinkela_wire_14294),
        .dout(new_Jinkela_wire_14295)
    );

    bfr new_Jinkela_buffer_11816 (
        .din(new_Jinkela_wire_14251),
        .dout(new_Jinkela_wire_14252)
    );

    bfr new_Jinkela_buffer_11848 (
        .din(_1182_),
        .dout(new_Jinkela_wire_14310)
    );

    bfr new_Jinkela_buffer_11817 (
        .din(new_Jinkela_wire_14252),
        .dout(new_Jinkela_wire_14253)
    );

    bfr new_Jinkela_buffer_11842 (
        .din(new_Jinkela_wire_14295),
        .dout(new_Jinkela_wire_14296)
    );

    bfr new_Jinkela_buffer_11818 (
        .din(new_Jinkela_wire_14253),
        .dout(new_Jinkela_wire_14254)
    );

    bfr new_Jinkela_buffer_11845 (
        .din(new_Jinkela_wire_14304),
        .dout(new_Jinkela_wire_14305)
    );

    bfr new_Jinkela_buffer_11819 (
        .din(new_Jinkela_wire_14254),
        .dout(new_Jinkela_wire_14255)
    );

    spl2 new_Jinkela_splitter_1076 (
        .a(new_Jinkela_wire_14296),
        .b(new_Jinkela_wire_14297),
        .c(new_Jinkela_wire_14298)
    );

    spl2 new_Jinkela_splitter_1067 (
        .a(new_Jinkela_wire_14255),
        .b(new_Jinkela_wire_14256),
        .c(new_Jinkela_wire_14257)
    );

    spl2 new_Jinkela_splitter_1081 (
        .a(_0797_),
        .b(new_Jinkela_wire_14317),
        .c(new_Jinkela_wire_14318)
    );

    bfr new_Jinkela_buffer_11849 (
        .din(new_Jinkela_wire_14312),
        .dout(new_Jinkela_wire_14313)
    );

    bfr new_Jinkela_buffer_11846 (
        .din(new_Jinkela_wire_14305),
        .dout(new_Jinkela_wire_14306)
    );

    spl2 new_Jinkela_splitter_1082 (
        .a(_1411_),
        .b(new_Jinkela_wire_14319),
        .c(new_Jinkela_wire_14320)
    );

    bfr new_Jinkela_buffer_11850 (
        .din(new_Jinkela_wire_14313),
        .dout(new_Jinkela_wire_14314)
    );

    spl2 new_Jinkela_splitter_1083 (
        .a(_1162_),
        .b(new_Jinkela_wire_14325),
        .c(new_Jinkela_wire_14326)
    );

    bfr new_Jinkela_buffer_11851 (
        .din(new_Jinkela_wire_14314),
        .dout(new_Jinkela_wire_14315)
    );

    bfr new_Jinkela_buffer_11853 (
        .din(new_Jinkela_wire_14320),
        .dout(new_Jinkela_wire_14321)
    );

    bfr new_Jinkela_buffer_11857 (
        .din(_1170_),
        .dout(new_Jinkela_wire_14327)
    );

    bfr new_Jinkela_buffer_11852 (
        .din(new_Jinkela_wire_14315),
        .dout(new_Jinkela_wire_14316)
    );

    spl2 new_Jinkela_splitter_1084 (
        .a(_0198_),
        .b(new_Jinkela_wire_14328),
        .c(new_Jinkela_wire_14329)
    );

    bfr new_Jinkela_buffer_11854 (
        .din(new_Jinkela_wire_14321),
        .dout(new_Jinkela_wire_14322)
    );

    bfr new_Jinkela_buffer_8313 (
        .din(new_Jinkela_wire_10240),
        .dout(new_Jinkela_wire_10241)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(new_Jinkela_wire_2091),
        .dout(new_Jinkela_wire_2092)
    );

    bfr new_Jinkela_buffer_8492 (
        .din(new_Jinkela_wire_10441),
        .dout(new_Jinkela_wire_10442)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(new_Jinkela_wire_2269),
        .dout(new_Jinkela_wire_2270)
    );

    bfr new_Jinkela_buffer_8314 (
        .din(new_Jinkela_wire_10241),
        .dout(new_Jinkela_wire_10242)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_2092),
        .dout(new_Jinkela_wire_2093)
    );

    bfr new_Jinkela_buffer_8347 (
        .din(new_Jinkela_wire_10288),
        .dout(new_Jinkela_wire_10289)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_2176),
        .dout(new_Jinkela_wire_2177)
    );

    bfr new_Jinkela_buffer_8315 (
        .din(new_Jinkela_wire_10242),
        .dout(new_Jinkela_wire_10243)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_2093),
        .dout(new_Jinkela_wire_2094)
    );

    bfr new_Jinkela_buffer_8453 (
        .din(new_Jinkela_wire_10402),
        .dout(new_Jinkela_wire_10403)
    );

    bfr new_Jinkela_buffer_8316 (
        .din(new_Jinkela_wire_10243),
        .dout(new_Jinkela_wire_10244)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_2094),
        .dout(new_Jinkela_wire_2095)
    );

    bfr new_Jinkela_buffer_8348 (
        .din(new_Jinkela_wire_10289),
        .dout(new_Jinkela_wire_10290)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_2177),
        .dout(new_Jinkela_wire_2178)
    );

    bfr new_Jinkela_buffer_8317 (
        .din(new_Jinkela_wire_10244),
        .dout(new_Jinkela_wire_10245)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(new_Jinkela_wire_2095),
        .dout(new_Jinkela_wire_2096)
    );

    spl2 new_Jinkela_splitter_826 (
        .a(_0328_),
        .b(new_Jinkela_wire_10558),
        .c(new_Jinkela_wire_10559)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_Jinkela_wire_2270),
        .dout(new_Jinkela_wire_2271)
    );

    bfr new_Jinkela_buffer_8318 (
        .din(new_Jinkela_wire_10245),
        .dout(new_Jinkela_wire_10246)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_2096),
        .dout(new_Jinkela_wire_2097)
    );

    bfr new_Jinkela_buffer_8349 (
        .din(new_Jinkela_wire_10290),
        .dout(new_Jinkela_wire_10291)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_2178),
        .dout(new_Jinkela_wire_2179)
    );

    bfr new_Jinkela_buffer_8319 (
        .din(new_Jinkela_wire_10246),
        .dout(new_Jinkela_wire_10247)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_2097),
        .dout(new_Jinkela_wire_2098)
    );

    bfr new_Jinkela_buffer_8454 (
        .din(new_Jinkela_wire_10403),
        .dout(new_Jinkela_wire_10404)
    );

    spl2 new_Jinkela_splitter_283 (
        .a(new_Jinkela_wire_2321),
        .b(new_Jinkela_wire_2322),
        .c(new_Jinkela_wire_2323)
    );

    bfr new_Jinkela_buffer_8320 (
        .din(new_Jinkela_wire_10247),
        .dout(new_Jinkela_wire_10248)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(new_Jinkela_wire_2098),
        .dout(new_Jinkela_wire_2099)
    );

    bfr new_Jinkela_buffer_8350 (
        .din(new_Jinkela_wire_10291),
        .dout(new_Jinkela_wire_10292)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_2179),
        .dout(new_Jinkela_wire_2180)
    );

    bfr new_Jinkela_buffer_8321 (
        .din(new_Jinkela_wire_10248),
        .dout(new_Jinkela_wire_10249)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_2099),
        .dout(new_Jinkela_wire_2100)
    );

    bfr new_Jinkela_buffer_8493 (
        .din(new_Jinkela_wire_10442),
        .dout(new_Jinkela_wire_10443)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_2271),
        .dout(new_Jinkela_wire_2272)
    );

    bfr new_Jinkela_buffer_8322 (
        .din(new_Jinkela_wire_10249),
        .dout(new_Jinkela_wire_10250)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_2100),
        .dout(new_Jinkela_wire_2101)
    );

    bfr new_Jinkela_buffer_8351 (
        .din(new_Jinkela_wire_10292),
        .dout(new_Jinkela_wire_10293)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_2180),
        .dout(new_Jinkela_wire_2181)
    );

    bfr new_Jinkela_buffer_8323 (
        .din(new_Jinkela_wire_10250),
        .dout(new_Jinkela_wire_10251)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_2101),
        .dout(new_Jinkela_wire_2102)
    );

    bfr new_Jinkela_buffer_8455 (
        .din(new_Jinkela_wire_10404),
        .dout(new_Jinkela_wire_10405)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(new_Jinkela_wire_2327),
        .dout(new_Jinkela_wire_2328)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(_0848_),
        .dout(new_Jinkela_wire_2342)
    );

    bfr new_Jinkela_buffer_8324 (
        .din(new_Jinkela_wire_10251),
        .dout(new_Jinkela_wire_10252)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_2102),
        .dout(new_Jinkela_wire_2103)
    );

    bfr new_Jinkela_buffer_8352 (
        .din(new_Jinkela_wire_10293),
        .dout(new_Jinkela_wire_10294)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_2181),
        .dout(new_Jinkela_wire_2182)
    );

    bfr new_Jinkela_buffer_8325 (
        .din(new_Jinkela_wire_10252),
        .dout(new_Jinkela_wire_10253)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(new_Jinkela_wire_2103),
        .dout(new_Jinkela_wire_2104)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_2272),
        .dout(new_Jinkela_wire_2273)
    );

    spl2 new_Jinkela_splitter_827 (
        .a(_0959_),
        .b(new_Jinkela_wire_10560),
        .c(new_Jinkela_wire_10561)
    );

    bfr new_Jinkela_buffer_8326 (
        .din(new_Jinkela_wire_10253),
        .dout(new_Jinkela_wire_10254)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(new_Jinkela_wire_2104),
        .dout(new_Jinkela_wire_2105)
    );

    bfr new_Jinkela_buffer_8353 (
        .din(new_Jinkela_wire_10294),
        .dout(new_Jinkela_wire_10295)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_2182),
        .dout(new_Jinkela_wire_2183)
    );

    spl2 new_Jinkela_splitter_813 (
        .a(new_Jinkela_wire_10254),
        .b(new_Jinkela_wire_10255),
        .c(new_Jinkela_wire_10256)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_2105),
        .dout(new_Jinkela_wire_2106)
    );

    bfr new_Jinkela_buffer_8354 (
        .din(new_Jinkela_wire_10295),
        .dout(new_Jinkela_wire_10296)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(_1476_),
        .dout(new_Jinkela_wire_2332)
    );

    bfr new_Jinkela_buffer_8456 (
        .din(new_Jinkela_wire_10405),
        .dout(new_Jinkela_wire_10406)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_2106),
        .dout(new_Jinkela_wire_2107)
    );

    bfr new_Jinkela_buffer_8494 (
        .din(new_Jinkela_wire_10443),
        .dout(new_Jinkela_wire_10444)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_2183),
        .dout(new_Jinkela_wire_2184)
    );

    bfr new_Jinkela_buffer_8355 (
        .din(new_Jinkela_wire_10296),
        .dout(new_Jinkela_wire_10297)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(new_Jinkela_wire_2107),
        .dout(new_Jinkela_wire_2108)
    );

    bfr new_Jinkela_buffer_8457 (
        .din(new_Jinkela_wire_10406),
        .dout(new_Jinkela_wire_10407)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_2273),
        .dout(new_Jinkela_wire_2274)
    );

    bfr new_Jinkela_buffer_8356 (
        .din(new_Jinkela_wire_10297),
        .dout(new_Jinkela_wire_10298)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_2108),
        .dout(new_Jinkela_wire_2109)
    );

    bfr new_Jinkela_buffer_8501 (
        .din(new_Jinkela_wire_10452),
        .dout(new_Jinkela_wire_10453)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_Jinkela_wire_2184),
        .dout(new_Jinkela_wire_2185)
    );

    bfr new_Jinkela_buffer_8357 (
        .din(new_Jinkela_wire_10298),
        .dout(new_Jinkela_wire_10299)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_2109),
        .dout(new_Jinkela_wire_2110)
    );

    bfr new_Jinkela_buffer_8458 (
        .din(new_Jinkela_wire_10407),
        .dout(new_Jinkela_wire_10408)
    );

    spl2 new_Jinkela_splitter_287 (
        .a(_0317_),
        .b(new_Jinkela_wire_2343),
        .c(new_Jinkela_wire_2344)
    );

    bfr new_Jinkela_buffer_8358 (
        .din(new_Jinkela_wire_10299),
        .dout(new_Jinkela_wire_10300)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(new_Jinkela_wire_2110),
        .dout(new_Jinkela_wire_2111)
    );

    bfr new_Jinkela_buffer_8495 (
        .din(new_Jinkela_wire_10444),
        .dout(new_Jinkela_wire_10445)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_2185),
        .dout(new_Jinkela_wire_2186)
    );

    bfr new_Jinkela_buffer_8359 (
        .din(new_Jinkela_wire_10300),
        .dout(new_Jinkela_wire_10301)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(new_Jinkela_wire_2111),
        .dout(new_Jinkela_wire_2112)
    );

    bfr new_Jinkela_buffer_8459 (
        .din(new_Jinkela_wire_10408),
        .dout(new_Jinkela_wire_10409)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_2274),
        .dout(new_Jinkela_wire_2275)
    );

    bfr new_Jinkela_buffer_4947 (
        .din(new_Jinkela_wire_6392),
        .dout(new_Jinkela_wire_6393)
    );

    bfr new_Jinkela_buffer_15349 (
        .din(new_Jinkela_wire_18299),
        .dout(new_Jinkela_wire_18300)
    );

    bfr new_Jinkela_buffer_4861 (
        .din(new_Jinkela_wire_6292),
        .dout(new_Jinkela_wire_6293)
    );

    bfr new_Jinkela_buffer_15234 (
        .din(new_Jinkela_wire_18168),
        .dout(new_Jinkela_wire_18169)
    );

    bfr new_Jinkela_buffer_15307 (
        .din(new_Jinkela_wire_18247),
        .dout(new_Jinkela_wire_18248)
    );

    bfr new_Jinkela_buffer_4862 (
        .din(new_Jinkela_wire_6293),
        .dout(new_Jinkela_wire_6294)
    );

    bfr new_Jinkela_buffer_15235 (
        .din(new_Jinkela_wire_18169),
        .dout(new_Jinkela_wire_18170)
    );

    bfr new_Jinkela_buffer_4948 (
        .din(new_Jinkela_wire_6393),
        .dout(new_Jinkela_wire_6394)
    );

    bfr new_Jinkela_buffer_15356 (
        .din(new_Jinkela_wire_18310),
        .dout(new_Jinkela_wire_18311)
    );

    bfr new_Jinkela_buffer_4863 (
        .din(new_Jinkela_wire_6294),
        .dout(new_Jinkela_wire_6295)
    );

    bfr new_Jinkela_buffer_15236 (
        .din(new_Jinkela_wire_18170),
        .dout(new_Jinkela_wire_18171)
    );

    bfr new_Jinkela_buffer_4964 (
        .din(new_Jinkela_wire_6423),
        .dout(new_Jinkela_wire_6424)
    );

    bfr new_Jinkela_buffer_15308 (
        .din(new_Jinkela_wire_18248),
        .dout(new_Jinkela_wire_18249)
    );

    bfr new_Jinkela_buffer_4864 (
        .din(new_Jinkela_wire_6295),
        .dout(new_Jinkela_wire_6296)
    );

    bfr new_Jinkela_buffer_15237 (
        .din(new_Jinkela_wire_18171),
        .dout(new_Jinkela_wire_18172)
    );

    bfr new_Jinkela_buffer_4949 (
        .din(new_Jinkela_wire_6394),
        .dout(new_Jinkela_wire_6395)
    );

    bfr new_Jinkela_buffer_15350 (
        .din(new_Jinkela_wire_18300),
        .dout(new_Jinkela_wire_18301)
    );

    bfr new_Jinkela_buffer_4865 (
        .din(new_Jinkela_wire_6296),
        .dout(new_Jinkela_wire_6297)
    );

    bfr new_Jinkela_buffer_15238 (
        .din(new_Jinkela_wire_18172),
        .dout(new_Jinkela_wire_18173)
    );

    bfr new_Jinkela_buffer_15309 (
        .din(new_Jinkela_wire_18249),
        .dout(new_Jinkela_wire_18250)
    );

    bfr new_Jinkela_buffer_4866 (
        .din(new_Jinkela_wire_6297),
        .dout(new_Jinkela_wire_6298)
    );

    bfr new_Jinkela_buffer_15239 (
        .din(new_Jinkela_wire_18173),
        .dout(new_Jinkela_wire_18174)
    );

    spl2 new_Jinkela_splitter_582 (
        .a(_1220_),
        .b(new_Jinkela_wire_6516),
        .c(new_Jinkela_wire_6517)
    );

    bfr new_Jinkela_buffer_4950 (
        .din(new_Jinkela_wire_6395),
        .dout(new_Jinkela_wire_6396)
    );

    bfr new_Jinkela_buffer_4867 (
        .din(new_Jinkela_wire_6298),
        .dout(new_Jinkela_wire_6299)
    );

    spl2 new_Jinkela_splitter_1327 (
        .a(_1780_),
        .b(new_Jinkela_wire_18375),
        .c(new_Jinkela_wire_18376)
    );

    bfr new_Jinkela_buffer_15240 (
        .din(new_Jinkela_wire_18174),
        .dout(new_Jinkela_wire_18175)
    );

    bfr new_Jinkela_buffer_4965 (
        .din(new_Jinkela_wire_6424),
        .dout(new_Jinkela_wire_6425)
    );

    bfr new_Jinkela_buffer_15310 (
        .din(new_Jinkela_wire_18250),
        .dout(new_Jinkela_wire_18251)
    );

    bfr new_Jinkela_buffer_4868 (
        .din(new_Jinkela_wire_6299),
        .dout(new_Jinkela_wire_6300)
    );

    bfr new_Jinkela_buffer_15241 (
        .din(new_Jinkela_wire_18175),
        .dout(new_Jinkela_wire_18176)
    );

    bfr new_Jinkela_buffer_4951 (
        .din(new_Jinkela_wire_6396),
        .dout(new_Jinkela_wire_6397)
    );

    bfr new_Jinkela_buffer_15351 (
        .din(new_Jinkela_wire_18301),
        .dout(new_Jinkela_wire_18302)
    );

    bfr new_Jinkela_buffer_4869 (
        .din(new_Jinkela_wire_6300),
        .dout(new_Jinkela_wire_6301)
    );

    bfr new_Jinkela_buffer_15242 (
        .din(new_Jinkela_wire_18176),
        .dout(new_Jinkela_wire_18177)
    );

    bfr new_Jinkela_buffer_15311 (
        .din(new_Jinkela_wire_18251),
        .dout(new_Jinkela_wire_18252)
    );

    bfr new_Jinkela_buffer_4870 (
        .din(new_Jinkela_wire_6301),
        .dout(new_Jinkela_wire_6302)
    );

    bfr new_Jinkela_buffer_15243 (
        .din(new_Jinkela_wire_18177),
        .dout(new_Jinkela_wire_18178)
    );

    bfr new_Jinkela_buffer_5050 (
        .din(_1500_),
        .dout(new_Jinkela_wire_6518)
    );

    bfr new_Jinkela_buffer_4952 (
        .din(new_Jinkela_wire_6397),
        .dout(new_Jinkela_wire_6398)
    );

    bfr new_Jinkela_buffer_4871 (
        .din(new_Jinkela_wire_6302),
        .dout(new_Jinkela_wire_6303)
    );

    spl2 new_Jinkela_splitter_1328 (
        .a(_0063_),
        .b(new_Jinkela_wire_18377),
        .c(new_Jinkela_wire_18378)
    );

    bfr new_Jinkela_buffer_15244 (
        .din(new_Jinkela_wire_18178),
        .dout(new_Jinkela_wire_18179)
    );

    bfr new_Jinkela_buffer_4966 (
        .din(new_Jinkela_wire_6425),
        .dout(new_Jinkela_wire_6426)
    );

    bfr new_Jinkela_buffer_15312 (
        .din(new_Jinkela_wire_18252),
        .dout(new_Jinkela_wire_18253)
    );

    bfr new_Jinkela_buffer_4872 (
        .din(new_Jinkela_wire_6303),
        .dout(new_Jinkela_wire_6304)
    );

    bfr new_Jinkela_buffer_15245 (
        .din(new_Jinkela_wire_18179),
        .dout(new_Jinkela_wire_18180)
    );

    bfr new_Jinkela_buffer_4953 (
        .din(new_Jinkela_wire_6398),
        .dout(new_Jinkela_wire_6399)
    );

    bfr new_Jinkela_buffer_15352 (
        .din(new_Jinkela_wire_18302),
        .dout(new_Jinkela_wire_18303)
    );

    bfr new_Jinkela_buffer_4873 (
        .din(new_Jinkela_wire_6304),
        .dout(new_Jinkela_wire_6305)
    );

    bfr new_Jinkela_buffer_15246 (
        .din(new_Jinkela_wire_18180),
        .dout(new_Jinkela_wire_18181)
    );

    spl2 new_Jinkela_splitter_584 (
        .a(_0890_),
        .b(new_Jinkela_wire_6521),
        .c(new_Jinkela_wire_6522)
    );

    bfr new_Jinkela_buffer_15313 (
        .din(new_Jinkela_wire_18253),
        .dout(new_Jinkela_wire_18254)
    );

    bfr new_Jinkela_buffer_4874 (
        .din(new_Jinkela_wire_6305),
        .dout(new_Jinkela_wire_6306)
    );

    bfr new_Jinkela_buffer_15247 (
        .din(new_Jinkela_wire_18181),
        .dout(new_Jinkela_wire_18182)
    );

    spl2 new_Jinkela_splitter_583 (
        .a(_1443_),
        .b(new_Jinkela_wire_6519),
        .c(new_Jinkela_wire_6520)
    );

    bfr new_Jinkela_buffer_4954 (
        .din(new_Jinkela_wire_6399),
        .dout(new_Jinkela_wire_6400)
    );

    bfr new_Jinkela_buffer_15357 (
        .din(new_Jinkela_wire_18311),
        .dout(new_Jinkela_wire_18312)
    );

    bfr new_Jinkela_buffer_4875 (
        .din(new_Jinkela_wire_6306),
        .dout(new_Jinkela_wire_6307)
    );

    bfr new_Jinkela_buffer_15248 (
        .din(new_Jinkela_wire_18182),
        .dout(new_Jinkela_wire_18183)
    );

    bfr new_Jinkela_buffer_4967 (
        .din(new_Jinkela_wire_6426),
        .dout(new_Jinkela_wire_6427)
    );

    bfr new_Jinkela_buffer_15314 (
        .din(new_Jinkela_wire_18254),
        .dout(new_Jinkela_wire_18255)
    );

    bfr new_Jinkela_buffer_4876 (
        .din(new_Jinkela_wire_6307),
        .dout(new_Jinkela_wire_6308)
    );

    bfr new_Jinkela_buffer_15249 (
        .din(new_Jinkela_wire_18183),
        .dout(new_Jinkela_wire_18184)
    );

    bfr new_Jinkela_buffer_4955 (
        .din(new_Jinkela_wire_6400),
        .dout(new_Jinkela_wire_6401)
    );

    bfr new_Jinkela_buffer_15353 (
        .din(new_Jinkela_wire_18303),
        .dout(new_Jinkela_wire_18304)
    );

    bfr new_Jinkela_buffer_4877 (
        .din(new_Jinkela_wire_6308),
        .dout(new_Jinkela_wire_6309)
    );

    bfr new_Jinkela_buffer_15250 (
        .din(new_Jinkela_wire_18184),
        .dout(new_Jinkela_wire_18185)
    );

    bfr new_Jinkela_buffer_5051 (
        .din(_1268_),
        .dout(new_Jinkela_wire_6523)
    );

    bfr new_Jinkela_buffer_15315 (
        .din(new_Jinkela_wire_18255),
        .dout(new_Jinkela_wire_18256)
    );

    bfr new_Jinkela_buffer_4878 (
        .din(new_Jinkela_wire_6309),
        .dout(new_Jinkela_wire_6310)
    );

    bfr new_Jinkela_buffer_15251 (
        .din(new_Jinkela_wire_18185),
        .dout(new_Jinkela_wire_18186)
    );

    bfr new_Jinkela_buffer_4956 (
        .din(new_Jinkela_wire_6401),
        .dout(new_Jinkela_wire_6402)
    );

    bfr new_Jinkela_buffer_15361 (
        .din(new_Jinkela_wire_18315),
        .dout(new_Jinkela_wire_18316)
    );

    bfr new_Jinkela_buffer_4879 (
        .din(new_Jinkela_wire_6310),
        .dout(new_Jinkela_wire_6311)
    );

    bfr new_Jinkela_buffer_15252 (
        .din(new_Jinkela_wire_18186),
        .dout(new_Jinkela_wire_18187)
    );

    bfr new_Jinkela_buffer_4968 (
        .din(new_Jinkela_wire_6427),
        .dout(new_Jinkela_wire_6428)
    );

    bfr new_Jinkela_buffer_15316 (
        .din(new_Jinkela_wire_18256),
        .dout(new_Jinkela_wire_18257)
    );

    bfr new_Jinkela_buffer_4880 (
        .din(new_Jinkela_wire_6311),
        .dout(new_Jinkela_wire_6312)
    );

    bfr new_Jinkela_buffer_15253 (
        .din(new_Jinkela_wire_18187),
        .dout(new_Jinkela_wire_18188)
    );

    spl2 new_Jinkela_splitter_572 (
        .a(new_Jinkela_wire_6402),
        .b(new_Jinkela_wire_6403),
        .c(new_Jinkela_wire_6404)
    );

    bfr new_Jinkela_buffer_15354 (
        .din(new_Jinkela_wire_18304),
        .dout(new_Jinkela_wire_18305)
    );

    bfr new_Jinkela_buffer_4881 (
        .din(new_Jinkela_wire_6312),
        .dout(new_Jinkela_wire_6313)
    );

    bfr new_Jinkela_buffer_15254 (
        .din(new_Jinkela_wire_18188),
        .dout(new_Jinkela_wire_18189)
    );

    bfr new_Jinkela_buffer_14381 (
        .din(new_Jinkela_wire_17195),
        .dout(new_Jinkela_wire_17196)
    );

    spl2 new_Jinkela_splitter_1266 (
        .a(_1313_),
        .b(new_Jinkela_wire_17534),
        .c(new_Jinkela_wire_17535)
    );

    bfr new_Jinkela_buffer_14521 (
        .din(new_Jinkela_wire_17337),
        .dout(new_Jinkela_wire_17338)
    );

    bfr new_Jinkela_buffer_14382 (
        .din(new_Jinkela_wire_17196),
        .dout(new_Jinkela_wire_17197)
    );

    bfr new_Jinkela_buffer_14544 (
        .din(new_Jinkela_wire_17368),
        .dout(new_Jinkela_wire_17369)
    );

    bfr new_Jinkela_buffer_14383 (
        .din(new_Jinkela_wire_17197),
        .dout(new_Jinkela_wire_17198)
    );

    bfr new_Jinkela_buffer_14522 (
        .din(new_Jinkela_wire_17338),
        .dout(new_Jinkela_wire_17339)
    );

    bfr new_Jinkela_buffer_14384 (
        .din(new_Jinkela_wire_17198),
        .dout(new_Jinkela_wire_17199)
    );

    bfr new_Jinkela_buffer_14549 (
        .din(new_Jinkela_wire_17375),
        .dout(new_Jinkela_wire_17376)
    );

    bfr new_Jinkela_buffer_14385 (
        .din(new_Jinkela_wire_17199),
        .dout(new_Jinkela_wire_17200)
    );

    bfr new_Jinkela_buffer_14523 (
        .din(new_Jinkela_wire_17339),
        .dout(new_Jinkela_wire_17340)
    );

    bfr new_Jinkela_buffer_14386 (
        .din(new_Jinkela_wire_17200),
        .dout(new_Jinkela_wire_17201)
    );

    bfr new_Jinkela_buffer_14545 (
        .din(new_Jinkela_wire_17369),
        .dout(new_Jinkela_wire_17370)
    );

    bfr new_Jinkela_buffer_14387 (
        .din(new_Jinkela_wire_17201),
        .dout(new_Jinkela_wire_17202)
    );

    bfr new_Jinkela_buffer_14524 (
        .din(new_Jinkela_wire_17340),
        .dout(new_Jinkela_wire_17341)
    );

    bfr new_Jinkela_buffer_14388 (
        .din(new_Jinkela_wire_17202),
        .dout(new_Jinkela_wire_17203)
    );

    bfr new_Jinkela_buffer_14389 (
        .din(new_Jinkela_wire_17203),
        .dout(new_Jinkela_wire_17204)
    );

    spl2 new_Jinkela_splitter_1265 (
        .a(_0935_),
        .b(new_Jinkela_wire_17532),
        .c(new_Jinkela_wire_17533)
    );

    bfr new_Jinkela_buffer_14525 (
        .din(new_Jinkela_wire_17341),
        .dout(new_Jinkela_wire_17342)
    );

    bfr new_Jinkela_buffer_14390 (
        .din(new_Jinkela_wire_17204),
        .dout(new_Jinkela_wire_17205)
    );

    spl2 new_Jinkela_splitter_1261 (
        .a(new_Jinkela_wire_17370),
        .b(new_Jinkela_wire_17371),
        .c(new_Jinkela_wire_17372)
    );

    bfr new_Jinkela_buffer_14391 (
        .din(new_Jinkela_wire_17205),
        .dout(new_Jinkela_wire_17206)
    );

    bfr new_Jinkela_buffer_14526 (
        .din(new_Jinkela_wire_17342),
        .dout(new_Jinkela_wire_17343)
    );

    bfr new_Jinkela_buffer_14392 (
        .din(new_Jinkela_wire_17206),
        .dout(new_Jinkela_wire_17207)
    );

    bfr new_Jinkela_buffer_14596 (
        .din(new_Jinkela_wire_17426),
        .dout(new_Jinkela_wire_17427)
    );

    bfr new_Jinkela_buffer_14393 (
        .din(new_Jinkela_wire_17207),
        .dout(new_Jinkela_wire_17208)
    );

    bfr new_Jinkela_buffer_14527 (
        .din(new_Jinkela_wire_17343),
        .dout(new_Jinkela_wire_17344)
    );

    bfr new_Jinkela_buffer_14394 (
        .din(new_Jinkela_wire_17208),
        .dout(new_Jinkela_wire_17209)
    );

    bfr new_Jinkela_buffer_14550 (
        .din(new_Jinkela_wire_17376),
        .dout(new_Jinkela_wire_17377)
    );

    bfr new_Jinkela_buffer_14395 (
        .din(new_Jinkela_wire_17209),
        .dout(new_Jinkela_wire_17210)
    );

    bfr new_Jinkela_buffer_14528 (
        .din(new_Jinkela_wire_17344),
        .dout(new_Jinkela_wire_17345)
    );

    bfr new_Jinkela_buffer_14396 (
        .din(new_Jinkela_wire_17210),
        .dout(new_Jinkela_wire_17211)
    );

    bfr new_Jinkela_buffer_14551 (
        .din(new_Jinkela_wire_17377),
        .dout(new_Jinkela_wire_17378)
    );

    bfr new_Jinkela_buffer_14397 (
        .din(new_Jinkela_wire_17211),
        .dout(new_Jinkela_wire_17212)
    );

    bfr new_Jinkela_buffer_14529 (
        .din(new_Jinkela_wire_17345),
        .dout(new_Jinkela_wire_17346)
    );

    bfr new_Jinkela_buffer_14398 (
        .din(new_Jinkela_wire_17212),
        .dout(new_Jinkela_wire_17213)
    );

    spl2 new_Jinkela_splitter_1267 (
        .a(_0973_),
        .b(new_Jinkela_wire_17536),
        .c(new_Jinkela_wire_17537)
    );

    bfr new_Jinkela_buffer_14399 (
        .din(new_Jinkela_wire_17213),
        .dout(new_Jinkela_wire_17214)
    );

    bfr new_Jinkela_buffer_14530 (
        .din(new_Jinkela_wire_17346),
        .dout(new_Jinkela_wire_17347)
    );

    bfr new_Jinkela_buffer_14400 (
        .din(new_Jinkela_wire_17214),
        .dout(new_Jinkela_wire_17215)
    );

    bfr new_Jinkela_buffer_14552 (
        .din(new_Jinkela_wire_17378),
        .dout(new_Jinkela_wire_17379)
    );

    bfr new_Jinkela_buffer_14401 (
        .din(new_Jinkela_wire_17215),
        .dout(new_Jinkela_wire_17216)
    );

    bfr new_Jinkela_buffer_7446 (
        .din(new_Jinkela_wire_9261),
        .dout(new_Jinkela_wire_9262)
    );

    bfr new_Jinkela_buffer_7551 (
        .din(new_Jinkela_wire_9374),
        .dout(new_Jinkela_wire_9375)
    );

    bfr new_Jinkela_buffer_7447 (
        .din(new_Jinkela_wire_9262),
        .dout(new_Jinkela_wire_9263)
    );

    bfr new_Jinkela_buffer_7519 (
        .din(new_Jinkela_wire_9336),
        .dout(new_Jinkela_wire_9337)
    );

    bfr new_Jinkela_buffer_7448 (
        .din(new_Jinkela_wire_9263),
        .dout(new_Jinkela_wire_9264)
    );

    spl2 new_Jinkela_splitter_767 (
        .a(_1447_),
        .b(new_Jinkela_wire_9544),
        .c(new_Jinkela_wire_9545)
    );

    bfr new_Jinkela_buffer_7449 (
        .din(new_Jinkela_wire_9264),
        .dout(new_Jinkela_wire_9265)
    );

    bfr new_Jinkela_buffer_7520 (
        .din(new_Jinkela_wire_9337),
        .dout(new_Jinkela_wire_9338)
    );

    bfr new_Jinkela_buffer_7450 (
        .din(new_Jinkela_wire_9265),
        .dout(new_Jinkela_wire_9266)
    );

    bfr new_Jinkela_buffer_7552 (
        .din(new_Jinkela_wire_9375),
        .dout(new_Jinkela_wire_9376)
    );

    bfr new_Jinkela_buffer_7451 (
        .din(new_Jinkela_wire_9266),
        .dout(new_Jinkela_wire_9267)
    );

    bfr new_Jinkela_buffer_7521 (
        .din(new_Jinkela_wire_9338),
        .dout(new_Jinkela_wire_9339)
    );

    bfr new_Jinkela_buffer_7452 (
        .din(new_Jinkela_wire_9267),
        .dout(new_Jinkela_wire_9268)
    );

    bfr new_Jinkela_buffer_7625 (
        .din(new_Jinkela_wire_9452),
        .dout(new_Jinkela_wire_9453)
    );

    bfr new_Jinkela_buffer_7453 (
        .din(new_Jinkela_wire_9268),
        .dout(new_Jinkela_wire_9269)
    );

    bfr new_Jinkela_buffer_7522 (
        .din(new_Jinkela_wire_9339),
        .dout(new_Jinkela_wire_9340)
    );

    bfr new_Jinkela_buffer_7454 (
        .din(new_Jinkela_wire_9269),
        .dout(new_Jinkela_wire_9270)
    );

    bfr new_Jinkela_buffer_7553 (
        .din(new_Jinkela_wire_9376),
        .dout(new_Jinkela_wire_9377)
    );

    bfr new_Jinkela_buffer_7455 (
        .din(new_Jinkela_wire_9270),
        .dout(new_Jinkela_wire_9271)
    );

    bfr new_Jinkela_buffer_7523 (
        .din(new_Jinkela_wire_9340),
        .dout(new_Jinkela_wire_9341)
    );

    bfr new_Jinkela_buffer_7456 (
        .din(new_Jinkela_wire_9271),
        .dout(new_Jinkela_wire_9272)
    );

    bfr new_Jinkela_buffer_7685 (
        .din(new_Jinkela_wire_9512),
        .dout(new_Jinkela_wire_9513)
    );

    bfr new_Jinkela_buffer_7457 (
        .din(new_Jinkela_wire_9272),
        .dout(new_Jinkela_wire_9273)
    );

    bfr new_Jinkela_buffer_7524 (
        .din(new_Jinkela_wire_9341),
        .dout(new_Jinkela_wire_9342)
    );

    bfr new_Jinkela_buffer_7458 (
        .din(new_Jinkela_wire_9273),
        .dout(new_Jinkela_wire_9274)
    );

    bfr new_Jinkela_buffer_7554 (
        .din(new_Jinkela_wire_9377),
        .dout(new_Jinkela_wire_9378)
    );

    bfr new_Jinkela_buffer_7459 (
        .din(new_Jinkela_wire_9274),
        .dout(new_Jinkela_wire_9275)
    );

    bfr new_Jinkela_buffer_7525 (
        .din(new_Jinkela_wire_9342),
        .dout(new_Jinkela_wire_9343)
    );

    bfr new_Jinkela_buffer_7460 (
        .din(new_Jinkela_wire_9275),
        .dout(new_Jinkela_wire_9276)
    );

    bfr new_Jinkela_buffer_7626 (
        .din(new_Jinkela_wire_9453),
        .dout(new_Jinkela_wire_9454)
    );

    bfr new_Jinkela_buffer_7461 (
        .din(new_Jinkela_wire_9276),
        .dout(new_Jinkela_wire_9277)
    );

    bfr new_Jinkela_buffer_7526 (
        .din(new_Jinkela_wire_9343),
        .dout(new_Jinkela_wire_9344)
    );

    bfr new_Jinkela_buffer_7462 (
        .din(new_Jinkela_wire_9277),
        .dout(new_Jinkela_wire_9278)
    );

    bfr new_Jinkela_buffer_7555 (
        .din(new_Jinkela_wire_9378),
        .dout(new_Jinkela_wire_9379)
    );

    bfr new_Jinkela_buffer_7463 (
        .din(new_Jinkela_wire_9278),
        .dout(new_Jinkela_wire_9279)
    );

    spl2 new_Jinkela_splitter_758 (
        .a(new_Jinkela_wire_9344),
        .b(new_Jinkela_wire_9345),
        .c(new_Jinkela_wire_9346)
    );

    bfr new_Jinkela_buffer_7464 (
        .din(new_Jinkela_wire_9279),
        .dout(new_Jinkela_wire_9280)
    );

    bfr new_Jinkela_buffer_7556 (
        .din(new_Jinkela_wire_9379),
        .dout(new_Jinkela_wire_9380)
    );

    bfr new_Jinkela_buffer_7465 (
        .din(new_Jinkela_wire_9280),
        .dout(new_Jinkela_wire_9281)
    );

    bfr new_Jinkela_buffer_7466 (
        .din(new_Jinkela_wire_9281),
        .dout(new_Jinkela_wire_9282)
    );

    bfr new_Jinkela_buffer_7627 (
        .din(new_Jinkela_wire_9454),
        .dout(new_Jinkela_wire_9455)
    );

    bfr new_Jinkela_buffer_4080 (
        .din(new_Jinkela_wire_5355),
        .dout(new_Jinkela_wire_5356)
    );

    bfr new_Jinkela_buffer_17815 (
        .din(new_Jinkela_wire_21247),
        .dout(new_Jinkela_wire_21248)
    );

    bfr new_Jinkela_buffer_4000 (
        .din(new_Jinkela_wire_5267),
        .dout(new_Jinkela_wire_5268)
    );

    bfr new_Jinkela_buffer_17816 (
        .din(new_Jinkela_wire_21248),
        .dout(new_Jinkela_wire_21249)
    );

    spl2 new_Jinkela_splitter_503 (
        .a(_0517_),
        .b(new_Jinkela_wire_5465),
        .c(new_Jinkela_wire_5466)
    );

    bfr new_Jinkela_buffer_4001 (
        .din(new_Jinkela_wire_5268),
        .dout(new_Jinkela_wire_5269)
    );

    bfr new_Jinkela_buffer_4081 (
        .din(new_Jinkela_wire_5356),
        .dout(new_Jinkela_wire_5357)
    );

    bfr new_Jinkela_buffer_17817 (
        .din(new_Jinkela_wire_21249),
        .dout(new_Jinkela_wire_21250)
    );

    bfr new_Jinkela_buffer_4002 (
        .din(new_Jinkela_wire_5269),
        .dout(new_Jinkela_wire_5270)
    );

    bfr new_Jinkela_buffer_17818 (
        .din(new_Jinkela_wire_21250),
        .dout(new_Jinkela_wire_21251)
    );

    bfr new_Jinkela_buffer_4003 (
        .din(new_Jinkela_wire_5270),
        .dout(new_Jinkela_wire_5271)
    );

    bfr new_Jinkela_buffer_4082 (
        .din(new_Jinkela_wire_5357),
        .dout(new_Jinkela_wire_5358)
    );

    bfr new_Jinkela_buffer_17819 (
        .din(new_Jinkela_wire_21251),
        .dout(new_Jinkela_wire_21252)
    );

    bfr new_Jinkela_buffer_4004 (
        .din(new_Jinkela_wire_5271),
        .dout(new_Jinkela_wire_5272)
    );

    bfr new_Jinkela_buffer_4154 (
        .din(new_Jinkela_wire_5459),
        .dout(new_Jinkela_wire_5460)
    );

    bfr new_Jinkela_buffer_17820 (
        .din(new_Jinkela_wire_21252),
        .dout(new_Jinkela_wire_21253)
    );

    bfr new_Jinkela_buffer_4005 (
        .din(new_Jinkela_wire_5272),
        .dout(new_Jinkela_wire_5273)
    );

    bfr new_Jinkela_buffer_4083 (
        .din(new_Jinkela_wire_5358),
        .dout(new_Jinkela_wire_5359)
    );

    bfr new_Jinkela_buffer_17821 (
        .din(new_Jinkela_wire_21253),
        .dout(new_Jinkela_wire_21254)
    );

    bfr new_Jinkela_buffer_4006 (
        .din(new_Jinkela_wire_5273),
        .dout(new_Jinkela_wire_5274)
    );

    bfr new_Jinkela_buffer_17822 (
        .din(new_Jinkela_wire_21254),
        .dout(new_Jinkela_wire_21255)
    );

    spl2 new_Jinkela_splitter_504 (
        .a(_0672_),
        .b(new_Jinkela_wire_5467),
        .c(new_Jinkela_wire_5468)
    );

    bfr new_Jinkela_buffer_4007 (
        .din(new_Jinkela_wire_5274),
        .dout(new_Jinkela_wire_5275)
    );

    bfr new_Jinkela_buffer_4084 (
        .din(new_Jinkela_wire_5359),
        .dout(new_Jinkela_wire_5360)
    );

    bfr new_Jinkela_buffer_17823 (
        .din(new_Jinkela_wire_21255),
        .dout(new_Jinkela_wire_21256)
    );

    bfr new_Jinkela_buffer_4008 (
        .din(new_Jinkela_wire_5275),
        .dout(new_Jinkela_wire_5276)
    );

    bfr new_Jinkela_buffer_4155 (
        .din(new_Jinkela_wire_5460),
        .dout(new_Jinkela_wire_5461)
    );

    bfr new_Jinkela_buffer_17824 (
        .din(new_Jinkela_wire_21256),
        .dout(new_Jinkela_wire_21257)
    );

    bfr new_Jinkela_buffer_4009 (
        .din(new_Jinkela_wire_5276),
        .dout(new_Jinkela_wire_5277)
    );

    bfr new_Jinkela_buffer_4085 (
        .din(new_Jinkela_wire_5360),
        .dout(new_Jinkela_wire_5361)
    );

    bfr new_Jinkela_buffer_17825 (
        .din(new_Jinkela_wire_21257),
        .dout(new_Jinkela_wire_21258)
    );

    bfr new_Jinkela_buffer_4010 (
        .din(new_Jinkela_wire_5277),
        .dout(new_Jinkela_wire_5278)
    );

    bfr new_Jinkela_buffer_4158 (
        .din(new_Jinkela_wire_5469),
        .dout(new_Jinkela_wire_5470)
    );

    bfr new_Jinkela_buffer_17826 (
        .din(new_Jinkela_wire_21258),
        .dout(new_Jinkela_wire_21259)
    );

    bfr new_Jinkela_buffer_4157 (
        .din(new_net_3942),
        .dout(new_Jinkela_wire_5469)
    );

    bfr new_Jinkela_buffer_4011 (
        .din(new_Jinkela_wire_5278),
        .dout(new_Jinkela_wire_5279)
    );

    bfr new_Jinkela_buffer_4086 (
        .din(new_Jinkela_wire_5361),
        .dout(new_Jinkela_wire_5362)
    );

    bfr new_Jinkela_buffer_17827 (
        .din(new_Jinkela_wire_21259),
        .dout(new_Jinkela_wire_21260)
    );

    spl2 new_Jinkela_splitter_483 (
        .a(new_Jinkela_wire_5279),
        .b(new_Jinkela_wire_5280),
        .c(new_Jinkela_wire_5281)
    );

    bfr new_Jinkela_buffer_4087 (
        .din(new_Jinkela_wire_5362),
        .dout(new_Jinkela_wire_5363)
    );

    bfr new_Jinkela_buffer_17828 (
        .din(new_Jinkela_wire_21260),
        .dout(new_Jinkela_wire_21261)
    );

    bfr new_Jinkela_buffer_4156 (
        .din(new_Jinkela_wire_5461),
        .dout(new_Jinkela_wire_5462)
    );

    bfr new_Jinkela_buffer_17829 (
        .din(new_Jinkela_wire_21261),
        .dout(new_Jinkela_wire_21262)
    );

    bfr new_Jinkela_buffer_4225 (
        .din(_0944_),
        .dout(new_Jinkela_wire_5537)
    );

    bfr new_Jinkela_buffer_4088 (
        .din(new_Jinkela_wire_5363),
        .dout(new_Jinkela_wire_5364)
    );

    bfr new_Jinkela_buffer_17830 (
        .din(new_Jinkela_wire_21262),
        .dout(new_Jinkela_wire_21263)
    );

    spl2 new_Jinkela_splitter_505 (
        .a(_0678_),
        .b(new_Jinkela_wire_5538),
        .c(new_Jinkela_wire_5539)
    );

    bfr new_Jinkela_buffer_4089 (
        .din(new_Jinkela_wire_5364),
        .dout(new_Jinkela_wire_5365)
    );

    spl2 new_Jinkela_splitter_506 (
        .a(_1661_),
        .b(new_Jinkela_wire_5540),
        .c(new_Jinkela_wire_5541)
    );

    bfr new_Jinkela_buffer_17831 (
        .din(new_Jinkela_wire_21263),
        .dout(new_Jinkela_wire_21264)
    );

    bfr new_Jinkela_buffer_4159 (
        .din(new_Jinkela_wire_5470),
        .dout(new_Jinkela_wire_5471)
    );

    bfr new_Jinkela_buffer_4090 (
        .din(new_Jinkela_wire_5365),
        .dout(new_Jinkela_wire_5366)
    );

    bfr new_Jinkela_buffer_17832 (
        .din(new_Jinkela_wire_21264),
        .dout(new_Jinkela_wire_21265)
    );

    spl2 new_Jinkela_splitter_507 (
        .a(_1610_),
        .b(new_Jinkela_wire_5542),
        .c(new_Jinkela_wire_5543)
    );

    bfr new_Jinkela_buffer_4091 (
        .din(new_Jinkela_wire_5366),
        .dout(new_Jinkela_wire_5367)
    );

    bfr new_Jinkela_buffer_17833 (
        .din(new_Jinkela_wire_21265),
        .dout(new_Jinkela_wire_21266)
    );

    bfr new_Jinkela_buffer_4160 (
        .din(new_Jinkela_wire_5471),
        .dout(new_Jinkela_wire_5472)
    );

    bfr new_Jinkela_buffer_4092 (
        .din(new_Jinkela_wire_5367),
        .dout(new_Jinkela_wire_5368)
    );

    bfr new_Jinkela_buffer_17834 (
        .din(new_Jinkela_wire_21266),
        .dout(new_Jinkela_wire_21267)
    );

    bfr new_Jinkela_buffer_4093 (
        .din(new_Jinkela_wire_5368),
        .dout(new_Jinkela_wire_5369)
    );

    bfr new_Jinkela_buffer_17835 (
        .din(new_Jinkela_wire_21267),
        .dout(new_Jinkela_wire_21268)
    );

    bfr new_Jinkela_buffer_4161 (
        .din(new_Jinkela_wire_5472),
        .dout(new_Jinkela_wire_5473)
    );

    bfr new_Jinkela_buffer_4094 (
        .din(new_Jinkela_wire_5369),
        .dout(new_Jinkela_wire_5370)
    );

    bfr new_Jinkela_buffer_11065 (
        .din(_0640_),
        .dout(new_Jinkela_wire_13341)
    );

    bfr new_Jinkela_buffer_10979 (
        .din(new_Jinkela_wire_13234),
        .dout(new_Jinkela_wire_13235)
    );

    bfr new_Jinkela_buffer_11058 (
        .din(new_Jinkela_wire_13327),
        .dout(new_Jinkela_wire_13328)
    );

    bfr new_Jinkela_buffer_10980 (
        .din(new_Jinkela_wire_13235),
        .dout(new_Jinkela_wire_13236)
    );

    bfr new_Jinkela_buffer_11066 (
        .din(new_Jinkela_wire_13343),
        .dout(new_Jinkela_wire_13344)
    );

    bfr new_Jinkela_buffer_10981 (
        .din(new_Jinkela_wire_13236),
        .dout(new_Jinkela_wire_13237)
    );

    bfr new_Jinkela_buffer_11059 (
        .din(new_Jinkela_wire_13328),
        .dout(new_Jinkela_wire_13329)
    );

    bfr new_Jinkela_buffer_10982 (
        .din(new_Jinkela_wire_13237),
        .dout(new_Jinkela_wire_13238)
    );

    bfr new_Jinkela_buffer_11062 (
        .din(new_Jinkela_wire_13335),
        .dout(new_Jinkela_wire_13336)
    );

    bfr new_Jinkela_buffer_10983 (
        .din(new_Jinkela_wire_13238),
        .dout(new_Jinkela_wire_13239)
    );

    bfr new_Jinkela_buffer_11060 (
        .din(new_Jinkela_wire_13329),
        .dout(new_Jinkela_wire_13330)
    );

    bfr new_Jinkela_buffer_10984 (
        .din(new_Jinkela_wire_13239),
        .dout(new_Jinkela_wire_13240)
    );

    bfr new_Jinkela_buffer_11070 (
        .din(_1663_),
        .dout(new_Jinkela_wire_13348)
    );

    spl2 new_Jinkela_splitter_987 (
        .a(_1554_),
        .b(new_Jinkela_wire_13342),
        .c(new_Jinkela_wire_13343)
    );

    bfr new_Jinkela_buffer_10985 (
        .din(new_Jinkela_wire_13240),
        .dout(new_Jinkela_wire_13241)
    );

    spl2 new_Jinkela_splitter_984 (
        .a(new_Jinkela_wire_13330),
        .b(new_Jinkela_wire_13331),
        .c(new_Jinkela_wire_13332)
    );

    bfr new_Jinkela_buffer_10986 (
        .din(new_Jinkela_wire_13241),
        .dout(new_Jinkela_wire_13242)
    );

    bfr new_Jinkela_buffer_10987 (
        .din(new_Jinkela_wire_13242),
        .dout(new_Jinkela_wire_13243)
    );

    bfr new_Jinkela_buffer_11063 (
        .din(new_Jinkela_wire_13336),
        .dout(new_Jinkela_wire_13337)
    );

    bfr new_Jinkela_buffer_10988 (
        .din(new_Jinkela_wire_13243),
        .dout(new_Jinkela_wire_13244)
    );

    bfr new_Jinkela_buffer_11064 (
        .din(new_Jinkela_wire_13337),
        .dout(new_Jinkela_wire_13338)
    );

    bfr new_Jinkela_buffer_10989 (
        .din(new_Jinkela_wire_13244),
        .dout(new_Jinkela_wire_13245)
    );

    bfr new_Jinkela_buffer_11071 (
        .din(new_net_3944),
        .dout(new_Jinkela_wire_13349)
    );

    bfr new_Jinkela_buffer_10990 (
        .din(new_Jinkela_wire_13245),
        .dout(new_Jinkela_wire_13246)
    );

    spl2 new_Jinkela_splitter_988 (
        .a(_1646_),
        .b(new_Jinkela_wire_13381),
        .c(new_Jinkela_wire_13382)
    );

    bfr new_Jinkela_buffer_10991 (
        .din(new_Jinkela_wire_13246),
        .dout(new_Jinkela_wire_13247)
    );

    bfr new_Jinkela_buffer_11067 (
        .din(new_Jinkela_wire_13344),
        .dout(new_Jinkela_wire_13345)
    );

    bfr new_Jinkela_buffer_10992 (
        .din(new_Jinkela_wire_13247),
        .dout(new_Jinkela_wire_13248)
    );

    spl2 new_Jinkela_splitter_989 (
        .a(_1468_),
        .b(new_Jinkela_wire_13387),
        .c(new_Jinkela_wire_13388)
    );

    bfr new_Jinkela_buffer_11072 (
        .din(new_Jinkela_wire_13349),
        .dout(new_Jinkela_wire_13350)
    );

    bfr new_Jinkela_buffer_10993 (
        .din(new_Jinkela_wire_13248),
        .dout(new_Jinkela_wire_13249)
    );

    bfr new_Jinkela_buffer_11068 (
        .din(new_Jinkela_wire_13345),
        .dout(new_Jinkela_wire_13346)
    );

    bfr new_Jinkela_buffer_10994 (
        .din(new_Jinkela_wire_13249),
        .dout(new_Jinkela_wire_13250)
    );

    bfr new_Jinkela_buffer_11103 (
        .din(new_Jinkela_wire_13382),
        .dout(new_Jinkela_wire_13383)
    );

    bfr new_Jinkela_buffer_10995 (
        .din(new_Jinkela_wire_13250),
        .dout(new_Jinkela_wire_13251)
    );

    bfr new_Jinkela_buffer_11069 (
        .din(new_Jinkela_wire_13346),
        .dout(new_Jinkela_wire_13347)
    );

    bfr new_Jinkela_buffer_10996 (
        .din(new_Jinkela_wire_13251),
        .dout(new_Jinkela_wire_13252)
    );

    bfr new_Jinkela_buffer_11073 (
        .din(new_Jinkela_wire_13350),
        .dout(new_Jinkela_wire_13351)
    );

    bfr new_Jinkela_buffer_10997 (
        .din(new_Jinkela_wire_13252),
        .dout(new_Jinkela_wire_13253)
    );

    bfr new_Jinkela_buffer_10998 (
        .din(new_Jinkela_wire_13253),
        .dout(new_Jinkela_wire_13254)
    );

    bfr new_Jinkela_buffer_11074 (
        .din(new_Jinkela_wire_13351),
        .dout(new_Jinkela_wire_13352)
    );

    bfr new_Jinkela_buffer_10999 (
        .din(new_Jinkela_wire_13254),
        .dout(new_Jinkela_wire_13255)
    );

    bfr new_Jinkela_buffer_14531 (
        .din(new_Jinkela_wire_17347),
        .dout(new_Jinkela_wire_17348)
    );

    bfr new_Jinkela_buffer_14402 (
        .din(new_Jinkela_wire_17216),
        .dout(new_Jinkela_wire_17217)
    );

    bfr new_Jinkela_buffer_14597 (
        .din(new_Jinkela_wire_17427),
        .dout(new_Jinkela_wire_17428)
    );

    bfr new_Jinkela_buffer_14403 (
        .din(new_Jinkela_wire_17217),
        .dout(new_Jinkela_wire_17218)
    );

    bfr new_Jinkela_buffer_14532 (
        .din(new_Jinkela_wire_17348),
        .dout(new_Jinkela_wire_17349)
    );

    bfr new_Jinkela_buffer_14404 (
        .din(new_Jinkela_wire_17218),
        .dout(new_Jinkela_wire_17219)
    );

    bfr new_Jinkela_buffer_14553 (
        .din(new_Jinkela_wire_17379),
        .dout(new_Jinkela_wire_17380)
    );

    bfr new_Jinkela_buffer_14405 (
        .din(new_Jinkela_wire_17219),
        .dout(new_Jinkela_wire_17220)
    );

    bfr new_Jinkela_buffer_14533 (
        .din(new_Jinkela_wire_17349),
        .dout(new_Jinkela_wire_17350)
    );

    bfr new_Jinkela_buffer_14406 (
        .din(new_Jinkela_wire_17220),
        .dout(new_Jinkela_wire_17221)
    );

    bfr new_Jinkela_buffer_14407 (
        .din(new_Jinkela_wire_17221),
        .dout(new_Jinkela_wire_17222)
    );

    bfr new_Jinkela_buffer_14534 (
        .din(new_Jinkela_wire_17350),
        .dout(new_Jinkela_wire_17351)
    );

    bfr new_Jinkela_buffer_14408 (
        .din(new_Jinkela_wire_17222),
        .dout(new_Jinkela_wire_17223)
    );

    bfr new_Jinkela_buffer_14554 (
        .din(new_Jinkela_wire_17380),
        .dout(new_Jinkela_wire_17381)
    );

    bfr new_Jinkela_buffer_14409 (
        .din(new_Jinkela_wire_17223),
        .dout(new_Jinkela_wire_17224)
    );

    bfr new_Jinkela_buffer_14535 (
        .din(new_Jinkela_wire_17351),
        .dout(new_Jinkela_wire_17352)
    );

    bfr new_Jinkela_buffer_14410 (
        .din(new_Jinkela_wire_17224),
        .dout(new_Jinkela_wire_17225)
    );

    bfr new_Jinkela_buffer_14598 (
        .din(new_Jinkela_wire_17428),
        .dout(new_Jinkela_wire_17429)
    );

    bfr new_Jinkela_buffer_14411 (
        .din(new_Jinkela_wire_17225),
        .dout(new_Jinkela_wire_17226)
    );

    bfr new_Jinkela_buffer_14536 (
        .din(new_Jinkela_wire_17352),
        .dout(new_Jinkela_wire_17353)
    );

    bfr new_Jinkela_buffer_14412 (
        .din(new_Jinkela_wire_17226),
        .dout(new_Jinkela_wire_17227)
    );

    bfr new_Jinkela_buffer_14555 (
        .din(new_Jinkela_wire_17381),
        .dout(new_Jinkela_wire_17382)
    );

    bfr new_Jinkela_buffer_14413 (
        .din(new_Jinkela_wire_17227),
        .dout(new_Jinkela_wire_17228)
    );

    bfr new_Jinkela_buffer_14537 (
        .din(new_Jinkela_wire_17353),
        .dout(new_Jinkela_wire_17354)
    );

    bfr new_Jinkela_buffer_14414 (
        .din(new_Jinkela_wire_17228),
        .dout(new_Jinkela_wire_17229)
    );

    bfr new_Jinkela_buffer_14415 (
        .din(new_Jinkela_wire_17229),
        .dout(new_Jinkela_wire_17230)
    );

    bfr new_Jinkela_buffer_14703 (
        .din(_1620_),
        .dout(new_Jinkela_wire_17542)
    );

    spl2 new_Jinkela_splitter_1257 (
        .a(new_Jinkela_wire_17354),
        .b(new_Jinkela_wire_17355),
        .c(new_Jinkela_wire_17356)
    );

    bfr new_Jinkela_buffer_14416 (
        .din(new_Jinkela_wire_17230),
        .dout(new_Jinkela_wire_17231)
    );

    bfr new_Jinkela_buffer_14599 (
        .din(new_Jinkela_wire_17429),
        .dout(new_Jinkela_wire_17430)
    );

    bfr new_Jinkela_buffer_14417 (
        .din(new_Jinkela_wire_17231),
        .dout(new_Jinkela_wire_17232)
    );

    bfr new_Jinkela_buffer_14556 (
        .din(new_Jinkela_wire_17382),
        .dout(new_Jinkela_wire_17383)
    );

    bfr new_Jinkela_buffer_14418 (
        .din(new_Jinkela_wire_17232),
        .dout(new_Jinkela_wire_17233)
    );

    bfr new_Jinkela_buffer_14557 (
        .din(new_Jinkela_wire_17383),
        .dout(new_Jinkela_wire_17384)
    );

    bfr new_Jinkela_buffer_14419 (
        .din(new_Jinkela_wire_17233),
        .dout(new_Jinkela_wire_17234)
    );

    bfr new_Jinkela_buffer_14699 (
        .din(new_Jinkela_wire_17537),
        .dout(new_Jinkela_wire_17538)
    );

    bfr new_Jinkela_buffer_14420 (
        .din(new_Jinkela_wire_17234),
        .dout(new_Jinkela_wire_17235)
    );

    spl2 new_Jinkela_splitter_1268 (
        .a(_1325_),
        .b(new_Jinkela_wire_17543),
        .c(new_Jinkela_wire_17544)
    );

    bfr new_Jinkela_buffer_14558 (
        .din(new_Jinkela_wire_17384),
        .dout(new_Jinkela_wire_17385)
    );

    bfr new_Jinkela_buffer_14421 (
        .din(new_Jinkela_wire_17235),
        .dout(new_Jinkela_wire_17236)
    );

    bfr new_Jinkela_buffer_14600 (
        .din(new_Jinkela_wire_17430),
        .dout(new_Jinkela_wire_17431)
    );

    bfr new_Jinkela_buffer_14422 (
        .din(new_Jinkela_wire_17236),
        .dout(new_Jinkela_wire_17237)
    );

    bfr new_Jinkela_buffer_7467 (
        .din(new_Jinkela_wire_9282),
        .dout(new_Jinkela_wire_9283)
    );

    bfr new_Jinkela_buffer_7557 (
        .din(new_Jinkela_wire_9380),
        .dout(new_Jinkela_wire_9381)
    );

    bfr new_Jinkela_buffer_7468 (
        .din(new_Jinkela_wire_9283),
        .dout(new_Jinkela_wire_9284)
    );

    bfr new_Jinkela_buffer_7686 (
        .din(new_Jinkela_wire_9513),
        .dout(new_Jinkela_wire_9514)
    );

    bfr new_Jinkela_buffer_7469 (
        .din(new_Jinkela_wire_9284),
        .dout(new_Jinkela_wire_9285)
    );

    bfr new_Jinkela_buffer_7558 (
        .din(new_Jinkela_wire_9381),
        .dout(new_Jinkela_wire_9382)
    );

    bfr new_Jinkela_buffer_7470 (
        .din(new_Jinkela_wire_9285),
        .dout(new_Jinkela_wire_9286)
    );

    bfr new_Jinkela_buffer_7628 (
        .din(new_Jinkela_wire_9455),
        .dout(new_Jinkela_wire_9456)
    );

    bfr new_Jinkela_buffer_7471 (
        .din(new_Jinkela_wire_9286),
        .dout(new_Jinkela_wire_9287)
    );

    bfr new_Jinkela_buffer_7559 (
        .din(new_Jinkela_wire_9382),
        .dout(new_Jinkela_wire_9383)
    );

    bfr new_Jinkela_buffer_7472 (
        .din(new_Jinkela_wire_9287),
        .dout(new_Jinkela_wire_9288)
    );

    bfr new_Jinkela_buffer_7692 (
        .din(new_Jinkela_wire_9523),
        .dout(new_Jinkela_wire_9524)
    );

    bfr new_Jinkela_buffer_7473 (
        .din(new_Jinkela_wire_9288),
        .dout(new_Jinkela_wire_9289)
    );

    bfr new_Jinkela_buffer_7560 (
        .din(new_Jinkela_wire_9383),
        .dout(new_Jinkela_wire_9384)
    );

    bfr new_Jinkela_buffer_7474 (
        .din(new_Jinkela_wire_9289),
        .dout(new_Jinkela_wire_9290)
    );

    bfr new_Jinkela_buffer_7629 (
        .din(new_Jinkela_wire_9456),
        .dout(new_Jinkela_wire_9457)
    );

    bfr new_Jinkela_buffer_7475 (
        .din(new_Jinkela_wire_9290),
        .dout(new_Jinkela_wire_9291)
    );

    bfr new_Jinkela_buffer_7561 (
        .din(new_Jinkela_wire_9384),
        .dout(new_Jinkela_wire_9385)
    );

    bfr new_Jinkela_buffer_7476 (
        .din(new_Jinkela_wire_9291),
        .dout(new_Jinkela_wire_9292)
    );

    bfr new_Jinkela_buffer_7687 (
        .din(new_Jinkela_wire_9514),
        .dout(new_Jinkela_wire_9515)
    );

    bfr new_Jinkela_buffer_7477 (
        .din(new_Jinkela_wire_9292),
        .dout(new_Jinkela_wire_9293)
    );

    bfr new_Jinkela_buffer_7562 (
        .din(new_Jinkela_wire_9385),
        .dout(new_Jinkela_wire_9386)
    );

    bfr new_Jinkela_buffer_7478 (
        .din(new_Jinkela_wire_9293),
        .dout(new_Jinkela_wire_9294)
    );

    bfr new_Jinkela_buffer_7630 (
        .din(new_Jinkela_wire_9457),
        .dout(new_Jinkela_wire_9458)
    );

    bfr new_Jinkela_buffer_7479 (
        .din(new_Jinkela_wire_9294),
        .dout(new_Jinkela_wire_9295)
    );

    bfr new_Jinkela_buffer_7563 (
        .din(new_Jinkela_wire_9386),
        .dout(new_Jinkela_wire_9387)
    );

    bfr new_Jinkela_buffer_7480 (
        .din(new_Jinkela_wire_9295),
        .dout(new_Jinkela_wire_9296)
    );

    bfr new_Jinkela_buffer_7707 (
        .din(_0757_),
        .dout(new_Jinkela_wire_9543)
    );

    spl2 new_Jinkela_splitter_766 (
        .a(_1407_),
        .b(new_Jinkela_wire_9541),
        .c(new_Jinkela_wire_9542)
    );

    spl2 new_Jinkela_splitter_757 (
        .a(new_Jinkela_wire_9296),
        .b(new_Jinkela_wire_9297),
        .c(new_Jinkela_wire_9298)
    );

    bfr new_Jinkela_buffer_7631 (
        .din(new_Jinkela_wire_9458),
        .dout(new_Jinkela_wire_9459)
    );

    bfr new_Jinkela_buffer_7564 (
        .din(new_Jinkela_wire_9387),
        .dout(new_Jinkela_wire_9388)
    );

    bfr new_Jinkela_buffer_7565 (
        .din(new_Jinkela_wire_9388),
        .dout(new_Jinkela_wire_9389)
    );

    bfr new_Jinkela_buffer_7688 (
        .din(new_Jinkela_wire_9515),
        .dout(new_Jinkela_wire_9516)
    );

    bfr new_Jinkela_buffer_7566 (
        .din(new_Jinkela_wire_9389),
        .dout(new_Jinkela_wire_9390)
    );

    bfr new_Jinkela_buffer_7632 (
        .din(new_Jinkela_wire_9459),
        .dout(new_Jinkela_wire_9460)
    );

    bfr new_Jinkela_buffer_7567 (
        .din(new_Jinkela_wire_9390),
        .dout(new_Jinkela_wire_9391)
    );

    bfr new_Jinkela_buffer_7693 (
        .din(new_Jinkela_wire_9524),
        .dout(new_Jinkela_wire_9525)
    );

    bfr new_Jinkela_buffer_7568 (
        .din(new_Jinkela_wire_9391),
        .dout(new_Jinkela_wire_9392)
    );

    bfr new_Jinkela_buffer_7633 (
        .din(new_Jinkela_wire_9460),
        .dout(new_Jinkela_wire_9461)
    );

    bfr new_Jinkela_buffer_7569 (
        .din(new_Jinkela_wire_9392),
        .dout(new_Jinkela_wire_9393)
    );

    bfr new_Jinkela_buffer_7689 (
        .din(new_Jinkela_wire_9516),
        .dout(new_Jinkela_wire_9517)
    );

    bfr new_Jinkela_buffer_7570 (
        .din(new_Jinkela_wire_9393),
        .dout(new_Jinkela_wire_9394)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_1393),
        .dout(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_17836 (
        .din(new_Jinkela_wire_21268),
        .dout(new_Jinkela_wire_21269)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_1181),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_11107 (
        .din(_1191_),
        .dout(new_Jinkela_wire_13389)
    );

    bfr new_Jinkela_buffer_11000 (
        .din(new_Jinkela_wire_13255),
        .dout(new_Jinkela_wire_13256)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_1296),
        .dout(new_Jinkela_wire_1297)
    );

    bfr new_Jinkela_buffer_17837 (
        .din(new_Jinkela_wire_21269),
        .dout(new_Jinkela_wire_21270)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_1182),
        .dout(new_Jinkela_wire_1183)
    );

    bfr new_Jinkela_buffer_11075 (
        .din(new_Jinkela_wire_13352),
        .dout(new_Jinkela_wire_13353)
    );

    bfr new_Jinkela_buffer_11001 (
        .din(new_Jinkela_wire_13256),
        .dout(new_Jinkela_wire_13257)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_1339),
        .dout(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_17838 (
        .din(new_Jinkela_wire_21270),
        .dout(new_Jinkela_wire_21271)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_1183),
        .dout(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_11002 (
        .din(new_Jinkela_wire_13257),
        .dout(new_Jinkela_wire_13258)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_1297),
        .dout(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_11104 (
        .din(new_Jinkela_wire_13383),
        .dout(new_Jinkela_wire_13384)
    );

    bfr new_Jinkela_buffer_17839 (
        .din(new_Jinkela_wire_21271),
        .dout(new_Jinkela_wire_21272)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_1184),
        .dout(new_Jinkela_wire_1185)
    );

    bfr new_Jinkela_buffer_11076 (
        .din(new_Jinkela_wire_13353),
        .dout(new_Jinkela_wire_13354)
    );

    bfr new_Jinkela_buffer_11003 (
        .din(new_Jinkela_wire_13258),
        .dout(new_Jinkela_wire_13259)
    );

    spl2 new_Jinkela_splitter_221 (
        .a(_0116_),
        .b(new_Jinkela_wire_1401),
        .c(new_Jinkela_wire_1402)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_net_3930),
        .dout(new_Jinkela_wire_1403)
    );

    bfr new_Jinkela_buffer_17840 (
        .din(new_Jinkela_wire_21272),
        .dout(new_Jinkela_wire_21273)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_1185),
        .dout(new_Jinkela_wire_1186)
    );

    bfr new_Jinkela_buffer_11004 (
        .din(new_Jinkela_wire_13259),
        .dout(new_Jinkela_wire_13260)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_1298),
        .dout(new_Jinkela_wire_1299)
    );

    spl2 new_Jinkela_splitter_991 (
        .a(_0224_),
        .b(new_Jinkela_wire_13392),
        .c(new_Jinkela_wire_13393)
    );

    bfr new_Jinkela_buffer_17841 (
        .din(new_Jinkela_wire_21273),
        .dout(new_Jinkela_wire_21274)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_1186),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_11077 (
        .din(new_Jinkela_wire_13354),
        .dout(new_Jinkela_wire_13355)
    );

    bfr new_Jinkela_buffer_11005 (
        .din(new_Jinkela_wire_13260),
        .dout(new_Jinkela_wire_13261)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_1340),
        .dout(new_Jinkela_wire_1341)
    );

    bfr new_Jinkela_buffer_17842 (
        .din(new_Jinkela_wire_21274),
        .dout(new_Jinkela_wire_21275)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_1187),
        .dout(new_Jinkela_wire_1188)
    );

    spl2 new_Jinkela_splitter_990 (
        .a(_0859_),
        .b(new_Jinkela_wire_13390),
        .c(new_Jinkela_wire_13391)
    );

    bfr new_Jinkela_buffer_11006 (
        .din(new_Jinkela_wire_13261),
        .dout(new_Jinkela_wire_13262)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_1299),
        .dout(new_Jinkela_wire_1300)
    );

    bfr new_Jinkela_buffer_11105 (
        .din(new_Jinkela_wire_13384),
        .dout(new_Jinkela_wire_13385)
    );

    bfr new_Jinkela_buffer_17843 (
        .din(new_Jinkela_wire_21275),
        .dout(new_Jinkela_wire_21276)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_1188),
        .dout(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_11078 (
        .din(new_Jinkela_wire_13355),
        .dout(new_Jinkela_wire_13356)
    );

    bfr new_Jinkela_buffer_11007 (
        .din(new_Jinkela_wire_13262),
        .dout(new_Jinkela_wire_13263)
    );

    bfr new_Jinkela_buffer_821 (
        .din(_1143_),
        .dout(new_Jinkela_wire_1567)
    );

    bfr new_Jinkela_buffer_17844 (
        .din(new_Jinkela_wire_21276),
        .dout(new_Jinkela_wire_21277)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_1189),
        .dout(new_Jinkela_wire_1190)
    );

    bfr new_Jinkela_buffer_11008 (
        .din(new_Jinkela_wire_13263),
        .dout(new_Jinkela_wire_13264)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_1300),
        .dout(new_Jinkela_wire_1301)
    );

    bfr new_Jinkela_buffer_17845 (
        .din(new_Jinkela_wire_21277),
        .dout(new_Jinkela_wire_21278)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_1190),
        .dout(new_Jinkela_wire_1191)
    );

    bfr new_Jinkela_buffer_11079 (
        .din(new_Jinkela_wire_13356),
        .dout(new_Jinkela_wire_13357)
    );

    bfr new_Jinkela_buffer_11009 (
        .din(new_Jinkela_wire_13264),
        .dout(new_Jinkela_wire_13265)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_1341),
        .dout(new_Jinkela_wire_1342)
    );

    bfr new_Jinkela_buffer_17846 (
        .din(new_Jinkela_wire_21278),
        .dout(new_Jinkela_wire_21279)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_1191),
        .dout(new_Jinkela_wire_1192)
    );

    bfr new_Jinkela_buffer_11010 (
        .din(new_Jinkela_wire_13265),
        .dout(new_Jinkela_wire_13266)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_1301),
        .dout(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_11106 (
        .din(new_Jinkela_wire_13385),
        .dout(new_Jinkela_wire_13386)
    );

    bfr new_Jinkela_buffer_17847 (
        .din(new_Jinkela_wire_21279),
        .dout(new_Jinkela_wire_21280)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_1192),
        .dout(new_Jinkela_wire_1193)
    );

    bfr new_Jinkela_buffer_11080 (
        .din(new_Jinkela_wire_13357),
        .dout(new_Jinkela_wire_13358)
    );

    bfr new_Jinkela_buffer_11011 (
        .din(new_Jinkela_wire_13266),
        .dout(new_Jinkela_wire_13267)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(_0850_),
        .b(new_Jinkela_wire_1570),
        .c(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_1394),
        .dout(new_Jinkela_wire_1395)
    );

    bfr new_Jinkela_buffer_17848 (
        .din(new_Jinkela_wire_21280),
        .dout(new_Jinkela_wire_21281)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_1193),
        .dout(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_11012 (
        .din(new_Jinkela_wire_13267),
        .dout(new_Jinkela_wire_13268)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_1302),
        .dout(new_Jinkela_wire_1303)
    );

    bfr new_Jinkela_buffer_17849 (
        .din(new_Jinkela_wire_21281),
        .dout(new_Jinkela_wire_21282)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_1194),
        .dout(new_Jinkela_wire_1195)
    );

    bfr new_Jinkela_buffer_11081 (
        .din(new_Jinkela_wire_13358),
        .dout(new_Jinkela_wire_13359)
    );

    bfr new_Jinkela_buffer_11013 (
        .din(new_Jinkela_wire_13268),
        .dout(new_Jinkela_wire_13269)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_1342),
        .dout(new_Jinkela_wire_1343)
    );

    bfr new_Jinkela_buffer_17850 (
        .din(new_Jinkela_wire_21282),
        .dout(new_Jinkela_wire_21283)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_1195),
        .dout(new_Jinkela_wire_1196)
    );

    spl2 new_Jinkela_splitter_992 (
        .a(_0295_),
        .b(new_Jinkela_wire_13394),
        .c(new_Jinkela_wire_13395)
    );

    bfr new_Jinkela_buffer_11014 (
        .din(new_Jinkela_wire_13269),
        .dout(new_Jinkela_wire_13270)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_1303),
        .dout(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_17851 (
        .din(new_Jinkela_wire_21283),
        .dout(new_Jinkela_wire_21284)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_1196),
        .dout(new_Jinkela_wire_1197)
    );

    bfr new_Jinkela_buffer_11082 (
        .din(new_Jinkela_wire_13359),
        .dout(new_Jinkela_wire_13360)
    );

    bfr new_Jinkela_buffer_11015 (
        .din(new_Jinkela_wire_13270),
        .dout(new_Jinkela_wire_13271)
    );

    bfr new_Jinkela_buffer_17852 (
        .din(new_Jinkela_wire_21284),
        .dout(new_Jinkela_wire_21285)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_1197),
        .dout(new_Jinkela_wire_1198)
    );

    spl2 new_Jinkela_splitter_993 (
        .a(_1480_),
        .b(new_Jinkela_wire_13396),
        .c(new_Jinkela_wire_13397)
    );

    bfr new_Jinkela_buffer_11016 (
        .din(new_Jinkela_wire_13271),
        .dout(new_Jinkela_wire_13272)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_1304),
        .dout(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_17853 (
        .din(new_Jinkela_wire_21285),
        .dout(new_Jinkela_wire_21286)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_1198),
        .dout(new_Jinkela_wire_1199)
    );

    bfr new_Jinkela_buffer_11083 (
        .din(new_Jinkela_wire_13360),
        .dout(new_Jinkela_wire_13361)
    );

    bfr new_Jinkela_buffer_11017 (
        .din(new_Jinkela_wire_13272),
        .dout(new_Jinkela_wire_13273)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_1343),
        .dout(new_Jinkela_wire_1344)
    );

    bfr new_Jinkela_buffer_17854 (
        .din(new_Jinkela_wire_21286),
        .dout(new_Jinkela_wire_21287)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_1199),
        .dout(new_Jinkela_wire_1200)
    );

    spl2 new_Jinkela_splitter_994 (
        .a(_0836_),
        .b(new_Jinkela_wire_13398),
        .c(new_Jinkela_wire_13399)
    );

    bfr new_Jinkela_buffer_11018 (
        .din(new_Jinkela_wire_13273),
        .dout(new_Jinkela_wire_13274)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_1305),
        .dout(new_Jinkela_wire_1306)
    );

    spl2 new_Jinkela_splitter_996 (
        .a(_0528_),
        .b(new_Jinkela_wire_13402),
        .c(new_Jinkela_wire_13403)
    );

    bfr new_Jinkela_buffer_17855 (
        .din(new_Jinkela_wire_21287),
        .dout(new_Jinkela_wire_21288)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_1200),
        .dout(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_11084 (
        .din(new_Jinkela_wire_13361),
        .dout(new_Jinkela_wire_13362)
    );

    bfr new_Jinkela_buffer_11019 (
        .din(new_Jinkela_wire_13274),
        .dout(new_Jinkela_wire_13275)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    bfr new_Jinkela_buffer_17856 (
        .din(new_Jinkela_wire_21288),
        .dout(new_Jinkela_wire_21289)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_1201),
        .dout(new_Jinkela_wire_1202)
    );

    spl2 new_Jinkela_splitter_995 (
        .a(_1434_),
        .b(new_Jinkela_wire_13400),
        .c(new_Jinkela_wire_13401)
    );

    bfr new_Jinkela_buffer_11020 (
        .din(new_Jinkela_wire_13275),
        .dout(new_Jinkela_wire_13276)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_1306),
        .dout(new_Jinkela_wire_1307)
    );

    bfr new_Jinkela_buffer_14559 (
        .din(new_Jinkela_wire_17385),
        .dout(new_Jinkela_wire_17386)
    );

    bfr new_Jinkela_buffer_14423 (
        .din(new_Jinkela_wire_17237),
        .dout(new_Jinkela_wire_17238)
    );

    spl2 new_Jinkela_splitter_1269 (
        .a(_1764_),
        .b(new_Jinkela_wire_17545),
        .c(new_Jinkela_wire_17546)
    );

    bfr new_Jinkela_buffer_14424 (
        .din(new_Jinkela_wire_17238),
        .dout(new_Jinkela_wire_17239)
    );

    spl2 new_Jinkela_splitter_1271 (
        .a(_0762_),
        .b(new_Jinkela_wire_17549),
        .c(new_Jinkela_wire_17550)
    );

    bfr new_Jinkela_buffer_14560 (
        .din(new_Jinkela_wire_17386),
        .dout(new_Jinkela_wire_17387)
    );

    bfr new_Jinkela_buffer_14425 (
        .din(new_Jinkela_wire_17239),
        .dout(new_Jinkela_wire_17240)
    );

    bfr new_Jinkela_buffer_14601 (
        .din(new_Jinkela_wire_17431),
        .dout(new_Jinkela_wire_17432)
    );

    bfr new_Jinkela_buffer_14426 (
        .din(new_Jinkela_wire_17240),
        .dout(new_Jinkela_wire_17241)
    );

    bfr new_Jinkela_buffer_14561 (
        .din(new_Jinkela_wire_17387),
        .dout(new_Jinkela_wire_17388)
    );

    bfr new_Jinkela_buffer_14427 (
        .din(new_Jinkela_wire_17241),
        .dout(new_Jinkela_wire_17242)
    );

    bfr new_Jinkela_buffer_14700 (
        .din(new_Jinkela_wire_17538),
        .dout(new_Jinkela_wire_17539)
    );

    bfr new_Jinkela_buffer_14428 (
        .din(new_Jinkela_wire_17242),
        .dout(new_Jinkela_wire_17243)
    );

    bfr new_Jinkela_buffer_14562 (
        .din(new_Jinkela_wire_17388),
        .dout(new_Jinkela_wire_17389)
    );

    bfr new_Jinkela_buffer_14429 (
        .din(new_Jinkela_wire_17243),
        .dout(new_Jinkela_wire_17244)
    );

    bfr new_Jinkela_buffer_14602 (
        .din(new_Jinkela_wire_17432),
        .dout(new_Jinkela_wire_17433)
    );

    bfr new_Jinkela_buffer_14430 (
        .din(new_Jinkela_wire_17244),
        .dout(new_Jinkela_wire_17245)
    );

    bfr new_Jinkela_buffer_14563 (
        .din(new_Jinkela_wire_17389),
        .dout(new_Jinkela_wire_17390)
    );

    bfr new_Jinkela_buffer_14431 (
        .din(new_Jinkela_wire_17245),
        .dout(new_Jinkela_wire_17246)
    );

    bfr new_Jinkela_buffer_14432 (
        .din(new_Jinkela_wire_17246),
        .dout(new_Jinkela_wire_17247)
    );

    bfr new_Jinkela_buffer_14564 (
        .din(new_Jinkela_wire_17390),
        .dout(new_Jinkela_wire_17391)
    );

    bfr new_Jinkela_buffer_14433 (
        .din(new_Jinkela_wire_17247),
        .dout(new_Jinkela_wire_17248)
    );

    bfr new_Jinkela_buffer_14603 (
        .din(new_Jinkela_wire_17433),
        .dout(new_Jinkela_wire_17434)
    );

    bfr new_Jinkela_buffer_14434 (
        .din(new_Jinkela_wire_17248),
        .dout(new_Jinkela_wire_17249)
    );

    bfr new_Jinkela_buffer_14565 (
        .din(new_Jinkela_wire_17391),
        .dout(new_Jinkela_wire_17392)
    );

    bfr new_Jinkela_buffer_14435 (
        .din(new_Jinkela_wire_17249),
        .dout(new_Jinkela_wire_17250)
    );

    bfr new_Jinkela_buffer_14701 (
        .din(new_Jinkela_wire_17539),
        .dout(new_Jinkela_wire_17540)
    );

    bfr new_Jinkela_buffer_14436 (
        .din(new_Jinkela_wire_17250),
        .dout(new_Jinkela_wire_17251)
    );

    bfr new_Jinkela_buffer_14566 (
        .din(new_Jinkela_wire_17392),
        .dout(new_Jinkela_wire_17393)
    );

    bfr new_Jinkela_buffer_14437 (
        .din(new_Jinkela_wire_17251),
        .dout(new_Jinkela_wire_17252)
    );

    bfr new_Jinkela_buffer_14604 (
        .din(new_Jinkela_wire_17434),
        .dout(new_Jinkela_wire_17435)
    );

    bfr new_Jinkela_buffer_14438 (
        .din(new_Jinkela_wire_17252),
        .dout(new_Jinkela_wire_17253)
    );

    bfr new_Jinkela_buffer_14567 (
        .din(new_Jinkela_wire_17393),
        .dout(new_Jinkela_wire_17394)
    );

    bfr new_Jinkela_buffer_14439 (
        .din(new_Jinkela_wire_17253),
        .dout(new_Jinkela_wire_17254)
    );

    bfr new_Jinkela_buffer_14440 (
        .din(new_Jinkela_wire_17254),
        .dout(new_Jinkela_wire_17255)
    );

    spl2 new_Jinkela_splitter_1270 (
        .a(_0289_),
        .b(new_Jinkela_wire_17547),
        .c(new_Jinkela_wire_17548)
    );

    bfr new_Jinkela_buffer_14568 (
        .din(new_Jinkela_wire_17394),
        .dout(new_Jinkela_wire_17395)
    );

    bfr new_Jinkela_buffer_14441 (
        .din(new_Jinkela_wire_17255),
        .dout(new_Jinkela_wire_17256)
    );

    bfr new_Jinkela_buffer_14605 (
        .din(new_Jinkela_wire_17435),
        .dout(new_Jinkela_wire_17436)
    );

    bfr new_Jinkela_buffer_14442 (
        .din(new_Jinkela_wire_17256),
        .dout(new_Jinkela_wire_17257)
    );

    bfr new_Jinkela_buffer_14569 (
        .din(new_Jinkela_wire_17395),
        .dout(new_Jinkela_wire_17396)
    );

    bfr new_Jinkela_buffer_14443 (
        .din(new_Jinkela_wire_17257),
        .dout(new_Jinkela_wire_17258)
    );

    bfr new_Jinkela_buffer_17857 (
        .din(new_Jinkela_wire_21289),
        .dout(new_Jinkela_wire_21290)
    );

    bfr new_Jinkela_buffer_17858 (
        .din(new_Jinkela_wire_21290),
        .dout(new_Jinkela_wire_21291)
    );

    bfr new_Jinkela_buffer_17859 (
        .din(new_Jinkela_wire_21291),
        .dout(new_Jinkela_wire_21292)
    );

    bfr new_Jinkela_buffer_17860 (
        .din(new_Jinkela_wire_21292),
        .dout(new_Jinkela_wire_21293)
    );

    bfr new_Jinkela_buffer_17861 (
        .din(new_Jinkela_wire_21293),
        .dout(new_Jinkela_wire_21294)
    );

    bfr new_Jinkela_buffer_17862 (
        .din(new_Jinkela_wire_21294),
        .dout(new_Jinkela_wire_21295)
    );

    bfr new_Jinkela_buffer_17863 (
        .din(new_Jinkela_wire_21295),
        .dout(new_Jinkela_wire_21296)
    );

    bfr new_Jinkela_buffer_17864 (
        .din(new_Jinkela_wire_21296),
        .dout(new_Jinkela_wire_21297)
    );

    bfr new_Jinkela_buffer_17865 (
        .din(new_Jinkela_wire_21297),
        .dout(new_Jinkela_wire_21298)
    );

    bfr new_Jinkela_buffer_17866 (
        .din(new_Jinkela_wire_21298),
        .dout(new_Jinkela_wire_21299)
    );

    bfr new_Jinkela_buffer_17867 (
        .din(new_Jinkela_wire_21299),
        .dout(new_Jinkela_wire_21300)
    );

    bfr new_Jinkela_buffer_17868 (
        .din(new_Jinkela_wire_21300),
        .dout(new_Jinkela_wire_21301)
    );

    bfr new_Jinkela_buffer_17869 (
        .din(new_Jinkela_wire_21301),
        .dout(new_Jinkela_wire_21302)
    );

    bfr new_Jinkela_buffer_17870 (
        .din(new_Jinkela_wire_21302),
        .dout(new_Jinkela_wire_21303)
    );

    bfr new_Jinkela_buffer_17871 (
        .din(new_Jinkela_wire_21303),
        .dout(new_Jinkela_wire_21304)
    );

    bfr new_Jinkela_buffer_17872 (
        .din(new_Jinkela_wire_21304),
        .dout(new_Jinkela_wire_21305)
    );

    bfr new_Jinkela_buffer_17873 (
        .din(new_Jinkela_wire_21305),
        .dout(new_Jinkela_wire_21306)
    );

    bfr new_Jinkela_buffer_17874 (
        .din(new_Jinkela_wire_21306),
        .dout(new_Jinkela_wire_21307)
    );

    bfr new_Jinkela_buffer_17875 (
        .din(new_Jinkela_wire_21307),
        .dout(new_Jinkela_wire_21308)
    );

    bfr new_Jinkela_buffer_17876 (
        .din(new_Jinkela_wire_21308),
        .dout(new_Jinkela_wire_21309)
    );

    bfr new_Jinkela_buffer_17877 (
        .din(new_Jinkela_wire_21309),
        .dout(new_Jinkela_wire_21310)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_1202),
        .dout(new_Jinkela_wire_1203)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_1344),
        .dout(new_Jinkela_wire_1345)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_1203),
        .dout(new_Jinkela_wire_1204)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_1307),
        .dout(new_Jinkela_wire_1308)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_1204),
        .dout(new_Jinkela_wire_1205)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_1403),
        .dout(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_1205),
        .dout(new_Jinkela_wire_1206)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_1308),
        .dout(new_Jinkela_wire_1309)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_1206),
        .dout(new_Jinkela_wire_1207)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_1345),
        .dout(new_Jinkela_wire_1346)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_1207),
        .dout(new_Jinkela_wire_1208)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_1309),
        .dout(new_Jinkela_wire_1310)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_1208),
        .dout(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_1396),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_1209),
        .dout(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_1310),
        .dout(new_Jinkela_wire_1311)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_1210),
        .dout(new_Jinkela_wire_1211)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_1346),
        .dout(new_Jinkela_wire_1347)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_1211),
        .dout(new_Jinkela_wire_1212)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_1311),
        .dout(new_Jinkela_wire_1312)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_1212),
        .dout(new_Jinkela_wire_1213)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_1213),
        .dout(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_1312),
        .dout(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_1214),
        .dout(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_1347),
        .dout(new_Jinkela_wire_1348)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_1215),
        .dout(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_1313),
        .dout(new_Jinkela_wire_1314)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_1217),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_1314),
        .dout(new_Jinkela_wire_1315)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_1218),
        .dout(new_Jinkela_wire_1219)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_1348),
        .dout(new_Jinkela_wire_1349)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_1219),
        .dout(new_Jinkela_wire_1220)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_1315),
        .dout(new_Jinkela_wire_1316)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_1404),
        .dout(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_1316),
        .dout(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_1222),
        .dout(new_Jinkela_wire_1223)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_1349),
        .dout(new_Jinkela_wire_1350)
    );

    bfr new_Jinkela_buffer_11085 (
        .din(new_Jinkela_wire_13362),
        .dout(new_Jinkela_wire_13363)
    );

    bfr new_Jinkela_buffer_11021 (
        .din(new_Jinkela_wire_13276),
        .dout(new_Jinkela_wire_13277)
    );

    bfr new_Jinkela_buffer_4095 (
        .din(new_Jinkela_wire_5370),
        .dout(new_Jinkela_wire_5371)
    );

    spl2 new_Jinkela_splitter_508 (
        .a(_1432_),
        .b(new_Jinkela_wire_5544),
        .c(new_Jinkela_wire_5545)
    );

    bfr new_Jinkela_buffer_4162 (
        .din(new_Jinkela_wire_5473),
        .dout(new_Jinkela_wire_5474)
    );

    bfr new_Jinkela_buffer_11022 (
        .din(new_Jinkela_wire_13277),
        .dout(new_Jinkela_wire_13278)
    );

    bfr new_Jinkela_buffer_4096 (
        .din(new_Jinkela_wire_5371),
        .dout(new_Jinkela_wire_5372)
    );

    bfr new_Jinkela_buffer_11086 (
        .din(new_Jinkela_wire_13363),
        .dout(new_Jinkela_wire_13364)
    );

    bfr new_Jinkela_buffer_11023 (
        .din(new_Jinkela_wire_13278),
        .dout(new_Jinkela_wire_13279)
    );

    bfr new_Jinkela_buffer_4097 (
        .din(new_Jinkela_wire_5372),
        .dout(new_Jinkela_wire_5373)
    );

    bfr new_Jinkela_buffer_4163 (
        .din(new_Jinkela_wire_5474),
        .dout(new_Jinkela_wire_5475)
    );

    spl2 new_Jinkela_splitter_997 (
        .a(_0114_),
        .b(new_Jinkela_wire_13404),
        .c(new_Jinkela_wire_13405)
    );

    bfr new_Jinkela_buffer_11024 (
        .din(new_Jinkela_wire_13279),
        .dout(new_Jinkela_wire_13280)
    );

    bfr new_Jinkela_buffer_4098 (
        .din(new_Jinkela_wire_5373),
        .dout(new_Jinkela_wire_5374)
    );

    spl2 new_Jinkela_splitter_509 (
        .a(_1035_),
        .b(new_Jinkela_wire_5546),
        .c(new_Jinkela_wire_5547)
    );

    bfr new_Jinkela_buffer_11087 (
        .din(new_Jinkela_wire_13364),
        .dout(new_Jinkela_wire_13365)
    );

    bfr new_Jinkela_buffer_11025 (
        .din(new_Jinkela_wire_13280),
        .dout(new_Jinkela_wire_13281)
    );

    bfr new_Jinkela_buffer_4099 (
        .din(new_Jinkela_wire_5374),
        .dout(new_Jinkela_wire_5375)
    );

    bfr new_Jinkela_buffer_4164 (
        .din(new_Jinkela_wire_5475),
        .dout(new_Jinkela_wire_5476)
    );

    bfr new_Jinkela_buffer_11112 (
        .din(_1729_),
        .dout(new_Jinkela_wire_13410)
    );

    bfr new_Jinkela_buffer_11026 (
        .din(new_Jinkela_wire_13281),
        .dout(new_Jinkela_wire_13282)
    );

    bfr new_Jinkela_buffer_4100 (
        .din(new_Jinkela_wire_5375),
        .dout(new_Jinkela_wire_5376)
    );

    bfr new_Jinkela_buffer_11108 (
        .din(new_Jinkela_wire_13405),
        .dout(new_Jinkela_wire_13406)
    );

    spl2 new_Jinkela_splitter_510 (
        .a(_0765_),
        .b(new_Jinkela_wire_5548),
        .c(new_Jinkela_wire_5549)
    );

    bfr new_Jinkela_buffer_11088 (
        .din(new_Jinkela_wire_13365),
        .dout(new_Jinkela_wire_13366)
    );

    bfr new_Jinkela_buffer_11027 (
        .din(new_Jinkela_wire_13282),
        .dout(new_Jinkela_wire_13283)
    );

    bfr new_Jinkela_buffer_4101 (
        .din(new_Jinkela_wire_5376),
        .dout(new_Jinkela_wire_5377)
    );

    spl2 new_Jinkela_splitter_512 (
        .a(_0545_),
        .b(new_Jinkela_wire_5665),
        .c(new_Jinkela_wire_5666)
    );

    bfr new_Jinkela_buffer_4165 (
        .din(new_Jinkela_wire_5476),
        .dout(new_Jinkela_wire_5477)
    );

    bfr new_Jinkela_buffer_11113 (
        .din(new_net_3934),
        .dout(new_Jinkela_wire_13411)
    );

    bfr new_Jinkela_buffer_11028 (
        .din(new_Jinkela_wire_13283),
        .dout(new_Jinkela_wire_13284)
    );

    bfr new_Jinkela_buffer_4102 (
        .din(new_Jinkela_wire_5377),
        .dout(new_Jinkela_wire_5378)
    );

    bfr new_Jinkela_buffer_4226 (
        .din(_0212_),
        .dout(new_Jinkela_wire_5550)
    );

    bfr new_Jinkela_buffer_11089 (
        .din(new_Jinkela_wire_13366),
        .dout(new_Jinkela_wire_13367)
    );

    bfr new_Jinkela_buffer_11029 (
        .din(new_Jinkela_wire_13284),
        .dout(new_Jinkela_wire_13285)
    );

    bfr new_Jinkela_buffer_4103 (
        .din(new_Jinkela_wire_5378),
        .dout(new_Jinkela_wire_5379)
    );

    bfr new_Jinkela_buffer_4166 (
        .din(new_Jinkela_wire_5477),
        .dout(new_Jinkela_wire_5478)
    );

    bfr new_Jinkela_buffer_11157 (
        .din(_0026_),
        .dout(new_Jinkela_wire_13455)
    );

    bfr new_Jinkela_buffer_11030 (
        .din(new_Jinkela_wire_13285),
        .dout(new_Jinkela_wire_13286)
    );

    bfr new_Jinkela_buffer_4104 (
        .din(new_Jinkela_wire_5379),
        .dout(new_Jinkela_wire_5380)
    );

    bfr new_Jinkela_buffer_11109 (
        .din(new_Jinkela_wire_13406),
        .dout(new_Jinkela_wire_13407)
    );

    bfr new_Jinkela_buffer_4338 (
        .din(_0046_),
        .dout(new_Jinkela_wire_5664)
    );

    bfr new_Jinkela_buffer_11090 (
        .din(new_Jinkela_wire_13367),
        .dout(new_Jinkela_wire_13368)
    );

    bfr new_Jinkela_buffer_11031 (
        .din(new_Jinkela_wire_13286),
        .dout(new_Jinkela_wire_13287)
    );

    bfr new_Jinkela_buffer_4105 (
        .din(new_Jinkela_wire_5380),
        .dout(new_Jinkela_wire_5381)
    );

    bfr new_Jinkela_buffer_4227 (
        .din(new_Jinkela_wire_5550),
        .dout(new_Jinkela_wire_5551)
    );

    bfr new_Jinkela_buffer_4167 (
        .din(new_Jinkela_wire_5478),
        .dout(new_Jinkela_wire_5479)
    );

    bfr new_Jinkela_buffer_11032 (
        .din(new_Jinkela_wire_13287),
        .dout(new_Jinkela_wire_13288)
    );

    bfr new_Jinkela_buffer_4106 (
        .din(new_Jinkela_wire_5381),
        .dout(new_Jinkela_wire_5382)
    );

    bfr new_Jinkela_buffer_11091 (
        .din(new_Jinkela_wire_13368),
        .dout(new_Jinkela_wire_13369)
    );

    bfr new_Jinkela_buffer_11033 (
        .din(new_Jinkela_wire_13288),
        .dout(new_Jinkela_wire_13289)
    );

    bfr new_Jinkela_buffer_4107 (
        .din(new_Jinkela_wire_5382),
        .dout(new_Jinkela_wire_5383)
    );

    spl2 new_Jinkela_splitter_513 (
        .a(_0424_),
        .b(new_Jinkela_wire_5667),
        .c(new_Jinkela_wire_5668)
    );

    bfr new_Jinkela_buffer_4168 (
        .din(new_Jinkela_wire_5479),
        .dout(new_Jinkela_wire_5480)
    );

    bfr new_Jinkela_buffer_11114 (
        .din(new_Jinkela_wire_13411),
        .dout(new_Jinkela_wire_13412)
    );

    bfr new_Jinkela_buffer_11034 (
        .din(new_Jinkela_wire_13289),
        .dout(new_Jinkela_wire_13290)
    );

    bfr new_Jinkela_buffer_4108 (
        .din(new_Jinkela_wire_5383),
        .dout(new_Jinkela_wire_5384)
    );

    bfr new_Jinkela_buffer_11110 (
        .din(new_Jinkela_wire_13407),
        .dout(new_Jinkela_wire_13408)
    );

    bfr new_Jinkela_buffer_11092 (
        .din(new_Jinkela_wire_13369),
        .dout(new_Jinkela_wire_13370)
    );

    bfr new_Jinkela_buffer_11035 (
        .din(new_Jinkela_wire_13290),
        .dout(new_Jinkela_wire_13291)
    );

    bfr new_Jinkela_buffer_4109 (
        .din(new_Jinkela_wire_5384),
        .dout(new_Jinkela_wire_5385)
    );

    bfr new_Jinkela_buffer_4228 (
        .din(new_Jinkela_wire_5551),
        .dout(new_Jinkela_wire_5552)
    );

    bfr new_Jinkela_buffer_4169 (
        .din(new_Jinkela_wire_5480),
        .dout(new_Jinkela_wire_5481)
    );

    bfr new_Jinkela_buffer_11036 (
        .din(new_Jinkela_wire_13291),
        .dout(new_Jinkela_wire_13292)
    );

    bfr new_Jinkela_buffer_4110 (
        .din(new_Jinkela_wire_5385),
        .dout(new_Jinkela_wire_5386)
    );

    bfr new_Jinkela_buffer_11093 (
        .din(new_Jinkela_wire_13370),
        .dout(new_Jinkela_wire_13371)
    );

    bfr new_Jinkela_buffer_11037 (
        .din(new_Jinkela_wire_13292),
        .dout(new_Jinkela_wire_13293)
    );

    bfr new_Jinkela_buffer_4111 (
        .din(new_Jinkela_wire_5386),
        .dout(new_Jinkela_wire_5387)
    );

    spl2 new_Jinkela_splitter_514 (
        .a(_1368_),
        .b(new_Jinkela_wire_5681),
        .c(new_Jinkela_wire_5682)
    );

    bfr new_Jinkela_buffer_4170 (
        .din(new_Jinkela_wire_5481),
        .dout(new_Jinkela_wire_5482)
    );

    bfr new_Jinkela_buffer_11158 (
        .din(_0240_),
        .dout(new_Jinkela_wire_13456)
    );

    bfr new_Jinkela_buffer_11038 (
        .din(new_Jinkela_wire_13293),
        .dout(new_Jinkela_wire_13294)
    );

    bfr new_Jinkela_buffer_4112 (
        .din(new_Jinkela_wire_5387),
        .dout(new_Jinkela_wire_5388)
    );

    bfr new_Jinkela_buffer_11111 (
        .din(new_Jinkela_wire_13408),
        .dout(new_Jinkela_wire_13409)
    );

    bfr new_Jinkela_buffer_11094 (
        .din(new_Jinkela_wire_13371),
        .dout(new_Jinkela_wire_13372)
    );

    bfr new_Jinkela_buffer_11039 (
        .din(new_Jinkela_wire_13294),
        .dout(new_Jinkela_wire_13295)
    );

    bfr new_Jinkela_buffer_4113 (
        .din(new_Jinkela_wire_5388),
        .dout(new_Jinkela_wire_5389)
    );

    bfr new_Jinkela_buffer_4229 (
        .din(new_Jinkela_wire_5552),
        .dout(new_Jinkela_wire_5553)
    );

    bfr new_Jinkela_buffer_4171 (
        .din(new_Jinkela_wire_5482),
        .dout(new_Jinkela_wire_5483)
    );

    bfr new_Jinkela_buffer_11040 (
        .din(new_Jinkela_wire_13295),
        .dout(new_Jinkela_wire_13296)
    );

    bfr new_Jinkela_buffer_4114 (
        .din(new_Jinkela_wire_5389),
        .dout(new_Jinkela_wire_5390)
    );

    bfr new_Jinkela_buffer_11095 (
        .din(new_Jinkela_wire_13372),
        .dout(new_Jinkela_wire_13373)
    );

    bfr new_Jinkela_buffer_11041 (
        .din(new_Jinkela_wire_13296),
        .dout(new_Jinkela_wire_13297)
    );

    bfr new_Jinkela_buffer_4115 (
        .din(new_Jinkela_wire_5390),
        .dout(new_Jinkela_wire_5391)
    );

    bfr new_Jinkela_buffer_14702 (
        .din(new_Jinkela_wire_17540),
        .dout(new_Jinkela_wire_17541)
    );

    bfr new_Jinkela_buffer_14444 (
        .din(new_Jinkela_wire_17258),
        .dout(new_Jinkela_wire_17259)
    );

    bfr new_Jinkela_buffer_14570 (
        .din(new_Jinkela_wire_17396),
        .dout(new_Jinkela_wire_17397)
    );

    bfr new_Jinkela_buffer_14445 (
        .din(new_Jinkela_wire_17259),
        .dout(new_Jinkela_wire_17260)
    );

    bfr new_Jinkela_buffer_14606 (
        .din(new_Jinkela_wire_17436),
        .dout(new_Jinkela_wire_17437)
    );

    bfr new_Jinkela_buffer_14446 (
        .din(new_Jinkela_wire_17260),
        .dout(new_Jinkela_wire_17261)
    );

    bfr new_Jinkela_buffer_14571 (
        .din(new_Jinkela_wire_17397),
        .dout(new_Jinkela_wire_17398)
    );

    bfr new_Jinkela_buffer_14447 (
        .din(new_Jinkela_wire_17261),
        .dout(new_Jinkela_wire_17262)
    );

    bfr new_Jinkela_buffer_14448 (
        .din(new_Jinkela_wire_17262),
        .dout(new_Jinkela_wire_17263)
    );

    bfr new_Jinkela_buffer_14572 (
        .din(new_Jinkela_wire_17398),
        .dout(new_Jinkela_wire_17399)
    );

    bfr new_Jinkela_buffer_14449 (
        .din(new_Jinkela_wire_17263),
        .dout(new_Jinkela_wire_17264)
    );

    bfr new_Jinkela_buffer_14607 (
        .din(new_Jinkela_wire_17437),
        .dout(new_Jinkela_wire_17438)
    );

    bfr new_Jinkela_buffer_14450 (
        .din(new_Jinkela_wire_17264),
        .dout(new_Jinkela_wire_17265)
    );

    bfr new_Jinkela_buffer_14573 (
        .din(new_Jinkela_wire_17399),
        .dout(new_Jinkela_wire_17400)
    );

    bfr new_Jinkela_buffer_14451 (
        .din(new_Jinkela_wire_17265),
        .dout(new_Jinkela_wire_17266)
    );

    bfr new_Jinkela_buffer_14452 (
        .din(new_Jinkela_wire_17266),
        .dout(new_Jinkela_wire_17267)
    );

    spl2 new_Jinkela_splitter_1272 (
        .a(_0864_),
        .b(new_Jinkela_wire_17551),
        .c(new_Jinkela_wire_17552)
    );

    bfr new_Jinkela_buffer_14574 (
        .din(new_Jinkela_wire_17400),
        .dout(new_Jinkela_wire_17401)
    );

    bfr new_Jinkela_buffer_14453 (
        .din(new_Jinkela_wire_17267),
        .dout(new_Jinkela_wire_17268)
    );

    bfr new_Jinkela_buffer_14608 (
        .din(new_Jinkela_wire_17438),
        .dout(new_Jinkela_wire_17439)
    );

    bfr new_Jinkela_buffer_14454 (
        .din(new_Jinkela_wire_17268),
        .dout(new_Jinkela_wire_17269)
    );

    bfr new_Jinkela_buffer_14575 (
        .din(new_Jinkela_wire_17401),
        .dout(new_Jinkela_wire_17402)
    );

    bfr new_Jinkela_buffer_14455 (
        .din(new_Jinkela_wire_17269),
        .dout(new_Jinkela_wire_17270)
    );

    bfr new_Jinkela_buffer_14456 (
        .din(new_Jinkela_wire_17270),
        .dout(new_Jinkela_wire_17271)
    );

    bfr new_Jinkela_buffer_14704 (
        .din(_1834_),
        .dout(new_Jinkela_wire_17553)
    );

    bfr new_Jinkela_buffer_14576 (
        .din(new_Jinkela_wire_17402),
        .dout(new_Jinkela_wire_17403)
    );

    bfr new_Jinkela_buffer_14457 (
        .din(new_Jinkela_wire_17271),
        .dout(new_Jinkela_wire_17272)
    );

    bfr new_Jinkela_buffer_14609 (
        .din(new_Jinkela_wire_17439),
        .dout(new_Jinkela_wire_17440)
    );

    bfr new_Jinkela_buffer_14458 (
        .din(new_Jinkela_wire_17272),
        .dout(new_Jinkela_wire_17273)
    );

    bfr new_Jinkela_buffer_14577 (
        .din(new_Jinkela_wire_17403),
        .dout(new_Jinkela_wire_17404)
    );

    bfr new_Jinkela_buffer_14459 (
        .din(new_Jinkela_wire_17273),
        .dout(new_Jinkela_wire_17274)
    );

    bfr new_Jinkela_buffer_14705 (
        .din(_0889_),
        .dout(new_Jinkela_wire_17556)
    );

    bfr new_Jinkela_buffer_14460 (
        .din(new_Jinkela_wire_17274),
        .dout(new_Jinkela_wire_17275)
    );

    spl2 new_Jinkela_splitter_1273 (
        .a(_0645_),
        .b(new_Jinkela_wire_17554),
        .c(new_Jinkela_wire_17555)
    );

    bfr new_Jinkela_buffer_14578 (
        .din(new_Jinkela_wire_17404),
        .dout(new_Jinkela_wire_17405)
    );

    bfr new_Jinkela_buffer_14461 (
        .din(new_Jinkela_wire_17275),
        .dout(new_Jinkela_wire_17276)
    );

    bfr new_Jinkela_buffer_14610 (
        .din(new_Jinkela_wire_17440),
        .dout(new_Jinkela_wire_17441)
    );

    bfr new_Jinkela_buffer_14462 (
        .din(new_Jinkela_wire_17276),
        .dout(new_Jinkela_wire_17277)
    );

    bfr new_Jinkela_buffer_14579 (
        .din(new_Jinkela_wire_17405),
        .dout(new_Jinkela_wire_17406)
    );

    bfr new_Jinkela_buffer_14463 (
        .din(new_Jinkela_wire_17277),
        .dout(new_Jinkela_wire_17278)
    );

    bfr new_Jinkela_buffer_14464 (
        .din(new_Jinkela_wire_17278),
        .dout(new_Jinkela_wire_17279)
    );

    bfr new_Jinkela_buffer_4339 (
        .din(new_Jinkela_wire_5668),
        .dout(new_Jinkela_wire_5669)
    );

    bfr new_Jinkela_buffer_17878 (
        .din(new_Jinkela_wire_21310),
        .dout(new_Jinkela_wire_21311)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_1223),
        .dout(new_Jinkela_wire_1224)
    );

    bfr new_Jinkela_buffer_4172 (
        .din(new_Jinkela_wire_5483),
        .dout(new_Jinkela_wire_5484)
    );

    bfr new_Jinkela_buffer_4116 (
        .din(new_Jinkela_wire_5391),
        .dout(new_Jinkela_wire_5392)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_1317),
        .dout(new_Jinkela_wire_1318)
    );

    bfr new_Jinkela_buffer_17879 (
        .din(new_Jinkela_wire_21311),
        .dout(new_Jinkela_wire_21312)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_1224),
        .dout(new_Jinkela_wire_1225)
    );

    bfr new_Jinkela_buffer_4117 (
        .din(new_Jinkela_wire_5392),
        .dout(new_Jinkela_wire_5393)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_1398),
        .dout(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_4230 (
        .din(new_Jinkela_wire_5553),
        .dout(new_Jinkela_wire_5554)
    );

    bfr new_Jinkela_buffer_17880 (
        .din(new_Jinkela_wire_21312),
        .dout(new_Jinkela_wire_21313)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_1225),
        .dout(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_4173 (
        .din(new_Jinkela_wire_5484),
        .dout(new_Jinkela_wire_5485)
    );

    bfr new_Jinkela_buffer_4118 (
        .din(new_Jinkela_wire_5393),
        .dout(new_Jinkela_wire_5394)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_1318),
        .dout(new_Jinkela_wire_1319)
    );

    bfr new_Jinkela_buffer_17881 (
        .din(new_Jinkela_wire_21313),
        .dout(new_Jinkela_wire_21314)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_1226),
        .dout(new_Jinkela_wire_1227)
    );

    bfr new_Jinkela_buffer_4119 (
        .din(new_Jinkela_wire_5394),
        .dout(new_Jinkela_wire_5395)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_1350),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_17882 (
        .din(new_Jinkela_wire_21314),
        .dout(new_Jinkela_wire_21315)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_1227),
        .dout(new_Jinkela_wire_1228)
    );

    bfr new_Jinkela_buffer_4174 (
        .din(new_Jinkela_wire_5485),
        .dout(new_Jinkela_wire_5486)
    );

    bfr new_Jinkela_buffer_4120 (
        .din(new_Jinkela_wire_5395),
        .dout(new_Jinkela_wire_5396)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_1319),
        .dout(new_Jinkela_wire_1320)
    );

    bfr new_Jinkela_buffer_17883 (
        .din(new_Jinkela_wire_21315),
        .dout(new_Jinkela_wire_21316)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_1228),
        .dout(new_Jinkela_wire_1229)
    );

    spl2 new_Jinkela_splitter_515 (
        .a(_1425_),
        .b(new_Jinkela_wire_5683),
        .c(new_Jinkela_wire_5684)
    );

    bfr new_Jinkela_buffer_4121 (
        .din(new_Jinkela_wire_5396),
        .dout(new_Jinkela_wire_5397)
    );

    bfr new_Jinkela_buffer_822 (
        .din(_1196_),
        .dout(new_Jinkela_wire_1572)
    );

    bfr new_Jinkela_buffer_4231 (
        .din(new_Jinkela_wire_5554),
        .dout(new_Jinkela_wire_5555)
    );

    bfr new_Jinkela_buffer_17884 (
        .din(new_Jinkela_wire_21316),
        .dout(new_Jinkela_wire_21317)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_1229),
        .dout(new_Jinkela_wire_1230)
    );

    bfr new_Jinkela_buffer_4175 (
        .din(new_Jinkela_wire_5486),
        .dout(new_Jinkela_wire_5487)
    );

    bfr new_Jinkela_buffer_4122 (
        .din(new_Jinkela_wire_5397),
        .dout(new_Jinkela_wire_5398)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_1320),
        .dout(new_Jinkela_wire_1321)
    );

    bfr new_Jinkela_buffer_17885 (
        .din(new_Jinkela_wire_21317),
        .dout(new_Jinkela_wire_21318)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_1230),
        .dout(new_Jinkela_wire_1231)
    );

    bfr new_Jinkela_buffer_4123 (
        .din(new_Jinkela_wire_5398),
        .dout(new_Jinkela_wire_5399)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_1351),
        .dout(new_Jinkela_wire_1352)
    );

    bfr new_Jinkela_buffer_17886 (
        .din(new_Jinkela_wire_21318),
        .dout(new_Jinkela_wire_21319)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_1231),
        .dout(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_4176 (
        .din(new_Jinkela_wire_5487),
        .dout(new_Jinkela_wire_5488)
    );

    bfr new_Jinkela_buffer_4124 (
        .din(new_Jinkela_wire_5399),
        .dout(new_Jinkela_wire_5400)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_1321),
        .dout(new_Jinkela_wire_1322)
    );

    bfr new_Jinkela_buffer_17887 (
        .din(new_Jinkela_wire_21319),
        .dout(new_Jinkela_wire_21320)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_1232),
        .dout(new_Jinkela_wire_1233)
    );

    bfr new_Jinkela_buffer_4125 (
        .din(new_Jinkela_wire_5400),
        .dout(new_Jinkela_wire_5401)
    );

    spl2 new_Jinkela_splitter_222 (
        .a(new_Jinkela_wire_1567),
        .b(new_Jinkela_wire_1568),
        .c(new_Jinkela_wire_1569)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_1399),
        .dout(new_Jinkela_wire_1400)
    );

    bfr new_Jinkela_buffer_4232 (
        .din(new_Jinkela_wire_5555),
        .dout(new_Jinkela_wire_5556)
    );

    bfr new_Jinkela_buffer_17888 (
        .din(new_Jinkela_wire_21320),
        .dout(new_Jinkela_wire_21321)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_1233),
        .dout(new_Jinkela_wire_1234)
    );

    bfr new_Jinkela_buffer_4177 (
        .din(new_Jinkela_wire_5488),
        .dout(new_Jinkela_wire_5489)
    );

    bfr new_Jinkela_buffer_4126 (
        .din(new_Jinkela_wire_5401),
        .dout(new_Jinkela_wire_5402)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_17889 (
        .din(new_Jinkela_wire_21321),
        .dout(new_Jinkela_wire_21322)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_1234),
        .dout(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_4127 (
        .din(new_Jinkela_wire_5402),
        .dout(new_Jinkela_wire_5403)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_1352),
        .dout(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_4340 (
        .din(new_Jinkela_wire_5669),
        .dout(new_Jinkela_wire_5670)
    );

    bfr new_Jinkela_buffer_17890 (
        .din(new_Jinkela_wire_21322),
        .dout(new_Jinkela_wire_21323)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_1235),
        .dout(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_4178 (
        .din(new_Jinkela_wire_5489),
        .dout(new_Jinkela_wire_5490)
    );

    bfr new_Jinkela_buffer_4128 (
        .din(new_Jinkela_wire_5403),
        .dout(new_Jinkela_wire_5404)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_1323),
        .dout(new_Jinkela_wire_1324)
    );

    spl2 new_Jinkela_splitter_1565 (
        .a(new_Jinkela_wire_21323),
        .b(new_Jinkela_wire_21324),
        .c(new_Jinkela_wire_21325)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_1236),
        .dout(new_Jinkela_wire_1237)
    );

    bfr new_Jinkela_buffer_4129 (
        .din(new_Jinkela_wire_5404),
        .dout(new_Jinkela_wire_5405)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_1405),
        .dout(new_Jinkela_wire_1406)
    );

    bfr new_Jinkela_buffer_4233 (
        .din(new_Jinkela_wire_5556),
        .dout(new_Jinkela_wire_5557)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_1237),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_4179 (
        .din(new_Jinkela_wire_5490),
        .dout(new_Jinkela_wire_5491)
    );

    bfr new_Jinkela_buffer_4130 (
        .din(new_Jinkela_wire_5405),
        .dout(new_Jinkela_wire_5406)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_1324),
        .dout(new_Jinkela_wire_1325)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_1238),
        .dout(new_Jinkela_wire_1239)
    );

    bfr new_Jinkela_buffer_4131 (
        .din(new_Jinkela_wire_5406),
        .dout(new_Jinkela_wire_5407)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_1353),
        .dout(new_Jinkela_wire_1354)
    );

    spl2 new_Jinkela_splitter_517 (
        .a(_1525_),
        .b(new_Jinkela_wire_5687),
        .c(new_Jinkela_wire_5688)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_1239),
        .dout(new_Jinkela_wire_1240)
    );

    bfr new_Jinkela_buffer_4180 (
        .din(new_Jinkela_wire_5491),
        .dout(new_Jinkela_wire_5492)
    );

    bfr new_Jinkela_buffer_4132 (
        .din(new_Jinkela_wire_5407),
        .dout(new_Jinkela_wire_5408)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_1325),
        .dout(new_Jinkela_wire_1326)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_1240),
        .dout(new_Jinkela_wire_1241)
    );

    spl2 new_Jinkela_splitter_516 (
        .a(_0969_),
        .b(new_Jinkela_wire_5685),
        .c(new_Jinkela_wire_5686)
    );

    bfr new_Jinkela_buffer_4133 (
        .din(new_Jinkela_wire_5408),
        .dout(new_Jinkela_wire_5409)
    );

    bfr new_Jinkela_buffer_4234 (
        .din(new_Jinkela_wire_5557),
        .dout(new_Jinkela_wire_5558)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_1241),
        .dout(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_4181 (
        .din(new_Jinkela_wire_5492),
        .dout(new_Jinkela_wire_5493)
    );

    bfr new_Jinkela_buffer_4134 (
        .din(new_Jinkela_wire_5409),
        .dout(new_Jinkela_wire_5410)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_1326),
        .dout(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_1242),
        .dout(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_4135 (
        .din(new_Jinkela_wire_5410),
        .dout(new_Jinkela_wire_5411)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_1354),
        .dout(new_Jinkela_wire_1355)
    );

    bfr new_Jinkela_buffer_4341 (
        .din(new_Jinkela_wire_5670),
        .dout(new_Jinkela_wire_5671)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_1243),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_4182 (
        .din(new_Jinkela_wire_5493),
        .dout(new_Jinkela_wire_5494)
    );

    bfr new_Jinkela_buffer_4136 (
        .din(new_Jinkela_wire_5411),
        .dout(new_Jinkela_wire_5412)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_1327),
        .dout(new_Jinkela_wire_1328)
    );

    bfr new_Jinkela_buffer_7634 (
        .din(new_Jinkela_wire_9461),
        .dout(new_Jinkela_wire_9462)
    );

    bfr new_Jinkela_buffer_11115 (
        .din(new_Jinkela_wire_13412),
        .dout(new_Jinkela_wire_13413)
    );

    bfr new_Jinkela_buffer_7571 (
        .din(new_Jinkela_wire_9394),
        .dout(new_Jinkela_wire_9395)
    );

    bfr new_Jinkela_buffer_11042 (
        .din(new_Jinkela_wire_13297),
        .dout(new_Jinkela_wire_13298)
    );

    spl2 new_Jinkela_splitter_768 (
        .a(_1112_),
        .b(new_Jinkela_wire_9550),
        .c(new_Jinkela_wire_9551)
    );

    bfr new_Jinkela_buffer_7708 (
        .din(new_Jinkela_wire_9545),
        .dout(new_Jinkela_wire_9546)
    );

    bfr new_Jinkela_buffer_11096 (
        .din(new_Jinkela_wire_13373),
        .dout(new_Jinkela_wire_13374)
    );

    bfr new_Jinkela_buffer_7572 (
        .din(new_Jinkela_wire_9395),
        .dout(new_Jinkela_wire_9396)
    );

    bfr new_Jinkela_buffer_11043 (
        .din(new_Jinkela_wire_13298),
        .dout(new_Jinkela_wire_13299)
    );

    bfr new_Jinkela_buffer_7635 (
        .din(new_Jinkela_wire_9462),
        .dout(new_Jinkela_wire_9463)
    );

    spl2 new_Jinkela_splitter_998 (
        .a(_0061_),
        .b(new_Jinkela_wire_13457),
        .c(new_Jinkela_wire_13458)
    );

    bfr new_Jinkela_buffer_7573 (
        .din(new_Jinkela_wire_9396),
        .dout(new_Jinkela_wire_9397)
    );

    bfr new_Jinkela_buffer_11044 (
        .din(new_Jinkela_wire_13299),
        .dout(new_Jinkela_wire_13300)
    );

    spl2 new_Jinkela_splitter_763 (
        .a(new_Jinkela_wire_9517),
        .b(new_Jinkela_wire_9518),
        .c(new_Jinkela_wire_9519)
    );

    spl2 new_Jinkela_splitter_999 (
        .a(_0446_),
        .b(new_Jinkela_wire_13459),
        .c(new_Jinkela_wire_13460)
    );

    bfr new_Jinkela_buffer_11097 (
        .din(new_Jinkela_wire_13374),
        .dout(new_Jinkela_wire_13375)
    );

    bfr new_Jinkela_buffer_7574 (
        .din(new_Jinkela_wire_9397),
        .dout(new_Jinkela_wire_9398)
    );

    bfr new_Jinkela_buffer_11045 (
        .din(new_Jinkela_wire_13300),
        .dout(new_Jinkela_wire_13301)
    );

    bfr new_Jinkela_buffer_7636 (
        .din(new_Jinkela_wire_9463),
        .dout(new_Jinkela_wire_9464)
    );

    bfr new_Jinkela_buffer_11116 (
        .din(new_Jinkela_wire_13413),
        .dout(new_Jinkela_wire_13414)
    );

    bfr new_Jinkela_buffer_7575 (
        .din(new_Jinkela_wire_9398),
        .dout(new_Jinkela_wire_9399)
    );

    bfr new_Jinkela_buffer_11046 (
        .din(new_Jinkela_wire_13301),
        .dout(new_Jinkela_wire_13302)
    );

    bfr new_Jinkela_buffer_11098 (
        .din(new_Jinkela_wire_13375),
        .dout(new_Jinkela_wire_13376)
    );

    bfr new_Jinkela_buffer_7576 (
        .din(new_Jinkela_wire_9399),
        .dout(new_Jinkela_wire_9400)
    );

    bfr new_Jinkela_buffer_11047 (
        .din(new_Jinkela_wire_13302),
        .dout(new_Jinkela_wire_13303)
    );

    bfr new_Jinkela_buffer_7637 (
        .din(new_Jinkela_wire_9464),
        .dout(new_Jinkela_wire_9465)
    );

    spl2 new_Jinkela_splitter_1004 (
        .a(_1178_),
        .b(new_Jinkela_wire_13574),
        .c(new_Jinkela_wire_13575)
    );

    bfr new_Jinkela_buffer_7577 (
        .din(new_Jinkela_wire_9400),
        .dout(new_Jinkela_wire_9401)
    );

    spl2 new_Jinkela_splitter_977 (
        .a(new_Jinkela_wire_13303),
        .b(new_Jinkela_wire_13304),
        .c(new_Jinkela_wire_13305)
    );

    bfr new_Jinkela_buffer_7694 (
        .din(new_Jinkela_wire_9525),
        .dout(new_Jinkela_wire_9526)
    );

    bfr new_Jinkela_buffer_11117 (
        .din(new_Jinkela_wire_13414),
        .dout(new_Jinkela_wire_13415)
    );

    bfr new_Jinkela_buffer_7578 (
        .din(new_Jinkela_wire_9401),
        .dout(new_Jinkela_wire_9402)
    );

    bfr new_Jinkela_buffer_11099 (
        .din(new_Jinkela_wire_13376),
        .dout(new_Jinkela_wire_13377)
    );

    bfr new_Jinkela_buffer_7638 (
        .din(new_Jinkela_wire_9465),
        .dout(new_Jinkela_wire_9466)
    );

    bfr new_Jinkela_buffer_11100 (
        .din(new_Jinkela_wire_13377),
        .dout(new_Jinkela_wire_13378)
    );

    bfr new_Jinkela_buffer_7579 (
        .din(new_Jinkela_wire_9402),
        .dout(new_Jinkela_wire_9403)
    );

    bfr new_Jinkela_buffer_7695 (
        .din(new_Jinkela_wire_9526),
        .dout(new_Jinkela_wire_9527)
    );

    bfr new_Jinkela_buffer_11101 (
        .din(new_Jinkela_wire_13378),
        .dout(new_Jinkela_wire_13379)
    );

    bfr new_Jinkela_buffer_7580 (
        .din(new_Jinkela_wire_9403),
        .dout(new_Jinkela_wire_9404)
    );

    bfr new_Jinkela_buffer_11118 (
        .din(new_Jinkela_wire_13415),
        .dout(new_Jinkela_wire_13416)
    );

    bfr new_Jinkela_buffer_7639 (
        .din(new_Jinkela_wire_9466),
        .dout(new_Jinkela_wire_9467)
    );

    bfr new_Jinkela_buffer_11102 (
        .din(new_Jinkela_wire_13379),
        .dout(new_Jinkela_wire_13380)
    );

    bfr new_Jinkela_buffer_7581 (
        .din(new_Jinkela_wire_9404),
        .dout(new_Jinkela_wire_9405)
    );

    bfr new_Jinkela_buffer_11159 (
        .din(_0643_),
        .dout(new_Jinkela_wire_13461)
    );

    spl2 new_Jinkela_splitter_1001 (
        .a(_0268_),
        .b(new_Jinkela_wire_13464),
        .c(new_Jinkela_wire_13465)
    );

    spl2 new_Jinkela_splitter_769 (
        .a(_1304_),
        .b(new_Jinkela_wire_9556),
        .c(new_Jinkela_wire_9557)
    );

    bfr new_Jinkela_buffer_11119 (
        .din(new_Jinkela_wire_13416),
        .dout(new_Jinkela_wire_13417)
    );

    bfr new_Jinkela_buffer_7582 (
        .din(new_Jinkela_wire_9405),
        .dout(new_Jinkela_wire_9406)
    );

    spl2 new_Jinkela_splitter_1000 (
        .a(_0394_),
        .b(new_Jinkela_wire_13462),
        .c(new_Jinkela_wire_13463)
    );

    bfr new_Jinkela_buffer_7640 (
        .din(new_Jinkela_wire_9467),
        .dout(new_Jinkela_wire_9468)
    );

    bfr new_Jinkela_buffer_11120 (
        .din(new_Jinkela_wire_13417),
        .dout(new_Jinkela_wire_13418)
    );

    bfr new_Jinkela_buffer_7583 (
        .din(new_Jinkela_wire_9406),
        .dout(new_Jinkela_wire_9407)
    );

    bfr new_Jinkela_buffer_7696 (
        .din(new_Jinkela_wire_9527),
        .dout(new_Jinkela_wire_9528)
    );

    bfr new_Jinkela_buffer_11121 (
        .din(new_Jinkela_wire_13418),
        .dout(new_Jinkela_wire_13419)
    );

    bfr new_Jinkela_buffer_7584 (
        .din(new_Jinkela_wire_9407),
        .dout(new_Jinkela_wire_9408)
    );

    bfr new_Jinkela_buffer_11160 (
        .din(_0531_),
        .dout(new_Jinkela_wire_13466)
    );

    bfr new_Jinkela_buffer_7641 (
        .din(new_Jinkela_wire_9468),
        .dout(new_Jinkela_wire_9469)
    );

    bfr new_Jinkela_buffer_11122 (
        .din(new_Jinkela_wire_13419),
        .dout(new_Jinkela_wire_13420)
    );

    bfr new_Jinkela_buffer_7585 (
        .din(new_Jinkela_wire_9408),
        .dout(new_Jinkela_wire_9409)
    );

    spl2 new_Jinkela_splitter_1003 (
        .a(_0343_),
        .b(new_Jinkela_wire_13572),
        .c(new_Jinkela_wire_13573)
    );

    bfr new_Jinkela_buffer_11161 (
        .din(new_Jinkela_wire_13466),
        .dout(new_Jinkela_wire_13467)
    );

    bfr new_Jinkela_buffer_7712 (
        .din(new_Jinkela_wire_9551),
        .dout(new_Jinkela_wire_9552)
    );

    bfr new_Jinkela_buffer_11123 (
        .din(new_Jinkela_wire_13420),
        .dout(new_Jinkela_wire_13421)
    );

    bfr new_Jinkela_buffer_7586 (
        .din(new_Jinkela_wire_9409),
        .dout(new_Jinkela_wire_9410)
    );

    bfr new_Jinkela_buffer_7642 (
        .din(new_Jinkela_wire_9469),
        .dout(new_Jinkela_wire_9470)
    );

    bfr new_Jinkela_buffer_11124 (
        .din(new_Jinkela_wire_13421),
        .dout(new_Jinkela_wire_13422)
    );

    bfr new_Jinkela_buffer_7587 (
        .din(new_Jinkela_wire_9410),
        .dout(new_Jinkela_wire_9411)
    );

    bfr new_Jinkela_buffer_7697 (
        .din(new_Jinkela_wire_9528),
        .dout(new_Jinkela_wire_9529)
    );

    bfr new_Jinkela_buffer_11162 (
        .din(new_Jinkela_wire_13467),
        .dout(new_Jinkela_wire_13468)
    );

    bfr new_Jinkela_buffer_11125 (
        .din(new_Jinkela_wire_13422),
        .dout(new_Jinkela_wire_13423)
    );

    bfr new_Jinkela_buffer_7588 (
        .din(new_Jinkela_wire_9411),
        .dout(new_Jinkela_wire_9412)
    );

    bfr new_Jinkela_buffer_7643 (
        .din(new_Jinkela_wire_9470),
        .dout(new_Jinkela_wire_9471)
    );

    bfr new_Jinkela_buffer_11126 (
        .din(new_Jinkela_wire_13423),
        .dout(new_Jinkela_wire_13424)
    );

    bfr new_Jinkela_buffer_7589 (
        .din(new_Jinkela_wire_9412),
        .dout(new_Jinkela_wire_9413)
    );

    spl2 new_Jinkela_splitter_1005 (
        .a(_0238_),
        .b(new_Jinkela_wire_13580),
        .c(new_Jinkela_wire_13581)
    );

    bfr new_Jinkela_buffer_7709 (
        .din(new_Jinkela_wire_9546),
        .dout(new_Jinkela_wire_9547)
    );

    bfr new_Jinkela_buffer_11163 (
        .din(new_Jinkela_wire_13468),
        .dout(new_Jinkela_wire_13469)
    );

    bfr new_Jinkela_buffer_11127 (
        .din(new_Jinkela_wire_13424),
        .dout(new_Jinkela_wire_13425)
    );

    bfr new_Jinkela_buffer_7590 (
        .din(new_Jinkela_wire_9413),
        .dout(new_Jinkela_wire_9414)
    );

    bfr new_Jinkela_buffer_7644 (
        .din(new_Jinkela_wire_9471),
        .dout(new_Jinkela_wire_9472)
    );

    bfr new_Jinkela_buffer_11264 (
        .din(new_Jinkela_wire_13575),
        .dout(new_Jinkela_wire_13576)
    );

    bfr new_Jinkela_buffer_11128 (
        .din(new_Jinkela_wire_13425),
        .dout(new_Jinkela_wire_13426)
    );

    bfr new_Jinkela_buffer_7591 (
        .din(new_Jinkela_wire_9414),
        .dout(new_Jinkela_wire_9415)
    );

    spl2 new_Jinkela_splitter_1006 (
        .a(_0408_),
        .b(new_Jinkela_wire_13582),
        .c(new_Jinkela_wire_13583)
    );

    bfr new_Jinkela_buffer_14783 (
        .din(_1704_),
        .dout(new_Jinkela_wire_17638)
    );

    bfr new_Jinkela_buffer_14580 (
        .din(new_Jinkela_wire_17406),
        .dout(new_Jinkela_wire_17407)
    );

    bfr new_Jinkela_buffer_14465 (
        .din(new_Jinkela_wire_17279),
        .dout(new_Jinkela_wire_17280)
    );

    bfr new_Jinkela_buffer_14611 (
        .din(new_Jinkela_wire_17441),
        .dout(new_Jinkela_wire_17442)
    );

    bfr new_Jinkela_buffer_14466 (
        .din(new_Jinkela_wire_17280),
        .dout(new_Jinkela_wire_17281)
    );

    bfr new_Jinkela_buffer_14581 (
        .din(new_Jinkela_wire_17407),
        .dout(new_Jinkela_wire_17408)
    );

    bfr new_Jinkela_buffer_14467 (
        .din(new_Jinkela_wire_17281),
        .dout(new_Jinkela_wire_17282)
    );

    spl2 new_Jinkela_splitter_1275 (
        .a(_0539_),
        .b(new_Jinkela_wire_17636),
        .c(new_Jinkela_wire_17637)
    );

    bfr new_Jinkela_buffer_14468 (
        .din(new_Jinkela_wire_17282),
        .dout(new_Jinkela_wire_17283)
    );

    bfr new_Jinkela_buffer_14582 (
        .din(new_Jinkela_wire_17408),
        .dout(new_Jinkela_wire_17409)
    );

    bfr new_Jinkela_buffer_14469 (
        .din(new_Jinkela_wire_17283),
        .dout(new_Jinkela_wire_17284)
    );

    bfr new_Jinkela_buffer_14612 (
        .din(new_Jinkela_wire_17442),
        .dout(new_Jinkela_wire_17443)
    );

    bfr new_Jinkela_buffer_14470 (
        .din(new_Jinkela_wire_17284),
        .dout(new_Jinkela_wire_17285)
    );

    bfr new_Jinkela_buffer_14583 (
        .din(new_Jinkela_wire_17409),
        .dout(new_Jinkela_wire_17410)
    );

    bfr new_Jinkela_buffer_14471 (
        .din(new_Jinkela_wire_17285),
        .dout(new_Jinkela_wire_17286)
    );

    bfr new_Jinkela_buffer_14706 (
        .din(new_Jinkela_wire_17556),
        .dout(new_Jinkela_wire_17557)
    );

    bfr new_Jinkela_buffer_14472 (
        .din(new_Jinkela_wire_17286),
        .dout(new_Jinkela_wire_17287)
    );

    bfr new_Jinkela_buffer_14584 (
        .din(new_Jinkela_wire_17410),
        .dout(new_Jinkela_wire_17411)
    );

    bfr new_Jinkela_buffer_14473 (
        .din(new_Jinkela_wire_17287),
        .dout(new_Jinkela_wire_17288)
    );

    bfr new_Jinkela_buffer_14613 (
        .din(new_Jinkela_wire_17443),
        .dout(new_Jinkela_wire_17444)
    );

    bfr new_Jinkela_buffer_14474 (
        .din(new_Jinkela_wire_17288),
        .dout(new_Jinkela_wire_17289)
    );

    bfr new_Jinkela_buffer_14585 (
        .din(new_Jinkela_wire_17411),
        .dout(new_Jinkela_wire_17412)
    );

    bfr new_Jinkela_buffer_14475 (
        .din(new_Jinkela_wire_17289),
        .dout(new_Jinkela_wire_17290)
    );

    spl2 new_Jinkela_splitter_1278 (
        .a(_1404_),
        .b(new_Jinkela_wire_17658),
        .c(new_Jinkela_wire_17659)
    );

    bfr new_Jinkela_buffer_14476 (
        .din(new_Jinkela_wire_17290),
        .dout(new_Jinkela_wire_17291)
    );

    bfr new_Jinkela_buffer_14586 (
        .din(new_Jinkela_wire_17412),
        .dout(new_Jinkela_wire_17413)
    );

    bfr new_Jinkela_buffer_14477 (
        .din(new_Jinkela_wire_17291),
        .dout(new_Jinkela_wire_17292)
    );

    bfr new_Jinkela_buffer_14614 (
        .din(new_Jinkela_wire_17444),
        .dout(new_Jinkela_wire_17445)
    );

    bfr new_Jinkela_buffer_14478 (
        .din(new_Jinkela_wire_17292),
        .dout(new_Jinkela_wire_17293)
    );

    bfr new_Jinkela_buffer_14587 (
        .din(new_Jinkela_wire_17413),
        .dout(new_Jinkela_wire_17414)
    );

    bfr new_Jinkela_buffer_14479 (
        .din(new_Jinkela_wire_17293),
        .dout(new_Jinkela_wire_17294)
    );

    bfr new_Jinkela_buffer_14707 (
        .din(new_Jinkela_wire_17557),
        .dout(new_Jinkela_wire_17558)
    );

    bfr new_Jinkela_buffer_14480 (
        .din(new_Jinkela_wire_17294),
        .dout(new_Jinkela_wire_17295)
    );

    bfr new_Jinkela_buffer_14588 (
        .din(new_Jinkela_wire_17414),
        .dout(new_Jinkela_wire_17415)
    );

    bfr new_Jinkela_buffer_14481 (
        .din(new_Jinkela_wire_17295),
        .dout(new_Jinkela_wire_17296)
    );

    bfr new_Jinkela_buffer_14615 (
        .din(new_Jinkela_wire_17445),
        .dout(new_Jinkela_wire_17446)
    );

    bfr new_Jinkela_buffer_14482 (
        .din(new_Jinkela_wire_17296),
        .dout(new_Jinkela_wire_17297)
    );

    bfr new_Jinkela_buffer_14589 (
        .din(new_Jinkela_wire_17415),
        .dout(new_Jinkela_wire_17416)
    );

    bfr new_Jinkela_buffer_14483 (
        .din(new_Jinkela_wire_17297),
        .dout(new_Jinkela_wire_17298)
    );

    bfr new_Jinkela_buffer_14484 (
        .din(new_Jinkela_wire_17298),
        .dout(new_Jinkela_wire_17299)
    );

    spl2 new_Jinkela_splitter_1277 (
        .a(_0189_),
        .b(new_Jinkela_wire_17656),
        .c(new_Jinkela_wire_17657)
    );

    bfr new_Jinkela_buffer_14590 (
        .din(new_Jinkela_wire_17416),
        .dout(new_Jinkela_wire_17417)
    );

    bfr new_Jinkela_buffer_14485 (
        .din(new_Jinkela_wire_17299),
        .dout(new_Jinkela_wire_17300)
    );

    bfr new_Jinkela_buffer_7698 (
        .din(new_Jinkela_wire_9529),
        .dout(new_Jinkela_wire_9530)
    );

    bfr new_Jinkela_buffer_7592 (
        .din(new_Jinkela_wire_9415),
        .dout(new_Jinkela_wire_9416)
    );

    bfr new_Jinkela_buffer_7645 (
        .din(new_Jinkela_wire_9472),
        .dout(new_Jinkela_wire_9473)
    );

    bfr new_Jinkela_buffer_7593 (
        .din(new_Jinkela_wire_9416),
        .dout(new_Jinkela_wire_9417)
    );

    spl2 new_Jinkela_splitter_770 (
        .a(_0501_),
        .b(new_Jinkela_wire_9558),
        .c(new_Jinkela_wire_9559)
    );

    bfr new_Jinkela_buffer_7594 (
        .din(new_Jinkela_wire_9417),
        .dout(new_Jinkela_wire_9418)
    );

    bfr new_Jinkela_buffer_7646 (
        .din(new_Jinkela_wire_9473),
        .dout(new_Jinkela_wire_9474)
    );

    bfr new_Jinkela_buffer_7595 (
        .din(new_Jinkela_wire_9418),
        .dout(new_Jinkela_wire_9419)
    );

    bfr new_Jinkela_buffer_7699 (
        .din(new_Jinkela_wire_9530),
        .dout(new_Jinkela_wire_9531)
    );

    bfr new_Jinkela_buffer_7596 (
        .din(new_Jinkela_wire_9419),
        .dout(new_Jinkela_wire_9420)
    );

    bfr new_Jinkela_buffer_7647 (
        .din(new_Jinkela_wire_9474),
        .dout(new_Jinkela_wire_9475)
    );

    bfr new_Jinkela_buffer_7597 (
        .din(new_Jinkela_wire_9420),
        .dout(new_Jinkela_wire_9421)
    );

    bfr new_Jinkela_buffer_7710 (
        .din(new_Jinkela_wire_9547),
        .dout(new_Jinkela_wire_9548)
    );

    bfr new_Jinkela_buffer_7598 (
        .din(new_Jinkela_wire_9421),
        .dout(new_Jinkela_wire_9422)
    );

    bfr new_Jinkela_buffer_7648 (
        .din(new_Jinkela_wire_9475),
        .dout(new_Jinkela_wire_9476)
    );

    bfr new_Jinkela_buffer_7599 (
        .din(new_Jinkela_wire_9422),
        .dout(new_Jinkela_wire_9423)
    );

    bfr new_Jinkela_buffer_7700 (
        .din(new_Jinkela_wire_9531),
        .dout(new_Jinkela_wire_9532)
    );

    bfr new_Jinkela_buffer_7600 (
        .din(new_Jinkela_wire_9423),
        .dout(new_Jinkela_wire_9424)
    );

    bfr new_Jinkela_buffer_7649 (
        .din(new_Jinkela_wire_9476),
        .dout(new_Jinkela_wire_9477)
    );

    bfr new_Jinkela_buffer_7601 (
        .din(new_Jinkela_wire_9424),
        .dout(new_Jinkela_wire_9425)
    );

    bfr new_Jinkela_buffer_7720 (
        .din(_0164_),
        .dout(new_Jinkela_wire_9564)
    );

    bfr new_Jinkela_buffer_7602 (
        .din(new_Jinkela_wire_9425),
        .dout(new_Jinkela_wire_9426)
    );

    bfr new_Jinkela_buffer_7650 (
        .din(new_Jinkela_wire_9477),
        .dout(new_Jinkela_wire_9478)
    );

    bfr new_Jinkela_buffer_7603 (
        .din(new_Jinkela_wire_9426),
        .dout(new_Jinkela_wire_9427)
    );

    bfr new_Jinkela_buffer_7701 (
        .din(new_Jinkela_wire_9532),
        .dout(new_Jinkela_wire_9533)
    );

    bfr new_Jinkela_buffer_7604 (
        .din(new_Jinkela_wire_9427),
        .dout(new_Jinkela_wire_9428)
    );

    bfr new_Jinkela_buffer_7651 (
        .din(new_Jinkela_wire_9478),
        .dout(new_Jinkela_wire_9479)
    );

    bfr new_Jinkela_buffer_7605 (
        .din(new_Jinkela_wire_9428),
        .dout(new_Jinkela_wire_9429)
    );

    bfr new_Jinkela_buffer_7711 (
        .din(new_Jinkela_wire_9548),
        .dout(new_Jinkela_wire_9549)
    );

    bfr new_Jinkela_buffer_7606 (
        .din(new_Jinkela_wire_9429),
        .dout(new_Jinkela_wire_9430)
    );

    bfr new_Jinkela_buffer_7652 (
        .din(new_Jinkela_wire_9479),
        .dout(new_Jinkela_wire_9480)
    );

    bfr new_Jinkela_buffer_7607 (
        .din(new_Jinkela_wire_9430),
        .dout(new_Jinkela_wire_9431)
    );

    bfr new_Jinkela_buffer_7702 (
        .din(new_Jinkela_wire_9533),
        .dout(new_Jinkela_wire_9534)
    );

    bfr new_Jinkela_buffer_7608 (
        .din(new_Jinkela_wire_9431),
        .dout(new_Jinkela_wire_9432)
    );

    bfr new_Jinkela_buffer_7653 (
        .din(new_Jinkela_wire_9480),
        .dout(new_Jinkela_wire_9481)
    );

    bfr new_Jinkela_buffer_7609 (
        .din(new_Jinkela_wire_9432),
        .dout(new_Jinkela_wire_9433)
    );

    bfr new_Jinkela_buffer_7713 (
        .din(new_Jinkela_wire_9552),
        .dout(new_Jinkela_wire_9553)
    );

    bfr new_Jinkela_buffer_7610 (
        .din(new_Jinkela_wire_9433),
        .dout(new_Jinkela_wire_9434)
    );

    bfr new_Jinkela_buffer_7654 (
        .din(new_Jinkela_wire_9481),
        .dout(new_Jinkela_wire_9482)
    );

    bfr new_Jinkela_buffer_7611 (
        .din(new_Jinkela_wire_9434),
        .dout(new_Jinkela_wire_9435)
    );

    bfr new_Jinkela_buffer_7703 (
        .din(new_Jinkela_wire_9534),
        .dout(new_Jinkela_wire_9535)
    );

    bfr new_Jinkela_buffer_7612 (
        .din(new_Jinkela_wire_9435),
        .dout(new_Jinkela_wire_9436)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    bfr new_Jinkela_buffer_4137 (
        .din(new_Jinkela_wire_5412),
        .dout(new_Jinkela_wire_5413)
    );

    bfr new_Jinkela_buffer_4235 (
        .din(new_Jinkela_wire_5558),
        .dout(new_Jinkela_wire_5559)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_1406),
        .dout(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_4183 (
        .din(new_Jinkela_wire_5494),
        .dout(new_Jinkela_wire_5495)
    );

    bfr new_Jinkela_buffer_4138 (
        .din(new_Jinkela_wire_5413),
        .dout(new_Jinkela_wire_5414)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_1328),
        .dout(new_Jinkela_wire_1329)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_1246),
        .dout(new_Jinkela_wire_1247)
    );

    bfr new_Jinkela_buffer_4139 (
        .din(new_Jinkela_wire_5414),
        .dout(new_Jinkela_wire_5415)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_1355),
        .dout(new_Jinkela_wire_1356)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_1247),
        .dout(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_4184 (
        .din(new_Jinkela_wire_5495),
        .dout(new_Jinkela_wire_5496)
    );

    spl2 new_Jinkela_splitter_487 (
        .a(new_Jinkela_wire_5415),
        .b(new_Jinkela_wire_5416),
        .c(new_Jinkela_wire_5417)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_1329),
        .dout(new_Jinkela_wire_1330)
    );

    bfr new_Jinkela_buffer_4236 (
        .din(new_Jinkela_wire_5559),
        .dout(new_Jinkela_wire_5560)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_1248),
        .dout(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_4185 (
        .din(new_Jinkela_wire_5496),
        .dout(new_Jinkela_wire_5497)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(_1622_),
        .b(new_Jinkela_wire_1573),
        .c(new_Jinkela_wire_1574)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    bfr new_Jinkela_buffer_4342 (
        .din(new_Jinkela_wire_5671),
        .dout(new_Jinkela_wire_5672)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_1330),
        .dout(new_Jinkela_wire_1331)
    );

    bfr new_Jinkela_buffer_4186 (
        .din(new_Jinkela_wire_5497),
        .dout(new_Jinkela_wire_5498)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_1250),
        .dout(new_Jinkela_wire_1251)
    );

    bfr new_Jinkela_buffer_4237 (
        .din(new_Jinkela_wire_5560),
        .dout(new_Jinkela_wire_5561)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_1356),
        .dout(new_Jinkela_wire_1357)
    );

    bfr new_Jinkela_buffer_4187 (
        .din(new_Jinkela_wire_5498),
        .dout(new_Jinkela_wire_5499)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(new_Jinkela_wire_1251),
        .b(new_Jinkela_wire_1252),
        .c(new_Jinkela_wire_1253)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_1357),
        .dout(new_Jinkela_wire_1358)
    );

    bfr new_Jinkela_buffer_4188 (
        .din(new_Jinkela_wire_5499),
        .dout(new_Jinkela_wire_5500)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(new_Jinkela_wire_1331),
        .b(new_Jinkela_wire_1332),
        .c(new_Jinkela_wire_1333)
    );

    spl2 new_Jinkela_splitter_518 (
        .a(_0887_),
        .b(new_Jinkela_wire_5689),
        .c(new_Jinkela_wire_5690)
    );

    bfr new_Jinkela_buffer_4238 (
        .din(new_Jinkela_wire_5561),
        .dout(new_Jinkela_wire_5562)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(_0834_),
        .b(new_Jinkela_wire_1575),
        .c(new_Jinkela_wire_1576)
    );

    bfr new_Jinkela_buffer_4189 (
        .din(new_Jinkela_wire_5500),
        .dout(new_Jinkela_wire_5501)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_1407),
        .dout(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_4343 (
        .din(new_Jinkela_wire_5672),
        .dout(new_Jinkela_wire_5673)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_1358),
        .dout(new_Jinkela_wire_1359)
    );

    bfr new_Jinkela_buffer_4190 (
        .din(new_Jinkela_wire_5501),
        .dout(new_Jinkela_wire_5502)
    );

    bfr new_Jinkela_buffer_4239 (
        .din(new_Jinkela_wire_5562),
        .dout(new_Jinkela_wire_5563)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_1359),
        .dout(new_Jinkela_wire_1360)
    );

    bfr new_Jinkela_buffer_4191 (
        .din(new_Jinkela_wire_5502),
        .dout(new_Jinkela_wire_5503)
    );

    bfr new_Jinkela_buffer_4359 (
        .din(_0290_),
        .dout(new_Jinkela_wire_5703)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_1360),
        .dout(new_Jinkela_wire_1361)
    );

    bfr new_Jinkela_buffer_4192 (
        .din(new_Jinkela_wire_5503),
        .dout(new_Jinkela_wire_5504)
    );

    bfr new_Jinkela_buffer_4351 (
        .din(_0787_),
        .dout(new_Jinkela_wire_5691)
    );

    bfr new_Jinkela_buffer_4240 (
        .din(new_Jinkela_wire_5563),
        .dout(new_Jinkela_wire_5564)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_1361),
        .dout(new_Jinkela_wire_1362)
    );

    bfr new_Jinkela_buffer_4193 (
        .din(new_Jinkela_wire_5504),
        .dout(new_Jinkela_wire_5505)
    );

    bfr new_Jinkela_buffer_4344 (
        .din(new_Jinkela_wire_5673),
        .dout(new_Jinkela_wire_5674)
    );

    spl2 new_Jinkela_splitter_226 (
        .a(_1509_),
        .b(new_Jinkela_wire_1577),
        .c(new_Jinkela_wire_1578)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_1362),
        .dout(new_Jinkela_wire_1363)
    );

    bfr new_Jinkela_buffer_4194 (
        .din(new_Jinkela_wire_5505),
        .dout(new_Jinkela_wire_5506)
    );

    bfr new_Jinkela_buffer_4241 (
        .din(new_Jinkela_wire_5564),
        .dout(new_Jinkela_wire_5565)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_1410),
        .dout(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_1363),
        .dout(new_Jinkela_wire_1364)
    );

    bfr new_Jinkela_buffer_4195 (
        .din(new_Jinkela_wire_5506),
        .dout(new_Jinkela_wire_5507)
    );

    bfr new_Jinkela_buffer_827 (
        .din(_1046_),
        .dout(new_Jinkela_wire_1583)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_1364),
        .dout(new_Jinkela_wire_1365)
    );

    bfr new_Jinkela_buffer_4196 (
        .din(new_Jinkela_wire_5507),
        .dout(new_Jinkela_wire_5508)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_1578),
        .dout(new_Jinkela_wire_1579)
    );

    spl2 new_Jinkela_splitter_520 (
        .a(_0656_),
        .b(new_Jinkela_wire_5697),
        .c(new_Jinkela_wire_5698)
    );

    bfr new_Jinkela_buffer_4242 (
        .din(new_Jinkela_wire_5565),
        .dout(new_Jinkela_wire_5566)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_1411),
        .dout(new_Jinkela_wire_1412)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_1365),
        .dout(new_Jinkela_wire_1366)
    );

    bfr new_Jinkela_buffer_4197 (
        .din(new_Jinkela_wire_5508),
        .dout(new_Jinkela_wire_5509)
    );

    bfr new_Jinkela_buffer_4345 (
        .din(new_Jinkela_wire_5674),
        .dout(new_Jinkela_wire_5675)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(_1570_),
        .b(new_Jinkela_wire_1584),
        .c(new_Jinkela_wire_1585)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_1366),
        .dout(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_4198 (
        .din(new_Jinkela_wire_5509),
        .dout(new_Jinkela_wire_5510)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(_0162_),
        .b(new_Jinkela_wire_1586),
        .c(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_4243 (
        .din(new_Jinkela_wire_5566),
        .dout(new_Jinkela_wire_5567)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_1412),
        .dout(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_1367),
        .dout(new_Jinkela_wire_1368)
    );

    bfr new_Jinkela_buffer_4199 (
        .din(new_Jinkela_wire_5510),
        .dout(new_Jinkela_wire_5511)
    );

    bfr new_Jinkela_buffer_4352 (
        .din(new_Jinkela_wire_5691),
        .dout(new_Jinkela_wire_5692)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_1368),
        .dout(new_Jinkela_wire_1369)
    );

    bfr new_Jinkela_buffer_4200 (
        .din(new_Jinkela_wire_5511),
        .dout(new_Jinkela_wire_5512)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_4244 (
        .din(new_Jinkela_wire_5567),
        .dout(new_Jinkela_wire_5568)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_1413),
        .dout(new_Jinkela_wire_1414)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_1369),
        .dout(new_Jinkela_wire_1370)
    );

    bfr new_Jinkela_buffer_4201 (
        .din(new_Jinkela_wire_5512),
        .dout(new_Jinkela_wire_5513)
    );

    bfr new_Jinkela_buffer_14616 (
        .din(new_Jinkela_wire_17446),
        .dout(new_Jinkela_wire_17447)
    );

    bfr new_Jinkela_buffer_14486 (
        .din(new_Jinkela_wire_17300),
        .dout(new_Jinkela_wire_17301)
    );

    bfr new_Jinkela_buffer_14591 (
        .din(new_Jinkela_wire_17417),
        .dout(new_Jinkela_wire_17418)
    );

    bfr new_Jinkela_buffer_14487 (
        .din(new_Jinkela_wire_17301),
        .dout(new_Jinkela_wire_17302)
    );

    bfr new_Jinkela_buffer_14708 (
        .din(new_Jinkela_wire_17558),
        .dout(new_Jinkela_wire_17559)
    );

    bfr new_Jinkela_buffer_14488 (
        .din(new_Jinkela_wire_17302),
        .dout(new_Jinkela_wire_17303)
    );

    bfr new_Jinkela_buffer_14592 (
        .din(new_Jinkela_wire_17418),
        .dout(new_Jinkela_wire_17419)
    );

    bfr new_Jinkela_buffer_14489 (
        .din(new_Jinkela_wire_17303),
        .dout(new_Jinkela_wire_17304)
    );

    bfr new_Jinkela_buffer_14617 (
        .din(new_Jinkela_wire_17447),
        .dout(new_Jinkela_wire_17448)
    );

    bfr new_Jinkela_buffer_14490 (
        .din(new_Jinkela_wire_17304),
        .dout(new_Jinkela_wire_17305)
    );

    bfr new_Jinkela_buffer_14593 (
        .din(new_Jinkela_wire_17419),
        .dout(new_Jinkela_wire_17420)
    );

    bfr new_Jinkela_buffer_14491 (
        .din(new_Jinkela_wire_17305),
        .dout(new_Jinkela_wire_17306)
    );

    bfr new_Jinkela_buffer_14784 (
        .din(new_Jinkela_wire_17638),
        .dout(new_Jinkela_wire_17639)
    );

    bfr new_Jinkela_buffer_14492 (
        .din(new_Jinkela_wire_17306),
        .dout(new_Jinkela_wire_17307)
    );

    spl2 new_Jinkela_splitter_1262 (
        .a(new_Jinkela_wire_17420),
        .b(new_Jinkela_wire_17421),
        .c(new_Jinkela_wire_17422)
    );

    bfr new_Jinkela_buffer_14493 (
        .din(new_Jinkela_wire_17307),
        .dout(new_Jinkela_wire_17308)
    );

    bfr new_Jinkela_buffer_14709 (
        .din(new_Jinkela_wire_17559),
        .dout(new_Jinkela_wire_17560)
    );

    bfr new_Jinkela_buffer_14494 (
        .din(new_Jinkela_wire_17308),
        .dout(new_Jinkela_wire_17309)
    );

    bfr new_Jinkela_buffer_14618 (
        .din(new_Jinkela_wire_17448),
        .dout(new_Jinkela_wire_17449)
    );

    bfr new_Jinkela_buffer_14495 (
        .din(new_Jinkela_wire_17309),
        .dout(new_Jinkela_wire_17310)
    );

    bfr new_Jinkela_buffer_14619 (
        .din(new_Jinkela_wire_17449),
        .dout(new_Jinkela_wire_17450)
    );

    bfr new_Jinkela_buffer_14496 (
        .din(new_Jinkela_wire_17310),
        .dout(new_Jinkela_wire_17311)
    );

    spl2 new_Jinkela_splitter_1280 (
        .a(_1633_),
        .b(new_Jinkela_wire_17662),
        .c(new_Jinkela_wire_17663)
    );

    bfr new_Jinkela_buffer_14497 (
        .din(new_Jinkela_wire_17311),
        .dout(new_Jinkela_wire_17312)
    );

    bfr new_Jinkela_buffer_14620 (
        .din(new_Jinkela_wire_17450),
        .dout(new_Jinkela_wire_17451)
    );

    bfr new_Jinkela_buffer_14498 (
        .din(new_Jinkela_wire_17312),
        .dout(new_Jinkela_wire_17313)
    );

    bfr new_Jinkela_buffer_14710 (
        .din(new_Jinkela_wire_17560),
        .dout(new_Jinkela_wire_17561)
    );

    bfr new_Jinkela_buffer_14499 (
        .din(new_Jinkela_wire_17313),
        .dout(new_Jinkela_wire_17314)
    );

    bfr new_Jinkela_buffer_14621 (
        .din(new_Jinkela_wire_17451),
        .dout(new_Jinkela_wire_17452)
    );

    bfr new_Jinkela_buffer_14500 (
        .din(new_Jinkela_wire_17314),
        .dout(new_Jinkela_wire_17315)
    );

    bfr new_Jinkela_buffer_14785 (
        .din(new_Jinkela_wire_17639),
        .dout(new_Jinkela_wire_17640)
    );

    bfr new_Jinkela_buffer_14501 (
        .din(new_Jinkela_wire_17315),
        .dout(new_Jinkela_wire_17316)
    );

    bfr new_Jinkela_buffer_14622 (
        .din(new_Jinkela_wire_17452),
        .dout(new_Jinkela_wire_17453)
    );

    bfr new_Jinkela_buffer_14711 (
        .din(new_Jinkela_wire_17561),
        .dout(new_Jinkela_wire_17562)
    );

    bfr new_Jinkela_buffer_14623 (
        .din(new_Jinkela_wire_17453),
        .dout(new_Jinkela_wire_17454)
    );

    spl2 new_Jinkela_splitter_1279 (
        .a(_0014_),
        .b(new_Jinkela_wire_17660),
        .c(new_Jinkela_wire_17661)
    );

    bfr new_Jinkela_buffer_14624 (
        .din(new_Jinkela_wire_17454),
        .dout(new_Jinkela_wire_17455)
    );

    bfr new_Jinkela_buffer_14712 (
        .din(new_Jinkela_wire_17562),
        .dout(new_Jinkela_wire_17563)
    );

    bfr new_Jinkela_buffer_14625 (
        .din(new_Jinkela_wire_17455),
        .dout(new_Jinkela_wire_17456)
    );

    bfr new_Jinkela_buffer_14786 (
        .din(new_Jinkela_wire_17640),
        .dout(new_Jinkela_wire_17641)
    );

    bfr new_Jinkela_buffer_14626 (
        .din(new_Jinkela_wire_17456),
        .dout(new_Jinkela_wire_17457)
    );

    bfr new_Jinkela_buffer_7655 (
        .din(new_Jinkela_wire_9482),
        .dout(new_Jinkela_wire_9483)
    );

    bfr new_Jinkela_buffer_7613 (
        .din(new_Jinkela_wire_9436),
        .dout(new_Jinkela_wire_9437)
    );

    bfr new_Jinkela_buffer_7716 (
        .din(new_Jinkela_wire_9559),
        .dout(new_Jinkela_wire_9560)
    );

    bfr new_Jinkela_buffer_7614 (
        .din(new_Jinkela_wire_9437),
        .dout(new_Jinkela_wire_9438)
    );

    bfr new_Jinkela_buffer_7656 (
        .din(new_Jinkela_wire_9483),
        .dout(new_Jinkela_wire_9484)
    );

    bfr new_Jinkela_buffer_7615 (
        .din(new_Jinkela_wire_9438),
        .dout(new_Jinkela_wire_9439)
    );

    bfr new_Jinkela_buffer_7704 (
        .din(new_Jinkela_wire_9535),
        .dout(new_Jinkela_wire_9536)
    );

    bfr new_Jinkela_buffer_7616 (
        .din(new_Jinkela_wire_9439),
        .dout(new_Jinkela_wire_9440)
    );

    bfr new_Jinkela_buffer_7657 (
        .din(new_Jinkela_wire_9484),
        .dout(new_Jinkela_wire_9485)
    );

    bfr new_Jinkela_buffer_7617 (
        .din(new_Jinkela_wire_9440),
        .dout(new_Jinkela_wire_9441)
    );

    bfr new_Jinkela_buffer_7714 (
        .din(new_Jinkela_wire_9553),
        .dout(new_Jinkela_wire_9554)
    );

    bfr new_Jinkela_buffer_7618 (
        .din(new_Jinkela_wire_9441),
        .dout(new_Jinkela_wire_9442)
    );

    bfr new_Jinkela_buffer_7658 (
        .din(new_Jinkela_wire_9485),
        .dout(new_Jinkela_wire_9486)
    );

    bfr new_Jinkela_buffer_7619 (
        .din(new_Jinkela_wire_9442),
        .dout(new_Jinkela_wire_9443)
    );

    bfr new_Jinkela_buffer_7705 (
        .din(new_Jinkela_wire_9536),
        .dout(new_Jinkela_wire_9537)
    );

    spl2 new_Jinkela_splitter_761 (
        .a(new_Jinkela_wire_9443),
        .b(new_Jinkela_wire_9444),
        .c(new_Jinkela_wire_9445)
    );

    bfr new_Jinkela_buffer_7721 (
        .din(_1024_),
        .dout(new_Jinkela_wire_9565)
    );

    bfr new_Jinkela_buffer_7659 (
        .din(new_Jinkela_wire_9486),
        .dout(new_Jinkela_wire_9487)
    );

    bfr new_Jinkela_buffer_7660 (
        .din(new_Jinkela_wire_9487),
        .dout(new_Jinkela_wire_9488)
    );

    bfr new_Jinkela_buffer_7706 (
        .din(new_Jinkela_wire_9537),
        .dout(new_Jinkela_wire_9538)
    );

    bfr new_Jinkela_buffer_7661 (
        .din(new_Jinkela_wire_9488),
        .dout(new_Jinkela_wire_9489)
    );

    bfr new_Jinkela_buffer_7715 (
        .din(new_Jinkela_wire_9554),
        .dout(new_Jinkela_wire_9555)
    );

    bfr new_Jinkela_buffer_7662 (
        .din(new_Jinkela_wire_9489),
        .dout(new_Jinkela_wire_9490)
    );

    spl2 new_Jinkela_splitter_765 (
        .a(new_Jinkela_wire_9538),
        .b(new_Jinkela_wire_9539),
        .c(new_Jinkela_wire_9540)
    );

    bfr new_Jinkela_buffer_7663 (
        .din(new_Jinkela_wire_9490),
        .dout(new_Jinkela_wire_9491)
    );

    bfr new_Jinkela_buffer_7717 (
        .din(new_Jinkela_wire_9560),
        .dout(new_Jinkela_wire_9561)
    );

    bfr new_Jinkela_buffer_7664 (
        .din(new_Jinkela_wire_9491),
        .dout(new_Jinkela_wire_9492)
    );

    spl2 new_Jinkela_splitter_772 (
        .a(_1359_),
        .b(new_Jinkela_wire_9599),
        .c(new_Jinkela_wire_9600)
    );

    bfr new_Jinkela_buffer_7665 (
        .din(new_Jinkela_wire_9492),
        .dout(new_Jinkela_wire_9493)
    );

    spl2 new_Jinkela_splitter_773 (
        .a(_1441_),
        .b(new_Jinkela_wire_9601),
        .c(new_Jinkela_wire_9602)
    );

    bfr new_Jinkela_buffer_7666 (
        .din(new_Jinkela_wire_9493),
        .dout(new_Jinkela_wire_9494)
    );

    bfr new_Jinkela_buffer_7718 (
        .din(new_Jinkela_wire_9561),
        .dout(new_Jinkela_wire_9562)
    );

    bfr new_Jinkela_buffer_7667 (
        .din(new_Jinkela_wire_9494),
        .dout(new_Jinkela_wire_9495)
    );

    bfr new_Jinkela_buffer_7722 (
        .din(new_Jinkela_wire_9565),
        .dout(new_Jinkela_wire_9566)
    );

    bfr new_Jinkela_buffer_7668 (
        .din(new_Jinkela_wire_9495),
        .dout(new_Jinkela_wire_9496)
    );

    bfr new_Jinkela_buffer_7719 (
        .din(new_Jinkela_wire_9562),
        .dout(new_Jinkela_wire_9563)
    );

    bfr new_Jinkela_buffer_7669 (
        .din(new_Jinkela_wire_9496),
        .dout(new_Jinkela_wire_9497)
    );

    bfr new_Jinkela_buffer_7753 (
        .din(new_Jinkela_wire_9602),
        .dout(new_Jinkela_wire_9603)
    );

    bfr new_Jinkela_buffer_7670 (
        .din(new_Jinkela_wire_9497),
        .dout(new_Jinkela_wire_9498)
    );

    bfr new_Jinkela_buffer_7723 (
        .din(new_Jinkela_wire_9566),
        .dout(new_Jinkela_wire_9567)
    );

    bfr new_Jinkela_buffer_7671 (
        .din(new_Jinkela_wire_9498),
        .dout(new_Jinkela_wire_9499)
    );

    spl2 new_Jinkela_splitter_774 (
        .a(_0121_),
        .b(new_Jinkela_wire_9607),
        .c(new_Jinkela_wire_9608)
    );

    bfr new_Jinkela_buffer_11164 (
        .din(new_Jinkela_wire_13469),
        .dout(new_Jinkela_wire_13470)
    );

    bfr new_Jinkela_buffer_11129 (
        .din(new_Jinkela_wire_13426),
        .dout(new_Jinkela_wire_13427)
    );

    bfr new_Jinkela_buffer_11130 (
        .din(new_Jinkela_wire_13427),
        .dout(new_Jinkela_wire_13428)
    );

    bfr new_Jinkela_buffer_11165 (
        .din(new_Jinkela_wire_13470),
        .dout(new_Jinkela_wire_13471)
    );

    bfr new_Jinkela_buffer_11131 (
        .din(new_Jinkela_wire_13428),
        .dout(new_Jinkela_wire_13429)
    );

    bfr new_Jinkela_buffer_11265 (
        .din(new_Jinkela_wire_13576),
        .dout(new_Jinkela_wire_13577)
    );

    bfr new_Jinkela_buffer_11132 (
        .din(new_Jinkela_wire_13429),
        .dout(new_Jinkela_wire_13430)
    );

    bfr new_Jinkela_buffer_11166 (
        .din(new_Jinkela_wire_13471),
        .dout(new_Jinkela_wire_13472)
    );

    bfr new_Jinkela_buffer_11133 (
        .din(new_Jinkela_wire_13430),
        .dout(new_Jinkela_wire_13431)
    );

    bfr new_Jinkela_buffer_11134 (
        .din(new_Jinkela_wire_13431),
        .dout(new_Jinkela_wire_13432)
    );

    spl2 new_Jinkela_splitter_1007 (
        .a(_1006_),
        .b(new_Jinkela_wire_13584),
        .c(new_Jinkela_wire_13585)
    );

    bfr new_Jinkela_buffer_11167 (
        .din(new_Jinkela_wire_13472),
        .dout(new_Jinkela_wire_13473)
    );

    bfr new_Jinkela_buffer_11135 (
        .din(new_Jinkela_wire_13432),
        .dout(new_Jinkela_wire_13433)
    );

    bfr new_Jinkela_buffer_11266 (
        .din(new_Jinkela_wire_13577),
        .dout(new_Jinkela_wire_13578)
    );

    bfr new_Jinkela_buffer_11136 (
        .din(new_Jinkela_wire_13433),
        .dout(new_Jinkela_wire_13434)
    );

    bfr new_Jinkela_buffer_11168 (
        .din(new_Jinkela_wire_13473),
        .dout(new_Jinkela_wire_13474)
    );

    bfr new_Jinkela_buffer_11137 (
        .din(new_Jinkela_wire_13434),
        .dout(new_Jinkela_wire_13435)
    );

    bfr new_Jinkela_buffer_11269 (
        .din(new_Jinkela_wire_13588),
        .dout(new_Jinkela_wire_13589)
    );

    bfr new_Jinkela_buffer_11138 (
        .din(new_Jinkela_wire_13435),
        .dout(new_Jinkela_wire_13436)
    );

    bfr new_Jinkela_buffer_11268 (
        .din(_1424_),
        .dout(new_Jinkela_wire_13586)
    );

    bfr new_Jinkela_buffer_11169 (
        .din(new_Jinkela_wire_13474),
        .dout(new_Jinkela_wire_13475)
    );

    bfr new_Jinkela_buffer_11139 (
        .din(new_Jinkela_wire_13436),
        .dout(new_Jinkela_wire_13437)
    );

    bfr new_Jinkela_buffer_11267 (
        .din(new_Jinkela_wire_13578),
        .dout(new_Jinkela_wire_13579)
    );

    bfr new_Jinkela_buffer_11140 (
        .din(new_Jinkela_wire_13437),
        .dout(new_Jinkela_wire_13438)
    );

    bfr new_Jinkela_buffer_11170 (
        .din(new_Jinkela_wire_13475),
        .dout(new_Jinkela_wire_13476)
    );

    bfr new_Jinkela_buffer_11141 (
        .din(new_Jinkela_wire_13438),
        .dout(new_Jinkela_wire_13439)
    );

    bfr new_Jinkela_buffer_11273 (
        .din(_0538_),
        .dout(new_Jinkela_wire_13593)
    );

    bfr new_Jinkela_buffer_11142 (
        .din(new_Jinkela_wire_13439),
        .dout(new_Jinkela_wire_13440)
    );

    spl2 new_Jinkela_splitter_1008 (
        .a(_0186_),
        .b(new_Jinkela_wire_13587),
        .c(new_Jinkela_wire_13588)
    );

    bfr new_Jinkela_buffer_11171 (
        .din(new_Jinkela_wire_13476),
        .dout(new_Jinkela_wire_13477)
    );

    bfr new_Jinkela_buffer_11143 (
        .din(new_Jinkela_wire_13440),
        .dout(new_Jinkela_wire_13441)
    );

    bfr new_Jinkela_buffer_11144 (
        .din(new_Jinkela_wire_13441),
        .dout(new_Jinkela_wire_13442)
    );

    bfr new_Jinkela_buffer_11172 (
        .din(new_Jinkela_wire_13477),
        .dout(new_Jinkela_wire_13478)
    );

    bfr new_Jinkela_buffer_11145 (
        .din(new_Jinkela_wire_13442),
        .dout(new_Jinkela_wire_13443)
    );

    bfr new_Jinkela_buffer_11146 (
        .din(new_Jinkela_wire_13443),
        .dout(new_Jinkela_wire_13444)
    );

    spl2 new_Jinkela_splitter_1010 (
        .a(_0048_),
        .b(new_Jinkela_wire_13675),
        .c(new_Jinkela_wire_13676)
    );

    bfr new_Jinkela_buffer_11173 (
        .din(new_Jinkela_wire_13478),
        .dout(new_Jinkela_wire_13479)
    );

    bfr new_Jinkela_buffer_11147 (
        .din(new_Jinkela_wire_13444),
        .dout(new_Jinkela_wire_13445)
    );

    bfr new_Jinkela_buffer_11148 (
        .din(new_Jinkela_wire_13445),
        .dout(new_Jinkela_wire_13446)
    );

    bfr new_Jinkela_buffer_11353 (
        .din(_0855_),
        .dout(new_Jinkela_wire_13677)
    );

    bfr new_Jinkela_buffer_11174 (
        .din(new_Jinkela_wire_13479),
        .dout(new_Jinkela_wire_13480)
    );

    bfr new_Jinkela_buffer_11149 (
        .din(new_Jinkela_wire_13446),
        .dout(new_Jinkela_wire_13447)
    );

    bfr new_Jinkela_buffer_11270 (
        .din(new_Jinkela_wire_13589),
        .dout(new_Jinkela_wire_13590)
    );

    bfr new_Jinkela_buffer_11150 (
        .din(new_Jinkela_wire_13447),
        .dout(new_Jinkela_wire_13448)
    );

    bfr new_Jinkela_buffer_4346 (
        .din(new_Jinkela_wire_5675),
        .dout(new_Jinkela_wire_5676)
    );

    bfr new_Jinkela_buffer_4202 (
        .din(new_Jinkela_wire_5513),
        .dout(new_Jinkela_wire_5514)
    );

    bfr new_Jinkela_buffer_11175 (
        .din(new_Jinkela_wire_13480),
        .dout(new_Jinkela_wire_13481)
    );

    bfr new_Jinkela_buffer_11151 (
        .din(new_Jinkela_wire_13448),
        .dout(new_Jinkela_wire_13449)
    );

    bfr new_Jinkela_buffer_4245 (
        .din(new_Jinkela_wire_5568),
        .dout(new_Jinkela_wire_5569)
    );

    bfr new_Jinkela_buffer_4203 (
        .din(new_Jinkela_wire_5514),
        .dout(new_Jinkela_wire_5515)
    );

    bfr new_Jinkela_buffer_11274 (
        .din(new_Jinkela_wire_13593),
        .dout(new_Jinkela_wire_13594)
    );

    bfr new_Jinkela_buffer_11152 (
        .din(new_Jinkela_wire_13449),
        .dout(new_Jinkela_wire_13450)
    );

    bfr new_Jinkela_buffer_4355 (
        .din(new_Jinkela_wire_5698),
        .dout(new_Jinkela_wire_5699)
    );

    bfr new_Jinkela_buffer_4204 (
        .din(new_Jinkela_wire_5515),
        .dout(new_Jinkela_wire_5516)
    );

    bfr new_Jinkela_buffer_11176 (
        .din(new_Jinkela_wire_13481),
        .dout(new_Jinkela_wire_13482)
    );

    bfr new_Jinkela_buffer_11153 (
        .din(new_Jinkela_wire_13450),
        .dout(new_Jinkela_wire_13451)
    );

    bfr new_Jinkela_buffer_4246 (
        .din(new_Jinkela_wire_5569),
        .dout(new_Jinkela_wire_5570)
    );

    bfr new_Jinkela_buffer_4205 (
        .din(new_Jinkela_wire_5516),
        .dout(new_Jinkela_wire_5517)
    );

    bfr new_Jinkela_buffer_11271 (
        .din(new_Jinkela_wire_13590),
        .dout(new_Jinkela_wire_13591)
    );

    bfr new_Jinkela_buffer_11154 (
        .din(new_Jinkela_wire_13451),
        .dout(new_Jinkela_wire_13452)
    );

    bfr new_Jinkela_buffer_4347 (
        .din(new_Jinkela_wire_5676),
        .dout(new_Jinkela_wire_5677)
    );

    bfr new_Jinkela_buffer_4206 (
        .din(new_Jinkela_wire_5517),
        .dout(new_Jinkela_wire_5518)
    );

    bfr new_Jinkela_buffer_11177 (
        .din(new_Jinkela_wire_13482),
        .dout(new_Jinkela_wire_13483)
    );

    bfr new_Jinkela_buffer_11155 (
        .din(new_Jinkela_wire_13452),
        .dout(new_Jinkela_wire_13453)
    );

    bfr new_Jinkela_buffer_4247 (
        .din(new_Jinkela_wire_5570),
        .dout(new_Jinkela_wire_5571)
    );

    bfr new_Jinkela_buffer_4207 (
        .din(new_Jinkela_wire_5518),
        .dout(new_Jinkela_wire_5519)
    );

    bfr new_Jinkela_buffer_11156 (
        .din(new_Jinkela_wire_13453),
        .dout(new_Jinkela_wire_13454)
    );

    bfr new_Jinkela_buffer_4353 (
        .din(new_Jinkela_wire_5692),
        .dout(new_Jinkela_wire_5693)
    );

    bfr new_Jinkela_buffer_4208 (
        .din(new_Jinkela_wire_5519),
        .dout(new_Jinkela_wire_5520)
    );

    spl2 new_Jinkela_splitter_1011 (
        .a(_0755_),
        .b(new_Jinkela_wire_13679),
        .c(new_Jinkela_wire_13680)
    );

    bfr new_Jinkela_buffer_11178 (
        .din(new_Jinkela_wire_13483),
        .dout(new_Jinkela_wire_13484)
    );

    bfr new_Jinkela_buffer_4248 (
        .din(new_Jinkela_wire_5571),
        .dout(new_Jinkela_wire_5572)
    );

    bfr new_Jinkela_buffer_11272 (
        .din(new_Jinkela_wire_13591),
        .dout(new_Jinkela_wire_13592)
    );

    bfr new_Jinkela_buffer_4209 (
        .din(new_Jinkela_wire_5520),
        .dout(new_Jinkela_wire_5521)
    );

    bfr new_Jinkela_buffer_11179 (
        .din(new_Jinkela_wire_13484),
        .dout(new_Jinkela_wire_13485)
    );

    bfr new_Jinkela_buffer_4348 (
        .din(new_Jinkela_wire_5677),
        .dout(new_Jinkela_wire_5678)
    );

    bfr new_Jinkela_buffer_11275 (
        .din(new_Jinkela_wire_13594),
        .dout(new_Jinkela_wire_13595)
    );

    bfr new_Jinkela_buffer_4210 (
        .din(new_Jinkela_wire_5521),
        .dout(new_Jinkela_wire_5522)
    );

    bfr new_Jinkela_buffer_11180 (
        .din(new_Jinkela_wire_13485),
        .dout(new_Jinkela_wire_13486)
    );

    bfr new_Jinkela_buffer_4249 (
        .din(new_Jinkela_wire_5572),
        .dout(new_Jinkela_wire_5573)
    );

    bfr new_Jinkela_buffer_4211 (
        .din(new_Jinkela_wire_5522),
        .dout(new_Jinkela_wire_5523)
    );

    bfr new_Jinkela_buffer_11354 (
        .din(_0724_),
        .dout(new_Jinkela_wire_13678)
    );

    bfr new_Jinkela_buffer_11181 (
        .din(new_Jinkela_wire_13486),
        .dout(new_Jinkela_wire_13487)
    );

    bfr new_Jinkela_buffer_11276 (
        .din(new_Jinkela_wire_13595),
        .dout(new_Jinkela_wire_13596)
    );

    bfr new_Jinkela_buffer_4212 (
        .din(new_Jinkela_wire_5523),
        .dout(new_Jinkela_wire_5524)
    );

    bfr new_Jinkela_buffer_11182 (
        .din(new_Jinkela_wire_13487),
        .dout(new_Jinkela_wire_13488)
    );

    bfr new_Jinkela_buffer_4360 (
        .din(_0718_),
        .dout(new_Jinkela_wire_5704)
    );

    bfr new_Jinkela_buffer_4250 (
        .din(new_Jinkela_wire_5573),
        .dout(new_Jinkela_wire_5574)
    );

    spl2 new_Jinkela_splitter_1012 (
        .a(_0695_),
        .b(new_Jinkela_wire_13681),
        .c(new_Jinkela_wire_13682)
    );

    bfr new_Jinkela_buffer_4213 (
        .din(new_Jinkela_wire_5524),
        .dout(new_Jinkela_wire_5525)
    );

    bfr new_Jinkela_buffer_11183 (
        .din(new_Jinkela_wire_13488),
        .dout(new_Jinkela_wire_13489)
    );

    bfr new_Jinkela_buffer_4349 (
        .din(new_Jinkela_wire_5678),
        .dout(new_Jinkela_wire_5679)
    );

    bfr new_Jinkela_buffer_11277 (
        .din(new_Jinkela_wire_13596),
        .dout(new_Jinkela_wire_13597)
    );

    bfr new_Jinkela_buffer_4214 (
        .din(new_Jinkela_wire_5525),
        .dout(new_Jinkela_wire_5526)
    );

    bfr new_Jinkela_buffer_11184 (
        .din(new_Jinkela_wire_13489),
        .dout(new_Jinkela_wire_13490)
    );

    bfr new_Jinkela_buffer_4251 (
        .din(new_Jinkela_wire_5574),
        .dout(new_Jinkela_wire_5575)
    );

    bfr new_Jinkela_buffer_4215 (
        .din(new_Jinkela_wire_5526),
        .dout(new_Jinkela_wire_5527)
    );

    bfr new_Jinkela_buffer_11185 (
        .din(new_Jinkela_wire_13490),
        .dout(new_Jinkela_wire_13491)
    );

    bfr new_Jinkela_buffer_4354 (
        .din(new_Jinkela_wire_5693),
        .dout(new_Jinkela_wire_5694)
    );

    bfr new_Jinkela_buffer_11278 (
        .din(new_Jinkela_wire_13597),
        .dout(new_Jinkela_wire_13598)
    );

    bfr new_Jinkela_buffer_4216 (
        .din(new_Jinkela_wire_5527),
        .dout(new_Jinkela_wire_5528)
    );

    bfr new_Jinkela_buffer_11186 (
        .din(new_Jinkela_wire_13491),
        .dout(new_Jinkela_wire_13492)
    );

    bfr new_Jinkela_buffer_4252 (
        .din(new_Jinkela_wire_5575),
        .dout(new_Jinkela_wire_5576)
    );

    bfr new_Jinkela_buffer_4217 (
        .din(new_Jinkela_wire_5528),
        .dout(new_Jinkela_wire_5529)
    );

    spl2 new_Jinkela_splitter_1013 (
        .a(_0593_),
        .b(new_Jinkela_wire_13683),
        .c(new_Jinkela_wire_13684)
    );

    bfr new_Jinkela_buffer_11187 (
        .din(new_Jinkela_wire_13492),
        .dout(new_Jinkela_wire_13493)
    );

    bfr new_Jinkela_buffer_4350 (
        .din(new_Jinkela_wire_5679),
        .dout(new_Jinkela_wire_5680)
    );

    bfr new_Jinkela_buffer_11279 (
        .din(new_Jinkela_wire_13598),
        .dout(new_Jinkela_wire_13599)
    );

    bfr new_Jinkela_buffer_4218 (
        .din(new_Jinkela_wire_5529),
        .dout(new_Jinkela_wire_5530)
    );

    bfr new_Jinkela_buffer_11188 (
        .din(new_Jinkela_wire_13493),
        .dout(new_Jinkela_wire_13494)
    );

    bfr new_Jinkela_buffer_4253 (
        .din(new_Jinkela_wire_5576),
        .dout(new_Jinkela_wire_5577)
    );

    bfr new_Jinkela_buffer_11355 (
        .din(new_Jinkela_wire_13686),
        .dout(new_Jinkela_wire_13687)
    );

    bfr new_Jinkela_buffer_4219 (
        .din(new_Jinkela_wire_5530),
        .dout(new_Jinkela_wire_5531)
    );

    spl2 new_Jinkela_splitter_1014 (
        .a(_1536_),
        .b(new_Jinkela_wire_13685),
        .c(new_Jinkela_wire_13686)
    );

    bfr new_Jinkela_buffer_11189 (
        .din(new_Jinkela_wire_13494),
        .dout(new_Jinkela_wire_13495)
    );

    bfr new_Jinkela_buffer_4364 (
        .din(_0793_),
        .dout(new_Jinkela_wire_5710)
    );

    bfr new_Jinkela_buffer_11280 (
        .din(new_Jinkela_wire_13599),
        .dout(new_Jinkela_wire_13600)
    );

    bfr new_Jinkela_buffer_4220 (
        .din(new_Jinkela_wire_5531),
        .dout(new_Jinkela_wire_5532)
    );

    bfr new_Jinkela_buffer_11190 (
        .din(new_Jinkela_wire_13495),
        .dout(new_Jinkela_wire_13496)
    );

    bfr new_Jinkela_buffer_4254 (
        .din(new_Jinkela_wire_5577),
        .dout(new_Jinkela_wire_5578)
    );

    bfr new_Jinkela_buffer_4221 (
        .din(new_Jinkela_wire_5532),
        .dout(new_Jinkela_wire_5533)
    );

    spl2 new_Jinkela_splitter_1015 (
        .a(_0766_),
        .b(new_Jinkela_wire_13691),
        .c(new_Jinkela_wire_13692)
    );

    bfr new_Jinkela_buffer_11191 (
        .din(new_Jinkela_wire_13496),
        .dout(new_Jinkela_wire_13497)
    );

    spl2 new_Jinkela_splitter_519 (
        .a(new_Jinkela_wire_5694),
        .b(new_Jinkela_wire_5695),
        .c(new_Jinkela_wire_5696)
    );

    bfr new_Jinkela_buffer_11281 (
        .din(new_Jinkela_wire_13600),
        .dout(new_Jinkela_wire_13601)
    );

    bfr new_Jinkela_buffer_4222 (
        .din(new_Jinkela_wire_5533),
        .dout(new_Jinkela_wire_5534)
    );

    bfr new_Jinkela_buffer_7672 (
        .din(new_Jinkela_wire_9499),
        .dout(new_Jinkela_wire_9500)
    );

    bfr new_Jinkela_buffer_7724 (
        .din(new_Jinkela_wire_9567),
        .dout(new_Jinkela_wire_9568)
    );

    bfr new_Jinkela_buffer_7673 (
        .din(new_Jinkela_wire_9500),
        .dout(new_Jinkela_wire_9501)
    );

    spl2 new_Jinkela_splitter_775 (
        .a(_0210_),
        .b(new_Jinkela_wire_9609),
        .c(new_Jinkela_wire_9610)
    );

    bfr new_Jinkela_buffer_7674 (
        .din(new_Jinkela_wire_9501),
        .dout(new_Jinkela_wire_9502)
    );

    bfr new_Jinkela_buffer_7725 (
        .din(new_Jinkela_wire_9568),
        .dout(new_Jinkela_wire_9569)
    );

    bfr new_Jinkela_buffer_7675 (
        .din(new_Jinkela_wire_9502),
        .dout(new_Jinkela_wire_9503)
    );

    bfr new_Jinkela_buffer_7676 (
        .din(new_Jinkela_wire_9503),
        .dout(new_Jinkela_wire_9504)
    );

    bfr new_Jinkela_buffer_7726 (
        .din(new_Jinkela_wire_9569),
        .dout(new_Jinkela_wire_9570)
    );

    bfr new_Jinkela_buffer_7677 (
        .din(new_Jinkela_wire_9504),
        .dout(new_Jinkela_wire_9505)
    );

    bfr new_Jinkela_buffer_7754 (
        .din(new_Jinkela_wire_9603),
        .dout(new_Jinkela_wire_9604)
    );

    bfr new_Jinkela_buffer_7678 (
        .din(new_Jinkela_wire_9505),
        .dout(new_Jinkela_wire_9506)
    );

    bfr new_Jinkela_buffer_7727 (
        .din(new_Jinkela_wire_9570),
        .dout(new_Jinkela_wire_9571)
    );

    bfr new_Jinkela_buffer_7679 (
        .din(new_Jinkela_wire_9506),
        .dout(new_Jinkela_wire_9507)
    );

    bfr new_Jinkela_buffer_7840 (
        .din(_0104_),
        .dout(new_Jinkela_wire_9696)
    );

    bfr new_Jinkela_buffer_7757 (
        .din(_0888_),
        .dout(new_Jinkela_wire_9611)
    );

    bfr new_Jinkela_buffer_7680 (
        .din(new_Jinkela_wire_9507),
        .dout(new_Jinkela_wire_9508)
    );

    bfr new_Jinkela_buffer_7728 (
        .din(new_Jinkela_wire_9571),
        .dout(new_Jinkela_wire_9572)
    );

    bfr new_Jinkela_buffer_7681 (
        .din(new_Jinkela_wire_9508),
        .dout(new_Jinkela_wire_9509)
    );

    bfr new_Jinkela_buffer_7755 (
        .din(new_Jinkela_wire_9604),
        .dout(new_Jinkela_wire_9605)
    );

    bfr new_Jinkela_buffer_7729 (
        .din(new_Jinkela_wire_9572),
        .dout(new_Jinkela_wire_9573)
    );

    bfr new_Jinkela_buffer_7839 (
        .din(_0750_),
        .dout(new_Jinkela_wire_9695)
    );

    bfr new_Jinkela_buffer_7730 (
        .din(new_Jinkela_wire_9573),
        .dout(new_Jinkela_wire_9574)
    );

    bfr new_Jinkela_buffer_7756 (
        .din(new_Jinkela_wire_9605),
        .dout(new_Jinkela_wire_9606)
    );

    bfr new_Jinkela_buffer_7731 (
        .din(new_Jinkela_wire_9574),
        .dout(new_Jinkela_wire_9575)
    );

    bfr new_Jinkela_buffer_7758 (
        .din(new_Jinkela_wire_9611),
        .dout(new_Jinkela_wire_9612)
    );

    bfr new_Jinkela_buffer_7732 (
        .din(new_Jinkela_wire_9575),
        .dout(new_Jinkela_wire_9576)
    );

    spl2 new_Jinkela_splitter_778 (
        .a(_0882_),
        .b(new_Jinkela_wire_9738),
        .c(new_Jinkela_wire_9739)
    );

    bfr new_Jinkela_buffer_7733 (
        .din(new_Jinkela_wire_9576),
        .dout(new_Jinkela_wire_9577)
    );

    bfr new_Jinkela_buffer_7759 (
        .din(new_Jinkela_wire_9612),
        .dout(new_Jinkela_wire_9613)
    );

    bfr new_Jinkela_buffer_7734 (
        .din(new_Jinkela_wire_9577),
        .dout(new_Jinkela_wire_9578)
    );

    spl2 new_Jinkela_splitter_779 (
        .a(_1224_),
        .b(new_Jinkela_wire_9740),
        .c(new_Jinkela_wire_9741)
    );

    bfr new_Jinkela_buffer_7735 (
        .din(new_Jinkela_wire_9578),
        .dout(new_Jinkela_wire_9579)
    );

    bfr new_Jinkela_buffer_7760 (
        .din(new_Jinkela_wire_9613),
        .dout(new_Jinkela_wire_9614)
    );

    bfr new_Jinkela_buffer_7736 (
        .din(new_Jinkela_wire_9579),
        .dout(new_Jinkela_wire_9580)
    );

    bfr new_Jinkela_buffer_7841 (
        .din(new_Jinkela_wire_9696),
        .dout(new_Jinkela_wire_9697)
    );

    bfr new_Jinkela_buffer_7737 (
        .din(new_Jinkela_wire_9580),
        .dout(new_Jinkela_wire_9581)
    );

    bfr new_Jinkela_buffer_7761 (
        .din(new_Jinkela_wire_9614),
        .dout(new_Jinkela_wire_9615)
    );

    bfr new_Jinkela_buffer_7738 (
        .din(new_Jinkela_wire_9581),
        .dout(new_Jinkela_wire_9582)
    );

    spl2 new_Jinkela_splitter_780 (
        .a(_0205_),
        .b(new_Jinkela_wire_9742),
        .c(new_Jinkela_wire_9743)
    );

    bfr new_Jinkela_buffer_7739 (
        .din(new_Jinkela_wire_9582),
        .dout(new_Jinkela_wire_9583)
    );

    bfr new_Jinkela_buffer_7762 (
        .din(new_Jinkela_wire_9615),
        .dout(new_Jinkela_wire_9616)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_1370),
        .dout(new_Jinkela_wire_1371)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(_1592_),
        .b(new_Jinkela_wire_1594),
        .c(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_1414),
        .dout(new_Jinkela_wire_1415)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_1371),
        .dout(new_Jinkela_wire_1372)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_1372),
        .dout(new_Jinkela_wire_1373)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_1373),
        .dout(new_Jinkela_wire_1374)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_1374),
        .dout(new_Jinkela_wire_1375)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_1375),
        .dout(new_Jinkela_wire_1376)
    );

    bfr new_Jinkela_buffer_828 (
        .din(_0126_),
        .dout(new_Jinkela_wire_1588)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_1376),
        .dout(new_Jinkela_wire_1377)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_1378),
        .dout(new_Jinkela_wire_1379)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    bfr new_Jinkela_buffer_644 (
        .din(new_Jinkela_wire_1379),
        .dout(new_Jinkela_wire_1380)
    );

    spl2 new_Jinkela_splitter_230 (
        .a(_1065_),
        .b(new_Jinkela_wire_1592),
        .c(new_Jinkela_wire_1593)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1588),
        .dout(new_Jinkela_wire_1589)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_1383),
        .dout(new_Jinkela_wire_1384)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(new_Jinkela_wire_1384),
        .b(new_Jinkela_wire_1385),
        .c(new_Jinkela_wire_1386)
    );

    spl2 new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_1589),
        .b(new_Jinkela_wire_1590),
        .c(new_Jinkela_wire_1591)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_1422),
        .dout(new_Jinkela_wire_1423)
    );

    spl2 new_Jinkela_splitter_233 (
        .a(_0167_),
        .b(new_Jinkela_wire_1602),
        .c(new_Jinkela_wire_1603)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(_0365_),
        .b(new_Jinkela_wire_1596),
        .c(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(_0841_),
        .b(new_Jinkela_wire_1608),
        .c(new_Jinkela_wire_1609)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_1426),
        .dout(new_Jinkela_wire_1427)
    );

    bfr new_Jinkela_buffer_4255 (
        .din(new_Jinkela_wire_5578),
        .dout(new_Jinkela_wire_5579)
    );

    bfr new_Jinkela_buffer_4223 (
        .din(new_Jinkela_wire_5534),
        .dout(new_Jinkela_wire_5535)
    );

    bfr new_Jinkela_buffer_4224 (
        .din(new_Jinkela_wire_5535),
        .dout(new_Jinkela_wire_5536)
    );

    spl2 new_Jinkela_splitter_523 (
        .a(_1485_),
        .b(new_Jinkela_wire_5714),
        .c(new_Jinkela_wire_5715)
    );

    bfr new_Jinkela_buffer_4256 (
        .din(new_Jinkela_wire_5579),
        .dout(new_Jinkela_wire_5580)
    );

    bfr new_Jinkela_buffer_4356 (
        .din(new_Jinkela_wire_5699),
        .dout(new_Jinkela_wire_5700)
    );

    bfr new_Jinkela_buffer_4257 (
        .din(new_Jinkela_wire_5580),
        .dout(new_Jinkela_wire_5581)
    );

    bfr new_Jinkela_buffer_4357 (
        .din(new_Jinkela_wire_5700),
        .dout(new_Jinkela_wire_5701)
    );

    bfr new_Jinkela_buffer_4258 (
        .din(new_Jinkela_wire_5581),
        .dout(new_Jinkela_wire_5582)
    );

    bfr new_Jinkela_buffer_4361 (
        .din(new_Jinkela_wire_5704),
        .dout(new_Jinkela_wire_5705)
    );

    bfr new_Jinkela_buffer_4259 (
        .din(new_Jinkela_wire_5582),
        .dout(new_Jinkela_wire_5583)
    );

    bfr new_Jinkela_buffer_4358 (
        .din(new_Jinkela_wire_5701),
        .dout(new_Jinkela_wire_5702)
    );

    bfr new_Jinkela_buffer_4260 (
        .din(new_Jinkela_wire_5583),
        .dout(new_Jinkela_wire_5584)
    );

    spl2 new_Jinkela_splitter_524 (
        .a(_1023_),
        .b(new_Jinkela_wire_5716),
        .c(new_Jinkela_wire_5717)
    );

    bfr new_Jinkela_buffer_4261 (
        .din(new_Jinkela_wire_5584),
        .dout(new_Jinkela_wire_5585)
    );

    bfr new_Jinkela_buffer_4362 (
        .din(new_Jinkela_wire_5705),
        .dout(new_Jinkela_wire_5706)
    );

    bfr new_Jinkela_buffer_4262 (
        .din(new_Jinkela_wire_5585),
        .dout(new_Jinkela_wire_5586)
    );

    bfr new_Jinkela_buffer_4365 (
        .din(new_Jinkela_wire_5710),
        .dout(new_Jinkela_wire_5711)
    );

    bfr new_Jinkela_buffer_4263 (
        .din(new_Jinkela_wire_5586),
        .dout(new_Jinkela_wire_5587)
    );

    bfr new_Jinkela_buffer_4363 (
        .din(new_Jinkela_wire_5706),
        .dout(new_Jinkela_wire_5707)
    );

    bfr new_Jinkela_buffer_4264 (
        .din(new_Jinkela_wire_5587),
        .dout(new_Jinkela_wire_5588)
    );

    bfr new_Jinkela_buffer_4265 (
        .din(new_Jinkela_wire_5588),
        .dout(new_Jinkela_wire_5589)
    );

    spl2 new_Jinkela_splitter_521 (
        .a(new_Jinkela_wire_5707),
        .b(new_Jinkela_wire_5708),
        .c(new_Jinkela_wire_5709)
    );

    bfr new_Jinkela_buffer_4266 (
        .din(new_Jinkela_wire_5589),
        .dout(new_Jinkela_wire_5590)
    );

    bfr new_Jinkela_buffer_4366 (
        .din(_1146_),
        .dout(new_Jinkela_wire_5720)
    );

    bfr new_Jinkela_buffer_4267 (
        .din(new_Jinkela_wire_5590),
        .dout(new_Jinkela_wire_5591)
    );

    spl2 new_Jinkela_splitter_522 (
        .a(new_Jinkela_wire_5711),
        .b(new_Jinkela_wire_5712),
        .c(new_Jinkela_wire_5713)
    );

    bfr new_Jinkela_buffer_4268 (
        .din(new_Jinkela_wire_5591),
        .dout(new_Jinkela_wire_5592)
    );

    spl2 new_Jinkela_splitter_525 (
        .a(_0790_),
        .b(new_Jinkela_wire_5718),
        .c(new_Jinkela_wire_5719)
    );

    bfr new_Jinkela_buffer_4269 (
        .din(new_Jinkela_wire_5592),
        .dout(new_Jinkela_wire_5593)
    );

    spl2 new_Jinkela_splitter_527 (
        .a(_1437_),
        .b(new_Jinkela_wire_5723),
        .c(new_Jinkela_wire_5724)
    );

    spl2 new_Jinkela_splitter_526 (
        .a(_0728_),
        .b(new_Jinkela_wire_5721),
        .c(new_Jinkela_wire_5722)
    );

    bfr new_Jinkela_buffer_4270 (
        .din(new_Jinkela_wire_5593),
        .dout(new_Jinkela_wire_5594)
    );

    bfr new_Jinkela_buffer_4271 (
        .din(new_Jinkela_wire_5594),
        .dout(new_Jinkela_wire_5595)
    );

    spl2 new_Jinkela_splitter_528 (
        .a(_0927_),
        .b(new_Jinkela_wire_5725),
        .c(new_Jinkela_wire_5726)
    );

    bfr new_Jinkela_buffer_4272 (
        .din(new_Jinkela_wire_5595),
        .dout(new_Jinkela_wire_5596)
    );

    spl2 new_Jinkela_splitter_529 (
        .a(_1466_),
        .b(new_Jinkela_wire_5727),
        .c(new_Jinkela_wire_5728)
    );

    bfr new_Jinkela_buffer_4273 (
        .din(new_Jinkela_wire_5596),
        .dout(new_Jinkela_wire_5597)
    );

    bfr new_Jinkela_buffer_4368 (
        .din(_1330_),
        .dout(new_Jinkela_wire_5730)
    );

    bfr new_Jinkela_buffer_4367 (
        .din(_0122_),
        .dout(new_Jinkela_wire_5729)
    );

    bfr new_Jinkela_buffer_4274 (
        .din(new_Jinkela_wire_5597),
        .dout(new_Jinkela_wire_5598)
    );

    bfr new_Jinkela_buffer_11192 (
        .din(new_Jinkela_wire_13497),
        .dout(new_Jinkela_wire_13498)
    );

    bfr new_Jinkela_buffer_11359 (
        .din(_1377_),
        .dout(new_Jinkela_wire_13693)
    );

    bfr new_Jinkela_buffer_11193 (
        .din(new_Jinkela_wire_13498),
        .dout(new_Jinkela_wire_13499)
    );

    bfr new_Jinkela_buffer_11282 (
        .din(new_Jinkela_wire_13601),
        .dout(new_Jinkela_wire_13602)
    );

    bfr new_Jinkela_buffer_11194 (
        .din(new_Jinkela_wire_13499),
        .dout(new_Jinkela_wire_13500)
    );

    spl2 new_Jinkela_splitter_1017 (
        .a(_0308_),
        .b(new_Jinkela_wire_13720),
        .c(new_Jinkela_wire_13721)
    );

    bfr new_Jinkela_buffer_11195 (
        .din(new_Jinkela_wire_13500),
        .dout(new_Jinkela_wire_13501)
    );

    bfr new_Jinkela_buffer_11283 (
        .din(new_Jinkela_wire_13602),
        .dout(new_Jinkela_wire_13603)
    );

    bfr new_Jinkela_buffer_11196 (
        .din(new_Jinkela_wire_13501),
        .dout(new_Jinkela_wire_13502)
    );

    bfr new_Jinkela_buffer_11356 (
        .din(new_Jinkela_wire_13687),
        .dout(new_Jinkela_wire_13688)
    );

    bfr new_Jinkela_buffer_11197 (
        .din(new_Jinkela_wire_13502),
        .dout(new_Jinkela_wire_13503)
    );

    bfr new_Jinkela_buffer_11284 (
        .din(new_Jinkela_wire_13603),
        .dout(new_Jinkela_wire_13604)
    );

    bfr new_Jinkela_buffer_11198 (
        .din(new_Jinkela_wire_13503),
        .dout(new_Jinkela_wire_13504)
    );

    bfr new_Jinkela_buffer_11383 (
        .din(_1126_),
        .dout(new_Jinkela_wire_13719)
    );

    bfr new_Jinkela_buffer_11199 (
        .din(new_Jinkela_wire_13504),
        .dout(new_Jinkela_wire_13505)
    );

    bfr new_Jinkela_buffer_11285 (
        .din(new_Jinkela_wire_13604),
        .dout(new_Jinkela_wire_13605)
    );

    bfr new_Jinkela_buffer_11200 (
        .din(new_Jinkela_wire_13505),
        .dout(new_Jinkela_wire_13506)
    );

    bfr new_Jinkela_buffer_11357 (
        .din(new_Jinkela_wire_13688),
        .dout(new_Jinkela_wire_13689)
    );

    bfr new_Jinkela_buffer_11201 (
        .din(new_Jinkela_wire_13506),
        .dout(new_Jinkela_wire_13507)
    );

    bfr new_Jinkela_buffer_11286 (
        .din(new_Jinkela_wire_13605),
        .dout(new_Jinkela_wire_13606)
    );

    bfr new_Jinkela_buffer_11202 (
        .din(new_Jinkela_wire_13507),
        .dout(new_Jinkela_wire_13508)
    );

    bfr new_Jinkela_buffer_11360 (
        .din(new_Jinkela_wire_13693),
        .dout(new_Jinkela_wire_13694)
    );

    bfr new_Jinkela_buffer_11203 (
        .din(new_Jinkela_wire_13508),
        .dout(new_Jinkela_wire_13509)
    );

    bfr new_Jinkela_buffer_11287 (
        .din(new_Jinkela_wire_13606),
        .dout(new_Jinkela_wire_13607)
    );

    bfr new_Jinkela_buffer_11204 (
        .din(new_Jinkela_wire_13509),
        .dout(new_Jinkela_wire_13510)
    );

    bfr new_Jinkela_buffer_11358 (
        .din(new_Jinkela_wire_13689),
        .dout(new_Jinkela_wire_13690)
    );

    bfr new_Jinkela_buffer_11205 (
        .din(new_Jinkela_wire_13510),
        .dout(new_Jinkela_wire_13511)
    );

    bfr new_Jinkela_buffer_11288 (
        .din(new_Jinkela_wire_13607),
        .dout(new_Jinkela_wire_13608)
    );

    bfr new_Jinkela_buffer_11206 (
        .din(new_Jinkela_wire_13511),
        .dout(new_Jinkela_wire_13512)
    );

    spl2 new_Jinkela_splitter_1018 (
        .a(_0420_),
        .b(new_Jinkela_wire_13722),
        .c(new_Jinkela_wire_13723)
    );

    bfr new_Jinkela_buffer_11207 (
        .din(new_Jinkela_wire_13512),
        .dout(new_Jinkela_wire_13513)
    );

    bfr new_Jinkela_buffer_11289 (
        .din(new_Jinkela_wire_13608),
        .dout(new_Jinkela_wire_13609)
    );

    bfr new_Jinkela_buffer_11208 (
        .din(new_Jinkela_wire_13513),
        .dout(new_Jinkela_wire_13514)
    );

    bfr new_Jinkela_buffer_11361 (
        .din(new_Jinkela_wire_13694),
        .dout(new_Jinkela_wire_13695)
    );

    bfr new_Jinkela_buffer_11209 (
        .din(new_Jinkela_wire_13514),
        .dout(new_Jinkela_wire_13515)
    );

    bfr new_Jinkela_buffer_11290 (
        .din(new_Jinkela_wire_13609),
        .dout(new_Jinkela_wire_13610)
    );

    bfr new_Jinkela_buffer_11210 (
        .din(new_Jinkela_wire_13515),
        .dout(new_Jinkela_wire_13516)
    );

    spl2 new_Jinkela_splitter_1019 (
        .a(_0292_),
        .b(new_Jinkela_wire_13724),
        .c(new_Jinkela_wire_13725)
    );

    bfr new_Jinkela_buffer_11211 (
        .din(new_Jinkela_wire_13516),
        .dout(new_Jinkela_wire_13517)
    );

    bfr new_Jinkela_buffer_11291 (
        .din(new_Jinkela_wire_13610),
        .dout(new_Jinkela_wire_13611)
    );

    bfr new_Jinkela_buffer_11212 (
        .din(new_Jinkela_wire_13517),
        .dout(new_Jinkela_wire_13518)
    );

    bfr new_Jinkela_buffer_11362 (
        .din(new_Jinkela_wire_13695),
        .dout(new_Jinkela_wire_13696)
    );

    bfr new_Jinkela_buffer_14713 (
        .din(new_Jinkela_wire_17563),
        .dout(new_Jinkela_wire_17564)
    );

    bfr new_Jinkela_buffer_14627 (
        .din(new_Jinkela_wire_17457),
        .dout(new_Jinkela_wire_17458)
    );

    bfr new_Jinkela_buffer_14628 (
        .din(new_Jinkela_wire_17458),
        .dout(new_Jinkela_wire_17459)
    );

    bfr new_Jinkela_buffer_14714 (
        .din(new_Jinkela_wire_17564),
        .dout(new_Jinkela_wire_17565)
    );

    bfr new_Jinkela_buffer_14629 (
        .din(new_Jinkela_wire_17459),
        .dout(new_Jinkela_wire_17460)
    );

    bfr new_Jinkela_buffer_14787 (
        .din(new_Jinkela_wire_17641),
        .dout(new_Jinkela_wire_17642)
    );

    bfr new_Jinkela_buffer_14630 (
        .din(new_Jinkela_wire_17460),
        .dout(new_Jinkela_wire_17461)
    );

    bfr new_Jinkela_buffer_14715 (
        .din(new_Jinkela_wire_17565),
        .dout(new_Jinkela_wire_17566)
    );

    bfr new_Jinkela_buffer_14631 (
        .din(new_Jinkela_wire_17461),
        .dout(new_Jinkela_wire_17462)
    );

    spl2 new_Jinkela_splitter_1281 (
        .a(_0288_),
        .b(new_Jinkela_wire_17668),
        .c(new_Jinkela_wire_17669)
    );

    bfr new_Jinkela_buffer_14632 (
        .din(new_Jinkela_wire_17462),
        .dout(new_Jinkela_wire_17463)
    );

    bfr new_Jinkela_buffer_14716 (
        .din(new_Jinkela_wire_17566),
        .dout(new_Jinkela_wire_17567)
    );

    bfr new_Jinkela_buffer_14633 (
        .din(new_Jinkela_wire_17463),
        .dout(new_Jinkela_wire_17464)
    );

    bfr new_Jinkela_buffer_14788 (
        .din(new_Jinkela_wire_17642),
        .dout(new_Jinkela_wire_17643)
    );

    bfr new_Jinkela_buffer_14634 (
        .din(new_Jinkela_wire_17464),
        .dout(new_Jinkela_wire_17465)
    );

    bfr new_Jinkela_buffer_14717 (
        .din(new_Jinkela_wire_17567),
        .dout(new_Jinkela_wire_17568)
    );

    bfr new_Jinkela_buffer_14635 (
        .din(new_Jinkela_wire_17465),
        .dout(new_Jinkela_wire_17466)
    );

    bfr new_Jinkela_buffer_14799 (
        .din(new_Jinkela_wire_17663),
        .dout(new_Jinkela_wire_17664)
    );

    bfr new_Jinkela_buffer_14803 (
        .din(_0366_),
        .dout(new_Jinkela_wire_17670)
    );

    bfr new_Jinkela_buffer_14636 (
        .din(new_Jinkela_wire_17466),
        .dout(new_Jinkela_wire_17467)
    );

    bfr new_Jinkela_buffer_14718 (
        .din(new_Jinkela_wire_17568),
        .dout(new_Jinkela_wire_17569)
    );

    bfr new_Jinkela_buffer_14637 (
        .din(new_Jinkela_wire_17467),
        .dout(new_Jinkela_wire_17468)
    );

    bfr new_Jinkela_buffer_14789 (
        .din(new_Jinkela_wire_17643),
        .dout(new_Jinkela_wire_17644)
    );

    bfr new_Jinkela_buffer_14638 (
        .din(new_Jinkela_wire_17468),
        .dout(new_Jinkela_wire_17469)
    );

    bfr new_Jinkela_buffer_14719 (
        .din(new_Jinkela_wire_17569),
        .dout(new_Jinkela_wire_17570)
    );

    bfr new_Jinkela_buffer_14639 (
        .din(new_Jinkela_wire_17469),
        .dout(new_Jinkela_wire_17470)
    );

    spl2 new_Jinkela_splitter_1282 (
        .a(_1252_),
        .b(new_Jinkela_wire_17671),
        .c(new_Jinkela_wire_17672)
    );

    bfr new_Jinkela_buffer_14640 (
        .din(new_Jinkela_wire_17470),
        .dout(new_Jinkela_wire_17471)
    );

    bfr new_Jinkela_buffer_14720 (
        .din(new_Jinkela_wire_17570),
        .dout(new_Jinkela_wire_17571)
    );

    bfr new_Jinkela_buffer_14641 (
        .din(new_Jinkela_wire_17471),
        .dout(new_Jinkela_wire_17472)
    );

    bfr new_Jinkela_buffer_14790 (
        .din(new_Jinkela_wire_17644),
        .dout(new_Jinkela_wire_17645)
    );

    bfr new_Jinkela_buffer_14642 (
        .din(new_Jinkela_wire_17472),
        .dout(new_Jinkela_wire_17473)
    );

    bfr new_Jinkela_buffer_14721 (
        .din(new_Jinkela_wire_17571),
        .dout(new_Jinkela_wire_17572)
    );

    bfr new_Jinkela_buffer_14643 (
        .din(new_Jinkela_wire_17473),
        .dout(new_Jinkela_wire_17474)
    );

    bfr new_Jinkela_buffer_14800 (
        .din(new_Jinkela_wire_17664),
        .dout(new_Jinkela_wire_17665)
    );

    bfr new_Jinkela_buffer_14644 (
        .din(new_Jinkela_wire_17474),
        .dout(new_Jinkela_wire_17475)
    );

    bfr new_Jinkela_buffer_14722 (
        .din(new_Jinkela_wire_17572),
        .dout(new_Jinkela_wire_17573)
    );

    bfr new_Jinkela_buffer_14645 (
        .din(new_Jinkela_wire_17475),
        .dout(new_Jinkela_wire_17476)
    );

    bfr new_Jinkela_buffer_14791 (
        .din(new_Jinkela_wire_17645),
        .dout(new_Jinkela_wire_17646)
    );

    bfr new_Jinkela_buffer_14646 (
        .din(new_Jinkela_wire_17476),
        .dout(new_Jinkela_wire_17477)
    );

    bfr new_Jinkela_buffer_14723 (
        .din(new_Jinkela_wire_17573),
        .dout(new_Jinkela_wire_17574)
    );

    bfr new_Jinkela_buffer_14647 (
        .din(new_Jinkela_wire_17477),
        .dout(new_Jinkela_wire_17478)
    );

    bfr new_Jinkela_buffer_7740 (
        .din(new_Jinkela_wire_9583),
        .dout(new_Jinkela_wire_9584)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_7842 (
        .din(new_Jinkela_wire_9697),
        .dout(new_Jinkela_wire_9698)
    );

    spl2 new_Jinkela_splitter_235 (
        .a(_1105_),
        .b(new_Jinkela_wire_1614),
        .c(new_Jinkela_wire_1615)
    );

    bfr new_Jinkela_buffer_7741 (
        .din(new_Jinkela_wire_9584),
        .dout(new_Jinkela_wire_9585)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_1428),
        .dout(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_7763 (
        .din(new_Jinkela_wire_9616),
        .dout(new_Jinkela_wire_9617)
    );

    bfr new_Jinkela_buffer_7742 (
        .din(new_Jinkela_wire_9585),
        .dout(new_Jinkela_wire_9586)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_7743 (
        .din(new_Jinkela_wire_9586),
        .dout(new_Jinkela_wire_9587)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    bfr new_Jinkela_buffer_7764 (
        .din(new_Jinkela_wire_9617),
        .dout(new_Jinkela_wire_9618)
    );

    bfr new_Jinkela_buffer_7744 (
        .din(new_Jinkela_wire_9587),
        .dout(new_Jinkela_wire_9588)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_7843 (
        .din(new_Jinkela_wire_9698),
        .dout(new_Jinkela_wire_9699)
    );

    bfr new_Jinkela_buffer_7745 (
        .din(new_Jinkela_wire_9588),
        .dout(new_Jinkela_wire_9589)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1609),
        .dout(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_7765 (
        .din(new_Jinkela_wire_9618),
        .dout(new_Jinkela_wire_9619)
    );

    spl2 new_Jinkela_splitter_236 (
        .a(_0183_),
        .b(new_Jinkela_wire_1616),
        .c(new_Jinkela_wire_1617)
    );

    bfr new_Jinkela_buffer_7746 (
        .din(new_Jinkela_wire_9589),
        .dout(new_Jinkela_wire_9590)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_1605),
        .dout(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    spl2 new_Jinkela_splitter_781 (
        .a(_1056_),
        .b(new_Jinkela_wire_9744),
        .c(new_Jinkela_wire_9745)
    );

    bfr new_Jinkela_buffer_7747 (
        .din(new_Jinkela_wire_9590),
        .dout(new_Jinkela_wire_9591)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_7766 (
        .din(new_Jinkela_wire_9619),
        .dout(new_Jinkela_wire_9620)
    );

    bfr new_Jinkela_buffer_7748 (
        .din(new_Jinkela_wire_9591),
        .dout(new_Jinkela_wire_9592)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1606),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_1435),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_7844 (
        .din(new_Jinkela_wire_9699),
        .dout(new_Jinkela_wire_9700)
    );

    bfr new_Jinkela_buffer_7749 (
        .din(new_Jinkela_wire_9592),
        .dout(new_Jinkela_wire_9593)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_1610),
        .dout(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    bfr new_Jinkela_buffer_7767 (
        .din(new_Jinkela_wire_9620),
        .dout(new_Jinkela_wire_9621)
    );

    bfr new_Jinkela_buffer_7750 (
        .din(new_Jinkela_wire_9593),
        .dout(new_Jinkela_wire_9594)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_net_3970),
        .dout(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_7880 (
        .din(_0293_),
        .dout(new_Jinkela_wire_9746)
    );

    bfr new_Jinkela_buffer_842 (
        .din(_0512_),
        .dout(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_7751 (
        .din(new_Jinkela_wire_9594),
        .dout(new_Jinkela_wire_9595)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1611),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_1438),
        .dout(new_Jinkela_wire_1439)
    );

    bfr new_Jinkela_buffer_7768 (
        .din(new_Jinkela_wire_9621),
        .dout(new_Jinkela_wire_9622)
    );

    bfr new_Jinkela_buffer_7752 (
        .din(new_Jinkela_wire_9595),
        .dout(new_Jinkela_wire_9596)
    );

    spl2 new_Jinkela_splitter_238 (
        .a(_1299_),
        .b(new_Jinkela_wire_1621),
        .c(new_Jinkela_wire_1622)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_1439),
        .dout(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_7845 (
        .din(new_Jinkela_wire_9700),
        .dout(new_Jinkela_wire_9701)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(_0325_),
        .b(new_Jinkela_wire_1619),
        .c(new_Jinkela_wire_1620)
    );

    spl2 new_Jinkela_splitter_771 (
        .a(new_Jinkela_wire_9596),
        .b(new_Jinkela_wire_9597),
        .c(new_Jinkela_wire_9598)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_1440),
        .dout(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_7881 (
        .din(_0342_),
        .dout(new_Jinkela_wire_9749)
    );

    spl2 new_Jinkela_splitter_782 (
        .a(_1364_),
        .b(new_Jinkela_wire_9747),
        .c(new_Jinkela_wire_9748)
    );

    bfr new_Jinkela_buffer_7769 (
        .din(new_Jinkela_wire_9622),
        .dout(new_Jinkela_wire_9623)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_7770 (
        .din(new_Jinkela_wire_9623),
        .dout(new_Jinkela_wire_9624)
    );

    bfr new_Jinkela_buffer_7846 (
        .din(new_Jinkela_wire_9701),
        .dout(new_Jinkela_wire_9702)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_1442),
        .dout(new_Jinkela_wire_1443)
    );

    bfr new_Jinkela_buffer_7771 (
        .din(new_Jinkela_wire_9624),
        .dout(new_Jinkela_wire_9625)
    );

    bfr new_Jinkela_buffer_843 (
        .din(_1385_),
        .dout(new_Jinkela_wire_1623)
    );

    bfr new_Jinkela_buffer_7937 (
        .din(_1209_),
        .dout(new_Jinkela_wire_9809)
    );

    bfr new_Jinkela_buffer_844 (
        .din(_1749_),
        .dout(new_Jinkela_wire_1626)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_1443),
        .dout(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_7772 (
        .din(new_Jinkela_wire_9625),
        .dout(new_Jinkela_wire_9626)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(_0113_),
        .b(new_Jinkela_wire_1624),
        .c(new_Jinkela_wire_1625)
    );

    bfr new_Jinkela_buffer_7847 (
        .din(new_Jinkela_wire_9702),
        .dout(new_Jinkela_wire_9703)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_1444),
        .dout(new_Jinkela_wire_1445)
    );

    bfr new_Jinkela_buffer_7773 (
        .din(new_Jinkela_wire_9626),
        .dout(new_Jinkela_wire_9627)
    );

    spl2 new_Jinkela_splitter_784 (
        .a(_0605_),
        .b(new_Jinkela_wire_9807),
        .c(new_Jinkela_wire_9808)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_1445),
        .dout(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_7774 (
        .din(new_Jinkela_wire_9627),
        .dout(new_Jinkela_wire_9628)
    );

    bfr new_Jinkela_buffer_845 (
        .din(_0972_),
        .dout(new_Jinkela_wire_1627)
    );

    bfr new_Jinkela_buffer_7848 (
        .din(new_Jinkela_wire_9703),
        .dout(new_Jinkela_wire_9704)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_1446),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_7775 (
        .din(new_Jinkela_wire_9628),
        .dout(new_Jinkela_wire_9629)
    );

    bfr new_Jinkela_buffer_889 (
        .din(_1361_),
        .dout(new_Jinkela_wire_1673)
    );

    bfr new_Jinkela_buffer_7882 (
        .din(new_Jinkela_wire_9749),
        .dout(new_Jinkela_wire_9750)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1627),
        .dout(new_Jinkela_wire_1628)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_1447),
        .dout(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_7776 (
        .din(new_Jinkela_wire_9629),
        .dout(new_Jinkela_wire_9630)
    );

    spl2 new_Jinkela_splitter_1283 (
        .a(_0975_),
        .b(new_Jinkela_wire_17673),
        .c(new_Jinkela_wire_17674)
    );

    spl2 new_Jinkela_splitter_530 (
        .a(_1323_),
        .b(new_Jinkela_wire_5731),
        .c(new_Jinkela_wire_5732)
    );

    bfr new_Jinkela_buffer_14804 (
        .din(new_Jinkela_wire_17676),
        .dout(new_Jinkela_wire_17677)
    );

    bfr new_Jinkela_buffer_4275 (
        .din(new_Jinkela_wire_5598),
        .dout(new_Jinkela_wire_5599)
    );

    bfr new_Jinkela_buffer_14648 (
        .din(new_Jinkela_wire_17478),
        .dout(new_Jinkela_wire_17479)
    );

    spl2 new_Jinkela_splitter_531 (
        .a(_1518_),
        .b(new_Jinkela_wire_5733),
        .c(new_Jinkela_wire_5734)
    );

    bfr new_Jinkela_buffer_14724 (
        .din(new_Jinkela_wire_17574),
        .dout(new_Jinkela_wire_17575)
    );

    bfr new_Jinkela_buffer_4276 (
        .din(new_Jinkela_wire_5599),
        .dout(new_Jinkela_wire_5600)
    );

    bfr new_Jinkela_buffer_14649 (
        .din(new_Jinkela_wire_17479),
        .dout(new_Jinkela_wire_17480)
    );

    bfr new_Jinkela_buffer_14792 (
        .din(new_Jinkela_wire_17646),
        .dout(new_Jinkela_wire_17647)
    );

    bfr new_Jinkela_buffer_4277 (
        .din(new_Jinkela_wire_5600),
        .dout(new_Jinkela_wire_5601)
    );

    bfr new_Jinkela_buffer_14650 (
        .din(new_Jinkela_wire_17480),
        .dout(new_Jinkela_wire_17481)
    );

    bfr new_Jinkela_buffer_14725 (
        .din(new_Jinkela_wire_17575),
        .dout(new_Jinkela_wire_17576)
    );

    spl2 new_Jinkela_splitter_532 (
        .a(_1062_),
        .b(new_Jinkela_wire_5735),
        .c(new_Jinkela_wire_5736)
    );

    bfr new_Jinkela_buffer_4278 (
        .din(new_Jinkela_wire_5601),
        .dout(new_Jinkela_wire_5602)
    );

    bfr new_Jinkela_buffer_14651 (
        .din(new_Jinkela_wire_17481),
        .dout(new_Jinkela_wire_17482)
    );

    bfr new_Jinkela_buffer_14801 (
        .din(new_Jinkela_wire_17665),
        .dout(new_Jinkela_wire_17666)
    );

    spl2 new_Jinkela_splitter_533 (
        .a(_1665_),
        .b(new_Jinkela_wire_5737),
        .c(new_Jinkela_wire_5738)
    );

    bfr new_Jinkela_buffer_4279 (
        .din(new_Jinkela_wire_5602),
        .dout(new_Jinkela_wire_5603)
    );

    bfr new_Jinkela_buffer_14652 (
        .din(new_Jinkela_wire_17482),
        .dout(new_Jinkela_wire_17483)
    );

    bfr new_Jinkela_buffer_14726 (
        .din(new_Jinkela_wire_17576),
        .dout(new_Jinkela_wire_17577)
    );

    bfr new_Jinkela_buffer_4369 (
        .din(_0280_),
        .dout(new_Jinkela_wire_5739)
    );

    bfr new_Jinkela_buffer_4280 (
        .din(new_Jinkela_wire_5603),
        .dout(new_Jinkela_wire_5604)
    );

    bfr new_Jinkela_buffer_14653 (
        .din(new_Jinkela_wire_17483),
        .dout(new_Jinkela_wire_17484)
    );

    bfr new_Jinkela_buffer_4370 (
        .din(_1463_),
        .dout(new_Jinkela_wire_5742)
    );

    bfr new_Jinkela_buffer_14793 (
        .din(new_Jinkela_wire_17647),
        .dout(new_Jinkela_wire_17648)
    );

    spl2 new_Jinkela_splitter_534 (
        .a(_1547_),
        .b(new_Jinkela_wire_5740),
        .c(new_Jinkela_wire_5741)
    );

    bfr new_Jinkela_buffer_4281 (
        .din(new_Jinkela_wire_5604),
        .dout(new_Jinkela_wire_5605)
    );

    bfr new_Jinkela_buffer_14654 (
        .din(new_Jinkela_wire_17484),
        .dout(new_Jinkela_wire_17485)
    );

    bfr new_Jinkela_buffer_4426 (
        .din(_0502_),
        .dout(new_Jinkela_wire_5802)
    );

    bfr new_Jinkela_buffer_14727 (
        .din(new_Jinkela_wire_17577),
        .dout(new_Jinkela_wire_17578)
    );

    bfr new_Jinkela_buffer_4282 (
        .din(new_Jinkela_wire_5605),
        .dout(new_Jinkela_wire_5606)
    );

    bfr new_Jinkela_buffer_14655 (
        .din(new_Jinkela_wire_17485),
        .dout(new_Jinkela_wire_17486)
    );

    spl2 new_Jinkela_splitter_536 (
        .a(_1705_),
        .b(new_Jinkela_wire_5800),
        .c(new_Jinkela_wire_5801)
    );

    bfr new_Jinkela_buffer_4283 (
        .din(new_Jinkela_wire_5606),
        .dout(new_Jinkela_wire_5607)
    );

    bfr new_Jinkela_buffer_14656 (
        .din(new_Jinkela_wire_17486),
        .dout(new_Jinkela_wire_17487)
    );

    bfr new_Jinkela_buffer_4371 (
        .din(new_Jinkela_wire_5742),
        .dout(new_Jinkela_wire_5743)
    );

    bfr new_Jinkela_buffer_14728 (
        .din(new_Jinkela_wire_17578),
        .dout(new_Jinkela_wire_17579)
    );

    bfr new_Jinkela_buffer_4284 (
        .din(new_Jinkela_wire_5607),
        .dout(new_Jinkela_wire_5608)
    );

    bfr new_Jinkela_buffer_14657 (
        .din(new_Jinkela_wire_17487),
        .dout(new_Jinkela_wire_17488)
    );

    spl2 new_Jinkela_splitter_537 (
        .a(_0117_),
        .b(new_Jinkela_wire_5804),
        .c(new_Jinkela_wire_5805)
    );

    bfr new_Jinkela_buffer_14794 (
        .din(new_Jinkela_wire_17648),
        .dout(new_Jinkela_wire_17649)
    );

    bfr new_Jinkela_buffer_4285 (
        .din(new_Jinkela_wire_5608),
        .dout(new_Jinkela_wire_5609)
    );

    bfr new_Jinkela_buffer_14658 (
        .din(new_Jinkela_wire_17488),
        .dout(new_Jinkela_wire_17489)
    );

    bfr new_Jinkela_buffer_4372 (
        .din(new_Jinkela_wire_5743),
        .dout(new_Jinkela_wire_5744)
    );

    bfr new_Jinkela_buffer_14729 (
        .din(new_Jinkela_wire_17579),
        .dout(new_Jinkela_wire_17580)
    );

    bfr new_Jinkela_buffer_4286 (
        .din(new_Jinkela_wire_5609),
        .dout(new_Jinkela_wire_5610)
    );

    bfr new_Jinkela_buffer_14659 (
        .din(new_Jinkela_wire_17489),
        .dout(new_Jinkela_wire_17490)
    );

    bfr new_Jinkela_buffer_14802 (
        .din(new_Jinkela_wire_17666),
        .dout(new_Jinkela_wire_17667)
    );

    bfr new_Jinkela_buffer_4427 (
        .din(_0551_),
        .dout(new_Jinkela_wire_5803)
    );

    bfr new_Jinkela_buffer_4287 (
        .din(new_Jinkela_wire_5610),
        .dout(new_Jinkela_wire_5611)
    );

    bfr new_Jinkela_buffer_14660 (
        .din(new_Jinkela_wire_17490),
        .dout(new_Jinkela_wire_17491)
    );

    bfr new_Jinkela_buffer_4373 (
        .din(new_Jinkela_wire_5744),
        .dout(new_Jinkela_wire_5745)
    );

    bfr new_Jinkela_buffer_14730 (
        .din(new_Jinkela_wire_17580),
        .dout(new_Jinkela_wire_17581)
    );

    bfr new_Jinkela_buffer_4288 (
        .din(new_Jinkela_wire_5611),
        .dout(new_Jinkela_wire_5612)
    );

    bfr new_Jinkela_buffer_14661 (
        .din(new_Jinkela_wire_17491),
        .dout(new_Jinkela_wire_17492)
    );

    spl2 new_Jinkela_splitter_538 (
        .a(_0352_),
        .b(new_Jinkela_wire_5806),
        .c(new_Jinkela_wire_5807)
    );

    bfr new_Jinkela_buffer_14795 (
        .din(new_Jinkela_wire_17649),
        .dout(new_Jinkela_wire_17650)
    );

    bfr new_Jinkela_buffer_4289 (
        .din(new_Jinkela_wire_5612),
        .dout(new_Jinkela_wire_5613)
    );

    bfr new_Jinkela_buffer_14662 (
        .din(new_Jinkela_wire_17492),
        .dout(new_Jinkela_wire_17493)
    );

    bfr new_Jinkela_buffer_4374 (
        .din(new_Jinkela_wire_5745),
        .dout(new_Jinkela_wire_5746)
    );

    bfr new_Jinkela_buffer_14731 (
        .din(new_Jinkela_wire_17581),
        .dout(new_Jinkela_wire_17582)
    );

    bfr new_Jinkela_buffer_4290 (
        .din(new_Jinkela_wire_5613),
        .dout(new_Jinkela_wire_5614)
    );

    bfr new_Jinkela_buffer_14663 (
        .din(new_Jinkela_wire_17493),
        .dout(new_Jinkela_wire_17494)
    );

    spl2 new_Jinkela_splitter_1284 (
        .a(_1771_),
        .b(new_Jinkela_wire_17675),
        .c(new_Jinkela_wire_17676)
    );

    bfr new_Jinkela_buffer_4291 (
        .din(new_Jinkela_wire_5614),
        .dout(new_Jinkela_wire_5615)
    );

    bfr new_Jinkela_buffer_14664 (
        .din(new_Jinkela_wire_17494),
        .dout(new_Jinkela_wire_17495)
    );

    bfr new_Jinkela_buffer_4375 (
        .din(new_Jinkela_wire_5746),
        .dout(new_Jinkela_wire_5747)
    );

    bfr new_Jinkela_buffer_14732 (
        .din(new_Jinkela_wire_17582),
        .dout(new_Jinkela_wire_17583)
    );

    bfr new_Jinkela_buffer_4292 (
        .din(new_Jinkela_wire_5615),
        .dout(new_Jinkela_wire_5616)
    );

    bfr new_Jinkela_buffer_14665 (
        .din(new_Jinkela_wire_17495),
        .dout(new_Jinkela_wire_17496)
    );

    bfr new_Jinkela_buffer_14796 (
        .din(new_Jinkela_wire_17650),
        .dout(new_Jinkela_wire_17651)
    );

    spl2 new_Jinkela_splitter_539 (
        .a(_1602_),
        .b(new_Jinkela_wire_5812),
        .c(new_Jinkela_wire_5813)
    );

    bfr new_Jinkela_buffer_4293 (
        .din(new_Jinkela_wire_5616),
        .dout(new_Jinkela_wire_5617)
    );

    bfr new_Jinkela_buffer_14666 (
        .din(new_Jinkela_wire_17496),
        .dout(new_Jinkela_wire_17497)
    );

    bfr new_Jinkela_buffer_4376 (
        .din(new_Jinkela_wire_5747),
        .dout(new_Jinkela_wire_5748)
    );

    bfr new_Jinkela_buffer_14733 (
        .din(new_Jinkela_wire_17583),
        .dout(new_Jinkela_wire_17584)
    );

    bfr new_Jinkela_buffer_4294 (
        .din(new_Jinkela_wire_5617),
        .dout(new_Jinkela_wire_5618)
    );

    bfr new_Jinkela_buffer_14667 (
        .din(new_Jinkela_wire_17497),
        .dout(new_Jinkela_wire_17498)
    );

    bfr new_Jinkela_buffer_4428 (
        .din(new_Jinkela_wire_5807),
        .dout(new_Jinkela_wire_5808)
    );

    bfr new_Jinkela_buffer_4432 (
        .din(_0542_),
        .dout(new_Jinkela_wire_5814)
    );

    spl2 new_Jinkela_splitter_1285 (
        .a(_1331_),
        .b(new_Jinkela_wire_17681),
        .c(new_Jinkela_wire_17682)
    );

    bfr new_Jinkela_buffer_4295 (
        .din(new_Jinkela_wire_5618),
        .dout(new_Jinkela_wire_5619)
    );

    bfr new_Jinkela_buffer_14668 (
        .din(new_Jinkela_wire_17498),
        .dout(new_Jinkela_wire_17499)
    );

    bfr new_Jinkela_buffer_11213 (
        .din(new_Jinkela_wire_13518),
        .dout(new_Jinkela_wire_13519)
    );

    bfr new_Jinkela_buffer_11292 (
        .din(new_Jinkela_wire_13611),
        .dout(new_Jinkela_wire_13612)
    );

    bfr new_Jinkela_buffer_11214 (
        .din(new_Jinkela_wire_13519),
        .dout(new_Jinkela_wire_13520)
    );

    bfr new_Jinkela_buffer_11215 (
        .din(new_Jinkela_wire_13520),
        .dout(new_Jinkela_wire_13521)
    );

    bfr new_Jinkela_buffer_11293 (
        .din(new_Jinkela_wire_13612),
        .dout(new_Jinkela_wire_13613)
    );

    bfr new_Jinkela_buffer_11216 (
        .din(new_Jinkela_wire_13521),
        .dout(new_Jinkela_wire_13522)
    );

    bfr new_Jinkela_buffer_11363 (
        .din(new_Jinkela_wire_13696),
        .dout(new_Jinkela_wire_13697)
    );

    bfr new_Jinkela_buffer_11217 (
        .din(new_Jinkela_wire_13522),
        .dout(new_Jinkela_wire_13523)
    );

    bfr new_Jinkela_buffer_11294 (
        .din(new_Jinkela_wire_13613),
        .dout(new_Jinkela_wire_13614)
    );

    bfr new_Jinkela_buffer_11218 (
        .din(new_Jinkela_wire_13523),
        .dout(new_Jinkela_wire_13524)
    );

    spl2 new_Jinkela_splitter_1020 (
        .a(_1426_),
        .b(new_Jinkela_wire_13730),
        .c(new_Jinkela_wire_13731)
    );

    bfr new_Jinkela_buffer_11219 (
        .din(new_Jinkela_wire_13524),
        .dout(new_Jinkela_wire_13525)
    );

    bfr new_Jinkela_buffer_11295 (
        .din(new_Jinkela_wire_13614),
        .dout(new_Jinkela_wire_13615)
    );

    bfr new_Jinkela_buffer_11220 (
        .din(new_Jinkela_wire_13525),
        .dout(new_Jinkela_wire_13526)
    );

    bfr new_Jinkela_buffer_11364 (
        .din(new_Jinkela_wire_13697),
        .dout(new_Jinkela_wire_13698)
    );

    bfr new_Jinkela_buffer_11221 (
        .din(new_Jinkela_wire_13526),
        .dout(new_Jinkela_wire_13527)
    );

    bfr new_Jinkela_buffer_11296 (
        .din(new_Jinkela_wire_13615),
        .dout(new_Jinkela_wire_13616)
    );

    bfr new_Jinkela_buffer_11222 (
        .din(new_Jinkela_wire_13527),
        .dout(new_Jinkela_wire_13528)
    );

    bfr new_Jinkela_buffer_11384 (
        .din(new_Jinkela_wire_13725),
        .dout(new_Jinkela_wire_13726)
    );

    bfr new_Jinkela_buffer_11388 (
        .din(_0079_),
        .dout(new_Jinkela_wire_13732)
    );

    bfr new_Jinkela_buffer_11223 (
        .din(new_Jinkela_wire_13528),
        .dout(new_Jinkela_wire_13529)
    );

    bfr new_Jinkela_buffer_11297 (
        .din(new_Jinkela_wire_13616),
        .dout(new_Jinkela_wire_13617)
    );

    bfr new_Jinkela_buffer_11224 (
        .din(new_Jinkela_wire_13529),
        .dout(new_Jinkela_wire_13530)
    );

    bfr new_Jinkela_buffer_11365 (
        .din(new_Jinkela_wire_13698),
        .dout(new_Jinkela_wire_13699)
    );

    bfr new_Jinkela_buffer_11225 (
        .din(new_Jinkela_wire_13530),
        .dout(new_Jinkela_wire_13531)
    );

    bfr new_Jinkela_buffer_11298 (
        .din(new_Jinkela_wire_13617),
        .dout(new_Jinkela_wire_13618)
    );

    bfr new_Jinkela_buffer_11226 (
        .din(new_Jinkela_wire_13531),
        .dout(new_Jinkela_wire_13532)
    );

    spl2 new_Jinkela_splitter_1022 (
        .a(_1770_),
        .b(new_Jinkela_wire_13846),
        .c(new_Jinkela_wire_13847)
    );

    bfr new_Jinkela_buffer_11227 (
        .din(new_Jinkela_wire_13532),
        .dout(new_Jinkela_wire_13533)
    );

    bfr new_Jinkela_buffer_11299 (
        .din(new_Jinkela_wire_13618),
        .dout(new_Jinkela_wire_13619)
    );

    bfr new_Jinkela_buffer_11228 (
        .din(new_Jinkela_wire_13533),
        .dout(new_Jinkela_wire_13534)
    );

    bfr new_Jinkela_buffer_11366 (
        .din(new_Jinkela_wire_13699),
        .dout(new_Jinkela_wire_13700)
    );

    bfr new_Jinkela_buffer_11229 (
        .din(new_Jinkela_wire_13534),
        .dout(new_Jinkela_wire_13535)
    );

    bfr new_Jinkela_buffer_11300 (
        .din(new_Jinkela_wire_13619),
        .dout(new_Jinkela_wire_13620)
    );

    bfr new_Jinkela_buffer_11230 (
        .din(new_Jinkela_wire_13535),
        .dout(new_Jinkela_wire_13536)
    );

    bfr new_Jinkela_buffer_11385 (
        .din(new_Jinkela_wire_13726),
        .dout(new_Jinkela_wire_13727)
    );

    bfr new_Jinkela_buffer_11231 (
        .din(new_Jinkela_wire_13536),
        .dout(new_Jinkela_wire_13537)
    );

    bfr new_Jinkela_buffer_11301 (
        .din(new_Jinkela_wire_13620),
        .dout(new_Jinkela_wire_13621)
    );

    bfr new_Jinkela_buffer_11232 (
        .din(new_Jinkela_wire_13537),
        .dout(new_Jinkela_wire_13538)
    );

    bfr new_Jinkela_buffer_11367 (
        .din(new_Jinkela_wire_13700),
        .dout(new_Jinkela_wire_13701)
    );

    bfr new_Jinkela_buffer_11233 (
        .din(new_Jinkela_wire_13538),
        .dout(new_Jinkela_wire_13539)
    );

    bfr new_Jinkela_buffer_11302 (
        .din(new_Jinkela_wire_13621),
        .dout(new_Jinkela_wire_13622)
    );

    spl2 new_Jinkela_splitter_242 (
        .a(_0431_),
        .b(new_Jinkela_wire_1763),
        .c(new_Jinkela_wire_1764)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_1448),
        .dout(new_Jinkela_wire_1449)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1628),
        .dout(new_Jinkela_wire_1629)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_1449),
        .dout(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_1450),
        .dout(new_Jinkela_wire_1451)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1629),
        .dout(new_Jinkela_wire_1630)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_1451),
        .dout(new_Jinkela_wire_1452)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_1452),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(new_Jinkela_wire_1630),
        .b(new_Jinkela_wire_1631),
        .c(new_Jinkela_wire_1632)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_1453),
        .dout(new_Jinkela_wire_1454)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1673),
        .dout(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1635),
        .dout(new_Jinkela_wire_1636)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    spl2 new_Jinkela_splitter_243 (
        .a(_1405_),
        .b(new_Jinkela_wire_1765),
        .c(new_Jinkela_wire_1766)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1636),
        .dout(new_Jinkela_wire_1637)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1674),
        .dout(new_Jinkela_wire_1675)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1637),
        .dout(new_Jinkela_wire_1638)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1638),
        .dout(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(_0883_),
        .b(new_Jinkela_wire_1771),
        .c(new_Jinkela_wire_1772)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1675),
        .dout(new_Jinkela_wire_1676)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1639),
        .dout(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1766),
        .dout(new_Jinkela_wire_1767)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_1465),
        .dout(new_Jinkela_wire_1466)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1640),
        .dout(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_1466),
        .dout(new_Jinkela_wire_1467)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(_0633_),
        .b(new_Jinkela_wire_1773),
        .c(new_Jinkela_wire_1774)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1676),
        .dout(new_Jinkela_wire_1677)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_1467),
        .dout(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1641),
        .dout(new_Jinkela_wire_1642)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_1468),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_14734 (
        .din(new_Jinkela_wire_17584),
        .dout(new_Jinkela_wire_17585)
    );

    bfr new_Jinkela_buffer_14669 (
        .din(new_Jinkela_wire_17499),
        .dout(new_Jinkela_wire_17500)
    );

    bfr new_Jinkela_buffer_14797 (
        .din(new_Jinkela_wire_17651),
        .dout(new_Jinkela_wire_17652)
    );

    bfr new_Jinkela_buffer_14670 (
        .din(new_Jinkela_wire_17500),
        .dout(new_Jinkela_wire_17501)
    );

    bfr new_Jinkela_buffer_14735 (
        .din(new_Jinkela_wire_17585),
        .dout(new_Jinkela_wire_17586)
    );

    bfr new_Jinkela_buffer_14671 (
        .din(new_Jinkela_wire_17501),
        .dout(new_Jinkela_wire_17502)
    );

    bfr new_Jinkela_buffer_14808 (
        .din(_0006_),
        .dout(new_Jinkela_wire_17683)
    );

    bfr new_Jinkela_buffer_14672 (
        .din(new_Jinkela_wire_17502),
        .dout(new_Jinkela_wire_17503)
    );

    bfr new_Jinkela_buffer_14736 (
        .din(new_Jinkela_wire_17586),
        .dout(new_Jinkela_wire_17587)
    );

    bfr new_Jinkela_buffer_14673 (
        .din(new_Jinkela_wire_17503),
        .dout(new_Jinkela_wire_17504)
    );

    bfr new_Jinkela_buffer_14798 (
        .din(new_Jinkela_wire_17652),
        .dout(new_Jinkela_wire_17653)
    );

    bfr new_Jinkela_buffer_14674 (
        .din(new_Jinkela_wire_17504),
        .dout(new_Jinkela_wire_17505)
    );

    bfr new_Jinkela_buffer_14737 (
        .din(new_Jinkela_wire_17587),
        .dout(new_Jinkela_wire_17588)
    );

    bfr new_Jinkela_buffer_14675 (
        .din(new_Jinkela_wire_17505),
        .dout(new_Jinkela_wire_17506)
    );

    bfr new_Jinkela_buffer_14676 (
        .din(new_Jinkela_wire_17506),
        .dout(new_Jinkela_wire_17507)
    );

    bfr new_Jinkela_buffer_14738 (
        .din(new_Jinkela_wire_17588),
        .dout(new_Jinkela_wire_17589)
    );

    bfr new_Jinkela_buffer_14677 (
        .din(new_Jinkela_wire_17507),
        .dout(new_Jinkela_wire_17508)
    );

    spl2 new_Jinkela_splitter_1276 (
        .a(new_Jinkela_wire_17653),
        .b(new_Jinkela_wire_17654),
        .c(new_Jinkela_wire_17655)
    );

    bfr new_Jinkela_buffer_14678 (
        .din(new_Jinkela_wire_17508),
        .dout(new_Jinkela_wire_17509)
    );

    bfr new_Jinkela_buffer_14739 (
        .din(new_Jinkela_wire_17589),
        .dout(new_Jinkela_wire_17590)
    );

    bfr new_Jinkela_buffer_14679 (
        .din(new_Jinkela_wire_17509),
        .dout(new_Jinkela_wire_17510)
    );

    bfr new_Jinkela_buffer_14849 (
        .din(_1284_),
        .dout(new_Jinkela_wire_17726)
    );

    bfr new_Jinkela_buffer_14809 (
        .din(_1373_),
        .dout(new_Jinkela_wire_17684)
    );

    bfr new_Jinkela_buffer_14680 (
        .din(new_Jinkela_wire_17510),
        .dout(new_Jinkela_wire_17511)
    );

    bfr new_Jinkela_buffer_14740 (
        .din(new_Jinkela_wire_17590),
        .dout(new_Jinkela_wire_17591)
    );

    bfr new_Jinkela_buffer_14681 (
        .din(new_Jinkela_wire_17511),
        .dout(new_Jinkela_wire_17512)
    );

    bfr new_Jinkela_buffer_14805 (
        .din(new_Jinkela_wire_17677),
        .dout(new_Jinkela_wire_17678)
    );

    bfr new_Jinkela_buffer_14682 (
        .din(new_Jinkela_wire_17512),
        .dout(new_Jinkela_wire_17513)
    );

    bfr new_Jinkela_buffer_14741 (
        .din(new_Jinkela_wire_17591),
        .dout(new_Jinkela_wire_17592)
    );

    bfr new_Jinkela_buffer_14683 (
        .din(new_Jinkela_wire_17513),
        .dout(new_Jinkela_wire_17514)
    );

    bfr new_Jinkela_buffer_14806 (
        .din(new_Jinkela_wire_17678),
        .dout(new_Jinkela_wire_17679)
    );

    bfr new_Jinkela_buffer_14684 (
        .din(new_Jinkela_wire_17514),
        .dout(new_Jinkela_wire_17515)
    );

    bfr new_Jinkela_buffer_14742 (
        .din(new_Jinkela_wire_17592),
        .dout(new_Jinkela_wire_17593)
    );

    bfr new_Jinkela_buffer_14685 (
        .din(new_Jinkela_wire_17515),
        .dout(new_Jinkela_wire_17516)
    );

    bfr new_Jinkela_buffer_14905 (
        .din(_1717_),
        .dout(new_Jinkela_wire_17784)
    );

    bfr new_Jinkela_buffer_14686 (
        .din(new_Jinkela_wire_17516),
        .dout(new_Jinkela_wire_17517)
    );

    bfr new_Jinkela_buffer_14743 (
        .din(new_Jinkela_wire_17593),
        .dout(new_Jinkela_wire_17594)
    );

    bfr new_Jinkela_buffer_14687 (
        .din(new_Jinkela_wire_17517),
        .dout(new_Jinkela_wire_17518)
    );

    bfr new_Jinkela_buffer_14807 (
        .din(new_Jinkela_wire_17679),
        .dout(new_Jinkela_wire_17680)
    );

    bfr new_Jinkela_buffer_14688 (
        .din(new_Jinkela_wire_17518),
        .dout(new_Jinkela_wire_17519)
    );

    bfr new_Jinkela_buffer_14744 (
        .din(new_Jinkela_wire_17594),
        .dout(new_Jinkela_wire_17595)
    );

    bfr new_Jinkela_buffer_14689 (
        .din(new_Jinkela_wire_17519),
        .dout(new_Jinkela_wire_17520)
    );

    bfr new_Jinkela_buffer_4377 (
        .din(new_Jinkela_wire_5748),
        .dout(new_Jinkela_wire_5749)
    );

    bfr new_Jinkela_buffer_4296 (
        .din(new_Jinkela_wire_5619),
        .dout(new_Jinkela_wire_5620)
    );

    spl2 new_Jinkela_splitter_542 (
        .a(_0370_),
        .b(new_Jinkela_wire_5882),
        .c(new_Jinkela_wire_5883)
    );

    bfr new_Jinkela_buffer_4297 (
        .din(new_Jinkela_wire_5620),
        .dout(new_Jinkela_wire_5621)
    );

    bfr new_Jinkela_buffer_4378 (
        .din(new_Jinkela_wire_5749),
        .dout(new_Jinkela_wire_5750)
    );

    bfr new_Jinkela_buffer_4298 (
        .din(new_Jinkela_wire_5621),
        .dout(new_Jinkela_wire_5622)
    );

    bfr new_Jinkela_buffer_4429 (
        .din(new_Jinkela_wire_5808),
        .dout(new_Jinkela_wire_5809)
    );

    bfr new_Jinkela_buffer_4299 (
        .din(new_Jinkela_wire_5622),
        .dout(new_Jinkela_wire_5623)
    );

    bfr new_Jinkela_buffer_4379 (
        .din(new_Jinkela_wire_5750),
        .dout(new_Jinkela_wire_5751)
    );

    bfr new_Jinkela_buffer_4300 (
        .din(new_Jinkela_wire_5623),
        .dout(new_Jinkela_wire_5624)
    );

    spl2 new_Jinkela_splitter_541 (
        .a(_1242_),
        .b(new_Jinkela_wire_5880),
        .c(new_Jinkela_wire_5881)
    );

    bfr new_Jinkela_buffer_4301 (
        .din(new_Jinkela_wire_5624),
        .dout(new_Jinkela_wire_5625)
    );

    bfr new_Jinkela_buffer_4380 (
        .din(new_Jinkela_wire_5751),
        .dout(new_Jinkela_wire_5752)
    );

    bfr new_Jinkela_buffer_4302 (
        .din(new_Jinkela_wire_5625),
        .dout(new_Jinkela_wire_5626)
    );

    bfr new_Jinkela_buffer_4430 (
        .din(new_Jinkela_wire_5809),
        .dout(new_Jinkela_wire_5810)
    );

    bfr new_Jinkela_buffer_4303 (
        .din(new_Jinkela_wire_5626),
        .dout(new_Jinkela_wire_5627)
    );

    bfr new_Jinkela_buffer_4381 (
        .din(new_Jinkela_wire_5752),
        .dout(new_Jinkela_wire_5753)
    );

    bfr new_Jinkela_buffer_4304 (
        .din(new_Jinkela_wire_5627),
        .dout(new_Jinkela_wire_5628)
    );

    bfr new_Jinkela_buffer_4433 (
        .din(new_Jinkela_wire_5814),
        .dout(new_Jinkela_wire_5815)
    );

    bfr new_Jinkela_buffer_4305 (
        .din(new_Jinkela_wire_5628),
        .dout(new_Jinkela_wire_5629)
    );

    bfr new_Jinkela_buffer_4382 (
        .din(new_Jinkela_wire_5753),
        .dout(new_Jinkela_wire_5754)
    );

    bfr new_Jinkela_buffer_4306 (
        .din(new_Jinkela_wire_5629),
        .dout(new_Jinkela_wire_5630)
    );

    bfr new_Jinkela_buffer_4431 (
        .din(new_Jinkela_wire_5810),
        .dout(new_Jinkela_wire_5811)
    );

    bfr new_Jinkela_buffer_4307 (
        .din(new_Jinkela_wire_5630),
        .dout(new_Jinkela_wire_5631)
    );

    bfr new_Jinkela_buffer_4383 (
        .din(new_Jinkela_wire_5754),
        .dout(new_Jinkela_wire_5755)
    );

    bfr new_Jinkela_buffer_4308 (
        .din(new_Jinkela_wire_5631),
        .dout(new_Jinkela_wire_5632)
    );

    bfr new_Jinkela_buffer_4309 (
        .din(new_Jinkela_wire_5632),
        .dout(new_Jinkela_wire_5633)
    );

    bfr new_Jinkela_buffer_4384 (
        .din(new_Jinkela_wire_5755),
        .dout(new_Jinkela_wire_5756)
    );

    bfr new_Jinkela_buffer_4310 (
        .din(new_Jinkela_wire_5633),
        .dout(new_Jinkela_wire_5634)
    );

    bfr new_Jinkela_buffer_4434 (
        .din(new_Jinkela_wire_5815),
        .dout(new_Jinkela_wire_5816)
    );

    bfr new_Jinkela_buffer_4311 (
        .din(new_Jinkela_wire_5634),
        .dout(new_Jinkela_wire_5635)
    );

    bfr new_Jinkela_buffer_4385 (
        .din(new_Jinkela_wire_5756),
        .dout(new_Jinkela_wire_5757)
    );

    bfr new_Jinkela_buffer_4312 (
        .din(new_Jinkela_wire_5635),
        .dout(new_Jinkela_wire_5636)
    );

    bfr new_Jinkela_buffer_4496 (
        .din(_0184_),
        .dout(new_Jinkela_wire_5886)
    );

    spl2 new_Jinkela_splitter_543 (
        .a(_0213_),
        .b(new_Jinkela_wire_5884),
        .c(new_Jinkela_wire_5885)
    );

    bfr new_Jinkela_buffer_4313 (
        .din(new_Jinkela_wire_5636),
        .dout(new_Jinkela_wire_5637)
    );

    bfr new_Jinkela_buffer_4386 (
        .din(new_Jinkela_wire_5757),
        .dout(new_Jinkela_wire_5758)
    );

    bfr new_Jinkela_buffer_4314 (
        .din(new_Jinkela_wire_5637),
        .dout(new_Jinkela_wire_5638)
    );

    bfr new_Jinkela_buffer_4435 (
        .din(new_Jinkela_wire_5816),
        .dout(new_Jinkela_wire_5817)
    );

    bfr new_Jinkela_buffer_4315 (
        .din(new_Jinkela_wire_5638),
        .dout(new_Jinkela_wire_5639)
    );

    bfr new_Jinkela_buffer_4387 (
        .din(new_Jinkela_wire_5758),
        .dout(new_Jinkela_wire_5759)
    );

    bfr new_Jinkela_buffer_4316 (
        .din(new_Jinkela_wire_5639),
        .dout(new_Jinkela_wire_5640)
    );

    bfr new_Jinkela_buffer_7849 (
        .din(new_Jinkela_wire_9704),
        .dout(new_Jinkela_wire_9705)
    );

    bfr new_Jinkela_buffer_11234 (
        .din(new_Jinkela_wire_13539),
        .dout(new_Jinkela_wire_13540)
    );

    bfr new_Jinkela_buffer_7777 (
        .din(new_Jinkela_wire_9630),
        .dout(new_Jinkela_wire_9631)
    );

    bfr new_Jinkela_buffer_11235 (
        .din(new_Jinkela_wire_13540),
        .dout(new_Jinkela_wire_13541)
    );

    spl2 new_Jinkela_splitter_786 (
        .a(_1370_),
        .b(new_Jinkela_wire_9860),
        .c(new_Jinkela_wire_9861)
    );

    bfr new_Jinkela_buffer_7778 (
        .din(new_Jinkela_wire_9631),
        .dout(new_Jinkela_wire_9632)
    );

    bfr new_Jinkela_buffer_11303 (
        .din(new_Jinkela_wire_13622),
        .dout(new_Jinkela_wire_13623)
    );

    bfr new_Jinkela_buffer_7850 (
        .din(new_Jinkela_wire_9705),
        .dout(new_Jinkela_wire_9706)
    );

    bfr new_Jinkela_buffer_11236 (
        .din(new_Jinkela_wire_13541),
        .dout(new_Jinkela_wire_13542)
    );

    bfr new_Jinkela_buffer_7779 (
        .din(new_Jinkela_wire_9632),
        .dout(new_Jinkela_wire_9633)
    );

    bfr new_Jinkela_buffer_11368 (
        .din(new_Jinkela_wire_13701),
        .dout(new_Jinkela_wire_13702)
    );

    bfr new_Jinkela_buffer_7883 (
        .din(new_Jinkela_wire_9750),
        .dout(new_Jinkela_wire_9751)
    );

    bfr new_Jinkela_buffer_11237 (
        .din(new_Jinkela_wire_13542),
        .dout(new_Jinkela_wire_13543)
    );

    bfr new_Jinkela_buffer_7780 (
        .din(new_Jinkela_wire_9633),
        .dout(new_Jinkela_wire_9634)
    );

    bfr new_Jinkela_buffer_11304 (
        .din(new_Jinkela_wire_13623),
        .dout(new_Jinkela_wire_13624)
    );

    bfr new_Jinkela_buffer_7851 (
        .din(new_Jinkela_wire_9706),
        .dout(new_Jinkela_wire_9707)
    );

    bfr new_Jinkela_buffer_11238 (
        .din(new_Jinkela_wire_13543),
        .dout(new_Jinkela_wire_13544)
    );

    bfr new_Jinkela_buffer_7781 (
        .din(new_Jinkela_wire_9634),
        .dout(new_Jinkela_wire_9635)
    );

    bfr new_Jinkela_buffer_11386 (
        .din(new_Jinkela_wire_13727),
        .dout(new_Jinkela_wire_13728)
    );

    bfr new_Jinkela_buffer_11239 (
        .din(new_Jinkela_wire_13544),
        .dout(new_Jinkela_wire_13545)
    );

    bfr new_Jinkela_buffer_7985 (
        .din(_0402_),
        .dout(new_Jinkela_wire_9859)
    );

    bfr new_Jinkela_buffer_7782 (
        .din(new_Jinkela_wire_9635),
        .dout(new_Jinkela_wire_9636)
    );

    bfr new_Jinkela_buffer_11305 (
        .din(new_Jinkela_wire_13624),
        .dout(new_Jinkela_wire_13625)
    );

    bfr new_Jinkela_buffer_7852 (
        .din(new_Jinkela_wire_9707),
        .dout(new_Jinkela_wire_9708)
    );

    bfr new_Jinkela_buffer_11240 (
        .din(new_Jinkela_wire_13545),
        .dout(new_Jinkela_wire_13546)
    );

    bfr new_Jinkela_buffer_7783 (
        .din(new_Jinkela_wire_9636),
        .dout(new_Jinkela_wire_9637)
    );

    bfr new_Jinkela_buffer_11369 (
        .din(new_Jinkela_wire_13702),
        .dout(new_Jinkela_wire_13703)
    );

    bfr new_Jinkela_buffer_7884 (
        .din(new_Jinkela_wire_9751),
        .dout(new_Jinkela_wire_9752)
    );

    bfr new_Jinkela_buffer_11241 (
        .din(new_Jinkela_wire_13546),
        .dout(new_Jinkela_wire_13547)
    );

    bfr new_Jinkela_buffer_7784 (
        .din(new_Jinkela_wire_9637),
        .dout(new_Jinkela_wire_9638)
    );

    bfr new_Jinkela_buffer_11306 (
        .din(new_Jinkela_wire_13625),
        .dout(new_Jinkela_wire_13626)
    );

    bfr new_Jinkela_buffer_7853 (
        .din(new_Jinkela_wire_9708),
        .dout(new_Jinkela_wire_9709)
    );

    bfr new_Jinkela_buffer_11242 (
        .din(new_Jinkela_wire_13547),
        .dout(new_Jinkela_wire_13548)
    );

    bfr new_Jinkela_buffer_7785 (
        .din(new_Jinkela_wire_9638),
        .dout(new_Jinkela_wire_9639)
    );

    bfr new_Jinkela_buffer_11389 (
        .din(new_Jinkela_wire_13732),
        .dout(new_Jinkela_wire_13733)
    );

    bfr new_Jinkela_buffer_7938 (
        .din(new_Jinkela_wire_9809),
        .dout(new_Jinkela_wire_9810)
    );

    bfr new_Jinkela_buffer_11243 (
        .din(new_Jinkela_wire_13548),
        .dout(new_Jinkela_wire_13549)
    );

    bfr new_Jinkela_buffer_7786 (
        .din(new_Jinkela_wire_9639),
        .dout(new_Jinkela_wire_9640)
    );

    bfr new_Jinkela_buffer_11307 (
        .din(new_Jinkela_wire_13626),
        .dout(new_Jinkela_wire_13627)
    );

    bfr new_Jinkela_buffer_7854 (
        .din(new_Jinkela_wire_9709),
        .dout(new_Jinkela_wire_9710)
    );

    bfr new_Jinkela_buffer_11244 (
        .din(new_Jinkela_wire_13549),
        .dout(new_Jinkela_wire_13550)
    );

    bfr new_Jinkela_buffer_7787 (
        .din(new_Jinkela_wire_9640),
        .dout(new_Jinkela_wire_9641)
    );

    bfr new_Jinkela_buffer_11370 (
        .din(new_Jinkela_wire_13703),
        .dout(new_Jinkela_wire_13704)
    );

    bfr new_Jinkela_buffer_7885 (
        .din(new_Jinkela_wire_9752),
        .dout(new_Jinkela_wire_9753)
    );

    bfr new_Jinkela_buffer_11245 (
        .din(new_Jinkela_wire_13550),
        .dout(new_Jinkela_wire_13551)
    );

    bfr new_Jinkela_buffer_7788 (
        .din(new_Jinkela_wire_9641),
        .dout(new_Jinkela_wire_9642)
    );

    bfr new_Jinkela_buffer_11308 (
        .din(new_Jinkela_wire_13627),
        .dout(new_Jinkela_wire_13628)
    );

    bfr new_Jinkela_buffer_7855 (
        .din(new_Jinkela_wire_9710),
        .dout(new_Jinkela_wire_9711)
    );

    bfr new_Jinkela_buffer_11246 (
        .din(new_Jinkela_wire_13551),
        .dout(new_Jinkela_wire_13552)
    );

    bfr new_Jinkela_buffer_7789 (
        .din(new_Jinkela_wire_9642),
        .dout(new_Jinkela_wire_9643)
    );

    bfr new_Jinkela_buffer_11387 (
        .din(new_Jinkela_wire_13728),
        .dout(new_Jinkela_wire_13729)
    );

    spl2 new_Jinkela_splitter_787 (
        .a(_0828_),
        .b(new_Jinkela_wire_9862),
        .c(new_Jinkela_wire_9863)
    );

    bfr new_Jinkela_buffer_11247 (
        .din(new_Jinkela_wire_13552),
        .dout(new_Jinkela_wire_13553)
    );

    bfr new_Jinkela_buffer_7790 (
        .din(new_Jinkela_wire_9643),
        .dout(new_Jinkela_wire_9644)
    );

    bfr new_Jinkela_buffer_11309 (
        .din(new_Jinkela_wire_13628),
        .dout(new_Jinkela_wire_13629)
    );

    bfr new_Jinkela_buffer_7856 (
        .din(new_Jinkela_wire_9711),
        .dout(new_Jinkela_wire_9712)
    );

    bfr new_Jinkela_buffer_11248 (
        .din(new_Jinkela_wire_13553),
        .dout(new_Jinkela_wire_13554)
    );

    bfr new_Jinkela_buffer_7791 (
        .din(new_Jinkela_wire_9644),
        .dout(new_Jinkela_wire_9645)
    );

    bfr new_Jinkela_buffer_11371 (
        .din(new_Jinkela_wire_13704),
        .dout(new_Jinkela_wire_13705)
    );

    bfr new_Jinkela_buffer_7886 (
        .din(new_Jinkela_wire_9753),
        .dout(new_Jinkela_wire_9754)
    );

    bfr new_Jinkela_buffer_11249 (
        .din(new_Jinkela_wire_13554),
        .dout(new_Jinkela_wire_13555)
    );

    bfr new_Jinkela_buffer_7792 (
        .din(new_Jinkela_wire_9645),
        .dout(new_Jinkela_wire_9646)
    );

    bfr new_Jinkela_buffer_11310 (
        .din(new_Jinkela_wire_13629),
        .dout(new_Jinkela_wire_13630)
    );

    bfr new_Jinkela_buffer_7857 (
        .din(new_Jinkela_wire_9712),
        .dout(new_Jinkela_wire_9713)
    );

    bfr new_Jinkela_buffer_11250 (
        .din(new_Jinkela_wire_13555),
        .dout(new_Jinkela_wire_13556)
    );

    bfr new_Jinkela_buffer_7793 (
        .din(new_Jinkela_wire_9646),
        .dout(new_Jinkela_wire_9647)
    );

    spl2 new_Jinkela_splitter_1032 (
        .a(_1503_),
        .b(new_Jinkela_wire_13990),
        .c(new_Jinkela_wire_13991)
    );

    spl2 new_Jinkela_splitter_1031 (
        .a(_0508_),
        .b(new_Jinkela_wire_13984),
        .c(new_Jinkela_wire_13985)
    );

    bfr new_Jinkela_buffer_7939 (
        .din(new_Jinkela_wire_9810),
        .dout(new_Jinkela_wire_9811)
    );

    bfr new_Jinkela_buffer_11251 (
        .din(new_Jinkela_wire_13556),
        .dout(new_Jinkela_wire_13557)
    );

    bfr new_Jinkela_buffer_7794 (
        .din(new_Jinkela_wire_9647),
        .dout(new_Jinkela_wire_9648)
    );

    bfr new_Jinkela_buffer_11311 (
        .din(new_Jinkela_wire_13630),
        .dout(new_Jinkela_wire_13631)
    );

    bfr new_Jinkela_buffer_7858 (
        .din(new_Jinkela_wire_9713),
        .dout(new_Jinkela_wire_9714)
    );

    bfr new_Jinkela_buffer_11252 (
        .din(new_Jinkela_wire_13557),
        .dout(new_Jinkela_wire_13558)
    );

    bfr new_Jinkela_buffer_7795 (
        .din(new_Jinkela_wire_9648),
        .dout(new_Jinkela_wire_9649)
    );

    bfr new_Jinkela_buffer_11372 (
        .din(new_Jinkela_wire_13705),
        .dout(new_Jinkela_wire_13706)
    );

    bfr new_Jinkela_buffer_7887 (
        .din(new_Jinkela_wire_9754),
        .dout(new_Jinkela_wire_9755)
    );

    bfr new_Jinkela_buffer_11253 (
        .din(new_Jinkela_wire_13558),
        .dout(new_Jinkela_wire_13559)
    );

    bfr new_Jinkela_buffer_7796 (
        .din(new_Jinkela_wire_9649),
        .dout(new_Jinkela_wire_9650)
    );

    bfr new_Jinkela_buffer_11312 (
        .din(new_Jinkela_wire_13631),
        .dout(new_Jinkela_wire_13632)
    );

    bfr new_Jinkela_buffer_7859 (
        .din(new_Jinkela_wire_9714),
        .dout(new_Jinkela_wire_9715)
    );

    bfr new_Jinkela_buffer_11254 (
        .din(new_Jinkela_wire_13559),
        .dout(new_Jinkela_wire_13560)
    );

    bfr new_Jinkela_buffer_7797 (
        .din(new_Jinkela_wire_9650),
        .dout(new_Jinkela_wire_9651)
    );

    bfr new_Jinkela_buffer_11390 (
        .din(new_Jinkela_wire_13733),
        .dout(new_Jinkela_wire_13734)
    );

    bfr new_Jinkela_buffer_14810 (
        .din(new_Jinkela_wire_17684),
        .dout(new_Jinkela_wire_17685)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_1469),
        .dout(new_Jinkela_wire_1470)
    );

    bfr new_Jinkela_buffer_14690 (
        .din(new_Jinkela_wire_17520),
        .dout(new_Jinkela_wire_17521)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1642),
        .dout(new_Jinkela_wire_1643)
    );

    bfr new_Jinkela_buffer_14745 (
        .din(new_Jinkela_wire_17595),
        .dout(new_Jinkela_wire_17596)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_1470),
        .dout(new_Jinkela_wire_1471)
    );

    bfr new_Jinkela_buffer_14691 (
        .din(new_Jinkela_wire_17521),
        .dout(new_Jinkela_wire_17522)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1677),
        .dout(new_Jinkela_wire_1678)
    );

    spl2 new_Jinkela_splitter_1289 (
        .a(_1267_),
        .b(new_Jinkela_wire_17788),
        .c(new_Jinkela_wire_17789)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_1471),
        .dout(new_Jinkela_wire_1472)
    );

    bfr new_Jinkela_buffer_14692 (
        .din(new_Jinkela_wire_17522),
        .dout(new_Jinkela_wire_17523)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    bfr new_Jinkela_buffer_14746 (
        .din(new_Jinkela_wire_17596),
        .dout(new_Jinkela_wire_17597)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_1472),
        .dout(new_Jinkela_wire_1473)
    );

    bfr new_Jinkela_buffer_14693 (
        .din(new_Jinkela_wire_17523),
        .dout(new_Jinkela_wire_17524)
    );

    bfr new_Jinkela_buffer_14811 (
        .din(new_Jinkela_wire_17685),
        .dout(new_Jinkela_wire_17686)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1767),
        .dout(new_Jinkela_wire_1768)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_1473),
        .dout(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_14694 (
        .din(new_Jinkela_wire_17524),
        .dout(new_Jinkela_wire_17525)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1644),
        .dout(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_14747 (
        .din(new_Jinkela_wire_17597),
        .dout(new_Jinkela_wire_17598)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_1474),
        .dout(new_Jinkela_wire_1475)
    );

    bfr new_Jinkela_buffer_14695 (
        .din(new_Jinkela_wire_17525),
        .dout(new_Jinkela_wire_17526)
    );

    bfr new_Jinkela_buffer_14850 (
        .din(new_Jinkela_wire_17726),
        .dout(new_Jinkela_wire_17727)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1678),
        .dout(new_Jinkela_wire_1679)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_1475),
        .dout(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_14696 (
        .din(new_Jinkela_wire_17526),
        .dout(new_Jinkela_wire_17527)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1645),
        .dout(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_14748 (
        .din(new_Jinkela_wire_17598),
        .dout(new_Jinkela_wire_17599)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_1476),
        .dout(new_Jinkela_wire_1477)
    );

    bfr new_Jinkela_buffer_14697 (
        .din(new_Jinkela_wire_17527),
        .dout(new_Jinkela_wire_17528)
    );

    bfr new_Jinkela_buffer_14812 (
        .din(new_Jinkela_wire_17686),
        .dout(new_Jinkela_wire_17687)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    bfr new_Jinkela_buffer_14698 (
        .din(new_Jinkela_wire_17528),
        .dout(new_Jinkela_wire_17529)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_14749 (
        .din(new_Jinkela_wire_17599),
        .dout(new_Jinkela_wire_17600)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    spl2 new_Jinkela_splitter_1264 (
        .a(new_Jinkela_wire_17529),
        .b(new_Jinkela_wire_17530),
        .c(new_Jinkela_wire_17531)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(_0613_),
        .b(new_Jinkela_wire_1775),
        .c(new_Jinkela_wire_1776)
    );

    bfr new_Jinkela_buffer_14750 (
        .din(new_Jinkela_wire_17600),
        .dout(new_Jinkela_wire_17601)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1679),
        .dout(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_1479),
        .dout(new_Jinkela_wire_1480)
    );

    bfr new_Jinkela_buffer_14911 (
        .din(_1098_),
        .dout(new_Jinkela_wire_17794)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_1647),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_14813 (
        .din(new_Jinkela_wire_17687),
        .dout(new_Jinkela_wire_17688)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_1480),
        .dout(new_Jinkela_wire_1481)
    );

    bfr new_Jinkela_buffer_14751 (
        .din(new_Jinkela_wire_17601),
        .dout(new_Jinkela_wire_17602)
    );

    bfr new_Jinkela_buffer_14851 (
        .din(new_Jinkela_wire_17727),
        .dout(new_Jinkela_wire_17728)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1768),
        .dout(new_Jinkela_wire_1769)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_1481),
        .dout(new_Jinkela_wire_1482)
    );

    bfr new_Jinkela_buffer_14752 (
        .din(new_Jinkela_wire_17602),
        .dout(new_Jinkela_wire_17603)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_14814 (
        .din(new_Jinkela_wire_17688),
        .dout(new_Jinkela_wire_17689)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_1482),
        .dout(new_Jinkela_wire_1483)
    );

    bfr new_Jinkela_buffer_14753 (
        .din(new_Jinkela_wire_17603),
        .dout(new_Jinkela_wire_17604)
    );

    bfr new_Jinkela_buffer_14906 (
        .din(new_Jinkela_wire_17784),
        .dout(new_Jinkela_wire_17785)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1680),
        .dout(new_Jinkela_wire_1681)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_1483),
        .dout(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_14754 (
        .din(new_Jinkela_wire_17604),
        .dout(new_Jinkela_wire_17605)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_14815 (
        .din(new_Jinkela_wire_17689),
        .dout(new_Jinkela_wire_17690)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_1484),
        .dout(new_Jinkela_wire_1485)
    );

    bfr new_Jinkela_buffer_14755 (
        .din(new_Jinkela_wire_17605),
        .dout(new_Jinkela_wire_17606)
    );

    bfr new_Jinkela_buffer_14852 (
        .din(new_Jinkela_wire_17728),
        .dout(new_Jinkela_wire_17729)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(_0137_),
        .b(new_Jinkela_wire_1779),
        .c(new_Jinkela_wire_1780)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_1485),
        .dout(new_Jinkela_wire_1486)
    );

    bfr new_Jinkela_buffer_14756 (
        .din(new_Jinkela_wire_17606),
        .dout(new_Jinkela_wire_17607)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1650),
        .dout(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_14816 (
        .din(new_Jinkela_wire_17690),
        .dout(new_Jinkela_wire_17691)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_14757 (
        .din(new_Jinkela_wire_17607),
        .dout(new_Jinkela_wire_17608)
    );

    spl2 new_Jinkela_splitter_247 (
        .a(_1464_),
        .b(new_Jinkela_wire_1777),
        .c(new_Jinkela_wire_1778)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_1681),
        .dout(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_14907 (
        .din(new_Jinkela_wire_17789),
        .dout(new_Jinkela_wire_17790)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_1487),
        .dout(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_14758 (
        .din(new_Jinkela_wire_17608),
        .dout(new_Jinkela_wire_17609)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1651),
        .dout(new_Jinkela_wire_1652)
    );

    bfr new_Jinkela_buffer_14817 (
        .din(new_Jinkela_wire_17691),
        .dout(new_Jinkela_wire_17692)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_1488),
        .dout(new_Jinkela_wire_1489)
    );

    bfr new_Jinkela_buffer_14759 (
        .din(new_Jinkela_wire_17609),
        .dout(new_Jinkela_wire_17610)
    );

    bfr new_Jinkela_buffer_14853 (
        .din(new_Jinkela_wire_17729),
        .dout(new_Jinkela_wire_17730)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1769),
        .dout(new_Jinkela_wire_1770)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_14760 (
        .din(new_Jinkela_wire_17610),
        .dout(new_Jinkela_wire_17611)
    );

    bfr new_Jinkela_buffer_4575 (
        .din(_1202_),
        .dout(new_Jinkela_wire_5967)
    );

    bfr new_Jinkela_buffer_7798 (
        .din(new_Jinkela_wire_9651),
        .dout(new_Jinkela_wire_9652)
    );

    bfr new_Jinkela_buffer_4317 (
        .din(new_Jinkela_wire_5640),
        .dout(new_Jinkela_wire_5641)
    );

    bfr new_Jinkela_buffer_7860 (
        .din(new_Jinkela_wire_9715),
        .dout(new_Jinkela_wire_9716)
    );

    bfr new_Jinkela_buffer_4388 (
        .din(new_Jinkela_wire_5759),
        .dout(new_Jinkela_wire_5760)
    );

    bfr new_Jinkela_buffer_7799 (
        .din(new_Jinkela_wire_9652),
        .dout(new_Jinkela_wire_9653)
    );

    bfr new_Jinkela_buffer_4318 (
        .din(new_Jinkela_wire_5641),
        .dout(new_Jinkela_wire_5642)
    );

    bfr new_Jinkela_buffer_7888 (
        .din(new_Jinkela_wire_9755),
        .dout(new_Jinkela_wire_9756)
    );

    bfr new_Jinkela_buffer_4436 (
        .din(new_Jinkela_wire_5817),
        .dout(new_Jinkela_wire_5818)
    );

    bfr new_Jinkela_buffer_7800 (
        .din(new_Jinkela_wire_9653),
        .dout(new_Jinkela_wire_9654)
    );

    bfr new_Jinkela_buffer_4319 (
        .din(new_Jinkela_wire_5642),
        .dout(new_Jinkela_wire_5643)
    );

    bfr new_Jinkela_buffer_7861 (
        .din(new_Jinkela_wire_9716),
        .dout(new_Jinkela_wire_9717)
    );

    bfr new_Jinkela_buffer_4389 (
        .din(new_Jinkela_wire_5760),
        .dout(new_Jinkela_wire_5761)
    );

    bfr new_Jinkela_buffer_7801 (
        .din(new_Jinkela_wire_9654),
        .dout(new_Jinkela_wire_9655)
    );

    bfr new_Jinkela_buffer_4320 (
        .din(new_Jinkela_wire_5643),
        .dout(new_Jinkela_wire_5644)
    );

    bfr new_Jinkela_buffer_7940 (
        .din(new_Jinkela_wire_9811),
        .dout(new_Jinkela_wire_9812)
    );

    bfr new_Jinkela_buffer_4497 (
        .din(_0776_),
        .dout(new_Jinkela_wire_5887)
    );

    bfr new_Jinkela_buffer_7802 (
        .din(new_Jinkela_wire_9655),
        .dout(new_Jinkela_wire_9656)
    );

    bfr new_Jinkela_buffer_4321 (
        .din(new_Jinkela_wire_5644),
        .dout(new_Jinkela_wire_5645)
    );

    bfr new_Jinkela_buffer_7862 (
        .din(new_Jinkela_wire_9717),
        .dout(new_Jinkela_wire_9718)
    );

    bfr new_Jinkela_buffer_4390 (
        .din(new_Jinkela_wire_5761),
        .dout(new_Jinkela_wire_5762)
    );

    bfr new_Jinkela_buffer_7803 (
        .din(new_Jinkela_wire_9656),
        .dout(new_Jinkela_wire_9657)
    );

    bfr new_Jinkela_buffer_4322 (
        .din(new_Jinkela_wire_5645),
        .dout(new_Jinkela_wire_5646)
    );

    bfr new_Jinkela_buffer_7889 (
        .din(new_Jinkela_wire_9756),
        .dout(new_Jinkela_wire_9757)
    );

    bfr new_Jinkela_buffer_4437 (
        .din(new_Jinkela_wire_5818),
        .dout(new_Jinkela_wire_5819)
    );

    bfr new_Jinkela_buffer_7804 (
        .din(new_Jinkela_wire_9657),
        .dout(new_Jinkela_wire_9658)
    );

    bfr new_Jinkela_buffer_4323 (
        .din(new_Jinkela_wire_5646),
        .dout(new_Jinkela_wire_5647)
    );

    bfr new_Jinkela_buffer_7863 (
        .din(new_Jinkela_wire_9718),
        .dout(new_Jinkela_wire_9719)
    );

    bfr new_Jinkela_buffer_4391 (
        .din(new_Jinkela_wire_5762),
        .dout(new_Jinkela_wire_5763)
    );

    bfr new_Jinkela_buffer_7805 (
        .din(new_Jinkela_wire_9658),
        .dout(new_Jinkela_wire_9659)
    );

    bfr new_Jinkela_buffer_4324 (
        .din(new_Jinkela_wire_5647),
        .dout(new_Jinkela_wire_5648)
    );

    spl2 new_Jinkela_splitter_545 (
        .a(_1289_),
        .b(new_Jinkela_wire_5968),
        .c(new_Jinkela_wire_5969)
    );

    spl2 new_Jinkela_splitter_788 (
        .a(_1553_),
        .b(new_Jinkela_wire_9864),
        .c(new_Jinkela_wire_9865)
    );

    bfr new_Jinkela_buffer_7806 (
        .din(new_Jinkela_wire_9659),
        .dout(new_Jinkela_wire_9660)
    );

    bfr new_Jinkela_buffer_4325 (
        .din(new_Jinkela_wire_5648),
        .dout(new_Jinkela_wire_5649)
    );

    bfr new_Jinkela_buffer_7864 (
        .din(new_Jinkela_wire_9719),
        .dout(new_Jinkela_wire_9720)
    );

    bfr new_Jinkela_buffer_4392 (
        .din(new_Jinkela_wire_5763),
        .dout(new_Jinkela_wire_5764)
    );

    bfr new_Jinkela_buffer_7807 (
        .din(new_Jinkela_wire_9660),
        .dout(new_Jinkela_wire_9661)
    );

    bfr new_Jinkela_buffer_4326 (
        .din(new_Jinkela_wire_5649),
        .dout(new_Jinkela_wire_5650)
    );

    bfr new_Jinkela_buffer_7890 (
        .din(new_Jinkela_wire_9757),
        .dout(new_Jinkela_wire_9758)
    );

    bfr new_Jinkela_buffer_4438 (
        .din(new_Jinkela_wire_5819),
        .dout(new_Jinkela_wire_5820)
    );

    bfr new_Jinkela_buffer_7808 (
        .din(new_Jinkela_wire_9661),
        .dout(new_Jinkela_wire_9662)
    );

    bfr new_Jinkela_buffer_4327 (
        .din(new_Jinkela_wire_5650),
        .dout(new_Jinkela_wire_5651)
    );

    bfr new_Jinkela_buffer_7865 (
        .din(new_Jinkela_wire_9720),
        .dout(new_Jinkela_wire_9721)
    );

    bfr new_Jinkela_buffer_4393 (
        .din(new_Jinkela_wire_5764),
        .dout(new_Jinkela_wire_5765)
    );

    bfr new_Jinkela_buffer_7809 (
        .din(new_Jinkela_wire_9662),
        .dout(new_Jinkela_wire_9663)
    );

    bfr new_Jinkela_buffer_4328 (
        .din(new_Jinkela_wire_5651),
        .dout(new_Jinkela_wire_5652)
    );

    bfr new_Jinkela_buffer_7941 (
        .din(new_Jinkela_wire_9812),
        .dout(new_Jinkela_wire_9813)
    );

    bfr new_Jinkela_buffer_4498 (
        .din(new_Jinkela_wire_5887),
        .dout(new_Jinkela_wire_5888)
    );

    bfr new_Jinkela_buffer_7810 (
        .din(new_Jinkela_wire_9663),
        .dout(new_Jinkela_wire_9664)
    );

    bfr new_Jinkela_buffer_4329 (
        .din(new_Jinkela_wire_5652),
        .dout(new_Jinkela_wire_5653)
    );

    bfr new_Jinkela_buffer_7866 (
        .din(new_Jinkela_wire_9721),
        .dout(new_Jinkela_wire_9722)
    );

    bfr new_Jinkela_buffer_4394 (
        .din(new_Jinkela_wire_5765),
        .dout(new_Jinkela_wire_5766)
    );

    bfr new_Jinkela_buffer_7811 (
        .din(new_Jinkela_wire_9664),
        .dout(new_Jinkela_wire_9665)
    );

    bfr new_Jinkela_buffer_4330 (
        .din(new_Jinkela_wire_5653),
        .dout(new_Jinkela_wire_5654)
    );

    bfr new_Jinkela_buffer_7891 (
        .din(new_Jinkela_wire_9758),
        .dout(new_Jinkela_wire_9759)
    );

    bfr new_Jinkela_buffer_4439 (
        .din(new_Jinkela_wire_5820),
        .dout(new_Jinkela_wire_5821)
    );

    bfr new_Jinkela_buffer_7812 (
        .din(new_Jinkela_wire_9665),
        .dout(new_Jinkela_wire_9666)
    );

    bfr new_Jinkela_buffer_4331 (
        .din(new_Jinkela_wire_5654),
        .dout(new_Jinkela_wire_5655)
    );

    bfr new_Jinkela_buffer_7867 (
        .din(new_Jinkela_wire_9722),
        .dout(new_Jinkela_wire_9723)
    );

    bfr new_Jinkela_buffer_4395 (
        .din(new_Jinkela_wire_5766),
        .dout(new_Jinkela_wire_5767)
    );

    bfr new_Jinkela_buffer_7813 (
        .din(new_Jinkela_wire_9666),
        .dout(new_Jinkela_wire_9667)
    );

    bfr new_Jinkela_buffer_4332 (
        .din(new_Jinkela_wire_5655),
        .dout(new_Jinkela_wire_5656)
    );

    bfr new_Jinkela_buffer_8026 (
        .din(new_net_3954),
        .dout(new_Jinkela_wire_9908)
    );

    bfr new_Jinkela_buffer_4576 (
        .din(_0611_),
        .dout(new_Jinkela_wire_5970)
    );

    bfr new_Jinkela_buffer_7986 (
        .din(_1467_),
        .dout(new_Jinkela_wire_9866)
    );

    bfr new_Jinkela_buffer_7814 (
        .din(new_Jinkela_wire_9667),
        .dout(new_Jinkela_wire_9668)
    );

    bfr new_Jinkela_buffer_4333 (
        .din(new_Jinkela_wire_5656),
        .dout(new_Jinkela_wire_5657)
    );

    bfr new_Jinkela_buffer_7868 (
        .din(new_Jinkela_wire_9723),
        .dout(new_Jinkela_wire_9724)
    );

    bfr new_Jinkela_buffer_4396 (
        .din(new_Jinkela_wire_5767),
        .dout(new_Jinkela_wire_5768)
    );

    bfr new_Jinkela_buffer_7815 (
        .din(new_Jinkela_wire_9668),
        .dout(new_Jinkela_wire_9669)
    );

    bfr new_Jinkela_buffer_4334 (
        .din(new_Jinkela_wire_5657),
        .dout(new_Jinkela_wire_5658)
    );

    bfr new_Jinkela_buffer_7892 (
        .din(new_Jinkela_wire_9759),
        .dout(new_Jinkela_wire_9760)
    );

    bfr new_Jinkela_buffer_4440 (
        .din(new_Jinkela_wire_5821),
        .dout(new_Jinkela_wire_5822)
    );

    bfr new_Jinkela_buffer_7816 (
        .din(new_Jinkela_wire_9669),
        .dout(new_Jinkela_wire_9670)
    );

    bfr new_Jinkela_buffer_4335 (
        .din(new_Jinkela_wire_5658),
        .dout(new_Jinkela_wire_5659)
    );

    bfr new_Jinkela_buffer_7869 (
        .din(new_Jinkela_wire_9724),
        .dout(new_Jinkela_wire_9725)
    );

    bfr new_Jinkela_buffer_4397 (
        .din(new_Jinkela_wire_5768),
        .dout(new_Jinkela_wire_5769)
    );

    bfr new_Jinkela_buffer_7817 (
        .din(new_Jinkela_wire_9670),
        .dout(new_Jinkela_wire_9671)
    );

    bfr new_Jinkela_buffer_4336 (
        .din(new_Jinkela_wire_5659),
        .dout(new_Jinkela_wire_5660)
    );

    bfr new_Jinkela_buffer_7942 (
        .din(new_Jinkela_wire_9813),
        .dout(new_Jinkela_wire_9814)
    );

    bfr new_Jinkela_buffer_4499 (
        .din(new_Jinkela_wire_5888),
        .dout(new_Jinkela_wire_5889)
    );

    bfr new_Jinkela_buffer_7818 (
        .din(new_Jinkela_wire_9671),
        .dout(new_Jinkela_wire_9672)
    );

    bfr new_Jinkela_buffer_4337 (
        .din(new_Jinkela_wire_5660),
        .dout(new_Jinkela_wire_5661)
    );

    bfr new_Jinkela_buffer_11255 (
        .din(new_Jinkela_wire_13560),
        .dout(new_Jinkela_wire_13561)
    );

    bfr new_Jinkela_buffer_11313 (
        .din(new_Jinkela_wire_13632),
        .dout(new_Jinkela_wire_13633)
    );

    bfr new_Jinkela_buffer_11256 (
        .din(new_Jinkela_wire_13561),
        .dout(new_Jinkela_wire_13562)
    );

    bfr new_Jinkela_buffer_11373 (
        .din(new_Jinkela_wire_13706),
        .dout(new_Jinkela_wire_13707)
    );

    bfr new_Jinkela_buffer_11257 (
        .din(new_Jinkela_wire_13562),
        .dout(new_Jinkela_wire_13563)
    );

    bfr new_Jinkela_buffer_11314 (
        .din(new_Jinkela_wire_13633),
        .dout(new_Jinkela_wire_13634)
    );

    bfr new_Jinkela_buffer_11258 (
        .din(new_Jinkela_wire_13563),
        .dout(new_Jinkela_wire_13564)
    );

    bfr new_Jinkela_buffer_11604 (
        .din(_0819_),
        .dout(new_Jinkela_wire_13954)
    );

    bfr new_Jinkela_buffer_11259 (
        .din(new_Jinkela_wire_13564),
        .dout(new_Jinkela_wire_13565)
    );

    bfr new_Jinkela_buffer_11315 (
        .din(new_Jinkela_wire_13634),
        .dout(new_Jinkela_wire_13635)
    );

    bfr new_Jinkela_buffer_11260 (
        .din(new_Jinkela_wire_13565),
        .dout(new_Jinkela_wire_13566)
    );

    bfr new_Jinkela_buffer_11374 (
        .din(new_Jinkela_wire_13707),
        .dout(new_Jinkela_wire_13708)
    );

    bfr new_Jinkela_buffer_11261 (
        .din(new_Jinkela_wire_13566),
        .dout(new_Jinkela_wire_13567)
    );

    bfr new_Jinkela_buffer_11316 (
        .din(new_Jinkela_wire_13635),
        .dout(new_Jinkela_wire_13636)
    );

    bfr new_Jinkela_buffer_11262 (
        .din(new_Jinkela_wire_13567),
        .dout(new_Jinkela_wire_13568)
    );

    bfr new_Jinkela_buffer_11391 (
        .din(new_Jinkela_wire_13734),
        .dout(new_Jinkela_wire_13735)
    );

    bfr new_Jinkela_buffer_11263 (
        .din(new_Jinkela_wire_13568),
        .dout(new_Jinkela_wire_13569)
    );

    bfr new_Jinkela_buffer_11317 (
        .din(new_Jinkela_wire_13636),
        .dout(new_Jinkela_wire_13637)
    );

    spl2 new_Jinkela_splitter_1002 (
        .a(new_Jinkela_wire_13569),
        .b(new_Jinkela_wire_13570),
        .c(new_Jinkela_wire_13571)
    );

    bfr new_Jinkela_buffer_11318 (
        .din(new_Jinkela_wire_13637),
        .dout(new_Jinkela_wire_13638)
    );

    bfr new_Jinkela_buffer_11375 (
        .din(new_Jinkela_wire_13708),
        .dout(new_Jinkela_wire_13709)
    );

    spl2 new_Jinkela_splitter_1024 (
        .a(_1128_),
        .b(new_Jinkela_wire_13955),
        .c(new_Jinkela_wire_13956)
    );

    bfr new_Jinkela_buffer_11319 (
        .din(new_Jinkela_wire_13638),
        .dout(new_Jinkela_wire_13639)
    );

    bfr new_Jinkela_buffer_11376 (
        .din(new_Jinkela_wire_13709),
        .dout(new_Jinkela_wire_13710)
    );

    bfr new_Jinkela_buffer_11320 (
        .din(new_Jinkela_wire_13639),
        .dout(new_Jinkela_wire_13640)
    );

    bfr new_Jinkela_buffer_11392 (
        .din(new_Jinkela_wire_13735),
        .dout(new_Jinkela_wire_13736)
    );

    bfr new_Jinkela_buffer_11321 (
        .din(new_Jinkela_wire_13640),
        .dout(new_Jinkela_wire_13641)
    );

    bfr new_Jinkela_buffer_11377 (
        .din(new_Jinkela_wire_13710),
        .dout(new_Jinkela_wire_13711)
    );

    bfr new_Jinkela_buffer_11322 (
        .din(new_Jinkela_wire_13641),
        .dout(new_Jinkela_wire_13642)
    );

    bfr new_Jinkela_buffer_11501 (
        .din(new_Jinkela_wire_13848),
        .dout(new_Jinkela_wire_13849)
    );

    bfr new_Jinkela_buffer_11323 (
        .din(new_Jinkela_wire_13642),
        .dout(new_Jinkela_wire_13643)
    );

    bfr new_Jinkela_buffer_11378 (
        .din(new_Jinkela_wire_13711),
        .dout(new_Jinkela_wire_13712)
    );

    bfr new_Jinkela_buffer_11324 (
        .din(new_Jinkela_wire_13643),
        .dout(new_Jinkela_wire_13644)
    );

    bfr new_Jinkela_buffer_11393 (
        .din(new_Jinkela_wire_13736),
        .dout(new_Jinkela_wire_13737)
    );

    bfr new_Jinkela_buffer_11325 (
        .din(new_Jinkela_wire_13644),
        .dout(new_Jinkela_wire_13645)
    );

    bfr new_Jinkela_buffer_11379 (
        .din(new_Jinkela_wire_13712),
        .dout(new_Jinkela_wire_13713)
    );

    bfr new_Jinkela_buffer_11326 (
        .din(new_Jinkela_wire_13645),
        .dout(new_Jinkela_wire_13646)
    );

    bfr new_Jinkela_buffer_11605 (
        .din(_0558_),
        .dout(new_Jinkela_wire_13957)
    );

    bfr new_Jinkela_buffer_11500 (
        .din(_0699_),
        .dout(new_Jinkela_wire_13848)
    );

    bfr new_Jinkela_buffer_11327 (
        .din(new_Jinkela_wire_13646),
        .dout(new_Jinkela_wire_13647)
    );

    bfr new_Jinkela_buffer_11380 (
        .din(new_Jinkela_wire_13713),
        .dout(new_Jinkela_wire_13714)
    );

    bfr new_Jinkela_buffer_11328 (
        .din(new_Jinkela_wire_13647),
        .dout(new_Jinkela_wire_13648)
    );

    bfr new_Jinkela_buffer_11394 (
        .din(new_Jinkela_wire_13737),
        .dout(new_Jinkela_wire_13738)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1652),
        .dout(new_Jinkela_wire_1653)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1682),
        .dout(new_Jinkela_wire_1683)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_1491),
        .dout(new_Jinkela_wire_1492)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1653),
        .dout(new_Jinkela_wire_1654)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_1492),
        .dout(new_Jinkela_wire_1493)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_1493),
        .dout(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1654),
        .dout(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_1494),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1683),
        .dout(new_Jinkela_wire_1684)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_1495),
        .dout(new_Jinkela_wire_1496)
    );

    bfr new_Jinkela_buffer_872 (
        .din(new_Jinkela_wire_1655),
        .dout(new_Jinkela_wire_1656)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_1496),
        .dout(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_1497),
        .dout(new_Jinkela_wire_1498)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_1656),
        .dout(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_1498),
        .dout(new_Jinkela_wire_1499)
    );

    bfr new_Jinkela_buffer_981 (
        .din(_0653_),
        .dout(new_Jinkela_wire_1781)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1684),
        .dout(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_1499),
        .dout(new_Jinkela_wire_1500)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_1657),
        .dout(new_Jinkela_wire_1658)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_1500),
        .dout(new_Jinkela_wire_1501)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(_1380_),
        .b(new_Jinkela_wire_1788),
        .c(new_Jinkela_wire_1789)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_1501),
        .dout(new_Jinkela_wire_1502)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_Jinkela_wire_1658),
        .dout(new_Jinkela_wire_1659)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_1502),
        .dout(new_Jinkela_wire_1503)
    );

    bfr new_Jinkela_buffer_982 (
        .din(_0555_),
        .dout(new_Jinkela_wire_1782)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_1503),
        .dout(new_Jinkela_wire_1504)
    );

    bfr new_Jinkela_buffer_876 (
        .din(new_Jinkela_wire_1659),
        .dout(new_Jinkela_wire_1660)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_1504),
        .dout(new_Jinkela_wire_1505)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_1505),
        .dout(new_Jinkela_wire_1506)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1660),
        .dout(new_Jinkela_wire_1661)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_1506),
        .dout(new_Jinkela_wire_1507)
    );

    bfr new_Jinkela_buffer_986 (
        .din(_0383_),
        .dout(new_Jinkela_wire_1790)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1686),
        .dout(new_Jinkela_wire_1687)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1661),
        .dout(new_Jinkela_wire_1662)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1782),
        .dout(new_Jinkela_wire_1783)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1662),
        .dout(new_Jinkela_wire_1663)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_7870 (
        .din(new_Jinkela_wire_9725),
        .dout(new_Jinkela_wire_9726)
    );

    bfr new_Jinkela_buffer_4398 (
        .din(new_Jinkela_wire_5769),
        .dout(new_Jinkela_wire_5770)
    );

    bfr new_Jinkela_buffer_7819 (
        .din(new_Jinkela_wire_9672),
        .dout(new_Jinkela_wire_9673)
    );

    spl2 new_Jinkela_splitter_511 (
        .a(new_Jinkela_wire_5661),
        .b(new_Jinkela_wire_5662),
        .c(new_Jinkela_wire_5663)
    );

    bfr new_Jinkela_buffer_7893 (
        .din(new_Jinkela_wire_9760),
        .dout(new_Jinkela_wire_9761)
    );

    bfr new_Jinkela_buffer_4399 (
        .din(new_Jinkela_wire_5770),
        .dout(new_Jinkela_wire_5771)
    );

    bfr new_Jinkela_buffer_7820 (
        .din(new_Jinkela_wire_9673),
        .dout(new_Jinkela_wire_9674)
    );

    bfr new_Jinkela_buffer_4441 (
        .din(new_Jinkela_wire_5822),
        .dout(new_Jinkela_wire_5823)
    );

    bfr new_Jinkela_buffer_7871 (
        .din(new_Jinkela_wire_9726),
        .dout(new_Jinkela_wire_9727)
    );

    bfr new_Jinkela_buffer_4592 (
        .din(_0567_),
        .dout(new_Jinkela_wire_5990)
    );

    bfr new_Jinkela_buffer_7821 (
        .din(new_Jinkela_wire_9674),
        .dout(new_Jinkela_wire_9675)
    );

    bfr new_Jinkela_buffer_4400 (
        .din(new_Jinkela_wire_5771),
        .dout(new_Jinkela_wire_5772)
    );

    bfr new_Jinkela_buffer_4442 (
        .din(new_Jinkela_wire_5823),
        .dout(new_Jinkela_wire_5824)
    );

    bfr new_Jinkela_buffer_8166 (
        .din(_0111_),
        .dout(new_Jinkela_wire_10048)
    );

    bfr new_Jinkela_buffer_7822 (
        .din(new_Jinkela_wire_9675),
        .dout(new_Jinkela_wire_9676)
    );

    bfr new_Jinkela_buffer_4401 (
        .din(new_Jinkela_wire_5772),
        .dout(new_Jinkela_wire_5773)
    );

    bfr new_Jinkela_buffer_7872 (
        .din(new_Jinkela_wire_9727),
        .dout(new_Jinkela_wire_9728)
    );

    bfr new_Jinkela_buffer_4500 (
        .din(new_Jinkela_wire_5889),
        .dout(new_Jinkela_wire_5890)
    );

    bfr new_Jinkela_buffer_7823 (
        .din(new_Jinkela_wire_9676),
        .dout(new_Jinkela_wire_9677)
    );

    bfr new_Jinkela_buffer_4402 (
        .din(new_Jinkela_wire_5773),
        .dout(new_Jinkela_wire_5774)
    );

    bfr new_Jinkela_buffer_7894 (
        .din(new_Jinkela_wire_9761),
        .dout(new_Jinkela_wire_9762)
    );

    bfr new_Jinkela_buffer_4443 (
        .din(new_Jinkela_wire_5824),
        .dout(new_Jinkela_wire_5825)
    );

    bfr new_Jinkela_buffer_7824 (
        .din(new_Jinkela_wire_9677),
        .dout(new_Jinkela_wire_9678)
    );

    bfr new_Jinkela_buffer_4403 (
        .din(new_Jinkela_wire_5774),
        .dout(new_Jinkela_wire_5775)
    );

    bfr new_Jinkela_buffer_7873 (
        .din(new_Jinkela_wire_9728),
        .dout(new_Jinkela_wire_9729)
    );

    spl2 new_Jinkela_splitter_547 (
        .a(_0635_),
        .b(new_Jinkela_wire_5988),
        .c(new_Jinkela_wire_5989)
    );

    bfr new_Jinkela_buffer_7825 (
        .din(new_Jinkela_wire_9678),
        .dout(new_Jinkela_wire_9679)
    );

    bfr new_Jinkela_buffer_4404 (
        .din(new_Jinkela_wire_5775),
        .dout(new_Jinkela_wire_5776)
    );

    bfr new_Jinkela_buffer_7943 (
        .din(new_Jinkela_wire_9814),
        .dout(new_Jinkela_wire_9815)
    );

    bfr new_Jinkela_buffer_4444 (
        .din(new_Jinkela_wire_5825),
        .dout(new_Jinkela_wire_5826)
    );

    bfr new_Jinkela_buffer_7826 (
        .din(new_Jinkela_wire_9679),
        .dout(new_Jinkela_wire_9680)
    );

    bfr new_Jinkela_buffer_4405 (
        .din(new_Jinkela_wire_5776),
        .dout(new_Jinkela_wire_5777)
    );

    bfr new_Jinkela_buffer_7874 (
        .din(new_Jinkela_wire_9729),
        .dout(new_Jinkela_wire_9730)
    );

    bfr new_Jinkela_buffer_4501 (
        .din(new_Jinkela_wire_5890),
        .dout(new_Jinkela_wire_5891)
    );

    bfr new_Jinkela_buffer_7827 (
        .din(new_Jinkela_wire_9680),
        .dout(new_Jinkela_wire_9681)
    );

    bfr new_Jinkela_buffer_4406 (
        .din(new_Jinkela_wire_5777),
        .dout(new_Jinkela_wire_5778)
    );

    bfr new_Jinkela_buffer_7895 (
        .din(new_Jinkela_wire_9762),
        .dout(new_Jinkela_wire_9763)
    );

    bfr new_Jinkela_buffer_4445 (
        .din(new_Jinkela_wire_5826),
        .dout(new_Jinkela_wire_5827)
    );

    bfr new_Jinkela_buffer_7828 (
        .din(new_Jinkela_wire_9681),
        .dout(new_Jinkela_wire_9682)
    );

    bfr new_Jinkela_buffer_4407 (
        .din(new_Jinkela_wire_5778),
        .dout(new_Jinkela_wire_5779)
    );

    bfr new_Jinkela_buffer_7875 (
        .din(new_Jinkela_wire_9730),
        .dout(new_Jinkela_wire_9731)
    );

    bfr new_Jinkela_buffer_4577 (
        .din(new_Jinkela_wire_5970),
        .dout(new_Jinkela_wire_5971)
    );

    bfr new_Jinkela_buffer_7829 (
        .din(new_Jinkela_wire_9682),
        .dout(new_Jinkela_wire_9683)
    );

    bfr new_Jinkela_buffer_4408 (
        .din(new_Jinkela_wire_5779),
        .dout(new_Jinkela_wire_5780)
    );

    bfr new_Jinkela_buffer_7987 (
        .din(new_Jinkela_wire_9866),
        .dout(new_Jinkela_wire_9867)
    );

    bfr new_Jinkela_buffer_4446 (
        .din(new_Jinkela_wire_5827),
        .dout(new_Jinkela_wire_5828)
    );

    bfr new_Jinkela_buffer_7830 (
        .din(new_Jinkela_wire_9683),
        .dout(new_Jinkela_wire_9684)
    );

    bfr new_Jinkela_buffer_4409 (
        .din(new_Jinkela_wire_5780),
        .dout(new_Jinkela_wire_5781)
    );

    bfr new_Jinkela_buffer_7876 (
        .din(new_Jinkela_wire_9731),
        .dout(new_Jinkela_wire_9732)
    );

    bfr new_Jinkela_buffer_4502 (
        .din(new_Jinkela_wire_5891),
        .dout(new_Jinkela_wire_5892)
    );

    bfr new_Jinkela_buffer_7831 (
        .din(new_Jinkela_wire_9684),
        .dout(new_Jinkela_wire_9685)
    );

    bfr new_Jinkela_buffer_4410 (
        .din(new_Jinkela_wire_5781),
        .dout(new_Jinkela_wire_5782)
    );

    bfr new_Jinkela_buffer_7896 (
        .din(new_Jinkela_wire_9763),
        .dout(new_Jinkela_wire_9764)
    );

    bfr new_Jinkela_buffer_4447 (
        .din(new_Jinkela_wire_5828),
        .dout(new_Jinkela_wire_5829)
    );

    bfr new_Jinkela_buffer_7832 (
        .din(new_Jinkela_wire_9685),
        .dout(new_Jinkela_wire_9686)
    );

    bfr new_Jinkela_buffer_4411 (
        .din(new_Jinkela_wire_5782),
        .dout(new_Jinkela_wire_5783)
    );

    bfr new_Jinkela_buffer_7877 (
        .din(new_Jinkela_wire_9732),
        .dout(new_Jinkela_wire_9733)
    );

    spl2 new_Jinkela_splitter_548 (
        .a(_0007_),
        .b(new_Jinkela_wire_5991),
        .c(new_Jinkela_wire_5992)
    );

    bfr new_Jinkela_buffer_7833 (
        .din(new_Jinkela_wire_9686),
        .dout(new_Jinkela_wire_9687)
    );

    bfr new_Jinkela_buffer_4412 (
        .din(new_Jinkela_wire_5783),
        .dout(new_Jinkela_wire_5784)
    );

    bfr new_Jinkela_buffer_7944 (
        .din(new_Jinkela_wire_9815),
        .dout(new_Jinkela_wire_9816)
    );

    bfr new_Jinkela_buffer_4448 (
        .din(new_Jinkela_wire_5829),
        .dout(new_Jinkela_wire_5830)
    );

    bfr new_Jinkela_buffer_7834 (
        .din(new_Jinkela_wire_9687),
        .dout(new_Jinkela_wire_9688)
    );

    bfr new_Jinkela_buffer_4413 (
        .din(new_Jinkela_wire_5784),
        .dout(new_Jinkela_wire_5785)
    );

    bfr new_Jinkela_buffer_7878 (
        .din(new_Jinkela_wire_9733),
        .dout(new_Jinkela_wire_9734)
    );

    bfr new_Jinkela_buffer_4503 (
        .din(new_Jinkela_wire_5892),
        .dout(new_Jinkela_wire_5893)
    );

    bfr new_Jinkela_buffer_7835 (
        .din(new_Jinkela_wire_9688),
        .dout(new_Jinkela_wire_9689)
    );

    bfr new_Jinkela_buffer_4414 (
        .din(new_Jinkela_wire_5785),
        .dout(new_Jinkela_wire_5786)
    );

    bfr new_Jinkela_buffer_7897 (
        .din(new_Jinkela_wire_9764),
        .dout(new_Jinkela_wire_9765)
    );

    bfr new_Jinkela_buffer_4449 (
        .din(new_Jinkela_wire_5830),
        .dout(new_Jinkela_wire_5831)
    );

    bfr new_Jinkela_buffer_7836 (
        .din(new_Jinkela_wire_9689),
        .dout(new_Jinkela_wire_9690)
    );

    bfr new_Jinkela_buffer_4415 (
        .din(new_Jinkela_wire_5786),
        .dout(new_Jinkela_wire_5787)
    );

    bfr new_Jinkela_buffer_7879 (
        .din(new_Jinkela_wire_9734),
        .dout(new_Jinkela_wire_9735)
    );

    bfr new_Jinkela_buffer_4578 (
        .din(new_Jinkela_wire_5971),
        .dout(new_Jinkela_wire_5972)
    );

    bfr new_Jinkela_buffer_7837 (
        .din(new_Jinkela_wire_9690),
        .dout(new_Jinkela_wire_9691)
    );

    bfr new_Jinkela_buffer_4416 (
        .din(new_Jinkela_wire_5787),
        .dout(new_Jinkela_wire_5788)
    );

    bfr new_Jinkela_buffer_8176 (
        .din(_0069_),
        .dout(new_Jinkela_wire_10060)
    );

    bfr new_Jinkela_buffer_4450 (
        .din(new_Jinkela_wire_5831),
        .dout(new_Jinkela_wire_5832)
    );

    bfr new_Jinkela_buffer_8027 (
        .din(new_Jinkela_wire_9908),
        .dout(new_Jinkela_wire_9909)
    );

    bfr new_Jinkela_buffer_7838 (
        .din(new_Jinkela_wire_9691),
        .dout(new_Jinkela_wire_9692)
    );

    bfr new_Jinkela_buffer_4417 (
        .din(new_Jinkela_wire_5788),
        .dout(new_Jinkela_wire_5789)
    );

    spl2 new_Jinkela_splitter_777 (
        .a(new_Jinkela_wire_9735),
        .b(new_Jinkela_wire_9736),
        .c(new_Jinkela_wire_9737)
    );

    bfr new_Jinkela_buffer_4504 (
        .din(new_Jinkela_wire_5893),
        .dout(new_Jinkela_wire_5894)
    );

    spl2 new_Jinkela_splitter_776 (
        .a(new_Jinkela_wire_9692),
        .b(new_Jinkela_wire_9693),
        .c(new_Jinkela_wire_9694)
    );

    bfr new_Jinkela_buffer_4418 (
        .din(new_Jinkela_wire_5789),
        .dout(new_Jinkela_wire_5790)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1687),
        .dout(new_Jinkela_wire_1688)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_1511),
        .dout(new_Jinkela_wire_1512)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1663),
        .dout(new_Jinkela_wire_1664)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_1512),
        .dout(new_Jinkela_wire_1513)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(_0455_),
        .b(new_Jinkela_wire_1797),
        .c(new_Jinkela_wire_1798)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_1513),
        .dout(new_Jinkela_wire_1514)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_1664),
        .dout(new_Jinkela_wire_1665)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_1514),
        .dout(new_Jinkela_wire_1515)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1792),
        .dout(new_Jinkela_wire_1793)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1688),
        .dout(new_Jinkela_wire_1689)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_1515),
        .dout(new_Jinkela_wire_1516)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_1665),
        .dout(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1516),
        .dout(new_Jinkela_wire_1517)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_1517),
        .dout(new_Jinkela_wire_1518)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1666),
        .dout(new_Jinkela_wire_1667)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1518),
        .dout(new_Jinkela_wire_1519)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1689),
        .dout(new_Jinkela_wire_1690)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1519),
        .dout(new_Jinkela_wire_1520)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1667),
        .dout(new_Jinkela_wire_1668)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1520),
        .dout(new_Jinkela_wire_1521)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1521),
        .dout(new_Jinkela_wire_1522)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1668),
        .dout(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1522),
        .dout(new_Jinkela_wire_1523)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(_0058_),
        .b(new_Jinkela_wire_1791),
        .c(new_Jinkela_wire_1792)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1690),
        .dout(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1523),
        .dout(new_Jinkela_wire_1524)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1524),
        .dout(new_Jinkela_wire_1525)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1670),
        .dout(new_Jinkela_wire_1671)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_1691),
        .dout(new_Jinkela_wire_1692)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1527),
        .dout(new_Jinkela_wire_1528)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1671),
        .dout(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1528),
        .dout(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1529),
        .dout(new_Jinkela_wire_1530)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1692),
        .dout(new_Jinkela_wire_1693)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1530),
        .dout(new_Jinkela_wire_1531)
    );

    spl2 new_Jinkela_splitter_249 (
        .a(new_Jinkela_wire_1785),
        .b(new_Jinkela_wire_1786),
        .c(new_Jinkela_wire_1787)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1531),
        .dout(new_Jinkela_wire_1532)
    );

    bfr new_Jinkela_buffer_14818 (
        .din(new_Jinkela_wire_17692),
        .dout(new_Jinkela_wire_17693)
    );

    bfr new_Jinkela_buffer_14761 (
        .din(new_Jinkela_wire_17611),
        .dout(new_Jinkela_wire_17612)
    );

    spl2 new_Jinkela_splitter_1288 (
        .a(new_Jinkela_wire_17785),
        .b(new_Jinkela_wire_17786),
        .c(new_Jinkela_wire_17787)
    );

    bfr new_Jinkela_buffer_14762 (
        .din(new_Jinkela_wire_17612),
        .dout(new_Jinkela_wire_17613)
    );

    bfr new_Jinkela_buffer_14819 (
        .din(new_Jinkela_wire_17693),
        .dout(new_Jinkela_wire_17694)
    );

    bfr new_Jinkela_buffer_14763 (
        .din(new_Jinkela_wire_17613),
        .dout(new_Jinkela_wire_17614)
    );

    bfr new_Jinkela_buffer_14854 (
        .din(new_Jinkela_wire_17730),
        .dout(new_Jinkela_wire_17731)
    );

    bfr new_Jinkela_buffer_14764 (
        .din(new_Jinkela_wire_17614),
        .dout(new_Jinkela_wire_17615)
    );

    bfr new_Jinkela_buffer_14820 (
        .din(new_Jinkela_wire_17694),
        .dout(new_Jinkela_wire_17695)
    );

    bfr new_Jinkela_buffer_14765 (
        .din(new_Jinkela_wire_17615),
        .dout(new_Jinkela_wire_17616)
    );

    bfr new_Jinkela_buffer_14912 (
        .din(_1436_),
        .dout(new_Jinkela_wire_17797)
    );

    bfr new_Jinkela_buffer_14766 (
        .din(new_Jinkela_wire_17616),
        .dout(new_Jinkela_wire_17617)
    );

    bfr new_Jinkela_buffer_14821 (
        .din(new_Jinkela_wire_17695),
        .dout(new_Jinkela_wire_17696)
    );

    bfr new_Jinkela_buffer_14767 (
        .din(new_Jinkela_wire_17617),
        .dout(new_Jinkela_wire_17618)
    );

    bfr new_Jinkela_buffer_14855 (
        .din(new_Jinkela_wire_17731),
        .dout(new_Jinkela_wire_17732)
    );

    bfr new_Jinkela_buffer_14768 (
        .din(new_Jinkela_wire_17618),
        .dout(new_Jinkela_wire_17619)
    );

    bfr new_Jinkela_buffer_14822 (
        .din(new_Jinkela_wire_17696),
        .dout(new_Jinkela_wire_17697)
    );

    bfr new_Jinkela_buffer_14769 (
        .din(new_Jinkela_wire_17619),
        .dout(new_Jinkela_wire_17620)
    );

    spl2 new_Jinkela_splitter_1290 (
        .a(_1561_),
        .b(new_Jinkela_wire_17795),
        .c(new_Jinkela_wire_17796)
    );

    bfr new_Jinkela_buffer_14770 (
        .din(new_Jinkela_wire_17620),
        .dout(new_Jinkela_wire_17621)
    );

    bfr new_Jinkela_buffer_14823 (
        .din(new_Jinkela_wire_17697),
        .dout(new_Jinkela_wire_17698)
    );

    bfr new_Jinkela_buffer_14771 (
        .din(new_Jinkela_wire_17621),
        .dout(new_Jinkela_wire_17622)
    );

    bfr new_Jinkela_buffer_14856 (
        .din(new_Jinkela_wire_17732),
        .dout(new_Jinkela_wire_17733)
    );

    bfr new_Jinkela_buffer_14772 (
        .din(new_Jinkela_wire_17622),
        .dout(new_Jinkela_wire_17623)
    );

    bfr new_Jinkela_buffer_14824 (
        .din(new_Jinkela_wire_17698),
        .dout(new_Jinkela_wire_17699)
    );

    bfr new_Jinkela_buffer_14773 (
        .din(new_Jinkela_wire_17623),
        .dout(new_Jinkela_wire_17624)
    );

    bfr new_Jinkela_buffer_14908 (
        .din(new_Jinkela_wire_17790),
        .dout(new_Jinkela_wire_17791)
    );

    bfr new_Jinkela_buffer_14774 (
        .din(new_Jinkela_wire_17624),
        .dout(new_Jinkela_wire_17625)
    );

    bfr new_Jinkela_buffer_14825 (
        .din(new_Jinkela_wire_17699),
        .dout(new_Jinkela_wire_17700)
    );

    bfr new_Jinkela_buffer_14775 (
        .din(new_Jinkela_wire_17625),
        .dout(new_Jinkela_wire_17626)
    );

    bfr new_Jinkela_buffer_14857 (
        .din(new_Jinkela_wire_17733),
        .dout(new_Jinkela_wire_17734)
    );

    bfr new_Jinkela_buffer_14776 (
        .din(new_Jinkela_wire_17626),
        .dout(new_Jinkela_wire_17627)
    );

    bfr new_Jinkela_buffer_14826 (
        .din(new_Jinkela_wire_17700),
        .dout(new_Jinkela_wire_17701)
    );

    bfr new_Jinkela_buffer_14777 (
        .din(new_Jinkela_wire_17627),
        .dout(new_Jinkela_wire_17628)
    );

    spl2 new_Jinkela_splitter_1291 (
        .a(_0291_),
        .b(new_Jinkela_wire_17798),
        .c(new_Jinkela_wire_17799)
    );

    bfr new_Jinkela_buffer_14778 (
        .din(new_Jinkela_wire_17628),
        .dout(new_Jinkela_wire_17629)
    );

    bfr new_Jinkela_buffer_14827 (
        .din(new_Jinkela_wire_17701),
        .dout(new_Jinkela_wire_17702)
    );

    bfr new_Jinkela_buffer_14779 (
        .din(new_Jinkela_wire_17629),
        .dout(new_Jinkela_wire_17630)
    );

    bfr new_Jinkela_buffer_14858 (
        .din(new_Jinkela_wire_17734),
        .dout(new_Jinkela_wire_17735)
    );

    bfr new_Jinkela_buffer_14780 (
        .din(new_Jinkela_wire_17630),
        .dout(new_Jinkela_wire_17631)
    );

    bfr new_Jinkela_buffer_14828 (
        .din(new_Jinkela_wire_17702),
        .dout(new_Jinkela_wire_17703)
    );

    bfr new_Jinkela_buffer_14781 (
        .din(new_Jinkela_wire_17631),
        .dout(new_Jinkela_wire_17632)
    );

    bfr new_Jinkela_buffer_11329 (
        .din(new_Jinkela_wire_13648),
        .dout(new_Jinkela_wire_13649)
    );

    bfr new_Jinkela_buffer_11381 (
        .din(new_Jinkela_wire_13714),
        .dout(new_Jinkela_wire_13715)
    );

    bfr new_Jinkela_buffer_11330 (
        .din(new_Jinkela_wire_13649),
        .dout(new_Jinkela_wire_13650)
    );

    bfr new_Jinkela_buffer_11502 (
        .din(new_Jinkela_wire_13849),
        .dout(new_Jinkela_wire_13850)
    );

    bfr new_Jinkela_buffer_11331 (
        .din(new_Jinkela_wire_13650),
        .dout(new_Jinkela_wire_13651)
    );

    bfr new_Jinkela_buffer_11382 (
        .din(new_Jinkela_wire_13715),
        .dout(new_Jinkela_wire_13716)
    );

    bfr new_Jinkela_buffer_11332 (
        .din(new_Jinkela_wire_13651),
        .dout(new_Jinkela_wire_13652)
    );

    bfr new_Jinkela_buffer_11395 (
        .din(new_Jinkela_wire_13738),
        .dout(new_Jinkela_wire_13739)
    );

    bfr new_Jinkela_buffer_11333 (
        .din(new_Jinkela_wire_13652),
        .dout(new_Jinkela_wire_13653)
    );

    spl2 new_Jinkela_splitter_1016 (
        .a(new_Jinkela_wire_13716),
        .b(new_Jinkela_wire_13717),
        .c(new_Jinkela_wire_13718)
    );

    bfr new_Jinkela_buffer_11334 (
        .din(new_Jinkela_wire_13653),
        .dout(new_Jinkela_wire_13654)
    );

    bfr new_Jinkela_buffer_11396 (
        .din(new_Jinkela_wire_13739),
        .dout(new_Jinkela_wire_13740)
    );

    bfr new_Jinkela_buffer_11335 (
        .din(new_Jinkela_wire_13654),
        .dout(new_Jinkela_wire_13655)
    );

    spl2 new_Jinkela_splitter_1026 (
        .a(_0127_),
        .b(new_Jinkela_wire_13960),
        .c(new_Jinkela_wire_13961)
    );

    bfr new_Jinkela_buffer_11336 (
        .din(new_Jinkela_wire_13655),
        .dout(new_Jinkela_wire_13656)
    );

    bfr new_Jinkela_buffer_11503 (
        .din(new_Jinkela_wire_13850),
        .dout(new_Jinkela_wire_13851)
    );

    bfr new_Jinkela_buffer_11337 (
        .din(new_Jinkela_wire_13656),
        .dout(new_Jinkela_wire_13657)
    );

    bfr new_Jinkela_buffer_11397 (
        .din(new_Jinkela_wire_13740),
        .dout(new_Jinkela_wire_13741)
    );

    bfr new_Jinkela_buffer_11338 (
        .din(new_Jinkela_wire_13657),
        .dout(new_Jinkela_wire_13658)
    );

    spl2 new_Jinkela_splitter_1025 (
        .a(_0285_),
        .b(new_Jinkela_wire_13958),
        .c(new_Jinkela_wire_13959)
    );

    bfr new_Jinkela_buffer_11339 (
        .din(new_Jinkela_wire_13658),
        .dout(new_Jinkela_wire_13659)
    );

    bfr new_Jinkela_buffer_11398 (
        .din(new_Jinkela_wire_13741),
        .dout(new_Jinkela_wire_13742)
    );

    bfr new_Jinkela_buffer_11340 (
        .din(new_Jinkela_wire_13659),
        .dout(new_Jinkela_wire_13660)
    );

    bfr new_Jinkela_buffer_11504 (
        .din(new_Jinkela_wire_13851),
        .dout(new_Jinkela_wire_13852)
    );

    bfr new_Jinkela_buffer_11341 (
        .din(new_Jinkela_wire_13660),
        .dout(new_Jinkela_wire_13661)
    );

    bfr new_Jinkela_buffer_11399 (
        .din(new_Jinkela_wire_13742),
        .dout(new_Jinkela_wire_13743)
    );

    bfr new_Jinkela_buffer_11342 (
        .din(new_Jinkela_wire_13661),
        .dout(new_Jinkela_wire_13662)
    );

    bfr new_Jinkela_buffer_11606 (
        .din(new_Jinkela_wire_13961),
        .dout(new_Jinkela_wire_13962)
    );

    bfr new_Jinkela_buffer_11343 (
        .din(new_Jinkela_wire_13662),
        .dout(new_Jinkela_wire_13663)
    );

    bfr new_Jinkela_buffer_11400 (
        .din(new_Jinkela_wire_13743),
        .dout(new_Jinkela_wire_13744)
    );

    bfr new_Jinkela_buffer_11344 (
        .din(new_Jinkela_wire_13663),
        .dout(new_Jinkela_wire_13664)
    );

    bfr new_Jinkela_buffer_11505 (
        .din(new_Jinkela_wire_13852),
        .dout(new_Jinkela_wire_13853)
    );

    bfr new_Jinkela_buffer_11345 (
        .din(new_Jinkela_wire_13664),
        .dout(new_Jinkela_wire_13665)
    );

    bfr new_Jinkela_buffer_11401 (
        .din(new_Jinkela_wire_13744),
        .dout(new_Jinkela_wire_13745)
    );

    bfr new_Jinkela_buffer_11346 (
        .din(new_Jinkela_wire_13665),
        .dout(new_Jinkela_wire_13666)
    );

    bfr new_Jinkela_buffer_11610 (
        .din(_0049_),
        .dout(new_Jinkela_wire_13966)
    );

    bfr new_Jinkela_buffer_11347 (
        .din(new_Jinkela_wire_13666),
        .dout(new_Jinkela_wire_13667)
    );

    bfr new_Jinkela_buffer_11402 (
        .din(new_Jinkela_wire_13745),
        .dout(new_Jinkela_wire_13746)
    );

    bfr new_Jinkela_buffer_11348 (
        .din(new_Jinkela_wire_13667),
        .dout(new_Jinkela_wire_13668)
    );

    bfr new_Jinkela_buffer_11506 (
        .din(new_Jinkela_wire_13853),
        .dout(new_Jinkela_wire_13854)
    );

    bfr new_Jinkela_buffer_11349 (
        .din(new_Jinkela_wire_13668),
        .dout(new_Jinkela_wire_13669)
    );

    bfr new_Jinkela_buffer_11403 (
        .din(new_Jinkela_wire_13746),
        .dout(new_Jinkela_wire_13747)
    );

    bfr new_Jinkela_buffer_14909 (
        .din(new_Jinkela_wire_17791),
        .dout(new_Jinkela_wire_17792)
    );

    bfr new_Jinkela_buffer_14782 (
        .din(new_Jinkela_wire_17632),
        .dout(new_Jinkela_wire_17633)
    );

    bfr new_Jinkela_buffer_14829 (
        .din(new_Jinkela_wire_17703),
        .dout(new_Jinkela_wire_17704)
    );

    spl2 new_Jinkela_splitter_1274 (
        .a(new_Jinkela_wire_17633),
        .b(new_Jinkela_wire_17634),
        .c(new_Jinkela_wire_17635)
    );

    bfr new_Jinkela_buffer_14830 (
        .din(new_Jinkela_wire_17704),
        .dout(new_Jinkela_wire_17705)
    );

    bfr new_Jinkela_buffer_14859 (
        .din(new_Jinkela_wire_17735),
        .dout(new_Jinkela_wire_17736)
    );

    bfr new_Jinkela_buffer_14913 (
        .din(_0227_),
        .dout(new_Jinkela_wire_17800)
    );

    bfr new_Jinkela_buffer_14831 (
        .din(new_Jinkela_wire_17705),
        .dout(new_Jinkela_wire_17706)
    );

    bfr new_Jinkela_buffer_14860 (
        .din(new_Jinkela_wire_17736),
        .dout(new_Jinkela_wire_17737)
    );

    bfr new_Jinkela_buffer_14832 (
        .din(new_Jinkela_wire_17706),
        .dout(new_Jinkela_wire_17707)
    );

    bfr new_Jinkela_buffer_14910 (
        .din(new_Jinkela_wire_17792),
        .dout(new_Jinkela_wire_17793)
    );

    bfr new_Jinkela_buffer_14833 (
        .din(new_Jinkela_wire_17707),
        .dout(new_Jinkela_wire_17708)
    );

    bfr new_Jinkela_buffer_14861 (
        .din(new_Jinkela_wire_17737),
        .dout(new_Jinkela_wire_17738)
    );

    bfr new_Jinkela_buffer_14834 (
        .din(new_Jinkela_wire_17708),
        .dout(new_Jinkela_wire_17709)
    );

    spl2 new_Jinkela_splitter_1294 (
        .a(_0756_),
        .b(new_Jinkela_wire_17860),
        .c(new_Jinkela_wire_17861)
    );

    bfr new_Jinkela_buffer_14835 (
        .din(new_Jinkela_wire_17709),
        .dout(new_Jinkela_wire_17710)
    );

    bfr new_Jinkela_buffer_14862 (
        .din(new_Jinkela_wire_17738),
        .dout(new_Jinkela_wire_17739)
    );

    bfr new_Jinkela_buffer_14836 (
        .din(new_Jinkela_wire_17710),
        .dout(new_Jinkela_wire_17711)
    );

    spl2 new_Jinkela_splitter_1293 (
        .a(_1019_),
        .b(new_Jinkela_wire_17858),
        .c(new_Jinkela_wire_17859)
    );

    bfr new_Jinkela_buffer_14837 (
        .din(new_Jinkela_wire_17711),
        .dout(new_Jinkela_wire_17712)
    );

    bfr new_Jinkela_buffer_14863 (
        .din(new_Jinkela_wire_17739),
        .dout(new_Jinkela_wire_17740)
    );

    bfr new_Jinkela_buffer_14838 (
        .din(new_Jinkela_wire_17712),
        .dout(new_Jinkela_wire_17713)
    );

    bfr new_Jinkela_buffer_14914 (
        .din(new_Jinkela_wire_17800),
        .dout(new_Jinkela_wire_17801)
    );

    bfr new_Jinkela_buffer_14839 (
        .din(new_Jinkela_wire_17713),
        .dout(new_Jinkela_wire_17714)
    );

    bfr new_Jinkela_buffer_14864 (
        .din(new_Jinkela_wire_17740),
        .dout(new_Jinkela_wire_17741)
    );

    bfr new_Jinkela_buffer_14840 (
        .din(new_Jinkela_wire_17714),
        .dout(new_Jinkela_wire_17715)
    );

    bfr new_Jinkela_buffer_14841 (
        .din(new_Jinkela_wire_17715),
        .dout(new_Jinkela_wire_17716)
    );

    bfr new_Jinkela_buffer_14865 (
        .din(new_Jinkela_wire_17741),
        .dout(new_Jinkela_wire_17742)
    );

    bfr new_Jinkela_buffer_14842 (
        .din(new_Jinkela_wire_17716),
        .dout(new_Jinkela_wire_17717)
    );

    bfr new_Jinkela_buffer_14915 (
        .din(new_Jinkela_wire_17801),
        .dout(new_Jinkela_wire_17802)
    );

    bfr new_Jinkela_buffer_14843 (
        .din(new_Jinkela_wire_17717),
        .dout(new_Jinkela_wire_17718)
    );

    bfr new_Jinkela_buffer_14866 (
        .din(new_Jinkela_wire_17742),
        .dout(new_Jinkela_wire_17743)
    );

    bfr new_Jinkela_buffer_14844 (
        .din(new_Jinkela_wire_17718),
        .dout(new_Jinkela_wire_17719)
    );

    bfr new_Jinkela_buffer_14969 (
        .din(_0657_),
        .dout(new_Jinkela_wire_17864)
    );

    spl2 new_Jinkela_splitter_1295 (
        .a(_1826_),
        .b(new_Jinkela_wire_17862),
        .c(new_Jinkela_wire_17863)
    );

    bfr new_Jinkela_buffer_14845 (
        .din(new_Jinkela_wire_17719),
        .dout(new_Jinkela_wire_17720)
    );

    bfr new_Jinkela_buffer_14867 (
        .din(new_Jinkela_wire_17743),
        .dout(new_Jinkela_wire_17744)
    );

    bfr new_Jinkela_buffer_14846 (
        .din(new_Jinkela_wire_17720),
        .dout(new_Jinkela_wire_17721)
    );

    bfr new_Jinkela_buffer_14916 (
        .din(new_Jinkela_wire_17802),
        .dout(new_Jinkela_wire_17803)
    );

    bfr new_Jinkela_buffer_14847 (
        .din(new_Jinkela_wire_17721),
        .dout(new_Jinkela_wire_17722)
    );

    bfr new_Jinkela_buffer_14868 (
        .din(new_Jinkela_wire_17744),
        .dout(new_Jinkela_wire_17745)
    );

    bfr new_Jinkela_buffer_14848 (
        .din(new_Jinkela_wire_17722),
        .dout(new_Jinkela_wire_17723)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1693),
        .dout(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1532),
        .dout(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1533),
        .dout(new_Jinkela_wire_1534)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1694),
        .dout(new_Jinkela_wire_1695)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(_1222_),
        .b(new_Jinkela_wire_1803),
        .c(new_Jinkela_wire_1804)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1695),
        .dout(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1536),
        .dout(new_Jinkela_wire_1537)
    );

    bfr new_Jinkela_buffer_988 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1537),
        .dout(new_Jinkela_wire_1538)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1696),
        .dout(new_Jinkela_wire_1697)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1538),
        .dout(new_Jinkela_wire_1539)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1798),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1539),
        .dout(new_Jinkela_wire_1540)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(_1060_),
        .b(new_Jinkela_wire_1805),
        .c(new_Jinkela_wire_1806)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1697),
        .dout(new_Jinkela_wire_1698)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_1540),
        .dout(new_Jinkela_wire_1541)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1794),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1541),
        .dout(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1698),
        .dout(new_Jinkela_wire_1699)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1542),
        .dout(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1806),
        .dout(new_Jinkela_wire_1807)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_1543),
        .dout(new_Jinkela_wire_1544)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1699),
        .dout(new_Jinkela_wire_1700)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1544),
        .dout(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1795),
        .dout(new_Jinkela_wire_1796)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1545),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1700),
        .dout(new_Jinkela_wire_1701)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1701),
        .dout(new_Jinkela_wire_1702)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1549),
        .dout(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_999 (
        .din(_1357_),
        .dout(new_Jinkela_wire_1811)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_1702),
        .dout(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1551),
        .dout(new_Jinkela_wire_1552)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1703),
        .dout(new_Jinkela_wire_1704)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1552),
        .dout(new_Jinkela_wire_1553)
    );

    bfr new_Jinkela_buffer_11350 (
        .din(new_Jinkela_wire_13669),
        .dout(new_Jinkela_wire_13670)
    );

    spl2 new_Jinkela_splitter_1027 (
        .a(_1642_),
        .b(new_Jinkela_wire_13967),
        .c(new_Jinkela_wire_13968)
    );

    bfr new_Jinkela_buffer_11351 (
        .din(new_Jinkela_wire_13670),
        .dout(new_Jinkela_wire_13671)
    );

    bfr new_Jinkela_buffer_11404 (
        .din(new_Jinkela_wire_13747),
        .dout(new_Jinkela_wire_13748)
    );

    bfr new_Jinkela_buffer_11352 (
        .din(new_Jinkela_wire_13671),
        .dout(new_Jinkela_wire_13672)
    );

    bfr new_Jinkela_buffer_11507 (
        .din(new_Jinkela_wire_13854),
        .dout(new_Jinkela_wire_13855)
    );

    spl2 new_Jinkela_splitter_1009 (
        .a(new_Jinkela_wire_13672),
        .b(new_Jinkela_wire_13673),
        .c(new_Jinkela_wire_13674)
    );

    bfr new_Jinkela_buffer_11611 (
        .din(_0003_),
        .dout(new_Jinkela_wire_13969)
    );

    spl2 new_Jinkela_splitter_1029 (
        .a(_1243_),
        .b(new_Jinkela_wire_13972),
        .c(new_Jinkela_wire_13973)
    );

    bfr new_Jinkela_buffer_11405 (
        .din(new_Jinkela_wire_13748),
        .dout(new_Jinkela_wire_13749)
    );

    bfr new_Jinkela_buffer_11406 (
        .din(new_Jinkela_wire_13749),
        .dout(new_Jinkela_wire_13750)
    );

    bfr new_Jinkela_buffer_11508 (
        .din(new_Jinkela_wire_13855),
        .dout(new_Jinkela_wire_13856)
    );

    bfr new_Jinkela_buffer_11407 (
        .din(new_Jinkela_wire_13750),
        .dout(new_Jinkela_wire_13751)
    );

    bfr new_Jinkela_buffer_11607 (
        .din(new_Jinkela_wire_13962),
        .dout(new_Jinkela_wire_13963)
    );

    bfr new_Jinkela_buffer_11408 (
        .din(new_Jinkela_wire_13751),
        .dout(new_Jinkela_wire_13752)
    );

    bfr new_Jinkela_buffer_11509 (
        .din(new_Jinkela_wire_13856),
        .dout(new_Jinkela_wire_13857)
    );

    bfr new_Jinkela_buffer_11409 (
        .din(new_Jinkela_wire_13752),
        .dout(new_Jinkela_wire_13753)
    );

    bfr new_Jinkela_buffer_11410 (
        .din(new_Jinkela_wire_13753),
        .dout(new_Jinkela_wire_13754)
    );

    bfr new_Jinkela_buffer_11510 (
        .din(new_Jinkela_wire_13857),
        .dout(new_Jinkela_wire_13858)
    );

    bfr new_Jinkela_buffer_11411 (
        .din(new_Jinkela_wire_13754),
        .dout(new_Jinkela_wire_13755)
    );

    bfr new_Jinkela_buffer_11608 (
        .din(new_Jinkela_wire_13963),
        .dout(new_Jinkela_wire_13964)
    );

    bfr new_Jinkela_buffer_11412 (
        .din(new_Jinkela_wire_13755),
        .dout(new_Jinkela_wire_13756)
    );

    bfr new_Jinkela_buffer_11511 (
        .din(new_Jinkela_wire_13858),
        .dout(new_Jinkela_wire_13859)
    );

    bfr new_Jinkela_buffer_11413 (
        .din(new_Jinkela_wire_13756),
        .dout(new_Jinkela_wire_13757)
    );

    spl2 new_Jinkela_splitter_1028 (
        .a(_1550_),
        .b(new_Jinkela_wire_13970),
        .c(new_Jinkela_wire_13971)
    );

    bfr new_Jinkela_buffer_11414 (
        .din(new_Jinkela_wire_13757),
        .dout(new_Jinkela_wire_13758)
    );

    bfr new_Jinkela_buffer_11512 (
        .din(new_Jinkela_wire_13859),
        .dout(new_Jinkela_wire_13860)
    );

    bfr new_Jinkela_buffer_11415 (
        .din(new_Jinkela_wire_13758),
        .dout(new_Jinkela_wire_13759)
    );

    bfr new_Jinkela_buffer_11609 (
        .din(new_Jinkela_wire_13964),
        .dout(new_Jinkela_wire_13965)
    );

    bfr new_Jinkela_buffer_11416 (
        .din(new_Jinkela_wire_13759),
        .dout(new_Jinkela_wire_13760)
    );

    bfr new_Jinkela_buffer_11513 (
        .din(new_Jinkela_wire_13860),
        .dout(new_Jinkela_wire_13861)
    );

    bfr new_Jinkela_buffer_11417 (
        .din(new_Jinkela_wire_13760),
        .dout(new_Jinkela_wire_13761)
    );

    bfr new_Jinkela_buffer_11418 (
        .din(new_Jinkela_wire_13761),
        .dout(new_Jinkela_wire_13762)
    );

    bfr new_Jinkela_buffer_11514 (
        .din(new_Jinkela_wire_13861),
        .dout(new_Jinkela_wire_13862)
    );

    bfr new_Jinkela_buffer_11419 (
        .din(new_Jinkela_wire_13762),
        .dout(new_Jinkela_wire_13763)
    );

    bfr new_Jinkela_buffer_11616 (
        .din(_1802_),
        .dout(new_Jinkela_wire_13978)
    );

    bfr new_Jinkela_buffer_11420 (
        .din(new_Jinkela_wire_13763),
        .dout(new_Jinkela_wire_13764)
    );

    bfr new_Jinkela_buffer_11515 (
        .din(new_Jinkela_wire_13862),
        .dout(new_Jinkela_wire_13863)
    );

    bfr new_Jinkela_buffer_11421 (
        .din(new_Jinkela_wire_13764),
        .dout(new_Jinkela_wire_13765)
    );

    bfr new_Jinkela_buffer_11612 (
        .din(new_Jinkela_wire_13973),
        .dout(new_Jinkela_wire_13974)
    );

    bfr new_Jinkela_buffer_11422 (
        .din(new_Jinkela_wire_13765),
        .dout(new_Jinkela_wire_13766)
    );

    bfr new_Jinkela_buffer_4451 (
        .din(new_Jinkela_wire_5832),
        .dout(new_Jinkela_wire_5833)
    );

    bfr new_Jinkela_buffer_7898 (
        .din(new_Jinkela_wire_9765),
        .dout(new_Jinkela_wire_9766)
    );

    bfr new_Jinkela_buffer_4419 (
        .din(new_Jinkela_wire_5790),
        .dout(new_Jinkela_wire_5791)
    );

    bfr new_Jinkela_buffer_7945 (
        .din(new_Jinkela_wire_9816),
        .dout(new_Jinkela_wire_9817)
    );

    spl2 new_Jinkela_splitter_549 (
        .a(_1696_),
        .b(new_Jinkela_wire_5993),
        .c(new_Jinkela_wire_5994)
    );

    bfr new_Jinkela_buffer_7899 (
        .din(new_Jinkela_wire_9766),
        .dout(new_Jinkela_wire_9767)
    );

    bfr new_Jinkela_buffer_4420 (
        .din(new_Jinkela_wire_5791),
        .dout(new_Jinkela_wire_5792)
    );

    bfr new_Jinkela_buffer_7988 (
        .din(new_Jinkela_wire_9867),
        .dout(new_Jinkela_wire_9868)
    );

    bfr new_Jinkela_buffer_4452 (
        .din(new_Jinkela_wire_5833),
        .dout(new_Jinkela_wire_5834)
    );

    bfr new_Jinkela_buffer_7900 (
        .din(new_Jinkela_wire_9767),
        .dout(new_Jinkela_wire_9768)
    );

    bfr new_Jinkela_buffer_4421 (
        .din(new_Jinkela_wire_5792),
        .dout(new_Jinkela_wire_5793)
    );

    bfr new_Jinkela_buffer_7946 (
        .din(new_Jinkela_wire_9817),
        .dout(new_Jinkela_wire_9818)
    );

    bfr new_Jinkela_buffer_4505 (
        .din(new_Jinkela_wire_5894),
        .dout(new_Jinkela_wire_5895)
    );

    bfr new_Jinkela_buffer_7901 (
        .din(new_Jinkela_wire_9768),
        .dout(new_Jinkela_wire_9769)
    );

    bfr new_Jinkela_buffer_4422 (
        .din(new_Jinkela_wire_5793),
        .dout(new_Jinkela_wire_5794)
    );

    bfr new_Jinkela_buffer_4453 (
        .din(new_Jinkela_wire_5834),
        .dout(new_Jinkela_wire_5835)
    );

    bfr new_Jinkela_buffer_7902 (
        .din(new_Jinkela_wire_9769),
        .dout(new_Jinkela_wire_9770)
    );

    bfr new_Jinkela_buffer_4423 (
        .din(new_Jinkela_wire_5794),
        .dout(new_Jinkela_wire_5795)
    );

    bfr new_Jinkela_buffer_7947 (
        .din(new_Jinkela_wire_9818),
        .dout(new_Jinkela_wire_9819)
    );

    bfr new_Jinkela_buffer_4579 (
        .din(new_Jinkela_wire_5972),
        .dout(new_Jinkela_wire_5973)
    );

    bfr new_Jinkela_buffer_7903 (
        .din(new_Jinkela_wire_9770),
        .dout(new_Jinkela_wire_9771)
    );

    bfr new_Jinkela_buffer_4424 (
        .din(new_Jinkela_wire_5795),
        .dout(new_Jinkela_wire_5796)
    );

    bfr new_Jinkela_buffer_7989 (
        .din(new_Jinkela_wire_9868),
        .dout(new_Jinkela_wire_9869)
    );

    bfr new_Jinkela_buffer_4454 (
        .din(new_Jinkela_wire_5835),
        .dout(new_Jinkela_wire_5836)
    );

    bfr new_Jinkela_buffer_7904 (
        .din(new_Jinkela_wire_9771),
        .dout(new_Jinkela_wire_9772)
    );

    bfr new_Jinkela_buffer_4425 (
        .din(new_Jinkela_wire_5796),
        .dout(new_Jinkela_wire_5797)
    );

    bfr new_Jinkela_buffer_7948 (
        .din(new_Jinkela_wire_9819),
        .dout(new_Jinkela_wire_9820)
    );

    bfr new_Jinkela_buffer_4506 (
        .din(new_Jinkela_wire_5895),
        .dout(new_Jinkela_wire_5896)
    );

    bfr new_Jinkela_buffer_7905 (
        .din(new_Jinkela_wire_9772),
        .dout(new_Jinkela_wire_9773)
    );

    spl2 new_Jinkela_splitter_535 (
        .a(new_Jinkela_wire_5797),
        .b(new_Jinkela_wire_5798),
        .c(new_Jinkela_wire_5799)
    );

    bfr new_Jinkela_buffer_8028 (
        .din(new_Jinkela_wire_9909),
        .dout(new_Jinkela_wire_9910)
    );

    bfr new_Jinkela_buffer_7906 (
        .din(new_Jinkela_wire_9773),
        .dout(new_Jinkela_wire_9774)
    );

    bfr new_Jinkela_buffer_4455 (
        .din(new_Jinkela_wire_5836),
        .dout(new_Jinkela_wire_5837)
    );

    bfr new_Jinkela_buffer_7949 (
        .din(new_Jinkela_wire_9820),
        .dout(new_Jinkela_wire_9821)
    );

    bfr new_Jinkela_buffer_4456 (
        .din(new_Jinkela_wire_5837),
        .dout(new_Jinkela_wire_5838)
    );

    bfr new_Jinkela_buffer_7907 (
        .din(new_Jinkela_wire_9774),
        .dout(new_Jinkela_wire_9775)
    );

    bfr new_Jinkela_buffer_4507 (
        .din(new_Jinkela_wire_5896),
        .dout(new_Jinkela_wire_5897)
    );

    bfr new_Jinkela_buffer_7990 (
        .din(new_Jinkela_wire_9869),
        .dout(new_Jinkela_wire_9870)
    );

    bfr new_Jinkela_buffer_4457 (
        .din(new_Jinkela_wire_5838),
        .dout(new_Jinkela_wire_5839)
    );

    bfr new_Jinkela_buffer_7908 (
        .din(new_Jinkela_wire_9775),
        .dout(new_Jinkela_wire_9776)
    );

    bfr new_Jinkela_buffer_4580 (
        .din(new_Jinkela_wire_5973),
        .dout(new_Jinkela_wire_5974)
    );

    bfr new_Jinkela_buffer_7950 (
        .din(new_Jinkela_wire_9821),
        .dout(new_Jinkela_wire_9822)
    );

    bfr new_Jinkela_buffer_4458 (
        .din(new_Jinkela_wire_5839),
        .dout(new_Jinkela_wire_5840)
    );

    bfr new_Jinkela_buffer_7909 (
        .din(new_Jinkela_wire_9776),
        .dout(new_Jinkela_wire_9777)
    );

    bfr new_Jinkela_buffer_4508 (
        .din(new_Jinkela_wire_5897),
        .dout(new_Jinkela_wire_5898)
    );

    bfr new_Jinkela_buffer_8177 (
        .din(_1226_),
        .dout(new_Jinkela_wire_10061)
    );

    bfr new_Jinkela_buffer_4459 (
        .din(new_Jinkela_wire_5840),
        .dout(new_Jinkela_wire_5841)
    );

    bfr new_Jinkela_buffer_7910 (
        .din(new_Jinkela_wire_9777),
        .dout(new_Jinkela_wire_9778)
    );

    bfr new_Jinkela_buffer_7951 (
        .din(new_Jinkela_wire_9822),
        .dout(new_Jinkela_wire_9823)
    );

    spl2 new_Jinkela_splitter_550 (
        .a(_1157_),
        .b(new_Jinkela_wire_5995),
        .c(new_Jinkela_wire_5996)
    );

    bfr new_Jinkela_buffer_4460 (
        .din(new_Jinkela_wire_5841),
        .dout(new_Jinkela_wire_5842)
    );

    bfr new_Jinkela_buffer_7911 (
        .din(new_Jinkela_wire_9778),
        .dout(new_Jinkela_wire_9779)
    );

    bfr new_Jinkela_buffer_4509 (
        .din(new_Jinkela_wire_5898),
        .dout(new_Jinkela_wire_5899)
    );

    bfr new_Jinkela_buffer_7991 (
        .din(new_Jinkela_wire_9870),
        .dout(new_Jinkela_wire_9871)
    );

    bfr new_Jinkela_buffer_4461 (
        .din(new_Jinkela_wire_5842),
        .dout(new_Jinkela_wire_5843)
    );

    bfr new_Jinkela_buffer_7912 (
        .din(new_Jinkela_wire_9779),
        .dout(new_Jinkela_wire_9780)
    );

    bfr new_Jinkela_buffer_4581 (
        .din(new_Jinkela_wire_5974),
        .dout(new_Jinkela_wire_5975)
    );

    bfr new_Jinkela_buffer_7952 (
        .din(new_Jinkela_wire_9823),
        .dout(new_Jinkela_wire_9824)
    );

    bfr new_Jinkela_buffer_4462 (
        .din(new_Jinkela_wire_5843),
        .dout(new_Jinkela_wire_5844)
    );

    bfr new_Jinkela_buffer_7913 (
        .din(new_Jinkela_wire_9780),
        .dout(new_Jinkela_wire_9781)
    );

    bfr new_Jinkela_buffer_4510 (
        .din(new_Jinkela_wire_5899),
        .dout(new_Jinkela_wire_5900)
    );

    bfr new_Jinkela_buffer_8167 (
        .din(new_Jinkela_wire_10048),
        .dout(new_Jinkela_wire_10049)
    );

    bfr new_Jinkela_buffer_8029 (
        .din(new_Jinkela_wire_9910),
        .dout(new_Jinkela_wire_9911)
    );

    bfr new_Jinkela_buffer_4463 (
        .din(new_Jinkela_wire_5844),
        .dout(new_Jinkela_wire_5845)
    );

    bfr new_Jinkela_buffer_7914 (
        .din(new_Jinkela_wire_9781),
        .dout(new_Jinkela_wire_9782)
    );

    spl2 new_Jinkela_splitter_551 (
        .a(_0074_),
        .b(new_Jinkela_wire_5999),
        .c(new_Jinkela_wire_6000)
    );

    bfr new_Jinkela_buffer_7953 (
        .din(new_Jinkela_wire_9824),
        .dout(new_Jinkela_wire_9825)
    );

    bfr new_Jinkela_buffer_4593 (
        .din(_0693_),
        .dout(new_Jinkela_wire_5997)
    );

    bfr new_Jinkela_buffer_4464 (
        .din(new_Jinkela_wire_5845),
        .dout(new_Jinkela_wire_5846)
    );

    bfr new_Jinkela_buffer_7915 (
        .din(new_Jinkela_wire_9782),
        .dout(new_Jinkela_wire_9783)
    );

    bfr new_Jinkela_buffer_4511 (
        .din(new_Jinkela_wire_5900),
        .dout(new_Jinkela_wire_5901)
    );

    bfr new_Jinkela_buffer_7992 (
        .din(new_Jinkela_wire_9871),
        .dout(new_Jinkela_wire_9872)
    );

    bfr new_Jinkela_buffer_4465 (
        .din(new_Jinkela_wire_5846),
        .dout(new_Jinkela_wire_5847)
    );

    bfr new_Jinkela_buffer_7916 (
        .din(new_Jinkela_wire_9783),
        .dout(new_Jinkela_wire_9784)
    );

    bfr new_Jinkela_buffer_4582 (
        .din(new_Jinkela_wire_5975),
        .dout(new_Jinkela_wire_5976)
    );

    bfr new_Jinkela_buffer_7954 (
        .din(new_Jinkela_wire_9825),
        .dout(new_Jinkela_wire_9826)
    );

    bfr new_Jinkela_buffer_4466 (
        .din(new_Jinkela_wire_5847),
        .dout(new_Jinkela_wire_5848)
    );

    bfr new_Jinkela_buffer_7917 (
        .din(new_Jinkela_wire_9784),
        .dout(new_Jinkela_wire_9785)
    );

    bfr new_Jinkela_buffer_4512 (
        .din(new_Jinkela_wire_5901),
        .dout(new_Jinkela_wire_5902)
    );

    bfr new_Jinkela_buffer_4467 (
        .din(new_Jinkela_wire_5848),
        .dout(new_Jinkela_wire_5849)
    );

    bfr new_Jinkela_buffer_7918 (
        .din(new_Jinkela_wire_9785),
        .dout(new_Jinkela_wire_9786)
    );

    bfr new_Jinkela_buffer_7955 (
        .din(new_Jinkela_wire_9826),
        .dout(new_Jinkela_wire_9827)
    );

    bfr new_Jinkela_buffer_4594 (
        .din(_1315_),
        .dout(new_Jinkela_wire_5998)
    );

endmodule
