module sorter48(a, b);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input a_8_;
  input a_9_;
  input a_10_;
  input a_11_;
  input a_12_;
  input a_13_;
  input a_14_;
  input a_15_;
  input a_16_;
  input a_17_;
  input a_18_;
  input a_19_;
  input a_20_;
  input a_21_;
  input a_22_;
  input a_23_;
  input a_24_;
  input a_25_;
  input a_26_;
  input a_27_;
  input a_28_;
  input a_29_;
  input a_30_;
  input a_31_;
  input a_32_;
  input a_33_;
  input a_34_;
  input a_35_;
  input a_36_;
  input a_37_;
  input a_38_;
  input a_39_;
  input a_40_;
  input a_41_;
  input a_42_;
  input a_43_;
  input a_44_;
  input a_45_;
  input a_46_;
  input a_47_;
  output b_0_;
  output b_1_;
  output b_2_;
  output b_3_;
  output b_4_;
  output b_5_;
  output b_6_;
  output b_7_;
  output b_8_;
  output b_9_;
  output b_10_;
  output b_11_;
  output b_12_;
  output b_13_;
  output b_14_;
  output b_15_;
  output b_16_;
  output b_17_;
  output b_18_;
  output b_19_;
  output b_20_;
  output b_21_;
  output b_22_;
  output b_23_;
  output b_24_;
  output b_25_;
  output b_26_;
  output b_27_;
  output b_28_;
  output b_29_;
  output b_30_;
  output b_31_;
  output b_32_;
  output b_33_;
  output b_34_;
  output b_35_;
  output b_36_;
  output b_37_;
  output b_38_;
  output b_39_;
  output b_40_;
  output b_41_;
  output b_42_;
  output b_43_;
  output b_44_;
  output b_45_;
  output b_46_;
  output b_47_;
  wire c_0_;
  wire c_1_;
  wire c_2_;
  wire c_3_;
  wire c_4_;
  wire c_5_;
  wire c_6_;
  wire c_7_;
  wire c_8_;
  wire c_9_;
  wire c_10_;
  wire c_11_;
  wire c_12_;
  wire c_13_;
  wire c_14_;
  wire c_15_;
  wire c_16_;
  wire c_17_;
  wire c_18_;
  wire c_19_;
  wire c_20_;
  wire c_21_;
  wire c_22_;
  wire c_23_;
  wire c_24_;
  wire c_25_;
  wire c_26_;
  wire c_27_;
  wire c_28_;
  wire c_29_;
  wire c_30_;
  wire c_31_;
  wire c_32_;
  wire c_33_;
  wire c_34_;
  wire c_35_;
  wire c_36_;
  wire c_37_;
  wire c_38_;
  wire c_39_;
  wire c_40_;
  wire c_41_;
  wire c_42_;
  wire c_43_;
  wire c_44_;
  wire c_45_;
  wire c_46_;
  wire c_47_;
  wire _g_0_c_0_;
  wire _g_0_c_1_;
  wire _g_0_c_2_;
  wire _g_0_c_3_;
  wire _g_0_c_4_;
  wire _g_0_c_5_;
  wire _g_0_c_6_;
  wire _g_0_c_7_;
  wire _g_0_c_8_;
  wire _g_0_c_9_;
  wire _g_0_c_10_;
  wire _g_0_c_11_;
  wire _g_0_c_12_;
  wire _g_0_c_13_;
  wire _g_0_c_14_;
  wire _g_0_c_15_;
  wire _g_0_c_16_;
  wire _g_0_c_17_;
  wire _g_0_c_18_;
  wire _g_0_c_19_;
  wire _g_0_c_20_;
  wire _g_0_c_21_;
  wire _g_0_c_22_;
  wire _g_0_c_23_;
  wire _g_0_g_0_c_0_;
  wire _g_0_g_0_c_1_;
  wire _g_0_g_0_c_2_;
  wire _g_0_g_0_c_3_;
  wire _g_0_g_0_c_4_;
  wire _g_0_g_0_c_5_;
  wire _g_0_g_0_c_6_;
  wire _g_0_g_0_c_7_;
  wire _g_0_g_0_c_8_;
  wire _g_0_g_0_c_9_;
  wire _g_0_g_0_c_10_;
  wire _g_0_g_0_c_11_;
  wire _g_0_g_0_g_0_c_0_;
  wire _g_0_g_0_g_0_c_1_;
  wire _g_0_g_0_g_0_c_2_;
  wire _g_0_g_0_g_0_c_3_;
  wire _g_0_g_0_g_0_c_4_;
  wire _g_0_g_0_g_0_c_5_;
  wire _g_0_g_0_g_0_g_3_c_0_;
  wire _g_0_g_0_g_0_g_3_c_1_;
  wire _g_0_g_0_g_0_g_3_c_2_;
  wire _g_0_g_0_g_0_g_3_c_3_;
  wire _g_0_g_0_g_0_g_3_c_4_;
  wire _g_0_g_0_g_0_g_3_c_5_;
  wire _g_0_g_0_g_1_c_0_;
  wire _g_0_g_0_g_1_c_1_;
  wire _g_0_g_0_g_1_c_2_;
  wire _g_0_g_0_g_1_c_3_;
  wire _g_0_g_0_g_1_c_4_;
  wire _g_0_g_0_g_1_c_5_;
  wire _g_0_g_0_g_1_g_3_c_0_;
  wire _g_0_g_0_g_1_g_3_c_1_;
  wire _g_0_g_0_g_1_g_3_c_2_;
  wire _g_0_g_0_g_1_g_3_c_3_;
  wire _g_0_g_0_g_1_g_3_c_4_;
  wire _g_0_g_0_g_1_g_3_c_5_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_0_g_1_c_0_;
  wire _g_0_g_1_c_1_;
  wire _g_0_g_1_c_2_;
  wire _g_0_g_1_c_3_;
  wire _g_0_g_1_c_4_;
  wire _g_0_g_1_c_5_;
  wire _g_0_g_1_c_6_;
  wire _g_0_g_1_c_7_;
  wire _g_0_g_1_c_8_;
  wire _g_0_g_1_c_9_;
  wire _g_0_g_1_c_10_;
  wire _g_0_g_1_c_11_;
  wire _g_0_g_1_g_0_c_0_;
  wire _g_0_g_1_g_0_c_1_;
  wire _g_0_g_1_g_0_c_2_;
  wire _g_0_g_1_g_0_c_3_;
  wire _g_0_g_1_g_0_c_4_;
  wire _g_0_g_1_g_0_c_5_;
  wire _g_0_g_1_g_0_g_3_c_0_;
  wire _g_0_g_1_g_0_g_3_c_1_;
  wire _g_0_g_1_g_0_g_3_c_2_;
  wire _g_0_g_1_g_0_g_3_c_3_;
  wire _g_0_g_1_g_0_g_3_c_4_;
  wire _g_0_g_1_g_0_g_3_c_5_;
  wire _g_0_g_1_g_1_c_0_;
  wire _g_0_g_1_g_1_c_1_;
  wire _g_0_g_1_g_1_c_2_;
  wire _g_0_g_1_g_1_c_3_;
  wire _g_0_g_1_g_1_c_4_;
  wire _g_0_g_1_g_1_c_5_;
  wire _g_0_g_1_g_1_g_3_c_0_;
  wire _g_0_g_1_g_1_g_3_c_1_;
  wire _g_0_g_1_g_1_g_3_c_2_;
  wire _g_0_g_1_g_1_g_3_c_3_;
  wire _g_0_g_1_g_1_g_3_c_4_;
  wire _g_0_g_1_g_1_g_3_c_5_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_1_c_0_;
  wire _g_1_c_1_;
  wire _g_1_c_2_;
  wire _g_1_c_3_;
  wire _g_1_c_4_;
  wire _g_1_c_5_;
  wire _g_1_c_6_;
  wire _g_1_c_7_;
  wire _g_1_c_8_;
  wire _g_1_c_9_;
  wire _g_1_c_10_;
  wire _g_1_c_11_;
  wire _g_1_c_12_;
  wire _g_1_c_13_;
  wire _g_1_c_14_;
  wire _g_1_c_15_;
  wire _g_1_c_16_;
  wire _g_1_c_17_;
  wire _g_1_c_18_;
  wire _g_1_c_19_;
  wire _g_1_c_20_;
  wire _g_1_c_21_;
  wire _g_1_c_22_;
  wire _g_1_c_23_;
  wire _g_1_g_0_c_0_;
  wire _g_1_g_0_c_1_;
  wire _g_1_g_0_c_2_;
  wire _g_1_g_0_c_3_;
  wire _g_1_g_0_c_4_;
  wire _g_1_g_0_c_5_;
  wire _g_1_g_0_c_6_;
  wire _g_1_g_0_c_7_;
  wire _g_1_g_0_c_8_;
  wire _g_1_g_0_c_9_;
  wire _g_1_g_0_c_10_;
  wire _g_1_g_0_c_11_;
  wire _g_1_g_0_g_0_c_0_;
  wire _g_1_g_0_g_0_c_1_;
  wire _g_1_g_0_g_0_c_2_;
  wire _g_1_g_0_g_0_c_3_;
  wire _g_1_g_0_g_0_c_4_;
  wire _g_1_g_0_g_0_c_5_;
  wire _g_1_g_0_g_0_g_3_c_0_;
  wire _g_1_g_0_g_0_g_3_c_1_;
  wire _g_1_g_0_g_0_g_3_c_2_;
  wire _g_1_g_0_g_0_g_3_c_3_;
  wire _g_1_g_0_g_0_g_3_c_4_;
  wire _g_1_g_0_g_0_g_3_c_5_;
  wire _g_1_g_0_g_1_c_0_;
  wire _g_1_g_0_g_1_c_1_;
  wire _g_1_g_0_g_1_c_2_;
  wire _g_1_g_0_g_1_c_3_;
  wire _g_1_g_0_g_1_c_4_;
  wire _g_1_g_0_g_1_c_5_;
  wire _g_1_g_0_g_1_g_3_c_0_;
  wire _g_1_g_0_g_1_g_3_c_1_;
  wire _g_1_g_0_g_1_g_3_c_2_;
  wire _g_1_g_0_g_1_g_3_c_3_;
  wire _g_1_g_0_g_1_g_3_c_4_;
  wire _g_1_g_0_g_1_g_3_c_5_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_1_g_1_c_0_;
  wire _g_1_g_1_c_1_;
  wire _g_1_g_1_c_2_;
  wire _g_1_g_1_c_3_;
  wire _g_1_g_1_c_4_;
  wire _g_1_g_1_c_5_;
  wire _g_1_g_1_c_6_;
  wire _g_1_g_1_c_7_;
  wire _g_1_g_1_c_8_;
  wire _g_1_g_1_c_9_;
  wire _g_1_g_1_c_10_;
  wire _g_1_g_1_c_11_;
  wire _g_1_g_1_g_0_c_0_;
  wire _g_1_g_1_g_0_c_1_;
  wire _g_1_g_1_g_0_c_2_;
  wire _g_1_g_1_g_0_c_3_;
  wire _g_1_g_1_g_0_c_4_;
  wire _g_1_g_1_g_0_c_5_;
  wire _g_1_g_1_g_0_g_3_c_0_;
  wire _g_1_g_1_g_0_g_3_c_1_;
  wire _g_1_g_1_g_0_g_3_c_2_;
  wire _g_1_g_1_g_0_g_3_c_3_;
  wire _g_1_g_1_g_0_g_3_c_4_;
  wire _g_1_g_1_g_0_g_3_c_5_;
  wire _g_1_g_1_g_1_c_0_;
  wire _g_1_g_1_g_1_c_1_;
  wire _g_1_g_1_g_1_c_2_;
  wire _g_1_g_1_g_1_c_3_;
  wire _g_1_g_1_g_1_c_4_;
  wire _g_1_g_1_g_1_c_5_;
  wire _g_1_g_1_g_1_g_3_c_0_;
  wire _g_1_g_1_g_1_g_3_c_1_;
  wire _g_1_g_1_g_1_g_3_c_2_;
  wire _g_1_g_1_g_1_g_3_c_3_;
  wire _g_1_g_1_g_1_g_3_c_4_;
  wire _g_1_g_1_g_1_g_3_c_5_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_10_23_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_23_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_24_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_24_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_25_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_25_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_26_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_26_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_27_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_27_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_28_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_28_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_29_6__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_29_6__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_30_7__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_30_7__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_31_8__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_31_8__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_32_9__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_32_9__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_33_10__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_33_10__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_34_11__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_34_11__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_35_12__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_35_12__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_36_13__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_36_13__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_37_14__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_37_14__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_38_15__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_38_15__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_39_16__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_39_16__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_40_17__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_40_17__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_41_18__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_41_18__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_42_19__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_42_19__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_43_20__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_43_20__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_44_21__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_44_21__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_45_22__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_45_22__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_10_46_23__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_10_46_23__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_;
  wire _m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_;
  or_bb _0160_ (
    .a(a_46_),
    .b(a_47_),
    .c(_0001_)
  );
  or_bb _0161_ (
    .a(_0001_),
    .b(a_45_),
    .c(_g_0_g_0_g_0_c_5_)
  );
  maj_bbb _0162_ (
    .a(a_45_),
    .b(a_46_),
    .c(a_47_),
    .d(_g_0_g_0_g_0_c_4_)
  );
  and_bb _0163_ (
    .a(a_46_),
    .b(a_47_),
    .c(_0000_)
  );
  and_bb _0164_ (
    .a(_0000_),
    .b(a_45_),
    .c(_g_0_g_0_g_0_c_3_)
  );
  or_bb _0165_ (
    .a(a_43_),
    .b(a_44_),
    .c(_0003_)
  );
  or_bb _0166_ (
    .a(_0003_),
    .b(a_42_),
    .c(_g_0_g_0_g_0_c_0_)
  );
  maj_bbb _0167_ (
    .a(a_42_),
    .b(a_43_),
    .c(a_44_),
    .d(_g_0_g_0_g_0_c_1_)
  );
  and_bb _0168_ (
    .a(a_43_),
    .b(a_44_),
    .c(_0002_)
  );
  and_bb _0169_ (
    .a(_0002_),
    .b(a_42_),
    .c(_g_0_g_0_g_0_c_2_)
  );
  or_bb _0170_ (
    .a(_g_0_g_0_g_0_c_2_),
    .b(_g_0_g_0_g_0_c_5_),
    .c(_g_0_g_0_g_0_g_3_c_5_)
  );
  and_bb _0171_ (
    .a(_g_0_g_0_g_0_c_2_),
    .b(_g_0_g_0_g_0_c_5_),
    .c(_g_0_g_0_g_0_g_3_c_2_)
  );
  or_bb _0172_ (
    .a(_g_0_g_0_g_0_c_1_),
    .b(_g_0_g_0_g_0_c_4_),
    .c(_g_0_g_0_g_0_g_3_c_4_)
  );
  and_bb _0173_ (
    .a(_g_0_g_0_g_0_c_1_),
    .b(_g_0_g_0_g_0_c_4_),
    .c(_g_0_g_0_g_0_g_3_c_1_)
  );
  or_bb _0174_ (
    .a(_g_0_g_0_g_0_c_0_),
    .b(_g_0_g_0_g_0_c_3_),
    .c(_g_0_g_0_g_0_g_3_c_3_)
  );
  and_bb _0175_ (
    .a(_g_0_g_0_g_0_c_0_),
    .b(_g_0_g_0_g_0_c_3_),
    .c(_g_0_g_0_g_0_g_3_c_0_)
  );
  or_bb _0176_ (
    .a(_g_0_g_0_g_0_g_3_c_4_),
    .b(_g_0_g_0_g_0_g_3_c_5_),
    .c(_0005_)
  );
  or_bb _0177_ (
    .a(_0005_),
    .b(_g_0_g_0_g_0_g_3_c_3_),
    .c(_g_0_g_0_c_11_)
  );
  maj_bbb _0178_ (
    .a(_g_0_g_0_g_0_g_3_c_3_),
    .b(_g_0_g_0_g_0_g_3_c_4_),
    .c(_g_0_g_0_g_0_g_3_c_5_),
    .d(_g_0_g_0_c_10_)
  );
  and_bb _0179_ (
    .a(_g_0_g_0_g_0_g_3_c_4_),
    .b(_g_0_g_0_g_0_g_3_c_5_),
    .c(_0004_)
  );
  and_bb _0180_ (
    .a(_0004_),
    .b(_g_0_g_0_g_0_g_3_c_3_),
    .c(_g_0_g_0_c_9_)
  );
  or_bb _0181_ (
    .a(_g_0_g_0_g_0_g_3_c_1_),
    .b(_g_0_g_0_g_0_g_3_c_2_),
    .c(_0007_)
  );
  or_bb _0182_ (
    .a(_0007_),
    .b(_g_0_g_0_g_0_g_3_c_0_),
    .c(_g_0_g_0_c_8_)
  );
  maj_bbb _0183_ (
    .a(_g_0_g_0_g_0_g_3_c_0_),
    .b(_g_0_g_0_g_0_g_3_c_1_),
    .c(_g_0_g_0_g_0_g_3_c_2_),
    .d(_g_0_g_0_c_7_)
  );
  and_bb _0184_ (
    .a(_g_0_g_0_g_0_g_3_c_1_),
    .b(_g_0_g_0_g_0_g_3_c_2_),
    .c(_0006_)
  );
  and_bb _0185_ (
    .a(_0006_),
    .b(_g_0_g_0_g_0_g_3_c_0_),
    .c(_g_0_g_0_c_6_)
  );
  or_bb _0186_ (
    .a(a_40_),
    .b(a_41_),
    .c(_0009_)
  );
  or_bb _0187_ (
    .a(_0009_),
    .b(a_39_),
    .c(_g_0_g_0_g_1_c_5_)
  );
  maj_bbb _0188_ (
    .a(a_39_),
    .b(a_40_),
    .c(a_41_),
    .d(_g_0_g_0_g_1_c_4_)
  );
  and_bb _0189_ (
    .a(a_40_),
    .b(a_41_),
    .c(_0008_)
  );
  and_bb _0190_ (
    .a(_0008_),
    .b(a_39_),
    .c(_g_0_g_0_g_1_c_3_)
  );
  or_bb _0191_ (
    .a(a_37_),
    .b(a_38_),
    .c(_0011_)
  );
  or_bb _0192_ (
    .a(_0011_),
    .b(a_36_),
    .c(_g_0_g_0_g_1_c_0_)
  );
  maj_bbb _0193_ (
    .a(a_36_),
    .b(a_37_),
    .c(a_38_),
    .d(_g_0_g_0_g_1_c_1_)
  );
  and_bb _0194_ (
    .a(a_37_),
    .b(a_38_),
    .c(_0010_)
  );
  and_bb _0195_ (
    .a(_0010_),
    .b(a_36_),
    .c(_g_0_g_0_g_1_c_2_)
  );
  or_bb _0196_ (
    .a(_g_0_g_0_g_1_c_2_),
    .b(_g_0_g_0_g_1_c_5_),
    .c(_g_0_g_0_g_1_g_3_c_5_)
  );
  and_bb _0197_ (
    .a(_g_0_g_0_g_1_c_2_),
    .b(_g_0_g_0_g_1_c_5_),
    .c(_g_0_g_0_g_1_g_3_c_2_)
  );
  or_bb _0198_ (
    .a(_g_0_g_0_g_1_c_1_),
    .b(_g_0_g_0_g_1_c_4_),
    .c(_g_0_g_0_g_1_g_3_c_4_)
  );
  and_bb _0199_ (
    .a(_g_0_g_0_g_1_c_1_),
    .b(_g_0_g_0_g_1_c_4_),
    .c(_g_0_g_0_g_1_g_3_c_1_)
  );
  or_bb _0200_ (
    .a(_g_0_g_0_g_1_c_0_),
    .b(_g_0_g_0_g_1_c_3_),
    .c(_g_0_g_0_g_1_g_3_c_3_)
  );
  and_bb _0201_ (
    .a(_g_0_g_0_g_1_c_0_),
    .b(_g_0_g_0_g_1_c_3_),
    .c(_g_0_g_0_g_1_g_3_c_0_)
  );
  or_bb _0202_ (
    .a(_g_0_g_0_g_1_g_3_c_4_),
    .b(_g_0_g_0_g_1_g_3_c_5_),
    .c(_0013_)
  );
  or_bb _0203_ (
    .a(_0013_),
    .b(_g_0_g_0_g_1_g_3_c_3_),
    .c(_g_0_g_0_c_0_)
  );
  maj_bbb _0204_ (
    .a(_g_0_g_0_g_1_g_3_c_3_),
    .b(_g_0_g_0_g_1_g_3_c_4_),
    .c(_g_0_g_0_g_1_g_3_c_5_),
    .d(_g_0_g_0_c_1_)
  );
  and_bb _0205_ (
    .a(_g_0_g_0_g_1_g_3_c_4_),
    .b(_g_0_g_0_g_1_g_3_c_5_),
    .c(_0012_)
  );
  and_bb _0206_ (
    .a(_0012_),
    .b(_g_0_g_0_g_1_g_3_c_3_),
    .c(_g_0_g_0_c_2_)
  );
  or_bb _0207_ (
    .a(_g_0_g_0_g_1_g_3_c_1_),
    .b(_g_0_g_0_g_1_g_3_c_2_),
    .c(_0015_)
  );
  or_bb _0208_ (
    .a(_0015_),
    .b(_g_0_g_0_g_1_g_3_c_0_),
    .c(_g_0_g_0_c_3_)
  );
  maj_bbb _0209_ (
    .a(_g_0_g_0_g_1_g_3_c_0_),
    .b(_g_0_g_0_g_1_g_3_c_1_),
    .c(_g_0_g_0_g_1_g_3_c_2_),
    .d(_g_0_g_0_c_4_)
  );
  and_bb _0210_ (
    .a(_g_0_g_0_g_1_g_3_c_1_),
    .b(_g_0_g_0_g_1_g_3_c_2_),
    .c(_0014_)
  );
  and_bb _0211_ (
    .a(_0014_),
    .b(_g_0_g_0_g_1_g_3_c_0_),
    .c(_g_0_g_0_c_5_)
  );
  or_bb _0212_ (
    .a(_g_0_g_0_c_0_),
    .b(_g_0_g_0_c_6_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0213_ (
    .a(_g_0_g_0_c_0_),
    .b(_g_0_g_0_c_6_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0214_ (
    .a(_g_0_g_0_c_1_),
    .b(_g_0_g_0_c_7_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0215_ (
    .a(_g_0_g_0_c_1_),
    .b(_g_0_g_0_c_7_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0216_ (
    .a(_g_0_g_0_c_2_),
    .b(_g_0_g_0_c_8_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0217_ (
    .a(_g_0_g_0_c_2_),
    .b(_g_0_g_0_c_8_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0218_ (
    .a(_g_0_g_0_c_3_),
    .b(_g_0_g_0_c_9_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0219_ (
    .a(_g_0_g_0_c_3_),
    .b(_g_0_g_0_c_9_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0220_ (
    .a(_g_0_g_0_c_4_),
    .b(_g_0_g_0_c_10_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0221_ (
    .a(_g_0_g_0_c_4_),
    .b(_g_0_g_0_c_10_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0222_ (
    .a(_g_0_g_0_c_5_),
    .b(_g_0_g_0_c_11_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0223_ (
    .a(_g_0_g_0_c_5_),
    .b(_g_0_g_0_c_11_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0224_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0225_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0226_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0227_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0228_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0229_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0230_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0017_)
  );
  or_bb _0231_ (
    .a(_0017_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_0_c_17_)
  );
  maj_bbb _0232_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(_g_0_c_16_)
  );
  and_bb _0233_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0016_)
  );
  and_bb _0234_ (
    .a(_0016_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_0_c_15_)
  );
  or_bb _0235_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0019_)
  );
  or_bb _0236_ (
    .a(_0019_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_0_c_14_)
  );
  maj_bbb _0237_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(_g_0_c_13_)
  );
  and_bb _0238_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0018_)
  );
  and_bb _0239_ (
    .a(_0018_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_0_c_12_)
  );
  or_bb _0240_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0241_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0242_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0243_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0244_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0245_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0246_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0021_)
  );
  or_bb _0247_ (
    .a(_0021_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_0_c_23_)
  );
  maj_bbb _0248_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(_g_0_c_22_)
  );
  and_bb _0249_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0020_)
  );
  and_bb _0250_ (
    .a(_0020_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_0_c_21_)
  );
  or_bb _0251_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0023_)
  );
  or_bb _0252_ (
    .a(_0023_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_0_c_20_)
  );
  maj_bbb _0253_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(_g_0_c_19_)
  );
  and_bb _0254_ (
    .a(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0022_)
  );
  and_bb _0255_ (
    .a(_0022_),
    .b(_g_0_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_0_c_18_)
  );
  or_bb _0256_ (
    .a(a_34_),
    .b(a_35_),
    .c(_0025_)
  );
  or_bb _0257_ (
    .a(_0025_),
    .b(a_33_),
    .c(_g_0_g_1_g_0_c_5_)
  );
  maj_bbb _0258_ (
    .a(a_33_),
    .b(a_34_),
    .c(a_35_),
    .d(_g_0_g_1_g_0_c_4_)
  );
  and_bb _0259_ (
    .a(a_34_),
    .b(a_35_),
    .c(_0024_)
  );
  and_bb _0260_ (
    .a(_0024_),
    .b(a_33_),
    .c(_g_0_g_1_g_0_c_3_)
  );
  or_bb _0261_ (
    .a(a_31_),
    .b(a_32_),
    .c(_0027_)
  );
  or_bb _0262_ (
    .a(_0027_),
    .b(a_30_),
    .c(_g_0_g_1_g_0_c_0_)
  );
  maj_bbb _0263_ (
    .a(a_30_),
    .b(a_31_),
    .c(a_32_),
    .d(_g_0_g_1_g_0_c_1_)
  );
  and_bb _0264_ (
    .a(a_31_),
    .b(a_32_),
    .c(_0026_)
  );
  and_bb _0265_ (
    .a(_0026_),
    .b(a_30_),
    .c(_g_0_g_1_g_0_c_2_)
  );
  or_bb _0266_ (
    .a(_g_0_g_1_g_0_c_2_),
    .b(_g_0_g_1_g_0_c_5_),
    .c(_g_0_g_1_g_0_g_3_c_5_)
  );
  and_bb _0267_ (
    .a(_g_0_g_1_g_0_c_2_),
    .b(_g_0_g_1_g_0_c_5_),
    .c(_g_0_g_1_g_0_g_3_c_2_)
  );
  or_bb _0268_ (
    .a(_g_0_g_1_g_0_c_1_),
    .b(_g_0_g_1_g_0_c_4_),
    .c(_g_0_g_1_g_0_g_3_c_4_)
  );
  and_bb _0269_ (
    .a(_g_0_g_1_g_0_c_1_),
    .b(_g_0_g_1_g_0_c_4_),
    .c(_g_0_g_1_g_0_g_3_c_1_)
  );
  or_bb _0270_ (
    .a(_g_0_g_1_g_0_c_0_),
    .b(_g_0_g_1_g_0_c_3_),
    .c(_g_0_g_1_g_0_g_3_c_3_)
  );
  and_bb _0271_ (
    .a(_g_0_g_1_g_0_c_0_),
    .b(_g_0_g_1_g_0_c_3_),
    .c(_g_0_g_1_g_0_g_3_c_0_)
  );
  or_bb _0272_ (
    .a(_g_0_g_1_g_0_g_3_c_4_),
    .b(_g_0_g_1_g_0_g_3_c_5_),
    .c(_0029_)
  );
  or_bb _0273_ (
    .a(_0029_),
    .b(_g_0_g_1_g_0_g_3_c_3_),
    .c(_g_0_g_1_c_11_)
  );
  maj_bbb _0274_ (
    .a(_g_0_g_1_g_0_g_3_c_3_),
    .b(_g_0_g_1_g_0_g_3_c_4_),
    .c(_g_0_g_1_g_0_g_3_c_5_),
    .d(_g_0_g_1_c_10_)
  );
  and_bb _0275_ (
    .a(_g_0_g_1_g_0_g_3_c_4_),
    .b(_g_0_g_1_g_0_g_3_c_5_),
    .c(_0028_)
  );
  and_bb _0276_ (
    .a(_0028_),
    .b(_g_0_g_1_g_0_g_3_c_3_),
    .c(_g_0_g_1_c_9_)
  );
  or_bb _0277_ (
    .a(_g_0_g_1_g_0_g_3_c_1_),
    .b(_g_0_g_1_g_0_g_3_c_2_),
    .c(_0031_)
  );
  or_bb _0278_ (
    .a(_0031_),
    .b(_g_0_g_1_g_0_g_3_c_0_),
    .c(_g_0_g_1_c_8_)
  );
  maj_bbb _0279_ (
    .a(_g_0_g_1_g_0_g_3_c_0_),
    .b(_g_0_g_1_g_0_g_3_c_1_),
    .c(_g_0_g_1_g_0_g_3_c_2_),
    .d(_g_0_g_1_c_7_)
  );
  and_bb _0280_ (
    .a(_g_0_g_1_g_0_g_3_c_1_),
    .b(_g_0_g_1_g_0_g_3_c_2_),
    .c(_0030_)
  );
  and_bb _0281_ (
    .a(_0030_),
    .b(_g_0_g_1_g_0_g_3_c_0_),
    .c(_g_0_g_1_c_6_)
  );
  or_bb _0282_ (
    .a(a_28_),
    .b(a_29_),
    .c(_0033_)
  );
  or_bb _0283_ (
    .a(_0033_),
    .b(a_27_),
    .c(_g_0_g_1_g_1_c_5_)
  );
  maj_bbb _0284_ (
    .a(a_27_),
    .b(a_28_),
    .c(a_29_),
    .d(_g_0_g_1_g_1_c_4_)
  );
  and_bb _0285_ (
    .a(a_28_),
    .b(a_29_),
    .c(_0032_)
  );
  and_bb _0286_ (
    .a(_0032_),
    .b(a_27_),
    .c(_g_0_g_1_g_1_c_3_)
  );
  or_bb _0287_ (
    .a(a_25_),
    .b(a_26_),
    .c(_0035_)
  );
  or_bb _0288_ (
    .a(_0035_),
    .b(a_24_),
    .c(_g_0_g_1_g_1_c_0_)
  );
  maj_bbb _0289_ (
    .a(a_24_),
    .b(a_25_),
    .c(a_26_),
    .d(_g_0_g_1_g_1_c_1_)
  );
  and_bb _0290_ (
    .a(a_25_),
    .b(a_26_),
    .c(_0034_)
  );
  and_bb _0291_ (
    .a(_0034_),
    .b(a_24_),
    .c(_g_0_g_1_g_1_c_2_)
  );
  or_bb _0292_ (
    .a(_g_0_g_1_g_1_c_2_),
    .b(_g_0_g_1_g_1_c_5_),
    .c(_g_0_g_1_g_1_g_3_c_5_)
  );
  and_bb _0293_ (
    .a(_g_0_g_1_g_1_c_2_),
    .b(_g_0_g_1_g_1_c_5_),
    .c(_g_0_g_1_g_1_g_3_c_2_)
  );
  or_bb _0294_ (
    .a(_g_0_g_1_g_1_c_1_),
    .b(_g_0_g_1_g_1_c_4_),
    .c(_g_0_g_1_g_1_g_3_c_4_)
  );
  and_bb _0295_ (
    .a(_g_0_g_1_g_1_c_1_),
    .b(_g_0_g_1_g_1_c_4_),
    .c(_g_0_g_1_g_1_g_3_c_1_)
  );
  or_bb _0296_ (
    .a(_g_0_g_1_g_1_c_0_),
    .b(_g_0_g_1_g_1_c_3_),
    .c(_g_0_g_1_g_1_g_3_c_3_)
  );
  and_bb _0297_ (
    .a(_g_0_g_1_g_1_c_0_),
    .b(_g_0_g_1_g_1_c_3_),
    .c(_g_0_g_1_g_1_g_3_c_0_)
  );
  or_bb _0298_ (
    .a(_g_0_g_1_g_1_g_3_c_4_),
    .b(_g_0_g_1_g_1_g_3_c_5_),
    .c(_0037_)
  );
  or_bb _0299_ (
    .a(_0037_),
    .b(_g_0_g_1_g_1_g_3_c_3_),
    .c(_g_0_g_1_c_0_)
  );
  maj_bbb _0300_ (
    .a(_g_0_g_1_g_1_g_3_c_3_),
    .b(_g_0_g_1_g_1_g_3_c_4_),
    .c(_g_0_g_1_g_1_g_3_c_5_),
    .d(_g_0_g_1_c_1_)
  );
  and_bb _0301_ (
    .a(_g_0_g_1_g_1_g_3_c_4_),
    .b(_g_0_g_1_g_1_g_3_c_5_),
    .c(_0036_)
  );
  and_bb _0302_ (
    .a(_0036_),
    .b(_g_0_g_1_g_1_g_3_c_3_),
    .c(_g_0_g_1_c_2_)
  );
  or_bb _0303_ (
    .a(_g_0_g_1_g_1_g_3_c_1_),
    .b(_g_0_g_1_g_1_g_3_c_2_),
    .c(_0039_)
  );
  or_bb _0304_ (
    .a(_0039_),
    .b(_g_0_g_1_g_1_g_3_c_0_),
    .c(_g_0_g_1_c_3_)
  );
  maj_bbb _0305_ (
    .a(_g_0_g_1_g_1_g_3_c_0_),
    .b(_g_0_g_1_g_1_g_3_c_1_),
    .c(_g_0_g_1_g_1_g_3_c_2_),
    .d(_g_0_g_1_c_4_)
  );
  and_bb _0306_ (
    .a(_g_0_g_1_g_1_g_3_c_1_),
    .b(_g_0_g_1_g_1_g_3_c_2_),
    .c(_0038_)
  );
  and_bb _0307_ (
    .a(_0038_),
    .b(_g_0_g_1_g_1_g_3_c_0_),
    .c(_g_0_g_1_c_5_)
  );
  or_bb _0308_ (
    .a(_g_0_g_1_c_0_),
    .b(_g_0_g_1_c_6_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0309_ (
    .a(_g_0_g_1_c_0_),
    .b(_g_0_g_1_c_6_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0310_ (
    .a(_g_0_g_1_c_1_),
    .b(_g_0_g_1_c_7_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0311_ (
    .a(_g_0_g_1_c_1_),
    .b(_g_0_g_1_c_7_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0312_ (
    .a(_g_0_g_1_c_2_),
    .b(_g_0_g_1_c_8_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0313_ (
    .a(_g_0_g_1_c_2_),
    .b(_g_0_g_1_c_8_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0314_ (
    .a(_g_0_g_1_c_3_),
    .b(_g_0_g_1_c_9_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0315_ (
    .a(_g_0_g_1_c_3_),
    .b(_g_0_g_1_c_9_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0316_ (
    .a(_g_0_g_1_c_4_),
    .b(_g_0_g_1_c_10_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0317_ (
    .a(_g_0_g_1_c_4_),
    .b(_g_0_g_1_c_10_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0318_ (
    .a(_g_0_g_1_c_5_),
    .b(_g_0_g_1_c_11_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0319_ (
    .a(_g_0_g_1_c_5_),
    .b(_g_0_g_1_c_11_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0320_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0321_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0322_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0323_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0324_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0325_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0326_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0041_)
  );
  or_bb _0327_ (
    .a(_0041_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_0_c_6_)
  );
  maj_bbb _0328_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(_g_0_c_7_)
  );
  and_bb _0329_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0040_)
  );
  and_bb _0330_ (
    .a(_0040_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_0_c_8_)
  );
  or_bb _0331_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0043_)
  );
  or_bb _0332_ (
    .a(_0043_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_0_c_9_)
  );
  maj_bbb _0333_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(_g_0_c_10_)
  );
  and_bb _0334_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0042_)
  );
  and_bb _0335_ (
    .a(_0042_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_0_c_11_)
  );
  or_bb _0336_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0337_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0338_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0339_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0340_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0341_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0342_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0045_)
  );
  or_bb _0343_ (
    .a(_0045_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_0_c_0_)
  );
  maj_bbb _0344_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(_g_0_c_1_)
  );
  and_bb _0345_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0044_)
  );
  and_bb _0346_ (
    .a(_0044_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_0_c_2_)
  );
  or_bb _0347_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0047_)
  );
  or_bb _0348_ (
    .a(_0047_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_0_c_3_)
  );
  maj_bbb _0349_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(_g_0_c_4_)
  );
  and_bb _0350_ (
    .a(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0046_)
  );
  and_bb _0351_ (
    .a(_0046_),
    .b(_g_0_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_0_c_5_)
  );
  or_bb _0352_ (
    .a(_g_0_c_1_),
    .b(_g_0_c_13_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_)
  );
  and_bb _0353_ (
    .a(_g_0_c_1_),
    .b(_g_0_c_13_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_)
  );
  or_bb _0354_ (
    .a(_g_0_c_2_),
    .b(_g_0_c_14_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_)
  );
  and_bb _0355_ (
    .a(_g_0_c_2_),
    .b(_g_0_c_14_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_)
  );
  or_bb _0356_ (
    .a(_g_0_c_3_),
    .b(_g_0_c_15_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_)
  );
  and_bb _0357_ (
    .a(_g_0_c_3_),
    .b(_g_0_c_15_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_)
  );
  or_bb _0358_ (
    .a(_g_0_c_4_),
    .b(_g_0_c_16_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_)
  );
  and_bb _0359_ (
    .a(_g_0_c_4_),
    .b(_g_0_c_16_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_)
  );
  or_bb _0360_ (
    .a(_g_0_c_5_),
    .b(_g_0_c_17_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_)
  );
  and_bb _0361_ (
    .a(_g_0_c_5_),
    .b(_g_0_c_17_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_)
  );
  or_bb _0362_ (
    .a(_g_0_c_6_),
    .b(_g_0_c_18_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_)
  );
  and_bb _0363_ (
    .a(_g_0_c_6_),
    .b(_g_0_c_18_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_)
  );
  or_bb _0364_ (
    .a(_g_0_c_7_),
    .b(_g_0_c_19_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_)
  );
  and_bb _0365_ (
    .a(_g_0_c_7_),
    .b(_g_0_c_19_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_)
  );
  or_bb _0366_ (
    .a(_g_0_c_8_),
    .b(_g_0_c_20_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_)
  );
  and_bb _0367_ (
    .a(_g_0_c_8_),
    .b(_g_0_c_20_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_)
  );
  or_bb _0368_ (
    .a(_g_0_c_9_),
    .b(_g_0_c_21_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_)
  );
  and_bb _0369_ (
    .a(_g_0_c_9_),
    .b(_g_0_c_21_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_)
  );
  or_bb _0370_ (
    .a(_g_0_c_10_),
    .b(_g_0_c_22_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_)
  );
  and_bb _0371_ (
    .a(_g_0_c_10_),
    .b(_g_0_c_22_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_)
  );
  or_bb _0372_ (
    .a(_g_0_c_11_),
    .b(_g_0_c_23_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_)
  );
  and_bb _0373_ (
    .a(_g_0_c_11_),
    .b(_g_0_c_23_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_)
  );
  or_bb _0374_ (
    .a(_g_0_c_0_),
    .b(_g_0_c_12_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_)
  );
  and_bb _0375_ (
    .a(_g_0_c_0_),
    .b(_g_0_c_12_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_)
  );
  or_bb _0376_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0377_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0378_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0379_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0380_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0381_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0382_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0383_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0384_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0385_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0386_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0387_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0388_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0389_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0390_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0391_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0392_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0393_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0394_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0049_)
  );
  or_bb _0395_ (
    .a(_0049_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_29_)
  );
  maj_bbb _0396_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(c_28_)
  );
  and_bb _0397_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0048_)
  );
  and_bb _0398_ (
    .a(_0048_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_27_)
  );
  or_bb _0399_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0051_)
  );
  or_bb _0400_ (
    .a(_0051_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_26_)
  );
  maj_bbb _0401_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(c_25_)
  );
  and_bb _0402_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0050_)
  );
  and_bb _0403_ (
    .a(_0050_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_24_)
  );
  or_bb _0404_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0405_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0406_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0407_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0408_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0409_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0410_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0053_)
  );
  or_bb _0411_ (
    .a(_0053_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_35_)
  );
  maj_bbb _0412_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(c_34_)
  );
  and_bb _0413_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0052_)
  );
  and_bb _0414_ (
    .a(_0052_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_33_)
  );
  or_bb _0415_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0055_)
  );
  or_bb _0416_ (
    .a(_0055_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_32_)
  );
  maj_bbb _0417_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(c_31_)
  );
  and_bb _0418_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0054_)
  );
  and_bb _0419_ (
    .a(_0054_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_30_)
  );
  or_bb _0420_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0421_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0422_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0423_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0424_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0425_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0426_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0427_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0428_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0429_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0430_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0431_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0432_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0433_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0434_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0435_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0436_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0437_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0438_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0057_)
  );
  or_bb _0439_ (
    .a(_0057_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_41_)
  );
  maj_bbb _0440_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(c_40_)
  );
  and_bb _0441_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0056_)
  );
  and_bb _0442_ (
    .a(_0056_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_39_)
  );
  or_bb _0443_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0059_)
  );
  or_bb _0444_ (
    .a(_0059_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_38_)
  );
  maj_bbb _0445_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(c_37_)
  );
  and_bb _0446_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0058_)
  );
  and_bb _0447_ (
    .a(_0058_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_36_)
  );
  or_bb _0448_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0449_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0450_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0451_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0452_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0453_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0454_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0061_)
  );
  or_bb _0455_ (
    .a(_0061_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_47_)
  );
  maj_bbb _0456_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(c_46_)
  );
  and_bb _0457_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0060_)
  );
  and_bb _0458_ (
    .a(_0060_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_45_)
  );
  or_bb _0459_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0063_)
  );
  or_bb _0460_ (
    .a(_0063_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_44_)
  );
  maj_bbb _0461_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(c_43_)
  );
  and_bb _0462_ (
    .a(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0062_)
  );
  and_bb _0463_ (
    .a(_0062_),
    .b(_g_0_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_42_)
  );
  or_bb _0464_ (
    .a(a_22_),
    .b(a_23_),
    .c(_0065_)
  );
  or_bb _0465_ (
    .a(_0065_),
    .b(a_21_),
    .c(_g_1_g_0_g_0_c_5_)
  );
  maj_bbb _0466_ (
    .a(a_21_),
    .b(a_22_),
    .c(a_23_),
    .d(_g_1_g_0_g_0_c_4_)
  );
  and_bb _0467_ (
    .a(a_22_),
    .b(a_23_),
    .c(_0064_)
  );
  and_bb _0468_ (
    .a(_0064_),
    .b(a_21_),
    .c(_g_1_g_0_g_0_c_3_)
  );
  or_bb _0469_ (
    .a(a_19_),
    .b(a_20_),
    .c(_0067_)
  );
  or_bb _0470_ (
    .a(_0067_),
    .b(a_18_),
    .c(_g_1_g_0_g_0_c_0_)
  );
  maj_bbb _0471_ (
    .a(a_18_),
    .b(a_19_),
    .c(a_20_),
    .d(_g_1_g_0_g_0_c_1_)
  );
  and_bb _0472_ (
    .a(a_19_),
    .b(a_20_),
    .c(_0066_)
  );
  and_bb _0473_ (
    .a(_0066_),
    .b(a_18_),
    .c(_g_1_g_0_g_0_c_2_)
  );
  or_bb _0474_ (
    .a(_g_1_g_0_g_0_c_2_),
    .b(_g_1_g_0_g_0_c_5_),
    .c(_g_1_g_0_g_0_g_3_c_5_)
  );
  and_bb _0475_ (
    .a(_g_1_g_0_g_0_c_2_),
    .b(_g_1_g_0_g_0_c_5_),
    .c(_g_1_g_0_g_0_g_3_c_2_)
  );
  or_bb _0476_ (
    .a(_g_1_g_0_g_0_c_1_),
    .b(_g_1_g_0_g_0_c_4_),
    .c(_g_1_g_0_g_0_g_3_c_4_)
  );
  and_bb _0477_ (
    .a(_g_1_g_0_g_0_c_1_),
    .b(_g_1_g_0_g_0_c_4_),
    .c(_g_1_g_0_g_0_g_3_c_1_)
  );
  or_bb _0478_ (
    .a(_g_1_g_0_g_0_c_0_),
    .b(_g_1_g_0_g_0_c_3_),
    .c(_g_1_g_0_g_0_g_3_c_3_)
  );
  and_bb _0479_ (
    .a(_g_1_g_0_g_0_c_0_),
    .b(_g_1_g_0_g_0_c_3_),
    .c(_g_1_g_0_g_0_g_3_c_0_)
  );
  or_bb _0480_ (
    .a(_g_1_g_0_g_0_g_3_c_4_),
    .b(_g_1_g_0_g_0_g_3_c_5_),
    .c(_0069_)
  );
  or_bb _0481_ (
    .a(_0069_),
    .b(_g_1_g_0_g_0_g_3_c_3_),
    .c(_g_1_g_0_c_11_)
  );
  maj_bbb _0482_ (
    .a(_g_1_g_0_g_0_g_3_c_3_),
    .b(_g_1_g_0_g_0_g_3_c_4_),
    .c(_g_1_g_0_g_0_g_3_c_5_),
    .d(_g_1_g_0_c_10_)
  );
  and_bb _0483_ (
    .a(_g_1_g_0_g_0_g_3_c_4_),
    .b(_g_1_g_0_g_0_g_3_c_5_),
    .c(_0068_)
  );
  and_bb _0484_ (
    .a(_0068_),
    .b(_g_1_g_0_g_0_g_3_c_3_),
    .c(_g_1_g_0_c_9_)
  );
  or_bb _0485_ (
    .a(_g_1_g_0_g_0_g_3_c_1_),
    .b(_g_1_g_0_g_0_g_3_c_2_),
    .c(_0071_)
  );
  or_bb _0486_ (
    .a(_0071_),
    .b(_g_1_g_0_g_0_g_3_c_0_),
    .c(_g_1_g_0_c_8_)
  );
  maj_bbb _0487_ (
    .a(_g_1_g_0_g_0_g_3_c_0_),
    .b(_g_1_g_0_g_0_g_3_c_1_),
    .c(_g_1_g_0_g_0_g_3_c_2_),
    .d(_g_1_g_0_c_7_)
  );
  and_bb _0488_ (
    .a(_g_1_g_0_g_0_g_3_c_1_),
    .b(_g_1_g_0_g_0_g_3_c_2_),
    .c(_0070_)
  );
  and_bb _0489_ (
    .a(_0070_),
    .b(_g_1_g_0_g_0_g_3_c_0_),
    .c(_g_1_g_0_c_6_)
  );
  or_bb _0490_ (
    .a(a_16_),
    .b(a_17_),
    .c(_0073_)
  );
  or_bb _0491_ (
    .a(_0073_),
    .b(a_15_),
    .c(_g_1_g_0_g_1_c_5_)
  );
  maj_bbb _0492_ (
    .a(a_15_),
    .b(a_16_),
    .c(a_17_),
    .d(_g_1_g_0_g_1_c_4_)
  );
  and_bb _0493_ (
    .a(a_16_),
    .b(a_17_),
    .c(_0072_)
  );
  and_bb _0494_ (
    .a(_0072_),
    .b(a_15_),
    .c(_g_1_g_0_g_1_c_3_)
  );
  or_bb _0495_ (
    .a(a_13_),
    .b(a_14_),
    .c(_0075_)
  );
  or_bb _0496_ (
    .a(_0075_),
    .b(a_12_),
    .c(_g_1_g_0_g_1_c_0_)
  );
  maj_bbb _0497_ (
    .a(a_12_),
    .b(a_13_),
    .c(a_14_),
    .d(_g_1_g_0_g_1_c_1_)
  );
  and_bb _0498_ (
    .a(a_13_),
    .b(a_14_),
    .c(_0074_)
  );
  and_bb _0499_ (
    .a(_0074_),
    .b(a_12_),
    .c(_g_1_g_0_g_1_c_2_)
  );
  or_bb _0500_ (
    .a(_g_1_g_0_g_1_c_2_),
    .b(_g_1_g_0_g_1_c_5_),
    .c(_g_1_g_0_g_1_g_3_c_5_)
  );
  and_bb _0501_ (
    .a(_g_1_g_0_g_1_c_2_),
    .b(_g_1_g_0_g_1_c_5_),
    .c(_g_1_g_0_g_1_g_3_c_2_)
  );
  or_bb _0502_ (
    .a(_g_1_g_0_g_1_c_1_),
    .b(_g_1_g_0_g_1_c_4_),
    .c(_g_1_g_0_g_1_g_3_c_4_)
  );
  and_bb _0503_ (
    .a(_g_1_g_0_g_1_c_1_),
    .b(_g_1_g_0_g_1_c_4_),
    .c(_g_1_g_0_g_1_g_3_c_1_)
  );
  or_bb _0504_ (
    .a(_g_1_g_0_g_1_c_0_),
    .b(_g_1_g_0_g_1_c_3_),
    .c(_g_1_g_0_g_1_g_3_c_3_)
  );
  and_bb _0505_ (
    .a(_g_1_g_0_g_1_c_0_),
    .b(_g_1_g_0_g_1_c_3_),
    .c(_g_1_g_0_g_1_g_3_c_0_)
  );
  or_bb _0506_ (
    .a(_g_1_g_0_g_1_g_3_c_4_),
    .b(_g_1_g_0_g_1_g_3_c_5_),
    .c(_0077_)
  );
  or_bb _0507_ (
    .a(_0077_),
    .b(_g_1_g_0_g_1_g_3_c_3_),
    .c(_g_1_g_0_c_0_)
  );
  maj_bbb _0508_ (
    .a(_g_1_g_0_g_1_g_3_c_3_),
    .b(_g_1_g_0_g_1_g_3_c_4_),
    .c(_g_1_g_0_g_1_g_3_c_5_),
    .d(_g_1_g_0_c_1_)
  );
  and_bb _0509_ (
    .a(_g_1_g_0_g_1_g_3_c_4_),
    .b(_g_1_g_0_g_1_g_3_c_5_),
    .c(_0076_)
  );
  and_bb _0510_ (
    .a(_0076_),
    .b(_g_1_g_0_g_1_g_3_c_3_),
    .c(_g_1_g_0_c_2_)
  );
  or_bb _0511_ (
    .a(_g_1_g_0_g_1_g_3_c_1_),
    .b(_g_1_g_0_g_1_g_3_c_2_),
    .c(_0079_)
  );
  or_bb _0512_ (
    .a(_0079_),
    .b(_g_1_g_0_g_1_g_3_c_0_),
    .c(_g_1_g_0_c_3_)
  );
  maj_bbb _0513_ (
    .a(_g_1_g_0_g_1_g_3_c_0_),
    .b(_g_1_g_0_g_1_g_3_c_1_),
    .c(_g_1_g_0_g_1_g_3_c_2_),
    .d(_g_1_g_0_c_4_)
  );
  and_bb _0514_ (
    .a(_g_1_g_0_g_1_g_3_c_1_),
    .b(_g_1_g_0_g_1_g_3_c_2_),
    .c(_0078_)
  );
  and_bb _0515_ (
    .a(_0078_),
    .b(_g_1_g_0_g_1_g_3_c_0_),
    .c(_g_1_g_0_c_5_)
  );
  or_bb _0516_ (
    .a(_g_1_g_0_c_0_),
    .b(_g_1_g_0_c_6_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0517_ (
    .a(_g_1_g_0_c_0_),
    .b(_g_1_g_0_c_6_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0518_ (
    .a(_g_1_g_0_c_1_),
    .b(_g_1_g_0_c_7_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0519_ (
    .a(_g_1_g_0_c_1_),
    .b(_g_1_g_0_c_7_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0520_ (
    .a(_g_1_g_0_c_2_),
    .b(_g_1_g_0_c_8_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0521_ (
    .a(_g_1_g_0_c_2_),
    .b(_g_1_g_0_c_8_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0522_ (
    .a(_g_1_g_0_c_3_),
    .b(_g_1_g_0_c_9_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0523_ (
    .a(_g_1_g_0_c_3_),
    .b(_g_1_g_0_c_9_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0524_ (
    .a(_g_1_g_0_c_4_),
    .b(_g_1_g_0_c_10_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0525_ (
    .a(_g_1_g_0_c_4_),
    .b(_g_1_g_0_c_10_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0526_ (
    .a(_g_1_g_0_c_5_),
    .b(_g_1_g_0_c_11_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0527_ (
    .a(_g_1_g_0_c_5_),
    .b(_g_1_g_0_c_11_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0528_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0529_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0530_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0531_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0532_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0533_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0534_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0081_)
  );
  or_bb _0535_ (
    .a(_0081_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_1_c_17_)
  );
  maj_bbb _0536_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(_g_1_c_16_)
  );
  and_bb _0537_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0080_)
  );
  and_bb _0538_ (
    .a(_0080_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_1_c_15_)
  );
  or_bb _0539_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0083_)
  );
  or_bb _0540_ (
    .a(_0083_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_1_c_14_)
  );
  maj_bbb _0541_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(_g_1_c_13_)
  );
  and_bb _0542_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0082_)
  );
  and_bb _0543_ (
    .a(_0082_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_1_c_12_)
  );
  or_bb _0544_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0545_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0546_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0547_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0548_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0549_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0550_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0085_)
  );
  or_bb _0551_ (
    .a(_0085_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_1_c_23_)
  );
  maj_bbb _0552_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(_g_1_c_22_)
  );
  and_bb _0553_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0084_)
  );
  and_bb _0554_ (
    .a(_0084_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_1_c_21_)
  );
  or_bb _0555_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0087_)
  );
  or_bb _0556_ (
    .a(_0087_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_1_c_20_)
  );
  maj_bbb _0557_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(_g_1_c_19_)
  );
  and_bb _0558_ (
    .a(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0086_)
  );
  and_bb _0559_ (
    .a(_0086_),
    .b(_g_1_g_0_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_1_c_18_)
  );
  or_bb _0560_ (
    .a(a_10_),
    .b(a_11_),
    .c(_0089_)
  );
  or_bb _0561_ (
    .a(_0089_),
    .b(a_9_),
    .c(_g_1_g_1_g_0_c_5_)
  );
  maj_bbb _0562_ (
    .a(a_9_),
    .b(a_10_),
    .c(a_11_),
    .d(_g_1_g_1_g_0_c_4_)
  );
  and_bb _0563_ (
    .a(a_10_),
    .b(a_11_),
    .c(_0088_)
  );
  and_bb _0564_ (
    .a(_0088_),
    .b(a_9_),
    .c(_g_1_g_1_g_0_c_3_)
  );
  or_bb _0565_ (
    .a(a_7_),
    .b(a_8_),
    .c(_0091_)
  );
  or_bb _0566_ (
    .a(_0091_),
    .b(a_6_),
    .c(_g_1_g_1_g_0_c_0_)
  );
  maj_bbb _0567_ (
    .a(a_6_),
    .b(a_7_),
    .c(a_8_),
    .d(_g_1_g_1_g_0_c_1_)
  );
  and_bb _0568_ (
    .a(a_7_),
    .b(a_8_),
    .c(_0090_)
  );
  and_bb _0569_ (
    .a(_0090_),
    .b(a_6_),
    .c(_g_1_g_1_g_0_c_2_)
  );
  or_bb _0570_ (
    .a(_g_1_g_1_g_0_c_2_),
    .b(_g_1_g_1_g_0_c_5_),
    .c(_g_1_g_1_g_0_g_3_c_5_)
  );
  and_bb _0571_ (
    .a(_g_1_g_1_g_0_c_2_),
    .b(_g_1_g_1_g_0_c_5_),
    .c(_g_1_g_1_g_0_g_3_c_2_)
  );
  or_bb _0572_ (
    .a(_g_1_g_1_g_0_c_1_),
    .b(_g_1_g_1_g_0_c_4_),
    .c(_g_1_g_1_g_0_g_3_c_4_)
  );
  and_bb _0573_ (
    .a(_g_1_g_1_g_0_c_1_),
    .b(_g_1_g_1_g_0_c_4_),
    .c(_g_1_g_1_g_0_g_3_c_1_)
  );
  or_bb _0574_ (
    .a(_g_1_g_1_g_0_c_0_),
    .b(_g_1_g_1_g_0_c_3_),
    .c(_g_1_g_1_g_0_g_3_c_3_)
  );
  and_bb _0575_ (
    .a(_g_1_g_1_g_0_c_0_),
    .b(_g_1_g_1_g_0_c_3_),
    .c(_g_1_g_1_g_0_g_3_c_0_)
  );
  or_bb _0576_ (
    .a(_g_1_g_1_g_0_g_3_c_4_),
    .b(_g_1_g_1_g_0_g_3_c_5_),
    .c(_0093_)
  );
  or_bb _0577_ (
    .a(_0093_),
    .b(_g_1_g_1_g_0_g_3_c_3_),
    .c(_g_1_g_1_c_11_)
  );
  maj_bbb _0578_ (
    .a(_g_1_g_1_g_0_g_3_c_3_),
    .b(_g_1_g_1_g_0_g_3_c_4_),
    .c(_g_1_g_1_g_0_g_3_c_5_),
    .d(_g_1_g_1_c_10_)
  );
  and_bb _0579_ (
    .a(_g_1_g_1_g_0_g_3_c_4_),
    .b(_g_1_g_1_g_0_g_3_c_5_),
    .c(_0092_)
  );
  and_bb _0580_ (
    .a(_0092_),
    .b(_g_1_g_1_g_0_g_3_c_3_),
    .c(_g_1_g_1_c_9_)
  );
  or_bb _0581_ (
    .a(_g_1_g_1_g_0_g_3_c_1_),
    .b(_g_1_g_1_g_0_g_3_c_2_),
    .c(_0095_)
  );
  or_bb _0582_ (
    .a(_0095_),
    .b(_g_1_g_1_g_0_g_3_c_0_),
    .c(_g_1_g_1_c_8_)
  );
  maj_bbb _0583_ (
    .a(_g_1_g_1_g_0_g_3_c_0_),
    .b(_g_1_g_1_g_0_g_3_c_1_),
    .c(_g_1_g_1_g_0_g_3_c_2_),
    .d(_g_1_g_1_c_7_)
  );
  and_bb _0584_ (
    .a(_g_1_g_1_g_0_g_3_c_1_),
    .b(_g_1_g_1_g_0_g_3_c_2_),
    .c(_0094_)
  );
  and_bb _0585_ (
    .a(_0094_),
    .b(_g_1_g_1_g_0_g_3_c_0_),
    .c(_g_1_g_1_c_6_)
  );
  or_bb _0586_ (
    .a(a_4_),
    .b(a_5_),
    .c(_0097_)
  );
  or_bb _0587_ (
    .a(_0097_),
    .b(a_3_),
    .c(_g_1_g_1_g_1_c_5_)
  );
  maj_bbb _0588_ (
    .a(a_3_),
    .b(a_4_),
    .c(a_5_),
    .d(_g_1_g_1_g_1_c_4_)
  );
  and_bb _0589_ (
    .a(a_4_),
    .b(a_5_),
    .c(_0096_)
  );
  and_bb _0590_ (
    .a(_0096_),
    .b(a_3_),
    .c(_g_1_g_1_g_1_c_3_)
  );
  or_bb _0591_ (
    .a(a_1_),
    .b(a_2_),
    .c(_0099_)
  );
  or_bb _0592_ (
    .a(_0099_),
    .b(a_0_),
    .c(_g_1_g_1_g_1_c_0_)
  );
  maj_bbb _0593_ (
    .a(a_0_),
    .b(a_1_),
    .c(a_2_),
    .d(_g_1_g_1_g_1_c_1_)
  );
  and_bb _0594_ (
    .a(a_1_),
    .b(a_2_),
    .c(_0098_)
  );
  and_bb _0595_ (
    .a(_0098_),
    .b(a_0_),
    .c(_g_1_g_1_g_1_c_2_)
  );
  or_bb _0596_ (
    .a(_g_1_g_1_g_1_c_2_),
    .b(_g_1_g_1_g_1_c_5_),
    .c(_g_1_g_1_g_1_g_3_c_5_)
  );
  and_bb _0597_ (
    .a(_g_1_g_1_g_1_c_2_),
    .b(_g_1_g_1_g_1_c_5_),
    .c(_g_1_g_1_g_1_g_3_c_2_)
  );
  or_bb _0598_ (
    .a(_g_1_g_1_g_1_c_1_),
    .b(_g_1_g_1_g_1_c_4_),
    .c(_g_1_g_1_g_1_g_3_c_4_)
  );
  and_bb _0599_ (
    .a(_g_1_g_1_g_1_c_1_),
    .b(_g_1_g_1_g_1_c_4_),
    .c(_g_1_g_1_g_1_g_3_c_1_)
  );
  or_bb _0600_ (
    .a(_g_1_g_1_g_1_c_0_),
    .b(_g_1_g_1_g_1_c_3_),
    .c(_g_1_g_1_g_1_g_3_c_3_)
  );
  and_bb _0601_ (
    .a(_g_1_g_1_g_1_c_0_),
    .b(_g_1_g_1_g_1_c_3_),
    .c(_g_1_g_1_g_1_g_3_c_0_)
  );
  or_bb _0602_ (
    .a(_g_1_g_1_g_1_g_3_c_4_),
    .b(_g_1_g_1_g_1_g_3_c_5_),
    .c(_0101_)
  );
  or_bb _0603_ (
    .a(_0101_),
    .b(_g_1_g_1_g_1_g_3_c_3_),
    .c(_g_1_g_1_c_0_)
  );
  maj_bbb _0604_ (
    .a(_g_1_g_1_g_1_g_3_c_3_),
    .b(_g_1_g_1_g_1_g_3_c_4_),
    .c(_g_1_g_1_g_1_g_3_c_5_),
    .d(_g_1_g_1_c_1_)
  );
  and_bb _0605_ (
    .a(_g_1_g_1_g_1_g_3_c_4_),
    .b(_g_1_g_1_g_1_g_3_c_5_),
    .c(_0100_)
  );
  and_bb _0606_ (
    .a(_0100_),
    .b(_g_1_g_1_g_1_g_3_c_3_),
    .c(_g_1_g_1_c_2_)
  );
  or_bb _0607_ (
    .a(_g_1_g_1_g_1_g_3_c_1_),
    .b(_g_1_g_1_g_1_g_3_c_2_),
    .c(_0103_)
  );
  or_bb _0608_ (
    .a(_0103_),
    .b(_g_1_g_1_g_1_g_3_c_0_),
    .c(_g_1_g_1_c_3_)
  );
  maj_bbb _0609_ (
    .a(_g_1_g_1_g_1_g_3_c_0_),
    .b(_g_1_g_1_g_1_g_3_c_1_),
    .c(_g_1_g_1_g_1_g_3_c_2_),
    .d(_g_1_g_1_c_4_)
  );
  and_bb _0610_ (
    .a(_g_1_g_1_g_1_g_3_c_1_),
    .b(_g_1_g_1_g_1_g_3_c_2_),
    .c(_0102_)
  );
  and_bb _0611_ (
    .a(_0102_),
    .b(_g_1_g_1_g_1_g_3_c_0_),
    .c(_g_1_g_1_c_5_)
  );
  or_bb _0612_ (
    .a(_g_1_g_1_c_0_),
    .b(_g_1_g_1_c_6_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0613_ (
    .a(_g_1_g_1_c_0_),
    .b(_g_1_g_1_c_6_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0614_ (
    .a(_g_1_g_1_c_1_),
    .b(_g_1_g_1_c_7_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0615_ (
    .a(_g_1_g_1_c_1_),
    .b(_g_1_g_1_c_7_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0616_ (
    .a(_g_1_g_1_c_2_),
    .b(_g_1_g_1_c_8_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0617_ (
    .a(_g_1_g_1_c_2_),
    .b(_g_1_g_1_c_8_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0618_ (
    .a(_g_1_g_1_c_3_),
    .b(_g_1_g_1_c_9_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0619_ (
    .a(_g_1_g_1_c_3_),
    .b(_g_1_g_1_c_9_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0620_ (
    .a(_g_1_g_1_c_4_),
    .b(_g_1_g_1_c_10_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0621_ (
    .a(_g_1_g_1_c_4_),
    .b(_g_1_g_1_c_10_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0622_ (
    .a(_g_1_g_1_c_5_),
    .b(_g_1_g_1_c_11_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0623_ (
    .a(_g_1_g_1_c_5_),
    .b(_g_1_g_1_c_11_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0624_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0625_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0626_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0627_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0628_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0629_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0630_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0105_)
  );
  or_bb _0631_ (
    .a(_0105_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_1_c_6_)
  );
  maj_bbb _0632_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(_g_1_c_7_)
  );
  and_bb _0633_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0104_)
  );
  and_bb _0634_ (
    .a(_0104_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(_g_1_c_8_)
  );
  or_bb _0635_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0107_)
  );
  or_bb _0636_ (
    .a(_0107_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_1_c_9_)
  );
  maj_bbb _0637_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(_g_1_c_10_)
  );
  and_bb _0638_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0106_)
  );
  and_bb _0639_ (
    .a(_0106_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(_g_1_c_11_)
  );
  or_bb _0640_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0641_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0642_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0643_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0644_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0645_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0646_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0109_)
  );
  or_bb _0647_ (
    .a(_0109_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_1_c_0_)
  );
  maj_bbb _0648_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(_g_1_c_1_)
  );
  and_bb _0649_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0108_)
  );
  and_bb _0650_ (
    .a(_0108_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(_g_1_c_2_)
  );
  or_bb _0651_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0111_)
  );
  or_bb _0652_ (
    .a(_0111_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_1_c_3_)
  );
  maj_bbb _0653_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(_g_1_c_4_)
  );
  and_bb _0654_ (
    .a(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0110_)
  );
  and_bb _0655_ (
    .a(_0110_),
    .b(_g_1_g_1_m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(_g_1_c_5_)
  );
  or_bb _0656_ (
    .a(_g_1_c_1_),
    .b(_g_1_c_13_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_)
  );
  and_bb _0657_ (
    .a(_g_1_c_1_),
    .b(_g_1_c_13_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_)
  );
  or_bb _0658_ (
    .a(_g_1_c_2_),
    .b(_g_1_c_14_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_)
  );
  and_bb _0659_ (
    .a(_g_1_c_2_),
    .b(_g_1_c_14_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_)
  );
  or_bb _0660_ (
    .a(_g_1_c_3_),
    .b(_g_1_c_15_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_)
  );
  and_bb _0661_ (
    .a(_g_1_c_3_),
    .b(_g_1_c_15_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_)
  );
  or_bb _0662_ (
    .a(_g_1_c_4_),
    .b(_g_1_c_16_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_)
  );
  and_bb _0663_ (
    .a(_g_1_c_4_),
    .b(_g_1_c_16_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_)
  );
  or_bb _0664_ (
    .a(_g_1_c_5_),
    .b(_g_1_c_17_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_)
  );
  and_bb _0665_ (
    .a(_g_1_c_5_),
    .b(_g_1_c_17_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_)
  );
  or_bb _0666_ (
    .a(_g_1_c_6_),
    .b(_g_1_c_18_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_)
  );
  and_bb _0667_ (
    .a(_g_1_c_6_),
    .b(_g_1_c_18_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_)
  );
  or_bb _0668_ (
    .a(_g_1_c_7_),
    .b(_g_1_c_19_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_)
  );
  and_bb _0669_ (
    .a(_g_1_c_7_),
    .b(_g_1_c_19_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_)
  );
  or_bb _0670_ (
    .a(_g_1_c_8_),
    .b(_g_1_c_20_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_)
  );
  and_bb _0671_ (
    .a(_g_1_c_8_),
    .b(_g_1_c_20_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_)
  );
  or_bb _0672_ (
    .a(_g_1_c_9_),
    .b(_g_1_c_21_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_)
  );
  and_bb _0673_ (
    .a(_g_1_c_9_),
    .b(_g_1_c_21_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_)
  );
  or_bb _0674_ (
    .a(_g_1_c_10_),
    .b(_g_1_c_22_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_)
  );
  and_bb _0675_ (
    .a(_g_1_c_10_),
    .b(_g_1_c_22_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_)
  );
  or_bb _0676_ (
    .a(_g_1_c_11_),
    .b(_g_1_c_23_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_)
  );
  and_bb _0677_ (
    .a(_g_1_c_11_),
    .b(_g_1_c_23_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_)
  );
  or_bb _0678_ (
    .a(_g_1_c_0_),
    .b(_g_1_c_12_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_)
  );
  and_bb _0679_ (
    .a(_g_1_c_0_),
    .b(_g_1_c_12_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_)
  );
  or_bb _0680_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0681_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0682_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0683_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0684_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0685_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0686_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0687_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0688_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0689_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0690_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0691_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0692_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0693_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0694_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0695_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0696_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0697_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0698_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0113_)
  );
  or_bb _0699_ (
    .a(_0113_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_18_)
  );
  maj_bbb _0700_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(c_19_)
  );
  and_bb _0701_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0112_)
  );
  and_bb _0702_ (
    .a(_0112_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_20_)
  );
  or_bb _0703_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0115_)
  );
  or_bb _0704_ (
    .a(_0115_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_21_)
  );
  maj_bbb _0705_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(c_22_)
  );
  and_bb _0706_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0114_)
  );
  and_bb _0707_ (
    .a(_0114_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_23_)
  );
  or_bb _0708_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0709_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0710_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0711_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0712_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0713_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0714_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0117_)
  );
  or_bb _0715_ (
    .a(_0117_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_12_)
  );
  maj_bbb _0716_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(c_13_)
  );
  and_bb _0717_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0116_)
  );
  and_bb _0718_ (
    .a(_0116_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_14_)
  );
  or_bb _0719_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0119_)
  );
  or_bb _0720_ (
    .a(_0119_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_15_)
  );
  maj_bbb _0721_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(c_16_)
  );
  and_bb _0722_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0118_)
  );
  and_bb _0723_ (
    .a(_0118_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_17_)
  );
  or_bb _0724_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0725_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0726_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0727_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0728_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0729_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0730_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0731_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0732_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0733_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0734_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0735_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0736_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0737_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0738_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0739_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0740_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0741_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0742_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0121_)
  );
  or_bb _0743_ (
    .a(_0121_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_6_)
  );
  maj_bbb _0744_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(c_7_)
  );
  and_bb _0745_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0120_)
  );
  and_bb _0746_ (
    .a(_0120_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(c_8_)
  );
  or_bb _0747_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0123_)
  );
  or_bb _0748_ (
    .a(_0123_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_9_)
  );
  maj_bbb _0749_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(c_10_)
  );
  and_bb _0750_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0122_)
  );
  and_bb _0751_ (
    .a(_0122_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(c_11_)
  );
  or_bb _0752_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0753_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0754_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0755_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0756_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0757_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0758_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0125_)
  );
  or_bb _0759_ (
    .a(_0125_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_0_)
  );
  maj_bbb _0760_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(c_1_)
  );
  and_bb _0761_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0124_)
  );
  and_bb _0762_ (
    .a(_0124_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(c_2_)
  );
  or_bb _0763_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0127_)
  );
  or_bb _0764_ (
    .a(_0127_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_3_)
  );
  maj_bbb _0765_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(c_4_)
  );
  and_bb _0766_ (
    .a(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0126_)
  );
  and_bb _0767_ (
    .a(_0126_),
    .b(_g_1_m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(c_5_)
  );
  or_bb _0768_ (
    .a(c_0_),
    .b(c_24_),
    .c(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_1_)
  );
  and_bb _0769_ (
    .a(c_0_),
    .b(c_24_),
    .c(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_0_)
  );
  or_bb _0770_ (
    .a(c_1_),
    .b(c_25_),
    .c(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_1_)
  );
  and_bb _0771_ (
    .a(c_1_),
    .b(c_25_),
    .c(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_0_)
  );
  or_bb _0772_ (
    .a(c_2_),
    .b(c_26_),
    .c(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_1_)
  );
  and_bb _0773_ (
    .a(c_2_),
    .b(c_26_),
    .c(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_0_)
  );
  or_bb _0774_ (
    .a(c_3_),
    .b(c_27_),
    .c(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_1_)
  );
  and_bb _0775_ (
    .a(c_3_),
    .b(c_27_),
    .c(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_0_)
  );
  or_bb _0776_ (
    .a(c_4_),
    .b(c_28_),
    .c(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_1_)
  );
  and_bb _0777_ (
    .a(c_4_),
    .b(c_28_),
    .c(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_0_)
  );
  or_bb _0778_ (
    .a(c_5_),
    .b(c_29_),
    .c(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_1_)
  );
  and_bb _0779_ (
    .a(c_5_),
    .b(c_29_),
    .c(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_0_)
  );
  or_bb _0780_ (
    .a(c_6_),
    .b(c_30_),
    .c(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_1_)
  );
  and_bb _0781_ (
    .a(c_6_),
    .b(c_30_),
    .c(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_0_)
  );
  or_bb _0782_ (
    .a(c_7_),
    .b(c_31_),
    .c(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_1_)
  );
  and_bb _0783_ (
    .a(c_7_),
    .b(c_31_),
    .c(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_0_)
  );
  or_bb _0784_ (
    .a(c_8_),
    .b(c_32_),
    .c(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_1_)
  );
  and_bb _0785_ (
    .a(c_8_),
    .b(c_32_),
    .c(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_0_)
  );
  or_bb _0786_ (
    .a(c_9_),
    .b(c_33_),
    .c(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_1_)
  );
  and_bb _0787_ (
    .a(c_9_),
    .b(c_33_),
    .c(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_0_)
  );
  or_bb _0788_ (
    .a(c_10_),
    .b(c_34_),
    .c(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_1_)
  );
  and_bb _0789_ (
    .a(c_10_),
    .b(c_34_),
    .c(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_0_)
  );
  or_bb _0790_ (
    .a(c_11_),
    .b(c_35_),
    .c(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_1_)
  );
  and_bb _0791_ (
    .a(c_11_),
    .b(c_35_),
    .c(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_0_)
  );
  or_bb _0792_ (
    .a(c_12_),
    .b(c_36_),
    .c(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_1_)
  );
  and_bb _0793_ (
    .a(c_12_),
    .b(c_36_),
    .c(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_0_)
  );
  or_bb _0794_ (
    .a(c_13_),
    .b(c_37_),
    .c(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_1_)
  );
  and_bb _0795_ (
    .a(c_13_),
    .b(c_37_),
    .c(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_0_)
  );
  or_bb _0796_ (
    .a(c_14_),
    .b(c_38_),
    .c(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_1_)
  );
  and_bb _0797_ (
    .a(c_14_),
    .b(c_38_),
    .c(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_0_)
  );
  or_bb _0798_ (
    .a(c_15_),
    .b(c_39_),
    .c(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_1_)
  );
  and_bb _0799_ (
    .a(c_15_),
    .b(c_39_),
    .c(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_0_)
  );
  or_bb _0800_ (
    .a(c_16_),
    .b(c_40_),
    .c(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_1_)
  );
  and_bb _0801_ (
    .a(c_16_),
    .b(c_40_),
    .c(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_0_)
  );
  or_bb _0802_ (
    .a(c_17_),
    .b(c_41_),
    .c(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_1_)
  );
  and_bb _0803_ (
    .a(c_17_),
    .b(c_41_),
    .c(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_0_)
  );
  or_bb _0804_ (
    .a(c_18_),
    .b(c_42_),
    .c(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_1_)
  );
  and_bb _0805_ (
    .a(c_18_),
    .b(c_42_),
    .c(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_0_)
  );
  or_bb _0806_ (
    .a(c_19_),
    .b(c_43_),
    .c(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_1_)
  );
  and_bb _0807_ (
    .a(c_19_),
    .b(c_43_),
    .c(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_0_)
  );
  or_bb _0808_ (
    .a(c_20_),
    .b(c_44_),
    .c(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_1_)
  );
  and_bb _0809_ (
    .a(c_20_),
    .b(c_44_),
    .c(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_0_)
  );
  or_bb _0810_ (
    .a(c_21_),
    .b(c_45_),
    .c(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_1_)
  );
  and_bb _0811_ (
    .a(c_21_),
    .b(c_45_),
    .c(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_0_)
  );
  or_bb _0812_ (
    .a(c_22_),
    .b(c_46_),
    .c(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_1_)
  );
  and_bb _0813_ (
    .a(c_22_),
    .b(c_46_),
    .c(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_0_)
  );
  or_bb _0814_ (
    .a(c_23_),
    .b(c_47_),
    .c(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_1_)
  );
  and_bb _0815_ (
    .a(c_23_),
    .b(c_47_),
    .c(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_0_)
  );
  or_bb _0816_ (
    .a(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_)
  );
  and_bb _0817_ (
    .a(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_)
  );
  or_bb _0818_ (
    .a(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_)
  );
  and_bb _0819_ (
    .a(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_)
  );
  or_bb _0820_ (
    .a(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_)
  );
  and_bb _0821_ (
    .a(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_)
  );
  or_bb _0822_ (
    .a(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_)
  );
  and_bb _0823_ (
    .a(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_)
  );
  or_bb _0824_ (
    .a(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_)
  );
  and_bb _0825_ (
    .a(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_)
  );
  or_bb _0826_ (
    .a(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_)
  );
  and_bb _0827_ (
    .a(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_)
  );
  or_bb _0828_ (
    .a(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_)
  );
  and_bb _0829_ (
    .a(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_)
  );
  or_bb _0830_ (
    .a(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_)
  );
  and_bb _0831_ (
    .a(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_)
  );
  or_bb _0832_ (
    .a(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_)
  );
  and_bb _0833_ (
    .a(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_)
  );
  or_bb _0834_ (
    .a(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_)
  );
  and_bb _0835_ (
    .a(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_)
  );
  or_bb _0836_ (
    .a(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_)
  );
  and_bb _0837_ (
    .a(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_)
  );
  or_bb _0838_ (
    .a(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_)
  );
  and_bb _0839_ (
    .a(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_)
  );
  or_bb _0840_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0841_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0842_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0843_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0844_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0845_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0846_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0847_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0848_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0849_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0850_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0851_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0852_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0853_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0854_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0855_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0856_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0857_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0858_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0129_)
  );
  or_bb _0859_ (
    .a(_0129_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_5_)
  );
  maj_bbb _0860_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(b_4_)
  );
  and_bb _0861_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0128_)
  );
  and_bb _0862_ (
    .a(_0128_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_3_)
  );
  or_bb _0863_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0131_)
  );
  or_bb _0864_ (
    .a(_0131_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_2_)
  );
  maj_bbb _0865_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(b_1_)
  );
  and_bb _0866_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0130_)
  );
  and_bb _0867_ (
    .a(_0130_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_0_)
  );
  or_bb _0868_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0869_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0870_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0871_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0872_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0873_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0874_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0133_)
  );
  or_bb _0875_ (
    .a(_0133_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_11_)
  );
  maj_bbb _0876_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(b_10_)
  );
  and_bb _0877_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0132_)
  );
  and_bb _0878_ (
    .a(_0132_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_9_)
  );
  or_bb _0879_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0135_)
  );
  or_bb _0880_ (
    .a(_0135_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_8_)
  );
  maj_bbb _0881_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(b_7_)
  );
  and_bb _0882_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0134_)
  );
  and_bb _0883_ (
    .a(_0134_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_6_)
  );
  or_bb _0884_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0885_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0886_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0887_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0888_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0889_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0890_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0891_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0892_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0893_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0894_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0895_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0896_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0897_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0898_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0899_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0900_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0901_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0902_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0137_)
  );
  or_bb _0903_ (
    .a(_0137_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_17_)
  );
  maj_bbb _0904_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(b_16_)
  );
  and_bb _0905_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0136_)
  );
  and_bb _0906_ (
    .a(_0136_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_15_)
  );
  or_bb _0907_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0139_)
  );
  or_bb _0908_ (
    .a(_0139_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_14_)
  );
  maj_bbb _0909_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(b_13_)
  );
  and_bb _0910_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0138_)
  );
  and_bb _0911_ (
    .a(_0138_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_12_)
  );
  or_bb _0912_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0913_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0914_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0915_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0916_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0917_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0918_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0141_)
  );
  or_bb _0919_ (
    .a(_0141_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_23_)
  );
  maj_bbb _0920_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(b_22_)
  );
  and_bb _0921_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0140_)
  );
  and_bb _0922_ (
    .a(_0140_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_21_)
  );
  or_bb _0923_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0143_)
  );
  or_bb _0924_ (
    .a(_0143_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_20_)
  );
  maj_bbb _0925_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(b_19_)
  );
  and_bb _0926_ (
    .a(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0142_)
  );
  and_bb _0927_ (
    .a(_0142_),
    .b(_m__genblock___src_b48s_merger48_v_13_47_0__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_18_)
  );
  or_bb _0928_ (
    .a(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_)
  );
  and_bb _0929_ (
    .a(_m__genblock___src_b48s_merger48_v_10_24_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_36_13__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_)
  );
  or_bb _0930_ (
    .a(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_)
  );
  and_bb _0931_ (
    .a(_m__genblock___src_b48s_merger48_v_10_25_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_37_14__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_)
  );
  or_bb _0932_ (
    .a(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_)
  );
  and_bb _0933_ (
    .a(_m__genblock___src_b48s_merger48_v_10_26_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_38_15__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_)
  );
  or_bb _0934_ (
    .a(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_)
  );
  and_bb _0935_ (
    .a(_m__genblock___src_b48s_merger48_v_10_27_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_39_16__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_)
  );
  or_bb _0936_ (
    .a(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_)
  );
  and_bb _0937_ (
    .a(_m__genblock___src_b48s_merger48_v_10_28_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_40_17__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_)
  );
  or_bb _0938_ (
    .a(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_)
  );
  and_bb _0939_ (
    .a(_m__genblock___src_b48s_merger48_v_10_29_6__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_41_18__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_)
  );
  or_bb _0940_ (
    .a(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_)
  );
  and_bb _0941_ (
    .a(_m__genblock___src_b48s_merger48_v_10_30_7__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_42_19__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_)
  );
  or_bb _0942_ (
    .a(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_)
  );
  and_bb _0943_ (
    .a(_m__genblock___src_b48s_merger48_v_10_31_8__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_43_20__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_)
  );
  or_bb _0944_ (
    .a(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_)
  );
  and_bb _0945_ (
    .a(_m__genblock___src_b48s_merger48_v_10_32_9__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_44_21__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_)
  );
  or_bb _0946_ (
    .a(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_)
  );
  and_bb _0947_ (
    .a(_m__genblock___src_b48s_merger48_v_10_33_10__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_45_22__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_)
  );
  or_bb _0948_ (
    .a(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_)
  );
  and_bb _0949_ (
    .a(_m__genblock___src_b48s_merger48_v_10_34_11__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_46_23__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_)
  );
  or_bb _0950_ (
    .a(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_)
  );
  and_bb _0951_ (
    .a(_m__genblock___src_b48s_merger48_v_10_23_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_10_35_12__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_)
  );
  or_bb _0952_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0953_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0954_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0955_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _0956_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _0957_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _0958_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _0959_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _0960_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _0961_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _0962_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _0963_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _0964_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _0965_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _0966_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _0967_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _0968_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _0969_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _0970_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0145_)
  );
  or_bb _0971_ (
    .a(_0145_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_29_)
  );
  maj_bbb _0972_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(b_28_)
  );
  and_bb _0973_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0144_)
  );
  and_bb _0974_ (
    .a(_0144_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_27_)
  );
  or_bb _0975_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0147_)
  );
  or_bb _0976_ (
    .a(_0147_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_26_)
  );
  maj_bbb _0977_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(b_25_)
  );
  and_bb _0978_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0146_)
  );
  and_bb _0979_ (
    .a(_0146_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_24_)
  );
  or_bb _0980_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _0981_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _0982_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _0983_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _0984_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _0985_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _0986_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0149_)
  );
  or_bb _0987_ (
    .a(_0149_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_35_)
  );
  maj_bbb _0988_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(b_34_)
  );
  and_bb _0989_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0148_)
  );
  and_bb _0990_ (
    .a(_0148_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_33_)
  );
  or_bb _0991_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0151_)
  );
  or_bb _0992_ (
    .a(_0151_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_32_)
  );
  maj_bbb _0993_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(b_31_)
  );
  and_bb _0994_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0150_)
  );
  and_bb _0995_ (
    .a(_0150_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_21_0__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_30_)
  );
  or_bb _0996_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_)
  );
  and_bb _0997_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_9_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_15_6__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_)
  );
  or_bb _0998_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_)
  );
  and_bb _0999_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_10_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_16_7__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_)
  );
  or_bb _1000_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_)
  );
  and_bb _1001_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_11_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_17_8__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_)
  );
  or_bb _1002_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_)
  );
  and_bb _1003_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_12_3__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_18_9__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_)
  );
  or_bb _1004_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_)
  );
  and_bb _1005_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_13_4__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_19_10__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_)
  );
  or_bb _1006_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_)
  );
  and_bb _1007_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_14_5__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_10_20_11__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_)
  );
  or_bb _1008_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_)
  );
  and_bb _1009_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_)
  );
  or_bb _1010_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_)
  );
  and_bb _1011_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_)
  );
  or_bb _1012_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_)
  );
  and_bb _1013_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_0_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_)
  );
  or_bb _1014_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0153_)
  );
  or_bb _1015_ (
    .a(_0153_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_41_)
  );
  maj_bbb _1016_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .d(b_40_)
  );
  and_bb _1017_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_5_),
    .c(_0152_)
  );
  and_bb _1018_ (
    .a(_0152_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_3_),
    .c(b_39_)
  );
  or_bb _1019_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0155_)
  );
  or_bb _1020_ (
    .a(_0155_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_38_)
  );
  maj_bbb _1021_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .d(b_37_)
  );
  and_bb _1022_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_2_),
    .c(_0154_)
  );
  and_bb _1023_ (
    .a(_0154_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_7_0__m_c_0_),
    .c(b_36_)
  );
  or_bb _1024_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_)
  );
  and_bb _1025_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_3_2__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_6_5__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_)
  );
  or_bb _1026_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_)
  );
  and_bb _1027_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_2_1__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_5_4__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_)
  );
  or_bb _1028_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_)
  );
  and_bb _1029_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_1_0__g_ord_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_10_4_3__g_ord_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_)
  );
  or_bb _1030_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0157_)
  );
  or_bb _1031_ (
    .a(_0157_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_47_)
  );
  maj_bbb _1032_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .d(b_46_)
  );
  and_bb _1033_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_4_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_5_),
    .c(_0156_)
  );
  and_bb _1034_ (
    .a(_0156_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_3_),
    .c(b_45_)
  );
  or_bb _1035_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0159_)
  );
  or_bb _1036_ (
    .a(_0159_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_44_)
  );
  maj_bbb _1037_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .c(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .d(b_43_)
  );
  and_bb _1038_ (
    .a(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_1_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_2_),
    .c(_0158_)
  );
  and_bb _1039_ (
    .a(_0158_),
    .b(_m__genblock___src_b48s_merger48_v_13_48_1__m__genblock___src_b48s_merger24_v_13_22_1__m__genblock___src_b48s_merger12_v_13_8_1__m_c_0_),
    .c(b_42_)
  );
endmodule
