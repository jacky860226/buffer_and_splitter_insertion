module c2670(G131,G26,G16,G30,G57,G12,G73,G147,G107,G75,G103,G141,G24,G62,G27,G76,G123,G4,G142,G118,G133,G150,G145,G39,G94,G19,G5,G152,G23,G96,G110,G120,G112,G47,G82,G157,G91,G106,G56,G13,G60,G148,G64,G20,G52,G8,G98,G11,G32,G66,G14,G143,G146,G28,G83,G108,G42,G3,G63,G144,G84,G87,G104,G132,G80,G36,G10,G54,G59,G92,G72,G79,G117,G31,G113,G116,G44,G1,G65,G154,G124,G55,G137,G38,G105,G61,G119,G90,G33,G22,G35,G115,G134,G40,G2,G25,G58,G111,G100,G126,G70,G9,G149,G121,G48,G78,G136,G43,G7,G81,G140,G89,G77,G95,G34,G99,G68,G67,G86,G15,G122,G45,G129,G18,G6,G93,G101,G125,G69,G114,G139,G97,G51,G109,G17,G74,G156,G153,G50,G138,G135,G71,G85,G155,G53,G37,G130,G46,G41,G49,G127,G102,G128,G151,G21,G88,G29);
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_2581;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_2742;
    wire new_Jinkela_wire_1987;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_1198;
    wire _0172_;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_1948;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_2354;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_1913;
    wire _0466_;
    wire _0166_;
    wire new_Jinkela_wire_2345;
    wire new_Jinkela_wire_2274;
    wire new_Jinkela_wire_2537;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_2098;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_2545;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_564;
    wire _0054_;
    wire new_Jinkela_wire_1892;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_2656;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_1886;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_505;
    wire _0149_;
    wire new_Jinkela_wire_1425;
    wire _0478_;
    wire new_Jinkela_wire_633;
    wire _0458_;
    wire new_Jinkela_wire_2306;
    wire new_Jinkela_wire_1273;
    wire _0137_;
    wire _0084_;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_1996;
    wire new_Jinkela_wire_2359;
    wire new_Jinkela_wire_531;
    wire _0385_;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_2367;
    wire _0322_;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_2129;
    wire new_Jinkela_wire_1840;
    wire _0118_;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_1702;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_1801;
    wire new_Jinkela_wire_2434;
    wire _0394_;
    wire new_Jinkela_wire_1945;
    wire new_Jinkela_wire_761;
    wire _0144_;
    wire new_Jinkela_wire_397;
    wire _0276_;
    wire new_Jinkela_wire_364;
    wire _0071_;
    wire _0354_;
    wire new_Jinkela_wire_516;
    wire _0160_;
    wire new_Jinkela_wire_1309;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_2170;
    wire new_Jinkela_wire_224;
    wire _0267_;
    wire new_Jinkela_wire_1417;
    wire _0482_;
    wire new_Jinkela_wire_1231;
    wire _0415_;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_2121;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_2270;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_2580;
    wire new_Jinkela_wire_1764;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_2163;
    wire new_Jinkela_wire_2741;
    wire new_Jinkela_wire_2125;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_2316;
    wire new_Jinkela_wire_2224;
    wire new_Jinkela_wire_2498;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_2207;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_2177;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_2086;
    wire new_Jinkela_wire_1871;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_1055;
    wire _0083_;
    wire new_Jinkela_wire_310;
    wire _0022_;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_2673;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_1246;
    wire _0079_;
    wire _0436_;
    wire _0465_;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_2171;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_1054;
    wire _0308_;
    wire new_Jinkela_wire_2501;
    wire new_Jinkela_wire_2607;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_775;
    wire _0437_;
    wire _0049_;
    wire new_Jinkela_wire_1815;
    wire _0368_;
    wire new_Jinkela_wire_2230;
    wire new_Jinkela_wire_2089;
    wire _0460_;
    wire new_Jinkela_wire_2495;
    wire _0377_;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_1073;
    wire _0027_;
    wire new_Jinkela_wire_2332;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_1722;
    wire _0113_;
    wire _0496_;
    wire new_Jinkela_wire_1530;
    wire _0375_;
    wire new_Jinkela_wire_2703;
    wire _0284_;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_1197;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_2078;
    wire _0185_;
    wire new_Jinkela_wire_1666;
    wire _0381_;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_1589;
    wire new_net_957;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_2720;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_2586;
    wire new_Jinkela_wire_1848;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_2167;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_2388;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_2470;
    wire _0090_;
    wire new_Jinkela_wire_1548;
    wire _0195_;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_596;
    wire _0074_;
    wire _0311_;
    wire new_Jinkela_wire_2410;
    wire new_Jinkela_wire_1951;
    wire new_Jinkela_wire_2382;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_2395;
    wire _0196_;
    wire _0175_;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_2540;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_2513;
    wire _0039_;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_1978;
    wire _0471_;
    wire new_Jinkela_wire_1866;
    wire _0259_;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_1757;
    wire new_Jinkela_wire_1906;
    wire new_Jinkela_wire_2408;
    wire new_Jinkela_wire_2261;
    wire new_Jinkela_wire_2642;
    wire _0101_;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_1469;
    wire _0213_;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_303;
    wire _0023_;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_2709;
    wire _0036_;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_247;
    wire _0016_;
    wire new_Jinkela_wire_1807;
    wire new_Jinkela_wire_1949;
    wire new_Jinkela_wire_2119;
    wire new_Jinkela_wire_2304;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_1994;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_2618;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_802;
    wire _0232_;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_1648;
    wire _0180_;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_199;
    wire new_net_12;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_2281;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_1426;
    wire _0307_;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_2605;
    wire new_Jinkela_wire_1234;
    wire new_Jinkela_wire_2360;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_2239;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_2533;
    wire _0491_;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_2530;
    wire new_Jinkela_wire_2363;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_2403;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_2471;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_1478;
    wire _0205_;
    wire _0064_;
    wire new_Jinkela_wire_1043;
    wire _0188_;
    wire new_Jinkela_wire_2362;
    wire new_Jinkela_wire_386;
    wire _0356_;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_1292;
    wire _0189_;
    wire new_Jinkela_wire_1299;
    wire _0461_;
    wire new_Jinkela_wire_1809;
    wire _0353_;
    wire new_Jinkela_wire_2223;
    wire new_Jinkela_wire_2600;
    wire new_Jinkela_wire_2227;
    wire new_Jinkela_wire_774;
    wire _0233_;
    wire new_Jinkela_wire_2191;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_2209;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_2241;
    wire new_Jinkela_wire_1045;
    wire _0382_;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_2014;
    wire _0085_;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_523;
    wire new_net_23;
    wire _0140_;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_430;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_1302;
    wire _0407_;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_2424;
    wire new_net_16;
    wire new_Jinkela_wire_2292;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_2494;
    wire new_Jinkela_wire_1832;
    wire new_Jinkela_wire_186;
    wire _0357_;
    wire new_Jinkela_wire_530;
    wire _0114_;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_2738;
    wire new_Jinkela_wire_2213;
    wire new_Jinkela_wire_2551;
    wire new_Jinkela_wire_1566;
    wire _0152_;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_2546;
    wire _0450_;
    wire _0141_;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_2111;
    wire new_Jinkela_wire_2100;
    wire new_Jinkela_wire_1693;
    wire new_Jinkela_wire_2131;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_2142;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_2390;
    wire new_Jinkela_wire_2257;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_2228;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_29;
    wire _0235_;
    wire _0402_;
    wire new_Jinkela_wire_1077;
    wire _0040_;
    wire new_Jinkela_wire_1148;
    wire _0475_;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_1286;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_2222;
    wire new_Jinkela_wire_2406;
    wire _0334_;
    wire _0319_;
    wire new_Jinkela_wire_714;
    wire _0246_;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_2597;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_2481;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_1859;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_2562;
    wire _0253_;
    wire new_Jinkela_wire_2601;
    wire new_Jinkela_wire_464;
    wire _0315_;
    wire _0431_;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_61;
    wire _0161_;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_2594;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_2187;
    wire _0147_;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_2611;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_1657;
    wire new_Jinkela_wire_2095;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_753;
    wire _0350_;
    wire new_Jinkela_wire_1057;
    wire _0058_;
    wire new_Jinkela_wire_2200;
    wire new_Jinkela_wire_1748;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_2476;
    wire new_Jinkela_wire_2739;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_2364;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_2589;
    wire new_Jinkela_wire_1408;
    wire new_net_19;
    wire new_Jinkela_wire_2330;
    wire new_Jinkela_wire_2030;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_2450;
    wire _0164_;
    wire new_Jinkela_wire_2500;
    wire _0265_;
    wire _0433_;
    wire new_Jinkela_wire_821;
    wire _0248_;
    wire new_Jinkela_wire_23;
    wire _0104_;
    wire new_Jinkela_wire_2287;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_1450;
    wire new_Jinkela_wire_2717;
    wire new_Jinkela_wire_2351;
    wire new_Jinkela_wire_1797;
    wire _0182_;
    wire new_Jinkela_wire_1874;
    wire _0229_;
    wire new_Jinkela_wire_2347;
    wire new_Jinkela_wire_282;
    wire _0223_;
    wire new_Jinkela_wire_1729;
    wire new_Jinkela_wire_2324;
    wire new_Jinkela_wire_1904;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_2457;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_1661;
    wire _0299_;
    wire new_Jinkela_wire_547;
    wire _0187_;
    wire new_Jinkela_wire_2454;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_2295;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_1855;
    wire _0449_;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_2103;
    wire _0048_;
    wire new_Jinkela_wire_2714;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_2320;
    wire new_Jinkela_wire_2381;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_2517;
    wire new_Jinkela_wire_2271;
    wire new_net_9;
    wire _0228_;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_284;
    wire _0176_;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_2389;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_2070;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_893;
    wire _0293_;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_2596;
    wire new_Jinkela_wire_2053;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_2458;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_2293;
    wire new_Jinkela_wire_215;
    wire new_net_963;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_1209;
    wire _0168_;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_2711;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_2196;
    wire new_Jinkela_wire_2352;
    wire new_Jinkela_wire_1498;
    wire _0279_;
    wire _0454_;
    wire new_Jinkela_wire_2158;
    wire new_Jinkela_wire_2083;
    wire _0111_;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_2299;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_2333;
    wire _0490_;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_2045;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_1063;
    wire _0287_;
    wire new_Jinkela_wire_453;
    wire _0224_;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_325;
    wire _0422_;
    wire new_Jinkela_wire_2743;
    wire _0328_;
    wire _0217_;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_2654;
    wire new_Jinkela_wire_2432;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_2521;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_2216;
    wire new_Jinkela_wire_33;
    wire _0183_;
    wire new_Jinkela_wire_2526;
    wire new_Jinkela_wire_1802;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_1297;
    wire _0405_;
    wire new_Jinkela_wire_2563;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_2604;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_1208;
    wire _0397_;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_2184;
    wire new_Jinkela_wire_2331;
    wire new_Jinkela_wire_1224;
    wire _0095_;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_2520;
    wire new_Jinkela_wire_2685;
    wire new_Jinkela_wire_2062;
    wire new_Jinkela_wire_2544;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_1655;
    wire _0102_;
    wire new_Jinkela_wire_2626;
    wire new_Jinkela_wire_2350;
    wire new_Jinkela_wire_2539;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_2164;
    wire _0121_;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_2523;
    wire _0480_;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_2181;
    wire new_Jinkela_wire_305;
    wire _0303_;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_425;
    wire _0272_;
    wire _0348_;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_1751;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_1037;
    wire _0236_;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_2679;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_2426;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_2559;
    wire new_Jinkela_wire_2116;
    wire new_Jinkela_wire_891;
    wire _0262_;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_2734;
    wire new_Jinkela_wire_2252;
    wire new_Jinkela_wire_2134;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_2578;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_1591;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_2620;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_2669;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_1930;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_1326;
    wire _0399_;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_2726;
    wire new_Jinkela_wire_133;
    wire _0212_;
    wire new_Jinkela_wire_111;
    wire _0295_;
    wire new_Jinkela_wire_1343;
    wire _0421_;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_1775;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_2250;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_137;
    wire _0379_;
    wire new_Jinkela_wire_2650;
    wire _0032_;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_1503;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_2197;
    wire new_Jinkela_wire_1400;
    wire _0179_;
    wire _0192_;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_273;
    wire _0283_;
    wire new_Jinkela_wire_610;
    wire _0139_;
    wire _0390_;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_2102;
    wire new_Jinkela_wire_2694;
    wire new_Jinkela_wire_2627;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_151;
    wire _0472_;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_2534;
    wire new_Jinkela_wire_2325;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_1626;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_1295;
    wire _0280_;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_490;
    wire _0004_;
    wire new_Jinkela_wire_2416;
    wire new_Jinkela_wire_651;
    wire _0477_;
    wire new_Jinkela_wire_2277;
    wire new_Jinkela_wire_2591;
    wire new_net_961;
    wire new_Jinkela_wire_1284;
    wire new_Jinkela_wire_1817;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_2297;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_1089;
    wire _0332_;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_617;
    wire _0369_;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_2254;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_1697;
    wire new_Jinkela_wire_2737;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_1856;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_2603;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_2629;
    wire _0474_;
    wire _0199_;
    wire new_Jinkela_wire_2017;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_2361;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_2397;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_2077;
    wire new_Jinkela_wire_2114;
    wire _0201_;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_2524;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_2641;
    wire _0252_;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_2074;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_2088;
    wire new_Jinkela_wire_1403;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_2161;
    wire new_Jinkela_wire_1819;
    wire new_Jinkela_wire_2051;
    wire new_Jinkela_wire_1585;
    wire _0157_;
    wire new_Jinkela_wire_2695;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_477;
    wire _0463_;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_2414;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_2508;
    wire new_Jinkela_wire_2689;
    wire new_Jinkela_wire_642;
    wire _0154_;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_1963;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_2326;
    wire _0202_;
    wire _0030_;
    wire _0070_;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_2391;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_559;
    wire _0414_;
    wire new_Jinkela_wire_1294;
    wire new_Jinkela_wire_2236;
    wire new_Jinkela_wire_2576;
    wire new_Jinkela_wire_1806;
    wire _0479_;
    wire new_Jinkela_wire_2282;
    wire new_Jinkela_wire_2154;
    wire _0150_;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_2725;
    wire _0026_;
    wire new_Jinkela_wire_2421;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_2674;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_2728;
    wire _0488_;
    wire new_Jinkela_wire_2105;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_2662;
    wire new_Jinkela_wire_1776;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_2305;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_2491;
    wire new_Jinkela_wire_264;
    wire _0301_;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_436;
    wire _0274_;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_1960;
    wire new_Jinkela_wire_2387;
    wire new_Jinkela_wire_327;
    wire _0258_;
    wire new_Jinkela_wire_345;
    wire _0062_;
    wire new_Jinkela_wire_2411;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_2251;
    wire new_Jinkela_wire_2335;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_1860;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_1066;
    wire _0204_;
    wire new_Jinkela_wire_2084;
    wire _0338_;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_2484;
    wire new_Jinkela_wire_2356;
    wire new_Jinkela_wire_1398;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_2379;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_2210;
    wire _0325_;
    wire new_Jinkela_wire_162;
    wire _0128_;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_1332;
    wire new_net_15;
    wire new_Jinkela_wire_1202;
    wire _0237_;
    wire new_Jinkela_wire_2489;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_26;
    wire _0041_;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_863;
    wire _0419_;
    wire new_Jinkela_wire_2380;
    wire new_Jinkela_wire_2211;
    wire new_Jinkela_wire_806;
    wire _0254_;
    wire _0126_;
    wire _0190_;
    wire new_Jinkela_wire_2465;
    wire _0193_;
    wire new_Jinkela_wire_1630;
    wire _0153_;
    wire new_Jinkela_wire_1262;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_1611;
    wire _0082_;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_2423;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_1531;
    wire _0124_;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_293;
    wire _0286_;
    wire new_Jinkela_wire_2401;
    wire new_Jinkela_wire_1880;
    wire _0309_;
    wire new_Jinkela_wire_2430;
    wire new_Jinkela_wire_2071;
    wire new_Jinkela_wire_2718;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_2055;
    wire new_Jinkela_wire_812;
    wire _0456_;
    wire new_Jinkela_wire_999;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_1166;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_2143;
    wire _0302_;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_1093;
    wire _0349_;
    wire new_Jinkela_wire_2355;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_2664;
    wire new_Jinkela_wire_1822;
    wire _0241_;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_2203;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_2182;
    wire new_Jinkela_wire_2038;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_1870;
    wire new_Jinkela_wire_2085;
    wire new_Jinkela_wire_2731;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_2001;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_1114;
    wire _0029_;
    wire new_Jinkela_wire_2366;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_2340;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_2640;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_2050;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_1938;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_2455;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_1749;
    wire _0194_;
    wire _0234_;
    wire new_Jinkela_wire_2740;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_263;
    wire _0266_;
    wire new_Jinkela_wire_2269;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_489;
    wire _0073_;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_2469;
    wire new_Jinkela_wire_2499;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_2291;
    wire new_Jinkela_wire_2561;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_1720;
    wire _0469_;
    wire new_Jinkela_wire_2686;
    wire new_Jinkela_wire_2486;
    wire new_Jinkela_wire_2516;
    wire new_Jinkela_wire_2173;
    wire _0365_;
    wire new_Jinkela_wire_959;
    wire _0197_;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_1725;
    wire _0052_;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_2464;
    wire new_Jinkela_wire_2623;
    wire _0094_;
    wire new_Jinkela_wire_1170;
    wire _0091_;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_2478;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_2374;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_2028;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_1853;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_2349;
    wire new_Jinkela_wire_2377;
    wire _0255_;
    wire new_Jinkela_wire_2612;
    wire new_Jinkela_wire_1600;
    wire _0010_;
    wire new_Jinkela_wire_2064;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_2052;
    wire _0015_;
    wire new_Jinkela_wire_2185;
    wire new_Jinkela_wire_2529;
    wire new_Jinkela_wire_790;
    wire _0467_;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_2599;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_1918;
    wire _0489_;
    wire new_Jinkela_wire_1553;
    wire _0412_;
    wire new_Jinkela_wire_2156;
    wire new_Jinkela_wire_1857;
    wire new_Jinkela_wire_955;
    wire _0420_;
    wire new_Jinkela_wire_739;
    wire _0416_;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_2487;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_1391;
    wire _0169_;
    wire _0392_;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_511;
    wire _0321_;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_2568;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_2592;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_2300;
    wire new_Jinkela_wire_1761;
    wire _0100_;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_2441;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_2420;
    wire new_Jinkela_wire_2730;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_2106;
    wire new_Jinkela_wire_2687;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_2059;
    wire new_Jinkela_wire_1997;
    wire new_net_1;
    wire new_Jinkela_wire_2643;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_2485;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_2547;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_913;
    wire _0323_;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_496;
    wire _0340_;
    wire new_Jinkela_wire_2567;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_2264;
    wire new_Jinkela_wire_1990;
    wire new_Jinkela_wire_2101;
    wire new_Jinkela_wire_2671;
    wire new_Jinkela_wire_1908;
    wire _0358_;
    wire new_Jinkela_wire_1675;
    wire _0317_;
    wire new_Jinkela_wire_2502;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_2370;
    wire new_net_950;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_2394;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_1485;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_1698;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_1358;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_1671;
    wire new_Jinkela_wire_1924;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_1746;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_2160;
    wire _0362_;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_480;
    wire _0186_;
    wire new_Jinkela_wire_2638;
    wire new_Jinkela_wire_1672;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_1888;
    wire new_Jinkela_wire_1544;
    wire _0441_;
    wire new_Jinkela_wire_2667;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_967;
    wire _0447_;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_1393;
    wire _0210_;
    wire new_net_6;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_2039;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_2268;
    wire new_Jinkela_wire_2091;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_2319;
    wire _0261_;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_2107;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_2194;
    wire new_Jinkela_wire_581;
    wire _0045_;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_1727;
    wire _0434_;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_2296;
    wire _0208_;
    wire _0438_;
    wire new_Jinkela_wire_1847;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_2698;
    wire new_Jinkela_wire_972;
    wire _0406_;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_1146;
    wire _0485_;
    wire new_Jinkela_wire_1097;
    wire _0002_;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_339;
    wire _0117_;
    wire new_Jinkela_wire_706;
    wire _0345_;
    wire _0427_;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_1967;
    wire new_Jinkela_wire_2063;
    wire new_Jinkela_wire_2564;
    wire new_Jinkela_wire_1771;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_1935;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_2453;
    wire new_Jinkela_wire_2385;
    wire _0214_;
    wire new_Jinkela_wire_2307;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_2445;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_2630;
    wire new_Jinkela_wire_2670;
    wire new_Jinkela_wire_2644;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_2602;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_2702;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_1737;
    wire new_Jinkela_wire_2309;
    wire _0296_;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_136;
    wire _0053_;
    wire new_Jinkela_wire_2721;
    wire new_Jinkela_wire_2384;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_1844;
    wire new_Jinkela_wire_2479;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_2637;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_930;
    wire _0359_;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_413;
    wire _0206_;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_1140;
    wire _0264_;
    wire new_Jinkela_wire_377;
    wire _0148_;
    wire new_Jinkela_wire_2249;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_1872;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_1741;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_2205;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_2049;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_1882;
    wire _0108_;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_1931;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_2691;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_1884;
    wire _0037_;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_1015;
    wire _0155_;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_2165;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_209;
    wire _0051_;
    wire new_Jinkela_wire_2214;
    wire new_Jinkela_wire_2127;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_2506;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_1647;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_2323;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_1972;
    wire new_Jinkela_wire_2536;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_2631;
    wire new_Jinkela_wire_2248;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_2431;
    wire _0231_;
    wire new_Jinkela_wire_2652;
    wire new_Jinkela_wire_2262;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_2066;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_2336;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_2449;
    wire new_Jinkela_wire_2183;
    wire new_Jinkela_wire_1705;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_1829;
    wire new_Jinkela_wire_2482;
    wire new_Jinkela_wire_2159;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_2727;
    wire new_Jinkela_wire_2120;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_2219;
    wire new_Jinkela_wire_2462;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_2505;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_178;
    wire new_net_7;
    wire new_Jinkela_wire_1099;
    wire _0209_;
    wire _0110_;
    wire _0336_;
    wire new_Jinkela_wire_1390;
    wire _0120_;
    wire new_Jinkela_wire_2619;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_2582;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_1567;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_2108;
    wire _0013_;
    wire _0138_;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_2697;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_2701;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_2609;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_2548;
    wire new_Jinkela_wire_2267;
    wire _0089_;
    wire new_Jinkela_wire_2090;
    wire new_Jinkela_wire_469;
    wire new_net_14;
    wire new_Jinkela_wire_1554;
    wire _0050_;
    wire new_Jinkela_wire_2079;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_2452;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_951;
    wire _0009_;
    wire new_Jinkela_wire_1656;
    wire new_Jinkela_wire_446;
    wire new_net_21;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_2735;
    wire new_Jinkela_wire_2338;
    wire _0446_;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_1490;
    wire _0351_;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_2369;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_1339;
    wire _0005_;
    wire new_Jinkela_wire_1421;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_2229;
    wire _0055_;
    wire new_Jinkela_wire_2456;
    wire _0203_;
    wire new_Jinkela_wire_2511;
    wire new_Jinkela_wire_2290;
    wire new_Jinkela_wire_2712;
    wire _0006_;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_2193;
    wire new_Jinkela_wire_329;
    wire _0271_;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_2719;
    wire new_Jinkela_wire_1207;
    wire _0256_;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_1515;
    wire _0318_;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_2443;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_2314;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_2005;
    wire _0035_;
    wire new_Jinkela_wire_2528;
    wire new_Jinkela_wire_2372;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_1346;
    wire _0355_;
    wire new_Jinkela_wire_2660;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_1230;
    wire _0484_;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_506;
    wire _0497_;
    wire new_Jinkela_wire_2556;
    wire _0398_;
    wire new_Jinkela_wire_850;
    wire _0268_;
    wire _0125_;
    wire new_Jinkela_wire_1915;
    wire _0207_;
    wire new_Jinkela_wire_2615;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_2075;
    wire new_Jinkela_wire_2146;
    wire _0245_;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_2035;
    wire new_Jinkela_wire_1726;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_2009;
    wire new_Jinkela_wire_2477;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_722;
    wire _0096_;
    wire new_Jinkela_wire_2118;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_2585;
    wire new_Jinkela_wire_2122;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_2301;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_2583;
    wire new_Jinkela_wire_1744;
    wire _0170_;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_2018;
    wire new_Jinkela_wire_1942;
    wire _0483_;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_2240;
    wire new_Jinkela_wire_1076;
    wire _0059_;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_79;
    wire _0000_;
    wire new_Jinkela_wire_2149;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_2393;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_2130;
    wire new_Jinkela_wire_1333;
    wire new_Jinkela_wire_1954;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_2375;
    wire _0285_;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_2696;
    wire _0165_;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_2099;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_665;
    wire _0393_;
    wire new_Jinkela_wire_2493;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_2560;
    wire _0078_;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_372;
    wire _0373_;
    wire new_Jinkela_wire_717;
    wire new_net_20;
    wire new_Jinkela_wire_835;
    wire _0320_;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_2418;
    wire new_Jinkela_wire_2202;
    wire new_net_959;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_1724;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_2004;
    wire new_Jinkela_wire_2398;
    wire new_Jinkela_wire_2234;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_2437;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_1468;
    wire _0352_;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_1895;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_2298;
    wire new_Jinkela_wire_1264;
    wire _0298_;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_2613;
    wire _0403_;
    wire _0076_;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_675;
    wire _0220_;
    wire _0065_;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_2598;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_56;
    wire _0281_;
    wire new_Jinkela_wire_2123;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_834;
    wire _0011_;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_135;
    wire _0107_;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_1975;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_760;
    wire new_net_954;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_2668;
    wire new_Jinkela_wire_2610;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_2273;
    wire new_Jinkela_wire_2634;
    wire new_Jinkela_wire_2557;
    wire new_Jinkela_wire_1156;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_2094;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_2247;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_2558;
    wire new_Jinkela_wire_1966;
    wire _0056_;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_2549;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_827;
    wire _0417_;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_647;
    wire _0097_;
    wire new_Jinkela_wire_2342;
    wire new_Jinkela_wire_894;
    wire new_net_5;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_1407;
    wire _0316_;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_1215;
    wire _0424_;
    wire new_Jinkela_wire_1178;
    wire new_Jinkela_wire_2115;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_1780;
    wire new_Jinkela_wire_1687;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_2082;
    wire _0495_;
    wire new_Jinkela_wire_2645;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_1068;
    wire _0343_;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_388;
    wire _0297_;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_2192;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_1627;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_2417;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_1020;
    wire new_net_948;
    wire _0443_;
    wire new_Jinkela_wire_2699;
    wire new_Jinkela_wire_1712;
    wire new_Jinkela_wire_41;
    wire _0230_;
    wire new_Jinkela_wire_627;
    wire _0198_;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_2136;
    wire new_Jinkela_wire_150;
    wire new_Jinkela_wire_705;
    wire _0386_;
    wire new_Jinkela_wire_2543;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_1955;
    wire new_Jinkela_wire_1717;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_2152;
    wire new_Jinkela_wire_2633;
    wire new_Jinkela_wire_2438;
    wire new_Jinkela_wire_2072;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_1767;
    wire new_Jinkela_wire_2334;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_2279;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_1878;
    wire _0003_;
    wire new_Jinkela_wire_2678;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_2665;
    wire new_Jinkela_wire_1939;
    wire new_Jinkela_wire_2683;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_1145;
    wire new_Jinkela_wire_1719;
    wire new_Jinkela_wire_1709;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_764;
    wire _0021_;
    wire new_Jinkela_wire_646;
    wire _0305_;
    wire new_Jinkela_wire_1800;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_13;
    wire _0388_;
    wire _0063_;
    wire new_Jinkela_wire_2276;
    wire _0270_;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_2724;
    wire new_Jinkela_wire_852;
    wire _0077_;
    wire _0314_;
    wire _0225_;
    wire new_Jinkela_wire_1893;
    wire _0292_;
    wire new_Jinkela_wire_2507;
    wire _0413_;
    wire new_Jinkela_wire_2413;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_2218;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_1713;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_2483;
    wire new_Jinkela_wire_2180;
    wire _0086_;
    wire new_Jinkela_wire_970;
    wire _0442_;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_895;
    wire new_Jinkela_wire_1921;
    wire _0163_;
    wire _0024_;
    wire _0012_;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_2068;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_1900;
    wire new_Jinkela_wire_2436;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_1379;
    wire _0017_;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_2343;
    wire new_Jinkela_wire_2056;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_2700;
    wire new_Jinkela_wire_2512;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_2392;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_981;
    wire new_net_18;
    wire new_Jinkela_wire_2407;
    wire new_Jinkela_wire_2373;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_1755;
    wire new_Jinkela_wire_692;
    wire _0075_;
    wire new_Jinkela_wire_1392;
    wire _0363_;
    wire new_Jinkela_wire_261;
    wire _0389_;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_2723;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_2310;
    wire new_Jinkela_wire_2303;
    wire new_Jinkela_wire_2172;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_2632;
    wire new_Jinkela_wire_2126;
    wire _0327_;
    wire new_Jinkela_wire_2624;
    wire new_Jinkela_wire_2117;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_1463;
    wire _0240_;
    wire new_Jinkela_wire_1036;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_1141;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_80;
    wire _0184_;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_2574;
    wire _0370_;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_2617;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_2327;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1438;
    wire _0360_;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_2571;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_1739;
    wire new_Jinkela_wire_2575;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_2628;
    wire _0429_;
    wire new_Jinkela_wire_2186;
    wire new_Jinkela_wire_76;
    wire _0300_;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_2584;
    wire new_Jinkela_wire_1506;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_1781;
    wire new_Jinkela_wire_2621;
    wire new_Jinkela_wire_2428;
    wire new_Jinkela_wire_2376;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_820;
    wire _0109_;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_2636;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_1754;
    wire _0033_;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_428;
    wire _0339_;
    wire _0131_;
    wire new_Jinkela_wire_2474;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_2729;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_2446;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_2015;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_2532;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_1605;
    wire _0066_;
    wire new_Jinkela_wire_2087;
    wire new_Jinkela_wire_2473;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_1792;
    wire new_Jinkela_wire_93;
    wire _0025_;
    wire _0409_;
    wire new_Jinkela_wire_2255;
    wire new_net_967;
    wire new_Jinkela_wire_2027;
    wire new_Jinkela_wire_2104;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_1957;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_678;
    wire _0167_;
    wire new_Jinkela_wire_2141;
    wire new_Jinkela_wire_2258;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_2308;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_708;
    wire _0344_;
    wire new_Jinkela_wire_2442;
    wire new_Jinkela_wire_2415;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_64;
    wire _0342_;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_1201;
    wire _0060_;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_2346;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_1514;
    wire _0331_;
    wire new_Jinkela_wire_2593;
    wire new_Jinkela_wire_1862;
    wire new_Jinkela_wire_1977;
    wire new_Jinkela_wire_1934;
    wire new_Jinkela_wire_2217;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_486;
    wire _0249_;
    wire new_Jinkela_wire_1549;
    wire new_net_952;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_2684;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_2672;
    wire new_Jinkela_wire_1786;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_1943;
    wire new_Jinkela_wire_1612;
    wire new_Jinkela_wire_2378;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_2080;
    wire new_Jinkela_wire_2402;
    wire new_Jinkela_wire_2448;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_2460;
    wire new_Jinkela_wire_2265;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_2317;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_2399;
    wire new_Jinkela_wire_2625;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_1258;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_1445;
    wire new_Jinkela_wire_976;
    wire _0239_;
    wire new_Jinkela_wire_2608;
    wire new_Jinkela_wire_2736;
    wire new_Jinkela_wire_1867;
    wire _0263_;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_2174;
    wire _0135_;
    wire new_Jinkela_wire_699;
    wire _0468_;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_2162;
    wire new_Jinkela_wire_1265;
    wire _0156_;
    wire new_Jinkela_wire_2368;
    wire new_Jinkela_wire_2409;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_1251;
    wire _0378_;
    wire new_Jinkela_wire_555;
    wire _0452_;
    wire new_Jinkela_wire_2463;
    wire new_Jinkela_wire_2033;
    wire _0238_;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_1691;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_2522;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_1823;
    wire new_Jinkela_wire_984;
    wire _0411_;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_2065;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_2677;
    wire new_Jinkela_wire_2212;
    wire new_Jinkela_wire_1135;
    wire _0435_;
    wire _0211_;
    wire _0067_;
    wire _0439_;
    wire new_Jinkela_wire_1419;
    wire _0068_;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_2461;
    wire _0455_;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_2034;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_2312;
    wire new_Jinkela_wire_440;
    wire _0008_;
    wire new_Jinkela_wire_2348;
    wire _0380_;
    wire new_net_3;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_2344;
    wire _0494_;
    wire _0423_;
    wire new_Jinkela_wire_2459;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_2266;
    wire new_Jinkela_wire_1843;
    wire new_Jinkela_wire_2412;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_861;
    wire _0127_;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_2383;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_2622;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_836;
    wire _0191_;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_558;
    wire _0451_;
    wire new_Jinkela_wire_1405;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_1984;
    wire _0219_;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_2515;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_241;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_2315;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_1916;
    wire new_Jinkela_wire_2693;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_814;
    wire _0115_;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_2480;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_1383;
    wire _0384_;
    wire _0313_;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_1953;
    wire new_Jinkela_wire_312;
    wire _0400_;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_2113;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_916;
    wire _0181_;
    wire new_Jinkela_wire_1050;
    wire new_net_965;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_2550;
    wire new_Jinkela_wire_1742;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_2708;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_1649;
    wire _0250_;
    wire new_net_13;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_2682;
    wire new_Jinkela_wire_2496;
    wire new_Jinkela_wire_2016;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_2244;
    wire new_Jinkela_wire_1969;
    wire new_Jinkela_wire_1187;
    wire new_net_4;
    wire new_Jinkela_wire_2444;
    wire new_Jinkela_wire_366;
    wire _0289_;
    wire new_Jinkela_wire_548;
    wire _0432_;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_2097;
    wire _0376_;
    wire new_Jinkela_wire_873;
    wire _0487_;
    wire _0290_;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_2043;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_1743;
    wire _0440_;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_2215;
    wire _0288_;
    wire new_Jinkela_wire_2488;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_2552;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_2490;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_2246;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_2339;
    wire _0444_;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_2124;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_28;
    wire _0244_;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_2541;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_2579;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_1723;
    wire _0282_;
    wire new_Jinkela_wire_2206;
    wire _0099_;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_174;
    wire _0069_;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_2358;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_1546;
    wire _0418_;
    wire _0047_;
    wire _0372_;
    wire new_Jinkela_wire_2144;
    wire new_Jinkela_wire_2566;
    wire new_Jinkela_wire_2337;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_1989;
    wire new_Jinkela_wire_1021;
    wire _0081_;
    wire new_Jinkela_wire_2048;
    wire new_Jinkela_wire_2318;
    wire _0106_;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_2658;
    wire new_Jinkela_wire_2577;
    wire new_Jinkela_wire_1266;
    wire _0080_;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_1803;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_2404;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_2733;
    wire _0291_;
    wire new_Jinkela_wire_1117;
    wire _0130_;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_1899;
    wire new_Jinkela_wire_2199;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_2073;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_2675;
    wire new_Jinkela_wire_2328;
    wire new_Jinkela_wire_2688;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_1413;
    wire _0178_;
    wire new_Jinkela_wire_1715;
    wire new_Jinkela_wire_825;
    wire _0018_;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_1040;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_2238;
    wire new_Jinkela_wire_1804;
    wire new_Jinkela_wire_1854;
    wire _0143_;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_2322;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_2427;
    wire _0457_;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_569;
    wire _0387_;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_1852;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_742;
    wire _0151_;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_2096;
    wire new_Jinkela_wire_2132;
    wire new_Jinkela_wire_498;
    wire new_net_11;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_2280;
    wire new_Jinkela_wire_2433;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_1779;
    wire new_Jinkela_wire_2286;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_1816;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_1110;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_1486;
    wire _0367_;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_2012;
    wire _0364_;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_886;
    wire _0014_;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_2663;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_2553;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_2157;
    wire new_Jinkela_wire_2357;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_2514;
    wire new_Jinkela_wire_2692;
    wire new_Jinkela_wire_1387;
    wire _0242_;
    wire new_Jinkela_wire_1765;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_1188;
    wire _0498_;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_2651;
    wire _0371_;
    wire new_Jinkela_wire_40;
    wire _0112_;
    wire new_Jinkela_wire_2329;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_1245;
    wire new_Jinkela_wire_2439;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_897;
    wire _0226_;
    wire new_Jinkela_wire_2590;
    wire new_Jinkela_wire_2151;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_427;
    wire _0374_;
    wire new_net_8;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_132;
    wire _0133_;
    wire new_Jinkela_wire_2635;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_1689;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_2195;
    wire new_Jinkela_wire_1889;
    wire new_Jinkela_wire_1003;
    wire _0116_;
    wire new_Jinkela_wire_121;
    wire _0326_;
    wire new_Jinkela_wire_1335;
    wire _0218_;
    wire _0044_;
    wire new_Jinkela_wire_2166;
    wire new_Jinkela_wire_925;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_1137;
    wire _0330_;
    wire new_Jinkela_wire_2647;
    wire new_Jinkela_wire_2176;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_2472;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_2289;
    wire new_Jinkela_wire_2067;
    wire new_Jinkela_wire_973;
    wire _0383_;
    wire new_Jinkela_wire_1051;
    wire _0142_;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_2288;
    wire new_Jinkela_wire_2178;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_586;
    wire _0088_;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_2659;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_2155;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_2242;
    wire new_Jinkela_wire_1907;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_2081;
    wire _0459_;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_2661;
    wire new_Jinkela_wire_1319;
    wire _0476_;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_2201;
    wire new_Jinkela_wire_2231;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_2150;
    wire _0257_;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_2278;
    wire new_Jinkela_wire_2648;
    wire _0404_;
    wire new_Jinkela_wire_1537;
    wire _0019_;
    wire new_Jinkela_wire_2093;
    wire new_Jinkela_wire_2497;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_2655;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_1420;
    wire new_Jinkela_wire_2371;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_2110;
    wire _0470_;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_2451;
    wire new_Jinkela_wire_1753;
    wire _0260_;
    wire new_Jinkela_wire_2396;
    wire _0173_;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_1973;
    wire new_Jinkela_wire_2565;
    wire new_Jinkela_wire_2706;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_83;
    wire _0247_;
    wire _0462_;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_2676;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_2168;
    wire _0007_;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_2527;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_2046;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_1151;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_2690;
    wire new_Jinkela_wire_1645;
    wire _0251_;
    wire _0277_;
    wire _0395_;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_2587;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_1883;
    wire new_Jinkela_wire_2208;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_1740;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_1436;
    wire new_Jinkela_wire_2284;
    wire new_Jinkela_wire_2226;
    wire new_net_17;
    wire new_Jinkela_wire_2057;
    wire new_Jinkela_wire_2225;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_172;
    wire _0473_;
    wire _0061_;
    wire _0042_;
    wire new_Jinkela_wire_2639;
    wire new_Jinkela_wire_1950;
    wire _0145_;
    wire new_Jinkela_wire_2135;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_2253;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_2419;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_1747;
    wire _0034_;
    wire _0273_;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_304;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_2002;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_2716;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_1896;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_1437;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_2353;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_2133;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_2148;
    wire new_Jinkela_wire_2681;
    wire new_Jinkela_wire_588;
    wire _0361_;
    wire new_Jinkela_wire_1243;
    wire _0092_;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_2710;
    wire new_Jinkela_wire_2572;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_1750;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_1125;
    wire _0425_;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_1833;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_2179;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_2147;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_2221;
    wire new_Jinkela_wire_2245;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_2569;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_2707;
    wire new_Jinkela_wire_2475;
    wire _0001_;
    wire new_Jinkela_wire_2145;
    wire new_Jinkela_wire_2243;
    wire new_Jinkela_wire_2235;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_2272;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_2010;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_869;
    wire _0132_;
    wire new_Jinkela_wire_1131;
    wire _0312_;
    wire _0492_;
    wire new_Jinkela_wire_2468;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_1570;
    wire _0410_;
    wire new_Jinkela_wire_2440;
    wire new_Jinkela_wire_124;
    wire _0129_;
    wire new_Jinkela_wire_2060;
    wire new_Jinkela_wire_2704;
    wire _0098_;
    wire new_Jinkela_wire_2237;
    wire _0119_;
    wire _0123_;
    wire _0174_;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_1252;
    wire new_Jinkela_wire_2666;
    wire _0408_;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_2732;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_1377;
    wire _0243_;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_1086;
    wire _0159_;
    wire new_Jinkela_wire_1861;
    wire _0493_;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_1660;
    wire _0333_;
    wire _0020_;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_2525;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_2061;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_2128;
    wire _0481_;
    wire new_Jinkela_wire_2275;
    wire new_Jinkela_wire_2233;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_1991;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_746;
    wire _0162_;
    wire new_Jinkela_wire_1517;
    wire _0426_;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_2535;
    wire new_Jinkela_wire_2510;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_2025;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_2519;
    wire new_Jinkela_wire_2538;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_2313;
    wire new_Jinkela_wire_1929;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_2058;
    wire _0093_;
    wire new_Jinkela_wire_1782;
    wire new_Jinkela_wire_2092;
    wire new_Jinkela_wire_823;
    wire _0329_;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_1688;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_1962;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_754;
    wire _0105_;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_1897;
    wire new_Jinkela_wire_2054;
    wire new_Jinkela_wire_1993;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_1818;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_843;
    wire _0136_;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_2256;
    wire new_Jinkela_wire_2680;
    wire _0158_;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_2503;
    wire new_Jinkela_wire_1941;
    wire _0448_;
    wire new_Jinkela_wire_2175;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_2188;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_2263;
    wire _0227_;
    wire _0401_;
    wire new_Jinkela_wire_924;
    wire _0269_;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_1439;
    wire new_Jinkela_wire_1788;
    wire _0122_;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_2139;
    wire new_Jinkela_wire_1865;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_2657;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_1360;
    wire _0171_;
    wire new_Jinkela_wire_1721;
    wire new_net_22;
    wire new_Jinkela_wire_2112;
    wire new_Jinkela_wire_2260;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_2531;
    wire new_Jinkela_wire_1947;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_1774;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_1728;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_2294;
    wire new_Jinkela_wire_2614;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_1540;
    wire new_net_0;
    wire new_Jinkela_wire_2646;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_279;
    wire _0038_;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_2422;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_956;
    wire _0310_;
    wire _0346_;
    wire new_Jinkela_wire_1971;
    wire _0428_;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_1344;
    wire _0430_;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_217;
    wire _0043_;
    wire new_Jinkela_wire_1617;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_2109;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_2606;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_1820;
    wire new_Jinkela_wire_1734;
    wire new_Jinkela_wire_1745;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_2573;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_2467;
    wire new_Jinkela_wire_2492;
    wire _0366_;
    wire _0396_;
    wire new_Jinkela_wire_86;
    wire new_Jinkela_wire_1475;
    wire _0306_;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_2595;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_2204;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_2044;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_2140;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_2283;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_2400;
    wire _0221_;
    wire _0453_;
    wire new_Jinkela_wire_1787;
    wire _0103_;
    wire new_Jinkela_wire_429;
    wire _0335_;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_1785;
    wire new_Jinkela_wire_82;
    wire _0275_;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_2365;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_1643;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_1583;
    wire new_Jinkela_wire_1315;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_2509;
    wire new_Jinkela_wire_2429;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_1773;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_1995;
    wire new_Jinkela_wire_2137;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_1869;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_2189;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_2649;
    wire new_Jinkela_wire_909;
    wire _0324_;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_2447;
    wire new_Jinkela_wire_2466;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_2570;
    wire new_Jinkela_wire_1607;
    wire _0087_;
    wire new_Jinkela_wire_1217;
    wire _0304_;
    wire new_Jinkela_wire_1985;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_52;
    wire _0200_;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_2542;
    wire new_Jinkela_wire_2588;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_2285;
    wire _0046_;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_1169;
    wire _0134_;
    wire new_Jinkela_wire_2169;
    wire new_Jinkela_wire_2554;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_2435;
    wire _0278_;
    wire new_Jinkela_wire_1404;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_2715;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_1557;
    wire _0215_;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_1828;
    wire new_Jinkela_wire_1763;
    wire _0072_;
    wire new_Jinkela_wire_2405;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_738;
    wire _0031_;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_1016;
    wire _0146_;
    wire new_Jinkela_wire_2713;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_2616;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_2386;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_2003;
    wire new_Jinkela_wire_2311;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_2198;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_205;
    wire _0391_;
    wire _0486_;
    wire new_Jinkela_wire_1477;
    wire _0294_;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_1375;
    wire _0464_;
    wire new_Jinkela_wire_1846;
    wire new_Jinkela_wire_2302;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_1911;
    wire new_Jinkela_wire_2153;
    wire _0177_;
    wire new_Jinkela_wire_1881;
    wire new_net_2;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_2220;
    wire new_Jinkela_wire_2722;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_1917;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_255;
    wire new_net_10;
    wire new_Jinkela_wire_2259;
    wire _0341_;
    wire new_Jinkela_wire_2037;
    wire new_Jinkela_wire_2653;
    wire _0057_;
    wire new_Jinkela_wire_1777;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_2425;
    wire _0347_;
    wire new_Jinkela_wire_2232;
    wire _0028_;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_1979;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_743;
    wire _0216_;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_2705;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_2069;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_2341;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_2504;
    wire new_Jinkela_wire_1356;
    wire _0445_;
    wire new_Jinkela_wire_2190;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_2076;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_2555;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_871;
    wire _0222_;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_2321;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_1115;
    wire _0337_;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_2138;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_2013;
    wire new_net_946;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_1759;
    wire new_Jinkela_wire_2518;
    wire new_Jinkela_wire_1296;
    input G131;
    input G26;
    input G16;
    input G30;
    input G57;
    input G12;
    input G73;
    input G147;
    input G107;
    input G75;
    input G103;
    input G141;
    input G24;
    input G62;
    input G27;
    input G76;
    input G123;
    input G4;
    input G142;
    input G118;
    input G133;
    input G150;
    input G145;
    input G39;
    input G94;
    input G19;
    input G5;
    input G152;
    input G23;
    input G96;
    input G110;
    input G120;
    input G112;
    input G47;
    input G82;
    input G157;
    input G91;
    input G106;
    input G56;
    input G13;
    input G60;
    input G148;
    input G64;
    input G20;
    input G52;
    input G8;
    input G98;
    input G11;
    input G32;
    input G66;
    input G14;
    input G143;
    input G146;
    input G28;
    input G83;
    input G108;
    input G42;
    input G3;
    input G63;
    input G144;
    input G84;
    input G87;
    input G104;
    input G132;
    input G80;
    input G36;
    input G10;
    input G54;
    input G59;
    input G92;
    input G72;
    input G79;
    input G117;
    input G31;
    input G113;
    input G116;
    input G44;
    input G1;
    input G65;
    input G154;
    input G124;
    input G55;
    input G137;
    input G38;
    input G105;
    input G61;
    input G119;
    input G90;
    input G33;
    input G22;
    input G35;
    input G115;
    input G134;
    input G40;
    input G2;
    input G25;
    input G58;
    input G111;
    input G100;
    input G126;
    input G70;
    input G9;
    input G149;
    input G121;
    input G48;
    input G78;
    input G136;
    input G43;
    input G7;
    input G81;
    input G140;
    input G89;
    input G77;
    input G95;
    input G34;
    input G99;
    input G68;
    input G67;
    input G86;
    input G15;
    input G122;
    input G45;
    input G129;
    input G18;
    input G6;
    input G93;
    input G101;
    input G125;
    input G69;
    input G114;
    input G139;
    input G97;
    input G51;
    input G109;
    input G17;
    input G74;
    input G156;
    input G153;
    input G50;
    input G138;
    input G135;
    input G71;
    input G85;
    input G155;
    input G53;
    input G37;
    input G130;
    input G46;
    input G41;
    input G49;
    input G127;
    input G102;
    input G128;
    input G151;
    input G21;
    input G88;
    input G29;
    output G2586;
    output G2567;
    output G2566;
    output G2546;
    output G2545;
    output G2549;
    output G2556;
    output G2590;
    output G2579;
    output G2591;
    output G2563;
    output G2569;
    output G2580;
    output G2571;
    output G2550;
    output G2531;
    output G2534;
    output G2570;
    output G2583;
    output G2557;
    output G2593;
    output G2535;
    output G2548;
    output G2532;
    output G2588;
    output G2587;
    output G2574;
    output G2577;
    output G2541;
    output G2543;
    output G2594;
    output G2576;
    output G2565;
    output G2582;
    output G2554;
    output G2558;
    output G2540;
    output G2572;
    output G2536;
    output G2562;
    output G2555;
    output G2552;
    output G2559;
    output G2573;
    output G2542;
    output G2578;
    output G2568;
    output G2539;
    output G2592;
    output G2537;
    output G2560;
    output G2581;
    output G2547;
    output G2544;
    output G2553;
    output G2561;
    output G2589;
    output G2564;
    output G2575;
    output G2585;
    output G2551;
    output G2538;
    output G2584;
    output G2533;

    bfr new_Jinkela_buffer_1605 (
        .din(new_Jinkela_wire_2178),
        .dout(new_Jinkela_wire_2179)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_2162),
        .dout(new_Jinkela_wire_2163)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(_0131_),
        .c(new_Jinkela_wire_2189),
        .b(new_Jinkela_wire_2190)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_2163),
        .dout(new_Jinkela_wire_2164)
    );

    bfr new_Jinkela_buffer_1606 (
        .din(new_Jinkela_wire_2179),
        .dout(new_Jinkela_wire_2180)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_2164),
        .dout(new_Jinkela_wire_2165)
    );

    spl2 new_Jinkela_splitter_219 (
        .a(_0339_),
        .c(new_Jinkela_wire_2187),
        .b(new_Jinkela_wire_2188)
    );

    bfr new_Jinkela_buffer_1596 (
        .din(new_Jinkela_wire_2165),
        .dout(new_Jinkela_wire_2166)
    );

    bfr new_Jinkela_buffer_1607 (
        .din(new_Jinkela_wire_2180),
        .dout(new_Jinkela_wire_2181)
    );

    bfr new_Jinkela_buffer_1597 (
        .din(new_Jinkela_wire_2166),
        .dout(new_Jinkela_wire_2167)
    );

    bfr new_Jinkela_buffer_1610 (
        .din(new_Jinkela_wire_2191),
        .dout(new_Jinkela_wire_2192)
    );

    bfr new_Jinkela_buffer_1598 (
        .din(new_Jinkela_wire_2167),
        .dout(new_Jinkela_wire_2168)
    );

    bfr new_Jinkela_buffer_1608 (
        .din(new_Jinkela_wire_2181),
        .dout(new_Jinkela_wire_2182)
    );

    bfr new_Jinkela_buffer_1599 (
        .din(new_Jinkela_wire_2168),
        .dout(new_Jinkela_wire_2169)
    );

    bfr new_Jinkela_buffer_1609 (
        .din(_0025_),
        .dout(new_Jinkela_wire_2191)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(new_Jinkela_wire_2169),
        .c(new_Jinkela_wire_2170),
        .b(new_Jinkela_wire_2171)
    );

    bfr new_Jinkela_buffer_1636 (
        .din(_0060_),
        .dout(new_Jinkela_wire_2218)
    );

    bfr new_Jinkela_buffer_1611 (
        .din(new_net_967),
        .dout(new_Jinkela_wire_2193)
    );

    bfr new_Jinkela_buffer_1612 (
        .din(new_Jinkela_wire_2193),
        .dout(new_Jinkela_wire_2194)
    );

    bfr new_Jinkela_buffer_1638 (
        .din(_0331_),
        .dout(new_Jinkela_wire_2220)
    );

    bfr new_Jinkela_buffer_1613 (
        .din(new_Jinkela_wire_2194),
        .dout(new_Jinkela_wire_2195)
    );

    bfr new_Jinkela_buffer_1637 (
        .din(new_Jinkela_wire_2218),
        .dout(new_Jinkela_wire_2219)
    );

    bfr new_Jinkela_buffer_1614 (
        .din(new_Jinkela_wire_2195),
        .dout(new_Jinkela_wire_2196)
    );

    bfr new_Jinkela_buffer_1644 (
        .din(new_net_952),
        .dout(new_Jinkela_wire_2226)
    );

    bfr new_Jinkela_buffer_1615 (
        .din(new_Jinkela_wire_2196),
        .dout(new_Jinkela_wire_2197)
    );

    bfr new_Jinkela_buffer_1639 (
        .din(new_Jinkela_wire_2220),
        .dout(new_Jinkela_wire_2221)
    );

    bfr new_Jinkela_buffer_1616 (
        .din(new_Jinkela_wire_2197),
        .dout(new_Jinkela_wire_2198)
    );

    bfr new_Jinkela_buffer_1670 (
        .din(_0468_),
        .dout(new_Jinkela_wire_2252)
    );

    bfr new_Jinkela_buffer_1617 (
        .din(new_Jinkela_wire_2198),
        .dout(new_Jinkela_wire_2199)
    );

    bfr new_Jinkela_buffer_1640 (
        .din(new_Jinkela_wire_2221),
        .dout(new_Jinkela_wire_2222)
    );

    bfr new_Jinkela_buffer_1618 (
        .din(new_Jinkela_wire_2199),
        .dout(new_Jinkela_wire_2200)
    );

    bfr new_Jinkela_buffer_1645 (
        .din(new_Jinkela_wire_2226),
        .dout(new_Jinkela_wire_2227)
    );

    bfr new_Jinkela_buffer_1619 (
        .din(new_Jinkela_wire_2200),
        .dout(new_Jinkela_wire_2201)
    );

    bfr new_Jinkela_buffer_1641 (
        .din(new_Jinkela_wire_2222),
        .dout(new_Jinkela_wire_2223)
    );

    bfr new_Jinkela_buffer_1620 (
        .din(new_Jinkela_wire_2201),
        .dout(new_Jinkela_wire_2202)
    );

    bfr new_Jinkela_buffer_2025 (
        .din(new_Jinkela_wire_2741),
        .dout(new_Jinkela_wire_2742)
    );

    bfr new_Jinkela_buffer_1673 (
        .din(_0156_),
        .dout(new_Jinkela_wire_2255)
    );

    bfr new_Jinkela_buffer_1676 (
        .din(_0378_),
        .dout(new_Jinkela_wire_2260)
    );

    bfr new_Jinkela_buffer_1621 (
        .din(new_Jinkela_wire_2202),
        .dout(new_Jinkela_wire_2203)
    );

    bfr new_Jinkela_buffer_1642 (
        .din(new_Jinkela_wire_2223),
        .dout(new_Jinkela_wire_2224)
    );

    bfr new_Jinkela_buffer_1622 (
        .din(new_Jinkela_wire_2203),
        .dout(new_Jinkela_wire_2204)
    );

    bfr new_Jinkela_buffer_1646 (
        .din(new_Jinkela_wire_2227),
        .dout(new_Jinkela_wire_2228)
    );

    bfr new_Jinkela_buffer_1623 (
        .din(new_Jinkela_wire_2204),
        .dout(new_Jinkela_wire_2205)
    );

    bfr new_Jinkela_buffer_1643 (
        .din(new_Jinkela_wire_2224),
        .dout(new_Jinkela_wire_2225)
    );

    and_bi _1032_ (
        .a(new_Jinkela_wire_1040),
        .b(new_Jinkela_wire_2451),
        .c(_0498_)
    );

    or_bb _1033_ (
        .a(new_Jinkela_wire_2447),
        .b(_0497_),
        .c(new_net_959)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_705),
        .dout(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    bfr new_Jinkela_buffer_1814 (
        .din(new_Jinkela_wire_2427),
        .dout(new_Jinkela_wire_2428)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(new_Jinkela_wire_1482),
        .dout(new_Jinkela_wire_1483)
    );

    spl4L new_Jinkela_splitter_130 (
        .a(new_Jinkela_wire_1503),
        .c(new_Jinkela_wire_1504),
        .e(new_Jinkela_wire_1505),
        .b(new_Jinkela_wire_1506),
        .d(new_Jinkela_wire_1507)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    spl4L new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_1498),
        .c(new_Jinkela_wire_1499),
        .e(new_Jinkela_wire_1500),
        .b(new_Jinkela_wire_1501),
        .d(new_Jinkela_wire_1502)
    );

    bfr new_Jinkela_buffer_1815 (
        .din(new_Jinkela_wire_2428),
        .dout(new_Jinkela_wire_2429)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_1483),
        .dout(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_1833 (
        .din(new_Jinkela_wire_2446),
        .dout(new_Jinkela_wire_2447)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(_0111_),
        .c(new_Jinkela_wire_1568),
        .b(new_Jinkela_wire_1569)
    );

    bfr new_Jinkela_buffer_1816 (
        .din(new_Jinkela_wire_2429),
        .dout(new_Jinkela_wire_2430)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_1484),
        .dout(new_Jinkela_wire_1485)
    );

    bfr new_Jinkela_buffer_1856 (
        .din(_0330_),
        .dout(new_Jinkela_wire_2490)
    );

    spl2 new_Jinkela_splitter_236 (
        .a(new_Jinkela_wire_2453),
        .c(new_Jinkela_wire_2454),
        .b(new_Jinkela_wire_2455)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_762),
        .dout(new_Jinkela_wire_763)
    );

    bfr new_Jinkela_buffer_1817 (
        .din(new_Jinkela_wire_2430),
        .dout(new_Jinkela_wire_2431)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_1485),
        .dout(new_Jinkela_wire_1486)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_1857 (
        .din(_0476_),
        .dout(new_Jinkela_wire_2493)
    );

    spl2 new_Jinkela_splitter_238 (
        .a(new_Jinkela_wire_2456),
        .c(new_Jinkela_wire_2457),
        .b(new_Jinkela_wire_2458)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_1818 (
        .din(new_Jinkela_wire_2431),
        .dout(new_Jinkela_wire_2432)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_764),
        .dout(new_Jinkela_wire_765)
    );

    spl3L new_Jinkela_splitter_134 (
        .a(new_net_9),
        .c(new_Jinkela_wire_1519),
        .b(new_Jinkela_wire_1520),
        .d(new_Jinkela_wire_1521)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(new_Jinkela_wire_1487),
        .dout(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    spl3L new_Jinkela_splitter_135 (
        .a(new_Jinkela_wire_1521),
        .c(new_Jinkela_wire_1522),
        .b(new_Jinkela_wire_1523),
        .d(new_Jinkela_wire_1524)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    spl4L new_Jinkela_splitter_239 (
        .a(new_Jinkela_wire_2459),
        .c(new_Jinkela_wire_2460),
        .e(new_Jinkela_wire_2461),
        .b(new_Jinkela_wire_2462),
        .d(new_Jinkela_wire_2463)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_1549),
        .dout(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_1488),
        .dout(new_Jinkela_wire_1489)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    spl2 new_Jinkela_splitter_243 (
        .a(_0088_),
        .c(new_Jinkela_wire_2491),
        .b(new_Jinkela_wire_2492)
    );

    bfr new_Jinkela_buffer_1854 (
        .din(new_Jinkela_wire_2485),
        .dout(new_Jinkela_wire_2486)
    );

    spl3L new_Jinkela_splitter_247 (
        .a(_0007_),
        .c(new_Jinkela_wire_2501),
        .b(new_Jinkela_wire_2503),
        .d(new_Jinkela_wire_2508)
    );

    bfr new_Jinkela_buffer_591 (
        .din(G119),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_1858 (
        .din(_0470_),
        .dout(new_Jinkela_wire_2496)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_1855 (
        .din(new_Jinkela_wire_2486),
        .dout(new_Jinkela_wire_2487)
    );

    bfr new_Jinkela_buffer_1838 (
        .din(new_Jinkela_wire_2464),
        .dout(new_Jinkela_wire_2465)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(_0293_),
        .c(new_Jinkela_wire_1547),
        .b(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_1839 (
        .din(new_Jinkela_wire_2465),
        .dout(new_Jinkela_wire_2466)
    );

    bfr new_Jinkela_buffer_594 (
        .din(G90),
        .dout(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_765),
        .dout(new_Jinkela_wire_766)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(new_Jinkela_wire_1491),
        .dout(new_Jinkela_wire_1492)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_1840 (
        .din(new_Jinkela_wire_2466),
        .dout(new_Jinkela_wire_2467)
    );

    bfr new_Jinkela_buffer_1837 (
        .din(new_Jinkela_wire_2463),
        .dout(new_Jinkela_wire_2464)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    spl2 new_Jinkela_splitter_242 (
        .a(new_Jinkela_wire_2487),
        .c(new_Jinkela_wire_2488),
        .b(new_Jinkela_wire_2489)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_1492),
        .dout(new_Jinkela_wire_1493)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    bfr new_Jinkela_buffer_1841 (
        .din(new_Jinkela_wire_2467),
        .dout(new_Jinkela_wire_2468)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_net_963),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_737),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_1493),
        .dout(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(_0173_),
        .c(new_Jinkela_wire_2499),
        .b(new_Jinkela_wire_2500)
    );

    bfr new_Jinkela_buffer_1842 (
        .din(new_Jinkela_wire_2468),
        .dout(new_Jinkela_wire_2469)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(_0454_),
        .c(new_Jinkela_wire_1566),
        .b(new_Jinkela_wire_1567)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(_0257_),
        .c(new_Jinkela_wire_2494),
        .b(new_Jinkela_wire_2495)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_1494),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_716),
        .dout(new_Jinkela_wire_717)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(new_Jinkela_wire_2496),
        .c(new_Jinkela_wire_2497),
        .b(new_Jinkela_wire_2498)
    );

    bfr new_Jinkela_buffer_1843 (
        .din(new_Jinkela_wire_2469),
        .dout(new_Jinkela_wire_2470)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    spl2 new_Jinkela_splitter_131 (
        .a(new_Jinkela_wire_1511),
        .c(new_Jinkela_wire_1512),
        .b(new_Jinkela_wire_1513)
    );

    spl4L new_Jinkela_splitter_249 (
        .a(new_Jinkela_wire_2508),
        .c(new_Jinkela_wire_2509),
        .e(new_Jinkela_wire_2510),
        .b(new_Jinkela_wire_2511),
        .d(new_Jinkela_wire_2512)
    );

    spl2 new_Jinkela_splitter_127 (
        .a(new_Jinkela_wire_1495),
        .c(new_Jinkela_wire_1496),
        .b(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_1844 (
        .din(new_Jinkela_wire_2470),
        .dout(new_Jinkela_wire_2471)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(_0251_),
        .c(new_Jinkela_wire_2513),
        .b(new_Jinkela_wire_2514)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_1524),
        .dout(new_Jinkela_wire_1525)
    );

    bfr new_Jinkela_buffer_1845 (
        .din(new_Jinkela_wire_2471),
        .dout(new_Jinkela_wire_2472)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_1859 (
        .din(new_Jinkela_wire_2501),
        .dout(new_Jinkela_wire_2502)
    );

    bfr new_Jinkela_buffer_1846 (
        .din(new_Jinkela_wire_2472),
        .dout(new_Jinkela_wire_2473)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_739),
        .dout(new_Jinkela_wire_740)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    bfr new_Jinkela_buffer_1860 (
        .din(new_net_17),
        .dout(new_Jinkela_wire_2515)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_1847 (
        .din(new_Jinkela_wire_2473),
        .dout(new_Jinkela_wire_2474)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_1527),
        .dout(new_Jinkela_wire_1528)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(new_Jinkela_wire_721),
        .c(new_Jinkela_wire_722),
        .b(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_1551),
        .dout(new_Jinkela_wire_1552)
    );

    bfr new_Jinkela_buffer_1848 (
        .din(new_Jinkela_wire_2474),
        .dout(new_Jinkela_wire_2475)
    );

    bfr new_Jinkela_buffer_598 (
        .din(G33),
        .dout(new_Jinkela_wire_783)
    );

    spl3L new_Jinkela_splitter_136 (
        .a(new_Jinkela_wire_1528),
        .c(new_Jinkela_wire_1529),
        .b(new_Jinkela_wire_1530),
        .d(new_Jinkela_wire_1531)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(_0287_),
        .dout(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_1849 (
        .din(new_Jinkela_wire_2475),
        .dout(new_Jinkela_wire_2476)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    spl3L new_Jinkela_splitter_137 (
        .a(new_Jinkela_wire_1531),
        .c(new_Jinkela_wire_1532),
        .b(new_Jinkela_wire_1533),
        .d(new_Jinkela_wire_1534)
    );

    spl4L new_Jinkela_splitter_248 (
        .a(new_Jinkela_wire_2503),
        .c(new_Jinkela_wire_2504),
        .e(new_Jinkela_wire_2505),
        .b(new_Jinkela_wire_2506),
        .d(new_Jinkela_wire_2507)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_770),
        .dout(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(new_Jinkela_wire_1552),
        .dout(new_Jinkela_wire_1553)
    );

    bfr new_Jinkela_buffer_1850 (
        .din(new_Jinkela_wire_2476),
        .dout(new_Jinkela_wire_2477)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_1883 (
        .din(_0473_),
        .dout(new_Jinkela_wire_2540)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(_0422_),
        .dout(new_Jinkela_wire_1579)
    );

    bfr new_Jinkela_buffer_1851 (
        .din(new_Jinkela_wire_2477),
        .dout(new_Jinkela_wire_2478)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1088),
        .dout(new_Jinkela_wire_1089)
    );

    and_bi _0864_ (
        .a(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_22),
        .c(_0337_)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_872 (
        .din(G97),
        .dout(new_Jinkela_wire_1127)
    );

    and_bi _0865_ (
        .a(new_Jinkela_wire_65),
        .b(new_Jinkela_wire_2060),
        .c(_0338_)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1089),
        .dout(new_Jinkela_wire_1090)
    );

    and_bi _0866_ (
        .a(new_Jinkela_wire_2724),
        .b(_0338_),
        .c(_0339_)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(G117),
        .c(new_Jinkela_wire_616),
        .b(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_473 (
        .din(G113),
        .dout(new_Jinkela_wire_649)
    );

    or_bb _0867_ (
        .a(new_Jinkela_wire_2187),
        .b(new_Jinkela_wire_16),
        .c(_0340_)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1090),
        .dout(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    and_bi _0868_ (
        .a(new_Jinkela_wire_15),
        .b(new_Jinkela_wire_2188),
        .c(_0341_)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    bfr new_Jinkela_buffer_470 (
        .din(G31),
        .dout(new_Jinkela_wire_646)
    );

    and_bi _0869_ (
        .a(_0340_),
        .b(_0341_),
        .c(_0342_)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1091),
        .dout(new_Jinkela_wire_1092)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    and_bi _0870_ (
        .a(new_Jinkela_wire_252),
        .b(new_Jinkela_wire_425),
        .c(_0343_)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    and_bi _0871_ (
        .a(new_Jinkela_wire_273),
        .b(new_Jinkela_wire_1969),
        .c(_0344_)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    and_bi _0872_ (
        .a(new_Jinkela_wire_2093),
        .b(_0344_),
        .c(_0345_)
    );

    or_bb _0873_ (
        .a(new_Jinkela_wire_1853),
        .b(new_Jinkela_wire_1169),
        .c(_0346_)
    );

    spl4L new_Jinkela_splitter_54 (
        .a(new_Jinkela_wire_625),
        .c(new_Jinkela_wire_626),
        .e(new_Jinkela_wire_631),
        .b(new_Jinkela_wire_636),
        .d(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_1093),
        .dout(new_Jinkela_wire_1094)
    );

    and_bi _0874_ (
        .a(new_Jinkela_wire_1170),
        .b(new_Jinkela_wire_1854),
        .c(_0347_)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_876 (
        .din(G51),
        .dout(new_Jinkela_wire_1131)
    );

    and_bi _0875_ (
        .a(_0346_),
        .b(_0347_),
        .c(_0348_)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    or_bb _0876_ (
        .a(new_Jinkela_wire_1599),
        .b(_0342_),
        .c(_0349_)
    );

    bfr new_Jinkela_buffer_477 (
        .din(G116),
        .dout(new_Jinkela_wire_653)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(new_Jinkela_wire_616),
        .c(new_Jinkela_wire_617),
        .b(new_Jinkela_wire_620)
    );

    or_bb _0877_ (
        .a(_0349_),
        .b(new_Jinkela_wire_1894),
        .c(_0350_)
    );

    spl4L new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_620),
        .c(new_Jinkela_wire_621),
        .e(new_Jinkela_wire_622),
        .b(new_Jinkela_wire_623),
        .d(new_Jinkela_wire_624)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1095),
        .dout(new_Jinkela_wire_1096)
    );

    and_bi _0878_ (
        .a(new_Jinkela_wire_259),
        .b(new_Jinkela_wire_848),
        .c(_0351_)
    );

    spl2 new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_617),
        .c(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_619)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_1128),
        .dout(new_Jinkela_wire_1129)
    );

    and_bi _0879_ (
        .a(new_Jinkela_wire_269),
        .b(new_Jinkela_wire_1517),
        .c(_0352_)
    );

    spl4L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_626),
        .c(new_Jinkela_wire_627),
        .e(new_Jinkela_wire_628),
        .b(new_Jinkela_wire_629),
        .d(new_Jinkela_wire_630)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    and_bi _0880_ (
        .a(new_Jinkela_wire_1929),
        .b(_0352_),
        .c(_0353_)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_1127),
        .dout(new_Jinkela_wire_1128)
    );

    and_bi _0881_ (
        .a(new_Jinkela_wire_1123),
        .b(new_Jinkela_wire_1444),
        .c(_0354_)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    spl4L new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_631),
        .c(new_Jinkela_wire_632),
        .e(new_Jinkela_wire_633),
        .b(new_Jinkela_wire_634),
        .d(new_Jinkela_wire_635)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1097),
        .dout(new_Jinkela_wire_1098)
    );

    and_bi _0882_ (
        .a(new_Jinkela_wire_1247),
        .b(new_Jinkela_wire_1548),
        .c(_0355_)
    );

    or_bb _0883_ (
        .a(_0355_),
        .b(new_Jinkela_wire_1343),
        .c(_0356_)
    );

    bfr new_Jinkela_buffer_484 (
        .din(G65),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_882 (
        .din(G109),
        .dout(new_Jinkela_wire_1137)
    );

    spl4L new_Jinkela_splitter_57 (
        .a(new_Jinkela_wire_636),
        .c(new_Jinkela_wire_637),
        .e(new_Jinkela_wire_638),
        .b(new_Jinkela_wire_639),
        .d(new_Jinkela_wire_640)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_1098),
        .c(new_Jinkela_wire_1099),
        .b(new_Jinkela_wire_1100)
    );

    and_bi _0884_ (
        .a(new_Jinkela_wire_880),
        .b(new_Jinkela_wire_1477),
        .c(_0357_)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_641),
        .c(new_Jinkela_wire_642),
        .e(new_Jinkela_wire_643),
        .b(new_Jinkela_wire_644),
        .d(new_Jinkela_wire_645)
    );

    spl2 new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_1100),
        .c(new_Jinkela_wire_1101),
        .b(new_Jinkela_wire_1102)
    );

    and_bi _0885_ (
        .a(new_Jinkela_wire_39),
        .b(new_Jinkela_wire_1074),
        .c(_0358_)
    );

    and_bi _0886_ (
        .a(new_Jinkela_wire_63),
        .b(new_Jinkela_wire_2273),
        .c(_0359_)
    );

    bfr new_Jinkela_buffer_478 (
        .din(G44),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    and_bi _0887_ (
        .a(new_Jinkela_wire_1786),
        .b(_0359_),
        .c(_0360_)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1131),
        .dout(new_Jinkela_wire_1132)
    );

    and_bi _0888_ (
        .a(new_Jinkela_wire_841),
        .b(new_Jinkela_wire_2183),
        .c(_0361_)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    or_bb _0889_ (
        .a(_0361_),
        .b(_0357_),
        .c(_0362_)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    or_bb _0890_ (
        .a(_0362_),
        .b(_0356_),
        .c(_0363_)
    );

    bfr new_Jinkela_buffer_487 (
        .din(1'b0),
        .dout(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1116),
        .dout(new_Jinkela_wire_1117)
    );

    and_bi _0891_ (
        .a(new_Jinkela_wire_48),
        .b(new_Jinkela_wire_1076),
        .c(_0364_)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_Jinkela_wire_1129),
        .dout(new_Jinkela_wire_1130)
    );

    and_bi _0892_ (
        .a(new_Jinkela_wire_61),
        .b(new_Jinkela_wire_2360),
        .c(_0365_)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_660),
        .dout(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    and_bi _0893_ (
        .a(new_Jinkela_wire_2440),
        .b(_0365_),
        .c(_0366_)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    bfr new_Jinkela_buffer_886 (
        .din(G17),
        .dout(new_Jinkela_wire_1141)
    );

    and_bi _0894_ (
        .a(new_Jinkela_wire_225),
        .b(new_Jinkela_wire_2601),
        .c(_0367_)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(G154),
        .c(new_Jinkela_wire_692),
        .b(new_Jinkela_wire_693)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    bfr new_Jinkela_buffer_516 (
        .din(G124),
        .dout(new_Jinkela_wire_694)
    );

    and_bi _0895_ (
        .a(new_Jinkela_wire_274),
        .b(new_Jinkela_wire_1654),
        .c(_0368_)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1132),
        .dout(new_Jinkela_wire_1133)
    );

    and_bi _0896_ (
        .a(new_Jinkela_wire_253),
        .b(new_Jinkela_wire_787),
        .c(_0369_)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    or_bb _0897_ (
        .a(_0369_),
        .b(new_Jinkela_wire_886),
        .c(_0370_)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1137),
        .dout(new_Jinkela_wire_1138)
    );

    or_bb _0898_ (
        .a(new_Jinkela_wire_2182),
        .b(_0368_),
        .c(_0371_)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    or_bb _0899_ (
        .a(new_Jinkela_wire_2450),
        .b(_0367_),
        .c(_0372_)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1133),
        .dout(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_550 (
        .din(G137),
        .dout(new_Jinkela_wire_730)
    );

    bfr new_Jinkela_buffer_1888 (
        .din(_0312_),
        .dout(new_Jinkela_wire_2549)
    );

    and_bi _0900_ (
        .a(new_Jinkela_wire_192),
        .b(new_Jinkela_wire_1366),
        .c(_0373_)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_664),
        .dout(new_Jinkela_wire_665)
    );

    spl3L new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_1121),
        .c(new_Jinkela_wire_1122),
        .b(new_Jinkela_wire_1123),
        .d(new_Jinkela_wire_1124)
    );

    and_bi _0901_ (
        .a(new_Jinkela_wire_226),
        .b(new_Jinkela_wire_2602),
        .c(_0374_)
    );

    bfr new_Jinkela_buffer_888 (
        .din(G74),
        .dout(new_Jinkela_wire_1143)
    );

    or_bb _0902_ (
        .a(_0374_),
        .b(new_Jinkela_wire_1991),
        .c(_0375_)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_665),
        .dout(new_Jinkela_wire_666)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    or_bb _0903_ (
        .a(_0375_),
        .b(_0372_),
        .c(_0376_)
    );

    bfr new_Jinkela_buffer_544 (
        .din(G55),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1134),
        .dout(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_694),
        .dout(new_Jinkela_wire_695)
    );

    or_bb _0904_ (
        .a(new_Jinkela_wire_2386),
        .b(_0363_),
        .c(_0377_)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_666),
        .dout(new_Jinkela_wire_667)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    and_bi _0905_ (
        .a(new_Jinkela_wire_102),
        .b(new_Jinkela_wire_2611),
        .c(_0378_)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1138),
        .dout(new_Jinkela_wire_1139)
    );

    and_bi _0696_ (
        .a(new_Jinkela_wire_858),
        .b(new_Jinkela_wire_2507),
        .c(_0184_)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_216),
        .dout(new_Jinkela_wire_217)
    );

    bfr new_Jinkela_buffer_2026 (
        .din(new_Jinkela_wire_2742),
        .dout(new_Jinkela_wire_2743)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_208),
        .dout(new_Jinkela_wire_209)
    );

    and_bi _0697_ (
        .a(new_Jinkela_wire_347),
        .b(new_Jinkela_wire_1849),
        .c(_0185_)
    );

    bfr new_Jinkela_buffer_172 (
        .din(G19),
        .dout(new_Jinkela_wire_243)
    );

    or_bb _0698_ (
        .a(_0185_),
        .b(_0184_),
        .c(_0186_)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_209),
        .dout(new_Jinkela_wire_210)
    );

    and_bi _0699_ (
        .a(_0183_),
        .b(_0186_),
        .c(_0187_)
    );

    and_bi _0700_ (
        .a(new_Jinkela_wire_1412),
        .b(new_Jinkela_wire_1516),
        .c(_0188_)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    and_bi _0701_ (
        .a(new_Jinkela_wire_1413),
        .b(new_Jinkela_wire_1518),
        .c(_0189_)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_237),
        .dout(new_Jinkela_wire_238)
    );

    and_bi _0702_ (
        .a(_0188_),
        .b(_0189_),
        .c(_0190_)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    and_bi _0703_ (
        .a(new_Jinkela_wire_2499),
        .b(new_Jinkela_wire_1700),
        .c(_0191_)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    and_bi _0704_ (
        .a(new_Jinkela_wire_2500),
        .b(new_Jinkela_wire_1701),
        .c(_0192_)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    and_bi _0705_ (
        .a(_0191_),
        .b(_0192_),
        .c(_0193_)
    );

    bfr new_Jinkela_buffer_174 (
        .din(G5),
        .dout(new_Jinkela_wire_245)
    );

    and_bi _0706_ (
        .a(new_Jinkela_wire_84),
        .b(new_Jinkela_wire_1983),
        .c(_0194_)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    and_bi _0707_ (
        .a(new_Jinkela_wire_1196),
        .b(new_Jinkela_wire_1842),
        .c(_0195_)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_240),
        .dout(new_Jinkela_wire_241)
    );

    and_bi _0708_ (
        .a(_0194_),
        .b(_0195_),
        .c(_0196_)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_221),
        .dout(new_Jinkela_wire_222)
    );

    and_bi _0709_ (
        .a(new_Jinkela_wire_984),
        .b(new_Jinkela_wire_1933),
        .c(_0197_)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    and_bi _0710_ (
        .a(new_Jinkela_wire_767),
        .b(new_Jinkela_wire_2504),
        .c(_0198_)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_222),
        .dout(new_Jinkela_wire_223)
    );

    or_bb _0711_ (
        .a(_0198_),
        .b(_0197_),
        .c(_0199_)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_241),
        .dout(new_Jinkela_wire_242)
    );

    and_bi _0712_ (
        .a(_0196_),
        .b(_0199_),
        .c(_0200_)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    and_bi _0713_ (
        .a(new_Jinkela_wire_2649),
        .b(new_Jinkela_wire_2619),
        .c(_0201_)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(G152),
        .c(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_248)
    );

    spl3L new_Jinkela_splitter_24 (
        .a(G23),
        .c(new_Jinkela_wire_249),
        .b(new_Jinkela_wire_251),
        .d(new_Jinkela_wire_256)
    );

    and_bi _0714_ (
        .a(new_Jinkela_wire_2648),
        .b(new_Jinkela_wire_2617),
        .c(_0202_)
    );

    spl3L new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_224),
        .c(new_Jinkela_wire_225),
        .b(new_Jinkela_wire_226),
        .d(new_Jinkela_wire_227)
    );

    and_bi _0715_ (
        .a(_0201_),
        .b(_0202_),
        .c(_0203_)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_245),
        .dout(new_Jinkela_wire_246)
    );

    and_bi _0716_ (
        .a(new_Jinkela_wire_1702),
        .b(new_Jinkela_wire_1945),
        .c(_0204_)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    and_bi _0717_ (
        .a(new_Jinkela_wire_1703),
        .b(new_Jinkela_wire_1946),
        .c(_0205_)
    );

    or_bb _0718_ (
        .a(_0205_),
        .b(_0204_),
        .c(_0206_)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    and_ii _0719_ (
        .a(new_Jinkela_wire_1858),
        .b(new_Jinkela_wire_2258),
        .c(_0207_)
    );

    and_bb _0720_ (
        .a(new_Jinkela_wire_1859),
        .b(new_Jinkela_wire_2259),
        .c(_0208_)
    );

    spl2 new_Jinkela_splitter_31 (
        .a(G96),
        .c(new_Jinkela_wire_276),
        .b(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_213 (
        .din(G120),
        .dout(new_Jinkela_wire_310)
    );

    or_bb _0721_ (
        .a(_0208_),
        .b(new_Jinkela_wire_1321),
        .c(_0209_)
    );

    spl4L new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_251),
        .c(new_Jinkela_wire_252),
        .e(new_Jinkela_wire_253),
        .b(new_Jinkela_wire_254),
        .d(new_Jinkela_wire_255)
    );

    and_bi _0722_ (
        .a(new_Jinkela_wire_1964),
        .b(_0209_),
        .c(new_net_15)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    and_bi _0723_ (
        .a(new_Jinkela_wire_2272),
        .b(new_Jinkela_wire_2363),
        .c(_0210_)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    and_bi _0724_ (
        .a(new_Jinkela_wire_2269),
        .b(new_Jinkela_wire_2362),
        .c(_0211_)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_278),
        .dout(new_Jinkela_wire_279)
    );

    and_bi _0725_ (
        .a(_0210_),
        .b(_0211_),
        .c(_0212_)
    );

    bfr new_Jinkela_buffer_209 (
        .din(G110),
        .dout(new_Jinkela_wire_306)
    );

    and_bi _0726_ (
        .a(new_Jinkela_wire_2062),
        .b(new_Jinkela_wire_1819),
        .c(_0213_)
    );

    and_bi _0727_ (
        .a(new_Jinkela_wire_1818),
        .b(new_Jinkela_wire_2063),
        .c(_0214_)
    );

    and_bi _0728_ (
        .a(_0213_),
        .b(_0214_),
        .c(_0215_)
    );

    bfr new_Jinkela_buffer_215 (
        .din(G112),
        .dout(new_Jinkela_wire_328)
    );

    spl4L new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_256),
        .c(new_Jinkela_wire_257),
        .e(new_Jinkela_wire_258),
        .b(new_Jinkela_wire_259),
        .d(new_Jinkela_wire_260)
    );

    and_bi _0729_ (
        .a(new_Jinkela_wire_1603),
        .b(new_Jinkela_wire_2634),
        .c(_0216_)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    and_bi _0730_ (
        .a(new_Jinkela_wire_1604),
        .b(new_Jinkela_wire_2635),
        .c(_0217_)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_net_19),
        .dout(new_Jinkela_wire_1481)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_279),
        .dout(new_Jinkela_wire_280)
    );

    and_bi _0731_ (
        .a(_0216_),
        .b(_0217_),
        .c(_0218_)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    and_bi _0732_ (
        .a(new_Jinkela_wire_627),
        .b(new_Jinkela_wire_1259),
        .c(_0219_)
    );

    spl2 new_Jinkela_splitter_132 (
        .a(_0299_),
        .c(new_Jinkela_wire_1514),
        .b(new_Jinkela_wire_1515)
    );

    bfr new_Jinkela_buffer_219 (
        .din(G47),
        .dout(new_Jinkela_wire_332)
    );

    and_bi _0733_ (
        .a(new_Jinkela_wire_639),
        .b(new_Jinkela_wire_71),
        .c(_0220_)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_307),
        .dout(new_Jinkela_wire_308)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_263),
        .dout(new_Jinkela_wire_264)
    );

    or_bb _0734_ (
        .a(_0220_),
        .b(new_Jinkela_wire_322),
        .c(_0221_)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_280),
        .dout(new_Jinkela_wire_281)
    );

    and_bi _0735_ (
        .a(new_Jinkela_wire_2308),
        .b(_0221_),
        .c(_0222_)
    );

    spl2 new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_264),
        .c(new_Jinkela_wire_265),
        .b(new_Jinkela_wire_268)
    );

    and_bi _0736_ (
        .a(new_Jinkela_wire_1136),
        .b(new_Jinkela_wire_1661),
        .c(_0223_)
    );

    spl4L new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_268),
        .c(new_Jinkela_wire_269),
        .e(new_Jinkela_wire_270),
        .b(new_Jinkela_wire_271),
        .d(new_Jinkela_wire_272)
    );

    and_bi _0737_ (
        .a(new_Jinkela_wire_115),
        .b(new_Jinkela_wire_2706),
        .c(_0224_)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_1925),
        .dout(new_Jinkela_wire_1926)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_1906),
        .dout(new_Jinkela_wire_1907)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_1553),
        .dout(new_Jinkela_wire_1554)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_1917),
        .dout(new_Jinkela_wire_1918)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_1536),
        .dout(new_Jinkela_wire_1537)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_1907),
        .dout(new_Jinkela_wire_1908)
    );

    spl2 new_Jinkela_splitter_141 (
        .a(_0405_),
        .c(new_Jinkela_wire_1582),
        .b(new_Jinkela_wire_1583)
    );

    spl2 new_Jinkela_splitter_142 (
        .a(_0102_),
        .c(new_Jinkela_wire_1584),
        .b(new_Jinkela_wire_1585)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_1537),
        .dout(new_Jinkela_wire_1538)
    );

    spl2 new_Jinkela_splitter_197 (
        .a(_0125_),
        .c(new_Jinkela_wire_1962),
        .b(new_Jinkela_wire_1963)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_1908),
        .dout(new_Jinkela_wire_1909)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(new_Jinkela_wire_1554),
        .dout(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(new_Jinkela_wire_1918),
        .dout(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_1538),
        .dout(new_Jinkela_wire_1539)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_1909),
        .dout(new_Jinkela_wire_1910)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_1571),
        .dout(new_Jinkela_wire_1572)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(new_Jinkela_wire_1539),
        .dout(new_Jinkela_wire_1540)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_1926),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_1910),
        .dout(new_Jinkela_wire_1911)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_1555),
        .dout(new_Jinkela_wire_1556)
    );

    spl2 new_Jinkela_splitter_190 (
        .a(new_Jinkela_wire_1919),
        .c(new_Jinkela_wire_1920),
        .b(new_Jinkela_wire_1921)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(new_Jinkela_wire_1540),
        .dout(new_Jinkela_wire_1541)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_1541),
        .dout(new_Jinkela_wire_1542)
    );

    spl4L new_Jinkela_splitter_194 (
        .a(new_Jinkela_wire_1937),
        .c(new_Jinkela_wire_1938),
        .e(new_Jinkela_wire_1939),
        .b(new_Jinkela_wire_1940),
        .d(new_Jinkela_wire_1941)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(new_Jinkela_wire_1556),
        .dout(new_Jinkela_wire_1557)
    );

    spl4L new_Jinkela_splitter_193 (
        .a(new_Jinkela_wire_1932),
        .c(new_Jinkela_wire_1933),
        .e(new_Jinkela_wire_1934),
        .b(new_Jinkela_wire_1935),
        .d(new_Jinkela_wire_1936)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(new_Jinkela_wire_1542),
        .dout(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(new_Jinkela_wire_1928),
        .dout(new_Jinkela_wire_1929)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(new_Jinkela_wire_1572),
        .dout(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(new_Jinkela_wire_1930),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_1543),
        .dout(new_Jinkela_wire_1544)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_1557),
        .dout(new_Jinkela_wire_1558)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(_0035_),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(new_Jinkela_wire_1942),
        .dout(new_Jinkela_wire_1943)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(new_Jinkela_wire_1544),
        .dout(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(new_Jinkela_wire_1943),
        .dout(new_Jinkela_wire_1944)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_1586),
        .dout(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_1545),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(_0398_),
        .dout(new_Jinkela_wire_1950)
    );

    spl2 new_Jinkela_splitter_195 (
        .a(new_Jinkela_wire_1944),
        .c(new_Jinkela_wire_1945),
        .b(new_Jinkela_wire_1946)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_1558),
        .dout(new_Jinkela_wire_1559)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_1573),
        .dout(new_Jinkela_wire_1574)
    );

    spl2 new_Jinkela_splitter_200 (
        .a(_0483_),
        .c(new_Jinkela_wire_1972),
        .b(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(_0207_),
        .dout(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_1559),
        .dout(new_Jinkela_wire_1560)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_1950),
        .dout(new_Jinkela_wire_1951)
    );

    spl3L new_Jinkela_splitter_201 (
        .a(_0000_),
        .c(new_Jinkela_wire_1974),
        .b(new_Jinkela_wire_1976),
        .d(new_Jinkela_wire_1981)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(new_Jinkela_wire_1951),
        .dout(new_Jinkela_wire_1952)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_1560),
        .dout(new_Jinkela_wire_1561)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_1574),
        .dout(new_Jinkela_wire_1575)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_1952),
        .dout(new_Jinkela_wire_1953)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(_0170_),
        .c(new_Jinkela_wire_1965),
        .b(new_Jinkela_wire_1967)
    );

    spl4L new_Jinkela_splitter_202 (
        .a(new_Jinkela_wire_1976),
        .c(new_Jinkela_wire_1977),
        .e(new_Jinkela_wire_1978),
        .b(new_Jinkela_wire_1979),
        .d(new_Jinkela_wire_1980)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_1953),
        .dout(new_Jinkela_wire_1954)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(_0480_),
        .dout(new_Jinkela_wire_1586)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    spl4L new_Jinkela_splitter_199 (
        .a(new_Jinkela_wire_1967),
        .c(new_Jinkela_wire_1968),
        .e(new_Jinkela_wire_1969),
        .b(new_Jinkela_wire_1970),
        .d(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_1575),
        .dout(new_Jinkela_wire_1576)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_1954),
        .dout(new_Jinkela_wire_1955)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(_0272_),
        .dout(new_Jinkela_wire_1590)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_1955),
        .dout(new_Jinkela_wire_1956)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(new_Jinkela_wire_1564),
        .dout(new_Jinkela_wire_1565)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_1576),
        .dout(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_1956),
        .dout(new_Jinkela_wire_1957)
    );

    spl2 new_Jinkela_splitter_143 (
        .a(_0303_),
        .c(new_Jinkela_wire_1588),
        .b(new_Jinkela_wire_1589)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(new_Jinkela_wire_1577),
        .dout(new_Jinkela_wire_1578)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(_0285_),
        .c(new_Jinkela_wire_1986),
        .b(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_1590),
        .dout(new_Jinkela_wire_1591)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(new_Jinkela_wire_1958),
        .dout(new_Jinkela_wire_1959)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(_0348_),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(new_Jinkela_wire_1974),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(_0399_),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_1959),
        .dout(new_Jinkela_wire_1960)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(_0212_),
        .c(new_Jinkela_wire_1603),
        .b(new_Jinkela_wire_1604)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(new_Jinkela_wire_1591),
        .dout(new_Jinkela_wire_1592)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(_0393_),
        .dout(new_Jinkela_wire_1988)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    spl2 new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_265),
        .c(new_Jinkela_wire_266),
        .b(new_Jinkela_wire_267)
    );

    and_bi _0525_ (
        .a(new_Jinkela_wire_628),
        .b(new_Jinkela_wire_1105),
        .c(_0023_)
    );

    bfr new_Jinkela_buffer_1624 (
        .din(new_Jinkela_wire_2205),
        .dout(new_Jinkela_wire_2206)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(_0425_),
        .c(new_Jinkela_wire_2546),
        .b(new_Jinkela_wire_2547)
    );

    spl3L new_Jinkela_splitter_30 (
        .a(new_Jinkela_wire_272),
        .c(new_Jinkela_wire_273),
        .b(new_Jinkela_wire_274),
        .d(new_Jinkela_wire_275)
    );

    or_bb _0526_ (
        .a(_0023_),
        .b(new_Jinkela_wire_321),
        .c(_0024_)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_1671 (
        .din(new_Jinkela_wire_2252),
        .dout(new_Jinkela_wire_2253)
    );

    bfr new_Jinkela_buffer_1852 (
        .din(new_Jinkela_wire_2478),
        .dout(new_Jinkela_wire_2479)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    and_bi _0527_ (
        .a(new_Jinkela_wire_1354),
        .b(_0024_),
        .c(_0025_)
    );

    bfr new_Jinkela_buffer_1625 (
        .din(new_Jinkela_wire_2206),
        .dout(new_Jinkela_wire_2207)
    );

    bfr new_Jinkela_buffer_1861 (
        .din(new_Jinkela_wire_2515),
        .dout(new_Jinkela_wire_2516)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(new_Jinkela_wire_2540),
        .c(new_Jinkela_wire_2541),
        .b(new_Jinkela_wire_2542)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_281),
        .dout(new_Jinkela_wire_282)
    );

    or_bb _0528_ (
        .a(new_Jinkela_wire_312),
        .b(new_Jinkela_wire_629),
        .c(_0026_)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_779),
        .dout(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_1647 (
        .din(new_Jinkela_wire_2228),
        .dout(new_Jinkela_wire_2229)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_310),
        .c(new_Jinkela_wire_311),
        .b(new_Jinkela_wire_313)
    );

    bfr new_Jinkela_buffer_1853 (
        .din(new_Jinkela_wire_2479),
        .dout(new_Jinkela_wire_2480)
    );

    and_bi _0529_ (
        .a(new_Jinkela_wire_337),
        .b(new_Jinkela_wire_1657),
        .c(_0027_)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_1626 (
        .din(new_Jinkela_wire_2207),
        .dout(new_Jinkela_wire_2208)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_775),
        .c(new_Jinkela_wire_776),
        .b(new_Jinkela_wire_777)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_282),
        .dout(new_Jinkela_wire_283)
    );

    bfr new_Jinkela_buffer_1862 (
        .din(new_Jinkela_wire_2516),
        .dout(new_Jinkela_wire_2517)
    );

    or_bb _0530_ (
        .a(new_Jinkela_wire_314),
        .b(new_Jinkela_wire_630),
        .c(_0028_)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(new_Jinkela_wire_2480),
        .c(new_Jinkela_wire_2481),
        .b(new_Jinkela_wire_2482)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    and_bi _0531_ (
        .a(new_Jinkela_wire_854),
        .b(new_Jinkela_wire_2707),
        .c(_0029_)
    );

    bfr new_Jinkela_buffer_225 (
        .din(G82),
        .dout(new_Jinkela_wire_338)
    );

    bfr new_Jinkela_buffer_1627 (
        .din(new_Jinkela_wire_2208),
        .dout(new_Jinkela_wire_2209)
    );

    bfr new_Jinkela_buffer_1863 (
        .din(new_Jinkela_wire_2517),
        .dout(new_Jinkela_wire_2518)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_283),
        .dout(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_1887 (
        .din(_0492_),
        .dout(new_Jinkela_wire_2548)
    );

    or_bb _0532_ (
        .a(_0029_),
        .b(_0027_),
        .c(_0030_)
    );

    bfr new_Jinkela_buffer_1648 (
        .din(new_Jinkela_wire_2229),
        .dout(new_Jinkela_wire_2230)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    and_bi _0533_ (
        .a(new_Jinkela_wire_2192),
        .b(_0030_),
        .c(new_net_8)
    );

    bfr new_Jinkela_buffer_1628 (
        .din(new_Jinkela_wire_2209),
        .dout(new_Jinkela_wire_2210)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_777),
        .dout(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_1884 (
        .din(new_Jinkela_wire_2542),
        .dout(new_Jinkela_wire_2543)
    );

    and_bi _0534_ (
        .a(new_Jinkela_wire_383),
        .b(new_Jinkela_wire_2703),
        .c(_0031_)
    );

    bfr new_Jinkela_buffer_1672 (
        .din(new_Jinkela_wire_2253),
        .dout(new_Jinkela_wire_2254)
    );

    bfr new_Jinkela_buffer_1864 (
        .din(new_Jinkela_wire_2518),
        .dout(new_Jinkela_wire_2519)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    or_bb _0535_ (
        .a(new_Jinkela_wire_790),
        .b(new_Jinkela_wire_633),
        .c(_0032_)
    );

    bfr new_Jinkela_buffer_1629 (
        .din(new_Jinkela_wire_2210),
        .dout(new_Jinkela_wire_2211)
    );

    spl3L new_Jinkela_splitter_254 (
        .a(_0410_),
        .c(new_Jinkela_wire_2550),
        .b(new_Jinkela_wire_2551),
        .d(new_Jinkela_wire_2552)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    and_bi _0536_ (
        .a(new_Jinkela_wire_637),
        .b(new_Jinkela_wire_997),
        .c(_0033_)
    );

    bfr new_Jinkela_buffer_601 (
        .din(G22),
        .dout(new_Jinkela_wire_786)
    );

    bfr new_Jinkela_buffer_1649 (
        .din(new_Jinkela_wire_2230),
        .dout(new_Jinkela_wire_2231)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_311),
        .dout(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_1865 (
        .din(new_Jinkela_wire_2519),
        .dout(new_Jinkela_wire_2520)
    );

    or_bb _0537_ (
        .a(_0033_),
        .b(new_Jinkela_wire_319),
        .c(_0034_)
    );

    spl4L new_Jinkela_splitter_33 (
        .a(new_Jinkela_wire_313),
        .c(new_Jinkela_wire_314),
        .e(new_Jinkela_wire_315),
        .b(new_Jinkela_wire_318),
        .d(new_Jinkela_wire_323)
    );

    bfr new_Jinkela_buffer_1630 (
        .din(new_Jinkela_wire_2211),
        .dout(new_Jinkela_wire_2212)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    and_bi _0538_ (
        .a(new_Jinkela_wire_1607),
        .b(_0034_),
        .c(_0035_)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    spl3L new_Jinkela_splitter_222 (
        .a(_0411_),
        .c(new_Jinkela_wire_2262),
        .b(new_Jinkela_wire_2263),
        .d(new_Jinkela_wire_2264)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    bfr new_Jinkela_buffer_1674 (
        .din(new_Jinkela_wire_2255),
        .dout(new_Jinkela_wire_2256)
    );

    and_bi _0539_ (
        .a(_0031_),
        .b(new_Jinkela_wire_1949),
        .c(new_net_6)
    );

    bfr new_Jinkela_buffer_1631 (
        .din(new_Jinkela_wire_2212),
        .dout(new_Jinkela_wire_2213)
    );

    bfr new_Jinkela_buffer_1866 (
        .din(new_Jinkela_wire_2520),
        .dout(new_Jinkela_wire_2521)
    );

    bfr new_Jinkela_buffer_1885 (
        .din(new_Jinkela_wire_2543),
        .dout(new_Jinkela_wire_2544)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    and_bi _0540_ (
        .a(new_Jinkela_wire_644),
        .b(new_Jinkela_wire_581),
        .c(_0036_)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_1650 (
        .din(new_Jinkela_wire_2231),
        .dout(new_Jinkela_wire_2232)
    );

    bfr new_Jinkela_buffer_1867 (
        .din(new_Jinkela_wire_2521),
        .dout(new_Jinkela_wire_2522)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    and_bi _0541_ (
        .a(new_Jinkela_wire_634),
        .b(new_Jinkela_wire_994),
        .c(_0037_)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_329),
        .dout(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_1632 (
        .din(new_Jinkela_wire_2213),
        .dout(new_Jinkela_wire_2214)
    );

    bfr new_Jinkela_buffer_1889 (
        .din(_0098_),
        .dout(new_Jinkela_wire_2553)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    or_bb _0542_ (
        .a(_0037_),
        .b(new_Jinkela_wire_326),
        .c(_0038_)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    spl2 new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_315),
        .c(new_Jinkela_wire_316),
        .b(new_Jinkela_wire_317)
    );

    bfr new_Jinkela_buffer_1678 (
        .din(_0067_),
        .dout(new_Jinkela_wire_2265)
    );

    and_bi _0543_ (
        .a(new_Jinkela_wire_1411),
        .b(_0038_),
        .c(_0039_)
    );

    bfr new_Jinkela_buffer_1633 (
        .din(new_Jinkela_wire_2214),
        .dout(new_Jinkela_wire_2215)
    );

    bfr new_Jinkela_buffer_1868 (
        .din(new_Jinkela_wire_2522),
        .dout(new_Jinkela_wire_2523)
    );

    bfr new_Jinkela_buffer_1886 (
        .din(new_Jinkela_wire_2544),
        .dout(new_Jinkela_wire_2545)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    and_bi _0544_ (
        .a(new_Jinkela_wire_1256),
        .b(new_Jinkela_wire_1662),
        .c(_0040_)
    );

    bfr new_Jinkela_buffer_603 (
        .din(G35),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_1651 (
        .din(new_Jinkela_wire_2232),
        .dout(new_Jinkela_wire_2233)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    spl4L new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_318),
        .c(new_Jinkela_wire_319),
        .e(new_Jinkela_wire_320),
        .b(new_Jinkela_wire_321),
        .d(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_1869 (
        .din(new_Jinkela_wire_2523),
        .dout(new_Jinkela_wire_2524)
    );

    and_bi _0548_ (
        .a(new_Jinkela_wire_643),
        .b(new_Jinkela_wire_785),
        .c(_0043_)
    );

    bfr new_Jinkela_buffer_1634 (
        .din(new_Jinkela_wire_2215),
        .dout(new_Jinkela_wire_2216)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(_0119_),
        .c(new_Jinkela_wire_2554),
        .b(new_Jinkela_wire_2555)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_290),
        .dout(new_Jinkela_wire_291)
    );

    and_bi _0549_ (
        .a(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_662),
        .c(_0044_)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_1677 (
        .din(new_Jinkela_wire_2260),
        .dout(new_Jinkela_wire_2261)
    );

    bfr new_Jinkela_buffer_1675 (
        .din(new_Jinkela_wire_2256),
        .dout(new_Jinkela_wire_2257)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_1870 (
        .din(new_Jinkela_wire_2524),
        .dout(new_Jinkela_wire_2525)
    );

    or_bb _0550_ (
        .a(_0044_),
        .b(new_Jinkela_wire_327),
        .c(_0045_)
    );

    spl2 new_Jinkela_splitter_37 (
        .a(G157),
        .c(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_1635 (
        .din(new_Jinkela_wire_2216),
        .dout(new_Jinkela_wire_2217)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(_0333_),
        .c(new_Jinkela_wire_2556),
        .b(new_Jinkela_wire_2557)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    and_bi _0551_ (
        .a(new_Jinkela_wire_2600),
        .b(_0045_),
        .c(_0046_)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_1652 (
        .din(new_Jinkela_wire_2233),
        .dout(new_Jinkela_wire_2234)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    spl4L new_Jinkela_splitter_36 (
        .a(new_Jinkela_wire_323),
        .c(new_Jinkela_wire_324),
        .e(new_Jinkela_wire_325),
        .b(new_Jinkela_wire_326),
        .d(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_1871 (
        .din(new_Jinkela_wire_2525),
        .dout(new_Jinkela_wire_2526)
    );

    and_bi _0552_ (
        .a(new_Jinkela_wire_659),
        .b(new_Jinkela_wire_1666),
        .c(_0047_)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    and_bi _0553_ (
        .a(new_Jinkela_wire_598),
        .b(new_Jinkela_wire_2702),
        .c(_0048_)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(G115),
        .c(new_Jinkela_wire_791),
        .b(new_Jinkela_wire_792)
    );

    bfr new_Jinkela_buffer_1653 (
        .din(new_Jinkela_wire_2234),
        .dout(new_Jinkela_wire_2235)
    );

    bfr new_Jinkela_buffer_1872 (
        .din(new_Jinkela_wire_2526),
        .dout(new_Jinkela_wire_2527)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    or_bb _0554_ (
        .a(_0048_),
        .b(_0047_),
        .c(_0049_)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    spl3L new_Jinkela_splitter_65 (
        .a(G134),
        .c(new_Jinkela_wire_824),
        .b(new_Jinkela_wire_825),
        .d(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    spl2 new_Jinkela_splitter_221 (
        .a(new_Jinkela_wire_2257),
        .c(new_Jinkela_wire_2258),
        .b(new_Jinkela_wire_2259)
    );

    and_bi _0555_ (
        .a(new_Jinkela_wire_2622),
        .b(_0049_),
        .c(new_net_3)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_1654 (
        .din(new_Jinkela_wire_2235),
        .dout(new_Jinkela_wire_2236)
    );

    bfr new_Jinkela_buffer_1873 (
        .din(new_Jinkela_wire_2527),
        .dout(new_Jinkela_wire_2528)
    );

    spl3L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_757),
        .c(new_Jinkela_wire_758),
        .b(new_Jinkela_wire_759),
        .d(new_Jinkela_wire_760)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(_0481_),
        .c(new_Jinkela_wire_2558),
        .b(new_Jinkela_wire_2559)
    );

    and_bi _0556_ (
        .a(new_Jinkela_wire_645),
        .b(new_Jinkela_wire_987),
        .c(_0050_)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_1891 (
        .din(_0426_),
        .dout(new_Jinkela_wire_2561)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    and_bi _0557_ (
        .a(new_Jinkela_wire_622),
        .b(new_Jinkela_wire_486),
        .c(_0051_)
    );

    bfr new_Jinkela_buffer_1655 (
        .din(new_Jinkela_wire_2236),
        .dout(new_Jinkela_wire_2237)
    );

    bfr new_Jinkela_buffer_1890 (
        .din(new_Jinkela_wire_2559),
        .dout(new_Jinkela_wire_2560)
    );

    bfr new_Jinkela_buffer_644 (
        .din(G40),
        .dout(new_Jinkela_wire_843)
    );

    bfr new_Jinkela_buffer_229 (
        .din(G91),
        .dout(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_1874 (
        .din(new_Jinkela_wire_2528),
        .dout(new_Jinkela_wire_2529)
    );

    or_bb _0558_ (
        .a(_0051_),
        .b(new_Jinkela_wire_325),
        .c(_0052_)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_1679 (
        .din(new_Jinkela_wire_2265),
        .dout(new_Jinkela_wire_2266)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    bfr new_Jinkela_buffer_1680 (
        .din(_0380_),
        .dout(new_Jinkela_wire_2267)
    );

    and_bi _0559_ (
        .a(new_Jinkela_wire_1912),
        .b(_0052_),
        .c(_0053_)
    );

    bfr new_Jinkela_buffer_1656 (
        .din(new_Jinkela_wire_2237),
        .dout(new_Jinkela_wire_2238)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(_0105_),
        .c(new_Jinkela_wire_2563),
        .b(new_Jinkela_wire_2564)
    );

    bfr new_Jinkela_buffer_1875 (
        .din(new_Jinkela_wire_2529),
        .dout(new_Jinkela_wire_2530)
    );

    and_bi _0560_ (
        .a(new_Jinkela_wire_1055),
        .b(new_Jinkela_wire_1665),
        .c(_0054_)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_338),
        .dout(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_647 (
        .din(G2),
        .dout(new_Jinkela_wire_846)
    );

    bfr new_Jinkela_buffer_648 (
        .din(G25),
        .dout(new_Jinkela_wire_847)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    bfr new_Jinkela_buffer_1893 (
        .din(_0448_),
        .dout(new_Jinkela_wire_2565)
    );

    and_bi _0561_ (
        .a(new_Jinkela_wire_729),
        .b(new_Jinkela_wire_2711),
        .c(_0055_)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_1657 (
        .din(new_Jinkela_wire_2238),
        .dout(new_Jinkela_wire_2239)
    );

    bfr new_Jinkela_buffer_1892 (
        .din(new_Jinkela_wire_2561),
        .dout(new_Jinkela_wire_2562)
    );

    bfr new_Jinkela_buffer_1876 (
        .din(new_Jinkela_wire_2530),
        .dout(new_Jinkela_wire_2531)
    );

    or_bb _0562_ (
        .a(_0055_),
        .b(_0054_),
        .c(_0056_)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(new_net_3),
        .c(new_Jinkela_wire_2268),
        .b(new_Jinkela_wire_2271)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_827),
        .dout(new_Jinkela_wire_828)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    and_bi _0563_ (
        .a(new_Jinkela_wire_1857),
        .b(_0056_),
        .c(new_net_4)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    bfr new_Jinkela_buffer_1658 (
        .din(new_Jinkela_wire_2239),
        .dout(new_Jinkela_wire_2240)
    );

    bfr new_Jinkela_buffer_1877 (
        .din(new_Jinkela_wire_2531),
        .dout(new_Jinkela_wire_2532)
    );

    or_bb _0564_ (
        .a(new_Jinkela_wire_238),
        .b(new_Jinkela_wire_635),
        .c(_0057_)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_843),
        .dout(new_Jinkela_wire_844)
    );

    bfr new_Jinkela_buffer_1699 (
        .din(_0494_),
        .dout(new_Jinkela_wire_2294)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(new_Jinkela_wire_2268),
        .c(new_Jinkela_wire_2269),
        .b(new_Jinkela_wire_2270)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    spl2 new_Jinkela_splitter_259 (
        .a(_0122_),
        .c(new_Jinkela_wire_2567),
        .b(new_Jinkela_wire_2568)
    );

    and_bi _0565_ (
        .a(new_Jinkela_wire_638),
        .b(new_Jinkela_wire_1192),
        .c(_0058_)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    bfr new_Jinkela_buffer_1659 (
        .din(new_Jinkela_wire_2240),
        .dout(new_Jinkela_wire_2241)
    );

    bfr new_Jinkela_buffer_1878 (
        .din(new_Jinkela_wire_2532),
        .dout(new_Jinkela_wire_2533)
    );

    or_bb _0566_ (
        .a(_0058_),
        .b(new_Jinkela_wire_317),
        .c(_0059_)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_335),
        .dout(new_Jinkela_wire_336)
    );

    spl4L new_Jinkela_splitter_225 (
        .a(new_Jinkela_wire_2271),
        .c(new_Jinkela_wire_2272),
        .e(new_Jinkela_wire_2273),
        .b(new_Jinkela_wire_2274),
        .d(new_Jinkela_wire_2275)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_299),
        .dout(new_Jinkela_wire_300)
    );

    and_bi _0567_ (
        .a(new_Jinkela_wire_2700),
        .b(_0059_),
        .c(_0060_)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_1660 (
        .din(new_Jinkela_wire_2241),
        .dout(new_Jinkela_wire_2242)
    );

    bfr new_Jinkela_buffer_1894 (
        .din(_0227_),
        .dout(new_Jinkela_wire_2566)
    );

    bfr new_Jinkela_buffer_1879 (
        .din(new_Jinkela_wire_2533),
        .dout(new_Jinkela_wire_2534)
    );

    and_bi _0568_ (
        .a(new_Jinkela_wire_1265),
        .b(new_Jinkela_wire_1667),
        .c(_0061_)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_1706 (
        .din(_0451_),
        .dout(new_Jinkela_wire_2301)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_1895 (
        .din(new_net_22),
        .dout(new_Jinkela_wire_2569)
    );

    and_bi _0569_ (
        .a(new_Jinkela_wire_391),
        .b(new_Jinkela_wire_2708),
        .c(_0062_)
    );

    bfr new_Jinkela_buffer_1661 (
        .din(new_Jinkela_wire_2242),
        .dout(new_Jinkela_wire_2243)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_1135),
        .dout(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1141),
        .dout(new_Jinkela_wire_1142)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1139),
        .dout(new_Jinkela_wire_1140)
    );

    spl2 new_Jinkela_splitter_90 (
        .a(G156),
        .c(new_Jinkela_wire_1144),
        .b(new_Jinkela_wire_1145)
    );

    spl2 new_Jinkela_splitter_91 (
        .a(G153),
        .c(new_Jinkela_wire_1146),
        .b(new_Jinkela_wire_1147)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1148),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_889 (
        .din(G50),
        .dout(new_Jinkela_wire_1148)
    );

    spl3L new_Jinkela_splitter_95 (
        .a(G135),
        .c(new_Jinkela_wire_1173),
        .b(new_Jinkela_wire_1174),
        .d(new_Jinkela_wire_1175)
    );

    spl3L new_Jinkela_splitter_92 (
        .a(G138),
        .c(new_Jinkela_wire_1154),
        .b(new_Jinkela_wire_1155),
        .d(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1190),
        .dout(new_Jinkela_wire_1191)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1156),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_914 (
        .din(G71),
        .dout(new_Jinkela_wire_1190)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1151),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1176),
        .dout(new_Jinkela_wire_1177)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1152),
        .dout(new_Jinkela_wire_1153)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(G155),
        .c(new_Jinkela_wire_1197),
        .b(new_Jinkela_wire_1198)
    );

    bfr new_Jinkela_buffer_917 (
        .din(G85),
        .dout(new_Jinkela_wire_1193)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_1159),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1191),
        .dout(new_Jinkela_wire_1192)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1175),
        .dout(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    spl2 new_Jinkela_splitter_99 (
        .a(G53),
        .c(new_Jinkela_wire_1199),
        .b(new_Jinkela_wire_1200)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1177),
        .dout(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_1178),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    spl3L new_Jinkela_splitter_93 (
        .a(new_Jinkela_wire_1163),
        .c(new_Jinkela_wire_1164),
        .b(new_Jinkela_wire_1165),
        .d(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1193),
        .dout(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1166),
        .dout(new_Jinkela_wire_1167)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1179),
        .dout(new_Jinkela_wire_1180)
    );

    bfr new_Jinkela_buffer_949 (
        .din(G37),
        .dout(new_Jinkela_wire_1229)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1167),
        .dout(new_Jinkela_wire_1168)
    );

    spl3L new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_1168),
        .c(new_Jinkela_wire_1169),
        .b(new_Jinkela_wire_1170),
        .d(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1200),
        .dout(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_1194),
        .dout(new_Jinkela_wire_1195)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1171),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1181),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1195),
        .dout(new_Jinkela_wire_1196)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_207),
        .dout(new_Jinkela_wire_208)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_Jinkela_wire_1592),
        .dout(new_Jinkela_wire_1593)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(_0421_),
        .c(new_Jinkela_wire_1605),
        .b(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_1593),
        .dout(new_Jinkela_wire_1594)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(_0390_),
        .c(new_Jinkela_wire_1615),
        .b(new_Jinkela_wire_1616)
    );

    spl2 new_Jinkela_splitter_144 (
        .a(new_Jinkela_wire_1600),
        .c(new_Jinkela_wire_1601),
        .b(new_Jinkela_wire_1602)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_1594),
        .dout(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(_0032_),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(_0283_),
        .dout(new_Jinkela_wire_1608)
    );

    spl2 new_Jinkela_splitter_148 (
        .a(_0472_),
        .c(new_Jinkela_wire_1617),
        .b(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_Jinkela_wire_1608),
        .dout(new_Jinkela_wire_1609)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_1609),
        .dout(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(new_net_961),
        .dout(new_Jinkela_wire_1622)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_1610),
        .dout(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_1618),
        .dout(new_Jinkela_wire_1619)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_Jinkela_wire_1611),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(_0414_),
        .dout(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(new_Jinkela_wire_1622),
        .dout(new_Jinkela_wire_1623)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_1619),
        .dout(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_1613),
        .dout(new_Jinkela_wire_1614)
    );

    spl2 new_Jinkela_splitter_149 (
        .a(_0150_),
        .c(new_Jinkela_wire_1649),
        .b(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(new_Jinkela_wire_1620),
        .dout(new_Jinkela_wire_1621)
    );

    spl3L new_Jinkela_splitter_151 (
        .a(_0026_),
        .c(new_Jinkela_wire_1656),
        .b(new_Jinkela_wire_1658),
        .d(new_Jinkela_wire_1663)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(new_Jinkela_wire_1623),
        .dout(new_Jinkela_wire_1624)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_1639),
        .dout(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(new_Jinkela_wire_1624),
        .dout(new_Jinkela_wire_1625)
    );

    spl4L new_Jinkela_splitter_152 (
        .a(new_Jinkela_wire_1658),
        .c(new_Jinkela_wire_1659),
        .e(new_Jinkela_wire_1660),
        .b(new_Jinkela_wire_1661),
        .d(new_Jinkela_wire_1662)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_1625),
        .dout(new_Jinkela_wire_1626)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_1640),
        .dout(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_1626),
        .dout(new_Jinkela_wire_1627)
    );

    spl3L new_Jinkela_splitter_0 (
        .a(G131),
        .c(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_1),
        .d(new_Jinkela_wire_2)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_2),
        .dout(new_Jinkela_wire_3)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_13 (
        .din(G26),
        .dout(new_Jinkela_wire_19)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_1627),
        .dout(new_Jinkela_wire_1628)
    );

    bfr new_Jinkela_buffer_15 (
        .din(G16),
        .dout(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_1641),
        .dout(new_Jinkela_wire_1642)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_5),
        .dout(new_Jinkela_wire_6)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(new_Jinkela_wire_1628),
        .dout(new_Jinkela_wire_1629)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_19),
        .dout(new_Jinkela_wire_20)
    );

    spl4L new_Jinkela_splitter_150 (
        .a(new_Jinkela_wire_1651),
        .c(new_Jinkela_wire_1652),
        .e(new_Jinkela_wire_1653),
        .b(new_Jinkela_wire_1654),
        .d(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_3),
        .dout(new_Jinkela_wire_4)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_1629),
        .dout(new_Jinkela_wire_1630)
    );

    bfr new_Jinkela_buffer_17 (
        .din(G30),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(new_Jinkela_wire_1642),
        .dout(new_Jinkela_wire_1643)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_4),
        .dout(new_Jinkela_wire_5)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_1630),
        .dout(new_Jinkela_wire_1631)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    spl3L new_Jinkela_splitter_96 (
        .a(new_Jinkela_wire_1182),
        .c(new_Jinkela_wire_1183),
        .b(new_Jinkela_wire_1184),
        .d(new_Jinkela_wire_1185)
    );

    and_bi _0906_ (
        .a(new_Jinkela_wire_1071),
        .b(new_Jinkela_wire_1515),
        .c(_0379_)
    );

    bfr new_Jinkela_buffer_25 (
        .din(G57),
        .dout(new_Jinkela_wire_31)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_336),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_1960),
        .dout(new_Jinkela_wire_1961)
    );

    bfr new_Jinkela_buffer_1711 (
        .din(_0219_),
        .dout(new_Jinkela_wire_2308)
    );

    or_bb _0907_ (
        .a(_0379_),
        .b(new_Jinkela_wire_2261),
        .c(_0380_)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    spl4L new_Jinkela_splitter_203 (
        .a(new_Jinkela_wire_1981),
        .c(new_Jinkela_wire_1982),
        .e(new_Jinkela_wire_1983),
        .b(new_Jinkela_wire_1984),
        .d(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1185),
        .dout(new_Jinkela_wire_1186)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(_0373_),
        .dout(new_Jinkela_wire_1990)
    );

    bfr new_Jinkela_buffer_1662 (
        .din(new_Jinkela_wire_2243),
        .dout(new_Jinkela_wire_2244)
    );

    and_bi _0908_ (
        .a(new_Jinkela_wire_1101),
        .b(new_Jinkela_wire_2385),
        .c(_0381_)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_23),
        .dout(new_Jinkela_wire_24)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_1988),
        .dout(new_Jinkela_wire_1989)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_net_20),
        .dout(new_Jinkela_wire_1992)
    );

    and_bi _0909_ (
        .a(new_Jinkela_wire_1294),
        .b(new_Jinkela_wire_1479),
        .c(_0382_)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    spl3L new_Jinkela_splitter_100 (
        .a(G130),
        .c(new_Jinkela_wire_1232),
        .b(new_Jinkela_wire_1233),
        .d(new_Jinkela_wire_1234)
    );

    spl2 new_Jinkela_splitter_38 (
        .a(G106),
        .c(new_Jinkela_wire_348),
        .b(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1186),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_1663 (
        .din(new_Jinkela_wire_2244),
        .dout(new_Jinkela_wire_2245)
    );

    or_bb _0910_ (
        .a(new_Jinkela_wire_1446),
        .b(_0381_),
        .c(_0383_)
    );

    spl3L new_Jinkela_splitter_2 (
        .a(G12),
        .c(new_Jinkela_wire_37),
        .b(new_Jinkela_wire_40),
        .d(new_Jinkela_wire_45)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_340),
        .dout(new_Jinkela_wire_341)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_965 (
        .din(G46),
        .dout(new_Jinkela_wire_1251)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(new_net_959),
        .dout(new_Jinkela_wire_2009)
    );

    or_bb _0911_ (
        .a(_0383_),
        .b(new_Jinkela_wire_2267),
        .c(_0384_)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1229),
        .dout(new_Jinkela_wire_1230)
    );

    spl2 new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_1187),
        .c(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_1990),
        .dout(new_Jinkela_wire_1991)
    );

    bfr new_Jinkela_buffer_1664 (
        .din(new_Jinkela_wire_2245),
        .dout(new_Jinkela_wire_2246)
    );

    and_bi _0912_ (
        .a(new_Jinkela_wire_842),
        .b(new_Jinkela_wire_2184),
        .c(_0385_)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_24),
        .dout(new_Jinkela_wire_25)
    );

    bfr new_Jinkela_buffer_261 (
        .din(G56),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    bfr new_Jinkela_buffer_1720 (
        .din(new_net_965),
        .dout(new_Jinkela_wire_2317)
    );

    and_bi _0913_ (
        .a(new_Jinkela_wire_1122),
        .b(new_Jinkela_wire_1445),
        .c(_0386_)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(_0076_),
        .c(new_Jinkela_wire_2019),
        .b(new_Jinkela_wire_2020)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1201),
        .dout(new_Jinkela_wire_1202)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    bfr new_Jinkela_buffer_1665 (
        .din(new_Jinkela_wire_2246),
        .dout(new_Jinkela_wire_2247)
    );

    or_bb _0914_ (
        .a(new_Jinkela_wire_2130),
        .b(_0385_),
        .c(_0387_)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_31),
        .dout(new_Jinkela_wire_32)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_1202),
        .dout(new_Jinkela_wire_1203)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(new_net_954),
        .dout(new_Jinkela_wire_2021)
    );

    bfr new_Jinkela_buffer_1682 (
        .din(new_Jinkela_wire_2276),
        .dout(new_Jinkela_wire_2277)
    );

    and_bi _0915_ (
        .a(new_Jinkela_wire_42),
        .b(new_Jinkela_wire_1142),
        .c(_0388_)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_10),
        .dout(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1234),
        .dout(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(new_Jinkela_wire_1993),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(new_Jinkela_wire_2009),
        .dout(new_Jinkela_wire_2010)
    );

    and_bi _0916_ (
        .a(new_Jinkela_wire_56),
        .b(new_Jinkela_wire_1815),
        .c(_0389_)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_25),
        .dout(new_Jinkela_wire_26)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1230),
        .dout(new_Jinkela_wire_1231)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1203),
        .dout(new_Jinkela_wire_1204)
    );

    and_bi _0917_ (
        .a(new_Jinkela_wire_2137),
        .b(_0389_),
        .c(_0390_)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_1667 (
        .din(new_Jinkela_wire_2248),
        .dout(new_Jinkela_wire_2249)
    );

    and_bi _0918_ (
        .a(new_Jinkela_wire_569),
        .b(new_Jinkela_wire_1615),
        .c(_0391_)
    );

    spl2 new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_37),
        .c(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_39)
    );

    bfr new_Jinkela_buffer_267 (
        .din(G13),
        .dout(new_Jinkela_wire_384)
    );

    spl4L new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_40),
        .c(new_Jinkela_wire_41),
        .e(new_Jinkela_wire_42),
        .b(new_Jinkela_wire_43),
        .d(new_Jinkela_wire_44)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_1204),
        .dout(new_Jinkela_wire_1205)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(new_Jinkela_wire_2021),
        .dout(new_Jinkela_wire_2022)
    );

    and_bi _0919_ (
        .a(new_Jinkela_wire_570),
        .b(new_Jinkela_wire_1616),
        .c(_0392_)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_350),
        .dout(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_971 (
        .din(G41),
        .dout(new_Jinkela_wire_1257)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    or_bb _0920_ (
        .a(_0392_),
        .b(_0391_),
        .c(_0393_)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_Jinkela_wire_2010),
        .dout(new_Jinkela_wire_2011)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1205),
        .dout(new_Jinkela_wire_1206)
    );

    bfr new_Jinkela_buffer_1707 (
        .din(new_Jinkela_wire_2301),
        .dout(new_Jinkela_wire_2302)
    );

    or_bb _0921_ (
        .a(new_Jinkela_wire_1989),
        .b(_0387_),
        .c(_0394_)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    bfr new_Jinkela_buffer_269 (
        .din(G60),
        .dout(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(new_Jinkela_wire_1996),
        .dout(new_Jinkela_wire_1997)
    );

    bfr new_Jinkela_buffer_1669 (
        .din(new_Jinkela_wire_2250),
        .dout(new_Jinkela_wire_2251)
    );

    or_bb _0922_ (
        .a(_0394_),
        .b(_0384_),
        .c(_0395_)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_32),
        .dout(new_Jinkela_wire_33)
    );

    bfr new_Jinkela_buffer_1702 (
        .din(new_Jinkela_wire_2296),
        .dout(new_Jinkela_wire_2297)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1206),
        .dout(new_Jinkela_wire_1207)
    );

    bfr new_Jinkela_buffer_1684 (
        .din(new_Jinkela_wire_2278),
        .dout(new_Jinkela_wire_2279)
    );

    or_bb _0923_ (
        .a(_0395_),
        .b(_0377_),
        .c(_0396_)
    );

    spl3L new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_14),
        .c(new_Jinkela_wire_15),
        .b(new_Jinkela_wire_16),
        .d(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1251),
        .dout(new_Jinkela_wire_1252)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(new_Jinkela_wire_1997),
        .dout(new_Jinkela_wire_1998)
    );

    or_bb _0924_ (
        .a(_0396_),
        .b(new_Jinkela_wire_1480),
        .c(_0397_)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1235),
        .dout(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1207),
        .dout(new_Jinkela_wire_1208)
    );

    bfr new_Jinkela_buffer_1685 (
        .din(new_Jinkela_wire_2279),
        .dout(new_Jinkela_wire_2280)
    );

    or_bb _0925_ (
        .a(_0397_),
        .b(new_Jinkela_wire_2490),
        .c(new_net_21)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(new_Jinkela_wire_1998),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(_0417_),
        .dout(new_Jinkela_wire_2048)
    );

    and_bi _0926_ (
        .a(new_Jinkela_wire_158),
        .b(new_Jinkela_wire_2452),
        .c(_0398_)
    );

    bfr new_Jinkela_buffer_974 (
        .din(G49),
        .dout(new_Jinkela_wire_1260)
    );

    bfr new_Jinkela_buffer_1703 (
        .din(new_Jinkela_wire_2297),
        .dout(new_Jinkela_wire_2298)
    );

    bfr new_Jinkela_buffer_45 (
        .din(G107),
        .dout(new_Jinkela_wire_77)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1208),
        .dout(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_1686 (
        .din(new_Jinkela_wire_2280),
        .dout(new_Jinkela_wire_2281)
    );

    and_bi _0927_ (
        .a(new_Jinkela_wire_210),
        .b(new_Jinkela_wire_1501),
        .c(_0399_)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_354),
        .dout(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(new_Jinkela_wire_2012),
        .dout(new_Jinkela_wire_2013)
    );

    and_bi _0928_ (
        .a(new_Jinkela_wire_1691),
        .b(new_Jinkela_wire_1601),
        .c(_0400_)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_33),
        .dout(new_Jinkela_wire_34)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1236),
        .dout(new_Jinkela_wire_1237)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1209),
        .dout(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_1687 (
        .din(new_Jinkela_wire_2281),
        .dout(new_Jinkela_wire_2282)
    );

    bfr new_Jinkela_buffer_1708 (
        .din(new_Jinkela_wire_2302),
        .dout(new_Jinkela_wire_2303)
    );

    and_bi _0929_ (
        .a(new_Jinkela_wire_1690),
        .b(new_Jinkela_wire_1602),
        .c(_0401_)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    spl2 new_Jinkela_splitter_39 (
        .a(G148),
        .c(new_Jinkela_wire_392),
        .b(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_2000),
        .dout(new_Jinkela_wire_2001)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(_0097_),
        .c(new_Jinkela_wire_2057),
        .b(new_Jinkela_wire_2058)
    );

    and_bi _0930_ (
        .a(_0400_),
        .b(_0401_),
        .c(_0402_)
    );

    bfr new_Jinkela_buffer_42 (
        .din(G147),
        .dout(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1252),
        .dout(new_Jinkela_wire_1253)
    );

    spl2 new_Jinkela_splitter_40 (
        .a(G64),
        .c(new_Jinkela_wire_394),
        .b(new_Jinkela_wire_395)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1210),
        .dout(new_Jinkela_wire_1211)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(new_net_5),
        .c(new_Jinkela_wire_2059),
        .b(new_Jinkela_wire_2061)
    );

    and_bi _0931_ (
        .a(new_Jinkela_wire_2484),
        .b(new_Jinkela_wire_1533),
        .c(_0403_)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_381),
        .dout(new_Jinkela_wire_382)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(new_Jinkela_wire_2001),
        .dout(new_Jinkela_wire_2002)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_2013),
        .dout(new_Jinkela_wire_2014)
    );

    and_bi _0932_ (
        .a(new_Jinkela_wire_1532),
        .b(new_Jinkela_wire_2483),
        .c(_0404_)
    );

    bfr new_Jinkela_buffer_39 (
        .din(G73),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1211),
        .dout(new_Jinkela_wire_1212)
    );

    bfr new_Jinkela_buffer_1689 (
        .din(new_Jinkela_wire_2283),
        .dout(new_Jinkela_wire_2284)
    );

    and_bi _0933_ (
        .a(_0403_),
        .b(_0404_),
        .c(_0405_)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_35),
        .dout(new_Jinkela_wire_36)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_386),
        .dout(new_Jinkela_wire_387)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_Jinkela_wire_2002),
        .dout(new_Jinkela_wire_2003)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    or_bb _0934_ (
        .a(new_Jinkela_wire_1582),
        .b(new_Jinkela_wire_1474),
        .c(_0406_)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1237),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1212),
        .dout(new_Jinkela_wire_1213)
    );

    bfr new_Jinkela_buffer_1690 (
        .din(new_Jinkela_wire_2284),
        .dout(new_Jinkela_wire_2285)
    );

    and_bi _0935_ (
        .a(new_Jinkela_wire_1475),
        .b(new_Jinkela_wire_1583),
        .c(_0407_)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(new_Jinkela_wire_2014),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(new_Jinkela_wire_2003),
        .dout(new_Jinkela_wire_2004)
    );

    and_bi _0936_ (
        .a(_0406_),
        .b(_0407_),
        .c(_0408_)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_70),
        .dout(new_Jinkela_wire_71)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1238),
        .dout(new_Jinkela_wire_1239)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1213),
        .dout(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_1691 (
        .din(new_Jinkela_wire_2285),
        .dout(new_Jinkela_wire_2286)
    );

    bfr new_Jinkela_buffer_1713 (
        .din(new_Jinkela_wire_2309),
        .dout(new_Jinkela_wire_2310)
    );

    and_bi _0937_ (
        .a(new_Jinkela_wire_176),
        .b(_0408_),
        .c(_0409_)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_Jinkela_wire_2048),
        .dout(new_Jinkela_wire_2049)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_50),
        .dout(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_359),
        .dout(new_Jinkela_wire_360)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1257),
        .dout(new_Jinkela_wire_1258)
    );

    or_bb _0938_ (
        .a(_0409_),
        .b(new_Jinkela_wire_1961),
        .c(new_net_22)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_49),
        .dout(new_Jinkela_wire_50)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1253),
        .dout(new_Jinkela_wire_1254)
    );

    spl4L new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_45),
        .c(new_Jinkela_wire_46),
        .e(new_Jinkela_wire_47),
        .b(new_Jinkela_wire_48),
        .d(new_Jinkela_wire_49)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1214),
        .dout(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_2004),
        .dout(new_Jinkela_wire_2005)
    );

    or_bb _0939_ (
        .a(new_Jinkela_wire_2645),
        .b(new_Jinkela_wire_1273),
        .c(_0410_)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_77),
        .dout(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_387),
        .dout(new_Jinkela_wire_388)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(new_Jinkela_wire_2005),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(new_Jinkela_wire_2015),
        .dout(new_Jinkela_wire_2016)
    );

    or_bb _0940_ (
        .a(new_Jinkela_wire_1752),
        .b(new_Jinkela_wire_30),
        .c(_0411_)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1239),
        .dout(new_Jinkela_wire_1240)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(new_net_13),
        .c(new_Jinkela_wire_2342),
        .b(new_Jinkela_wire_2343)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1215),
        .dout(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_1693 (
        .din(new_Jinkela_wire_2287),
        .dout(new_Jinkela_wire_2288)
    );

    and_ii _0941_ (
        .a(new_Jinkela_wire_2262),
        .b(new_Jinkela_wire_2550),
        .c(_0412_)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_2023),
        .dout(new_Jinkela_wire_2024)
    );

    bfr new_Jinkela_buffer_49 (
        .din(G75),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(new_Jinkela_wire_2006),
        .c(new_Jinkela_wire_2007),
        .b(new_Jinkela_wire_2008)
    );

    or_bb _0942_ (
        .a(new_Jinkela_wire_1743),
        .b(new_Jinkela_wire_446),
        .c(_0413_)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_980 (
        .din(G127),
        .dout(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_1694 (
        .din(new_Jinkela_wire_2288),
        .dout(new_Jinkela_wire_2289)
    );

    bfr new_Jinkela_buffer_1710 (
        .din(new_Jinkela_wire_2304),
        .dout(new_Jinkela_wire_2305)
    );

    or_bb _0943_ (
        .a(new_Jinkela_wire_2143),
        .b(new_Jinkela_wire_229),
        .c(_0414_)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_388),
        .dout(new_Jinkela_wire_389)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(new_Jinkela_wire_73),
        .c(new_Jinkela_wire_74),
        .b(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(new_net_4),
        .c(new_Jinkela_wire_2360),
        .b(new_Jinkela_wire_2361)
    );

    or_bb _0944_ (
        .a(new_Jinkela_wire_2263),
        .b(new_Jinkela_wire_2551),
        .c(_0415_)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1240),
        .dout(new_Jinkela_wire_1241)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_2016),
        .dout(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1217),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_1695 (
        .din(new_Jinkela_wire_2289),
        .dout(new_Jinkela_wire_2290)
    );

    or_bb _0945_ (
        .a(new_Jinkela_wire_1352),
        .b(new_Jinkela_wire_447),
        .c(_0416_)
    );

    bfr new_Jinkela_buffer_303 (
        .din(G20),
        .dout(new_Jinkela_wire_424)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(new_Jinkela_wire_2017),
        .dout(new_Jinkela_wire_2018)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_75),
        .dout(new_Jinkela_wire_76)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_363),
        .dout(new_Jinkela_wire_364)
    );

    spl2 new_Jinkela_splitter_226 (
        .a(new_Jinkela_wire_2305),
        .c(new_Jinkela_wire_2306),
        .b(new_Jinkela_wire_2307)
    );

    or_bb _0946_ (
        .a(new_Jinkela_wire_1746),
        .b(new_Jinkela_wire_2368),
        .c(_0417_)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1254),
        .dout(new_Jinkela_wire_1255)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_2024),
        .dout(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1218),
        .dout(new_Jinkela_wire_1219)
    );

    or_bb _0947_ (
        .a(new_Jinkela_wire_2144),
        .b(new_Jinkela_wire_574),
        .c(_0418_)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_2049),
        .dout(new_Jinkela_wire_2050)
    );

    bfr new_Jinkela_buffer_1696 (
        .din(new_Jinkela_wire_2290),
        .dout(new_Jinkela_wire_2291)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_844),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_650 (
        .din(G58),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_829),
        .dout(new_Jinkela_wire_830)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_830),
        .dout(new_Jinkela_wire_831)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_803),
        .dout(new_Jinkela_wire_804)
    );

    bfr new_Jinkela_buffer_656 (
        .din(G111),
        .dout(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_831),
        .dout(new_Jinkela_wire_832)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_804),
        .dout(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_832),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_660 (
        .din(G100),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    spl3L new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_835),
        .c(new_Jinkela_wire_836),
        .b(new_Jinkela_wire_837),
        .d(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_838),
        .dout(new_Jinkela_wire_839)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    spl3L new_Jinkela_splitter_68 (
        .a(G126),
        .c(new_Jinkela_wire_863),
        .b(new_Jinkela_wire_864),
        .d(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_675 (
        .din(G70),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_1880 (
        .din(new_Jinkela_wire_2534),
        .dout(new_Jinkela_wire_2535)
    );

    or_bb _0738_ (
        .a(_0224_),
        .b(_0223_),
        .c(_0225_)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(_0082_),
        .dout(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(_0309_),
        .dout(new_Jinkela_wire_1714)
    );

    and_bi _0739_ (
        .a(new_Jinkela_wire_2715),
        .b(_0225_),
        .c(_0226_)
    );

    spl3L new_Jinkela_splitter_262 (
        .a(new_Jinkela_wire_2576),
        .c(new_Jinkela_wire_2577),
        .b(new_Jinkela_wire_2578),
        .d(new_Jinkela_wire_2579)
    );

    bfr new_Jinkela_buffer_1881 (
        .din(new_Jinkela_wire_2535),
        .dout(new_Jinkela_wire_2536)
    );

    and_bi _0740_ (
        .a(new_Jinkela_wire_623),
        .b(new_Jinkela_wire_648),
        .c(_0227_)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(new_net_0),
        .c(new_Jinkela_wire_2575),
        .b(new_Jinkela_wire_2576)
    );

    and_bi _0741_ (
        .a(new_Jinkela_wire_640),
        .b(new_Jinkela_wire_530),
        .c(_0228_)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(_0286_),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_1920 (
        .din(_0306_),
        .dout(new_Jinkela_wire_2603)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_1706),
        .dout(new_Jinkela_wire_1707)
    );

    bfr new_Jinkela_buffer_1882 (
        .din(new_Jinkela_wire_2536),
        .dout(new_Jinkela_wire_2537)
    );

    or_bb _0742_ (
        .a(_0228_),
        .b(new_Jinkela_wire_324),
        .c(_0229_)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_1711),
        .dout(new_Jinkela_wire_1712)
    );

    bfr new_Jinkela_buffer_1896 (
        .din(new_Jinkela_wire_2569),
        .dout(new_Jinkela_wire_2570)
    );

    and_bi _0743_ (
        .a(new_Jinkela_wire_2566),
        .b(_0229_),
        .c(_0230_)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_1707),
        .dout(new_Jinkela_wire_1708)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(new_Jinkela_wire_2537),
        .c(new_Jinkela_wire_2538),
        .b(new_Jinkela_wire_2539)
    );

    and_bi _0744_ (
        .a(new_Jinkela_wire_527),
        .b(new_Jinkela_wire_1660),
        .c(_0231_)
    );

    bfr new_Jinkela_buffer_1897 (
        .din(new_Jinkela_wire_2570),
        .dout(new_Jinkela_wire_2571)
    );

    and_bi _0745_ (
        .a(new_Jinkela_wire_431),
        .b(new_Jinkela_wire_2712),
        .c(_0232_)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(_0456_),
        .dout(new_Jinkela_wire_1715)
    );

    spl2 new_Jinkela_splitter_162 (
        .a(new_Jinkela_wire_1708),
        .c(new_Jinkela_wire_1709),
        .b(new_Jinkela_wire_1710)
    );

    or_bb _0746_ (
        .a(_0232_),
        .b(_0231_),
        .c(_0233_)
    );

    and_bi _0747_ (
        .a(new_Jinkela_wire_2127),
        .b(_0233_),
        .c(_0234_)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(_0241_),
        .dout(new_Jinkela_wire_1717)
    );

    bfr new_Jinkela_buffer_1919 (
        .din(_0043_),
        .dout(new_Jinkela_wire_2600)
    );

    bfr new_Jinkela_buffer_1898 (
        .din(new_Jinkela_wire_2571),
        .dout(new_Jinkela_wire_2572)
    );

    and_bi _0748_ (
        .a(new_Jinkela_wire_2454),
        .b(new_Jinkela_wire_1723),
        .c(_0235_)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_1712),
        .dout(new_Jinkela_wire_1713)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(_0366_),
        .c(new_Jinkela_wire_2601),
        .b(new_Jinkela_wire_2602)
    );

    and_bi _0749_ (
        .a(new_Jinkela_wire_2455),
        .b(new_Jinkela_wire_1724),
        .c(_0236_)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_1715),
        .dout(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_1921 (
        .din(new_Jinkela_wire_2603),
        .dout(new_Jinkela_wire_2604)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(new_Jinkela_wire_2572),
        .c(new_Jinkela_wire_2573),
        .b(new_Jinkela_wire_2574)
    );

    and_bi _0750_ (
        .a(_0235_),
        .b(_0236_),
        .c(_0237_)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(_0234_),
        .c(new_Jinkela_wire_1718),
        .b(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(_0094_),
        .dout(new_Jinkela_wire_1732)
    );

    and_ii _0751_ (
        .a(new_Jinkela_wire_1868),
        .b(new_Jinkela_wire_2458),
        .c(_0238_)
    );

    spl2 new_Jinkela_splitter_166 (
        .a(_0073_),
        .c(new_Jinkela_wire_1730),
        .b(new_Jinkela_wire_1731)
    );

    and_bb _0752_ (
        .a(new_Jinkela_wire_1867),
        .b(new_Jinkela_wire_2461),
        .c(_0239_)
    );

    bfr new_Jinkela_buffer_1899 (
        .din(new_Jinkela_wire_2579),
        .dout(new_Jinkela_wire_2580)
    );

    or_bb _0753_ (
        .a(_0239_),
        .b(_0238_),
        .c(_0240_)
    );

    bfr new_Jinkela_buffer_1900 (
        .din(new_Jinkela_wire_2580),
        .dout(new_Jinkela_wire_2581)
    );

    spl2 new_Jinkela_splitter_169 (
        .a(_0412_),
        .c(new_Jinkela_wire_1739),
        .b(new_Jinkela_wire_1741)
    );

    and_bi _0754_ (
        .a(new_Jinkela_wire_642),
        .b(new_Jinkela_wire_845),
        .c(_0241_)
    );

    spl2 new_Jinkela_splitter_164 (
        .a(new_Jinkela_wire_1718),
        .c(new_Jinkela_wire_1719),
        .b(new_Jinkela_wire_1720)
    );

    bfr new_Jinkela_buffer_1926 (
        .din(_0275_),
        .dout(new_Jinkela_wire_2609)
    );

    and_bi _0755_ (
        .a(new_Jinkela_wire_621),
        .b(new_Jinkela_wire_611),
        .c(_0242_)
    );

    spl4L new_Jinkela_splitter_165 (
        .a(new_Jinkela_wire_1721),
        .c(new_Jinkela_wire_1722),
        .e(new_Jinkela_wire_1723),
        .b(new_Jinkela_wire_1724),
        .d(new_Jinkela_wire_1725)
    );

    bfr new_Jinkela_buffer_1901 (
        .din(new_Jinkela_wire_2581),
        .dout(new_Jinkela_wire_2582)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(new_Jinkela_wire_1725),
        .dout(new_Jinkela_wire_1726)
    );

    or_bb _0756_ (
        .a(_0242_),
        .b(new_Jinkela_wire_320),
        .c(_0243_)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(_0324_),
        .c(new_Jinkela_wire_2610),
        .b(new_Jinkela_wire_2611)
    );

    spl2 new_Jinkela_splitter_168 (
        .a(_0091_),
        .c(new_Jinkela_wire_1737),
        .b(new_Jinkela_wire_1738)
    );

    bfr new_Jinkela_buffer_1927 (
        .din(_0304_),
        .dout(new_Jinkela_wire_2612)
    );

    and_bi _0757_ (
        .a(new_Jinkela_wire_1717),
        .b(_0243_),
        .c(_0244_)
    );

    bfr new_Jinkela_buffer_1902 (
        .din(new_Jinkela_wire_2582),
        .dout(new_Jinkela_wire_2583)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(new_Jinkela_wire_1732),
        .dout(new_Jinkela_wire_1733)
    );

    and_bi _0758_ (
        .a(new_Jinkela_wire_1153),
        .b(new_Jinkela_wire_1659),
        .c(_0245_)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_1739),
        .dout(new_Jinkela_wire_1740)
    );

    bfr new_Jinkela_buffer_1922 (
        .din(new_Jinkela_wire_2604),
        .dout(new_Jinkela_wire_2605)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(new_Jinkela_wire_1726),
        .dout(new_Jinkela_wire_1727)
    );

    and_bi _0759_ (
        .a(new_Jinkela_wire_773),
        .b(new_Jinkela_wire_2713),
        .c(_0246_)
    );

    bfr new_Jinkela_buffer_1903 (
        .din(new_Jinkela_wire_2583),
        .dout(new_Jinkela_wire_2584)
    );

    or_bb _0760_ (
        .a(_0246_),
        .b(_0245_),
        .c(_0247_)
    );

    spl4L new_Jinkela_splitter_171 (
        .a(_0416_),
        .c(new_Jinkela_wire_1746),
        .e(new_Jinkela_wire_1747),
        .b(new_Jinkela_wire_1748),
        .d(new_Jinkela_wire_1749)
    );

    bfr new_Jinkela_buffer_1930 (
        .din(_0046_),
        .dout(new_Jinkela_wire_2621)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(new_Jinkela_wire_1727),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_1928 (
        .din(new_Jinkela_wire_2612),
        .dout(new_Jinkela_wire_2613)
    );

    and_bi _0761_ (
        .a(new_Jinkela_wire_2388),
        .b(_0247_),
        .c(_0248_)
    );

    bfr new_Jinkela_buffer_1904 (
        .din(new_Jinkela_wire_2584),
        .dout(new_Jinkela_wire_2585)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(new_Jinkela_wire_1733),
        .dout(new_Jinkela_wire_1734)
    );

    and_ii _0762_ (
        .a(new_Jinkela_wire_1504),
        .b(new_Jinkela_wire_1522),
        .c(_0249_)
    );

    bfr new_Jinkela_buffer_1923 (
        .din(new_Jinkela_wire_2605),
        .dout(new_Jinkela_wire_2606)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(new_Jinkela_wire_1728),
        .dout(new_Jinkela_wire_1729)
    );

    and_bb _0763_ (
        .a(new_Jinkela_wire_1500),
        .b(new_Jinkela_wire_1523),
        .c(_0250_)
    );

    bfr new_Jinkela_buffer_1905 (
        .din(new_Jinkela_wire_2585),
        .dout(new_Jinkela_wire_2586)
    );

    and_bi _0764_ (
        .a(_0249_),
        .b(_0250_),
        .c(_0251_)
    );

    spl3L new_Jinkela_splitter_173 (
        .a(new_net_1),
        .c(new_Jinkela_wire_1752),
        .b(new_Jinkela_wire_1753),
        .d(new_Jinkela_wire_1754)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(new_Jinkela_wire_1734),
        .c(new_Jinkela_wire_1735),
        .b(new_Jinkela_wire_1736)
    );

    or_bb _0765_ (
        .a(new_Jinkela_wire_2513),
        .b(new_Jinkela_wire_2175),
        .c(_0252_)
    );

    bfr new_Jinkela_buffer_1906 (
        .din(new_Jinkela_wire_2586),
        .dout(new_Jinkela_wire_2587)
    );

    and_bi _0766_ (
        .a(new_Jinkela_wire_2176),
        .b(new_Jinkela_wire_2514),
        .c(_0253_)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(_0100_),
        .c(new_Jinkela_wire_1750),
        .b(new_Jinkela_wire_1751)
    );

    bfr new_Jinkela_buffer_1924 (
        .din(new_Jinkela_wire_2606),
        .dout(new_Jinkela_wire_2607)
    );

    spl4L new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_1741),
        .c(new_Jinkela_wire_1742),
        .e(new_Jinkela_wire_1743),
        .b(new_Jinkela_wire_1744),
        .d(new_Jinkela_wire_1745)
    );

    and_bi _0767_ (
        .a(_0252_),
        .b(_0253_),
        .c(_0254_)
    );

    bfr new_Jinkela_buffer_1907 (
        .din(new_Jinkela_wire_2587),
        .dout(new_Jinkela_wire_2588)
    );

    or_bb _0768_ (
        .a(new_Jinkela_wire_1697),
        .b(new_Jinkela_wire_1695),
        .c(_0255_)
    );

    spl2 new_Jinkela_splitter_265 (
        .a(_0200_),
        .c(new_Jinkela_wire_2614),
        .b(new_Jinkela_wire_2616)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(new_Jinkela_wire_1754),
        .dout(new_Jinkela_wire_1755)
    );

    and_bb _0769_ (
        .a(new_Jinkela_wire_1698),
        .b(new_Jinkela_wire_1696),
        .c(_0256_)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(_0358_),
        .dout(new_Jinkela_wire_1778)
    );

    bfr new_Jinkela_buffer_1908 (
        .din(new_Jinkela_wire_2588),
        .dout(new_Jinkela_wire_2589)
    );

    and_bi _0770_ (
        .a(_0255_),
        .b(_0256_),
        .c(_0257_)
    );

    bfr new_Jinkela_buffer_1925 (
        .din(new_Jinkela_wire_2607),
        .dout(new_Jinkela_wire_2608)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_1755),
        .dout(new_Jinkela_wire_1756)
    );

    and_bi _0771_ (
        .a(new_Jinkela_wire_2488),
        .b(new_Jinkela_wire_2494),
        .c(_0258_)
    );

    bfr new_Jinkela_buffer_1909 (
        .din(new_Jinkela_wire_2589),
        .dout(new_Jinkela_wire_2590)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_1778),
        .dout(new_Jinkela_wire_1779)
    );

    and_bi _0772_ (
        .a(new_Jinkela_wire_2495),
        .b(new_Jinkela_wire_2489),
        .c(_0259_)
    );

    bfr new_Jinkela_buffer_1932 (
        .din(_0278_),
        .dout(new_Jinkela_wire_2625)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(_0317_),
        .dout(new_Jinkela_wire_1787)
    );

    or_bb _0773_ (
        .a(_0259_),
        .b(new_Jinkela_wire_1324),
        .c(_0260_)
    );

    bfr new_Jinkela_buffer_1910 (
        .din(new_Jinkela_wire_2590),
        .dout(new_Jinkela_wire_2591)
    );

    and_bi _0774_ (
        .a(new_Jinkela_wire_1675),
        .b(_0260_),
        .c(new_net_16)
    );

    spl4L new_Jinkela_splitter_266 (
        .a(new_Jinkela_wire_2616),
        .c(new_Jinkela_wire_2617),
        .e(new_Jinkela_wire_2618),
        .b(new_Jinkela_wire_2619),
        .d(new_Jinkela_wire_2620)
    );

    or_bb _0775_ (
        .a(new_Jinkela_wire_1751),
        .b(new_Jinkela_wire_2058),
        .c(new_net_965)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    bfr new_Jinkela_buffer_1911 (
        .din(new_Jinkela_wire_2591),
        .dout(new_Jinkela_wire_2592)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_net_950),
        .dout(new_Jinkela_wire_1796)
    );

    or_bb _0776_ (
        .a(new_Jinkela_wire_846),
        .b(new_Jinkela_wire_889),
        .c(_0261_)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_1779),
        .dout(new_Jinkela_wire_1780)
    );

    spl2 new_Jinkela_splitter_267 (
        .a(_0134_),
        .c(new_Jinkela_wire_2623),
        .b(new_Jinkela_wire_2624)
    );

    or_bb _0777_ (
        .a(_0261_),
        .b(new_Jinkela_wire_453),
        .c(new_net_952)
    );

    spl3L new_Jinkela_splitter_174 (
        .a(new_Jinkela_wire_1757),
        .c(new_Jinkela_wire_1758),
        .b(new_Jinkela_wire_1759),
        .d(new_Jinkela_wire_1760)
    );

    bfr new_Jinkela_buffer_1912 (
        .din(new_Jinkela_wire_2592),
        .dout(new_Jinkela_wire_2593)
    );

    or_bb _0778_ (
        .a(new_Jinkela_wire_951),
        .b(new_Jinkela_wire_891),
        .c(new_net_10)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_1787),
        .dout(new_Jinkela_wire_1788)
    );

    bfr new_Jinkela_buffer_1929 (
        .din(new_Jinkela_wire_2614),
        .dout(new_Jinkela_wire_2615)
    );

    or_bb _0779_ (
        .a(new_Jinkela_wire_2672),
        .b(new_Jinkela_wire_776),
        .c(new_net_957)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_1760),
        .dout(new_Jinkela_wire_1761)
    );

    bfr new_Jinkela_buffer_1913 (
        .din(new_Jinkela_wire_2593),
        .dout(new_Jinkela_wire_2594)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(_0301_),
        .dout(new_Jinkela_wire_1668)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_1631),
        .dout(new_Jinkela_wire_1632)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(new_Jinkela_wire_1632),
        .dout(new_Jinkela_wire_1633)
    );

    spl4L new_Jinkela_splitter_153 (
        .a(new_Jinkela_wire_1663),
        .c(new_Jinkela_wire_1664),
        .e(new_Jinkela_wire_1665),
        .b(new_Jinkela_wire_1666),
        .d(new_Jinkela_wire_1667)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(new_Jinkela_wire_1644),
        .dout(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(new_Jinkela_wire_1635),
        .dout(new_Jinkela_wire_1636)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_1645),
        .dout(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(new_Jinkela_wire_1636),
        .dout(new_Jinkela_wire_1637)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_1637),
        .dout(new_Jinkela_wire_1638)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_1647),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(_0274_),
        .dout(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_1656),
        .dout(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_1668),
        .dout(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(_0258_),
        .dout(new_Jinkela_wire_1675)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(_0128_),
        .dout(new_Jinkela_wire_1676)
    );

    spl2 new_Jinkela_splitter_155 (
        .a(new_net_15),
        .c(new_Jinkela_wire_1681),
        .b(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(new_Jinkela_wire_1670),
        .dout(new_Jinkela_wire_1671)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_1671),
        .dout(new_Jinkela_wire_1672)
    );

    spl3L new_Jinkela_splitter_156 (
        .a(_0237_),
        .c(new_Jinkela_wire_1690),
        .b(new_Jinkela_wire_1691),
        .d(new_Jinkela_wire_1692)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_1676),
        .dout(new_Jinkela_wire_1677)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_1672),
        .dout(new_Jinkela_wire_1673)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_1677),
        .dout(new_Jinkela_wire_1678)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_1682),
        .dout(new_Jinkela_wire_1683)
    );

    spl2 new_Jinkela_splitter_158 (
        .a(_0254_),
        .c(new_Jinkela_wire_1697),
        .b(new_Jinkela_wire_1698)
    );

    spl2 new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_1678),
        .c(new_Jinkela_wire_1679),
        .b(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(new_Jinkela_wire_1683),
        .dout(new_Jinkela_wire_1684)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_1692),
        .dout(new_Jinkela_wire_1693)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(_0190_),
        .dout(new_Jinkela_wire_1699)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(_0153_),
        .c(new_Jinkela_wire_1704),
        .b(new_Jinkela_wire_1705)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_1684),
        .dout(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_1693),
        .dout(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(new_Jinkela_wire_1686),
        .dout(new_Jinkela_wire_1687)
    );

    spl2 new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_1699),
        .c(new_Jinkela_wire_1700),
        .b(new_Jinkela_wire_1701)
    );

    spl2 new_Jinkela_splitter_160 (
        .a(_0193_),
        .c(new_Jinkela_wire_1702),
        .b(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_1687),
        .dout(new_Jinkela_wire_1688)
    );

    spl2 new_Jinkela_splitter_157 (
        .a(new_Jinkela_wire_1694),
        .c(new_Jinkela_wire_1695),
        .b(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_1688),
        .dout(new_Jinkela_wire_1689)
    );

    spl2 new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_840),
        .c(new_Jinkela_wire_841),
        .b(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    or_bb _0570_ (
        .a(_0062_),
        .b(_0061_),
        .c(_0063_)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1241),
        .dout(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1219),
        .dout(new_Jinkela_wire_1220)
    );

    or_bb _0571_ (
        .a(_0063_),
        .b(new_Jinkela_wire_2219),
        .c(new_net_9)
    );

    bfr new_Jinkela_buffer_305 (
        .din(G52),
        .dout(new_Jinkela_wire_426)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    and_bi _0572_ (
        .a(new_Jinkela_wire_624),
        .b(new_Jinkela_wire_763),
        .c(_0064_)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_819),
        .c(new_Jinkela_wire_820),
        .e(new_Jinkela_wire_821),
        .b(new_Jinkela_wire_822),
        .d(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1258),
        .dout(new_Jinkela_wire_1259)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    and_bi _0573_ (
        .a(new_Jinkela_wire_619),
        .b(new_Jinkela_wire_883),
        .c(_0065_)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_390),
        .dout(new_Jinkela_wire_391)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    or_bb _0574_ (
        .a(_0065_),
        .b(new_Jinkela_wire_316),
        .c(_0066_)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1242),
        .dout(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    and_bi _0575_ (
        .a(new_Jinkela_wire_1443),
        .b(_0066_),
        .c(_0067_)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_424),
        .dout(new_Jinkela_wire_425)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    and_bi _0576_ (
        .a(new_Jinkela_wire_897),
        .b(new_Jinkela_wire_1664),
        .c(_0068_)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1255),
        .dout(new_Jinkela_wire_1256)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1222),
        .dout(new_Jinkela_wire_1223)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    and_bi _0577_ (
        .a(new_Jinkela_wire_604),
        .b(new_Jinkela_wire_2705),
        .c(_0069_)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    or_bb _0578_ (
        .a(_0069_),
        .b(_0068_),
        .c(_0070_)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1243),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1223),
        .dout(new_Jinkela_wire_1224)
    );

    and_bi _0579_ (
        .a(new_Jinkela_wire_2266),
        .b(_0070_),
        .c(new_net_7)
    );

    bfr new_Jinkela_buffer_311 (
        .din(G8),
        .dout(new_Jinkela_wire_432)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    and_bi _0580_ (
        .a(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_557),
        .c(_0071_)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1260),
        .dout(new_Jinkela_wire_1261)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1224),
        .dout(new_Jinkela_wire_1225)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    and_bi _0581_ (
        .a(new_Jinkela_wire_1),
        .b(new_Jinkela_wire_556),
        .c(_0072_)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_370),
        .dout(new_Jinkela_wire_371)
    );

    and_bi _0582_ (
        .a(_0071_),
        .b(_0072_),
        .c(_0073_)
    );

    bfr new_Jinkela_buffer_678 (
        .din(G9),
        .dout(new_Jinkela_wire_884)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1225),
        .dout(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_322 (
        .din(G98),
        .dout(new_Jinkela_wire_448)
    );

    and_bi _0583_ (
        .a(new_Jinkela_wire_1144),
        .b(new_Jinkela_wire_1278),
        .c(_0074_)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_426),
        .dout(new_Jinkela_wire_427)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(G149),
        .c(new_Jinkela_wire_887),
        .b(new_Jinkela_wire_888)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    and_bi _0584_ (
        .a(new_Jinkela_wire_1145),
        .b(new_Jinkela_wire_1279),
        .c(_0075_)
    );

    bfr new_Jinkela_buffer_988 (
        .din(G102),
        .dout(new_Jinkela_wire_1274)
    );

    spl3L new_Jinkela_splitter_72 (
        .a(G121),
        .c(new_Jinkela_wire_889),
        .b(new_Jinkela_wire_890),
        .d(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1226),
        .dout(new_Jinkela_wire_1227)
    );

    and_bi _0585_ (
        .a(_0074_),
        .b(_0075_),
        .c(_0076_)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    and_bi _0586_ (
        .a(new_Jinkela_wire_1730),
        .b(new_Jinkela_wire_2019),
        .c(_0077_)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1227),
        .dout(new_Jinkela_wire_1228)
    );

    and_bi _0587_ (
        .a(new_Jinkela_wire_1731),
        .b(new_Jinkela_wire_2020),
        .c(_0078_)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    and_bi _0588_ (
        .a(_0077_),
        .b(_0078_),
        .c(_0079_)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1261),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_687 (
        .din(G78),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_399),
        .dout(new_Jinkela_wire_400)
    );

    and_bi _0589_ (
        .a(new_Jinkela_wire_1173),
        .b(new_Jinkela_wire_902),
        .c(_0080_)
    );

    spl3L new_Jinkela_splitter_101 (
        .a(new_Jinkela_wire_1246),
        .c(new_Jinkela_wire_1247),
        .b(new_Jinkela_wire_1248),
        .d(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    and_bi _0590_ (
        .a(new_Jinkela_wire_1174),
        .b(new_Jinkela_wire_903),
        .c(_0081_)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1266),
        .dout(new_Jinkela_wire_1267)
    );

    and_bi _0591_ (
        .a(_0080_),
        .b(_0081_),
        .c(_0082_)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_427),
        .dout(new_Jinkela_wire_428)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    and_bi _0592_ (
        .a(new_Jinkela_wire_1355),
        .b(new_Jinkela_wire_1709),
        .c(_0083_)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_400),
        .dout(new_Jinkela_wire_401)
    );

    and_bi _0593_ (
        .a(new_Jinkela_wire_1356),
        .b(new_Jinkela_wire_1710),
        .c(_0084_)
    );

    spl3L new_Jinkela_splitter_102 (
        .a(G128),
        .c(new_Jinkela_wire_1278),
        .b(new_Jinkela_wire_1279),
        .d(new_Jinkela_wire_1280)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_871),
        .dout(new_Jinkela_wire_872)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    spl2 new_Jinkela_splitter_104 (
        .a(G151),
        .c(new_Jinkela_wire_1295),
        .b(new_Jinkela_wire_1296)
    );

    and_bi _0594_ (
        .a(_0083_),
        .b(_0084_),
        .c(_0085_)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    and_bi _0595_ (
        .a(new_Jinkela_wire_1056),
        .b(new_Jinkela_wire_1232),
        .c(_0086_)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_432),
        .dout(new_Jinkela_wire_433)
    );

    bfr new_Jinkela_buffer_681 (
        .din(G48),
        .dout(new_Jinkela_wire_892)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1267),
        .dout(new_Jinkela_wire_1268)
    );

    and_bi _0596_ (
        .a(new_Jinkela_wire_1057),
        .b(new_Jinkela_wire_1233),
        .c(_0087_)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1264),
        .dout(new_Jinkela_wire_1265)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    and_bi _0597_ (
        .a(_0086_),
        .b(_0087_),
        .c(_0088_)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    spl3L new_Jinkela_splitter_73 (
        .a(G136),
        .c(new_Jinkela_wire_902),
        .b(new_Jinkela_wire_903),
        .d(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1274),
        .dout(new_Jinkela_wire_1275)
    );

    and_bi _0598_ (
        .a(new_Jinkela_wire_212),
        .b(new_Jinkela_wire_825),
        .c(_0089_)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1268),
        .dout(new_Jinkela_wire_1269)
    );

    and_bi _0599_ (
        .a(new_Jinkela_wire_211),
        .b(new_Jinkela_wire_824),
        .c(_0090_)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(G21),
        .dout(new_Jinkela_wire_1297)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_403),
        .dout(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1280),
        .dout(new_Jinkela_wire_1281)
    );

    and_bi _0600_ (
        .a(_0089_),
        .b(_0090_),
        .c(_0091_)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1269),
        .dout(new_Jinkela_wire_1270)
    );

    spl2 new_Jinkela_splitter_76 (
        .a(G43),
        .c(new_Jinkela_wire_921),
        .b(new_Jinkela_wire_922)
    );

    and_bi _0601_ (
        .a(new_Jinkela_wire_2491),
        .b(new_Jinkela_wire_1737),
        .c(_0092_)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_404),
        .dout(new_Jinkela_wire_405)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1275),
        .dout(new_Jinkela_wire_1276)
    );

    and_bi _0602_ (
        .a(new_Jinkela_wire_2492),
        .b(new_Jinkela_wire_1738),
        .c(_0093_)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1270),
        .dout(new_Jinkela_wire_1271)
    );

    and_bi _0603_ (
        .a(_0092_),
        .b(_0093_),
        .c(_0094_)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_433),
        .dout(new_Jinkela_wire_434)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(new_Jinkela_wire_876),
        .c(new_Jinkela_wire_877),
        .b(new_Jinkela_wire_878)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_405),
        .dout(new_Jinkela_wire_406)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(G88),
        .dout(new_Jinkela_wire_1299)
    );

    and_bi _0604_ (
        .a(new_Jinkela_wire_1447),
        .b(new_Jinkela_wire_1735),
        .c(_0095_)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1271),
        .dout(new_Jinkela_wire_1272)
    );

    spl2 new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_878),
        .c(new_Jinkela_wire_879),
        .b(new_Jinkela_wire_880)
    );

    and_bi _0605_ (
        .a(new_Jinkela_wire_1448),
        .b(new_Jinkela_wire_1736),
        .c(_0096_)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_430),
        .dout(new_Jinkela_wire_431)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1276),
        .dout(new_Jinkela_wire_1277)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_406),
        .dout(new_Jinkela_wire_407)
    );

    or_bb _0606_ (
        .a(_0096_),
        .b(_0095_),
        .c(new_net_13)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1272),
        .dout(new_Jinkela_wire_1273)
    );

    or_bb _0607_ (
        .a(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_89),
        .c(_0097_)
    );

    spl2 new_Jinkela_splitter_43 (
        .a(G32),
        .c(new_Jinkela_wire_454),
        .b(new_Jinkela_wire_455)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1282),
        .dout(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_407),
        .dout(new_Jinkela_wire_408)
    );

    and_bi _0608_ (
        .a(new_Jinkela_wire_90),
        .b(new_Jinkela_wire_180),
        .c(_0098_)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_1435),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_356 (
        .din(G66),
        .dout(new_Jinkela_wire_484)
    );

    and_bi _0609_ (
        .a(new_Jinkela_wire_2057),
        .b(new_Jinkela_wire_2553),
        .c(_0099_)
    );

    bfr new_Jinkela_buffer_326 (
        .din(G11),
        .dout(new_Jinkela_wire_452)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    and_bi _0545_ (
        .a(new_Jinkela_wire_36),
        .b(new_Jinkela_wire_2710),
        .c(_0041_)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1281),
        .dout(new_Jinkela_wire_1282)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    or_bb _0610_ (
        .a(new_Jinkela_wire_957),
        .b(new_Jinkela_wire_1111),
        .c(_0100_)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1297),
        .dout(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_434),
        .dout(new_Jinkela_wire_435)
    );

    and_bi _0611_ (
        .a(new_Jinkela_wire_1110),
        .b(new_Jinkela_wire_956),
        .c(_0101_)
    );

    and_bi _0524_ (
        .a(new_Jinkela_wire_632),
        .b(new_Jinkela_wire_1231),
        .c(_0022_)
    );

    and_bi _0502_ (
        .a(new_Jinkela_wire_782),
        .b(new_Jinkela_wire_1845),
        .c(_0003_)
    );

    or_bb _0500_ (
        .a(new_Jinkela_wire_1977),
        .b(new_Jinkela_wire_578),
        .c(_0001_)
    );

    or_bb _0501_ (
        .a(new_Jinkela_wire_503),
        .b(new_Jinkela_wire_235),
        .c(_0002_)
    );

    or_bb _0499_ (
        .a(new_Jinkela_wire_501),
        .b(new_Jinkela_wire_232),
        .c(_0000_)
    );

    and_bi _0503_ (
        .a(_0001_),
        .b(_0003_),
        .c(_0004_)
    );

    and_bi _0507_ (
        .a(new_Jinkela_wire_309),
        .b(new_Jinkela_wire_2506),
        .c(_0008_)
    );

    or_bb _0506_ (
        .a(new_Jinkela_wire_504),
        .b(new_Jinkela_wire_233),
        .c(_0007_)
    );

    or_bb _0504_ (
        .a(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_234),
        .c(_0005_)
    );

    and_bi _0516_ (
        .a(_0012_),
        .b(_0015_),
        .c(new_net_0)
    );

    and_bi _0505_ (
        .a(new_Jinkela_wire_862),
        .b(new_Jinkela_wire_1934),
        .c(_0006_)
    );

    or_bb _0508_ (
        .a(_0008_),
        .b(_0006_),
        .c(_0009_)
    );

    and_bi _0509_ (
        .a(_0004_),
        .b(_0009_),
        .c(new_net_2)
    );

    or_bb _0510_ (
        .a(new_Jinkela_wire_2505),
        .b(new_Jinkela_wire_521),
        .c(_0010_)
    );

    and_bi _0511_ (
        .a(new_Jinkela_wire_451),
        .b(new_Jinkela_wire_1936),
        .c(_0011_)
    );

    and_bi _0512_ (
        .a(_0010_),
        .b(_0011_),
        .c(_0012_)
    );

    and_bi _0513_ (
        .a(new_Jinkela_wire_1302),
        .b(new_Jinkela_wire_1850),
        .c(_0013_)
    );

    and_bi _0514_ (
        .a(new_Jinkela_wire_901),
        .b(new_Jinkela_wire_1982),
        .c(_0014_)
    );

    or_bb _0515_ (
        .a(_0014_),
        .b(_0013_),
        .c(_0015_)
    );

    and_bi _0517_ (
        .a(new_Jinkela_wire_1140),
        .b(new_Jinkela_wire_2509),
        .c(_0016_)
    );

    and_bi _0518_ (
        .a(new_Jinkela_wire_615),
        .b(new_Jinkela_wire_1980),
        .c(_0017_)
    );

    or_bb _0519_ (
        .a(_0017_),
        .b(_0016_),
        .c(_0018_)
    );

    and_bi _0520_ (
        .a(new_Jinkela_wire_976),
        .b(new_Jinkela_wire_1852),
        .c(_0019_)
    );

    and_bi _0521_ (
        .a(new_Jinkela_wire_991),
        .b(new_Jinkela_wire_1935),
        .c(_0020_)
    );

    or_bb _0522_ (
        .a(_0020_),
        .b(_0019_),
        .c(_0021_)
    );

    or_bb _0523_ (
        .a(_0021_),
        .b(_0018_),
        .c(new_net_1)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(new_Jinkela_wire_2025),
        .dout(new_Jinkela_wire_2026)
    );

    bfr new_Jinkela_buffer_1715 (
        .din(new_Jinkela_wire_2311),
        .dout(new_Jinkela_wire_2312)
    );

    bfr new_Jinkela_buffer_1697 (
        .din(new_Jinkela_wire_2291),
        .dout(new_Jinkela_wire_2292)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_2065),
        .dout(new_Jinkela_wire_2066)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(_0316_),
        .dout(new_Jinkela_wire_2085)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_1721 (
        .din(new_Jinkela_wire_2317),
        .dout(new_Jinkela_wire_2318)
    );

    bfr new_Jinkela_buffer_1698 (
        .din(new_Jinkela_wire_2292),
        .dout(new_Jinkela_wire_2293)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_2050),
        .dout(new_Jinkela_wire_2051)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_2027),
        .dout(new_Jinkela_wire_2028)
    );

    bfr new_Jinkela_buffer_1745 (
        .din(new_Jinkela_wire_2343),
        .dout(new_Jinkela_wire_2344)
    );

    bfr new_Jinkela_buffer_1716 (
        .din(new_Jinkela_wire_2312),
        .dout(new_Jinkela_wire_2313)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(new_Jinkela_wire_2028),
        .dout(new_Jinkela_wire_2029)
    );

    bfr new_Jinkela_buffer_1722 (
        .din(new_Jinkela_wire_2318),
        .dout(new_Jinkela_wire_2319)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_2051),
        .dout(new_Jinkela_wire_2052)
    );

    bfr new_Jinkela_buffer_1717 (
        .din(new_Jinkela_wire_2313),
        .dout(new_Jinkela_wire_2314)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(new_Jinkela_wire_2029),
        .dout(new_Jinkela_wire_2030)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_2059),
        .dout(new_Jinkela_wire_2060)
    );

    bfr new_Jinkela_buffer_1718 (
        .din(new_Jinkela_wire_2314),
        .dout(new_Jinkela_wire_2315)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(new_Jinkela_wire_2030),
        .dout(new_Jinkela_wire_2031)
    );

    bfr new_Jinkela_buffer_1723 (
        .din(new_Jinkela_wire_2319),
        .dout(new_Jinkela_wire_2320)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(new_Jinkela_wire_2052),
        .dout(new_Jinkela_wire_2053)
    );

    bfr new_Jinkela_buffer_1719 (
        .din(new_Jinkela_wire_2315),
        .dout(new_Jinkela_wire_2316)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_2031),
        .dout(new_Jinkela_wire_2032)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(_0343_),
        .dout(new_Jinkela_wire_2087)
    );

    bfr new_Jinkela_buffer_1724 (
        .din(new_Jinkela_wire_2320),
        .dout(new_Jinkela_wire_2321)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(new_Jinkela_wire_2032),
        .dout(new_Jinkela_wire_2033)
    );

    bfr new_Jinkela_buffer_1779 (
        .din(_0244_),
        .dout(new_Jinkela_wire_2387)
    );

    bfr new_Jinkela_buffer_1746 (
        .din(new_Jinkela_wire_2344),
        .dout(new_Jinkela_wire_2345)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(new_Jinkela_wire_2053),
        .dout(new_Jinkela_wire_2054)
    );

    bfr new_Jinkela_buffer_1725 (
        .din(new_Jinkela_wire_2321),
        .dout(new_Jinkela_wire_2322)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(new_Jinkela_wire_2033),
        .dout(new_Jinkela_wire_2034)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(_0289_),
        .c(new_Jinkela_wire_2384),
        .b(new_Jinkela_wire_2385)
    );

    spl4L new_Jinkela_splitter_209 (
        .a(new_Jinkela_wire_2061),
        .c(new_Jinkela_wire_2062),
        .e(new_Jinkela_wire_2063),
        .b(new_Jinkela_wire_2064),
        .d(new_Jinkela_wire_2065)
    );

    bfr new_Jinkela_buffer_1726 (
        .din(new_Jinkela_wire_2322),
        .dout(new_Jinkela_wire_2323)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(new_Jinkela_wire_2034),
        .dout(new_Jinkela_wire_2035)
    );

    spl3L new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_2361),
        .c(new_Jinkela_wire_2362),
        .b(new_Jinkela_wire_2363),
        .d(new_Jinkela_wire_2364)
    );

    bfr new_Jinkela_buffer_1747 (
        .din(new_Jinkela_wire_2345),
        .dout(new_Jinkela_wire_2346)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_2054),
        .dout(new_Jinkela_wire_2055)
    );

    bfr new_Jinkela_buffer_1727 (
        .din(new_Jinkela_wire_2323),
        .dout(new_Jinkela_wire_2324)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(new_Jinkela_wire_2035),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_1778 (
        .din(_0376_),
        .dout(new_Jinkela_wire_2386)
    );

    bfr new_Jinkela_buffer_1728 (
        .din(new_Jinkela_wire_2324),
        .dout(new_Jinkela_wire_2325)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_2036),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1761 (
        .din(new_Jinkela_wire_2364),
        .dout(new_Jinkela_wire_2365)
    );

    bfr new_Jinkela_buffer_1748 (
        .din(new_Jinkela_wire_2346),
        .dout(new_Jinkela_wire_2347)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_2055),
        .dout(new_Jinkela_wire_2056)
    );

    bfr new_Jinkela_buffer_1729 (
        .din(new_Jinkela_wire_2325),
        .dout(new_Jinkela_wire_2326)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(_0099_),
        .c(new_Jinkela_wire_2389),
        .b(new_Jinkela_wire_2390)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(_0297_),
        .dout(new_Jinkela_wire_2094)
    );

    bfr new_Jinkela_buffer_1730 (
        .din(new_Jinkela_wire_2326),
        .dout(new_Jinkela_wire_2327)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1781 (
        .din(_0418_),
        .dout(new_Jinkela_wire_2391)
    );

    bfr new_Jinkela_buffer_1749 (
        .din(new_Jinkela_wire_2347),
        .dout(new_Jinkela_wire_2348)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(new_Jinkela_wire_2087),
        .dout(new_Jinkela_wire_2088)
    );

    bfr new_Jinkela_buffer_1731 (
        .din(new_Jinkela_wire_2327),
        .dout(new_Jinkela_wire_2328)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_2066),
        .dout(new_Jinkela_wire_2067)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1780 (
        .din(new_Jinkela_wire_2387),
        .dout(new_Jinkela_wire_2388)
    );

    bfr new_Jinkela_buffer_1732 (
        .din(new_Jinkela_wire_2328),
        .dout(new_Jinkela_wire_2329)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1750 (
        .din(new_Jinkela_wire_2348),
        .dout(new_Jinkela_wire_2349)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_net_948),
        .dout(new_Jinkela_wire_2102)
    );

    bfr new_Jinkela_buffer_1733 (
        .din(new_Jinkela_wire_2329),
        .dout(new_Jinkela_wire_2330)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_2067),
        .dout(new_Jinkela_wire_2068)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(new_Jinkela_wire_2041),
        .dout(new_Jinkela_wire_2042)
    );

    bfr new_Jinkela_buffer_1734 (
        .din(new_Jinkela_wire_2330),
        .dout(new_Jinkela_wire_2331)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(new_Jinkela_wire_2042),
        .dout(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_1762 (
        .din(new_Jinkela_wire_2365),
        .dout(new_Jinkela_wire_2366)
    );

    bfr new_Jinkela_buffer_1751 (
        .din(new_Jinkela_wire_2349),
        .dout(new_Jinkela_wire_2350)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(new_Jinkela_wire_2088),
        .dout(new_Jinkela_wire_2089)
    );

    bfr new_Jinkela_buffer_1735 (
        .din(new_Jinkela_wire_2331),
        .dout(new_Jinkela_wire_2332)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_2068),
        .dout(new_Jinkela_wire_2069)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    bfr new_Jinkela_buffer_1736 (
        .din(new_Jinkela_wire_2332),
        .dout(new_Jinkela_wire_2333)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(_0495_),
        .dout(new_Jinkela_wire_2086)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_2044),
        .dout(new_Jinkela_wire_2045)
    );

    bfr new_Jinkela_buffer_1752 (
        .din(new_Jinkela_wire_2350),
        .dout(new_Jinkela_wire_2351)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_2094),
        .dout(new_Jinkela_wire_2095)
    );

    bfr new_Jinkela_buffer_1737 (
        .din(new_Jinkela_wire_2333),
        .dout(new_Jinkela_wire_2334)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_2069),
        .dout(new_Jinkela_wire_2070)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_1738 (
        .din(new_Jinkela_wire_2334),
        .dout(new_Jinkela_wire_2335)
    );

    and_bi _0948_ (
        .a(new_Jinkela_wire_1072),
        .b(new_Jinkela_wire_1745),
        .c(_0419_)
    );

    and_bi _0949_ (
        .a(new_Jinkela_wire_972),
        .b(new_Jinkela_wire_1353),
        .c(_0420_)
    );

    and_bi _0950_ (
        .a(_0419_),
        .b(_0420_),
        .c(_0421_)
    );

    and_bi _0951_ (
        .a(new_Jinkela_wire_1875),
        .b(new_Jinkela_wire_1605),
        .c(_0422_)
    );

    or_bb _0952_ (
        .a(new_Jinkela_wire_1742),
        .b(new_Jinkela_wire_1292),
        .c(_0423_)
    );

    and_bi _0953_ (
        .a(new_Jinkela_wire_1126),
        .b(new_Jinkela_wire_1348),
        .c(_0424_)
    );

    and_bi _0954_ (
        .a(_0423_),
        .b(_0424_),
        .c(_0425_)
    );

    or_bb _0955_ (
        .a(new_Jinkela_wire_2546),
        .b(new_Jinkela_wire_1530),
        .c(_0426_)
    );

    or_bb _0956_ (
        .a(new_Jinkela_wire_1744),
        .b(new_Jinkela_wire_877),
        .c(_0427_)
    );

    and_bi _0957_ (
        .a(new_Jinkela_wire_1172),
        .b(new_Jinkela_wire_1350),
        .c(_0428_)
    );

    and_bi _0958_ (
        .a(_0427_),
        .b(_0428_),
        .c(_0429_)
    );

    and_bi _0959_ (
        .a(new_Jinkela_wire_2185),
        .b(new_Jinkela_wire_1512),
        .c(_0430_)
    );

    or_bb _0960_ (
        .a(new_Jinkela_wire_1740),
        .b(new_Jinkela_wire_1099),
        .c(_0431_)
    );

    and_bi _0961_ (
        .a(new_Jinkela_wire_920),
        .b(new_Jinkela_wire_1351),
        .c(_0432_)
    );

    and_bi _0962_ (
        .a(_0431_),
        .b(_0432_),
        .c(_0433_)
    );

    or_bb _0963_ (
        .a(_0433_),
        .b(new_Jinkela_wire_1729),
        .c(_0434_)
    );

    or_bb _0964_ (
        .a(new_Jinkela_wire_1840),
        .b(_0430_),
        .c(_0435_)
    );

    and_bi _0965_ (
        .a(new_Jinkela_wire_1513),
        .b(new_Jinkela_wire_2186),
        .c(_0436_)
    );

    and_bi _0966_ (
        .a(new_Jinkela_wire_1529),
        .b(new_Jinkela_wire_2547),
        .c(_0437_)
    );

    or_bb _0967_ (
        .a(_0437_),
        .b(_0436_),
        .c(_0438_)
    );

    and_bi _0968_ (
        .a(_0435_),
        .b(_0438_),
        .c(_0439_)
    );

    and_bi _0969_ (
        .a(new_Jinkela_wire_2562),
        .b(_0439_),
        .c(_0440_)
    );

    or_bb _0970_ (
        .a(_0440_),
        .b(new_Jinkela_wire_1581),
        .c(_0441_)
    );

    and_bi _0971_ (
        .a(new_Jinkela_wire_1874),
        .b(new_Jinkela_wire_1606),
        .c(_0442_)
    );

    and_bi _0972_ (
        .a(new_Jinkela_wire_442),
        .b(new_Jinkela_wire_2462),
        .c(_0443_)
    );

    and_bi _0973_ (
        .a(new_Jinkela_wire_1250),
        .b(new_Jinkela_wire_2146),
        .c(_0444_)
    );

    and_bi _0974_ (
        .a(new_Jinkela_wire_107),
        .b(new_Jinkela_wire_1748),
        .c(_0445_)
    );

    and_bi _0975_ (
        .a(_0444_),
        .b(_0445_),
        .c(_0446_)
    );

    and_bi _0976_ (
        .a(new_Jinkela_wire_2124),
        .b(new_Jinkela_wire_1922),
        .c(_0447_)
    );

    or_bb _0977_ (
        .a(_0447_),
        .b(new_Jinkela_wire_2148),
        .c(_0448_)
    );

    and_bi _0978_ (
        .a(_0441_),
        .b(new_Jinkela_wire_2565),
        .c(_0449_)
    );

    and_bi _0979_ (
        .a(new_Jinkela_wire_2125),
        .b(new_Jinkela_wire_1923),
        .c(_0450_)
    );

    and_bi _0980_ (
        .a(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_2064),
        .c(_0451_)
    );

    and_bi _0981_ (
        .a(new_Jinkela_wire_18),
        .b(new_Jinkela_wire_2145),
        .c(_0452_)
    );

    and_bi _0982_ (
        .a(new_Jinkela_wire_197),
        .b(new_Jinkela_wire_1747),
        .c(_0453_)
    );

    and_bi _0983_ (
        .a(_0452_),
        .b(_0453_),
        .c(_0454_)
    );

    and_bi _0984_ (
        .a(new_Jinkela_wire_2306),
        .b(new_Jinkela_wire_1566),
        .c(_0455_)
    );

    or_bb _0985_ (
        .a(_0455_),
        .b(_0450_),
        .c(_0456_)
    );

    or_bb _0986_ (
        .a(new_Jinkela_wire_1716),
        .b(_0449_),
        .c(_0457_)
    );

    and_bi _0987_ (
        .a(new_Jinkela_wire_1824),
        .b(new_Jinkela_wire_1749),
        .c(_0458_)
    );

    and_bi _0988_ (
        .a(new_Jinkela_wire_2307),
        .b(new_Jinkela_wire_1567),
        .c(_0459_)
    );

    or_bb _0989_ (
        .a(_0459_),
        .b(new_Jinkela_wire_1332),
        .c(_0460_)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_409),
        .dout(new_Jinkela_wire_410)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(G29),
        .dout(new_Jinkela_wire_1303)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(_0466_),
        .dout(new_Jinkela_wire_1325)
    );

    bfr new_Jinkela_buffer_1941 (
        .din(_0486_),
        .dout(new_Jinkela_wire_2636)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_1914 (
        .din(new_Jinkela_wire_2594),
        .dout(new_Jinkela_wire_2595)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1299),
        .dout(new_Jinkela_wire_1300)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1284),
        .dout(new_Jinkela_wire_1285)
    );

    bfr new_Jinkela_buffer_1931 (
        .din(new_Jinkela_wire_2621),
        .dout(new_Jinkela_wire_2622)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1283),
        .dout(new_Jinkela_wire_1284)
    );

    bfr new_Jinkela_buffer_1915 (
        .din(new_Jinkela_wire_2595),
        .dout(new_Jinkela_wire_2596)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_411),
        .dout(new_Jinkela_wire_412)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1307),
        .dout(new_Jinkela_wire_1308)
    );

    bfr new_Jinkela_buffer_1933 (
        .din(new_Jinkela_wire_2625),
        .dout(new_Jinkela_wire_2626)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1285),
        .dout(new_Jinkela_wire_1286)
    );

    bfr new_Jinkela_buffer_1916 (
        .din(new_Jinkela_wire_2596),
        .dout(new_Jinkela_wire_2597)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_412),
        .dout(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(new_Jinkela_wire_1300),
        .dout(new_Jinkela_wire_1301)
    );

    spl2 new_Jinkela_splitter_268 (
        .a(_0215_),
        .c(new_Jinkela_wire_2634),
        .b(new_Jinkela_wire_2635)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_436),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1286),
        .dout(new_Jinkela_wire_1287)
    );

    bfr new_Jinkela_buffer_1917 (
        .din(new_Jinkela_wire_2597),
        .dout(new_Jinkela_wire_2598)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_413),
        .dout(new_Jinkela_wire_414)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(_0478_),
        .dout(new_Jinkela_wire_1329)
    );

    spl3L new_Jinkela_splitter_271 (
        .a(new_net_10),
        .c(new_Jinkela_wire_2671),
        .b(new_Jinkela_wire_2672),
        .d(new_Jinkela_wire_2673)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1303),
        .dout(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_1942 (
        .din(new_Jinkela_wire_2636),
        .dout(new_Jinkela_wire_2637)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1287),
        .dout(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_1918 (
        .din(new_Jinkela_wire_2598),
        .dout(new_Jinkela_wire_2599)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1301),
        .dout(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_1934 (
        .din(new_Jinkela_wire_2626),
        .dout(new_Jinkela_wire_2627)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_437),
        .dout(new_Jinkela_wire_438)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1288),
        .dout(new_Jinkela_wire_1289)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    bfr new_Jinkela_buffer_1935 (
        .din(new_Jinkela_wire_2627),
        .dout(new_Jinkela_wire_2628)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1289),
        .dout(new_Jinkela_wire_1290)
    );

    spl3L new_Jinkela_splitter_269 (
        .a(new_net_2),
        .c(new_Jinkela_wire_2645),
        .b(new_Jinkela_wire_2646),
        .d(new_Jinkela_wire_2647)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_416),
        .dout(new_Jinkela_wire_417)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1325),
        .dout(new_Jinkela_wire_1326)
    );

    bfr new_Jinkela_buffer_1936 (
        .din(new_Jinkela_wire_2628),
        .dout(new_Jinkela_wire_2629)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1304),
        .dout(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_438),
        .dout(new_Jinkela_wire_439)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1290),
        .dout(new_Jinkela_wire_1291)
    );

    bfr new_Jinkela_buffer_1996 (
        .din(_0057_),
        .dout(new_Jinkela_wire_2700)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_417),
        .dout(new_Jinkela_wire_418)
    );

    spl3L new_Jinkela_splitter_270 (
        .a(new_Jinkela_wire_2647),
        .c(new_Jinkela_wire_2648),
        .b(new_Jinkela_wire_2649),
        .d(new_Jinkela_wire_2650)
    );

    bfr new_Jinkela_buffer_1937 (
        .din(new_Jinkela_wire_2629),
        .dout(new_Jinkela_wire_2630)
    );

    spl3L new_Jinkela_splitter_103 (
        .a(new_Jinkela_wire_1291),
        .c(new_Jinkela_wire_1292),
        .b(new_Jinkela_wire_1293),
        .d(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_1943 (
        .din(new_Jinkela_wire_2637),
        .dout(new_Jinkela_wire_2638)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_418),
        .dout(new_Jinkela_wire_419)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(_0458_),
        .dout(new_Jinkela_wire_1330)
    );

    bfr new_Jinkela_buffer_1938 (
        .din(new_Jinkela_wire_2630),
        .dout(new_Jinkela_wire_2631)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1305),
        .dout(new_Jinkela_wire_1306)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_419),
        .dout(new_Jinkela_wire_420)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1326),
        .dout(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_1939 (
        .din(new_Jinkela_wire_2631),
        .dout(new_Jinkela_wire_2632)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1306),
        .dout(new_Jinkela_wire_1307)
    );

    bfr new_Jinkela_buffer_359 (
        .din(G14),
        .dout(new_Jinkela_wire_487)
    );

    bfr new_Jinkela_buffer_1944 (
        .din(new_Jinkela_wire_2638),
        .dout(new_Jinkela_wire_2639)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_420),
        .dout(new_Jinkela_wire_421)
    );

    spl2 new_Jinkela_splitter_106 (
        .a(_0137_),
        .c(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1334)
    );

    bfr new_Jinkela_buffer_1940 (
        .din(new_Jinkela_wire_2632),
        .dout(new_Jinkela_wire_2633)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_421),
        .dout(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(_0322_),
        .dout(new_Jinkela_wire_1335)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1327),
        .dout(new_Jinkela_wire_1328)
    );

    bfr new_Jinkela_buffer_1945 (
        .din(new_Jinkela_wire_2639),
        .dout(new_Jinkela_wire_2640)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1308),
        .dout(new_Jinkela_wire_1309)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_484),
        .dout(new_Jinkela_wire_485)
    );

    bfr new_Jinkela_buffer_1970 (
        .din(new_Jinkela_wire_2673),
        .dout(new_Jinkela_wire_2674)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_422),
        .dout(new_Jinkela_wire_423)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1330),
        .dout(new_Jinkela_wire_1331)
    );

    bfr new_Jinkela_buffer_1946 (
        .din(new_Jinkela_wire_2640),
        .dout(new_Jinkela_wire_2641)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1309),
        .dout(new_Jinkela_wire_1310)
    );

    spl3L new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_441),
        .c(new_Jinkela_wire_442),
        .b(new_Jinkela_wire_443),
        .d(new_Jinkela_wire_444)
    );

    bfr new_Jinkela_buffer_1950 (
        .din(new_Jinkela_wire_2650),
        .dout(new_Jinkela_wire_2651)
    );

    bfr new_Jinkela_buffer_1947 (
        .din(new_Jinkela_wire_2641),
        .dout(new_Jinkela_wire_2642)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1310),
        .dout(new_Jinkela_wire_1311)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_444),
        .dout(new_Jinkela_wire_445)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1335),
        .dout(new_Jinkela_wire_1336)
    );

    bfr new_Jinkela_buffer_1971 (
        .din(new_Jinkela_wire_2674),
        .dout(new_Jinkela_wire_2675)
    );

    spl3L new_Jinkela_splitter_44 (
        .a(G143),
        .c(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_490),
        .d(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(new_Jinkela_wire_1331),
        .dout(new_Jinkela_wire_1332)
    );

    bfr new_Jinkela_buffer_1948 (
        .din(new_Jinkela_wire_2642),
        .dout(new_Jinkela_wire_2643)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_Jinkela_wire_1311),
        .dout(new_Jinkela_wire_1312)
    );

    spl2 new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_445),
        .c(new_Jinkela_wire_446),
        .b(new_Jinkela_wire_447)
    );

    bfr new_Jinkela_buffer_1951 (
        .din(new_Jinkela_wire_2651),
        .dout(new_Jinkela_wire_2652)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_485),
        .dout(new_Jinkela_wire_486)
    );

    bfr new_Jinkela_buffer_1949 (
        .din(new_Jinkela_wire_2643),
        .dout(new_Jinkela_wire_2644)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1312),
        .dout(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_1999 (
        .din(_0337_),
        .dout(new_Jinkela_wire_2716)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(G146),
        .c(new_Jinkela_wire_501),
        .e(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_503),
        .d(new_Jinkela_wire_504)
    );

    spl3L new_Jinkela_splitter_272 (
        .a(_0028_),
        .c(new_Jinkela_wire_2701),
        .b(new_Jinkela_wire_2704),
        .d(new_Jinkela_wire_2709)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(_0354_),
        .dout(new_Jinkela_wire_1341)
    );

    bfr new_Jinkela_buffer_1952 (
        .din(new_Jinkela_wire_2652),
        .dout(new_Jinkela_wire_2653)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1313),
        .dout(new_Jinkela_wire_1314)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(_0267_),
        .c(new_Jinkela_wire_1344),
        .b(new_Jinkela_wire_1345)
    );

    bfr new_Jinkela_buffer_1953 (
        .din(new_Jinkela_wire_2653),
        .dout(new_Jinkela_wire_2654)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1314),
        .dout(new_Jinkela_wire_1315)
    );

    bfr new_Jinkela_buffer_368 (
        .din(G28),
        .dout(new_Jinkela_wire_505)
    );

    spl4L new_Jinkela_splitter_274 (
        .a(new_Jinkela_wire_2704),
        .c(new_Jinkela_wire_2705),
        .e(new_Jinkela_wire_2706),
        .b(new_Jinkela_wire_2707),
        .d(new_Jinkela_wire_2708)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(_0482_),
        .dout(new_Jinkela_wire_1346)
    );

    bfr new_Jinkela_buffer_1972 (
        .din(new_Jinkela_wire_2675),
        .dout(new_Jinkela_wire_2676)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1336),
        .dout(new_Jinkela_wire_1337)
    );

    bfr new_Jinkela_buffer_1954 (
        .din(new_Jinkela_wire_2654),
        .dout(new_Jinkela_wire_2655)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1315),
        .dout(new_Jinkela_wire_1316)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    bfr new_Jinkela_buffer_1997 (
        .din(_0222_),
        .dout(new_Jinkela_wire_2714)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1341),
        .dout(new_Jinkela_wire_1342)
    );

    bfr new_Jinkela_buffer_1955 (
        .din(new_Jinkela_wire_2655),
        .dout(new_Jinkela_wire_2656)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1316),
        .dout(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_729 (
        .din(G7),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    spl3L new_Jinkela_splitter_77 (
        .a(G140),
        .c(new_Jinkela_wire_956),
        .b(new_Jinkela_wire_957),
        .d(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_730 (
        .din(G81),
        .dout(new_Jinkela_wire_952)
    );

    bfr new_Jinkela_buffer_745 (
        .din(G89),
        .dout(new_Jinkela_wire_973)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_952),
        .dout(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    spl3L new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_910),
        .c(new_Jinkela_wire_911),
        .b(new_Jinkela_wire_912),
        .d(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_953),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    spl3L new_Jinkela_splitter_75 (
        .a(new_Jinkela_wire_915),
        .c(new_Jinkela_wire_916),
        .b(new_Jinkela_wire_917),
        .d(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_749 (
        .din(G77),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_753 (
        .din(G95),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_960),
        .dout(new_Jinkela_wire_961)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_961),
        .dout(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    or_bb _0780_ (
        .a(new_Jinkela_wire_2671),
        .b(new_Jinkela_wire_74),
        .c(new_net_967)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(new_Jinkela_wire_1780),
        .dout(new_Jinkela_wire_1781)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(new_Jinkela_wire_2046),
        .dout(new_Jinkela_wire_2047)
    );

    or_bb _0546_ (
        .a(_0041_),
        .b(_0040_),
        .c(_0042_)
    );

    and_bi _0781_ (
        .a(new_Jinkela_wire_1199),
        .b(new_Jinkela_wire_276),
        .c(_0262_)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(new_Jinkela_wire_1761),
        .dout(new_Jinkela_wire_1762)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(new_Jinkela_wire_2089),
        .dout(new_Jinkela_wire_2090)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_2070),
        .dout(new_Jinkela_wire_2071)
    );

    or_bb _0782_ (
        .a(new_Jinkela_wire_998),
        .b(new_Jinkela_wire_921),
        .c(_0263_)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(new_net_6),
        .c(new_Jinkela_wire_1815),
        .b(new_Jinkela_wire_1816)
    );

    spl3L new_Jinkela_splitter_178 (
        .a(_0002_),
        .c(new_Jinkela_wire_1841),
        .b(new_Jinkela_wire_1843),
        .d(new_Jinkela_wire_1848)
    );

    and_bi _0783_ (
        .a(_0262_),
        .b(_0263_),
        .c(_0264_)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(new_Jinkela_wire_1762),
        .dout(new_Jinkela_wire_1763)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(_0443_),
        .dout(new_Jinkela_wire_2119)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_2071),
        .dout(new_Jinkela_wire_2072)
    );

    and_bi _0784_ (
        .a(new_Jinkela_wire_454),
        .b(new_Jinkela_wire_348),
        .c(_0265_)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(new_Jinkela_wire_1781),
        .dout(new_Jinkela_wire_1782)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(_0230_),
        .dout(new_Jinkela_wire_2126)
    );

    or_bb _0785_ (
        .a(new_Jinkela_wire_118),
        .b(new_Jinkela_wire_394),
        .c(_0266_)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_Jinkela_wire_1763),
        .dout(new_Jinkela_wire_1764)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_2090),
        .dout(new_Jinkela_wire_2091)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_2072),
        .dout(new_Jinkela_wire_2073)
    );

    and_bi _0786_ (
        .a(_0265_),
        .b(_0266_),
        .c(_0267_)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_1788),
        .dout(new_Jinkela_wire_1789)
    );

    or_bb _0787_ (
        .a(new_Jinkela_wire_1344),
        .b(new_Jinkela_wire_1860),
        .c(new_net_17)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_1764),
        .dout(new_Jinkela_wire_1765)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_2095),
        .dout(new_Jinkela_wire_2096)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_2073),
        .dout(new_Jinkela_wire_2074)
    );

    and_bi _0788_ (
        .a(new_Jinkela_wire_76),
        .b(new_Jinkela_wire_1345),
        .c(_0268_)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_1782),
        .dout(new_Jinkela_wire_1783)
    );

    and_bi _0789_ (
        .a(new_Jinkela_wire_778),
        .b(new_Jinkela_wire_1861),
        .c(_0269_)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_1765),
        .dout(new_Jinkela_wire_1766)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_2091),
        .dout(new_Jinkela_wire_2092)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(new_Jinkela_wire_2074),
        .dout(new_Jinkela_wire_2075)
    );

    or_bb _0790_ (
        .a(_0269_),
        .b(_0268_),
        .c(new_net_11)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_1796),
        .dout(new_Jinkela_wire_1797)
    );

    or_bb _0791_ (
        .a(new_Jinkela_wire_653),
        .b(new_Jinkela_wire_890),
        .c(_0270_)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_1766),
        .dout(new_Jinkela_wire_1767)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(new_Jinkela_wire_2102),
        .dout(new_Jinkela_wire_2103)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_2075),
        .dout(new_Jinkela_wire_2076)
    );

    or_bb _0792_ (
        .a(new_Jinkela_wire_2142),
        .b(new_Jinkela_wire_2408),
        .c(_0271_)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    or_bb _0793_ (
        .a(new_Jinkela_wire_1947),
        .b(new_Jinkela_wire_513),
        .c(new_net_950)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(new_Jinkela_wire_1767),
        .dout(new_Jinkela_wire_1768)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_2092),
        .dout(new_Jinkela_wire_2093)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_2076),
        .dout(new_Jinkela_wire_2077)
    );

    and_bi _0794_ (
        .a(G1),
        .b(G3),
        .c(_0272_)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_1789),
        .dout(new_Jinkela_wire_1790)
    );

    or_bb _0795_ (
        .a(new_Jinkela_wire_1597),
        .b(new_Jinkela_wire_1948),
        .c(new_net_946)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(new_Jinkela_wire_1768),
        .dout(new_Jinkela_wire_1769)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(new_Jinkela_wire_2096),
        .dout(new_Jinkela_wire_2097)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_2077),
        .dout(new_Jinkela_wire_2078)
    );

    or_bb _0796_ (
        .a(new_Jinkela_wire_1499),
        .b(new_Jinkela_wire_164),
        .c(_0273_)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    and_bi _0797_ (
        .a(new_Jinkela_wire_160),
        .b(new_Jinkela_wire_1864),
        .c(_0274_)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_1769),
        .dout(new_Jinkela_wire_1770)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_2126),
        .dout(new_Jinkela_wire_2127)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_2078),
        .dout(new_Jinkela_wire_2079)
    );

    and_bi _0798_ (
        .a(_0273_),
        .b(new_Jinkela_wire_1674),
        .c(new_net_18)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    or_bb _0799_ (
        .a(new_Jinkela_wire_1520),
        .b(new_Jinkela_wire_159),
        .c(_0275_)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_1770),
        .dout(new_Jinkela_wire_1771)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(new_Jinkela_wire_2097),
        .dout(new_Jinkela_wire_2098)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_2079),
        .dout(new_Jinkela_wire_2080)
    );

    and_bi _0800_ (
        .a(new_Jinkela_wire_2460),
        .b(new_Jinkela_wire_163),
        .c(_0276_)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_1785),
        .dout(new_Jinkela_wire_1786)
    );

    and_bi _0801_ (
        .a(new_Jinkela_wire_2609),
        .b(_0276_),
        .c(new_net_19)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_1771),
        .dout(new_Jinkela_wire_1772)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_2103),
        .dout(new_Jinkela_wire_2104)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_2080),
        .dout(new_Jinkela_wire_2081)
    );

    and_bi _0802_ (
        .a(new_Jinkela_wire_162),
        .b(new_Jinkela_wire_1720),
        .c(_0277_)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_1790),
        .dout(new_Jinkela_wire_1791)
    );

    or_bb _0803_ (
        .a(new_Jinkela_wire_148),
        .b(new_Jinkela_wire_198),
        .c(_0278_)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(new_Jinkela_wire_1772),
        .dout(new_Jinkela_wire_1773)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(new_Jinkela_wire_2098),
        .dout(new_Jinkela_wire_2099)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_2081),
        .dout(new_Jinkela_wire_2082)
    );

    and_bi _0804_ (
        .a(new_Jinkela_wire_1505),
        .b(new_Jinkela_wire_2633),
        .c(_0279_)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_1797),
        .dout(new_Jinkela_wire_1798)
    );

    or_bb _0805_ (
        .a(_0279_),
        .b(_0277_),
        .c(new_net_20)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(new_Jinkela_wire_1773),
        .dout(new_Jinkela_wire_1774)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(_0386_),
        .dout(new_Jinkela_wire_2128)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(new_Jinkela_wire_2082),
        .c(new_Jinkela_wire_2083),
        .b(new_Jinkela_wire_2084)
    );

    or_bb _0806_ (
        .a(new_Jinkela_wire_1650),
        .b(new_Jinkela_wire_500),
        .c(_0280_)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_1791),
        .dout(new_Jinkela_wire_1792)
    );

    and_bi _0807_ (
        .a(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_1652),
        .c(_0281_)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(new_Jinkela_wire_1774),
        .dout(new_Jinkela_wire_1775)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_2104),
        .dout(new_Jinkela_wire_2105)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(new_Jinkela_wire_2119),
        .dout(new_Jinkela_wire_2120)
    );

    and_bi _0808_ (
        .a(_0280_),
        .b(_0281_),
        .c(_0282_)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(_0434_),
        .dout(new_Jinkela_wire_1840)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(new_Jinkela_wire_2099),
        .dout(new_Jinkela_wire_2100)
    );

    or_bb _0809_ (
        .a(_0282_),
        .b(new_Jinkela_wire_543),
        .c(new_net_963)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(new_Jinkela_wire_1775),
        .dout(new_Jinkela_wire_1776)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_2100),
        .dout(new_Jinkela_wire_2101)
    );

    and_bi _0810_ (
        .a(new_Jinkela_wire_250),
        .b(new_Jinkela_wire_244),
        .c(_0283_)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_1792),
        .dout(new_Jinkela_wire_1793)
    );

    and_bi _0811_ (
        .a(new_Jinkela_wire_275),
        .b(new_Jinkela_wire_2620),
        .c(_0284_)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_1776),
        .dout(new_Jinkela_wire_1777)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_2105),
        .dout(new_Jinkela_wire_2106)
    );

    and_bi _0812_ (
        .a(new_Jinkela_wire_1614),
        .b(_0284_),
        .c(_0285_)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_1798),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_2120),
        .dout(new_Jinkela_wire_2121)
    );

    and_bi _0813_ (
        .a(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_1986),
        .c(_0286_)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_2106),
        .dout(new_Jinkela_wire_2107)
    );

    and_bi _0814_ (
        .a(new_Jinkela_wire_44),
        .b(new_Jinkela_wire_385),
        .c(_0287_)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(_0296_),
        .dout(new_Jinkela_wire_1855)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(_0345_),
        .c(new_Jinkela_wire_1853),
        .b(new_Jinkela_wire_1854)
    );

    and_bi _0815_ (
        .a(new_Jinkela_wire_67),
        .b(new_Jinkela_wire_1722),
        .c(_0288_)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_1794),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_2107),
        .dout(new_Jinkela_wire_2108)
    );

    and_bi _0816_ (
        .a(new_Jinkela_wire_1578),
        .b(_0288_),
        .c(_0289_)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(_0388_),
        .dout(new_Jinkela_wire_2131)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_2121),
        .dout(new_Jinkela_wire_2122)
    );

    and_bi _0817_ (
        .a(new_Jinkela_wire_1102),
        .b(new_Jinkela_wire_2384),
        .c(_0290_)
    );

    spl3L new_Jinkela_splitter_176 (
        .a(new_Jinkela_wire_1817),
        .c(new_Jinkela_wire_1818),
        .b(new_Jinkela_wire_1819),
        .d(new_Jinkela_wire_1820)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_2108),
        .dout(new_Jinkela_wire_2109)
    );

    and_bi _0818_ (
        .a(new_Jinkela_wire_46),
        .b(new_Jinkela_wire_1029),
        .c(_0291_)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    and_bi _0819_ (
        .a(new_Jinkela_wire_2457),
        .b(new_Jinkela_wire_68),
        .c(_0292_)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_2109),
        .dout(new_Jinkela_wire_2110)
    );

    and_bi _0820_ (
        .a(new_Jinkela_wire_2407),
        .b(_0292_),
        .c(_0293_)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_2128),
        .dout(new_Jinkela_wire_2129)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_2122),
        .dout(new_Jinkela_wire_2123)
    );

    and_bi _0821_ (
        .a(new_Jinkela_wire_1248),
        .b(new_Jinkela_wire_1547),
        .c(_0294_)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_2110),
        .dout(new_Jinkela_wire_2111)
    );

    bfr new_Jinkela_buffer_1681 (
        .din(new_Jinkela_wire_2275),
        .dout(new_Jinkela_wire_2276)
    );

    bfr new_Jinkela_buffer_1700 (
        .din(new_Jinkela_wire_2294),
        .dout(new_Jinkela_wire_2295)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    and_bi _0612_ (
        .a(new_Jinkela_wire_1750),
        .b(new_Jinkela_wire_1410),
        .c(_0102_)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1337),
        .dout(new_Jinkela_wire_1338)
    );

    bfr new_Jinkela_buffer_1753 (
        .din(new_Jinkela_wire_2351),
        .dout(new_Jinkela_wire_2352)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1317),
        .dout(new_Jinkela_wire_1318)
    );

    and_bi _0613_ (
        .a(new_Jinkela_wire_2389),
        .b(new_Jinkela_wire_1584),
        .c(_0103_)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    bfr new_Jinkela_buffer_1739 (
        .din(new_Jinkela_wire_2335),
        .dout(new_Jinkela_wire_2336)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_937),
        .dout(new_Jinkela_wire_938)
    );

    and_bi _0614_ (
        .a(new_Jinkela_wire_2390),
        .b(new_Jinkela_wire_1585),
        .c(_0104_)
    );

    bfr new_Jinkela_buffer_1763 (
        .din(new_Jinkela_wire_2366),
        .dout(new_Jinkela_wire_2367)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1318),
        .dout(new_Jinkela_wire_1319)
    );

    and_bi _0615_ (
        .a(_0103_),
        .b(_0104_),
        .c(_0105_)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_1740 (
        .din(new_Jinkela_wire_2336),
        .dout(new_Jinkela_wire_2337)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(_0022_),
        .dout(new_Jinkela_wire_1354)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    and_bi _0616_ (
        .a(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_1154),
        .c(_0106_)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1338),
        .dout(new_Jinkela_wire_1339)
    );

    bfr new_Jinkela_buffer_1754 (
        .din(new_Jinkela_wire_2352),
        .dout(new_Jinkela_wire_2353)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1319),
        .dout(new_Jinkela_wire_1320)
    );

    and_bi _0617_ (
        .a(new_Jinkela_wire_490),
        .b(new_Jinkela_wire_1155),
        .c(_0107_)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_1741 (
        .din(new_Jinkela_wire_2337),
        .dout(new_Jinkela_wire_2338)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    and_bi _0618_ (
        .a(_0106_),
        .b(_0107_),
        .c(_0108_)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1342),
        .dout(new_Jinkela_wire_1343)
    );

    spl2 new_Jinkela_splitter_105 (
        .a(new_Jinkela_wire_1320),
        .c(new_Jinkela_wire_1321),
        .b(new_Jinkela_wire_1322)
    );

    and_bi _0619_ (
        .a(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_531),
        .c(_0109_)
    );

    bfr new_Jinkela_buffer_757 (
        .din(G34),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_1742 (
        .din(new_Jinkela_wire_2338),
        .dout(new_Jinkela_wire_2339)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    and_bi _0620_ (
        .a(new_Jinkela_wire_343),
        .b(new_Jinkela_wire_532),
        .c(_0110_)
    );

    bfr new_Jinkela_buffer_1782 (
        .din(new_Jinkela_wire_2391),
        .dout(new_Jinkela_wire_2392)
    );

    bfr new_Jinkela_buffer_1755 (
        .din(new_Jinkela_wire_2353),
        .dout(new_Jinkela_wire_2354)
    );

    and_bi _0621_ (
        .a(_0109_),
        .b(_0110_),
        .c(_0111_)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1339),
        .dout(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_1743 (
        .din(new_Jinkela_wire_2339),
        .dout(new_Jinkela_wire_2340)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    and_bi _0622_ (
        .a(new_Jinkela_wire_1862),
        .b(new_Jinkela_wire_1568),
        .c(_0112_)
    );

    spl2 new_Jinkela_splitter_111 (
        .a(_0465_),
        .c(new_Jinkela_wire_1357),
        .b(new_Jinkela_wire_1360)
    );

    spl2 new_Jinkela_splitter_230 (
        .a(new_Jinkela_wire_2367),
        .c(new_Jinkela_wire_2368),
        .b(new_Jinkela_wire_2369)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1323),
        .dout(new_Jinkela_wire_1324)
    );

    and_bi _0623_ (
        .a(new_Jinkela_wire_1863),
        .b(new_Jinkela_wire_1569),
        .c(_0113_)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_1744 (
        .din(new_Jinkela_wire_2340),
        .dout(new_Jinkela_wire_2341)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    and_bi _0624_ (
        .a(_0112_),
        .b(_0113_),
        .c(_0114_)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(_0415_),
        .c(new_Jinkela_wire_1347),
        .b(new_Jinkela_wire_1349)
    );

    bfr new_Jinkela_buffer_1756 (
        .din(new_Jinkela_wire_2354),
        .dout(new_Jinkela_wire_2355)
    );

    and_bi _0625_ (
        .a(new_Jinkela_wire_2563),
        .b(new_Jinkela_wire_1467),
        .c(_0115_)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1347),
        .dout(new_Jinkela_wire_1348)
    );

    spl4L new_Jinkela_splitter_109 (
        .a(new_Jinkela_wire_1349),
        .c(new_Jinkela_wire_1350),
        .e(new_Jinkela_wire_1351),
        .b(new_Jinkela_wire_1352),
        .d(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    and_bi _0626_ (
        .a(new_Jinkela_wire_2564),
        .b(new_Jinkela_wire_1468),
        .c(_0116_)
    );

    spl2 new_Jinkela_splitter_110 (
        .a(_0079_),
        .c(new_Jinkela_wire_1355),
        .b(new_Jinkela_wire_1356)
    );

    bfr new_Jinkela_buffer_1764 (
        .din(new_Jinkela_wire_2369),
        .dout(new_Jinkela_wire_2370)
    );

    bfr new_Jinkela_buffer_1757 (
        .din(new_Jinkela_wire_2355),
        .dout(new_Jinkela_wire_2356)
    );

    or_bb _0627_ (
        .a(_0116_),
        .b(_0115_),
        .c(new_net_12)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    and_bi _0628_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_1146),
        .c(_0117_)
    );

    bfr new_Jinkela_buffer_1701 (
        .din(new_Jinkela_wire_2295),
        .dout(new_Jinkela_wire_2296)
    );

    bfr new_Jinkela_buffer_1789 (
        .din(_0291_),
        .dout(new_Jinkela_wire_2399)
    );

    bfr new_Jinkela_buffer_1758 (
        .din(new_Jinkela_wire_2356),
        .dout(new_Jinkela_wire_2357)
    );

    and_bi _0629_ (
        .a(new_Jinkela_wire_248),
        .b(new_Jinkela_wire_1147),
        .c(_0118_)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(_0308_),
        .c(new_Jinkela_wire_1365),
        .b(new_Jinkela_wire_1366)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    and_bi _0630_ (
        .a(_0117_),
        .b(_0118_),
        .c(_0119_)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_net_957),
        .dout(new_Jinkela_wire_1379)
    );

    spl2 new_Jinkela_splitter_233 (
        .a(new_net_11),
        .c(new_Jinkela_wire_2408),
        .b(new_Jinkela_wire_2409)
    );

    bfr new_Jinkela_buffer_1759 (
        .din(new_Jinkela_wire_2357),
        .dout(new_Jinkela_wire_2358)
    );

    and_bi _0631_ (
        .a(new_Jinkela_wire_392),
        .b(new_Jinkela_wire_887),
        .c(_0120_)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(new_Jinkela_wire_1367),
        .dout(new_Jinkela_wire_1368)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    and_bi _0632_ (
        .a(new_Jinkela_wire_393),
        .b(new_Jinkela_wire_888),
        .c(_0121_)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(new_Jinkela_wire_1357),
        .c(new_Jinkela_wire_1358),
        .b(new_Jinkela_wire_1359)
    );

    bfr new_Jinkela_buffer_1765 (
        .din(new_Jinkela_wire_2370),
        .dout(new_Jinkela_wire_2371)
    );

    bfr new_Jinkela_buffer_1760 (
        .din(new_Jinkela_wire_2358),
        .dout(new_Jinkela_wire_2359)
    );

    bfr new_Jinkela_buffer_1666 (
        .din(new_Jinkela_wire_2247),
        .dout(new_Jinkela_wire_2248)
    );

    and_bi _0633_ (
        .a(_0120_),
        .b(_0121_),
        .c(_0122_)
    );

    spl3L new_Jinkela_splitter_78 (
        .a(new_Jinkela_wire_967),
        .c(new_Jinkela_wire_968),
        .b(new_Jinkela_wire_969),
        .d(new_Jinkela_wire_970)
    );

    spl4L new_Jinkela_splitter_113 (
        .a(new_Jinkela_wire_1360),
        .c(new_Jinkela_wire_1361),
        .e(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_1363),
        .d(new_Jinkela_wire_1364)
    );

    bfr new_Jinkela_buffer_1819 (
        .din(_0364_),
        .dout(new_Jinkela_wire_2433)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    and_bi _0634_ (
        .a(new_Jinkela_wire_2554),
        .b(new_Jinkela_wire_2567),
        .c(_0123_)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(_0460_),
        .dout(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_1783 (
        .din(new_Jinkela_wire_2392),
        .dout(new_Jinkela_wire_2393)
    );

    bfr new_Jinkela_buffer_1766 (
        .din(new_Jinkela_wire_2371),
        .dout(new_Jinkela_wire_2372)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(_0496_),
        .dout(new_Jinkela_wire_1370)
    );

    and_bi _0635_ (
        .a(new_Jinkela_wire_2555),
        .b(new_Jinkela_wire_2568),
        .c(_0124_)
    );

    bfr new_Jinkela_buffer_760 (
        .din(G99),
        .dout(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_948),
        .dout(new_Jinkela_wire_949)
    );

    and_bi _0636_ (
        .a(_0123_),
        .b(_0124_),
        .c(_0125_)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1368),
        .dout(new_Jinkela_wire_1369)
    );

    bfr new_Jinkela_buffer_1790 (
        .din(new_Jinkela_wire_2399),
        .dout(new_Jinkela_wire_2400)
    );

    bfr new_Jinkela_buffer_1767 (
        .din(new_Jinkela_wire_2372),
        .dout(new_Jinkela_wire_2373)
    );

    and_bi _0637_ (
        .a(new_Jinkela_wire_230),
        .b(new_Jinkela_wire_1295),
        .c(_0126_)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1370),
        .dout(new_Jinkela_wire_1371)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    and_bi _0638_ (
        .a(new_Jinkela_wire_231),
        .b(new_Jinkela_wire_1296),
        .c(_0127_)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(_0311_),
        .dout(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_1784 (
        .din(new_Jinkela_wire_2393),
        .dout(new_Jinkela_wire_2394)
    );

    bfr new_Jinkela_buffer_1768 (
        .din(new_Jinkela_wire_2373),
        .dout(new_Jinkela_wire_2374)
    );

    and_bi _0639_ (
        .a(_0126_),
        .b(_0127_),
        .c(_0128_)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(new_Jinkela_wire_1371),
        .dout(new_Jinkela_wire_1372)
    );

    and_bi _0640_ (
        .a(new_Jinkela_wire_1962),
        .b(new_Jinkela_wire_1679),
        .c(_0129_)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1379),
        .dout(new_Jinkela_wire_1380)
    );

    bfr new_Jinkela_buffer_1769 (
        .din(new_Jinkela_wire_2374),
        .dout(new_Jinkela_wire_2375)
    );

    and_bi _0641_ (
        .a(new_Jinkela_wire_1963),
        .b(new_Jinkela_wire_1680),
        .c(_0130_)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1372),
        .dout(new_Jinkela_wire_1373)
    );

    bfr new_Jinkela_buffer_1798 (
        .din(new_Jinkela_wire_2409),
        .dout(new_Jinkela_wire_2410)
    );

    or_bb _0642_ (
        .a(_0130_),
        .b(_0129_),
        .c(_0131_)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(_0039_),
        .dout(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_1785 (
        .din(new_Jinkela_wire_2394),
        .dout(new_Jinkela_wire_2395)
    );

    bfr new_Jinkela_buffer_1770 (
        .din(new_Jinkela_wire_2375),
        .dout(new_Jinkela_wire_2376)
    );

    or_bb _0643_ (
        .a(new_Jinkela_wire_863),
        .b(new_Jinkela_wire_1085),
        .c(_0132_)
    );

    bfr new_Jinkela_buffer_764 (
        .din(G68),
        .dout(new_Jinkela_wire_992)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1373),
        .dout(new_Jinkela_wire_1374)
    );

    and_bi _0644_ (
        .a(new_Jinkela_wire_1086),
        .b(new_Jinkela_wire_864),
        .c(_0133_)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    bfr new_Jinkela_buffer_1791 (
        .din(new_Jinkela_wire_2400),
        .dout(new_Jinkela_wire_2401)
    );

    bfr new_Jinkela_buffer_1771 (
        .din(new_Jinkela_wire_2376),
        .dout(new_Jinkela_wire_2377)
    );

    and_bi _0645_ (
        .a(_0132_),
        .b(_0133_),
        .c(_0134_)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_Jinkela_wire_1374),
        .dout(new_Jinkela_wire_1375)
    );

    and_bi _0646_ (
        .a(new_Jinkela_wire_692),
        .b(new_Jinkela_wire_1197),
        .c(_0135_)
    );

    bfr new_Jinkela_buffer_767 (
        .din(G67),
        .dout(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(_0471_),
        .dout(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_1786 (
        .din(new_Jinkela_wire_2395),
        .dout(new_Jinkela_wire_2396)
    );

    bfr new_Jinkela_buffer_1772 (
        .din(new_Jinkela_wire_2377),
        .dout(new_Jinkela_wire_2378)
    );

    and_bi _0647_ (
        .a(new_Jinkela_wire_693),
        .b(new_Jinkela_wire_1198),
        .c(_0136_)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(new_Jinkela_wire_1375),
        .dout(new_Jinkela_wire_1376)
    );

    and_bi _0648_ (
        .a(_0135_),
        .b(_0136_),
        .c(_0137_)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    bfr new_Jinkela_buffer_1773 (
        .din(new_Jinkela_wire_2378),
        .dout(new_Jinkela_wire_2379)
    );

    bfr new_Jinkela_buffer_1712 (
        .din(_0313_),
        .dout(new_Jinkela_wire_2309)
    );

    or_bb _0649_ (
        .a(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_2623),
        .c(_0138_)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1376),
        .dout(new_Jinkela_wire_1377)
    );

    and_bi _0650_ (
        .a(new_Jinkela_wire_2624),
        .b(new_Jinkela_wire_1334),
        .c(_0139_)
    );

    spl2 new_Jinkela_splitter_79 (
        .a(G86),
        .c(new_Jinkela_wire_998),
        .b(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(new_Jinkela_wire_1405),
        .dout(new_Jinkela_wire_1406)
    );

    bfr new_Jinkela_buffer_1683 (
        .din(new_Jinkela_wire_2277),
        .dout(new_Jinkela_wire_2278)
    );

    bfr new_Jinkela_buffer_798 (
        .din(G15),
        .dout(new_Jinkela_wire_1028)
    );

    bfr new_Jinkela_buffer_1774 (
        .din(new_Jinkela_wire_2379),
        .dout(new_Jinkela_wire_2380)
    );

    and_bi _0651_ (
        .a(_0138_),
        .b(_0139_),
        .c(_0140_)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    bfr new_Jinkela_buffer_1787 (
        .din(new_Jinkela_wire_2396),
        .dout(new_Jinkela_wire_2397)
    );

    and_ii _0652_ (
        .a(new_Jinkela_wire_1457),
        .b(new_Jinkela_wire_2189),
        .c(_0141_)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_1792 (
        .din(new_Jinkela_wire_2401),
        .dout(new_Jinkela_wire_2402)
    );

    bfr new_Jinkela_buffer_1775 (
        .din(new_Jinkela_wire_2380),
        .dout(new_Jinkela_wire_2381)
    );

    bfr new_Jinkela_buffer_1668 (
        .din(new_Jinkela_wire_2249),
        .dout(new_Jinkela_wire_2250)
    );

    and_bb _0653_ (
        .a(new_Jinkela_wire_1458),
        .b(new_Jinkela_wire_2190),
        .c(_0142_)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(_0101_),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    bfr new_Jinkela_buffer_53 (
        .din(G103),
        .dout(new_Jinkela_wire_85)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    spl3L new_Jinkela_splitter_6 (
        .a(new_Jinkela_wire_55),
        .c(new_Jinkela_wire_56),
        .b(new_Jinkela_wire_57),
        .d(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_377 (
        .din(G83),
        .dout(new_Jinkela_wire_514)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_492),
        .dout(new_Jinkela_wire_493)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    spl4L new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_59),
        .c(new_Jinkela_wire_60),
        .e(new_Jinkela_wire_61),
        .b(new_Jinkela_wire_62),
        .d(new_Jinkela_wire_64)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    spl4L new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_64),
        .c(new_Jinkela_wire_65),
        .e(new_Jinkela_wire_66),
        .b(new_Jinkela_wire_67),
        .d(new_Jinkela_wire_68)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_493),
        .dout(new_Jinkela_wire_494)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_79),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_70 (
        .din(G24),
        .dout(new_Jinkela_wire_108)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    bfr new_Jinkela_buffer_381 (
        .din(G108),
        .dout(new_Jinkela_wire_518)
    );

    spl3L new_Jinkela_splitter_10 (
        .a(G141),
        .c(new_Jinkela_wire_89),
        .b(new_Jinkela_wire_90),
        .d(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_494),
        .dout(new_Jinkela_wire_495)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_468),
        .dout(new_Jinkela_wire_469)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_469),
        .dout(new_Jinkela_wire_470)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_91),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_495),
        .dout(new_Jinkela_wire_496)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_470),
        .dout(new_Jinkela_wire_471)
    );

    bfr new_Jinkela_buffer_72 (
        .din(G62),
        .dout(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_87),
        .dout(new_Jinkela_wire_88)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_514),
        .dout(new_Jinkela_wire_515)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_496),
        .dout(new_Jinkela_wire_497)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_108),
        .dout(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_472),
        .dout(new_Jinkela_wire_473)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    bfr new_Jinkela_buffer_78 (
        .din(G27),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_93),
        .dout(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_94),
        .dout(new_Jinkela_wire_95)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_497),
        .dout(new_Jinkela_wire_498)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_474),
        .dout(new_Jinkela_wire_475)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(G76),
        .c(new_Jinkela_wire_118),
        .b(new_Jinkela_wire_119)
    );

    bfr new_Jinkela_buffer_385 (
        .din(G42),
        .dout(new_Jinkela_wire_522)
    );

    spl2 new_Jinkela_splitter_13 (
        .a(G123),
        .c(new_Jinkela_wire_148),
        .b(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_475),
        .dout(new_Jinkela_wire_476)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_95),
        .dout(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(new_Jinkela_wire_498),
        .c(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_500)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_515),
        .dout(new_Jinkela_wire_516)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_112),
        .dout(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    spl3L new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_100),
        .c(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_102),
        .d(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_104),
        .dout(new_Jinkela_wire_105)
    );

    bfr new_Jinkela_buffer_127 (
        .din(G4),
        .dout(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    bfr new_Jinkela_buffer_1704 (
        .din(new_Jinkela_wire_2298),
        .dout(new_Jinkela_wire_2299)
    );

    bfr new_Jinkela_buffer_1688 (
        .din(new_Jinkela_wire_2282),
        .dout(new_Jinkela_wire_2283)
    );

    bfr new_Jinkela_buffer_1705 (
        .din(new_Jinkela_wire_2299),
        .dout(new_Jinkela_wire_2300)
    );

    bfr new_Jinkela_buffer_1973 (
        .din(new_Jinkela_wire_2676),
        .dout(new_Jinkela_wire_2677)
    );

    and_bi _0990_ (
        .a(_0457_),
        .b(new_Jinkela_wire_1369),
        .c(_0461_)
    );

    bfr new_Jinkela_buffer_1956 (
        .din(new_Jinkela_wire_2656),
        .dout(new_Jinkela_wire_2657)
    );

    and_bi _0991_ (
        .a(new_Jinkela_wire_2398),
        .b(_0461_),
        .c(_0462_)
    );

    spl2 new_Jinkela_splitter_273 (
        .a(new_Jinkela_wire_2701),
        .c(new_Jinkela_wire_2702),
        .b(new_Jinkela_wire_2703)
    );

    and_bi _0992_ (
        .a(new_Jinkela_wire_2056),
        .b(_0462_),
        .c(_0463_)
    );

    bfr new_Jinkela_buffer_1957 (
        .din(new_Jinkela_wire_2657),
        .dout(new_Jinkela_wire_2658)
    );

    and_bi _0993_ (
        .a(new_Jinkela_wire_1648),
        .b(_0463_),
        .c(_0464_)
    );

    bfr new_Jinkela_buffer_1974 (
        .din(new_Jinkela_wire_2677),
        .dout(new_Jinkela_wire_2678)
    );

    and_bi _0994_ (
        .a(new_Jinkela_wire_2552),
        .b(new_Jinkela_wire_2264),
        .c(_0465_)
    );

    bfr new_Jinkela_buffer_1958 (
        .din(new_Jinkela_wire_2658),
        .dout(new_Jinkela_wire_2659)
    );

    or_bb _0995_ (
        .a(new_Jinkela_wire_2151),
        .b(new_Jinkela_wire_911),
        .c(_0466_)
    );

    bfr new_Jinkela_buffer_2000 (
        .din(new_Jinkela_wire_2716),
        .dout(new_Jinkela_wire_2717)
    );

    and_bi _0996_ (
        .a(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_1328),
        .c(_0467_)
    );

    bfr new_Jinkela_buffer_1709 (
        .din(new_Jinkela_wire_2303),
        .dout(new_Jinkela_wire_2304)
    );

    bfr new_Jinkela_buffer_1959 (
        .din(new_Jinkela_wire_2659),
        .dout(new_Jinkela_wire_2660)
    );

    or_bb _0997_ (
        .a(new_Jinkela_wire_1970),
        .b(new_Jinkela_wire_1164),
        .c(_0468_)
    );

    bfr new_Jinkela_buffer_1975 (
        .din(new_Jinkela_wire_2678),
        .dout(new_Jinkela_wire_2679)
    );

    and_bi _0998_ (
        .a(new_Jinkela_wire_1364),
        .b(new_Jinkela_wire_2254),
        .c(_0469_)
    );

    bfr new_Jinkela_buffer_1960 (
        .din(new_Jinkela_wire_2660),
        .dout(new_Jinkela_wire_2661)
    );

    and_bi _0999_ (
        .a(_0467_),
        .b(_0469_),
        .c(_0470_)
    );

    or_bb _1000_ (
        .a(new_Jinkela_wire_1968),
        .b(new_Jinkela_wire_1165),
        .c(_0471_)
    );

    bfr new_Jinkela_buffer_1961 (
        .din(new_Jinkela_wire_2661),
        .dout(new_Jinkela_wire_2662)
    );

    and_bi _1001_ (
        .a(new_Jinkela_wire_1359),
        .b(new_Jinkela_wire_1409),
        .c(_0472_)
    );

    bfr new_Jinkela_buffer_1692 (
        .din(new_Jinkela_wire_2286),
        .dout(new_Jinkela_wire_2287)
    );

    spl4L new_Jinkela_splitter_275 (
        .a(new_Jinkela_wire_2709),
        .c(new_Jinkela_wire_2710),
        .e(new_Jinkela_wire_2711),
        .b(new_Jinkela_wire_2712),
        .d(new_Jinkela_wire_2713)
    );

    bfr new_Jinkela_buffer_1976 (
        .din(new_Jinkela_wire_2679),
        .dout(new_Jinkela_wire_2680)
    );

    or_bb _1002_ (
        .a(new_Jinkela_wire_2618),
        .b(new_Jinkela_wire_1184),
        .c(_0473_)
    );

    bfr new_Jinkela_buffer_1962 (
        .din(new_Jinkela_wire_2662),
        .dout(new_Jinkela_wire_2663)
    );

    and_bi _1003_ (
        .a(new_Jinkela_wire_836),
        .b(new_Jinkela_wire_2270),
        .c(_0474_)
    );

    and_bi _1004_ (
        .a(new_Jinkela_wire_2541),
        .b(_0474_),
        .c(_0475_)
    );

    bfr new_Jinkela_buffer_1963 (
        .din(new_Jinkela_wire_2663),
        .dout(new_Jinkela_wire_2664)
    );

    and_bi _1005_ (
        .a(new_Jinkela_wire_1358),
        .b(_0475_),
        .c(_0476_)
    );

    bfr new_Jinkela_buffer_1998 (
        .din(new_Jinkela_wire_2714),
        .dout(new_Jinkela_wire_2715)
    );

    bfr new_Jinkela_buffer_1977 (
        .din(new_Jinkela_wire_2680),
        .dout(new_Jinkela_wire_2681)
    );

    and_ii _1006_ (
        .a(new_Jinkela_wire_2493),
        .b(new_Jinkela_wire_1617),
        .c(_0477_)
    );

    bfr new_Jinkela_buffer_1964 (
        .din(new_Jinkela_wire_2664),
        .dout(new_Jinkela_wire_2665)
    );

    or_bb _1007_ (
        .a(new_Jinkela_wire_2150),
        .b(new_Jinkela_wire_912),
        .c(_0478_)
    );

    and_bi _1008_ (
        .a(new_Jinkela_wire_1183),
        .b(new_Jinkela_wire_2615),
        .c(_0479_)
    );

    bfr new_Jinkela_buffer_1965 (
        .din(new_Jinkela_wire_2665),
        .dout(new_Jinkela_wire_2666)
    );

    and_bi _1009_ (
        .a(new_Jinkela_wire_1329),
        .b(_0479_),
        .c(_0480_)
    );

    bfr new_Jinkela_buffer_2008 (
        .din(new_net_946),
        .dout(new_Jinkela_wire_2725)
    );

    bfr new_Jinkela_buffer_1978 (
        .din(new_Jinkela_wire_2681),
        .dout(new_Jinkela_wire_2682)
    );

    and_bi _1010_ (
        .a(new_Jinkela_wire_1363),
        .b(new_Jinkela_wire_1587),
        .c(_0481_)
    );

    bfr new_Jinkela_buffer_1966 (
        .din(new_Jinkela_wire_2666),
        .dout(new_Jinkela_wire_2667)
    );

    or_bb _1011_ (
        .a(new_Jinkela_wire_2274),
        .b(new_Jinkela_wire_837),
        .c(_0482_)
    );

    and_bi _1012_ (
        .a(new_Jinkela_wire_1361),
        .b(new_Jinkela_wire_1346),
        .c(_0483_)
    );

    bfr new_Jinkela_buffer_1967 (
        .din(new_Jinkela_wire_2667),
        .dout(new_Jinkela_wire_2668)
    );

    or_bb _1013_ (
        .a(new_Jinkela_wire_1972),
        .b(new_Jinkela_wire_2558),
        .c(_0484_)
    );

    bfr new_Jinkela_buffer_1979 (
        .din(new_Jinkela_wire_2682),
        .dout(new_Jinkela_wire_2683)
    );

    and_bi _1014_ (
        .a(_0477_),
        .b(_0484_),
        .c(_0485_)
    );

    bfr new_Jinkela_buffer_1968 (
        .din(new_Jinkela_wire_2668),
        .dout(new_Jinkela_wire_2669)
    );

    or_ii _1015_ (
        .a(_0485_),
        .b(new_Jinkela_wire_2497),
        .c(_0486_)
    );

    or_bb _1016_ (
        .a(new_Jinkela_wire_2644),
        .b(_0464_),
        .c(_0487_)
    );

    bfr new_Jinkela_buffer_1969 (
        .din(new_Jinkela_wire_2669),
        .dout(new_Jinkela_wire_2670)
    );

    and_bi _1017_ (
        .a(new_Jinkela_wire_2545),
        .b(new_Jinkela_wire_1973),
        .c(_0488_)
    );

    bfr new_Jinkela_buffer_2001 (
        .din(new_Jinkela_wire_2717),
        .dout(new_Jinkela_wire_2718)
    );

    bfr new_Jinkela_buffer_1980 (
        .din(new_Jinkela_wire_2683),
        .dout(new_Jinkela_wire_2684)
    );

    and_bi _1018_ (
        .a(new_Jinkela_wire_2560),
        .b(_0488_),
        .c(_0489_)
    );

    and_bi _1019_ (
        .a(new_Jinkela_wire_2498),
        .b(_0489_),
        .c(_0490_)
    );

    bfr new_Jinkela_buffer_2009 (
        .din(new_Jinkela_wire_2725),
        .dout(new_Jinkela_wire_2726)
    );

    bfr new_Jinkela_buffer_1981 (
        .din(new_Jinkela_wire_2684),
        .dout(new_Jinkela_wire_2685)
    );

    or_bb _1020_ (
        .a(_0490_),
        .b(new_Jinkela_wire_1621),
        .c(_0491_)
    );

    and_bi _1021_ (
        .a(_0487_),
        .b(new_Jinkela_wire_1442),
        .c(G2591)
    );

    bfr new_Jinkela_buffer_2002 (
        .din(new_Jinkela_wire_2718),
        .dout(new_Jinkela_wire_2719)
    );

    bfr new_Jinkela_buffer_1982 (
        .din(new_Jinkela_wire_2685),
        .dout(new_Jinkela_wire_2686)
    );

    or_bb _1022_ (
        .a(new_Jinkela_wire_2413),
        .b(new_Jinkela_wire_1414),
        .c(_0492_)
    );

    or_bb _1023_ (
        .a(new_Jinkela_wire_2548),
        .b(new_Jinkela_wire_2342),
        .c(_0493_)
    );

    bfr new_Jinkela_buffer_1983 (
        .din(new_Jinkela_wire_2686),
        .dout(new_Jinkela_wire_2687)
    );

    or_bb _1024_ (
        .a(_0493_),
        .b(new_Jinkela_wire_1895),
        .c(_0494_)
    );

    or_bb _1025_ (
        .a(new_Jinkela_wire_2300),
        .b(new_Jinkela_wire_1681),
        .c(_0495_)
    );

    bfr new_Jinkela_buffer_2003 (
        .din(new_Jinkela_wire_2719),
        .dout(new_Jinkela_wire_2720)
    );

    bfr new_Jinkela_buffer_1984 (
        .din(new_Jinkela_wire_2687),
        .dout(new_Jinkela_wire_2688)
    );

    or_bb _1026_ (
        .a(new_Jinkela_wire_2086),
        .b(new_Jinkela_wire_1459),
        .c(new_net_23)
    );

    and_bi _1027_ (
        .a(new_Jinkela_wire_791),
        .b(new_Jinkela_wire_1143),
        .c(new_net_954)
    );

    bfr new_Jinkela_buffer_2010 (
        .din(new_Jinkela_wire_2726),
        .dout(new_Jinkela_wire_2727)
    );

    bfr new_Jinkela_buffer_1985 (
        .din(new_Jinkela_wire_2688),
        .dout(new_Jinkela_wire_2689)
    );

    or_bb _1028_ (
        .a(new_Jinkela_wire_1719),
        .b(new_Jinkela_wire_1042),
        .c(new_net_948)
    );

    bfr new_Jinkela_buffer_1714 (
        .din(new_Jinkela_wire_2310),
        .dout(new_Jinkela_wire_2311)
    );

    and_bi _1029_ (
        .a(new_Jinkela_wire_199),
        .b(new_Jinkela_wire_1030),
        .c(_0496_)
    );

    bfr new_Jinkela_buffer_2004 (
        .din(new_Jinkela_wire_2720),
        .dout(new_Jinkela_wire_2721)
    );

    bfr new_Jinkela_buffer_1986 (
        .din(new_Jinkela_wire_2689),
        .dout(new_Jinkela_wire_2690)
    );

    or_bb _1030_ (
        .a(new_Jinkela_wire_1378),
        .b(new_Jinkela_wire_1502),
        .c(new_net_961)
    );

    and_bi _1031_ (
        .a(new_Jinkela_wire_1049),
        .b(new_Jinkela_wire_1470),
        .c(_0497_)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    spl2 new_Jinkela_splitter_183 (
        .a(_0264_),
        .c(new_Jinkela_wire_1860),
        .b(new_Jinkela_wire_1861)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_105),
        .dout(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_Jinkela_wire_1802),
        .dout(new_Jinkela_wire_1803)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    spl4L new_Jinkela_splitter_180 (
        .a(new_Jinkela_wire_1848),
        .c(new_Jinkela_wire_1849),
        .e(new_Jinkela_wire_1850),
        .b(new_Jinkela_wire_1851),
        .d(new_Jinkela_wire_1852)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_2111),
        .dout(new_Jinkela_wire_2112)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_1820),
        .dout(new_Jinkela_wire_1821)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_106),
        .dout(new_Jinkela_wire_107)
    );

    spl2 new_Jinkela_splitter_80 (
        .a(G122),
        .c(new_Jinkela_wire_1030),
        .b(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_1803),
        .dout(new_Jinkela_wire_1804)
    );

    spl3L new_Jinkela_splitter_83 (
        .a(G129),
        .c(new_Jinkela_wire_1056),
        .b(new_Jinkela_wire_1057),
        .d(new_Jinkela_wire_1058)
    );

    spl2 new_Jinkela_splitter_211 (
        .a(new_Jinkela_wire_2123),
        .c(new_Jinkela_wire_2124),
        .b(new_Jinkela_wire_2125)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(_0270_),
        .dout(new_Jinkela_wire_2138)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_2112),
        .dout(new_Jinkela_wire_2113)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_1804),
        .dout(new_Jinkela_wire_1805)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    spl4L new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_1843),
        .c(new_Jinkela_wire_1844),
        .e(new_Jinkela_wire_1845),
        .b(new_Jinkela_wire_1846),
        .d(new_Jinkela_wire_1847)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_2113),
        .dout(new_Jinkela_wire_2114)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    spl3L new_Jinkela_splitter_18 (
        .a(G118),
        .c(new_Jinkela_wire_198),
        .b(new_Jinkela_wire_199),
        .d(new_Jinkela_wire_200)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_1805),
        .dout(new_Jinkela_wire_1806)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_Jinkela_wire_2131),
        .dout(new_Jinkela_wire_2132)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_1051),
        .dout(new_Jinkela_wire_1052)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_2114),
        .dout(new_Jinkela_wire_2115)
    );

    spl3L new_Jinkela_splitter_19 (
        .a(G133),
        .c(new_Jinkela_wire_211),
        .b(new_Jinkela_wire_212),
        .d(new_Jinkela_wire_213)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_1806),
        .dout(new_Jinkela_wire_1807)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(new_Jinkela_wire_2129),
        .dout(new_Jinkela_wire_2130)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_831 (
        .din(G18),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_2115),
        .dout(new_Jinkela_wire_2116)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_1822),
        .dout(new_Jinkela_wire_1823)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    spl4L new_Jinkela_splitter_212 (
        .a(_0413_),
        .c(new_Jinkela_wire_2143),
        .e(new_Jinkela_wire_2144),
        .b(new_Jinkela_wire_2145),
        .d(new_Jinkela_wire_2146)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(_0442_),
        .dout(new_Jinkela_wire_2147)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1050),
        .dout(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_2116),
        .dout(new_Jinkela_wire_2117)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(G150),
        .c(new_Jinkela_wire_230),
        .b(new_Jinkela_wire_231)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_1841),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(new_Jinkela_wire_2132),
        .dout(new_Jinkela_wire_2133)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(new_Jinkela_wire_1856),
        .dout(new_Jinkela_wire_1857)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_2117),
        .dout(new_Jinkela_wire_2118)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    spl2 new_Jinkela_splitter_177 (
        .a(new_Jinkela_wire_1823),
        .c(new_Jinkela_wire_1824),
        .b(new_Jinkela_wire_1825)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_2138),
        .dout(new_Jinkela_wire_2139)
    );

    and_bi _0547_ (
        .a(new_Jinkela_wire_1406),
        .b(_0042_),
        .c(new_net_5)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(new_Jinkela_wire_2133),
        .dout(new_Jinkela_wire_2134)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_1810),
        .dout(new_Jinkela_wire_1811)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_net_18),
        .dout(new_Jinkela_wire_2155)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1058),
        .dout(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_814 (
        .din(G45),
        .dout(new_Jinkela_wire_1050)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(new_Jinkela_wire_2134),
        .dout(new_Jinkela_wire_2135)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_1811),
        .dout(new_Jinkela_wire_1812)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(new_Jinkela_wire_2139),
        .dout(new_Jinkela_wire_2140)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(new_Jinkela_wire_2011),
        .dout(new_Jinkela_wire_2012)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(_0206_),
        .c(new_Jinkela_wire_1858),
        .b(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(new_Jinkela_wire_2135),
        .dout(new_Jinkela_wire_2136)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    spl3L new_Jinkela_splitter_16 (
        .a(G142),
        .c(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_180),
        .d(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(new_Jinkela_wire_2152),
        .c(new_Jinkela_wire_2153),
        .b(new_Jinkela_wire_2154)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_Jinkela_wire_2147),
        .dout(new_Jinkela_wire_2148)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(_0053_),
        .dout(new_Jinkela_wire_1856)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(new_Jinkela_wire_2136),
        .dout(new_Jinkela_wire_2137)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(new_Jinkela_wire_1826),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_2140),
        .dout(new_Jinkela_wire_2141)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    spl4L new_Jinkela_splitter_213 (
        .a(_0163_),
        .c(new_Jinkela_wire_2149),
        .e(new_Jinkela_wire_2150),
        .b(new_Jinkela_wire_2151),
        .d(new_Jinkela_wire_2152)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_2141),
        .dout(new_Jinkela_wire_2142)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_833 (
        .din(G6),
        .dout(new_Jinkela_wire_1075)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1052),
        .dout(new_Jinkela_wire_1053)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_154),
        .dout(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1011),
        .dout(new_Jinkela_wire_1012)
    );

    spl3L new_Jinkela_splitter_185 (
        .a(new_net_7),
        .c(new_Jinkela_wire_1864),
        .b(new_Jinkela_wire_1865),
        .d(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_1600 (
        .din(_0327_),
        .dout(new_Jinkela_wire_2172)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    bfr new_Jinkela_buffer_1603 (
        .din(_0370_),
        .dout(new_Jinkela_wire_2177)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    spl4L new_Jinkela_splitter_22 (
        .a(G145),
        .c(new_Jinkela_wire_232),
        .e(new_Jinkela_wire_233),
        .b(new_Jinkela_wire_234),
        .d(new_Jinkela_wire_235)
    );

    spl2 new_Jinkela_splitter_184 (
        .a(_0108_),
        .c(new_Jinkela_wire_1862),
        .b(new_Jinkela_wire_1863)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(_0240_),
        .c(new_Jinkela_wire_2175),
        .b(new_Jinkela_wire_2176)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_155),
        .dout(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1013),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_2155),
        .dout(new_Jinkela_wire_2156)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_1891),
        .dout(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_1601 (
        .din(new_Jinkela_wire_2172),
        .dout(new_Jinkela_wire_2173)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(new_Jinkela_wire_1830),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_2156),
        .dout(new_Jinkela_wire_2157)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(_0336_),
        .dout(new_Jinkela_wire_1891)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    spl2 new_Jinkela_splitter_218 (
        .a(_0429_),
        .c(new_Jinkela_wire_2185),
        .b(new_Jinkela_wire_2186)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1073),
        .dout(new_Jinkela_wire_1074)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_1053),
        .dout(new_Jinkela_wire_1054)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_2157),
        .dout(new_Jinkela_wire_2158)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    bfr new_Jinkela_buffer_1604 (
        .din(new_Jinkela_wire_2177),
        .dout(new_Jinkela_wire_2178)
    );

    spl3L new_Jinkela_splitter_186 (
        .a(new_Jinkela_wire_1866),
        .c(new_Jinkela_wire_1867),
        .b(new_Jinkela_wire_1868),
        .d(new_Jinkela_wire_1869)
    );

    bfr new_Jinkela_buffer_1602 (
        .din(new_Jinkela_wire_2173),
        .dout(new_Jinkela_wire_2174)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_136),
        .dout(new_Jinkela_wire_137)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_1832),
        .dout(new_Jinkela_wire_1833)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(new_Jinkela_wire_2158),
        .dout(new_Jinkela_wire_2159)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1016),
        .dout(new_Jinkela_wire_1017)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_Jinkela_wire_1869),
        .dout(new_Jinkela_wire_1870)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_137),
        .dout(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_1833),
        .dout(new_Jinkela_wire_1834)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(new_Jinkela_wire_2159),
        .dout(new_Jinkela_wire_2160)
    );

    spl4L new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_157),
        .c(new_Jinkela_wire_158),
        .e(new_Jinkela_wire_159),
        .b(new_Jinkela_wire_160),
        .d(new_Jinkela_wire_161)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1017),
        .dout(new_Jinkela_wire_1018)
    );

    spl2 new_Jinkela_splitter_189 (
        .a(new_net_14),
        .c(new_Jinkela_wire_1895),
        .b(new_Jinkela_wire_1896)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(_0360_),
        .c(new_Jinkela_wire_2183),
        .b(new_Jinkela_wire_2184)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(new_Jinkela_wire_1834),
        .dout(new_Jinkela_wire_1835)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(new_Jinkela_wire_2160),
        .dout(new_Jinkela_wire_2161)
    );

    spl4L new_Jinkela_splitter_15 (
        .a(new_Jinkela_wire_161),
        .c(new_Jinkela_wire_162),
        .e(new_Jinkela_wire_163),
        .b(new_Jinkela_wire_164),
        .d(new_Jinkela_wire_165)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_1018),
        .dout(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_1896),
        .dout(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(_0050_),
        .dout(new_Jinkela_wire_1912)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_2161),
        .dout(new_Jinkela_wire_2162)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1054),
        .dout(new_Jinkela_wire_1055)
    );

    or_bb _0822_ (
        .a(_0294_),
        .b(_0290_),
        .c(_0295_)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1383),
        .dout(new_Jinkela_wire_1384)
    );

    bfr new_Jinkela_buffer_391 (
        .din(G63),
        .dout(new_Jinkela_wire_528)
    );

    or_bb _0823_ (
        .a(_0295_),
        .b(new_Jinkela_wire_1713),
        .c(_0296_)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_1407),
        .dout(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    and_bi _0824_ (
        .a(new_Jinkela_wire_41),
        .b(new_Jinkela_wire_246),
        .c(_0297_)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(new_Jinkela_wire_1384),
        .dout(new_Jinkela_wire_1385)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_519),
        .dout(new_Jinkela_wire_520)
    );

    and_bi _0825_ (
        .a(new_Jinkela_wire_60),
        .b(new_Jinkela_wire_1865),
        .c(_0298_)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(_0036_),
        .dout(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_522),
        .dout(new_Jinkela_wire_523)
    );

    and_bi _0826_ (
        .a(new_Jinkela_wire_2101),
        .b(_0298_),
        .c(_0299_)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1385),
        .dout(new_Jinkela_wire_1386)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_520),
        .dout(new_Jinkela_wire_521)
    );

    and_bi _0827_ (
        .a(new_Jinkela_wire_1070),
        .b(new_Jinkela_wire_1514),
        .c(_0300_)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_404 (
        .din(G84),
        .dout(new_Jinkela_wire_544)
    );

    spl3L new_Jinkela_splitter_47 (
        .a(G144),
        .c(new_Jinkela_wire_531),
        .b(new_Jinkela_wire_532),
        .d(new_Jinkela_wire_533)
    );

    and_bi _0828_ (
        .a(new_Jinkela_wire_257),
        .b(new_Jinkela_wire_1298),
        .c(_0301_)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1386),
        .dout(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_523),
        .dout(new_Jinkela_wire_524)
    );

    and_bi _0829_ (
        .a(new_Jinkela_wire_267),
        .b(new_Jinkela_wire_2646),
        .c(_0302_)
    );

    spl2 new_Jinkela_splitter_115 (
        .a(_0180_),
        .c(new_Jinkela_wire_1412),
        .b(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(new_net_12),
        .c(new_Jinkela_wire_1414),
        .b(new_Jinkela_wire_1415)
    );

    and_bi _0830_ (
        .a(new_Jinkela_wire_1673),
        .b(_0302_),
        .c(_0303_)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1387),
        .dout(new_Jinkela_wire_1388)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_524),
        .dout(new_Jinkela_wire_525)
    );

    and_bi _0831_ (
        .a(new_Jinkela_wire_969),
        .b(new_Jinkela_wire_1588),
        .c(_0304_)
    );

    bfr new_Jinkela_buffer_408 (
        .din(G87),
        .dout(new_Jinkela_wire_548)
    );

    or_bb _0832_ (
        .a(new_Jinkela_wire_2613),
        .b(_0300_),
        .c(_0305_)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_Jinkela_wire_1388),
        .dout(new_Jinkela_wire_1389)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_525),
        .dout(new_Jinkela_wire_526)
    );

    and_bi _0833_ (
        .a(new_Jinkela_wire_258),
        .b(new_Jinkela_wire_117),
        .c(_0306_)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    and_bi _0834_ (
        .a(new_Jinkela_wire_266),
        .b(new_Jinkela_wire_2575),
        .c(_0307_)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1389),
        .dout(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_526),
        .dout(new_Jinkela_wire_527)
    );

    and_bi _0835_ (
        .a(new_Jinkela_wire_2608),
        .b(_0307_),
        .c(_0308_)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(_0491_),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    and_bi _0836_ (
        .a(new_Jinkela_wire_191),
        .b(new_Jinkela_wire_1365),
        .c(_0309_)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_1390),
        .dout(new_Jinkela_wire_1391)
    );

    and_bi _0837_ (
        .a(new_Jinkela_wire_1189),
        .b(new_Jinkela_wire_1987),
        .c(_0310_)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(_0064_),
        .dout(new_Jinkela_wire_1443)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_534),
        .dout(new_Jinkela_wire_535)
    );

    or_bb _0838_ (
        .a(_0310_),
        .b(new_Jinkela_wire_1714),
        .c(_0311_)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_1391),
        .dout(new_Jinkela_wire_1392)
    );

    or_bb _0839_ (
        .a(new_Jinkela_wire_1404),
        .b(_0305_),
        .c(_0312_)
    );

    bfr new_Jinkela_buffer_412 (
        .din(G104),
        .dout(new_Jinkela_wire_552)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_535),
        .dout(new_Jinkela_wire_536)
    );

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    and_bi _0840_ (
        .a(new_Jinkela_wire_43),
        .b(new_Jinkela_wire_488),
        .c(_0313_)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_1392),
        .dout(new_Jinkela_wire_1393)
    );

    and_bi _0841_ (
        .a(new_Jinkela_wire_1519),
        .b(new_Jinkela_wire_58),
        .c(_0314_)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    and_bi _0842_ (
        .a(new_Jinkela_wire_2316),
        .b(_0314_),
        .c(_0315_)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(new_Jinkela_wire_1393),
        .dout(new_Jinkela_wire_1394)
    );

    and_bi _0843_ (
        .a(new_Jinkela_wire_1293),
        .b(new_Jinkela_wire_1478),
        .c(_0316_)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_537),
        .dout(new_Jinkela_wire_538)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    and_bi _0844_ (
        .a(new_Jinkela_wire_47),
        .b(new_Jinkela_wire_178),
        .c(_0317_)
    );

    spl2 new_Jinkela_splitter_117 (
        .a(_0353_),
        .c(new_Jinkela_wire_1444),
        .b(new_Jinkela_wire_1445)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_Jinkela_wire_1394),
        .dout(new_Jinkela_wire_1395)
    );

    and_bi _0845_ (
        .a(new_Jinkela_wire_66),
        .b(new_Jinkela_wire_1506),
        .c(_0318_)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_546),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(_0382_),
        .dout(new_Jinkela_wire_1446)
    );

    and_bi _0846_ (
        .a(new_Jinkela_wire_1795),
        .b(_0318_),
        .c(_0319_)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    and_bi _0847_ (
        .a(new_Jinkela_wire_879),
        .b(new_Jinkela_wire_1476),
        .c(_0320_)
    );

    spl3L new_Jinkela_splitter_48 (
        .a(G132),
        .c(new_Jinkela_wire_556),
        .b(new_Jinkela_wire_557),
        .d(new_Jinkela_wire_558)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_539),
        .dout(new_Jinkela_wire_540)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    or_bb _0848_ (
        .a(_0320_),
        .b(new_Jinkela_wire_2085),
        .c(_0321_)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_1396),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_429 (
        .din(G80),
        .dout(new_Jinkela_wire_575)
    );

    and_bi _0849_ (
        .a(new_Jinkela_wire_255),
        .b(new_Jinkela_wire_20),
        .c(_0322_)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_540),
        .dout(new_Jinkela_wire_541)
    );

    and_bi _0850_ (
        .a(new_Jinkela_wire_271),
        .b(new_Jinkela_wire_1753),
        .c(_0323_)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    and_bi _0851_ (
        .a(new_Jinkela_wire_1340),
        .b(_0323_),
        .c(_0324_)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    and_bi _0852_ (
        .a(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_2610),
        .c(_0325_)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(_0085_),
        .c(new_Jinkela_wire_1447),
        .b(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_1398),
        .dout(new_Jinkela_wire_1399)
    );

    and_bi _0853_ (
        .a(new_Jinkela_wire_968),
        .b(new_Jinkela_wire_1589),
        .c(_0326_)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_net_23),
        .dout(new_Jinkela_wire_1449)
    );

    or_bb _0854_ (
        .a(_0326_),
        .b(_0325_),
        .c(_0327_)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_1399),
        .dout(new_Jinkela_wire_1400)
    );

    or_bb _0855_ (
        .a(new_Jinkela_wire_2174),
        .b(_0321_),
        .c(_0328_)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_558),
        .dout(new_Jinkela_wire_559)
    );

    or_bb _0856_ (
        .a(_0328_),
        .b(new_Jinkela_wire_2549),
        .c(_0329_)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_1400),
        .dout(new_Jinkela_wire_1401)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    or_bb _0857_ (
        .a(_0329_),
        .b(new_Jinkela_wire_1855),
        .c(_0330_)
    );

    bfr new_Jinkela_buffer_433 (
        .din(G36),
        .dout(new_Jinkela_wire_579)
    );

    and_bi _0858_ (
        .a(new_Jinkela_wire_254),
        .b(new_Jinkela_wire_109),
        .c(_0331_)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_1401),
        .dout(new_Jinkela_wire_1402)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    and_bi _0859_ (
        .a(new_Jinkela_wire_270),
        .b(new_Jinkela_wire_2149),
        .c(_0332_)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    and_bi _0860_ (
        .a(new_Jinkela_wire_2225),
        .b(_0332_),
        .c(_0333_)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_1402),
        .dout(new_Jinkela_wire_1403)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    or_bb _0861_ (
        .a(new_Jinkela_wire_2556),
        .b(new_Jinkela_wire_916),
        .c(_0334_)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    and_bi _0862_ (
        .a(new_Jinkela_wire_917),
        .b(new_Jinkela_wire_2557),
        .c(_0335_)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_1422),
        .dout(new_Jinkela_wire_1423)
    );

    bfr new_Jinkela_buffer_436 (
        .din(G10),
        .dout(new_Jinkela_wire_582)
    );

    and_bi _0863_ (
        .a(_0334_),
        .b(_0335_),
        .c(_0336_)
    );

    bfr new_Jinkela_buffer_578 (
        .din(G38),
        .dout(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_667),
        .dout(new_Jinkela_wire_668)
    );

    bfr new_Jinkela_buffer_1788 (
        .din(new_Jinkela_wire_2397),
        .dout(new_Jinkela_wire_2398)
    );

    bfr new_Jinkela_buffer_1776 (
        .din(new_Jinkela_wire_2381),
        .dout(new_Jinkela_wire_2382)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_695),
        .dout(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_668),
        .dout(new_Jinkela_wire_669)
    );

    bfr new_Jinkela_buffer_1827 (
        .din(_0498_),
        .dout(new_Jinkela_wire_2441)
    );

    bfr new_Jinkela_buffer_1777 (
        .din(new_Jinkela_wire_2382),
        .dout(new_Jinkela_wire_2383)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_669),
        .dout(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_1793 (
        .din(new_Jinkela_wire_2402),
        .dout(new_Jinkela_wire_2403)
    );

    bfr new_Jinkela_buffer_585 (
        .din(G61),
        .dout(new_Jinkela_wire_768)
    );

    bfr new_Jinkela_buffer_1820 (
        .din(new_Jinkela_wire_2433),
        .dout(new_Jinkela_wire_2434)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_696),
        .dout(new_Jinkela_wire_697)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_670),
        .dout(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_1794 (
        .din(new_Jinkela_wire_2403),
        .dout(new_Jinkela_wire_2404)
    );

    bfr new_Jinkela_buffer_1799 (
        .din(new_Jinkela_wire_2410),
        .dout(new_Jinkela_wire_2411)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    bfr new_Jinkela_buffer_1795 (
        .din(new_Jinkela_wire_2404),
        .dout(new_Jinkela_wire_2405)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_1834 (
        .din(_0371_),
        .dout(new_Jinkela_wire_2448)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_697),
        .dout(new_Jinkela_wire_698)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_1796 (
        .din(new_Jinkela_wire_2405),
        .dout(new_Jinkela_wire_2406)
    );

    bfr new_Jinkela_buffer_1800 (
        .din(new_Jinkela_wire_2411),
        .dout(new_Jinkela_wire_2412)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    bfr new_Jinkela_buffer_1797 (
        .din(new_Jinkela_wire_2406),
        .dout(new_Jinkela_wire_2407)
    );

    bfr new_Jinkela_buffer_1821 (
        .din(new_Jinkela_wire_2434),
        .dout(new_Jinkela_wire_2435)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_698),
        .dout(new_Jinkela_wire_699)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(new_Jinkela_wire_2412),
        .c(new_Jinkela_wire_2413),
        .b(new_Jinkela_wire_2414)
    );

    bfr new_Jinkela_buffer_1801 (
        .din(new_Jinkela_wire_2414),
        .dout(new_Jinkela_wire_2415)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_1828 (
        .din(new_Jinkela_wire_2441),
        .dout(new_Jinkela_wire_2442)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_726),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_1822 (
        .din(new_Jinkela_wire_2435),
        .dout(new_Jinkela_wire_2436)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_676),
        .dout(new_Jinkela_wire_677)
    );

    bfr new_Jinkela_buffer_1802 (
        .din(new_Jinkela_wire_2415),
        .dout(new_Jinkela_wire_2416)
    );

    spl3L new_Jinkela_splitter_235 (
        .a(_0226_),
        .c(new_Jinkela_wire_2451),
        .b(new_Jinkela_wire_2452),
        .d(new_Jinkela_wire_2453)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(new_net_8),
        .c(new_Jinkela_wire_2456),
        .b(new_Jinkela_wire_2459)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    bfr new_Jinkela_buffer_1803 (
        .din(new_Jinkela_wire_2416),
        .dout(new_Jinkela_wire_2417)
    );

    bfr new_Jinkela_buffer_1823 (
        .din(new_Jinkela_wire_2436),
        .dout(new_Jinkela_wire_2437)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_678),
        .dout(new_Jinkela_wire_679)
    );

    bfr new_Jinkela_buffer_1804 (
        .din(new_Jinkela_wire_2417),
        .dout(new_Jinkela_wire_2418)
    );

    bfr new_Jinkela_buffer_1829 (
        .din(new_Jinkela_wire_2442),
        .dout(new_Jinkela_wire_2443)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_1805 (
        .din(new_Jinkela_wire_2418),
        .dout(new_Jinkela_wire_2419)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_1824 (
        .din(new_Jinkela_wire_2437),
        .dout(new_Jinkela_wire_2438)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_1806 (
        .din(new_Jinkela_wire_2419),
        .dout(new_Jinkela_wire_2420)
    );

    bfr new_Jinkela_buffer_1835 (
        .din(new_Jinkela_wire_2448),
        .dout(new_Jinkela_wire_2449)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    bfr new_Jinkela_buffer_1807 (
        .din(new_Jinkela_wire_2420),
        .dout(new_Jinkela_wire_2421)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    bfr new_Jinkela_buffer_1825 (
        .din(new_Jinkela_wire_2438),
        .dout(new_Jinkela_wire_2439)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_702),
        .dout(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_682),
        .dout(new_Jinkela_wire_683)
    );

    bfr new_Jinkela_buffer_1808 (
        .din(new_Jinkela_wire_2421),
        .dout(new_Jinkela_wire_2422)
    );

    bfr new_Jinkela_buffer_1830 (
        .din(new_Jinkela_wire_2443),
        .dout(new_Jinkela_wire_2444)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_731),
        .dout(new_Jinkela_wire_732)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_1809 (
        .din(new_Jinkela_wire_2422),
        .dout(new_Jinkela_wire_2423)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_1826 (
        .din(new_Jinkela_wire_2439),
        .dout(new_Jinkela_wire_2440)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_1810 (
        .din(new_Jinkela_wire_2423),
        .dout(new_Jinkela_wire_2424)
    );

    spl3L new_Jinkela_splitter_241 (
        .a(_0218_),
        .c(new_Jinkela_wire_2483),
        .b(new_Jinkela_wire_2484),
        .d(new_Jinkela_wire_2485)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    bfr new_Jinkela_buffer_1811 (
        .din(new_Jinkela_wire_2424),
        .dout(new_Jinkela_wire_2425)
    );

    bfr new_Jinkela_buffer_1831 (
        .din(new_Jinkela_wire_2444),
        .dout(new_Jinkela_wire_2445)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_704),
        .dout(new_Jinkela_wire_705)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_686),
        .dout(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_1812 (
        .din(new_Jinkela_wire_2425),
        .dout(new_Jinkela_wire_2426)
    );

    bfr new_Jinkela_buffer_1836 (
        .din(new_Jinkela_wire_2449),
        .dout(new_Jinkela_wire_2450)
    );

    bfr new_Jinkela_buffer_581 (
        .din(G105),
        .dout(new_Jinkela_wire_764)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_1813 (
        .din(new_Jinkela_wire_2426),
        .dout(new_Jinkela_wire_2427)
    );

    bfr new_Jinkela_buffer_1832 (
        .din(new_Jinkela_wire_2445),
        .dout(new_Jinkela_wire_2446)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    or_bb _0654_ (
        .a(_0142_),
        .b(new_Jinkela_wire_592),
        .c(_0143_)
    );

    spl2 new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_1039),
        .c(new_Jinkela_wire_1040),
        .b(new_Jinkela_wire_1041)
    );

    and_bi _0655_ (
        .a(new_Jinkela_wire_1469),
        .b(_0143_),
        .c(new_net_14)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    and_bi _0656_ (
        .a(new_Jinkela_wire_980),
        .b(new_Jinkela_wire_1979),
        .c(_0144_)
    );

    spl2 new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_1041),
        .c(new_Jinkela_wire_1042),
        .b(new_Jinkela_wire_1043)
    );

    and_bi _0657_ (
        .a(new_Jinkela_wire_1130),
        .b(new_Jinkela_wire_1941),
        .c(_0145_)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    and_bi _0658_ (
        .a(_0144_),
        .b(_0145_),
        .c(_0146_)
    );

    and_bi _0659_ (
        .a(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_2511),
        .c(_0147_)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_1059),
        .dout(new_Jinkela_wire_1060)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1022),
        .dout(new_Jinkela_wire_1023)
    );

    and_bi _0660_ (
        .a(new_Jinkela_wire_551),
        .b(new_Jinkela_wire_1844),
        .c(_0148_)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    or_bb _0661_ (
        .a(_0148_),
        .b(_0147_),
        .c(_0149_)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1023),
        .dout(new_Jinkela_wire_1024)
    );

    and_bi _0662_ (
        .a(_0146_),
        .b(_0149_),
        .c(_0150_)
    );

    or_bb _0663_ (
        .a(new_Jinkela_wire_1655),
        .b(new_Jinkela_wire_2578),
        .c(_0151_)
    );

    bfr new_Jinkela_buffer_835 (
        .din(G93),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    and_bi _0664_ (
        .a(new_Jinkela_wire_2577),
        .b(new_Jinkela_wire_1653),
        .c(_0152_)
    );

    and_bi _0665_ (
        .a(_0151_),
        .b(_0152_),
        .c(_0153_)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_1060),
        .dout(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    or_bb _0666_ (
        .a(new_Jinkela_wire_1704),
        .b(new_Jinkela_wire_1758),
        .c(_0154_)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1044),
        .dout(new_Jinkela_wire_1045)
    );

    and_bi _0667_ (
        .a(new_Jinkela_wire_1705),
        .b(new_Jinkela_wire_1759),
        .c(_0155_)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    and_bi _0668_ (
        .a(_0154_),
        .b(_0155_),
        .c(_0156_)
    );

    and_bi _0669_ (
        .a(new_Jinkela_wire_1080),
        .b(new_Jinkela_wire_1851),
        .c(_0157_)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1075),
        .dout(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1045),
        .dout(new_Jinkela_wire_1046)
    );

    and_bi _0670_ (
        .a(new_Jinkela_wire_88),
        .b(new_Jinkela_wire_1939),
        .c(_0158_)
    );

    and_bi _0671_ (
        .a(_0157_),
        .b(_0158_),
        .c(_0159_)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1046),
        .dout(new_Jinkela_wire_1047)
    );

    and_bi _0672_ (
        .a(new_Jinkela_wire_652),
        .b(new_Jinkela_wire_2502),
        .c(_0160_)
    );

    bfr new_Jinkela_buffer_839 (
        .din(G101),
        .dout(new_Jinkela_wire_1081)
    );

    and_bi _0673_ (
        .a(new_Jinkela_wire_517),
        .b(new_Jinkela_wire_1984),
        .c(_0161_)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1062),
        .dout(new_Jinkela_wire_1063)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1047),
        .dout(new_Jinkela_wire_1048)
    );

    or_bb _0674_ (
        .a(_0161_),
        .b(_0160_),
        .c(_0162_)
    );

    and_bi _0675_ (
        .a(_0159_),
        .b(_0162_),
        .c(_0163_)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_1061),
        .dout(new_Jinkela_wire_1062)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1048),
        .dout(new_Jinkela_wire_1049)
    );

    and_bi _0676_ (
        .a(new_Jinkela_wire_341),
        .b(new_Jinkela_wire_1978),
        .c(_0164_)
    );

    and_bi _0677_ (
        .a(new_Jinkela_wire_1277),
        .b(new_Jinkela_wire_1940),
        .c(_0165_)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    and_bi _0678_ (
        .a(_0164_),
        .b(_0165_),
        .c(_0166_)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    and_bi _0679_ (
        .a(new_Jinkela_wire_331),
        .b(new_Jinkela_wire_2512),
        .c(_0167_)
    );

    spl3L new_Jinkela_splitter_85 (
        .a(G125),
        .c(new_Jinkela_wire_1085),
        .b(new_Jinkela_wire_1086),
        .d(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_854 (
        .din(G69),
        .dout(new_Jinkela_wire_1103)
    );

    and_bi _0680_ (
        .a(new_Jinkela_wire_608),
        .b(new_Jinkela_wire_1846),
        .c(_0168_)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    or_bb _0681_ (
        .a(_0168_),
        .b(_0167_),
        .c(_0169_)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    and_bi _0682_ (
        .a(_0166_),
        .b(_0169_),
        .c(_0170_)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    and_bi _0683_ (
        .a(new_Jinkela_wire_2154),
        .b(new_Jinkela_wire_1971),
        .c(_0171_)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    and_bi _0684_ (
        .a(new_Jinkela_wire_2153),
        .b(new_Jinkela_wire_1966),
        .c(_0172_)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    and_bi _0685_ (
        .a(_0171_),
        .b(_0172_),
        .c(_0173_)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    and_bi _0686_ (
        .a(new_Jinkela_wire_547),
        .b(new_Jinkela_wire_1985),
        .c(_0174_)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    and_bi _0687_ (
        .a(new_Jinkela_wire_242),
        .b(new_Jinkela_wire_1847),
        .c(_0175_)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    and_bi _0688_ (
        .a(_0174_),
        .b(_0175_),
        .c(_0176_)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1068),
        .dout(new_Jinkela_wire_1069)
    );

    and_bi _0689_ (
        .a(new_Jinkela_wire_555),
        .b(new_Jinkela_wire_1931),
        .c(_0177_)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    and_bi _0690_ (
        .a(new_Jinkela_wire_1109),
        .b(new_Jinkela_wire_2510),
        .c(_0178_)
    );

    spl3L new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_1069),
        .c(new_Jinkela_wire_1070),
        .b(new_Jinkela_wire_1071),
        .d(new_Jinkela_wire_1072)
    );

    or_bb _0691_ (
        .a(_0178_),
        .b(_0177_),
        .c(_0179_)
    );

    bfr new_Jinkela_buffer_857 (
        .din(G114),
        .dout(new_Jinkela_wire_1106)
    );

    and_bi _0692_ (
        .a(_0176_),
        .b(_0179_),
        .c(_0180_)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    and_bi _0693_ (
        .a(new_Jinkela_wire_955),
        .b(new_Jinkela_wire_1975),
        .c(_0181_)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1087),
        .dout(new_Jinkela_wire_1088)
    );

    spl3L new_Jinkela_splitter_88 (
        .a(G139),
        .c(new_Jinkela_wire_1110),
        .b(new_Jinkela_wire_1111),
        .d(new_Jinkela_wire_1112)
    );

    and_bi _0694_ (
        .a(new_Jinkela_wire_1084),
        .b(new_Jinkela_wire_1938),
        .c(_0182_)
    );

    and_bi _0695_ (
        .a(_0181_),
        .b(_0182_),
        .c(_0183_)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_1892),
        .dout(new_Jinkela_wire_1893)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_1870),
        .dout(new_Jinkela_wire_1871)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(new_Jinkela_wire_1838),
        .dout(new_Jinkela_wire_1839)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_1897),
        .dout(new_Jinkela_wire_1898)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_1871),
        .dout(new_Jinkela_wire_1872)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_1893),
        .dout(new_Jinkela_wire_1894)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(new_Jinkela_wire_1872),
        .dout(new_Jinkela_wire_1873)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_net_21),
        .dout(new_Jinkela_wire_1913)
    );

    spl2 new_Jinkela_splitter_191 (
        .a(_0446_),
        .c(new_Jinkela_wire_1922),
        .b(new_Jinkela_wire_1923)
    );

    spl3L new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_1873),
        .c(new_Jinkela_wire_1874),
        .b(new_Jinkela_wire_1875),
        .d(new_Jinkela_wire_1876)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_1876),
        .dout(new_Jinkela_wire_1877)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_1877),
        .dout(new_Jinkela_wire_1878)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(_0351_),
        .dout(new_Jinkela_wire_1924)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_1898),
        .dout(new_Jinkela_wire_1899)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_1878),
        .dout(new_Jinkela_wire_1879)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_1913),
        .dout(new_Jinkela_wire_1914)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_1879),
        .dout(new_Jinkela_wire_1880)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_1899),
        .dout(new_Jinkela_wire_1900)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_1880),
        .dout(new_Jinkela_wire_1881)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_1924),
        .dout(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_1881),
        .dout(new_Jinkela_wire_1882)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_1882),
        .dout(new_Jinkela_wire_1883)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_1914),
        .dout(new_Jinkela_wire_1915)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_1883),
        .dout(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(_0203_),
        .dout(new_Jinkela_wire_1942)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_1884),
        .dout(new_Jinkela_wire_1885)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_1885),
        .dout(new_Jinkela_wire_1886)
    );

    spl3L new_Jinkela_splitter_192 (
        .a(_0005_),
        .c(new_Jinkela_wire_1930),
        .b(new_Jinkela_wire_1932),
        .d(new_Jinkela_wire_1937)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_1886),
        .dout(new_Jinkela_wire_1887)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_1915),
        .dout(new_Jinkela_wire_1916)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_1887),
        .dout(new_Jinkela_wire_1888)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(new_Jinkela_wire_1903),
        .dout(new_Jinkela_wire_1904)
    );

    spl2 new_Jinkela_splitter_188 (
        .a(new_Jinkela_wire_1888),
        .c(new_Jinkela_wire_1889),
        .b(new_Jinkela_wire_1890)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(_0271_),
        .c(new_Jinkela_wire_1947),
        .b(new_Jinkela_wire_1948)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_1904),
        .dout(new_Jinkela_wire_1905)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_1916),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_Jinkela_wire_1905),
        .dout(new_Jinkela_wire_1906)
    );

    bfr new_Jinkela_buffer_1987 (
        .din(new_Jinkela_wire_2690),
        .dout(new_Jinkela_wire_2691)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_561),
        .dout(new_Jinkela_wire_562)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    bfr new_Jinkela_buffer_2005 (
        .din(new_Jinkela_wire_2721),
        .dout(new_Jinkela_wire_2722)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_1988 (
        .din(new_Jinkela_wire_2691),
        .dout(new_Jinkela_wire_2692)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_1438),
        .dout(new_Jinkela_wire_1439)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_562),
        .dout(new_Jinkela_wire_563)
    );

    bfr new_Jinkela_buffer_2011 (
        .din(new_Jinkela_wire_2727),
        .dout(new_Jinkela_wire_2728)
    );

    bfr new_Jinkela_buffer_1989 (
        .din(new_Jinkela_wire_2692),
        .dout(new_Jinkela_wire_2693)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(new_net_16),
        .c(new_Jinkela_wire_1459),
        .b(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_142),
        .dout(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_563),
        .dout(new_Jinkela_wire_564)
    );

    bfr new_Jinkela_buffer_2006 (
        .din(new_Jinkela_wire_2722),
        .dout(new_Jinkela_wire_2723)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_1990 (
        .din(new_Jinkela_wire_2693),
        .dout(new_Jinkela_wire_2694)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_447 (
        .din(G54),
        .dout(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_1439),
        .dout(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_1426),
        .dout(new_Jinkela_wire_1427)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_564),
        .dout(new_Jinkela_wire_565)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_166),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_1991 (
        .din(new_Jinkela_wire_2694),
        .dout(new_Jinkela_wire_2695)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(_0140_),
        .dout(new_Jinkela_wire_1454)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_565),
        .dout(new_Jinkela_wire_566)
    );

    bfr new_Jinkela_buffer_2007 (
        .din(new_Jinkela_wire_2723),
        .dout(new_Jinkela_wire_2724)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_1449),
        .dout(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_1992 (
        .din(new_Jinkela_wire_2695),
        .dout(new_Jinkela_wire_2696)
    );

    bfr new_Jinkela_buffer_165 (
        .din(G39),
        .dout(new_Jinkela_wire_236)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_1440),
        .dout(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_145),
        .dout(new_Jinkela_wire_146)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_1428),
        .dout(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_566),
        .dout(new_Jinkela_wire_567)
    );

    bfr new_Jinkela_buffer_2012 (
        .din(new_Jinkela_wire_2728),
        .dout(new_Jinkela_wire_2729)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_167),
        .dout(new_Jinkela_wire_168)
    );

    bfr new_Jinkela_buffer_1993 (
        .din(new_Jinkela_wire_2696),
        .dout(new_Jinkela_wire_2697)
    );

    bfr new_Jinkela_buffer_453 (
        .din(G59),
        .dout(new_Jinkela_wire_599)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_146),
        .dout(new_Jinkela_wire_147)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_567),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_1994 (
        .din(new_Jinkela_wire_2697),
        .dout(new_Jinkela_wire_2698)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_168),
        .dout(new_Jinkela_wire_169)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    spl3L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_568),
        .c(new_Jinkela_wire_569),
        .b(new_Jinkela_wire_570),
        .d(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_2013 (
        .din(new_Jinkela_wire_2729),
        .dout(new_Jinkela_wire_2730)
    );

    bfr new_Jinkela_buffer_1995 (
        .din(new_Jinkela_wire_2698),
        .dout(new_Jinkela_wire_2699)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_593),
        .dout(new_Jinkela_wire_594)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_169),
        .dout(new_Jinkela_wire_170)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_1450),
        .dout(new_Jinkela_wire_1451)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_584),
        .dout(new_Jinkela_wire_585)
    );

    bfr new_Jinkela_buffer_2014 (
        .din(new_Jinkela_wire_2730),
        .dout(new_Jinkela_wire_2731)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_170),
        .dout(new_Jinkela_wire_171)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_168 (
        .din(G94),
        .dout(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_459 (
        .din(G92),
        .dout(new_Jinkela_wire_605)
    );

    bfr new_Jinkela_buffer_2015 (
        .din(new_Jinkela_wire_2731),
        .dout(new_Jinkela_wire_2732)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    spl2 new_Jinkela_splitter_119 (
        .a(new_Jinkela_wire_1451),
        .c(new_Jinkela_wire_1452),
        .b(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_203),
        .dout(new_Jinkela_wire_204)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    bfr new_Jinkela_buffer_2016 (
        .din(new_Jinkela_wire_2732),
        .dout(new_Jinkela_wire_2733)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_172),
        .dout(new_Jinkela_wire_173)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_594),
        .dout(new_Jinkela_wire_595)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(_0114_),
        .dout(new_Jinkela_wire_1466)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(_0141_),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_586),
        .dout(new_Jinkela_wire_587)
    );

    spl2 new_Jinkela_splitter_123 (
        .a(_0402_),
        .c(new_Jinkela_wire_1470),
        .b(new_Jinkela_wire_1471)
    );

    bfr new_Jinkela_buffer_2017 (
        .din(new_Jinkela_wire_2733),
        .dout(new_Jinkela_wire_2734)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_173),
        .dout(new_Jinkela_wire_174)
    );

    spl2 new_Jinkela_splitter_120 (
        .a(new_Jinkela_wire_1456),
        .c(new_Jinkela_wire_1457),
        .b(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_599),
        .dout(new_Jinkela_wire_600)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    bfr new_Jinkela_buffer_2018 (
        .din(new_Jinkela_wire_2734),
        .dout(new_Jinkela_wire_2735)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_595),
        .dout(new_Jinkela_wire_596)
    );

    spl2 new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_1466),
        .c(new_Jinkela_wire_1467),
        .b(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_588),
        .dout(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_2019 (
        .din(new_Jinkela_wire_2735),
        .dout(new_Jinkela_wire_2736)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    bfr new_Jinkela_buffer_463 (
        .din(G72),
        .dout(new_Jinkela_wire_609)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_204),
        .dout(new_Jinkela_wire_205)
    );

    spl3L new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_190),
        .c(new_Jinkela_wire_191),
        .b(new_Jinkela_wire_192),
        .d(new_Jinkela_wire_193)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_589),
        .dout(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_2020 (
        .din(new_Jinkela_wire_2736),
        .dout(new_Jinkela_wire_2737)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_596),
        .dout(new_Jinkela_wire_597)
    );

    spl2 new_Jinkela_splitter_125 (
        .a(_0319_),
        .c(new_Jinkela_wire_1476),
        .b(new_Jinkela_wire_1477)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_193),
        .dout(new_Jinkela_wire_194)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_590),
        .dout(new_Jinkela_wire_591)
    );

    spl2 new_Jinkela_splitter_126 (
        .a(_0315_),
        .c(new_Jinkela_wire_1478),
        .b(new_Jinkela_wire_1479)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_2021 (
        .din(new_Jinkela_wire_2737),
        .dout(new_Jinkela_wire_2738)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_600),
        .dout(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_205),
        .dout(new_Jinkela_wire_206)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_194),
        .dout(new_Jinkela_wire_195)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_1471),
        .dout(new_Jinkela_wire_1472)
    );

    bfr new_Jinkela_buffer_2022 (
        .din(new_Jinkela_wire_2738),
        .dout(new_Jinkela_wire_2739)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_597),
        .dout(new_Jinkela_wire_598)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(_0350_),
        .dout(new_Jinkela_wire_1480)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_195),
        .dout(new_Jinkela_wire_196)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_1472),
        .dout(new_Jinkela_wire_1473)
    );

    bfr new_Jinkela_buffer_2023 (
        .din(new_Jinkela_wire_2739),
        .dout(new_Jinkela_wire_2740)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_215),
        .dout(new_Jinkela_wire_216)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    spl2 new_Jinkela_splitter_128 (
        .a(_0248_),
        .c(new_Jinkela_wire_1498),
        .b(new_Jinkela_wire_1503)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_206),
        .dout(new_Jinkela_wire_207)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_196),
        .dout(new_Jinkela_wire_197)
    );

    bfr new_Jinkela_buffer_466 (
        .din(G79),
        .dout(new_Jinkela_wire_612)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(new_Jinkela_wire_1473),
        .c(new_Jinkela_wire_1474),
        .b(new_Jinkela_wire_1475)
    );

    bfr new_Jinkela_buffer_2024 (
        .din(new_Jinkela_wire_2740),
        .dout(new_Jinkela_wire_2741)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    spl3L new_Jinkela_splitter_133 (
        .a(_0187_),
        .c(new_Jinkela_wire_1516),
        .b(new_Jinkela_wire_1517),
        .d(new_Jinkela_wire_1518)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_213),
        .dout(new_Jinkela_wire_214)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(new_Jinkela_wire_1481),
        .dout(new_Jinkela_wire_1482)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

endmodule
