module c2670(G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G2531, G2532, G2533, G2534, G2535, G2536, G2537, G2538, G2539, G2540, G2541, G2542, G2543, G2544, G2545, G2546, G2547, G2548, G2549, G2550, G2551, G2552, G2553, G2554, G2555, G2556, G2557, G2558, G2559, G2560, G2561, G2562, G2563, G2564, G2565, G2566, G2567, G2568, G2569, G2570, G2571, G2572, G2573, G2574, G2575, G2576, G2577, G2578, G2579, G2580, G2581, G2582, G2583, G2584, G2585, G2586, G2587, G2588, G2589, G2590, G2591, G2592, G2593, G2594, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G52, G53, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99);
	wire new_net_1545;
	wire new_net_2436;
	wire new_net_2739;
	wire new_net_875;
	wire new_net_1060;
	wire new_net_1639;
	wire new_net_1799;
	wire new_net_2482;
	wire new_net_1890;
	wire new_net_2571;
	wire new_net_323;
	wire new_net_152;
	wire new_net_356;
	wire new_net_569;
	wire new_net_730;
	wire new_net_758;
	wire new_net_779;
	wire new_net_884;
	wire new_net_926;
	wire new_net_1191;
	wire new_net_2723;
	wire new_net_906;
	wire new_net_2650;
	wire new_net_776;
	wire new_net_1578;
	wire new_net_1740;
	wire new_net_306;
	wire new_net_411;
	wire new_net_480;
	wire new_net_1367;
	wire new_net_1379;
	wire new_net_1807;
	wire new_net_1819;
	wire new_net_1885;
	wire new_net_1991;
	wire new_net_2044;
	wire new_net_2579;
	wire new_net_1090;
	wire new_net_1548;
	wire new_net_2035;
	wire new_net_2292;
	wire new_net_937;
	wire new_net_1471;
	wire new_net_1513;
	wire new_net_2559;
	wire new_net_807;
	wire new_net_49;
	wire new_net_517;
	wire new_net_223;
	wire new_net_813;
	wire new_net_1292;
	wire new_net_1647;
	wire new_net_1907;
	wire new_net_1968;
	wire new_net_1980;
	wire new_net_2073;
	wire new_net_2683;
	wire new_net_2450;
	wire new_net_2681;
	wire new_net_1484;
	wire new_net_1403;
	wire new_net_2568;
	wire new_net_2494;
	wire new_net_83;
	wire new_net_134;
	wire new_net_605;
	wire new_net_838;
	wire new_net_1010;
	wire new_net_1040;
	wire new_net_1212;
	wire new_net_1489;
	wire new_net_1732;
	wire new_net_1830;
	wire new_net_2243;
	wire _0324_;
	wire new_net_2618;
	wire new_net_1123;
	wire new_net_2543;
	wire new_net_2172;
	wire new_net_2465;
	wire new_net_2432;
	wire _0365_;
	wire new_net_1297;
	wire new_net_570;
	wire new_net_732;
	wire new_net_687;
	wire new_net_273;
	wire new_net_621;
	wire new_net_357;
	wire new_net_853;
	wire new_net_895;
	wire new_net_916;
	wire new_net_961;
	wire new_net_2438;
	wire new_net_869;
	wire _0406_;
	wire new_net_1062;
	wire _0399_;
	wire new_net_1439;
	wire new_net_2792;
	wire _0423_;
	wire new_net_456;
	wire new_net_100;
	wire new_net_307;
	wire new_net_391;
	wire new_net_412;
	wire new_net_481;
	wire new_net_1102;
	wire new_net_1111;
	wire new_net_1130;
	wire new_net_1260;
	wire new_net_1275;
	wire new_net_1211;
	wire new_net_1895;
	wire new_net_1406;
	wire new_net_2763;
	wire new_net_2315;
	wire new_net_2275;
	wire new_net_2728;
	wire new_net_1148;
	wire new_net_682;
	wire new_net_50;
	wire new_net_518;
	wire new_net_1195;
	wire new_net_1228;
	wire new_net_1348;
	wire new_net_1396;
	wire new_net_1410;
	wire new_net_1422;
	wire new_net_1585;
	wire new_net_1993;
	wire new_net_2361;
	wire new_net_1915;
	wire new_net_2297;
	wire new_net_2224;
	wire new_net_84;
	wire new_net_135;
	wire new_net_153;
	wire new_net_324;
	wire new_net_606;
	wire new_net_654;
	wire new_net_1233;
	wire new_net_1291;
	wire new_net_1324;
	wire new_net_1518;
	wire new_net_2376;
	wire new_net_2641;
	wire new_net_2268;
	wire new_net_2610;
	wire new_net_2455;
	wire new_net_1009;
	wire new_net_2690;
	wire new_net_622;
	wire new_net_652;
	wire new_net_651;
	wire new_net_274;
	wire new_net_759;
	wire new_net_780;
	wire new_net_885;
	wire new_net_927;
	wire new_net_1298;
	wire new_net_1368;
	wire new_net_2099;
	wire new_net_2428;
	wire new_net_2731;
	wire new_net_2623;
	wire new_net_1504;
	wire new_net_2588;
	wire new_net_1127;
	wire new_net_1711;
	wire new_net_101;
	wire new_net_224;
	wire new_net_739;
	wire new_net_392;
	wire new_net_992;
	wire new_net_1427;
	wire new_net_1648;
	wire new_net_1908;
	wire new_net_1981;
	wire new_net_2067;
	wire new_net_1305;
	wire new_net_2369;
	wire new_net_2146;
	wire new_net_2256;
	wire new_net_1071;
	wire new_net_1605;
	wire new_net_51;
	wire new_net_1041;
	wire new_net_1213;
	wire new_net_1309;
	wire new_net_1490;
	wire new_net_1733;
	wire new_net_1831;
	wire new_net_1843;
	wire new_net_1875;
	wire new_net_2311;
	wire new_net_772;
	wire new_net_2309;
	wire _0447_;
	wire new_net_2386;
	wire new_net_1287;
	wire new_net_2355;
	wire new_net_2065;
	wire new_net_2322;
	wire _0464_;
	wire new_net_214;
	wire new_net_2063;
	wire new_net_2320;
	wire _0488_;
	wire new_net_85;
	wire new_net_136;
	wire new_net_154;
	wire new_net_325;
	wire new_net_358;
	wire new_net_571;
	wire new_net_979;
	wire new_net_1671;
	wire new_net_1825;
	wire new_net_1919;
	wire new_net_2507;
	wire new_net_803;
	wire new_net_1155;
	wire new_net_1590;
	wire new_net_2220;
	wire new_net_1998;
	wire new_net_1922;
	wire new_net_1956;
	wire new_net_2405;
	wire new_net_413;
	wire new_net_482;
	wire new_net_854;
	wire new_net_896;
	wire new_net_917;
	wire new_net_1103;
	wire new_net_1112;
	wire new_net_1131;
	wire new_net_1261;
	wire new_net_1276;
	wire new_net_1724;
	wire new_net_1924;
	wire new_net_2264;
	wire new_net_2754;
	wire new_net_1524;
	wire new_net_1693;
	wire new_net_1281;
	wire new_net_1522;
	wire new_net_834;
	wire new_net_2160;
	wire new_net_2420;
	wire new_net_2646;
	wire new_net_2095;
	wire new_net_2202;
	wire new_net_1978;
	wire new_net_225;
	wire new_net_309;
	wire new_net_393;
	wire new_net_519;
	wire new_net_1179;
	wire new_net_1196;
	wire new_net_1349;
	wire new_net_1397;
	wire new_net_1411;
	wire _0040_;
	wire new_net_1616;
	wire new_net_1777;
	wire new_net_2802;
	wire _0325_;
	wire new_net_2584;
	wire new_net_2365;
	wire _0366_;
	wire new_net_865;
	wire new_net_2740;
	wire new_net_607;
	wire new_net_722;
	wire new_net_998;
	wire new_net_1234;
	wire new_net_1267;
	wire new_net_1325;
	wire new_net_1755;
	wire new_net_1853;
	wire new_net_1940;
	wire new_net_1509;
	wire new_net_2142;
	wire new_net_2252;
	wire new_net_1716;
	wire new_net_2006;
	wire _0407_;
	wire new_net_1337;
	wire new_net_1558;
	wire new_net_1964;
	wire new_net_2188;
	wire new_net_1810;
	wire _0424_;
	wire new_net_1768;
	wire new_net_623;
	wire new_net_572;
	wire new_net_86;
	wire new_net_137;
	wire new_net_275;
	wire new_net_359;
	wire new_net_1369;
	wire new_net_1453;
	wire new_net_1809;
	wire new_net_1610;
	wire new_net_1069;
	wire new_net_1344;
	wire new_net_1038;
	wire new_net_2490;
	wire new_net_1118;
	wire new_net_2766;
	wire new_net_414;
	wire new_net_483;
	wire new_net_102;
	wire new_net_760;
	wire new_net_781;
	wire new_net_886;
	wire new_net_928;
	wire new_net_1381;
	wire new_net_1649;
	wire new_net_1909;
	wire new_net_2327;
	wire new_net_2592;
	wire new_net_2512;
	wire new_net_797;
	wire new_net_1597;
	wire new_net_2260;
	wire new_net_2525;
	wire new_net_52;
	wire new_net_394;
	wire new_net_520;
	wire new_net_727;
	wire new_net_1042;
	wire new_net_1491;
	wire new_net_1734;
	wire new_net_1832;
	wire new_net_1844;
	wire new_net_2613;
	wire new_net_1479;
	wire new_net_954;
	wire _0285_;
	wire new_net_2342;
	wire new_net_2154;
	wire new_net_2414;
	wire new_net_959;
	wire new_net_2351;
	wire new_net_127;
	wire new_net_828;
	wire new_net_1529;
	wire new_net_1698;
	wire new_net_2759;
	wire new_net_2719;
	wire new_net_326;
	wire new_net_608;
	wire new_net_155;
	wire new_net_963;
	wire new_net_980;
	wire new_net_1027;
	wire new_net_1615;
	wire new_net_1672;
	wire new_net_1920;
	wire new_net_2345;
	wire new_net_1745;
	wire new_net_2207;
	wire new_net_1628;
	wire new_net_1789;
	wire new_net_2471;
	wire new_net_2774;
	wire new_net_1621;
	wire new_net_1782;
	wire new_net_2213;
	wire new_net_87;
	wire new_net_138;
	wire new_net_276;
	wire new_net_360;
	wire new_net_573;
	wire new_net_624;
	wire new_net_1104;
	wire new_net_1113;
	wire new_net_1132;
	wire new_net_1277;
	wire new_net_2745;
	wire new_net_2114;
	wire new_net_1272;
	wire _0122_;
	wire new_net_1685;
	wire new_net_11;
	wire new_net_2193;
	wire new_net_2486;
	wire new_net_1563;
	wire new_net_484;
	wire new_net_103;
	wire new_net_226;
	wire new_net_855;
	wire new_net_897;
	wire new_net_918;
	wire new_net_1197;
	wire new_net_1350;
	wire new_net_1412;
	wire new_net_1424;
	wire _0163_;
	wire _0448_;
	wire new_net_1458;
	wire new_net_1737;
	wire new_net_1079;
	wire new_net_1820;
	wire new_net_2694;
	wire _0465_;
	wire new_net_1867;
	wire new_net_2548;
	wire new_net_638;
	wire new_net_53;
	wire _0489_;
	wire new_net_395;
	wire new_net_521;
	wire new_net_1240;
	wire new_net_1326;
	wire new_net_1495;
	wire new_net_1756;
	wire new_net_1854;
	wire new_net_915;
	wire new_net_1464;
	wire new_net_1323;
	wire new_net_1753;
	wire new_net_2665;
	wire new_net_1549;
	wire new_net_2332;
	wire new_net_2514;
	wire new_net_1837;
	wire new_net_2373;
	wire new_net_327;
	wire new_net_156;
	wire new_net_506;
	wire new_net_248;
	wire new_net_717;
	wire new_net_1031;
	wire new_net_1370;
	wire new_net_1167;
	wire new_net_1390;
	wire new_net_1602;
	wire new_net_2150;
	wire new_net_2338;
	wire new_net_257;
	wire new_net_2319;
	wire new_net_2347;
	wire new_net_1003;
	wire new_net_2523;
	wire new_net_1248;
	wire new_net_2605;
	wire new_net_1900;
	wire new_net_139;
	wire new_net_664;
	wire new_net_361;
	wire new_net_415;
	wire new_net_625;
	wire new_net_679;
	wire new_net_1092;
	wire new_net_1536;
	wire new_net_1650;
	wire new_net_1910;
	wire new_net_1534;
	wire new_net_1703;
	wire _0326_;
	wire new_net_1946;
	wire new_net_553;
	wire new_net_268;
	wire _0058_;
	wire new_net_1708;
	wire _0367_;
	wire new_net_2178;
	wire new_net_227;
	wire new_net_485;
	wire new_net_761;
	wire new_net_782;
	wire new_net_887;
	wire new_net_929;
	wire new_net_1043;
	wire new_net_1241;
	wire new_net_1466;
	wire new_net_1633;
	wire new_net_2010;
	wire new_net_2476;
	wire new_net_2045;
	wire _0384_;
	wire new_net_1884;
	wire _0408_;
	wire new_net_1237;
	wire new_net_2442;
	wire new_net_2750;
	wire _0425_;
	wire new_net_457;
	wire new_net_396;
	wire new_net_522;
	wire new_net_690;
	wire new_net_609;
	wire new_net_1391;
	wire new_net_1673;
	wire new_net_1921;
	wire new_net_2054;
	wire new_net_466;
	wire new_net_2233;
	wire new_net_1106;
	wire new_net_1570;
	wire new_net_2383;
	wire new_net_1568;
	wire new_net_2798;
	wire new_net_1081;
	wire new_net_2281;
	wire new_net_277;
	wire new_net_88;
	wire new_net_750;
	wire new_net_744;
	wire new_net_574;
	wire new_net_751;
	wire new_net_1093;
	wire new_net_1105;
	wire new_net_1114;
	wire new_net_1133;
	wire new_net_2029;
	wire new_net_2136;
	wire new_net_793;
	wire new_net_2703;
	wire new_net_2553;
	wire new_net_1231;
	wire new_net_2402;
	wire new_net_1023;
	wire new_net_2672;
	wire new_net_2670;
	wire new_net_1554;
	wire new_net_104;
	wire new_net_140;
	wire new_net_362;
	wire new_net_416;
	wire new_net_626;
	wire new_net_997;
	wire new_net_1198;
	wire new_net_1351;
	wire new_net_1366;
	wire new_net_1413;
	wire new_net_1925;
	wire new_net_2519;
	wire new_net_2711;
	wire new_net_1430;
	wire new_net_824;
	wire new_net_1449;
	wire new_net_2122;
	wire new_net_2380;
	wire new_net_2535;
	wire new_net_2090;
	wire new_net_1253;
	wire new_net_54;
	wire new_net_228;
	wire new_net_486;
	wire new_net_856;
	wire new_net_898;
	wire new_net_919;
	wire new_net_1327;
	wire new_net_1757;
	wire new_net_1855;
	wire new_net_1658;
	wire new_net_1416;
	wire new_net_1705;
	wire new_net_849;
	wire new_net_1541;
	wire new_net_2139;
	wire new_net_2249;
	wire new_net_2735;
	wire new_net_610;
	wire new_net_657;
	wire new_net_157;
	wire new_net_328;
	wire new_net_397;
	wire new_net_523;
	wire new_net_995;
	wire new_net_1056;
	wire new_net_1371;
	wire _0082_;
	wire new_net_1709;
	wire new_net_173;
	wire _0099_;
	wire new_net_1886;
	wire new_net_2302;
	wire new_net_880;
	wire new_net_2633;
	wire new_net_2050;
	wire new_net_726;
	wire new_net_575;
	wire new_net_89;
	wire new_net_745;
	wire new_net_981;
	wire new_net_1651;
	wire new_net_1911;
	wire new_net_1984;
	wire new_net_2103;
	wire new_net_2141;
	wire new_net_1689;
	wire new_net_2447;
	wire new_net_2056;
	wire _0164_;
	wire new_net_2013;
	wire new_net_1983;
	wire _0449_;
	wire new_net_1316;
	wire new_net_1575;
	wire _0466_;
	wire new_net_215;
	wire new_net_911;
	wire new_net_2655;
	wire new_net_0;
	wire new_net_105;
	wire new_net_141;
	wire new_net_312;
	wire new_net_627;
	wire _0490_;
	wire new_net_1032;
	wire new_net_1044;
	wire new_net_1214;
	wire new_net_1242;
	wire new_net_2359;
	wire new_net_1321;
	wire new_net_2286;
	wire new_net_714;
	wire new_net_229;
	wire new_net_487;
	wire new_net_55;
	wire new_net_762;
	wire new_net_783;
	wire new_net_668;
	wire new_net_888;
	wire new_net_930;
	wire new_net_942;
	wire new_net_965;
	wire new_net_2677;
	wire new_net_17;
	wire new_net_1480;
	wire new_net_2564;
	wire new_net_1932;
	wire new_net_2086;
	wire new_net_2789;
	wire new_net_386;
	wire new_net_818;
	wire new_net_158;
	wire new_net_329;
	wire new_net_398;
	wire new_net_678;
	wire new_net_996;
	wire new_net_1094;
	wire new_net_1115;
	wire new_net_1134;
	wire new_net_1279;
	wire new_net_1444;
	wire new_net_2391;
	wire _0042_;
	wire new_net_2539;
	wire new_net_1258;
	wire _0327_;
	wire new_net_2168;
	wire new_net_2461;
	wire new_net_2499;
	wire new_net_2248;
	wire _0344_;
	wire new_net_1546;
	wire new_net_90;
	wire new_net_417;
	wire new_net_363;
	wire _0368_;
	wire new_net_576;
	wire new_net_752;
	wire new_net_1199;
	wire new_net_1352;
	wire new_net_1399;
	wire new_net_1414;
	wire new_net_2437;
	wire new_net_670;
	wire _0385_;
	wire new_net_1435;
	wire new_net_1640;
	wire new_net_1800;
	wire _0409_;
	wire new_net_2483;
	wire new_net_2698;
	wire new_net_1643;
	wire new_net_142;
	wire _0426_;
	wire new_net_313;
	wire new_net_716;
	wire new_net_1215;
	wire new_net_1328;
	wire new_net_1758;
	wire new_net_1856;
	wire new_net_2077;
	wire new_net_2203;
	wire new_net_2572;
	wire new_net_1654;
	wire new_net_2724;
	wire new_net_2651;
	wire new_net_2236;
	wire new_net_1224;
	wire new_net_1581;
	wire new_net_1988;
	wire new_net_56;
	wire new_net_611;
	wire new_net_12;
	wire new_net_488;
	wire new_net_749;
	wire new_net_857;
	wire new_net_899;
	wire new_net_920;
	wire new_net_988;
	wire new_net_1372;
	wire new_net_1579;
	wire new_net_1741;
	wire new_net_16;
	wire new_net_1091;
	wire new_net_2036;
	wire new_net_2293;
	wire new_net_2596;
	wire new_net_2706;
	wire new_net_2781;
	wire new_net_1514;
	wire new_net_159;
	wire new_net_279;
	wire new_net_399;
	wire new_net_1652;
	wire new_net_1137;
	wire new_net_1985;
	wire new_net_2059;
	wire new_net_2104;
	wire new_net_2560;
	wire new_net_2583;
	wire new_net_2637;
	wire new_net_2785;
	wire new_net_2682;
	wire _0287_;
	wire new_net_2451;
	wire new_net_535;
	wire new_net_128;
	wire new_net_106;
	wire new_net_641;
	wire new_net_418;
	wire new_net_628;
	wire new_net_364;
	wire new_net_1033;
	wire new_net_1045;
	wire new_net_845;
	wire new_net_1243;
	wire new_net_1468;
	wire new_net_1941;
	wire new_net_2495;
	wire new_net_2062;
	wire new_net_30;
	wire new_net_1500;
	wire new_net_1124;
	wire new_net_2544;
	wire new_net_2688;
	wire new_net_1423;
	wire new_net_2173;
	wire new_net_2466;
	wire new_net_1294;
	wire new_net_2433;
	wire new_net_143;
	wire new_net_230;
	wire new_net_982;
	wire new_net_1668;
	wire new_net_1675;
	wire new_net_1923;
	wire new_net_2124;
	wire new_net_2348;
	wire new_net_2367;
	wire new_net_2398;
	wire new_net_876;
	wire new_net_2439;
	wire _0100_;
	wire _0124_;
	wire new_net_593;
	wire new_net_2118;
	wire new_net_191;
	wire new_net_2793;
	wire new_net_57;
	wire new_net_330;
	wire new_net_612;
	wire _0000_;
	wire new_net_65;
	wire new_net_763;
	wire new_net_784;
	wire new_net_889;
	wire new_net_931;
	wire new_net_1095;
	wire _0141_;
	wire new_net_198;
	wire new_net_2795;
	wire _0165_;
	wire new_net_1896;
	wire new_net_1950;
	wire _0450_;
	wire new_net_907;
	wire new_net_2316;
	wire new_net_1821;
	wire new_net_79;
	wire new_net_777;
	wire new_net_2276;
	wire new_net_2503;
	wire new_net_2729;
	wire new_net_685;
	wire _0467_;
	wire new_net_577;
	wire new_net_677;
	wire new_net_91;
	wire new_net_160;
	wire new_net_280;
	wire new_net_400;
	wire new_net_1200;
	wire new_net_1299;
	wire _0491_;
	wire new_net_1307;
	wire new_net_1586;
	wire new_net_1994;
	wire new_net_1918;
	wire new_net_1952;
	wire new_net_2012;
	wire new_net_2362;
	wire new_net_938;
	wire _0001_;
	wire new_net_419;
	wire new_net_629;
	wire new_net_365;
	wire new_net_107;
	wire new_net_314;
	wire new_net_645;
	wire new_net_808;
	wire new_net_1216;
	wire new_net_1329;
	wire new_net_2041;
	wire new_net_2225;
	wire new_net_2298;
	wire new_net_814;
	wire new_net_1400;
	wire new_net_1519;
	wire new_net_2377;
	wire new_net_2642;
	wire new_net_1938;
	wire new_net_2198;
	wire new_net_1974;
	wire new_net_1175;
	wire new_net_2611;
	wire new_net_1936;
	wire new_net_2456;
	wire new_net_144;
	wire new_net_231;
	wire new_net_646;
	wire new_net_489;
	wire new_net_1373;
	wire new_net_1813;
	wire new_net_1879;
	wire new_net_1891;
	wire new_net_1943;
	wire new_net_1997;
	wire new_net_2691;
	wire new_net_2580;
	wire new_net_839;
	wire new_net_2100;
	wire new_net_2429;
	wire new_net_2624;
	wire new_net_1505;
	wire _0002_;
	wire new_net_331;
	wire new_net_753;
	wire new_net_58;
	wire _0369_;
	wire new_net_858;
	wire new_net_900;
	wire new_net_921;
	wire new_net_1128;
	wire new_net_1308;
	wire new_net_1467;
	wire new_net_1712;
	wire new_net_2002;
	wire new_net_2660;
	wire new_net_2370;
	wire new_net_1306;
	wire _0386_;
	wire new_net_870;
	wire new_net_2147;
	wire _0410_;
	wire new_net_1606;
	wire new_net_92;
	wire new_net_281;
	wire new_net_401;
	wire new_net_578;
	wire new_net_1004;
	wire new_net_1011;
	wire new_net_1034;
	wire new_net_1065;
	wire new_net_1300;
	wire new_net_1469;
	wire new_net_2312;
	wire new_net_2021;
	wire new_net_2024;
	wire new_net_2387;
	wire new_net_2356;
	wire new_net_2066;
	wire new_net_2323;
	wire new_net_315;
	wire _0003_;
	wire new_net_420;
	wire new_net_630;
	wire new_net_366;
	wire new_net_967;
	wire new_net_983;
	wire new_net_1676;
	wire new_net_2064;
	wire new_net_2125;
	wire new_net_2321;
	wire new_net_2508;
	wire _0206_;
	wire new_net_2771;
	wire new_net_1264;
	wire new_net_1593;
	wire new_net_1591;
	wire new_net_1999;
	wire new_net_1957;
	wire new_net_145;
	wire new_net_490;
	wire new_net_526;
	wire new_net_713;
	wire new_net_733;
	wire new_net_613;
	wire new_net_950;
	wire new_net_1096;
	wire new_net_1117;
	wire new_net_1136;
	wire new_net_2406;
	wire new_net_1725;
	wire new_net_2081;
	wire _0264_;
	wire new_net_2755;
	wire new_net_1525;
	wire new_net_1694;
	wire new_net_1282;
	wire new_net_2687;
	wire new_net_2647;
	wire new_net_2421;
	wire _0004_;
	wire new_net_681;
	wire new_net_728;
	wire new_net_332;
	wire new_net_161;
	wire new_net_648;
	wire new_net_764;
	wire new_net_785;
	wire new_net_890;
	wire new_net_932;
	wire new_net_946;
	wire new_net_2126;
	wire new_net_1617;
	wire new_net_1778;
	wire new_net_2803;
	wire new_net_696;
	wire new_net_108;
	wire new_net_282;
	wire new_net_402;
	wire new_net_691;
	wire new_net_1217;
	wire new_net_1330;
	wire new_net_1858;
	wire new_net_2143;
	wire new_net_2205;
	wire new_net_2366;
	wire new_net_2741;
	wire _0084_;
	wire new_net_1268;
	wire new_net_2253;
	wire new_net_1510;
	wire new_net_2222;
	wire new_net_2218;
	wire new_net_1717;
	wire new_net_2189;
	wire new_net_1965;
	wire new_net_1559;
	wire _0125_;
	wire new_net_1304;
	wire new_net_1811;
	wire new_net_232;
	wire new_net_421;
	wire _0005_;
	wire new_net_367;
	wire new_net_316;
	wire new_net_631;
	wire new_net_1374;
	wire new_net_1376;
	wire new_net_1814;
	wire new_net_1880;
	wire new_net_2306;
	wire new_net_1454;
	wire new_net_1611;
	wire _0166_;
	wire new_net_773;
	wire new_net_1039;
	wire new_net_1863;
	wire new_net_2060;
	wire _0183_;
	wire new_net_2019;
	wire new_net_614;
	wire new_net_13;
	wire new_net_680;
	wire new_net_146;
	wire new_net_527;
	wire new_net_1263;
	wire new_net_1963;
	wire new_net_1987;
	wire new_net_2106;
	wire new_net_2716;
	wire new_net_2767;
	wire new_net_2661;
	wire new_net_2699;
	wire new_net_2328;
	wire new_net_2760;
	wire new_net_1833;
	wire new_net_804;
	wire new_net_1440;
	wire new_net_2107;
	wire new_net_2334;
	wire new_net_1598;
	wire new_net_333;
	wire _0006_;
	wire new_net_162;
	wire new_net_579;
	wire new_net_754;
	wire new_net_859;
	wire new_net_901;
	wire new_net_922;
	wire new_net_1005;
	wire new_net_1035;
	wire new_net_1161;
	wire new_net_2261;
	wire new_net_2601;
	wire new_net_516;
	wire new_net_948;
	wire new_net_2155;
	wire new_net_2415;
	wire new_net_2092;
	wire new_net_835;
	wire new_net_2352;
	wire new_net_109;
	wire new_net_283;
	wire new_net_403;
	wire new_net_746;
	wire new_net_984;
	wire new_net_1392;
	wire new_net_1530;
	wire new_net_1677;
	wire new_net_1699;
	wire new_net_1913;
	wire new_net_1942;
	wire new_net_1488;
	wire new_net_1903;
	wire _0329_;
	wire new_net_1187;
	wire new_net_1746;
	wire new_net_2208;
	wire new_net_2395;
	wire new_net_1629;
	wire new_net_1790;
	wire new_net_976;
	wire new_net_2472;
	wire new_net_1783;
	wire new_net_2775;
	wire _0346_;
	wire new_net_317;
	wire _0007_;
	wire new_net_738;
	wire new_net_233;
	wire new_net_422;
	wire new_net_491;
	wire new_net_632;
	wire _0370_;
	wire new_net_368;
	wire new_net_866;
	wire new_net_2214;
	wire new_net_2183;
	wire new_net_2746;
	wire new_net_1273;
	wire _0411_;
	wire new_net_60;
	wire new_net_528;
	wire new_net_615;
	wire new_net_1028;
	wire new_net_1202;
	wire new_net_1355;
	wire new_net_1382;
	wire new_net_1417;
	wire new_net_1620;
	wire new_net_1564;
	wire new_net_2194;
	wire new_net_2487;
	wire new_net_1816;
	wire new_net_2576;
	wire new_net_1459;
	wire new_net_2025;
	wire new_net_2132;
	wire new_net_2695;
	wire new_net_580;
	wire _0008_;
	wire new_net_334;
	wire new_net_765;
	wire new_net_786;
	wire new_net_891;
	wire new_net_933;
	wire new_net_1218;
	wire new_net_1331;
	wire new_net_1653;
	wire new_net_2549;
	wire new_net_2589;
	wire new_net_1496;
	wire new_net_2069;
	wire new_net_1019;
	wire new_net_985;
	wire new_net_1754;
	wire new_net_2666;
	wire new_net_1550;
	wire new_net_798;
	wire new_net_2515;
	wire new_net_1838;
	wire new_net_1362;
	wire new_net_404;
	wire new_net_695;
	wire new_net_1046;
	wire _0248_;
	wire new_net_1236;
	wire new_net_1375;
	wire new_net_1576;
	wire new_net_1815;
	wire new_net_1881;
	wire new_net_1893;
	wire new_net_2374;
	wire new_net_1445;
	wire new_net_2339;
	wire new_net_1603;
	wire new_net_2411;
	wire new_net_999;
	wire new_net_2531;
	wire new_net_2524;
	wire new_net_22;
	wire new_net_536;
	wire new_net_1249;
	wire new_net_1901;
	wire new_net_423;
	wire new_net_492;
	wire new_net_633;
	wire new_net_369;
	wire _0009_;
	wire new_net_318;
	wire _0306_;
	wire new_net_147;
	wire new_net_24;
	wire new_net_829;
	wire new_net_2537;
	wire new_net_1537;
	wire new_net_2424;
	wire new_net_1947;
	wire new_net_1052;
	wire new_net_2;
	wire new_net_163;
	wire new_net_616;
	wire new_net_1006;
	wire new_net_1012;
	wire new_net_1029;
	wire new_net_1036;
	wire new_net_1302;
	wire new_net_1320;
	wire new_net_1826;
	wire new_net_1634;
	wire new_net_2477;
	wire new_net_2629;
	wire new_net_2046;
	wire new_net_587;
	wire new_net_2443;
	wire _0126_;
	wire new_net_1;
	wire new_net_639;
	wire _0010_;
	wire new_net_110;
	wire new_net_581;
	wire new_net_755;
	wire new_net_860;
	wire new_net_902;
	wire new_net_923;
	wire new_net_66;
	wire new_net_769;
	wire new_net_2011;
	wire new_net_2269;
	wire new_net_2055;
	wire new_net_2384;
	wire new_net_1571;
	wire _0167_;
	wire new_net_1569;
	wire _0184_;
	wire new_net_234;
	wire new_net_405;
	wire new_net_683;
	wire new_net_1098;
	wire _0469_;
	wire new_net_1107;
	wire new_net_1119;
	wire new_net_1138;
	wire new_net_1289;
	wire new_net_1150;
	wire new_net_2282;
	wire _0493_;
	wire new_net_800;
	wire new_net_2704;
	wire new_net_1873;
	wire new_net_2554;
	wire new_net_709;
	wire new_net_243;
	wire new_net_2673;
	wire new_net_1678;
	wire new_net_61;
	wire new_net_529;
	wire new_net_370;
	wire _0011_;
	wire new_net_493;
	wire new_net_319;
	wire new_net_634;
	wire new_net_148;
	wire new_net_1203;
	wire new_net_1356;
	wire new_net_1555;
	wire new_net_1845;
	wire new_net_1928;
	wire new_net_508;
	wire new_net_2520;
	wire new_net_1926;
	wire new_net_2712;
	wire new_net_259;
	wire new_net_2684;
	wire new_net_1401;
	wire new_net_1729;
	wire new_net_2536;
	wire new_net_164;
	wire new_net_335;
	wire new_net_644;
	wire new_net_1219;
	wire new_net_1332;
	wire new_net_1345;
	wire new_net_1860;
	wire new_net_1859;
	wire new_net_1935;
	wire new_net_1254;
	wire new_net_2615;
	wire new_net_973;
	wire _0330_;
	wire new_net_1706;
	wire new_net_291;
	wire new_net_555;
	wire new_net_1542;
	wire _0062_;
	wire new_net_111;
	wire new_net_582;
	wire _0347_;
	wire _0012_;
	wire new_net_285;
	wire new_net_562;
	wire new_net_766;
	wire new_net_787;
	wire new_net_892;
	wire new_net_934;
	wire _0371_;
	wire new_net_1232;
	wire _0388_;
	wire new_net_41;
	wire _0412_;
	wire new_net_1887;
	wire new_net_2303;
	wire new_net_235;
	wire new_net_406;
	wire new_net_424;
	wire new_net_675;
	wire new_net_1244;
	wire new_net_1295;
	wire new_net_1644;
	wire new_net_1761;
	wire new_net_1804;
	wire new_net_1933;
	wire _0429_;
	wire new_net_2720;
	wire _0473_;
	wire new_net_1690;
	wire new_net_2057;
	wire new_net_1144;
	wire new_net_2527;
	wire new_net_1317;
	wire new_net_2764;
	wire new_net_14;
	wire new_net_494;
	wire new_net_635;
	wire new_net_689;
	wire new_net_62;
	wire new_net_530;
	wire _0013_;
	wire new_net_617;
	wire new_net_1007;
	wire new_net_1030;
	wire new_net_2656;
	wire new_net_1087;
	wire new_net_794;
	wire new_net_1048;
	wire new_net_2287;
	wire new_net_2074;
	wire new_net_723;
	wire new_net_96;
	wire new_net_165;
	wire new_net_647;
	wire new_net_684;
	wire new_net_729;
	wire new_net_986;
	wire new_net_1238;
	wire new_net_1313;
	wire new_net_1655;
	wire new_net_2678;
	wire new_net_2565;
	wire new_net_2087;
	wire _0290_;
	wire new_net_825;
	wire new_net_1431;
	wire new_net_2790;
	wire new_net_2491;
	wire new_net_2717;
	wire new_net_286;
	wire new_net_583;
	wire _0014_;
	wire new_net_756;
	wire new_net_861;
	wire new_net_903;
	wire _0307_;
	wire new_net_924;
	wire new_net_1013;
	wire new_net_1099;
	wire new_net_2392;
	wire new_net_2540;
	wire new_net_1259;
	wire new_net_2169;
	wire new_net_2462;
	wire new_net_2500;
	wire new_net_850;
	wire new_net_1664;
	wire new_net_236;
	wire new_net_371;
	wire new_net_407;
	wire new_net_425;
	wire new_net_1204;
	wire new_net_1296;
	wire new_net_1357;
	wire new_net_1394;
	wire new_net_1419;
	wire new_net_1622;
	wire new_net_2657;
	wire new_net_1301;
	wire new_net_1641;
	wire new_net_1801;
	wire new_net_2257;
	wire new_net_2484;
	wire new_net_700;
	wire new_net_881;
	wire new_net_531;
	wire new_net_618;
	wire new_net_636;
	wire _0015_;
	wire new_net_1220;
	wire new_net_1333;
	wire new_net_1849;
	wire new_net_731;
	wire new_net_1861;
	wire new_net_1812;
	wire new_net_1892;
	wire new_net_2573;
	wire _0168_;
	wire new_net_2272;
	wire new_net_2725;
	wire _0453_;
	wire new_net_2652;
	wire new_net_2237;
	wire new_net_97;
	wire new_net_112;
	wire new_net_166;
	wire _0185_;
	wire new_net_1377;
	wire new_net_1520;
	wire new_net_1582;
	wire _0470_;
	wire new_net_217;
	wire new_net_912;
	wire new_net_1989;
	wire new_net_1315;
	wire new_net_1580;
	wire new_net_1742;
	wire _0494_;
	wire new_net_2037;
	wire new_net_2294;
	wire new_net_1473;
	wire new_net_287;
	wire _0016_;
	wire new_net_767;
	wire new_net_374;
	wire new_net_788;
	wire new_net_893;
	wire new_net_935;
	wire new_net_1393;
	wire new_net_1645;
	wire new_net_1762;
	wire new_net_1515;
	wire new_net_2561;
	wire new_net_2083;
	wire new_net_2638;
	wire new_net_943;
	wire new_net_2786;
	wire new_net_1970;
	wire new_net_2265;
	wire new_net_2452;
	wire new_net_819;
	wire new_net_63;
	wire new_net_150;
	wire new_net_237;
	wire new_net_321;
	wire new_net_372;
	wire new_net_408;
	wire new_net_426;
	wire new_net_495;
	wire new_net_697;
	wire new_net_1008;
	wire new_net_2161;
	wire new_net_2096;
	wire new_net_2496;
	wire new_net_2245;
	wire new_net_2336;
	wire _0331_;
	wire new_net_2192;
	wire new_net_2620;
	wire new_net_1501;
	wire new_net_2585;
	wire new_net_1125;
	wire _0063_;
	wire new_net_2545;
	wire new_net_532;
	wire new_net_337;
	wire _0017_;
	wire _0348_;
	wire new_net_987;
	wire new_net_1239;
	wire new_net_1341;
	wire new_net_1656;
	wire new_net_1680;
	wire new_net_1916;
	wire new_net_2174;
	wire new_net_2434;
	wire _0372_;
	wire new_net_435;
	wire new_net_2779;
	wire new_net_33;
	wire _0389_;
	wire new_net_442;
	wire new_net_710;
	wire _0413_;
	wire new_net_584;
	wire new_net_113;
	wire new_net_167;
	wire new_net_1014;
	wire new_net_1100;
	wire new_net_1109;
	wire new_net_1140;
	wire new_net_1246;
	wire new_net_1314;
	wire new_net_1450;
	wire new_net_2119;
	wire new_net_2794;
	wire _0430_;
	wire new_net_1108;
	wire new_net_1245;
	wire new_net_2130;
	wire new_net_1408;
	wire new_net_474;
	wire new_net_2317;
	wire new_net_2109;
	wire _0018_;
	wire new_net_288;
	wire new_net_757;
	wire new_net_862;
	wire new_net_904;
	wire new_net_925;
	wire new_net_1310;
	wire new_net_1358;
	wire new_net_1420;
	wire new_net_790;
	wire new_net_1822;
	wire new_net_2504;
	wire new_net_1230;
	wire new_net_1587;
	wire new_net_2593;
	wire new_net_1995;
	wire new_net_1917;
	wire new_net_64;
	wire new_net_238;
	wire new_net_409;
	wire new_net_427;
	wire new_net_659;
	wire new_net_496;
	wire new_net_619;
	wire new_net_1221;
	wire new_net_1322;
	wire new_net_1334;
	wire new_net_2782;
	wire new_net_2042;
	wire new_net_2299;
	wire new_net_2226;
	wire new_net_821;
	wire new_net_2448;
	wire new_net_2751;
	wire new_net_1278;
	wire new_net_2378;
	wire new_net_2643;
	wire new_net_537;
	wire new_net_1939;
	wire new_net_2199;
	wire new_net_2148;
	wire new_net_338;
	wire new_net_721;
	wire new_net_98;
	wire _0019_;
	wire new_net_1176;
	wire new_net_1303;
	wire new_net_1378;
	wire new_net_1720;
	wire new_net_1806;
	wire new_net_130;
	wire new_net_1937;
	wire new_net_2241;
	wire new_net_1774;
	wire new_net_2612;
	wire new_net_25;
	wire new_net_2799;
	wire new_net_846;
	wire new_net_2581;
	wire new_net_585;
	wire new_net_674;
	wire new_net_1646;
	wire new_net_1763;
	wire new_net_1967;
	wire new_net_2072;
	wire new_net_2091;
	wire new_net_2110;
	wire new_net_2310;
	wire new_net_1506;
	wire new_net_2488;
	wire new_net_1129;
	wire new_net_1794;
	wire new_net_1713;
	wire new_net_994;
	wire new_net_877;
	wire new_net_2371;
	wire new_net_2115;
	wire _0104_;
	wire new_net_322;
	wire new_net_736;
	wire new_net_151;
	wire new_net_373;
	wire _0020_;
	wire new_net_595;
	wire new_net_768;
	wire new_net_789;
	wire new_net_894;
	wire new_net_936;
	wire new_net_1073;
	wire new_net_1607;
	wire new_net_67;
	wire new_net_2313;
	wire new_net_2015;
	wire _0454_;
	wire new_net_908;
	wire new_net_2388;
	wire new_net_533;
	wire new_net_620;
	wire new_net_10;
	wire new_net_15;
	wire new_net_239;
	wire new_net_81;
	wire new_net_410;
	wire new_net_428;
	wire new_net_778;
	wire new_net_1395;
	wire _0471_;
	wire new_net_2324;
	wire _0495_;
	wire new_net_1827;
	wire new_net_2509;
	wire new_net_2772;
	wire new_net_1594;
	wire new_net_1157;
	wire new_net_1592;
	wire new_net_2333;
	wire new_net_114;
	wire new_net_99;
	wire new_net_168;
	wire _0021_;
	wire new_net_244;
	wire new_net_939;
	wire new_net_1101;
	wire new_net_1110;
	wire new_net_1141;
	wire new_net_1247;
	wire new_net_2000;
	wire new_net_1697;
	wire new_net_809;
	wire new_net_2407;
	wire new_net_509;
	wire new_net_815;
	wire new_net_1726;
	wire new_net_2082;
	wire new_net_1526;
	wire new_net_1695;
	wire new_net_2606;
	wire new_net_289;
	wire new_net_712;
	wire new_net_1347;
	wire new_net_1421;
	wire new_net_1624;
	wire new_net_1636;
	wire new_net_1710;
	wire new_net_1785;
	wire new_net_1796;
	wire new_net_1927;
	wire new_net_2648;
	wire new_net_2127;
	wire new_net_2204;
	wire new_net_840;
	wire new_net_1181;
	wire new_net_2164;
	wire new_net_1625;
	wire new_net_1786;
	wire new_net_1353;
	wire new_net_1618;
	wire new_net_1779;
	wire _0332_;
	wire new_net_556;
	wire new_net_292;
	wire new_net_2210;
	wire new_net_1876;
	wire _0349_;
	wire _0373_;
	wire new_net_2179;
	wire new_net_2742;
	wire new_net_2144;
	wire new_net_1269;
	wire new_net_2254;
	wire new_net_1511;
	wire _0390_;
	wire new_net_871;
	wire new_net_2008;
	wire _0414_;
	wire new_net_1339;
	wire new_net_1560;
	wire new_net_1966;
	wire new_net_2190;
	wire new_net_1805;
	wire _0022_;
	wire _0064_;
	wire _0106_;
	wire _0190_;
	wire _0232_;
	wire _0274_;
	wire _0148_;
	wire _0316_;
	wire _0358_;
	wire _0400_;
	wire new_net_1455;
	wire new_net_2307;
	wire new_net_1612;
	wire new_net_1770;
	wire new_net_1120;
	wire new_net_2768;
	wire new_net_240;
	wire new_net_655;
	wire new_net_650;
	wire new_net_1470;
	wire new_net_1721;
	wire new_net_1897;
	wire new_net_1949;
	wire new_net_2001;
	wire new_net_2032;
	wire new_net_2289;
	wire new_net_1547;
	wire new_net_2662;
	wire new_net_2329;
	wire _0210_;
	wire new_net_1834;
	wire new_net_2108;
	wire new_net_1441;
	wire new_net_2335;
	wire new_net_1599;
	wire new_net_2078;
	wire _0023_;
	wire _0065_;
	wire _0107_;
	wire _0191_;
	wire _0233_;
	wire _0275_;
	wire _0149_;
	wire _0317_;
	wire _0359_;
	wire _0401_;
	wire new_net_115;
	wire new_net_2344;
	wire new_net_2602;
	wire new_net_2123;
	wire new_net_2156;
	wire new_net_2416;
	wire new_net_842;
	wire new_net_2353;
	wire _0309_;
	wire new_net_2761;
	wire new_net_1531;
	wire new_net_1700;
	wire new_net_206;
	wire new_net_290;
	wire new_net_1164;
	wire new_net_1404;
	wire new_net_2240;
	wire new_net_2502;
	wire new_net_2569;
	wire new_net_1384;
	wire new_net_1747;
	wire new_net_2209;
	wire new_net_2363;
	wire new_net_1630;
	wire new_net_1791;
	wire new_net_2473;
	wire new_net_2776;
	wire new_net_1623;
	wire new_net_1784;
	wire new_net_2140;
	wire new_net_2215;
	wire _0192_;
	wire _0234_;
	wire _0276_;
	wire _0024_;
	wire _0066_;
	wire _0108_;
	wire _0150_;
	wire _0318_;
	wire _0360_;
	wire _0402_;
	wire new_net_2747;
	wire _0105_;
	wire new_net_1274;
	wire new_net_2051;
	wire new_net_2230;
	wire new_net_1687;
	wire new_net_241;
	wire new_net_640;
	wire _0153_;
	wire new_net_969;
	wire new_net_1049;
	wire new_net_1061;
	wire new_net_1070;
	wire new_net_1080;
	wire new_net_1172;
	wire new_net_1184;
	wire new_net_1565;
	wire new_net_1817;
	wire new_net_774;
	wire new_net_2577;
	wire new_net_2278;
	wire new_net_2696;
	wire _0187_;
	wire _0487_;
	wire new_net_554;
	wire _0193_;
	wire _0235_;
	wire _0277_;
	wire _0025_;
	wire _0067_;
	wire _0109_;
	wire _0151_;
	wire _0319_;
	wire new_net_1497;
	wire new_net_1869;
	wire new_net_2550;
	wire new_net_1912;
	wire new_net_2070;
	wire new_net_1674;
	wire new_net_2667;
	wire new_net_805;
	wire new_net_1551;
	wire new_net_2516;
	wire new_net_1839;
	wire new_net_811;
	wire new_net_1201;
	wire new_net_207;
	wire new_net_375;
	wire new_net_1223;
	wire new_net_1336;
	wire new_net_1681;
	wire new_net_1864;
	wire new_net_2022;
	wire new_net_1477;
	wire new_net_2111;
	wire new_net_1446;
	wire new_net_1169;
	wire new_net_2152;
	wire new_net_2412;
	wire new_net_2349;
	wire new_net_836;
	wire new_net_1902;
	wire new_net_970;
	wire _0446_;
	wire _0194_;
	wire _0236_;
	wire _0278_;
	wire _0152_;
	wire _0026_;
	wire _0068_;
	wire _0110_;
	wire _0320_;
	wire _0362_;
	wire new_net_1538;
	wire new_net_2177;
	wire new_net_2425;
	wire _0333_;
	wire new_net_1948;
	wire new_net_2732;
	wire new_net_1958;
	wire new_net_711;
	wire new_net_242;
	wire new_net_1002;
	wire new_net_1604;
	wire _0374_;
	wire new_net_867;
	wire new_net_1635;
	wire new_net_1765;
	wire new_net_1795;
	wire new_net_1969;
	wire new_net_2112;
	wire new_net_2478;
	wire new_net_2047;
	wire _0391_;
	wire _0415_;
	wire new_net_2444;
	wire new_net_117;
	wire new_net_189;
	wire new_net_258;
	wire new_net_465;
	wire _0027_;
	wire _0069_;
	wire _0111_;
	wire _0195_;
	wire _0237_;
	wire _0279_;
	wire new_net_1311;
	wire new_net_1572;
	wire new_net_2231;
	wire new_net_2692;
	wire new_net_1083;
	wire new_net_448;
	wire new_net_208;
	wire new_net_376;
	wire new_net_499;
	wire new_net_989;
	wire new_net_1145;
	wire new_net_1472;
	wire new_net_1659;
	wire new_net_1682;
	wire new_net_2003;
	wire new_net_2031;
	wire new_net_2283;
	wire new_net_2555;
	wire new_net_5;
	wire new_net_799;
	wire new_net_1025;
	wire new_net_1679;
	wire new_net_2597;
	wire new_net_2674;
	wire new_net_725;
	wire _0196_;
	wire _0238_;
	wire _0280_;
	wire _0028_;
	wire _0070_;
	wire _0112_;
	wire _0154_;
	wire _0322_;
	wire _0364_;
	wire new_net_1001;
	wire new_net_1556;
	wire new_net_1929;
	wire new_net_2713;
	wire new_net_1451;
	wire _0310_;
	wire new_net_830;
	wire new_net_1016;
	wire new_net_1383;
	wire new_net_2159;
	wire new_net_26;
	wire new_net_1255;
	wire new_net_2221;
	wire new_net_2458;
	wire new_net_2526;
	wire new_net_2616;
	wire new_net_1660;
	wire new_net_1418;
	wire new_net_1543;
	wire new_net_1387;
	wire new_net_2737;
	wire new_net_34;
	wire new_net_172;
	wire _0029_;
	wire _0071_;
	wire _0113_;
	wire _0155_;
	wire _0239_;
	wire _0281_;
	wire _0197_;
	wire _0323_;
	wire new_net_1058;
	wire new_net_1637;
	wire new_net_1797;
	wire new_net_2440;
	wire new_net_1888;
	wire new_net_2304;
	wire new_net_2635;
	wire new_net_2381;
	wire new_net_596;
	wire new_net_742;
	wire new_net_68;
	wire new_net_209;
	wire new_net_449;
	wire new_net_500;
	wire new_net_701;
	wire new_net_770;
	wire new_net_1481;
	wire new_net_1723;
	wire new_net_1899;
	wire new_net_2721;
	wire _0147_;
	wire new_net_1691;
	wire new_net_2058;
	wire new_net_1318;
	wire new_net_1492;
	wire new_net_2277;
	wire new_net_2730;
	wire new_net_342;
	wire _0492_;
	wire new_net_665;
	wire new_net_432;
	wire _0156_;
	wire _0030_;
	wire _0072_;
	wire _0114_;
	wire _0198_;
	wire _0240_;
	wire new_net_2701;
	wire new_net_801;
	wire new_net_2033;
	wire new_net_2290;
	wire new_net_2288;
	wire new_net_1342;
	wire new_net_118;
	wire new_net_589;
	wire new_net_666;
	wire new_net_715;
	wire new_net_1121;
	wire new_net_1154;
	wire new_net_1166;
	wire new_net_2149;
	wire new_net_2628;
	wire new_net_510;
	wire new_net_2679;
	wire new_net_1482;
	wire new_net_1848;
	wire new_net_2566;
	wire new_net_832;
	wire new_net_2343;
	wire new_net_2791;
	wire new_net_2718;
	wire new_net_2492;
	wire new_net_467;
	wire _0451_;
	wire new_net_706;
	wire _0283_;
	wire _0157_;
	wire _0031_;
	wire _0073_;
	wire _0115_;
	wire _0199_;
	wire _0241_;
	wire new_net_2052;
	wire new_net_1905;
	wire new_net_2393;
	wire new_net_2541;
	wire _0334_;
	wire new_net_2170;
	wire new_net_1346;
	wire new_net_1707;
	wire new_net_2430;
	wire new_net_557;
	wire new_net_2463;
	wire new_net_2501;
	wire new_net_863;
	wire _0351_;
	wire new_net_1751;
	wire new_net_2625;
	wire new_net_69;
	wire new_net_450;
	wire new_net_1051;
	wire new_net_1072;
	wire new_net_1082;
	wire new_net_1149;
	wire _0375_;
	wire new_net_1174;
	wire new_net_1186;
	wire new_net_1250;
	wire _0392_;
	wire new_net_1437;
	wire new_net_1642;
	wire new_net_1802;
	wire _0416_;
	wire new_net_433;
	wire new_net_538;
	wire _0452_;
	wire _0032_;
	wire _0074_;
	wire _0116_;
	wire _0158_;
	wire _0242_;
	wire _0284_;
	wire _0200_;
	wire new_net_2736;
	wire new_net_2273;
	wire new_net_2726;
	wire new_net_2238;
	wire new_net_1226;
	wire new_net_2357;
	wire new_net_1583;
	wire new_net_708;
	wire new_net_734;
	wire new_net_590;
	wire new_net_119;
	wire new_net_260;
	wire new_net_293;
	wire new_net_1015;
	wire new_net_1205;
	wire new_net_1225;
	wire new_net_1338;
	wire new_net_2101;
	wire new_net_795;
	wire new_net_2295;
	wire new_net_1474;
	wire new_net_2708;
	wire new_net_36;
	wire new_net_501;
	wire new_net_378;
	wire new_net_192;
	wire _0075_;
	wire _0033_;
	wire _0117_;
	wire _0159_;
	wire _0201_;
	wire _0243_;
	wire new_net_1139;
	wire new_net_1209;
	wire new_net_116;
	wire new_net_1516;
	wire new_net_2084;
	wire new_net_2639;
	wire new_net_2266;
	wire new_net_2608;
	wire _0294_;
	wire new_net_826;
	wire new_net_2453;
	wire new_net_1283;
	wire new_net_2162;
	wire new_net_656;
	wire new_net_451;
	wire new_net_702;
	wire _0311_;
	wire new_net_1265;
	wire new_net_1385;
	wire new_net_1971;
	wire new_net_2271;
	wire new_net_2619;
	wire new_net_2097;
	wire new_net_2621;
	wire new_net_851;
	wire new_net_1502;
	wire new_net_2586;
	wire new_net_1425;
	wire new_net_990;
	wire _0496_;
	wire new_net_434;
	wire _0034_;
	wire _0076_;
	wire _0118_;
	wire _0160_;
	wire _0202_;
	wire _0244_;
	wire _0286_;
	wire _0328_;
	wire new_net_2780;
	wire new_net_882;
	wire new_net_2570;
	wire new_net_737;
	wire new_net_120;
	wire new_net_174;
	wire new_net_261;
	wire new_net_294;
	wire new_net_468;
	wire new_net_558;
	wire new_net_971;
	wire new_net_991;
	wire new_net_1147;
	wire new_net_2234;
	wire new_net_1077;
	wire new_net_341;
	wire new_net_2061;
	wire new_net_2318;
	wire new_net_1823;
	wire _0189_;
	wire new_net_2505;
	wire new_net_70;
	wire _0455_;
	wire new_net_211;
	wire _0497_;
	wire _0035_;
	wire _0077_;
	wire _0119_;
	wire _0161_;
	wire _0203_;
	wire _0245_;
	wire _0474_;
	wire new_net_348;
	wire new_net_913;
	wire new_net_1588;
	wire new_net_2594;
	wire new_net_1996;
	wire new_net_1954;
	wire new_net_2403;
	wire new_net_502;
	wire new_net_2783;
	wire new_net_1722;
	wire new_net_452;
	wire new_net_1018;
	wire new_net_1142;
	wire new_net_1206;
	wire new_net_1286;
	wire new_net_2223;
	wire new_net_2262;
	wire new_net_2528;
	wire new_net_2043;
	wire new_net_2300;
	wire new_net_251;
	wire new_net_944;
	wire new_net_2227;
	wire new_net_2449;
	wire new_net_2752;
	wire new_net_2158;
	wire new_net_2644;
	wire new_net_2654;
	wire new_net_820;
	wire new_net_2093;
	wire new_net_2200;
	wire new_net_267;
	wire new_net_1976;
	wire new_net_1177;
	wire new_net_540;
	wire _0456_;
	wire _0498_;
	wire _0204_;
	wire _0246_;
	wire _0288_;
	wire _0036_;
	wire _0078_;
	wire _0120_;
	wire _0162_;
	wire new_net_1775;
	wire new_net_2242;
	wire new_net_2800;
	wire new_net_2582;
	wire _0335_;
	wire new_net_2675;
	wire _0352_;
	wire new_net_559;
	wire new_net_673;
	wire new_net_7;
	wire new_net_121;
	wire new_net_175;
	wire new_net_193;
	wire new_net_379;
	wire new_net_469;
	wire new_net_1483;
	wire _0376_;
	wire new_net_1507;
	wire new_net_1714;
	wire new_net_35;
	wire new_net_2004;
	wire new_net_446;
	wire new_net_1335;
	wire new_net_2186;
	wire _0393_;
	wire new_net_1808;
	wire new_net_2116;
	wire _0417_;
	wire new_net_38;
	wire new_net_503;
	wire new_net_71;
	wire _0457_;
	wire _0205_;
	wire _0247_;
	wire _0289_;
	wire _0037_;
	wire _0079_;
	wire _0121_;
	wire _0434_;
	wire new_net_460;
	wire new_net_1067;
	wire new_net_1608;
	wire new_net_1405;
	wire new_net_2314;
	wire new_net_2023;
	wire new_net_2016;
	wire new_net_1116;
	wire new_net_2389;
	wire new_net_476;
	wire new_net_978;
	wire new_net_637;
	wire new_net_1156;
	wire new_net_1168;
	wire new_net_2151;
	wire new_net_2325;
	wire new_net_791;
	wire new_net_2375;
	wire new_net_2394;
	wire new_net_2590;
	wire new_net_2630;
	wire new_net_1828;
	wire new_net_2360;
	wire new_net_2510;
	wire new_net_1595;
	wire new_net_1840;
	wire new_net_2258;
	wire new_net_295;
	wire new_net_436;
	wire new_net_699;
	wire new_net_592;
	wire new_net_262;
	wire new_net_693;
	wire new_net_23;
	wire new_net_541;
	wire _0038_;
	wire _0080_;
	wire new_net_952;
	wire new_net_822;
	wire new_net_2340;
	wire new_net_957;
	wire new_net_2757;
	wire new_net_1527;
	wire new_net_1696;
	wire new_net_539;
	wire new_net_122;
	wire new_net_176;
	wire new_net_194;
	wire new_net_212;
	wire new_net_380;
	wire new_net_707;
	wire new_net_1000;
	wire new_net_1053;
	wire new_net_1074;
	wire new_net_1084;
	wire new_net_546;
	wire new_net_661;
	wire new_net_1743;
	wire new_net_2128;
	wire new_net_847;
	wire new_net_1182;
	wire new_net_2165;
	wire new_net_1626;
	wire new_net_1787;
	wire new_net_2469;
	wire new_net_1354;
	wire new_net_1619;
	wire new_net_1780;
	wire new_net_2211;
	wire new_net_1877;
	wire _0459_;
	wire new_net_39;
	wire new_net_504;
	wire new_net_453;
	wire _0039_;
	wire _0081_;
	wire _0123_;
	wire _0207_;
	wire _0249_;
	wire _0291_;
	wire new_net_169;
	wire new_net_2180;
	wire new_net_2368;
	wire new_net_2743;
	wire new_net_1270;
	wire new_net_878;
	wire new_net_1683;
	wire new_net_2009;
	wire new_net_1561;
	wire new_net_1227;
	wire new_net_597;
	wire new_net_1340;
	wire new_net_1868;
	wire new_net_2014;
	wire new_net_2191;
	wire new_net_2250;
	wire new_net_2756;
	wire new_net_1284;
	wire new_net_2270;
	wire new_net_2308;
	wire new_net_2385;
	wire new_net_1456;
	wire new_net_1735;
	wire new_net_1613;
	wire _0458_;
	wire new_net_909;
	wire new_net_1865;
	wire new_net_1738;
	wire new_net_2546;
	wire new_net_1493;
	wire new_net_263;
	wire new_net_470;
	wire new_net_542;
	wire _0460_;
	wire new_net_296;
	wire new_net_560;
	wire new_net_698;
	wire _0208_;
	wire _0250_;
	wire _0292_;
	wire _0475_;
	wire new_net_1389;
	wire new_net_1462;
	wire new_net_1670;
	wire new_net_2769;
	wire new_net_2663;
	wire new_net_2330;
	wire new_net_1835;
	wire new_net_940;
	wire new_net_1442;
	wire new_net_72;
	wire new_net_123;
	wire new_net_177;
	wire new_net_195;
	wire new_net_718;
	wire new_net_972;
	wire new_net_1165;
	wire new_net_1600;
	wire new_net_1766;
	wire new_net_1973;
	wire new_net_2079;
	wire new_net_810;
	wire new_net_1163;
	wire new_net_2521;
	wire new_net_1851;
	wire new_net_382;
	wire new_net_816;
	wire new_net_2603;
	wire new_net_2685;
	wire new_net_1898;
	wire new_net_389;
	wire new_net_2157;
	wire new_net_2417;
	wire new_net_40;
	wire new_net_247;
	wire new_net_505;
	wire new_net_454;
	wire _0461_;
	wire _0209_;
	wire _0251_;
	wire _0293_;
	wire _0041_;
	wire _0083_;
	wire new_net_1532;
	wire new_net_1701;
	wire new_net_1944;
	wire new_net_841;
	wire _0336_;
	wire new_net_1748;
	wire new_net_429;
	wire new_net_2176;
	wire new_net_1631;
	wire new_net_1792;
	wire new_net_2474;
	wire new_net_2777;
	wire new_net_8;
	wire new_net_347;
	wire _0353_;
	wire new_net_437;
	wire new_net_993;
	wire new_net_1476;
	wire new_net_1663;
	wire new_net_1686;
	wire new_net_1951;
	wire new_net_2007;
	wire new_net_2216;
	wire new_net_2251;
	wire _0377_;
	wire new_net_1882;
	wire new_net_1764;
	wire _0394_;
	wire new_net_872;
	wire new_net_2185;
	wire new_net_2748;
	wire _0418_;
	wire new_net_381;
	wire new_net_561;
	wire new_net_543;
	wire _0420_;
	wire new_net_18;
	wire new_net_471;
	wire _0462_;
	wire new_net_594;
	wire new_net_9;
	wire _0252_;
	wire new_net_1688;
	wire _0435_;
	wire new_net_2196;
	wire new_net_1566;
	wire new_net_1380;
	wire new_net_2489;
	wire new_net_1818;
	wire new_net_2796;
	wire new_net_2765;
	wire new_net_748;
	wire new_net_2279;
	wire new_net_2027;
	wire new_net_2134;
	wire new_net_743;
	wire new_net_73;
	wire new_net_124;
	wire new_net_178;
	wire new_net_196;
	wire new_net_1020;
	wire new_net_1428;
	wire new_net_1767;
	wire new_net_2244;
	wire new_net_2530;
	wire new_net_2551;
	wire new_net_1498;
	wire new_net_2400;
	wire new_net_1021;
	wire new_net_2075;
	wire new_net_1842;
	wire new_net_1552;
	wire new_net_1857;
	wire new_net_2517;
	wire _0043_;
	wire _0085_;
	wire _0127_;
	wire _0211_;
	wire _0253_;
	wire _0169_;
	wire _0295_;
	wire _0337_;
	wire _0379_;
	wire _0463_;
	wire new_net_1364;
	wire new_net_1759;
	wire new_net_2599;
	wire new_net_1447;
	wire new_net_2120;
	wire new_net_2413;
	wire new_net_2533;
	wire new_net_2088;
	wire new_net_2350;
	wire new_net_1251;
	wire new_net_843;
	wire new_net_264;
	wire new_net_438;
	wire new_net_703;
	wire new_net_1361;
	wire new_net_1727;
	wire new_net_2026;
	wire new_net_2038;
	wire new_net_2133;
	wire _0313_;
	wire new_net_2171;
	wire new_net_1539;
	wire new_net_2426;
	wire new_net_2773;
	wire new_net_2733;
	wire new_net_1054;
	wire new_net_692;
	wire _0212_;
	wire _0254_;
	wire _0296_;
	wire _0044_;
	wire _0086_;
	wire _0128_;
	wire _0170_;
	wire _0338_;
	wire _0380_;
	wire new_net_874;
	wire new_net_1959;
	wire new_net_2479;
	wire new_net_1962;
	wire new_net_2631;
	wire new_net_2048;
	wire new_net_2485;
	wire new_net_74;
	wire new_net_125;
	wire new_net_179;
	wire new_net_197;
	wire new_net_1151;
	wire new_net_1158;
	wire new_net_1188;
	wire new_net_1208;
	wire new_net_1432;
	wire new_net_1961;
	wire new_net_2445;
	wire new_net_2574;
	wire _0442_;
	wire new_net_905;
	wire new_net_1573;
	wire new_net_2693;
	wire new_net_775;
	wire new_net_2653;
	wire new_net_507;
	wire _0213_;
	wire _0255_;
	wire _0297_;
	wire _0045_;
	wire _0087_;
	wire _0129_;
	wire _0171_;
	wire _0339_;
	wire _0381_;
	wire new_net_2284;
	wire new_net_1153;
	wire new_net_2556;
	wire new_net_806;
	wire new_net_2598;
	wire new_net_265;
	wire new_net_298;
	wire new_net_439;
	wire new_net_472;
	wire new_net_544;
	wire new_net_812;
	wire new_net_1055;
	wire new_net_1064;
	wire new_net_1076;
	wire new_net_1086;
	wire new_net_2409;
	wire new_net_1847;
	wire new_net_2562;
	wire new_net_1557;
	wire new_net_1930;
	wire new_net_2787;
	wire new_net_663;
	wire new_net_2714;
	wire new_net_1731;
	wire _0214_;
	wire _0256_;
	wire _0298_;
	wire _0172_;
	wire _0046_;
	wire _0088_;
	wire _0130_;
	wire _0340_;
	wire _0382_;
	wire new_net_667;
	wire new_net_837;
	wire new_net_2422;
	wire new_net_2459;
	wire new_net_2497;
	wire new_net_1661;
	wire new_net_975;
	wire new_net_2246;
	wire new_net_2804;
	wire new_net_1544;
	wire _0361_;
	wire new_net_42;
	wire new_net_75;
	wire new_net_126;
	wire new_net_180;
	wire new_net_249;
	wire _0354_;
	wire new_net_1193;
	wire new_net_1229;
	wire new_net_1386;
	wire new_net_1870;
	wire new_net_2175;
	wire new_net_2435;
	wire new_net_2468;
	wire new_net_2627;
	wire new_net_2738;
	wire _0378_;
	wire new_net_868;
	wire new_net_1638;
	wire new_net_1798;
	wire new_net_447;
	wire new_net_2481;
	wire new_net_1990;
	wire new_net_2219;
	wire new_net_2441;
	wire _0395_;
	wire _0419_;
	wire new_net_1207;
	wire new_net_1889;
	wire new_net_2305;
	wire new_net_349;
	wire _0173_;
	wire _0047_;
	wire _0089_;
	wire _0131_;
	wire _0215_;
	wire _0257_;
	wire _0299_;
	wire _0341_;
	wire _0383_;
	wire new_net_2382;
	wire new_net_2722;
	wire new_net_2649;
	wire new_net_1146;
	wire new_net_1222;
	wire new_net_1986;
	wire new_net_1319;
	wire new_net_1577;
	wire new_net_1739;
	wire new_net_299;
	wire new_net_440;
	wire new_net_563;
	wire new_net_694;
	wire new_net_545;
	wire new_net_1434;
	wire new_net_1975;
	wire new_net_2163;
	wire new_net_2182;
	wire new_net_2604;
	wire new_net_1047;
	wire new_net_2700;
	wire new_net_1089;
	wire new_net_2034;
	wire new_net_2291;
	wire new_net_1512;
	wire new_net_2558;
	wire new_net_1135;
	wire _0468_;
	wire new_net_216;
	wire _0048_;
	wire _0090_;
	wire _0132_;
	wire _0174_;
	wire _0216_;
	wire _0258_;
	wire _0300_;
	wire _0342_;
	wire new_net_2710;
	wire _0273_;
	wire new_net_2567;
	wire new_net_1846;
	wire new_net_2493;
	wire new_net_3;
	wire new_net_43;
	wire new_net_76;
	wire new_net_181;
	wire new_net_250;
	wire new_net_658;
	wire new_net_974;
	wire new_net_1429;
	wire new_net_1478;
	wire new_net_1665;
	wire _0314_;
	wire new_net_831;
	wire new_net_2617;
	wire new_net_1122;
	wire new_net_2542;
	wire new_net_2464;
	wire new_net_2431;
	wire new_net_1666;
	wire _0427_;
	wire new_net_19;
	wire _0049_;
	wire _0091_;
	wire _0133_;
	wire _0175_;
	wire _0217_;
	wire _0259_;
	wire _0301_;
	wire _0343_;
	wire new_net_643;
	wire new_net_1438;
	wire new_net_1803;
	wire new_net_441;
	wire new_net_564;
	wire new_net_688;
	wire new_net_1022;
	wire new_net_1190;
	wire new_net_1460;
	wire new_net_1769;
	wire new_net_1953;
	wire new_net_2396;
	wire new_net_2532;
	wire new_net_771;
	wire new_net_1285;
	wire new_net_1894;
	wire _0443_;
	wire new_net_705;
	wire new_net_1657;
	wire new_net_2131;
	wire new_net_2274;
	wire new_net_2727;
	wire new_net_2239;
	wire _0428_;
	wire new_net_385;
	wire new_net_598;
	wire _0050_;
	wire _0092_;
	wire _0134_;
	wire _0176_;
	wire _0218_;
	wire _0260_;
	wire _0302_;
	wire _0484_;
	wire new_net_1584;
	wire new_net_1992;
	wire new_net_2102;
	wire new_net_1152;
	wire new_net_802;
	wire new_net_1914;
	wire new_net_1359;
	wire new_net_2039;
	wire new_net_2296;
	wire new_net_182;
	wire new_net_350;
	wire new_net_458;
	wire new_net_660;
	wire new_net_1363;
	wire new_net_1388;
	wire new_net_1475;
	wire new_net_2028;
	wire new_net_2040;
	wire new_net_2135;
	wire new_net_1760;
	wire new_net_1517;
	wire new_net_2640;
	wire new_net_383;
	wire new_net_1972;
	wire new_net_2267;
	wire new_net_833;
	wire new_net_1173;
	wire new_net_1934;
	wire new_net_2609;
	wire new_net_2454;
	wire new_net_1171;
	wire new_net_2607;
	wire new_net_300;
	wire _0051_;
	wire _0093_;
	wire _0135_;
	wire _0177_;
	wire _0219_;
	wire _0261_;
	wire _0303_;
	wire _0345_;
	wire _0387_;
	wire new_net_2578;
	wire new_net_2689;
	wire _0321_;
	wire new_net_2167;
	wire new_net_2098;
	wire new_net_2427;
	wire new_net_2622;
	wire new_net_1503;
	wire new_net_2587;
	wire new_net_864;
	wire new_net_1160;
	wire new_net_1461;
	wire new_net_2117;
	wire new_net_2255;
	wire new_net_2379;
	wire new_net_2634;
	wire new_net_1426;
	wire new_net_2707;
	wire _0355_;
	wire new_net_2145;
	wire _0403_;
	wire _0396_;
	wire new_net_77;
	wire _0472_;
	wire new_net_218;
	wire _0220_;
	wire _0262_;
	wire _0304_;
	wire _0052_;
	wire _0094_;
	wire _0136_;
	wire _0178_;
	wire new_net_2235;
	wire new_net_2354;
	wire new_net_27;
	wire new_net_351;
	wire new_net_459;
	wire new_net_1057;
	wire new_net_1066;
	wire new_net_1088;
	wire new_net_1180;
	wire new_net_1256;
	wire new_net_1271;
	wire new_net_1436;
	wire new_net_1824;
	wire new_net_2506;
	wire new_net_1589;
	wire new_net_796;
	wire new_net_2595;
	wire new_net_2705;
	wire new_net_6;
	wire new_net_511;
	wire new_net_475;
	wire new_net_547;
	wire _0221_;
	wire _0263_;
	wire _0305_;
	wire _0053_;
	wire _0095_;
	wire _0137_;
	wire _0179_;
	wire new_net_2404;
	wire new_net_2784;
	wire new_net_2263;
	wire new_net_2753;
	wire new_net_1523;
	wire new_net_1692;
	wire new_net_1280;
	wire new_net_1521;
	wire new_net_2645;
	wire new_net_2419;
	wire new_net_827;
	wire new_net_4;
	wire new_net_200;
	wire new_net_1485;
	wire new_net_1728;
	wire new_net_1872;
	wire new_net_2018;
	wire new_net_2094;
	wire new_net_2195;
	wire new_net_2201;
	wire new_net_1178;
	wire new_net_2614;
	wire _0315_;
	wire new_net_1776;
	wire new_net_2801;
	wire new_net_852;
	wire new_net_2364;
	wire new_net_45;
	wire new_net_252;
	wire _0432_;
	wire new_net_129;
	wire new_net_78;
	wire _0180_;
	wire _0054_;
	wire _0096_;
	wire _0138_;
	wire _0222_;
	wire new_net_1266;
	wire new_net_1508;
	wire new_net_1715;
	wire new_net_2005;
	wire new_net_2187;
	wire new_net_1718;
	wire new_net_188;
	wire new_net_28;
	wire new_net_1126;
	wire new_net_1288;
	wire new_net_1904;
	wire new_net_1977;
	wire new_net_883;
	wire new_net_2184;
	wire new_net_2575;
	wire new_net_2668;
	wire new_net_2680;
	wire new_net_1452;
	wire new_net_1075;
	wire new_net_1609;
	wire new_net_1037;
	wire _0444_;
	wire new_net_2017;
	wire new_net_2390;
	wire new_net_302;
	wire new_net_443;
	wire new_net_512;
	wire _0433_;
	wire _0181_;
	wire _0055_;
	wire _0097_;
	wire _0139_;
	wire _0223_;
	wire _0265_;
	wire _0485_;
	wire new_net_1312;
	wire new_net_2659;
	wire new_net_2326;
	wire new_net_2697;
	wire new_net_914;
	wire new_net_2591;
	wire new_net_1829;
	wire new_net_2511;
	wire new_net_2071;
	wire new_net_2105;
	wire new_net_1596;
	wire new_net_2259;
	wire new_net_201;
	wire new_net_219;
	wire new_net_387;
	wire new_net_600;
	wire new_net_1159;
	wire new_net_1667;
	wire new_net_1750;
	wire new_net_2228;
	wire new_net_2247;
	wire new_net_2397;
	wire new_net_945;
	wire new_net_2341;
	wire new_net_2153;
	wire new_net_2758;
	wire new_net_1528;
	wire _0476_;
	wire new_net_352;
	wire _0224_;
	wire _0266_;
	wire _0056_;
	wire _0098_;
	wire _0140_;
	wire _0182_;
	wire _0308_;
	wire _0350_;
	wire new_net_269;
	wire new_net_1486;
	wire new_net_2129;
	wire new_net_1185;
	wire new_net_1744;
	wire new_net_2206;
	wire new_net_1183;
	wire new_net_2166;
	wire new_net_1627;
	wire new_net_1788;
	wire new_net_2470;
	wire new_net_1781;
	wire new_net_1398;
	wire new_net_2212;
	wire new_net_720;
	wire new_net_653;
	wire _0363_;
	wire new_net_1024;
	wire new_net_1192;
	wire new_net_1407;
	wire new_net_1771;
	wire new_net_1955;
	wire new_net_2467;
	wire new_net_1878;
	wire _0356_;
	wire new_net_301;
	wire new_net_2181;
	wire new_net_2744;
	wire new_net_37;
	wire new_net_2113;
	wire _0404_;
	wire _0397_;
	wire new_net_1684;
	wire new_net_44;
	wire new_net_270;
	wire new_net_686;
	wire new_net_477;
	wire new_net_549;
	wire new_net_455;
	wire _0477_;
	wire new_net_303;
	wire _0225_;
	wire _0267_;
	wire _0057_;
	wire _0421_;
	wire _0431_;
	wire new_net_649;
	wire new_net_1562;
	wire new_net_1210;
	wire new_net_1772;
	wire new_net_1457;
	wire new_net_1736;
	wire new_net_1078;
	wire new_net_1614;
	wire new_net_601;
	wire new_net_46;
	wire new_net_202;
	wire new_net_220;
	wire new_net_253;
	wire new_net_388;
	wire new_net_1365;
	wire new_net_1866;
	wire new_net_2030;
	wire new_net_1494;
	wire new_net_2547;
	wire new_net_792;
	wire new_net_1017;
	wire new_net_2770;
	wire new_net_2664;
	wire new_net_2331;
	wire new_net_2513;
	wire new_net_1836;
	wire new_net_1360;
	wire _0436_;
	wire new_net_461;
	wire new_net_719;
	wire new_net_29;
	wire new_net_80;
	wire _0478_;
	wire new_net_353;
	wire _0226_;
	wire _0268_;
	wire _0142_;
	wire new_net_1443;
	wire new_net_2337;
	wire new_net_2372;
	wire new_net_1601;
	wire new_net_2080;
	wire new_net_2529;
	wire new_net_2346;
	wire new_net_2522;
	wire _0282_;
	wire new_net_823;
	wire new_net_1852;
	wire new_net_2686;
	wire new_net_1402;
	wire new_net_1850;
	wire new_net_567;
	wire new_net_669;
	wire new_net_444;
	wire new_net_1162;
	wire new_net_1463;
	wire new_net_1487;
	wire new_net_1730;
	wire new_net_2418;
	wire new_net_2457;
	wire new_net_2636;
	wire new_net_1535;
	wire new_net_1533;
	wire new_net_1702;
	wire new_net_548;
	wire new_net_1945;
	wire new_net_848;
	wire new_net_1050;
	wire new_net_1749;
	wire new_net_304;
	wire new_net_747;
	wire new_net_550;
	wire new_net_514;
	wire _0437_;
	wire _0059_;
	wire _0101_;
	wire _0227_;
	wire _0269_;
	wire _0143_;
	wire new_net_1465;
	wire new_net_1632;
	wire new_net_1793;
	wire new_net_2475;
	wire new_net_2778;
	wire new_net_171;
	wire new_net_1097;
	wire new_net_2217;
	wire new_net_1883;
	wire new_net_879;
	wire new_net_2749;
	wire new_net_602;
	wire new_net_47;
	wire new_net_131;
	wire new_net_185;
	wire new_net_203;
	wire new_net_221;
	wire new_net_254;
	wire new_net_740;
	wire new_net_1059;
	wire new_net_1068;
	wire new_net_2053;
	wire new_net_2232;
	wire new_net_599;
	wire new_net_1567;
	wire _0445_;
	wire new_net_2797;
	wire new_net_910;
	wire _0480_;
	wire new_net_354;
	wire _0438_;
	wire _0228_;
	wire _0270_;
	wire _0060_;
	wire _0102_;
	wire _0144_;
	wire _0186_;
	wire _0312_;
	wire _0486_;
	wire new_net_2280;
	wire _0479_;
	wire new_net_2658;
	wire new_net_2702;
	wire new_net_1871;
	wire new_net_1262;
	wire new_net_2552;
	wire new_net_1499;
	wire new_net_2401;
	wire new_net_2671;
	wire new_net_2076;
	wire new_net_2669;
	wire new_net_271;
	wire new_net_478;
	wire new_net_568;
	wire new_net_1752;
	wire new_net_1553;
	wire new_net_1874;
	wire new_net_2020;
	wire new_net_2197;
	wire new_net_2762;
	wire new_net_941;
	wire new_net_2518;
	wire new_net_1841;
	wire new_net_377;
	wire new_net_2600;
	wire new_net_513;
	wire new_net_1448;
	wire new_net_2121;
	wire new_net_384;
	wire new_net_817;
	wire new_net_2534;
	wire new_net_2089;
	wire new_net_676;
	wire new_net_704;
	wire new_net_551;
	wire _0481_;
	wire new_net_515;
	wire _0229_;
	wire _0271_;
	wire _0061_;
	wire _0103_;
	wire _0145_;
	wire new_net_20;
	wire new_net_1252;
	wire new_net_1415;
	wire new_net_1704;
	wire new_net_1540;
	wire new_net_2138;
	wire new_net_1189;
	wire new_net_2734;
	wire new_net_132;
	wire new_net_186;
	wire new_net_204;
	wire new_net_1143;
	wire new_net_1170;
	wire new_net_1290;
	wire new_net_1343;
	wire new_net_1906;
	wire new_net_1979;
	wire new_net_2229;
	wire _0357_;
	wire new_net_2626;
	wire new_net_1960;
	wire new_net_2480;
	wire _0405_;
	wire new_net_2301;
	wire new_net_2632;
	wire new_net_2049;
	wire _0398_;
	wire new_net_873;
	wire new_net_1719;
	wire new_net_671;
	wire _0440_;
	wire new_net_642;
	wire new_net_82;
	wire _0482_;
	wire new_net_355;
	wire _0230_;
	wire _0272_;
	wire _0146_;
	wire _0188_;
	wire _0422_;
	wire new_net_1063;
	wire new_net_2446;
	wire _0439_;
	wire new_net_1982;
	wire new_net_1574;
	wire new_net_672;
	wire new_net_724;
	wire new_net_272;
	wire new_net_305;
	wire new_net_479;
	wire new_net_977;
	wire new_net_1235;
	wire new_net_1669;
	wire new_net_2137;
	wire new_net_2399;
	wire new_net_1085;
	wire new_net_2358;
	wire new_net_2068;
	wire new_net_2285;
	wire new_net_2557;
	wire new_net_48;
	wire new_net_255;
	wire _0441_;
	wire new_net_390;
	wire new_net_21;
	wire new_net_552;
	wire new_net_735;
	wire _0483_;
	wire new_net_222;
	wire _0231_;
	wire new_net_2676;
	wire new_net_2709;
	wire new_net_2410;
	wire new_net_2563;
	wire new_net_1931;
	wire new_net_2085;
	wire new_net_2408;
	wire new_net_2788;
	wire new_net_2715;
	wire new_net_31;
	wire new_net_133;
	wire new_net_205;
	wire new_net_662;
	wire new_net_741;
	wire new_net_1026;
	wire new_net_1194;
	wire new_net_1409;
	wire new_net_1433;
	wire new_net_1773;
	wire new_net_844;
	wire new_net_2423;
	wire new_net_2538;
	wire new_net_1862;
	wire new_net_1257;
	wire new_net_2460;
	wire new_net_2498;
	wire new_net_1662;
	wire new_net_2805;
	wire new_net_1293;
	input G1;
	input G10;
	input G100;
	input G101;
	input G102;
	input G103;
	input G104;
	input G105;
	input G106;
	input G107;
	input G108;
	input G109;
	input G11;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G12;
	input G120;
	input G121;
	input G122;
	input G123;
	input G124;
	input G125;
	input G126;
	input G127;
	input G128;
	input G129;
	input G13;
	input G130;
	input G131;
	input G132;
	input G133;
	input G134;
	input G135;
	input G136;
	input G137;
	input G138;
	input G139;
	input G14;
	input G140;
	input G141;
	input G142;
	input G143;
	input G144;
	input G145;
	input G146;
	input G147;
	input G148;
	input G149;
	input G15;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G16;
	input G17;
	input G18;
	input G19;
	input G2;
	input G20;
	input G21;
	input G22;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G28;
	input G29;
	input G3;
	input G30;
	input G31;
	input G32;
	input G33;
	input G34;
	input G35;
	input G36;
	input G37;
	input G38;
	input G39;
	input G4;
	input G40;
	input G41;
	input G42;
	input G43;
	input G44;
	input G45;
	input G46;
	input G47;
	input G48;
	input G49;
	input G5;
	input G50;
	input G51;
	input G52;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G6;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G67;
	input G68;
	input G69;
	input G7;
	input G70;
	input G71;
	input G72;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G8;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G9;
	input G90;
	input G91;
	input G92;
	input G93;
	input G94;
	input G95;
	input G96;
	input G97;
	input G98;
	input G99;
	output G2531;
	output G2532;
	output G2533;
	output G2534;
	output G2535;
	output G2536;
	output G2537;
	output G2538;
	output G2539;
	output G2540;
	output G2541;
	output G2542;
	output G2543;
	output G2544;
	output G2545;
	output G2546;
	output G2547;
	output G2548;
	output G2549;
	output G2550;
	output G2551;
	output G2552;
	output G2553;
	output G2554;
	output G2555;
	output G2556;
	output G2557;
	output G2558;
	output G2559;
	output G2560;
	output G2561;
	output G2562;
	output G2563;
	output G2564;
	output G2565;
	output G2566;
	output G2567;
	output G2568;
	output G2569;
	output G2570;
	output G2571;
	output G2572;
	output G2573;
	output G2574;
	output G2575;
	output G2576;
	output G2577;
	output G2578;
	output G2579;
	output G2580;
	output G2581;
	output G2582;
	output G2583;
	output G2584;
	output G2585;
	output G2586;
	output G2587;
	output G2588;
	output G2589;
	output G2590;
	output G2591;
	output G2592;
	output G2593;
	output G2594;

	or_bb _0499_ (
		.a(new_net_114),
		.b(new_net_157),
		.c(_0000_)
	);

	or_bb _0500_ (
		.a(new_net_632),
		.b(new_net_750),
		.c(_0001_)
	);

	or_bb _0501_ (
		.a(new_net_115),
		.b(new_net_159),
		.c(_0002_)
	);

	and_bi _0502_ (
		.a(new_net_751),
		.b(new_net_538),
		.c(_0003_)
	);

	and_bi _0503_ (
		.a(_0001_),
		.b(_0003_),
		.c(_0004_)
	);

	or_bb _0504_ (
		.a(new_net_116),
		.b(new_net_160),
		.c(_0005_)
	);

	and_bi _0505_ (
		.a(new_net_752),
		.b(new_net_118),
		.c(_0006_)
	);

	or_bb _0506_ (
		.a(new_net_117),
		.b(new_net_158),
		.c(_0007_)
	);

	and_bi _0507_ (
		.a(new_net_753),
		.b(new_net_174),
		.c(_0008_)
	);

	or_bb _0508_ (
		.a(_0008_),
		.b(_0006_),
		.c(_0009_)
	);

	and_bi _0509_ (
		.a(_0004_),
		.b(_0009_),
		.c(new_net_2)
	);

	or_bb _0510_ (
		.a(new_net_180),
		.b(new_net_754),
		.c(_0010_)
	);

	and_bi _0511_ (
		.a(new_net_755),
		.b(new_net_121),
		.c(_0011_)
	);

	and_bi _0512_ (
		.a(_0010_),
		.b(_0011_),
		.c(_0012_)
	);

	and_bi _0513_ (
		.a(new_net_756),
		.b(new_net_536),
		.c(_0013_)
	);

	and_bi _0514_ (
		.a(new_net_757),
		.b(new_net_635),
		.c(_0014_)
	);

	or_bb _0515_ (
		.a(_0014_),
		.b(_0013_),
		.c(_0015_)
	);

	and_bi _0516_ (
		.a(_0012_),
		.b(_0015_),
		.c(new_net_0)
	);

	and_bi _0517_ (
		.a(new_net_758),
		.b(new_net_175),
		.c(_0016_)
	);

	and_bi _0518_ (
		.a(new_net_759),
		.b(new_net_634),
		.c(_0017_)
	);

	or_bb _0519_ (
		.a(_0017_),
		.b(_0016_),
		.c(_0018_)
	);

	and_bi _0520_ (
		.a(new_net_760),
		.b(new_net_540),
		.c(_0019_)
	);

	and_bi _0521_ (
		.a(new_net_761),
		.b(new_net_119),
		.c(_0020_)
	);

	or_bb _0522_ (
		.a(_0020_),
		.b(_0019_),
		.c(_0021_)
	);

	or_bb _0523_ (
		.a(_0021_),
		.b(_0018_),
		.c(new_net_1)
	);

	and_bi _0524_ (
		.a(new_net_404),
		.b(new_net_762),
		.c(_0022_)
	);

	and_bi _0525_ (
		.a(new_net_391),
		.b(new_net_763),
		.c(_0023_)
	);

	or_bb _0526_ (
		.a(_0023_),
		.b(new_net_550),
		.c(_0024_)
	);

	and_bi _0527_ (
		.a(new_net_764),
		.b(_0024_),
		.c(_0025_)
	);

	or_bb _0528_ (
		.a(new_net_552),
		.b(new_net_399),
		.c(_0026_)
	);

	and_bi _0529_ (
		.a(new_net_765),
		.b(new_net_33),
		.c(_0027_)
	);

	or_bb _0530_ (
		.a(new_net_553),
		.b(new_net_405),
		.c(_0028_)
	);

	and_bi _0531_ (
		.a(new_net_766),
		.b(new_net_200),
		.c(_0029_)
	);

	or_bb _0532_ (
		.a(_0029_),
		.b(_0027_),
		.c(_0030_)
	);

	and_bi _0533_ (
		.a(new_net_767),
		.b(_0030_),
		.c(new_net_8)
	);

	and_bi _0534_ (
		.a(new_net_768),
		.b(new_net_206),
		.c(_0031_)
	);

	or_bb _0535_ (
		.a(new_net_769),
		.b(new_net_396),
		.c(_0032_)
	);

	and_bi _0536_ (
		.a(new_net_406),
		.b(new_net_770),
		.c(_0033_)
	);

	or_bb _0537_ (
		.a(_0033_),
		.b(new_net_546),
		.c(_0034_)
	);

	and_bi _0538_ (
		.a(new_net_771),
		.b(_0034_),
		.c(_0035_)
	);

	and_bi _0539_ (
		.a(_0031_),
		.b(new_net_772),
		.c(new_net_6)
	);

	and_bi _0540_ (
		.a(new_net_407),
		.b(new_net_773),
		.c(_0036_)
	);

	and_bi _0541_ (
		.a(new_net_392),
		.b(new_net_774),
		.c(_0037_)
	);

	or_bb _0542_ (
		.a(_0037_),
		.b(new_net_551),
		.c(_0038_)
	);

	and_bi _0543_ (
		.a(new_net_775),
		.b(_0038_),
		.c(_0039_)
	);

	and_bi _0544_ (
		.a(new_net_776),
		.b(new_net_40),
		.c(_0040_)
	);

	and_bi _0545_ (
		.a(new_net_777),
		.b(new_net_201),
		.c(_0041_)
	);

	or_bb _0546_ (
		.a(_0041_),
		.b(_0040_),
		.c(_0042_)
	);

	and_bi _0547_ (
		.a(new_net_778),
		.b(_0042_),
		.c(new_net_5)
	);

	and_bi _0548_ (
		.a(new_net_408),
		.b(new_net_779),
		.c(_0043_)
	);

	and_bi _0549_ (
		.a(new_net_393),
		.b(new_net_780),
		.c(_0044_)
	);

	or_bb _0550_ (
		.a(_0044_),
		.b(new_net_554),
		.c(_0045_)
	);

	and_bi _0551_ (
		.a(new_net_781),
		.b(_0045_),
		.c(_0046_)
	);

	and_bi _0552_ (
		.a(new_net_782),
		.b(new_net_39),
		.c(_0047_)
	);

	and_bi _0553_ (
		.a(new_net_783),
		.b(new_net_202),
		.c(_0048_)
	);

	or_bb _0554_ (
		.a(_0048_),
		.b(_0047_),
		.c(_0049_)
	);

	and_bi _0555_ (
		.a(new_net_784),
		.b(_0049_),
		.c(new_net_3)
	);

	and_bi _0556_ (
		.a(new_net_411),
		.b(new_net_785),
		.c(_0050_)
	);

	and_bi _0557_ (
		.a(new_net_397),
		.b(new_net_786),
		.c(_0051_)
	);

	or_bb _0558_ (
		.a(_0051_),
		.b(new_net_555),
		.c(_0052_)
	);

	and_bi _0559_ (
		.a(new_net_787),
		.b(_0052_),
		.c(_0053_)
	);

	and_bi _0560_ (
		.a(new_net_788),
		.b(new_net_37),
		.c(_0054_)
	);

	and_bi _0561_ (
		.a(new_net_789),
		.b(new_net_203),
		.c(_0055_)
	);

	or_bb _0562_ (
		.a(_0055_),
		.b(_0054_),
		.c(_0056_)
	);

	and_bi _0563_ (
		.a(new_net_790),
		.b(_0056_),
		.c(new_net_4)
	);

	or_bb _0564_ (
		.a(new_net_791),
		.b(new_net_400),
		.c(_0057_)
	);

	and_bi _0565_ (
		.a(new_net_394),
		.b(new_net_792),
		.c(_0058_)
	);

	or_bb _0566_ (
		.a(_0058_),
		.b(new_net_556),
		.c(_0059_)
	);

	and_bi _0567_ (
		.a(new_net_793),
		.b(_0059_),
		.c(_0060_)
	);

	and_bi _0568_ (
		.a(new_net_794),
		.b(new_net_38),
		.c(_0061_)
	);

	and_bi _0569_ (
		.a(new_net_795),
		.b(new_net_204),
		.c(_0062_)
	);

	or_bb _0570_ (
		.a(_0062_),
		.b(_0061_),
		.c(_0063_)
	);

	or_bb _0571_ (
		.a(_0063_),
		.b(new_net_796),
		.c(new_net_9)
	);

	and_bi _0572_ (
		.a(new_net_409),
		.b(new_net_797),
		.c(_0064_)
	);

	and_bi _0573_ (
		.a(new_net_395),
		.b(new_net_798),
		.c(_0065_)
	);

	or_bb _0574_ (
		.a(_0065_),
		.b(new_net_557),
		.c(_0066_)
	);

	and_bi _0575_ (
		.a(new_net_799),
		.b(_0066_),
		.c(_0067_)
	);

	and_bi _0576_ (
		.a(new_net_800),
		.b(new_net_41),
		.c(_0068_)
	);

	and_bi _0577_ (
		.a(new_net_801),
		.b(new_net_205),
		.c(_0069_)
	);

	or_bb _0578_ (
		.a(_0069_),
		.b(_0068_),
		.c(_0070_)
	);

	and_bi _0579_ (
		.a(new_net_802),
		.b(_0070_),
		.c(new_net_7)
	);

	and_bi _0580_ (
		.a(new_net_439),
		.b(new_net_302),
		.c(_0071_)
	);

	and_bi _0581_ (
		.a(new_net_438),
		.b(new_net_300),
		.c(_0072_)
	);

	and_bi _0582_ (
		.a(_0071_),
		.b(_0072_),
		.c(_0073_)
	);

	and_bi _0583_ (
		.a(new_net_442),
		.b(new_net_163),
		.c(_0074_)
	);

	and_bi _0584_ (
		.a(new_net_443),
		.b(new_net_165),
		.c(_0075_)
	);

	and_bi _0585_ (
		.a(_0074_),
		.b(_0075_),
		.c(_0076_)
	);

	and_bi _0586_ (
		.a(new_net_273),
		.b(new_net_350),
		.c(_0077_)
	);

	and_bi _0587_ (
		.a(new_net_274),
		.b(new_net_351),
		.c(_0078_)
	);

	and_bi _0588_ (
		.a(_0077_),
		.b(_0078_),
		.c(_0079_)
	);

	and_bi _0589_ (
		.a(new_net_381),
		.b(new_net_417),
		.c(_0080_)
	);

	and_bi _0590_ (
		.a(new_net_386),
		.b(new_net_419),
		.c(_0081_)
	);

	and_bi _0591_ (
		.a(_0080_),
		.b(_0081_),
		.c(_0082_)
	);

	and_bi _0592_ (
		.a(new_net_458),
		.b(new_net_567),
		.c(_0083_)
	);

	and_bi _0593_ (
		.a(new_net_459),
		.b(new_net_568),
		.c(_0084_)
	);

	and_bi _0594_ (
		.a(_0083_),
		.b(_0084_),
		.c(_0085_)
	);

	and_bi _0595_ (
		.a(new_net_214),
		.b(new_net_279),
		.c(_0086_)
	);

	and_bi _0596_ (
		.a(new_net_218),
		.b(new_net_281),
		.c(_0087_)
	);

	and_bi _0597_ (
		.a(_0086_),
		.b(_0087_),
		.c(_0088_)
	);

	and_bi _0598_ (
		.a(new_net_332),
		.b(new_net_355),
		.c(_0089_)
	);

	and_bi _0599_ (
		.a(new_net_331),
		.b(new_net_352),
		.c(_0090_)
	);

	and_bi _0600_ (
		.a(_0089_),
		.b(_0090_),
		.c(_0091_)
	);

	and_bi _0601_ (
		.a(new_net_102),
		.b(new_net_185),
		.c(_0092_)
	);

	and_bi _0602_ (
		.a(new_net_103),
		.b(new_net_186),
		.c(_0093_)
	);

	and_bi _0603_ (
		.a(_0092_),
		.b(_0093_),
		.c(_0094_)
	);

	and_bi _0604_ (
		.a(new_net_260),
		.b(new_net_328),
		.c(_0095_)
	);

	and_bi _0605_ (
		.a(new_net_261),
		.b(new_net_329),
		.c(_0096_)
	);

	or_bb _0606_ (
		.a(_0096_),
		.b(_0095_),
		.c(new_net_13)
	);

	or_bb _0607_ (
		.a(new_net_24),
		.b(new_net_623),
		.c(_0097_)
	);

	and_bi _0608_ (
		.a(new_net_627),
		.b(new_net_28),
		.c(_0098_)
	);

	and_bi _0609_ (
		.a(new_net_348),
		.b(new_net_803),
		.c(_0099_)
	);

	or_bb _0610_ (
		.a(new_net_580),
		.b(new_net_520),
		.c(_0100_)
	);

	and_bi _0611_ (
		.a(new_net_519),
		.b(new_net_579),
		.c(_0101_)
	);

	and_bi _0612_ (
		.a(new_net_619),
		.b(new_net_804),
		.c(_0102_)
	);

	and_bi _0613_ (
		.a(new_net_446),
		.b(new_net_262),
		.c(_0103_)
	);

	and_bi _0614_ (
		.a(new_net_447),
		.b(new_net_263),
		.c(_0104_)
	);

	and_bi _0615_ (
		.a(_0103_),
		.b(_0104_),
		.c(_0105_)
	);

	and_bi _0616_ (
		.a(new_net_48),
		.b(new_net_485),
		.c(_0106_)
	);

	and_bi _0617_ (
		.a(new_net_51),
		.b(new_net_483),
		.c(_0107_)
	);

	and_bi _0618_ (
		.a(_0106_),
		.b(_0107_),
		.c(_0108_)
	);

	and_bi _0619_ (
		.a(new_net_470),
		.b(new_net_65),
		.c(_0109_)
	);

	and_bi _0620_ (
		.a(new_net_471),
		.b(new_net_66),
		.c(_0110_)
	);

	and_bi _0621_ (
		.a(_0109_),
		.b(_0110_),
		.c(_0111_)
	);

	and_bi _0622_ (
		.a(new_net_108),
		.b(new_net_161),
		.c(_0112_)
	);

	and_bi _0623_ (
		.a(new_net_109),
		.b(new_net_162),
		.c(_0113_)
	);

	and_bi _0624_ (
		.a(_0112_),
		.b(_0113_),
		.c(_0114_)
	);

	and_bi _0625_ (
		.a(new_net_96),
		.b(new_net_371),
		.c(_0115_)
	);

	and_bi _0626_ (
		.a(new_net_97),
		.b(new_net_372),
		.c(_0116_)
	);

	or_bb _0627_ (
		.a(_0116_),
		.b(_0115_),
		.c(new_net_12)
	);

	and_bi _0628_ (
		.a(new_net_98),
		.b(new_net_341),
		.c(_0117_)
	);

	and_bi _0629_ (
		.a(new_net_99),
		.b(new_net_342),
		.c(_0118_)
	);

	and_bi _0630_ (
		.a(_0117_),
		.b(_0118_),
		.c(_0119_)
	);

	and_bi _0631_ (
		.a(new_net_621),
		.b(new_net_232),
		.c(_0120_)
	);

	and_bi _0632_ (
		.a(new_net_622),
		.b(new_net_233),
		.c(_0121_)
	);

	and_bi _0633_ (
		.a(_0120_),
		.b(_0121_),
		.c(_0122_)
	);

	and_bi _0634_ (
		.a(new_net_495),
		.b(new_net_489),
		.c(_0123_)
	);

	and_bi _0635_ (
		.a(new_net_496),
		.b(new_net_490),
		.c(_0124_)
	);

	and_bi _0636_ (
		.a(_0123_),
		.b(_0124_),
		.c(_0125_)
	);

	and_bi _0637_ (
		.a(new_net_264),
		.b(new_net_291),
		.c(_0126_)
	);

	and_bi _0638_ (
		.a(new_net_265),
		.b(new_net_292),
		.c(_0127_)
	);

	and_bi _0639_ (
		.a(_0126_),
		.b(_0127_),
		.c(_0128_)
	);

	and_bi _0640_ (
		.a(new_net_110),
		.b(new_net_52),
		.c(_0129_)
	);

	and_bi _0641_ (
		.a(new_net_111),
		.b(new_net_53),
		.c(_0130_)
	);

	or_bb _0642_ (
		.a(_0130_),
		.b(_0129_),
		.c(_0131_)
	);

	or_bb _0643_ (
		.a(new_net_193),
		.b(new_net_72),
		.c(_0132_)
	);

	and_bi _0644_ (
		.a(new_net_75),
		.b(new_net_195),
		.c(_0133_)
	);

	and_bi _0645_ (
		.a(_0132_),
		.b(_0133_),
		.c(_0134_)
	);

	and_bi _0646_ (
		.a(new_net_377),
		.b(new_net_413),
		.c(_0135_)
	);

	and_bi _0647_ (
		.a(new_net_378),
		.b(new_net_414),
		.c(_0136_)
	);

	and_bi _0648_ (
		.a(_0135_),
		.b(_0136_),
		.c(_0137_)
	);

	or_bb _0649_ (
		.a(new_net_289),
		.b(new_net_222),
		.c(_0138_)
	);

	and_bi _0650_ (
		.a(new_net_223),
		.b(new_net_290),
		.c(_0139_)
	);

	and_bi _0651_ (
		.a(_0138_),
		.b(_0139_),
		.c(_0140_)
	);

	and_ii _0652_ (
		.a(new_net_379),
		.b(new_net_373),
		.c(_0141_)
	);

	and_bb _0653_ (
		.a(new_net_380),
		.b(new_net_374),
		.c(_0142_)
	);

	or_bb _0654_ (
		.a(_0142_),
		.b(new_net_805),
		.c(_0143_)
	);

	and_bi _0655_ (
		.a(new_net_806),
		.b(_0143_),
		.c(new_net_14)
	);

	and_bi _0656_ (
		.a(new_net_807),
		.b(new_net_628),
		.c(_0144_)
	);

	and_bi _0657_ (
		.a(new_net_808),
		.b(new_net_123),
		.c(_0145_)
	);

	and_bi _0658_ (
		.a(_0144_),
		.b(_0145_),
		.c(_0146_)
	);

	and_bi _0659_ (
		.a(new_net_809),
		.b(new_net_181),
		.c(_0147_)
	);

	and_bi _0660_ (
		.a(new_net_810),
		.b(new_net_535),
		.c(_0148_)
	);

	or_bb _0661_ (
		.a(_0148_),
		.b(_0147_),
		.c(_0149_)
	);

	and_bi _0662_ (
		.a(_0146_),
		.b(_0149_),
		.c(_0150_)
	);

	or_bb _0663_ (
		.a(new_net_85),
		.b(new_net_467),
		.c(_0151_)
	);

	and_bi _0664_ (
		.a(new_net_465),
		.b(new_net_84),
		.c(_0152_)
	);

	and_bi _0665_ (
		.a(_0151_),
		.b(_0152_),
		.c(_0153_)
	);

	or_bb _0666_ (
		.a(new_net_100),
		.b(new_net_267),
		.c(_0154_)
	);

	and_bi _0667_ (
		.a(new_net_101),
		.b(new_net_270),
		.c(_0155_)
	);

	and_bi _0668_ (
		.a(_0154_),
		.b(_0155_),
		.c(_0156_)
	);

	and_bi _0669_ (
		.a(new_net_811),
		.b(new_net_539),
		.c(_0157_)
	);

	and_bi _0670_ (
		.a(new_net_812),
		.b(new_net_120),
		.c(_0158_)
	);

	and_bi _0671_ (
		.a(_0157_),
		.b(_0158_),
		.c(_0159_)
	);

	and_bi _0672_ (
		.a(new_net_813),
		.b(new_net_176),
		.c(_0160_)
	);

	and_bi _0673_ (
		.a(new_net_814),
		.b(new_net_633),
		.c(_0161_)
	);

	or_bb _0674_ (
		.a(_0161_),
		.b(_0160_),
		.c(_0162_)
	);

	and_bi _0675_ (
		.a(_0159_),
		.b(_0162_),
		.c(_0163_)
	);

	and_bi _0676_ (
		.a(new_net_815),
		.b(new_net_629),
		.c(_0164_)
	);

	and_bi _0677_ (
		.a(new_net_816),
		.b(new_net_124),
		.c(_0165_)
	);

	and_bi _0678_ (
		.a(_0164_),
		.b(_0165_),
		.c(_0166_)
	);

	and_bi _0679_ (
		.a(new_net_817),
		.b(new_net_182),
		.c(_0167_)
	);

	and_bi _0680_ (
		.a(new_net_818),
		.b(new_net_537),
		.c(_0168_)
	);

	or_bb _0681_ (
		.a(_0168_),
		.b(_0167_),
		.c(_0169_)
	);

	and_bi _0682_ (
		.a(_0166_),
		.b(_0169_),
		.c(_0170_)
	);

	and_bi _0683_ (
		.a(new_net_449),
		.b(new_net_56),
		.c(_0171_)
	);

	and_bi _0684_ (
		.a(new_net_448),
		.b(new_net_55),
		.c(_0172_)
	);

	and_bi _0685_ (
		.a(_0171_),
		.b(_0172_),
		.c(_0173_)
	);

	and_bi _0686_ (
		.a(new_net_819),
		.b(new_net_630),
		.c(_0174_)
	);

	and_bi _0687_ (
		.a(new_net_820),
		.b(new_net_541),
		.c(_0175_)
	);

	and_bi _0688_ (
		.a(_0174_),
		.b(_0175_),
		.c(_0176_)
	);

	and_bi _0689_ (
		.a(new_net_821),
		.b(new_net_125),
		.c(_0177_)
	);

	and_bi _0690_ (
		.a(new_net_822),
		.b(new_net_177),
		.c(_0178_)
	);

	or_bb _0691_ (
		.a(_0178_),
		.b(_0177_),
		.c(_0179_)
	);

	and_bi _0692_ (
		.a(_0176_),
		.b(_0179_),
		.c(_0180_)
	);

	and_bi _0693_ (
		.a(new_net_823),
		.b(new_net_636),
		.c(_0181_)
	);

	and_bi _0694_ (
		.a(new_net_824),
		.b(new_net_122),
		.c(_0182_)
	);

	and_bi _0695_ (
		.a(_0181_),
		.b(_0182_),
		.c(_0183_)
	);

	and_bi _0696_ (
		.a(new_net_825),
		.b(new_net_178),
		.c(_0184_)
	);

	and_bi _0697_ (
		.a(new_net_826),
		.b(new_net_542),
		.c(_0185_)
	);

	or_bb _0698_ (
		.a(_0185_),
		.b(_0184_),
		.c(_0186_)
	);

	and_bi _0699_ (
		.a(_0183_),
		.b(_0186_),
		.c(_0187_)
	);

	and_bi _0700_ (
		.a(new_net_312),
		.b(new_net_560),
		.c(_0188_)
	);

	and_bi _0701_ (
		.a(new_net_313),
		.b(new_net_562),
		.c(_0189_)
	);

	and_bi _0702_ (
		.a(_0188_),
		.b(_0189_),
		.c(_0190_)
	);

	and_bi _0703_ (
		.a(new_net_112),
		.b(new_net_29),
		.c(_0191_)
	);

	and_bi _0704_ (
		.a(new_net_113),
		.b(new_net_30),
		.c(_0192_)
	);

	and_bi _0705_ (
		.a(_0191_),
		.b(_0192_),
		.c(_0193_)
	);

	and_bi _0706_ (
		.a(new_net_827),
		.b(new_net_631),
		.c(_0194_)
	);

	and_bi _0707_ (
		.a(new_net_828),
		.b(new_net_543),
		.c(_0195_)
	);

	and_bi _0708_ (
		.a(_0194_),
		.b(_0195_),
		.c(_0196_)
	);

	and_bi _0709_ (
		.a(new_net_829),
		.b(new_net_126),
		.c(_0197_)
	);

	and_bi _0710_ (
		.a(new_net_830),
		.b(new_net_179),
		.c(_0198_)
	);

	or_bb _0711_ (
		.a(_0198_),
		.b(_0197_),
		.c(_0199_)
	);

	and_bi _0712_ (
		.a(_0196_),
		.b(_0199_),
		.c(_0200_)
	);

	and_bi _0713_ (
		.a(new_net_258),
		.b(new_net_427),
		.c(_0201_)
	);

	and_bi _0714_ (
		.a(new_net_255),
		.b(new_net_425),
		.c(_0202_)
	);

	and_bi _0715_ (
		.a(_0201_),
		.b(_0202_),
		.c(_0203_)
	);

	and_bi _0716_ (
		.a(new_net_42),
		.b(new_net_387),
		.c(_0204_)
	);

	and_bi _0717_ (
		.a(new_net_43),
		.b(new_net_388),
		.c(_0205_)
	);

	or_bb _0718_ (
		.a(_0205_),
		.b(_0204_),
		.c(_0206_)
	);

	and_ii _0719_ (
		.a(new_net_70),
		.b(new_net_544),
		.c(_0207_)
	);

	and_bb _0720_ (
		.a(new_net_71),
		.b(new_net_545),
		.c(_0208_)
	);

	or_bb _0721_ (
		.a(_0208_),
		.b(new_net_324),
		.c(_0209_)
	);

	and_bi _0722_ (
		.a(new_net_831),
		.b(_0209_),
		.c(new_net_15)
	);

	and_bi _0723_ (
		.a(new_net_172),
		.b(new_net_309),
		.c(_0210_)
	);

	and_bi _0724_ (
		.a(new_net_168),
		.b(new_net_307),
		.c(_0211_)
	);

	and_bi _0725_ (
		.a(_0210_),
		.b(_0211_),
		.c(_0212_)
	);

	and_bi _0726_ (
		.a(new_net_188),
		.b(new_net_286),
		.c(_0213_)
	);

	and_bi _0727_ (
		.a(new_net_287),
		.b(new_net_192),
		.c(_0214_)
	);

	and_bi _0728_ (
		.a(_0213_),
		.b(_0214_),
		.c(_0215_)
	);

	and_bi _0729_ (
		.a(new_net_46),
		.b(new_net_153),
		.c(_0216_)
	);

	and_bi _0730_ (
		.a(new_net_47),
		.b(new_net_154),
		.c(_0217_)
	);

	and_bi _0731_ (
		.a(_0216_),
		.b(_0217_),
		.c(_0218_)
	);

	and_bi _0732_ (
		.a(new_net_403),
		.b(new_net_832),
		.c(_0219_)
	);

	and_bi _0733_ (
		.a(new_net_410),
		.b(new_net_833),
		.c(_0220_)
	);

	or_bb _0734_ (
		.a(_0220_),
		.b(new_net_547),
		.c(_0221_)
	);

	and_bi _0735_ (
		.a(new_net_834),
		.b(_0221_),
		.c(_0222_)
	);

	and_bi _0736_ (
		.a(new_net_835),
		.b(new_net_34),
		.c(_0223_)
	);

	and_bi _0737_ (
		.a(new_net_836),
		.b(new_net_207),
		.c(_0224_)
	);

	or_bb _0738_ (
		.a(_0224_),
		.b(_0223_),
		.c(_0225_)
	);

	and_bi _0739_ (
		.a(new_net_837),
		.b(_0225_),
		.c(_0226_)
	);

	and_bi _0740_ (
		.a(new_net_402),
		.b(new_net_838),
		.c(_0227_)
	);

	and_bi _0741_ (
		.a(new_net_412),
		.b(new_net_839),
		.c(_0228_)
	);

	or_bb _0742_ (
		.a(_0228_),
		.b(new_net_548),
		.c(_0229_)
	);

	and_bi _0743_ (
		.a(new_net_840),
		.b(_0229_),
		.c(_0230_)
	);

	and_bi _0744_ (
		.a(new_net_841),
		.b(new_net_35),
		.c(_0231_)
	);

	and_bi _0745_ (
		.a(new_net_842),
		.b(new_net_208),
		.c(_0232_)
	);

	or_bb _0746_ (
		.a(_0232_),
		.b(_0231_),
		.c(_0233_)
	);

	and_bi _0747_ (
		.a(new_net_843),
		.b(_0233_),
		.c(_0234_)
	);

	and_bi _0748_ (
		.a(new_net_529),
		.b(new_net_77),
		.c(_0235_)
	);

	and_bi _0749_ (
		.a(new_net_532),
		.b(new_net_80),
		.c(_0236_)
	);

	and_bi _0750_ (
		.a(_0235_),
		.b(_0236_),
		.c(_0237_)
	);

	and_ii _0751_ (
		.a(new_net_432),
		.b(new_net_605),
		.c(_0238_)
	);

	and_bb _0752_ (
		.a(new_net_429),
		.b(new_net_600),
		.c(_0239_)
	);

	or_bb _0753_ (
		.a(_0239_),
		.b(_0238_),
		.c(_0240_)
	);

	and_bi _0754_ (
		.a(new_net_398),
		.b(new_net_844),
		.c(_0241_)
	);

	and_bi _0755_ (
		.a(new_net_401),
		.b(new_net_845),
		.c(_0242_)
	);

	or_bb _0756_ (
		.a(_0242_),
		.b(new_net_549),
		.c(_0243_)
	);

	and_bi _0757_ (
		.a(new_net_846),
		.b(_0243_),
		.c(_0244_)
	);

	and_bi _0758_ (
		.a(new_net_847),
		.b(new_net_36),
		.c(_0245_)
	);

	and_bi _0759_ (
		.a(new_net_848),
		.b(new_net_209),
		.c(_0246_)
	);

	or_bb _0760_ (
		.a(_0246_),
		.b(_0245_),
		.c(_0247_)
	);

	and_bi _0761_ (
		.a(new_net_849),
		.b(_0247_),
		.c(_0248_)
	);

	and_ii _0762_ (
		.a(new_net_234),
		.b(new_net_592),
		.c(_0249_)
	);

	and_bb _0763_ (
		.a(new_net_239),
		.b(new_net_595),
		.c(_0250_)
	);

	and_bi _0764_ (
		.a(_0249_),
		.b(_0250_),
		.c(_0251_)
	);

	or_bb _0765_ (
		.a(new_net_577),
		.b(new_net_253),
		.c(_0252_)
	);

	and_bi _0766_ (
		.a(new_net_254),
		.b(new_net_578),
		.c(_0253_)
	);

	and_bi _0767_ (
		.a(_0252_),
		.b(_0253_),
		.c(_0254_)
	);

	or_bb _0768_ (
		.a(new_net_44),
		.b(new_net_474),
		.c(_0255_)
	);

	and_bb _0769_ (
		.a(new_net_45),
		.b(new_net_476),
		.c(_0256_)
	);

	and_bi _0770_ (
		.a(_0255_),
		.b(_0256_),
		.c(_0257_)
	);

	and_bi _0771_ (
		.a(new_net_226),
		.b(new_net_295),
		.c(_0258_)
	);

	and_bi _0772_ (
		.a(new_net_296),
		.b(new_net_227),
		.c(_0259_)
	);

	or_bb _0773_ (
		.a(_0259_),
		.b(new_net_325),
		.c(_0260_)
	);

	and_bi _0774_ (
		.a(new_net_850),
		.b(_0260_),
		.c(new_net_16)
	);

	or_bb _0775_ (
		.a(new_net_620),
		.b(new_net_349),
		.c(new_net_965)
	);

	or_bb _0776_ (
		.a(new_net_851),
		.b(new_net_571),
		.c(_0261_)
	);

	or_bb _0777_ (
		.a(_0261_),
		.b(new_net_852),
		.c(new_net_952)
	);

	or_bb _0778_ (
		.a(new_net_853),
		.b(new_net_572),
		.c(new_net_10)
	);

	or_bb _0779_ (
		.a(new_net_589),
		.b(new_net_468),
		.c(new_net_957)
	);

	or_bb _0780_ (
		.a(new_net_590),
		.b(new_net_155),
		.c(new_net_967)
	);

	and_bi _0781_ (
		.a(new_net_277),
		.b(new_net_31),
		.c(_0262_)
	);

	or_bb _0782_ (
		.a(new_net_335),
		.b(new_net_212),
		.c(_0263_)
	);

	and_bi _0783_ (
		.a(_0262_),
		.b(_0263_),
		.c(_0264_)
	);

	and_bi _0784_ (
		.a(new_net_444),
		.b(new_net_472),
		.c(_0265_)
	);

	or_bb _0785_ (
		.a(new_net_533),
		.b(new_net_198),
		.c(_0266_)
	);

	and_bi _0786_ (
		.a(_0265_),
		.b(_0266_),
		.c(_0267_)
	);

	or_bb _0787_ (
		.a(new_net_389),
		.b(new_net_326),
		.c(new_net_17)
	);

	and_bi _0788_ (
		.a(new_net_156),
		.b(new_net_390),
		.c(_0268_)
	);

	and_bi _0789_ (
		.a(new_net_469),
		.b(new_net_327),
		.c(_0269_)
	);

	or_bb _0790_ (
		.a(_0269_),
		.b(_0268_),
		.c(new_net_11)
	);

	or_bb _0791_ (
		.a(new_net_854),
		.b(new_net_573),
		.c(_0270_)
	);

	or_bb _0792_ (
		.a(new_net_855),
		.b(new_net_299),
		.c(_0271_)
	);

	or_bb _0793_ (
		.a(new_net_499),
		.b(new_net_856),
		.c(new_net_950)
	);

	and_bi _0794_ (
		.a(G1),
		.b(G3),
		.c(_0272_)
	);

	or_bb _0795_ (
		.a(new_net_857),
		.b(new_net_500),
		.c(new_net_946)
	);

	or_bb _0796_ (
		.a(new_net_235),
		.b(new_net_363),
		.c(_0273_)
	);

	and_bi _0797_ (
		.a(new_net_367),
		.b(new_net_433),
		.c(_0274_)
	);

	and_bi _0798_ (
		.a(_0273_),
		.b(new_net_858),
		.c(new_net_18)
	);

	or_bb _0799_ (
		.a(new_net_597),
		.b(new_net_368),
		.c(_0275_)
	);

	and_bi _0800_ (
		.a(new_net_601),
		.b(new_net_365),
		.c(_0276_)
	);

	and_bi _0801_ (
		.a(new_net_859),
		.b(_0276_),
		.c(new_net_19)
	);

	and_bi _0802_ (
		.a(new_net_364),
		.b(new_net_78),
		.c(_0277_)
	);

	or_bb _0803_ (
		.a(new_net_369),
		.b(new_net_526),
		.c(_0278_)
	);

	and_bi _0804_ (
		.a(new_net_236),
		.b(new_net_860),
		.c(_0279_)
	);

	or_bb _0805_ (
		.a(_0279_),
		.b(_0277_),
		.c(new_net_20)
	);

	or_bb _0806_ (
		.a(new_net_83),
		.b(new_net_50),
		.c(_0280_)
	);

	and_bi _0807_ (
		.a(new_net_49),
		.b(new_net_87),
		.c(_0281_)
	);

	and_bi _0808_ (
		.a(_0280_),
		.b(_0281_),
		.c(_0282_)
	);

	or_bb _0809_ (
		.a(_0282_),
		.b(new_net_67),
		.c(new_net_963)
	);

	and_bi _0810_ (
		.a(new_net_131),
		.b(new_net_861),
		.c(_0283_)
	);

	and_bi _0811_ (
		.a(new_net_137),
		.b(new_net_428),
		.c(_0284_)
	);

	and_bi _0812_ (
		.a(new_net_862),
		.b(_0284_),
		.c(_0285_)
	);

	and_bi _0813_ (
		.a(new_net_385),
		.b(new_net_271),
		.c(_0286_)
	);

	and_bi _0814_ (
		.a(new_net_501),
		.b(new_net_863),
		.c(_0287_)
	);

	and_bi _0815_ (
		.a(new_net_504),
		.b(new_net_82),
		.c(_0288_)
	);

	and_bi _0816_ (
		.a(new_net_864),
		.b(_0288_),
		.c(_0289_)
	);

	and_bi _0817_ (
		.a(new_net_76),
		.b(new_net_243),
		.c(_0290_)
	);

	and_bi _0818_ (
		.a(new_net_502),
		.b(new_net_865),
		.c(_0291_)
	);

	and_bi _0819_ (
		.a(new_net_606),
		.b(new_net_514),
		.c(_0292_)
	);

	and_bi _0820_ (
		.a(new_net_866),
		.b(_0292_),
		.c(_0293_)
	);

	and_bi _0821_ (
		.a(new_net_282),
		.b(new_net_224),
		.c(_0294_)
	);

	or_bb _0822_ (
		.a(_0294_),
		.b(_0290_),
		.c(_0295_)
	);

	or_bb _0823_ (
		.a(_0295_),
		.b(new_net_867),
		.c(_0296_)
	);

	and_bi _0824_ (
		.a(new_net_508),
		.b(new_net_868),
		.c(_0297_)
	);

	and_bi _0825_ (
		.a(new_net_515),
		.b(new_net_434),
		.c(_0298_)
	);

	and_bi _0826_ (
		.a(new_net_869),
		.b(_0298_),
		.c(_0299_)
	);

	and_bi _0827_ (
		.a(new_net_217),
		.b(new_net_460),
		.c(_0300_)
	);

	and_bi _0828_ (
		.a(new_net_142),
		.b(new_net_870),
		.c(_0301_)
	);

	and_bi _0829_ (
		.a(new_net_144),
		.b(new_net_257),
		.c(_0302_)
	);

	and_bi _0830_ (
		.a(new_net_871),
		.b(_0302_),
		.c(_0303_)
	);

	and_bi _0831_ (
		.a(new_net_582),
		.b(new_net_247),
		.c(_0304_)
	);

	or_bb _0832_ (
		.a(new_net_872),
		.b(_0300_),
		.c(_0305_)
	);

	and_bi _0833_ (
		.a(new_net_145),
		.b(new_net_873),
		.c(_0306_)
	);

	and_bi _0834_ (
		.a(new_net_132),
		.b(new_net_466),
		.c(_0307_)
	);

	and_bi _0835_ (
		.a(new_net_874),
		.b(_0307_),
		.c(_0308_)
	);

	and_bi _0836_ (
		.a(new_net_25),
		.b(new_net_563),
		.c(_0309_)
	);

	and_bi _0837_ (
		.a(new_net_384),
		.b(new_net_272),
		.c(_0310_)
	);

	or_bb _0838_ (
		.a(_0310_),
		.b(new_net_875),
		.c(_0311_)
	);

	or_bb _0839_ (
		.a(new_net_876),
		.b(_0305_),
		.c(_0312_)
	);

	and_bi _0840_ (
		.a(new_net_509),
		.b(new_net_877),
		.c(_0313_)
	);

	and_bi _0841_ (
		.a(new_net_596),
		.b(new_net_505),
		.c(_0314_)
	);

	and_bi _0842_ (
		.a(new_net_878),
		.b(_0314_),
		.c(_0315_)
	);

	and_bi _0843_ (
		.a(new_net_167),
		.b(new_net_611),
		.c(_0316_)
	);

	and_bi _0844_ (
		.a(new_net_510),
		.b(new_net_879),
		.c(_0317_)
	);

	and_bi _0845_ (
		.a(new_net_516),
		.b(new_net_238),
		.c(_0318_)
	);

	and_bi _0846_ (
		.a(new_net_880),
		.b(_0318_),
		.c(_0319_)
	);

	and_bi _0847_ (
		.a(new_net_197),
		.b(new_net_106),
		.c(_0320_)
	);

	or_bb _0848_ (
		.a(_0320_),
		.b(new_net_881),
		.c(_0321_)
	);

	and_bi _0849_ (
		.a(new_net_146),
		.b(new_net_882),
		.c(_0322_)
	);

	and_bi _0850_ (
		.a(new_net_133),
		.b(new_net_268),
		.c(_0323_)
	);

	and_bi _0851_ (
		.a(new_net_883),
		.b(_0323_),
		.c(_0324_)
	);

	and_bi _0852_ (
		.a(new_net_625),
		.b(new_net_63),
		.c(_0325_)
	);

	and_bi _0853_ (
		.a(new_net_581),
		.b(new_net_248),
		.c(_0326_)
	);

	or_bb _0854_ (
		.a(_0326_),
		.b(_0325_),
		.c(_0327_)
	);

	or_bb _0855_ (
		.a(new_net_884),
		.b(_0321_),
		.c(_0328_)
	);

	or_bb _0856_ (
		.a(_0328_),
		.b(new_net_885),
		.c(_0329_)
	);

	or_bb _0857_ (
		.a(_0329_),
		.b(new_net_886),
		.c(_0330_)
	);

	and_bi _0858_ (
		.a(new_net_134),
		.b(new_net_887),
		.c(_0331_)
	);

	and_bi _0859_ (
		.a(new_net_138),
		.b(new_net_450),
		.c(_0332_)
	);

	and_bi _0860_ (
		.a(new_net_888),
		.b(_0332_),
		.c(_0333_)
	);

	or_bb _0861_ (
		.a(new_net_151),
		.b(new_net_421),
		.c(_0334_)
	);

	and_bi _0862_ (
		.a(new_net_418),
		.b(new_net_152),
		.c(_0335_)
	);

	and_bi _0863_ (
		.a(_0334_),
		.b(_0335_),
		.c(_0336_)
	);

	and_bi _0864_ (
		.a(new_net_511),
		.b(new_net_889),
		.c(_0337_)
	);

	and_bi _0865_ (
		.a(new_net_517),
		.b(new_net_191),
		.c(_0338_)
	);

	and_bi _0866_ (
		.a(new_net_890),
		.b(_0338_),
		.c(_0339_)
	);

	or_bb _0867_ (
		.a(new_net_68),
		.b(new_net_441),
		.c(_0340_)
	);

	and_bi _0868_ (
		.a(new_net_437),
		.b(new_net_69),
		.c(_0341_)
	);

	and_bi _0869_ (
		.a(_0340_),
		.b(_0341_),
		.c(_0342_)
	);

	and_bi _0870_ (
		.a(new_net_135),
		.b(new_net_891),
		.c(_0343_)
	);

	and_bi _0871_ (
		.a(new_net_139),
		.b(new_net_57),
		.c(_0344_)
	);

	and_bi _0872_ (
		.a(new_net_892),
		.b(_0344_),
		.c(_0345_)
	);

	or_bb _0873_ (
		.a(new_net_249),
		.b(new_net_487),
		.c(_0346_)
	);

	and_bi _0874_ (
		.a(new_net_482),
		.b(new_net_250),
		.c(_0347_)
	);

	and_bi _0875_ (
		.a(_0346_),
		.b(_0347_),
		.c(_0348_)
	);

	or_bb _0876_ (
		.a(new_net_893),
		.b(_0342_),
		.c(_0349_)
	);

	or_bb _0877_ (
		.a(_0349_),
		.b(new_net_894),
		.c(_0350_)
	);

	and_bi _0878_ (
		.a(new_net_136),
		.b(new_net_895),
		.c(_0351_)
	);

	and_bi _0879_ (
		.a(new_net_140),
		.b(new_net_561),
		.c(_0352_)
	);

	and_bi _0880_ (
		.a(new_net_896),
		.b(_0352_),
		.c(_0353_)
	);

	and_bi _0881_ (
		.a(new_net_522),
		.b(new_net_607),
		.c(_0354_)
	);

	and_bi _0882_ (
		.a(new_net_280),
		.b(new_net_225),
		.c(_0355_)
	);

	or_bb _0883_ (
		.a(_0355_),
		.b(new_net_897),
		.c(_0356_)
	);

	and_bi _0884_ (
		.a(new_net_194),
		.b(new_net_107),
		.c(_0357_)
	);

	and_bi _0885_ (
		.a(new_net_518),
		.b(new_net_898),
		.c(_0358_)
	);

	and_bi _0886_ (
		.a(new_net_503),
		.b(new_net_169),
		.c(_0359_)
	);

	and_bi _0887_ (
		.a(new_net_899),
		.b(_0359_),
		.c(_0360_)
	);

	and_bi _0888_ (
		.a(new_net_353),
		.b(new_net_91),
		.c(_0361_)
	);

	or_bb _0889_ (
		.a(_0361_),
		.b(_0357_),
		.c(_0362_)
	);

	or_bb _0890_ (
		.a(_0362_),
		.b(_0356_),
		.c(_0363_)
	);

	and_bi _0891_ (
		.a(new_net_506),
		.b(new_net_900),
		.c(_0364_)
	);

	and_bi _0892_ (
		.a(new_net_512),
		.b(new_net_305),
		.c(_0365_)
	);

	and_bi _0893_ (
		.a(new_net_901),
		.b(_0365_),
		.c(_0366_)
	);

	and_bi _0894_ (
		.a(new_net_330),
		.b(new_net_251),
		.c(_0367_)
	);

	and_bi _0895_ (
		.a(new_net_141),
		.b(new_net_86),
		.c(_0368_)
	);

	and_bi _0896_ (
		.a(new_net_143),
		.b(new_net_902),
		.c(_0369_)
	);

	or_bb _0897_ (
		.a(_0369_),
		.b(new_net_903),
		.c(_0370_)
	);

	or_bb _0898_ (
		.a(new_net_904),
		.b(_0368_),
		.c(_0371_)
	);

	or_bb _0899_ (
		.a(new_net_905),
		.b(_0367_),
		.c(_0372_)
	);

	and_bi _0900_ (
		.a(new_net_27),
		.b(new_net_564),
		.c(_0373_)
	);

	and_bi _0901_ (
		.a(new_net_334),
		.b(new_net_252),
		.c(_0374_)
	);

	or_bb _0902_ (
		.a(_0374_),
		.b(new_net_906),
		.c(_0375_)
	);

	or_bb _0903_ (
		.a(_0375_),
		.b(_0372_),
		.c(_0376_)
	);

	or_bb _0904_ (
		.a(new_net_907),
		.b(_0363_),
		.c(_0377_)
	);

	and_bi _0905_ (
		.a(new_net_626),
		.b(new_net_64),
		.c(_0378_)
	);

	and_bi _0906_ (
		.a(new_net_215),
		.b(new_net_461),
		.c(_0379_)
	);

	or_bb _0907_ (
		.a(_0379_),
		.b(new_net_908),
		.c(_0380_)
	);

	and_bi _0908_ (
		.a(new_net_74),
		.b(new_net_244),
		.c(_0381_)
	);

	and_bi _0909_ (
		.a(new_net_166),
		.b(new_net_612),
		.c(_0382_)
	);

	or_bb _0910_ (
		.a(new_net_909),
		.b(_0381_),
		.c(_0383_)
	);

	or_bb _0911_ (
		.a(_0383_),
		.b(new_net_910),
		.c(_0384_)
	);

	and_bi _0912_ (
		.a(new_net_354),
		.b(new_net_92),
		.c(_0385_)
	);

	and_bi _0913_ (
		.a(new_net_523),
		.b(new_net_608),
		.c(_0386_)
	);

	or_bb _0914_ (
		.a(new_net_911),
		.b(_0385_),
		.c(_0387_)
	);

	and_bi _0915_ (
		.a(new_net_507),
		.b(new_net_912),
		.c(_0388_)
	);

	and_bi _0916_ (
		.a(new_net_513),
		.b(new_net_285),
		.c(_0389_)
	);

	and_bi _0917_ (
		.a(new_net_913),
		.b(_0389_),
		.c(_0390_)
	);

	and_bi _0918_ (
		.a(new_net_301),
		.b(new_net_322),
		.c(_0391_)
	);

	and_bi _0919_ (
		.a(new_net_304),
		.b(new_net_323),
		.c(_0392_)
	);

	or_bb _0920_ (
		.a(_0392_),
		.b(_0391_),
		.c(_0393_)
	);

	or_bb _0921_ (
		.a(new_net_914),
		.b(_0387_),
		.c(_0394_)
	);

	or_bb _0922_ (
		.a(_0394_),
		.b(_0384_),
		.c(_0395_)
	);

	or_bb _0923_ (
		.a(_0395_),
		.b(_0377_),
		.c(_0396_)
	);

	or_bb _0924_ (
		.a(_0396_),
		.b(new_net_915),
		.c(_0397_)
	);

	or_bb _0925_ (
		.a(_0397_),
		.b(new_net_916),
		.c(new_net_21)
	);

	and_bi _0926_ (
		.a(new_net_366),
		.b(new_net_530),
		.c(_0398_)
	);

	and_bi _0927_ (
		.a(new_net_528),
		.b(new_net_240),
		.c(_0399_)
	);

	and_bi _0928_ (
		.a(new_net_477),
		.b(new_net_609),
		.c(_0400_)
	);

	and_bi _0929_ (
		.a(new_net_475),
		.b(new_net_610),
		.c(_0401_)
	);

	and_bi _0930_ (
		.a(_0400_),
		.b(_0401_),
		.c(_0402_)
	);

	and_bi _0931_ (
		.a(new_net_229),
		.b(new_net_598),
		.c(_0403_)
	);

	and_bi _0932_ (
		.a(new_net_593),
		.b(new_net_228),
		.c(_0404_)
	);

	and_bi _0933_ (
		.a(_0403_),
		.b(_0404_),
		.c(_0405_)
	);

	or_bb _0934_ (
		.a(new_net_569),
		.b(new_net_88),
		.c(_0406_)
	);

	and_bi _0935_ (
		.a(new_net_90),
		.b(new_net_570),
		.c(_0407_)
	);

	and_bi _0936_ (
		.a(_0406_),
		.b(_0407_),
		.c(_0408_)
	);

	and_bi _0937_ (
		.a(new_net_370),
		.b(_0408_),
		.c(_0409_)
	);

	or_bb _0938_ (
		.a(_0409_),
		.b(new_net_917),
		.c(new_net_22)
	);

	or_bb _0939_ (
		.a(new_net_259),
		.b(new_net_918),
		.c(_0410_)
	);

	or_bb _0940_ (
		.a(new_net_269),
		.b(new_net_919),
		.c(_0411_)
	);

	and_ii _0941_ (
		.a(new_net_219),
		.b(new_net_574),
		.c(_0412_)
	);

	or_bb _0942_ (
		.a(new_net_358),
		.b(new_net_127),
		.c(_0413_)
	);

	or_bb _0943_ (
		.a(new_net_491),
		.b(new_net_333),
		.c(_0414_)
	);

	or_bb _0944_ (
		.a(new_net_220),
		.b(new_net_576),
		.c(_0415_)
	);

	or_bb _0945_ (
		.a(new_net_453),
		.b(new_net_130),
		.c(_0416_)
	);

	or_bb _0946_ (
		.a(new_net_478),
		.b(new_net_306),
		.c(_0417_)
	);

	or_bb _0947_ (
		.a(new_net_492),
		.b(new_net_303),
		.c(_0418_)
	);

	and_bi _0948_ (
		.a(new_net_216),
		.b(new_net_359),
		.c(_0419_)
	);

	and_bi _0949_ (
		.a(new_net_583),
		.b(new_net_455),
		.c(_0420_)
	);

	and_bi _0950_ (
		.a(_0419_),
		.b(_0420_),
		.c(_0421_)
	);

	and_bi _0951_ (
		.a(new_net_435),
		.b(new_net_415),
		.c(_0422_)
	);

	or_bb _0952_ (
		.a(new_net_362),
		.b(new_net_164),
		.c(_0423_)
	);

	and_bi _0953_ (
		.a(new_net_521),
		.b(new_net_456),
		.c(_0424_)
	);

	and_bi _0954_ (
		.a(_0423_),
		.b(_0424_),
		.c(_0425_)
	);

	or_bb _0955_ (
		.a(new_net_375),
		.b(new_net_599),
		.c(_0426_)
	);

	or_bb _0956_ (
		.a(new_net_360),
		.b(new_net_196),
		.c(_0427_)
	);

	and_bi _0957_ (
		.a(new_net_486),
		.b(new_net_457),
		.c(_0428_)
	);

	and_bi _0958_ (
		.a(_0427_),
		.b(_0428_),
		.c(_0429_)
	);

	and_bi _0959_ (
		.a(new_net_337),
		.b(new_net_241),
		.c(_0430_)
	);

	or_bb _0960_ (
		.a(new_net_361),
		.b(new_net_73),
		.c(_0431_)
	);

	and_bi _0961_ (
		.a(new_net_420),
		.b(new_net_454),
		.c(_0432_)
	);

	and_bi _0962_ (
		.a(_0431_),
		.b(_0432_),
		.c(_0433_)
	);

	or_bb _0963_ (
		.a(_0433_),
		.b(new_net_81),
		.c(_0434_)
	);

	or_bb _0964_ (
		.a(new_net_920),
		.b(_0430_),
		.c(_0435_)
	);

	and_bi _0965_ (
		.a(new_net_242),
		.b(new_net_338),
		.c(_0436_)
	);

	and_bi _0966_ (
		.a(new_net_594),
		.b(new_net_376),
		.c(_0437_)
	);

	or_bb _0967_ (
		.a(_0437_),
		.b(_0436_),
		.c(_0438_)
	);

	and_bi _0968_ (
		.a(_0435_),
		.b(_0438_),
		.c(_0439_)
	);

	and_bi _0969_ (
		.a(new_net_921),
		.b(_0439_),
		.c(_0440_)
	);

	or_bb _0970_ (
		.a(_0440_),
		.b(new_net_922),
		.c(_0441_)
	);

	and_bi _0971_ (
		.a(new_net_436),
		.b(new_net_416),
		.c(_0442_)
	);

	and_bi _0972_ (
		.a(new_net_129),
		.b(new_net_602),
		.c(_0443_)
	);

	and_bi _0973_ (
		.a(new_net_283),
		.b(new_net_493),
		.c(_0444_)
	);

	and_bi _0974_ (
		.a(new_net_624),
		.b(new_net_480),
		.c(_0445_)
	);

	and_bi _0975_ (
		.a(_0444_),
		.b(_0445_),
		.c(_0446_)
	);

	and_bi _0976_ (
		.a(new_net_61),
		.b(new_net_147),
		.c(_0447_)
	);

	or_bb _0977_ (
		.a(_0447_),
		.b(new_net_923),
		.c(_0448_)
	);

	and_bi _0978_ (
		.a(_0441_),
		.b(new_net_924),
		.c(_0449_)
	);

	and_bi _0979_ (
		.a(new_net_62),
		.b(new_net_148),
		.c(_0450_)
	);

	and_bi _0980_ (
		.a(new_net_128),
		.b(new_net_189),
		.c(_0451_)
	);

	and_bi _0981_ (
		.a(new_net_440),
		.b(new_net_494),
		.c(_0452_)
	);

	and_bi _0982_ (
		.a(new_net_26),
		.b(new_net_479),
		.c(_0453_)
	);

	and_bi _0983_ (
		.a(_0452_),
		.b(_0453_),
		.c(_0454_)
	);

	and_bi _0984_ (
		.a(new_net_275),
		.b(new_net_584),
		.c(_0455_)
	);

	or_bb _0985_ (
		.a(_0455_),
		.b(_0450_),
		.c(_0456_)
	);

	or_bb _0986_ (
		.a(new_net_925),
		.b(_0449_),
		.c(_0457_)
	);

	and_bi _0987_ (
		.a(new_net_288),
		.b(new_net_481),
		.c(_0458_)
	);

	and_bi _0988_ (
		.a(new_net_276),
		.b(new_net_585),
		.c(_0459_)
	);

	or_bb _0989_ (
		.a(_0459_),
		.b(new_net_926),
		.c(_0460_)
	);

	and_bi _0990_ (
		.a(_0457_),
		.b(new_net_927),
		.c(_0461_)
	);

	and_bi _0991_ (
		.a(new_net_928),
		.b(_0461_),
		.c(_0462_)
	);

	and_bi _0992_ (
		.a(new_net_929),
		.b(_0462_),
		.c(_0463_)
	);

	and_bi _0993_ (
		.a(new_net_930),
		.b(_0463_),
		.c(_0464_)
	);

	and_bi _0994_ (
		.a(new_net_575),
		.b(new_net_221),
		.c(_0465_)
	);

	or_bb _0995_ (
		.a(new_net_451),
		.b(new_net_422),
		.c(_0466_)
	);

	and_bi _0996_ (
		.a(new_net_314),
		.b(new_net_931),
		.c(_0467_)
	);

	or_bb _0997_ (
		.a(new_net_58),
		.b(new_net_488),
		.c(_0468_)
	);

	and_bi _0998_ (
		.a(new_net_316),
		.b(new_net_932),
		.c(_0469_)
	);

	and_bi _0999_ (
		.a(_0467_),
		.b(_0469_),
		.c(_0470_)
	);

	or_bb _1000_ (
		.a(new_net_54),
		.b(new_net_484),
		.c(_0471_)
	);

	and_bi _1001_ (
		.a(new_net_318),
		.b(new_net_933),
		.c(_0472_)
	);

	or_bb _1002_ (
		.a(new_net_426),
		.b(new_net_382),
		.c(_0473_)
	);

	and_bi _1003_ (
		.a(new_net_356),
		.b(new_net_171),
		.c(_0474_)
	);

	and_bi _1004_ (
		.a(new_net_293),
		.b(_0474_),
		.c(_0475_)
	);

	and_bi _1005_ (
		.a(new_net_319),
		.b(_0475_),
		.c(_0476_)
	);

	and_ii _1006_ (
		.a(new_net_934),
		.b(new_net_104),
		.c(_0477_)
	);

	or_bb _1007_ (
		.a(new_net_452),
		.b(new_net_423),
		.c(_0478_)
	);

	and_bi _1008_ (
		.a(new_net_383),
		.b(new_net_424),
		.c(_0479_)
	);

	and_bi _1009_ (
		.a(new_net_935),
		.b(_0479_),
		.c(_0480_)
	);

	and_bi _1010_ (
		.a(new_net_315),
		.b(new_net_936),
		.c(_0481_)
	);

	or_bb _1011_ (
		.a(new_net_173),
		.b(new_net_357),
		.c(_0482_)
	);

	and_bi _1012_ (
		.a(new_net_317),
		.b(new_net_937),
		.c(_0483_)
	);

	or_bb _1013_ (
		.a(new_net_617),
		.b(new_net_558),
		.c(_0484_)
	);

	and_bi _1014_ (
		.a(_0477_),
		.b(_0484_),
		.c(_0485_)
	);

	or_ii _1015_ (
		.a(_0485_),
		.b(new_net_230),
		.c(_0486_)
	);

	or_bb _1016_ (
		.a(new_net_938),
		.b(_0464_),
		.c(_0487_)
	);

	and_bi _1017_ (
		.a(new_net_294),
		.b(new_net_618),
		.c(_0488_)
	);

	and_bi _1018_ (
		.a(new_net_559),
		.b(_0488_),
		.c(_0489_)
	);

	and_bi _1019_ (
		.a(new_net_231),
		.b(_0489_),
		.c(_0490_)
	);

	or_bb _1020_ (
		.a(_0490_),
		.b(new_net_105),
		.c(_0491_)
	);

	and_bi _1021_ (
		.a(_0487_),
		.b(new_net_939),
		.c(G2591)
	);

	or_bb _1022_ (
		.a(new_net_298),
		.b(new_net_321),
		.c(_0492_)
	);

	or_bb _1023_ (
		.a(new_net_940),
		.b(new_net_150),
		.c(_0493_)
	);

	or_bb _1024_ (
		.a(_0493_),
		.b(new_net_60),
		.c(_0494_)
	);

	or_bb _1025_ (
		.a(new_net_941),
		.b(new_net_587),
		.c(_0495_)
	);

	or_bb _1026_ (
		.a(new_net_942),
		.b(new_net_211),
		.c(new_net_23)
	);

	and_bi _1027_ (
		.a(new_net_347),
		.b(new_net_943),
		.c(new_net_954)
	);

	or_bb _1028_ (
		.a(new_net_79),
		.b(new_net_613),
		.c(new_net_948)
	);

	and_bi _1029_ (
		.a(new_net_527),
		.b(new_net_615),
		.c(_0496_)
	);

	or_bb _1030_ (
		.a(new_net_944),
		.b(new_net_237),
		.c(new_net_961)
	);

	and_bi _1031_ (
		.a(new_net_616),
		.b(new_net_89),
		.c(_0497_)
	);

	and_bi _1032_ (
		.a(new_net_614),
		.b(new_net_531),
		.c(_0498_)
	);

	or_bb _1033_ (
		.a(new_net_945),
		.b(_0497_),
		.c(new_net_959)
	);

	spl2 new_net_724_v_fanout (
		.a(new_net_724),
		.b(G2569),
		.c(G2560)
	);

	spl2 new_net_733_v_fanout (
		.a(new_net_733),
		.b(G2561),
		.c(G2568)
	);

	spl2 new_net_738_v_fanout (
		.a(new_net_738),
		.b(G2562),
		.c(G2567)
	);

	spl4L new_net_672_v_fanout (
		.a(new_net_672),
		.b(G2533),
		.c(G2549),
		.d(G2532),
		.e(G2531)
	);

	bfr new_net_969_bfr_after (
		.din(new_net_23),
		.dout(new_net_969)
	);

	bfr new_net_970_bfr_after (
		.din(new_net_969),
		.dout(new_net_970)
	);

	bfr new_net_971_bfr_after (
		.din(new_net_970),
		.dout(new_net_971)
	);

	spl2 new_net_23_v_fanout (
		.a(new_net_971),
		.b(G2594),
		.c(G2593)
	);

	bfr new_net_972_bfr_after (
		.din(new_net_22),
		.dout(new_net_972)
	);

	bfr new_net_973_bfr_after (
		.din(new_net_972),
		.dout(new_net_973)
	);

	bfr new_net_974_bfr_after (
		.din(new_net_973),
		.dout(new_net_974)
	);

	bfr new_net_975_bfr_after (
		.din(new_net_974),
		.dout(new_net_975)
	);

	spl2 new_net_22_v_fanout (
		.a(new_net_975),
		.b(G2589),
		.c(G2588)
	);

	bfr new_net_976_bfr_before (
		.din(new_net_976),
		.dout(G2590)
	);

	bfr new_net_977_bfr_before (
		.din(new_net_977),
		.dout(new_net_976)
	);

	bfr new_net_978_bfr_before (
		.din(new_net_978),
		.dout(new_net_977)
	);

	bfr new_net_979_bfr_before (
		.din(new_net_979),
		.dout(new_net_978)
	);

	bfr new_net_980_bfr_before (
		.din(new_net_980),
		.dout(new_net_979)
	);

	spl2 new_net_16_v_fanout (
		.a(new_net_16),
		.b(new_net_211),
		.c(new_net_980)
	);

	bfr new_net_981_bfr_after (
		.din(new_net_21),
		.dout(new_net_981)
	);

	bfr new_net_982_bfr_after (
		.din(new_net_981),
		.dout(new_net_982)
	);

	bfr new_net_983_bfr_after (
		.din(new_net_982),
		.dout(new_net_983)
	);

	bfr new_net_984_bfr_after (
		.din(new_net_983),
		.dout(new_net_984)
	);

	bfr new_net_985_bfr_after (
		.din(new_net_984),
		.dout(new_net_985)
	);

	bfr new_net_986_bfr_after (
		.din(new_net_985),
		.dout(new_net_986)
	);

	bfr new_net_987_bfr_after (
		.din(new_net_986),
		.dout(new_net_987)
	);

	spl2 new_net_21_v_fanout (
		.a(new_net_987),
		.b(G2585),
		.c(G2584)
	);

	bfr new_net_988_bfr_before (
		.din(new_net_988),
		.dout(G2587)
	);

	bfr new_net_989_bfr_before (
		.din(new_net_989),
		.dout(new_net_988)
	);

	bfr new_net_990_bfr_before (
		.din(new_net_990),
		.dout(new_net_989)
	);

	bfr new_net_991_bfr_before (
		.din(new_net_991),
		.dout(new_net_990)
	);

	bfr new_net_992_bfr_before (
		.din(new_net_992),
		.dout(new_net_991)
	);

	bfr new_net_993_bfr_before (
		.din(new_net_993),
		.dout(new_net_992)
	);

	bfr new_net_994_bfr_before (
		.din(new_net_994),
		.dout(new_net_993)
	);

	spl2 new_net_15_v_fanout (
		.a(new_net_15),
		.b(new_net_587),
		.c(new_net_994)
	);

	spl2 new_net_749_v_fanout (
		.a(new_net_749),
		.b(new_net_227),
		.c(new_net_226)
	);

	spl2 _0257__v_fanout (
		.a(_0257_),
		.b(new_net_296),
		.c(new_net_295)
	);

	spl2 new_net_748_v_fanout (
		.a(new_net_748),
		.b(new_net_90),
		.c(new_net_88)
	);

	spl2 _0405__v_fanout (
		.a(_0405_),
		.b(new_net_570),
		.c(new_net_569)
	);

	spl2 _0446__v_fanout (
		.a(_0446_),
		.b(new_net_148),
		.c(new_net_147)
	);

	spl2 _0206__v_fanout (
		.a(_0206_),
		.b(new_net_71),
		.c(new_net_70)
	);

	spl2 _0454__v_fanout (
		.a(_0454_),
		.b(new_net_585),
		.c(new_net_584)
	);

	bfr new_net_995_bfr_before (
		.din(new_net_995),
		.dout(new_net_748)
	);

	bfr new_net_996_bfr_before (
		.din(new_net_996),
		.dout(new_net_995)
	);

	spl2 _0402__v_fanout (
		.a(_0402_),
		.b(new_net_996),
		.c(new_net_89)
	);

	spl2 _0254__v_fanout (
		.a(_0254_),
		.b(new_net_45),
		.c(new_net_44)
	);

	bfr new_net_997_bfr_before (
		.din(new_net_997),
		.dout(new_net_749)
	);

	bfr new_net_998_bfr_before (
		.din(new_net_998),
		.dout(new_net_997)
	);

	spl3L _0218__v_fanout (
		.a(_0218_),
		.b(new_net_228),
		.c(new_net_998),
		.d(new_net_229)
	);

	bfr new_net_999_bfr_before (
		.din(new_net_999),
		.dout(G2566)
	);

	bfr new_net_1000_bfr_before (
		.din(new_net_1000),
		.dout(new_net_999)
	);

	bfr new_net_1001_bfr_before (
		.din(new_net_1001),
		.dout(new_net_1000)
	);

	bfr new_net_1002_bfr_before (
		.din(new_net_1002),
		.dout(new_net_1001)
	);

	bfr new_net_1003_bfr_before (
		.din(new_net_1003),
		.dout(new_net_1002)
	);

	bfr new_net_1004_bfr_before (
		.din(new_net_1004),
		.dout(new_net_1003)
	);

	bfr new_net_1005_bfr_before (
		.din(new_net_1005),
		.dout(new_net_1004)
	);

	bfr new_net_1006_bfr_before (
		.din(new_net_1006),
		.dout(new_net_1005)
	);

	bfr new_net_1007_bfr_before (
		.din(new_net_1007),
		.dout(new_net_1006)
	);

	bfr new_net_1008_bfr_before (
		.din(new_net_1008),
		.dout(new_net_1007)
	);

	bfr new_net_1009_bfr_before (
		.din(new_net_1009),
		.dout(new_net_1008)
	);

	bfr new_net_1010_bfr_before (
		.din(new_net_1010),
		.dout(new_net_1009)
	);

	spl3L new_net_729_v_fanout (
		.a(new_net_729),
		.b(new_net_593),
		.c(new_net_1010),
		.d(new_net_598)
	);

	spl2 new_net_747_v_fanout (
		.a(new_net_747),
		.b(new_net_476),
		.c(new_net_474)
	);

	spl2 _0425__v_fanout (
		.a(_0425_),
		.b(new_net_376),
		.c(new_net_375)
	);

	spl2 _0429__v_fanout (
		.a(_0429_),
		.b(new_net_338),
		.c(new_net_337)
	);

	spl2 _0421__v_fanout (
		.a(_0421_),
		.b(new_net_416),
		.c(new_net_415)
	);

	bfr new_net_1011_bfr_after (
		.din(_0470_),
		.dout(new_net_1011)
	);

	spl2 _0470__v_fanout (
		.a(new_net_1011),
		.b(new_net_231),
		.c(new_net_230)
	);

	bfr new_net_1012_bfr_after (
		.din(_0156_),
		.dout(new_net_1012)
	);

	bfr new_net_1013_bfr_after (
		.din(new_net_1012),
		.dout(new_net_1013)
	);

	bfr new_net_1014_bfr_after (
		.din(new_net_1013),
		.dout(new_net_1014)
	);

	spl2 _0156__v_fanout (
		.a(new_net_1014),
		.b(new_net_545),
		.c(new_net_544)
	);

	bfr new_net_1015_bfr_before (
		.din(new_net_1015),
		.dout(new_net_738)
	);

	bfr new_net_1016_bfr_before (
		.din(new_net_1016),
		.dout(new_net_1015)
	);

	bfr new_net_1017_bfr_before (
		.din(new_net_1017),
		.dout(new_net_1016)
	);

	bfr new_net_1018_bfr_before (
		.din(new_net_1018),
		.dout(new_net_1017)
	);

	bfr new_net_1019_bfr_before (
		.din(new_net_1019),
		.dout(new_net_1018)
	);

	bfr new_net_1020_bfr_before (
		.din(new_net_1020),
		.dout(new_net_1019)
	);

	bfr new_net_1021_bfr_before (
		.din(new_net_1021),
		.dout(new_net_1020)
	);

	bfr new_net_1022_bfr_before (
		.din(new_net_1022),
		.dout(new_net_1021)
	);

	bfr new_net_1023_bfr_before (
		.din(new_net_1023),
		.dout(new_net_1022)
	);

	bfr new_net_1024_bfr_before (
		.din(new_net_1024),
		.dout(new_net_1023)
	);

	bfr new_net_1025_bfr_before (
		.din(new_net_1025),
		.dout(new_net_1024)
	);

	bfr new_net_1026_bfr_before (
		.din(new_net_1026),
		.dout(new_net_1025)
	);

	spl3L new_net_737_v_fanout (
		.a(new_net_737),
		.b(new_net_435),
		.c(new_net_436),
		.d(new_net_1026)
	);

	bfr new_net_1027_bfr_before (
		.din(new_net_1027),
		.dout(new_net_559)
	);

	spl2 _0481__v_fanout (
		.a(_0481_),
		.b(new_net_1027),
		.c(new_net_558)
	);

	spl3L new_net_728_v_fanout (
		.a(new_net_728),
		.b(new_net_599),
		.c(new_net_594),
		.d(new_net_729)
	);

	spl2 _0193__v_fanout (
		.a(_0193_),
		.b(new_net_43),
		.c(new_net_42)
	);

	spl2 new_net_721_v_fanout (
		.a(new_net_721),
		.b(new_net_242),
		.c(new_net_241)
	);

	bfr new_net_1028_bfr_before (
		.din(new_net_1028),
		.dout(new_net_105)
	);

	bfr new_net_1029_bfr_before (
		.din(new_net_1029),
		.dout(new_net_1028)
	);

	bfr new_net_1030_bfr_before (
		.din(new_net_1030),
		.dout(new_net_1029)
	);

	spl2 _0472__v_fanout (
		.a(_0472_),
		.b(new_net_1030),
		.c(new_net_104)
	);

	spl4L _0416__v_fanout (
		.a(_0416_),
		.b(new_net_480),
		.c(new_net_478),
		.d(new_net_481),
		.e(new_net_479)
	);

	spl4L _0413__v_fanout (
		.a(_0413_),
		.b(new_net_494),
		.c(new_net_491),
		.d(new_net_493),
		.e(new_net_492)
	);

	spl2 _0483__v_fanout (
		.a(_0483_),
		.b(new_net_618),
		.c(new_net_617)
	);

	bfr new_net_1031_bfr_after (
		.din(new_net_18),
		.dout(new_net_1031)
	);

	bfr new_net_1032_bfr_after (
		.din(new_net_1031),
		.dout(new_net_1032)
	);

	bfr new_net_1033_bfr_after (
		.din(new_net_1032),
		.dout(new_net_1033)
	);

	bfr new_net_1034_bfr_after (
		.din(new_net_1033),
		.dout(new_net_1034)
	);

	bfr new_net_1035_bfr_after (
		.din(new_net_1034),
		.dout(new_net_1035)
	);

	bfr new_net_1036_bfr_after (
		.din(new_net_1035),
		.dout(new_net_1036)
	);

	bfr new_net_1037_bfr_after (
		.din(new_net_1036),
		.dout(new_net_1037)
	);

	bfr new_net_1038_bfr_after (
		.din(new_net_1037),
		.dout(new_net_1038)
	);

	bfr new_net_1039_bfr_after (
		.din(new_net_1038),
		.dout(new_net_1039)
	);

	bfr new_net_1040_bfr_after (
		.din(new_net_1039),
		.dout(new_net_1040)
	);

	bfr new_net_1041_bfr_after (
		.din(new_net_1040),
		.dout(new_net_1041)
	);

	bfr new_net_1042_bfr_after (
		.din(new_net_1041),
		.dout(new_net_1042)
	);

	bfr new_net_1043_bfr_after (
		.din(new_net_1042),
		.dout(new_net_1043)
	);

	bfr new_net_1044_bfr_after (
		.din(new_net_1043),
		.dout(new_net_1044)
	);

	bfr new_net_1045_bfr_after (
		.din(new_net_1044),
		.dout(new_net_1045)
	);

	spl2 new_net_18_v_fanout (
		.a(new_net_1045),
		.b(G2574),
		.c(G2573)
	);

	bfr new_net_1046_bfr_before (
		.din(new_net_1046),
		.dout(new_net_747)
	);

	bfr new_net_1047_bfr_before (
		.din(new_net_1047),
		.dout(new_net_1046)
	);

	spl3L _0237__v_fanout (
		.a(_0237_),
		.b(new_net_477),
		.c(new_net_475),
		.d(new_net_1047)
	);

	spl2 _0240__v_fanout (
		.a(_0240_),
		.b(new_net_254),
		.c(new_net_253)
	);

	bfr new_net_1048_bfr_after (
		.din(new_net_20),
		.dout(new_net_1048)
	);

	bfr new_net_1049_bfr_after (
		.din(new_net_1048),
		.dout(new_net_1049)
	);

	bfr new_net_1050_bfr_after (
		.din(new_net_1049),
		.dout(new_net_1050)
	);

	bfr new_net_1051_bfr_after (
		.din(new_net_1050),
		.dout(new_net_1051)
	);

	bfr new_net_1052_bfr_after (
		.din(new_net_1051),
		.dout(new_net_1052)
	);

	bfr new_net_1053_bfr_after (
		.din(new_net_1052),
		.dout(new_net_1053)
	);

	bfr new_net_1054_bfr_after (
		.din(new_net_1053),
		.dout(new_net_1054)
	);

	bfr new_net_1055_bfr_after (
		.din(new_net_1054),
		.dout(new_net_1055)
	);

	bfr new_net_1056_bfr_after (
		.din(new_net_1055),
		.dout(new_net_1056)
	);

	bfr new_net_1057_bfr_after (
		.din(new_net_1056),
		.dout(new_net_1057)
	);

	bfr new_net_1058_bfr_after (
		.din(new_net_1057),
		.dout(new_net_1058)
	);

	bfr new_net_1059_bfr_after (
		.din(new_net_1058),
		.dout(new_net_1059)
	);

	bfr new_net_1060_bfr_after (
		.din(new_net_1059),
		.dout(new_net_1060)
	);

	bfr new_net_1061_bfr_after (
		.din(new_net_1060),
		.dout(new_net_1061)
	);

	bfr new_net_1062_bfr_after (
		.din(new_net_1061),
		.dout(new_net_1062)
	);

	spl2 new_net_20_v_fanout (
		.a(new_net_1062),
		.b(G2579),
		.c(G2578)
	);

	spl2 _0251__v_fanout (
		.a(_0251_),
		.b(new_net_578),
		.c(new_net_577)
	);

	spl2 _0319__v_fanout (
		.a(_0319_),
		.b(new_net_107),
		.c(new_net_106)
	);

	bfr new_net_1063_bfr_before (
		.din(new_net_1063),
		.dout(G2571)
	);

	bfr new_net_1064_bfr_before (
		.din(new_net_1064),
		.dout(new_net_1063)
	);

	bfr new_net_1065_bfr_before (
		.din(new_net_1065),
		.dout(new_net_1064)
	);

	bfr new_net_1066_bfr_before (
		.din(new_net_1066),
		.dout(new_net_1065)
	);

	bfr new_net_1067_bfr_before (
		.din(new_net_1067),
		.dout(new_net_1066)
	);

	bfr new_net_1068_bfr_before (
		.din(new_net_1068),
		.dout(new_net_1067)
	);

	bfr new_net_1069_bfr_before (
		.din(new_net_1069),
		.dout(new_net_1068)
	);

	bfr new_net_1070_bfr_before (
		.din(new_net_1070),
		.dout(new_net_1069)
	);

	bfr new_net_1071_bfr_before (
		.din(new_net_1071),
		.dout(new_net_1070)
	);

	bfr new_net_1072_bfr_before (
		.din(new_net_1072),
		.dout(new_net_1071)
	);

	bfr new_net_1073_bfr_before (
		.din(new_net_1073),
		.dout(new_net_1072)
	);

	bfr new_net_1074_bfr_before (
		.din(new_net_1074),
		.dout(new_net_1073)
	);

	bfr new_net_1075_bfr_before (
		.din(new_net_1075),
		.dout(new_net_1074)
	);

	bfr new_net_1076_bfr_before (
		.din(new_net_1076),
		.dout(new_net_1075)
	);

	spl2 new_net_730_v_fanout (
		.a(new_net_730),
		.b(new_net_306),
		.c(new_net_1076)
	);

	spl2 _0289__v_fanout (
		.a(_0289_),
		.b(new_net_244),
		.c(new_net_243)
	);

	bfr new_net_1077_bfr_after (
		.din(new_net_19),
		.dout(new_net_1077)
	);

	bfr new_net_1078_bfr_after (
		.din(new_net_1077),
		.dout(new_net_1078)
	);

	bfr new_net_1079_bfr_after (
		.din(new_net_1078),
		.dout(new_net_1079)
	);

	bfr new_net_1080_bfr_after (
		.din(new_net_1079),
		.dout(new_net_1080)
	);

	bfr new_net_1081_bfr_after (
		.din(new_net_1080),
		.dout(new_net_1081)
	);

	bfr new_net_1082_bfr_after (
		.din(new_net_1081),
		.dout(new_net_1082)
	);

	bfr new_net_1083_bfr_after (
		.din(new_net_1082),
		.dout(new_net_1083)
	);

	bfr new_net_1084_bfr_after (
		.din(new_net_1083),
		.dout(new_net_1084)
	);

	bfr new_net_1085_bfr_after (
		.din(new_net_1084),
		.dout(new_net_1085)
	);

	bfr new_net_1086_bfr_after (
		.din(new_net_1085),
		.dout(new_net_1086)
	);

	bfr new_net_1087_bfr_after (
		.din(new_net_1086),
		.dout(new_net_1087)
	);

	bfr new_net_1088_bfr_after (
		.din(new_net_1087),
		.dout(new_net_1088)
	);

	bfr new_net_1089_bfr_after (
		.din(new_net_1088),
		.dout(new_net_1089)
	);

	bfr new_net_1090_bfr_after (
		.din(new_net_1089),
		.dout(new_net_1090)
	);

	bfr new_net_1091_bfr_after (
		.din(new_net_1090),
		.dout(new_net_1091)
	);

	spl2 new_net_19_v_fanout (
		.a(new_net_1091),
		.b(G2576),
		.c(G2575)
	);

	spl2 _0339__v_fanout (
		.a(_0339_),
		.b(new_net_69),
		.c(new_net_68)
	);

	bfr new_net_1092_bfr_before (
		.din(new_net_1092),
		.dout(G2570)
	);

	bfr new_net_1093_bfr_before (
		.din(new_net_1093),
		.dout(new_net_1092)
	);

	bfr new_net_1094_bfr_before (
		.din(new_net_1094),
		.dout(new_net_1093)
	);

	bfr new_net_1095_bfr_before (
		.din(new_net_1095),
		.dout(new_net_1094)
	);

	bfr new_net_1096_bfr_before (
		.din(new_net_1096),
		.dout(new_net_1095)
	);

	bfr new_net_1097_bfr_before (
		.din(new_net_1097),
		.dout(new_net_1096)
	);

	bfr new_net_1098_bfr_before (
		.din(new_net_1098),
		.dout(new_net_1097)
	);

	bfr new_net_1099_bfr_before (
		.din(new_net_1099),
		.dout(new_net_1098)
	);

	bfr new_net_1100_bfr_before (
		.din(new_net_1100),
		.dout(new_net_1099)
	);

	bfr new_net_1101_bfr_before (
		.din(new_net_1101),
		.dout(new_net_1100)
	);

	bfr new_net_1102_bfr_before (
		.din(new_net_1102),
		.dout(new_net_1101)
	);

	bfr new_net_1103_bfr_before (
		.din(new_net_1103),
		.dout(new_net_1102)
	);

	bfr new_net_1104_bfr_before (
		.din(new_net_1104),
		.dout(new_net_1103)
	);

	bfr new_net_1105_bfr_before (
		.din(new_net_1105),
		.dout(new_net_1104)
	);

	spl2 new_net_720_v_fanout (
		.a(new_net_720),
		.b(new_net_288),
		.c(new_net_1105)
	);

	spl2 _0360__v_fanout (
		.a(_0360_),
		.b(new_net_92),
		.c(new_net_91)
	);

	spl2 _0293__v_fanout (
		.a(_0293_),
		.b(new_net_225),
		.c(new_net_224)
	);

	bfr new_net_1106_bfr_before (
		.din(new_net_1106),
		.dout(G2581)
	);

	bfr new_net_1107_bfr_before (
		.din(new_net_1107),
		.dout(new_net_1106)
	);

	bfr new_net_1108_bfr_before (
		.din(new_net_1108),
		.dout(new_net_1107)
	);

	bfr new_net_1109_bfr_before (
		.din(new_net_1109),
		.dout(new_net_1108)
	);

	bfr new_net_1110_bfr_before (
		.din(new_net_1110),
		.dout(new_net_1109)
	);

	bfr new_net_1111_bfr_before (
		.din(new_net_1111),
		.dout(new_net_1110)
	);

	bfr new_net_1112_bfr_before (
		.din(new_net_1112),
		.dout(new_net_1111)
	);

	bfr new_net_1113_bfr_before (
		.din(new_net_1113),
		.dout(new_net_1112)
	);

	bfr new_net_1114_bfr_before (
		.din(new_net_1114),
		.dout(new_net_1113)
	);

	bfr new_net_1115_bfr_before (
		.din(new_net_1115),
		.dout(new_net_1114)
	);

	bfr new_net_1116_bfr_before (
		.din(new_net_1116),
		.dout(new_net_1115)
	);

	bfr new_net_1117_bfr_before (
		.din(new_net_1117),
		.dout(new_net_1116)
	);

	bfr new_net_1118_bfr_before (
		.din(new_net_1118),
		.dout(new_net_1117)
	);

	bfr new_net_1119_bfr_before (
		.din(new_net_1119),
		.dout(new_net_1118)
	);

	bfr new_net_1120_bfr_before (
		.din(new_net_1120),
		.dout(new_net_1119)
	);

	spl2 new_net_14_v_fanout (
		.a(new_net_14),
		.b(new_net_60),
		.c(new_net_1120)
	);

	spl2 _0215__v_fanout (
		.a(_0215_),
		.b(new_net_154),
		.c(new_net_153)
	);

	spl2 _0212__v_fanout (
		.a(_0212_),
		.b(new_net_47),
		.c(new_net_46)
	);

	spl2 _0299__v_fanout (
		.a(_0299_),
		.b(new_net_461),
		.c(new_net_460)
	);

	bfr new_net_1121_bfr_after (
		.din(_0451_),
		.dout(new_net_1121)
	);

	bfr new_net_1122_bfr_after (
		.din(new_net_1121),
		.dout(new_net_1122)
	);

	bfr new_net_1123_bfr_after (
		.din(new_net_1122),
		.dout(new_net_1123)
	);

	bfr new_net_1124_bfr_after (
		.din(new_net_1123),
		.dout(new_net_1124)
	);

	bfr new_net_1125_bfr_after (
		.din(new_net_1124),
		.dout(new_net_1125)
	);

	spl2 _0451__v_fanout (
		.a(new_net_1125),
		.b(new_net_276),
		.c(new_net_275)
	);

	bfr new_net_1126_bfr_before (
		.din(new_net_1126),
		.dout(G2583)
	);

	bfr new_net_1127_bfr_before (
		.din(new_net_1127),
		.dout(new_net_1126)
	);

	bfr new_net_1128_bfr_before (
		.din(new_net_1128),
		.dout(new_net_1127)
	);

	bfr new_net_1129_bfr_before (
		.din(new_net_1129),
		.dout(new_net_1128)
	);

	bfr new_net_1130_bfr_before (
		.din(new_net_1130),
		.dout(new_net_1129)
	);

	bfr new_net_1131_bfr_before (
		.din(new_net_1131),
		.dout(new_net_1130)
	);

	bfr new_net_1132_bfr_before (
		.din(new_net_1132),
		.dout(new_net_1131)
	);

	bfr new_net_1133_bfr_before (
		.din(new_net_1133),
		.dout(new_net_1132)
	);

	bfr new_net_1134_bfr_before (
		.din(new_net_1134),
		.dout(new_net_1133)
	);

	bfr new_net_1135_bfr_before (
		.din(new_net_1135),
		.dout(new_net_1134)
	);

	bfr new_net_1136_bfr_before (
		.din(new_net_1136),
		.dout(new_net_1135)
	);

	bfr new_net_1137_bfr_before (
		.din(new_net_1137),
		.dout(new_net_1136)
	);

	bfr new_net_1138_bfr_before (
		.din(new_net_1138),
		.dout(new_net_1137)
	);

	bfr new_net_1139_bfr_before (
		.din(new_net_1139),
		.dout(new_net_1138)
	);

	bfr new_net_1140_bfr_before (
		.din(new_net_1140),
		.dout(new_net_1139)
	);

	bfr new_net_1141_bfr_before (
		.din(new_net_1141),
		.dout(new_net_1140)
	);

	spl2 new_net_13_v_fanout (
		.a(new_net_13),
		.b(new_net_150),
		.c(new_net_1141)
	);

	spl4L new_net_746_v_fanout (
		.a(new_net_746),
		.b(new_net_317),
		.c(new_net_319),
		.d(new_net_314),
		.e(new_net_318)
	);

	spl3L new_net_742_v_fanout (
		.a(new_net_742),
		.b(new_net_453),
		.c(new_net_454),
		.d(new_net_455)
	);

	bfr new_net_1142_bfr_after (
		.din(_0399_),
		.dout(new_net_1142)
	);

	spl2 _0399__v_fanout (
		.a(new_net_1142),
		.b(new_net_610),
		.c(new_net_609)
	);

	spl2 new_net_741_v_fanout (
		.a(new_net_741),
		.b(new_net_457),
		.c(new_net_456)
	);

	spl2 new_net_743_v_fanout (
		.a(new_net_743),
		.b(new_net_362),
		.c(new_net_361)
	);

	spl2 new_net_745_v_fanout (
		.a(new_net_745),
		.b(new_net_316),
		.c(new_net_315)
	);

	spl2 _0315__v_fanout (
		.a(_0315_),
		.b(new_net_612),
		.c(new_net_611)
	);

	spl2 _0366__v_fanout (
		.a(_0366_),
		.b(new_net_252),
		.c(new_net_251)
	);

	bfr new_net_1143_bfr_after (
		.din(_0443_),
		.dout(new_net_1143)
	);

	bfr new_net_1144_bfr_after (
		.din(new_net_1143),
		.dout(new_net_1144)
	);

	bfr new_net_1145_bfr_after (
		.din(new_net_1144),
		.dout(new_net_1145)
	);

	bfr new_net_1146_bfr_after (
		.din(new_net_1145),
		.dout(new_net_1146)
	);

	bfr new_net_1147_bfr_after (
		.din(new_net_1146),
		.dout(new_net_1147)
	);

	spl2 _0443__v_fanout (
		.a(new_net_1147),
		.b(new_net_62),
		.c(new_net_61)
	);

	spl3L new_net_744_v_fanout (
		.a(new_net_744),
		.b(new_net_360),
		.c(new_net_358),
		.d(new_net_359)
	);

	spl2 _0345__v_fanout (
		.a(_0345_),
		.b(new_net_250),
		.c(new_net_249)
	);

	bfr new_net_1148_bfr_before (
		.din(new_net_1148),
		.dout(new_net_440)
	);

	spl3L new_net_659_v_fanout (
		.a(new_net_659),
		.b(new_net_441),
		.c(new_net_437),
		.d(new_net_1148)
	);

	spl2 _0390__v_fanout (
		.a(_0390_),
		.b(new_net_323),
		.c(new_net_322)
	);

	spl2 new_net_690_v_fanout (
		.a(new_net_690),
		.b(new_net_194),
		.c(new_net_197)
	);

	spl2 _0415__v_fanout (
		.a(_0415_),
		.b(new_net_742),
		.c(new_net_741)
	);

	spl2 new_net_681_v_fanout (
		.a(new_net_681),
		.b(new_net_354),
		.c(new_net_353)
	);

	bfr new_net_1149_bfr_before (
		.din(new_net_1149),
		.dout(new_net_283)
	);

	spl3L new_net_679_v_fanout (
		.a(new_net_679),
		.b(new_net_1149),
		.c(new_net_280),
		.d(new_net_282)
	);

	spl2 _0412__v_fanout (
		.a(_0412_),
		.b(new_net_744),
		.c(new_net_743)
	);

	bfr new_net_1150_bfr_after (
		.din(_0203_),
		.dout(new_net_1150)
	);

	bfr new_net_1151_bfr_after (
		.din(new_net_1150),
		.dout(new_net_1151)
	);

	bfr new_net_1152_bfr_after (
		.din(new_net_1151),
		.dout(new_net_1152)
	);

	spl2 _0203__v_fanout (
		.a(new_net_1152),
		.b(new_net_388),
		.c(new_net_387)
	);

	spl2 new_net_687_v_fanout (
		.a(new_net_687),
		.b(new_net_76),
		.c(new_net_74)
	);

	spl2 _0465__v_fanout (
		.a(_0465_),
		.b(new_net_745),
		.c(new_net_746)
	);

	spl2 _0285__v_fanout (
		.a(_0285_),
		.b(new_net_272),
		.c(new_net_271)
	);

	spl2 new_net_658_v_fanout (
		.a(new_net_658),
		.b(new_net_166),
		.c(new_net_167)
	);

	bfr new_net_1153_bfr_before (
		.din(new_net_1153),
		.dout(G2557)
	);

	bfr new_net_1154_bfr_before (
		.din(new_net_1154),
		.dout(new_net_1153)
	);

	bfr new_net_1155_bfr_before (
		.din(new_net_1155),
		.dout(new_net_1154)
	);

	bfr new_net_1156_bfr_before (
		.din(new_net_1156),
		.dout(new_net_1155)
	);

	bfr new_net_1157_bfr_before (
		.din(new_net_1157),
		.dout(new_net_1156)
	);

	bfr new_net_1158_bfr_before (
		.din(new_net_1158),
		.dout(new_net_1157)
	);

	bfr new_net_1159_bfr_before (
		.din(new_net_1159),
		.dout(new_net_1158)
	);

	bfr new_net_1160_bfr_before (
		.din(new_net_1160),
		.dout(new_net_1159)
	);

	bfr new_net_1161_bfr_before (
		.din(new_net_1161),
		.dout(new_net_1160)
	);

	bfr new_net_1162_bfr_before (
		.din(new_net_1162),
		.dout(new_net_1161)
	);

	bfr new_net_1163_bfr_before (
		.din(new_net_1163),
		.dout(new_net_1162)
	);

	bfr new_net_1164_bfr_before (
		.din(new_net_1164),
		.dout(new_net_1163)
	);

	bfr new_net_1165_bfr_before (
		.din(new_net_1165),
		.dout(new_net_1164)
	);

	bfr new_net_1166_bfr_before (
		.din(new_net_1166),
		.dout(new_net_1165)
	);

	bfr new_net_1167_bfr_before (
		.din(new_net_1167),
		.dout(new_net_1166)
	);

	bfr new_net_1168_bfr_before (
		.din(new_net_1168),
		.dout(new_net_1167)
	);

	bfr new_net_1169_bfr_before (
		.din(new_net_1169),
		.dout(new_net_1168)
	);

	spl3L new_net_718_v_fanout (
		.a(new_net_718),
		.b(new_net_267),
		.c(new_net_1169),
		.d(new_net_270)
	);

	spl2 _0153__v_fanout (
		.a(_0153_),
		.b(new_net_101),
		.c(new_net_100)
	);

	spl2 _0173__v_fanout (
		.a(_0173_),
		.b(new_net_113),
		.c(new_net_112)
	);

	spl2 new_net_684_v_fanout (
		.a(new_net_684),
		.b(new_net_215),
		.c(new_net_217)
	);

	bfr new_net_1170_bfr_before (
		.din(new_net_1170),
		.dout(G2556)
	);

	bfr new_net_1171_bfr_before (
		.din(new_net_1171),
		.dout(new_net_1170)
	);

	bfr new_net_1172_bfr_before (
		.din(new_net_1172),
		.dout(new_net_1171)
	);

	bfr new_net_1173_bfr_before (
		.din(new_net_1173),
		.dout(new_net_1172)
	);

	bfr new_net_1174_bfr_before (
		.din(new_net_1174),
		.dout(new_net_1173)
	);

	bfr new_net_1175_bfr_before (
		.din(new_net_1175),
		.dout(new_net_1174)
	);

	bfr new_net_1176_bfr_before (
		.din(new_net_1176),
		.dout(new_net_1175)
	);

	bfr new_net_1177_bfr_before (
		.din(new_net_1177),
		.dout(new_net_1176)
	);

	bfr new_net_1178_bfr_before (
		.din(new_net_1178),
		.dout(new_net_1177)
	);

	bfr new_net_1179_bfr_before (
		.din(new_net_1179),
		.dout(new_net_1178)
	);

	bfr new_net_1180_bfr_before (
		.din(new_net_1180),
		.dout(new_net_1179)
	);

	bfr new_net_1181_bfr_before (
		.din(new_net_1181),
		.dout(new_net_1180)
	);

	bfr new_net_1182_bfr_before (
		.din(new_net_1182),
		.dout(new_net_1181)
	);

	bfr new_net_1183_bfr_before (
		.din(new_net_1183),
		.dout(new_net_1182)
	);

	bfr new_net_1184_bfr_before (
		.din(new_net_1184),
		.dout(new_net_1183)
	);

	bfr new_net_1185_bfr_before (
		.din(new_net_1185),
		.dout(new_net_1184)
	);

	bfr new_net_1186_bfr_before (
		.din(new_net_1186),
		.dout(new_net_1185)
	);

	bfr new_net_1187_bfr_before (
		.din(new_net_1187),
		.dout(new_net_1186)
	);

	spl2 new_net_709_v_fanout (
		.a(new_net_709),
		.b(new_net_298),
		.c(new_net_1187)
	);

	bfr new_net_1188_bfr_before (
		.din(new_net_1188),
		.dout(new_net_733)
	);

	bfr new_net_1189_bfr_before (
		.din(new_net_1189),
		.dout(new_net_1188)
	);

	bfr new_net_1190_bfr_before (
		.din(new_net_1190),
		.dout(new_net_1189)
	);

	bfr new_net_1191_bfr_before (
		.din(new_net_1191),
		.dout(new_net_1190)
	);

	bfr new_net_1192_bfr_before (
		.din(new_net_1192),
		.dout(new_net_1191)
	);

	bfr new_net_1193_bfr_before (
		.din(new_net_1193),
		.dout(new_net_1192)
	);

	bfr new_net_1194_bfr_before (
		.din(new_net_1194),
		.dout(new_net_1193)
	);

	bfr new_net_1195_bfr_before (
		.din(new_net_1195),
		.dout(new_net_1194)
	);

	bfr new_net_1196_bfr_before (
		.din(new_net_1196),
		.dout(new_net_1195)
	);

	bfr new_net_1197_bfr_before (
		.din(new_net_1197),
		.dout(new_net_1196)
	);

	bfr new_net_1198_bfr_before (
		.din(new_net_1198),
		.dout(new_net_1197)
	);

	bfr new_net_1199_bfr_before (
		.din(new_net_1199),
		.dout(new_net_1198)
	);

	bfr new_net_1200_bfr_before (
		.din(new_net_1200),
		.dout(new_net_1199)
	);

	bfr new_net_1201_bfr_before (
		.din(new_net_1201),
		.dout(new_net_1200)
	);

	bfr new_net_1202_bfr_before (
		.din(new_net_1202),
		.dout(new_net_1201)
	);

	bfr new_net_1203_bfr_before (
		.din(new_net_1203),
		.dout(new_net_1202)
	);

	bfr new_net_1204_bfr_before (
		.din(new_net_1204),
		.dout(new_net_1203)
	);

	spl4L new_net_735_v_fanout (
		.a(new_net_735),
		.b(new_net_601),
		.c(new_net_606),
		.d(new_net_1204),
		.e(new_net_605)
	);

	spl2 new_net_685_v_fanout (
		.a(new_net_685),
		.b(new_net_130),
		.c(new_net_127)
	);

	spl2 new_net_734_v_fanout (
		.a(new_net_734),
		.b(new_net_602),
		.c(new_net_600)
	);

	spl2 new_net_731_v_fanout (
		.a(new_net_731),
		.b(new_net_173),
		.c(new_net_169)
	);

	bfr new_net_1205_bfr_after (
		.din(_0473_),
		.dout(new_net_1205)
	);

	bfr new_net_1206_bfr_before (
		.din(new_net_1206),
		.dout(new_net_294)
	);

	bfr new_net_1207_bfr_before (
		.din(new_net_1207),
		.dout(new_net_1206)
	);

	bfr new_net_1208_bfr_before (
		.din(new_net_1208),
		.dout(new_net_1207)
	);

	spl2 _0473__v_fanout (
		.a(new_net_1205),
		.b(new_net_1208),
		.c(new_net_293)
	);

	bfr new_net_1209_bfr_before (
		.din(new_net_1209),
		.dout(new_net_216)
	);

	spl2 new_net_683_v_fanout (
		.a(new_net_683),
		.b(new_net_1209),
		.c(new_net_684)
	);

	bfr new_net_1210_bfr_before (
		.din(new_net_1210),
		.dout(new_net_81)
	);

	bfr new_net_1211_bfr_before (
		.din(new_net_1211),
		.dout(new_net_1210)
	);

	bfr new_net_1212_bfr_before (
		.din(new_net_1212),
		.dout(new_net_1211)
	);

	bfr new_net_1213_bfr_before (
		.din(new_net_1213),
		.dout(new_net_1212)
	);

	spl4L new_net_740_v_fanout (
		.a(new_net_740),
		.b(new_net_1213),
		.c(new_net_82),
		.d(new_net_80),
		.e(new_net_77)
	);

	bfr new_net_1214_bfr_before (
		.din(new_net_1214),
		.dout(new_net_724)
	);

	bfr new_net_1215_bfr_before (
		.din(new_net_1215),
		.dout(new_net_1214)
	);

	bfr new_net_1216_bfr_before (
		.din(new_net_1216),
		.dout(new_net_1215)
	);

	bfr new_net_1217_bfr_before (
		.din(new_net_1217),
		.dout(new_net_1216)
	);

	bfr new_net_1218_bfr_before (
		.din(new_net_1218),
		.dout(new_net_1217)
	);

	bfr new_net_1219_bfr_before (
		.din(new_net_1219),
		.dout(new_net_1218)
	);

	bfr new_net_1220_bfr_before (
		.din(new_net_1220),
		.dout(new_net_1219)
	);

	bfr new_net_1221_bfr_before (
		.din(new_net_1221),
		.dout(new_net_1220)
	);

	bfr new_net_1222_bfr_before (
		.din(new_net_1222),
		.dout(new_net_1221)
	);

	bfr new_net_1223_bfr_before (
		.din(new_net_1223),
		.dout(new_net_1222)
	);

	bfr new_net_1224_bfr_before (
		.din(new_net_1224),
		.dout(new_net_1223)
	);

	bfr new_net_1225_bfr_before (
		.din(new_net_1225),
		.dout(new_net_1224)
	);

	bfr new_net_1226_bfr_before (
		.din(new_net_1226),
		.dout(new_net_1225)
	);

	bfr new_net_1227_bfr_before (
		.din(new_net_1227),
		.dout(new_net_1226)
	);

	bfr new_net_1228_bfr_before (
		.din(new_net_1228),
		.dout(new_net_1227)
	);

	bfr new_net_1229_bfr_before (
		.din(new_net_1229),
		.dout(new_net_1228)
	);

	bfr new_net_1230_bfr_before (
		.din(new_net_1230),
		.dout(new_net_1229)
	);

	spl2 new_net_725_v_fanout (
		.a(new_net_725),
		.b(new_net_1230),
		.c(new_net_189)
	);

	spl2 _0303__v_fanout (
		.a(_0303_),
		.b(new_net_248),
		.c(new_net_247)
	);

	bfr new_net_1231_bfr_before (
		.din(new_net_1231),
		.dout(new_net_721)
	);

	bfr new_net_1232_bfr_before (
		.din(new_net_1232),
		.dout(new_net_1231)
	);

	bfr new_net_1233_bfr_before (
		.din(new_net_1233),
		.dout(new_net_1232)
	);

	bfr new_net_1234_bfr_before (
		.din(new_net_1234),
		.dout(new_net_1233)
	);

	spl4L new_net_723_v_fanout (
		.a(new_net_723),
		.b(new_net_1234),
		.c(new_net_235),
		.d(new_net_240),
		.e(new_net_239)
	);

	bfr new_net_1235_bfr_before (
		.din(new_net_1235),
		.dout(new_net_164)
	);

	spl2 new_net_657_v_fanout (
		.a(new_net_657),
		.b(new_net_658),
		.c(new_net_1235)
	);

	spl2 _0324__v_fanout (
		.a(_0324_),
		.b(new_net_64),
		.c(new_net_63)
	);

	bfr new_net_1236_bfr_before (
		.din(new_net_1236),
		.dout(new_net_728)
	);

	bfr new_net_1237_bfr_before (
		.din(new_net_1237),
		.dout(new_net_1236)
	);

	bfr new_net_1238_bfr_before (
		.din(new_net_1238),
		.dout(new_net_1237)
	);

	bfr new_net_1239_bfr_before (
		.din(new_net_1239),
		.dout(new_net_1238)
	);

	spl3L new_net_727_v_fanout (
		.a(new_net_727),
		.b(new_net_595),
		.c(new_net_592),
		.d(new_net_1239)
	);

	spl4L new_net_722_v_fanout (
		.a(new_net_722),
		.b(new_net_236),
		.c(new_net_237),
		.d(new_net_238),
		.e(new_net_234)
	);

	bfr new_net_1240_bfr_before (
		.din(new_net_1240),
		.dout(new_net_737)
	);

	bfr new_net_1241_bfr_before (
		.din(new_net_1241),
		.dout(new_net_1240)
	);

	bfr new_net_1242_bfr_before (
		.din(new_net_1242),
		.dout(new_net_1241)
	);

	bfr new_net_1243_bfr_before (
		.din(new_net_1243),
		.dout(new_net_1242)
	);

	spl3L new_net_736_v_fanout (
		.a(new_net_736),
		.b(new_net_432),
		.c(new_net_429),
		.d(new_net_1243)
	);

	spl2 _0333__v_fanout (
		.a(_0333_),
		.b(new_net_152),
		.c(new_net_151)
	);

	bfr new_net_1244_bfr_before (
		.din(new_net_1244),
		.dout(G2572)
	);

	bfr new_net_1245_bfr_before (
		.din(new_net_1245),
		.dout(new_net_1244)
	);

	bfr new_net_1246_bfr_before (
		.din(new_net_1246),
		.dout(new_net_1245)
	);

	bfr new_net_1247_bfr_before (
		.din(new_net_1247),
		.dout(new_net_1246)
	);

	bfr new_net_1248_bfr_before (
		.din(new_net_1248),
		.dout(new_net_1247)
	);

	bfr new_net_1249_bfr_before (
		.din(new_net_1249),
		.dout(new_net_1248)
	);

	bfr new_net_1250_bfr_before (
		.din(new_net_1250),
		.dout(new_net_1249)
	);

	bfr new_net_1251_bfr_before (
		.din(new_net_1251),
		.dout(new_net_1250)
	);

	bfr new_net_1252_bfr_before (
		.din(new_net_1252),
		.dout(new_net_1251)
	);

	bfr new_net_1253_bfr_before (
		.din(new_net_1253),
		.dout(new_net_1252)
	);

	bfr new_net_1254_bfr_before (
		.din(new_net_1254),
		.dout(new_net_1253)
	);

	bfr new_net_1255_bfr_before (
		.din(new_net_1255),
		.dout(new_net_1254)
	);

	bfr new_net_1256_bfr_before (
		.din(new_net_1256),
		.dout(new_net_1255)
	);

	bfr new_net_1257_bfr_before (
		.din(new_net_1257),
		.dout(new_net_1256)
	);

	bfr new_net_1258_bfr_before (
		.din(new_net_1258),
		.dout(new_net_1257)
	);

	bfr new_net_1259_bfr_before (
		.din(new_net_1259),
		.dout(new_net_1258)
	);

	bfr new_net_1260_bfr_before (
		.din(new_net_1260),
		.dout(new_net_1259)
	);

	bfr new_net_1261_bfr_before (
		.din(new_net_1261),
		.dout(new_net_1260)
	);

	spl4L new_net_732_v_fanout (
		.a(new_net_732),
		.b(new_net_172),
		.c(new_net_168),
		.d(new_net_1261),
		.e(new_net_171)
	);

	spl2 _0353__v_fanout (
		.a(_0353_),
		.b(new_net_608),
		.c(new_net_607)
	);

	spl2 new_net_689_v_fanout (
		.a(new_net_689),
		.b(new_net_690),
		.c(new_net_196)
	);

	bfr new_net_1262_bfr_before (
		.din(new_net_1262),
		.dout(new_net_303)
	);

	bfr new_net_1263_bfr_before (
		.din(new_net_1263),
		.dout(new_net_1262)
	);

	bfr new_net_1264_bfr_before (
		.din(new_net_1264),
		.dout(new_net_1263)
	);

	spl3L new_net_669_v_fanout (
		.a(new_net_669),
		.b(new_net_1264),
		.c(new_net_301),
		.d(new_net_304)
	);

	spl2 new_net_739_v_fanout (
		.a(new_net_739),
		.b(new_net_78),
		.c(new_net_79)
	);

	spl3L new_net_726_v_fanout (
		.a(new_net_726),
		.b(new_net_188),
		.c(new_net_191),
		.d(new_net_192)
	);

	spl2 _0308__v_fanout (
		.a(_0308_),
		.b(new_net_564),
		.c(new_net_563)
	);

	spl2 new_net_686_v_fanout (
		.a(new_net_686),
		.b(new_net_687),
		.c(new_net_73)
	);

	bfr new_net_1265_bfr_before (
		.din(new_net_1265),
		.dout(G2582)
	);

	bfr new_net_1266_bfr_before (
		.din(new_net_1266),
		.dout(new_net_1265)
	);

	bfr new_net_1267_bfr_before (
		.din(new_net_1267),
		.dout(new_net_1266)
	);

	bfr new_net_1268_bfr_before (
		.din(new_net_1268),
		.dout(new_net_1267)
	);

	bfr new_net_1269_bfr_before (
		.din(new_net_1269),
		.dout(new_net_1268)
	);

	bfr new_net_1270_bfr_before (
		.din(new_net_1270),
		.dout(new_net_1269)
	);

	bfr new_net_1271_bfr_before (
		.din(new_net_1271),
		.dout(new_net_1270)
	);

	bfr new_net_1272_bfr_before (
		.din(new_net_1272),
		.dout(new_net_1271)
	);

	bfr new_net_1273_bfr_before (
		.din(new_net_1273),
		.dout(new_net_1272)
	);

	bfr new_net_1274_bfr_before (
		.din(new_net_1274),
		.dout(new_net_1273)
	);

	bfr new_net_1275_bfr_before (
		.din(new_net_1275),
		.dout(new_net_1274)
	);

	bfr new_net_1276_bfr_before (
		.din(new_net_1276),
		.dout(new_net_1275)
	);

	bfr new_net_1277_bfr_before (
		.din(new_net_1277),
		.dout(new_net_1276)
	);

	bfr new_net_1278_bfr_before (
		.din(new_net_1278),
		.dout(new_net_1277)
	);

	bfr new_net_1279_bfr_before (
		.din(new_net_1279),
		.dout(new_net_1278)
	);

	bfr new_net_1280_bfr_before (
		.din(new_net_1280),
		.dout(new_net_1279)
	);

	bfr new_net_1281_bfr_before (
		.din(new_net_1281),
		.dout(new_net_1280)
	);

	bfr new_net_1282_bfr_before (
		.din(new_net_1282),
		.dout(new_net_1281)
	);

	spl2 new_net_12_v_fanout (
		.a(new_net_12),
		.b(new_net_321),
		.c(new_net_1282)
	);

	bfr new_net_1283_bfr_after (
		.din(_0190_),
		.dout(new_net_1283)
	);

	spl2 _0190__v_fanout (
		.a(new_net_1283),
		.b(new_net_30),
		.c(new_net_29)
	);

	spl2 _0085__v_fanout (
		.a(_0085_),
		.b(new_net_261),
		.c(new_net_260)
	);

	spl2 _0248__v_fanout (
		.a(_0248_),
		.b(new_net_722),
		.c(new_net_723)
	);

	bfr new_net_1284_bfr_before (
		.din(new_net_1284),
		.dout(new_net_720)
	);

	bfr new_net_1285_bfr_before (
		.din(new_net_1285),
		.dout(new_net_1284)
	);

	bfr new_net_1286_bfr_before (
		.din(new_net_1286),
		.dout(new_net_1285)
	);

	spl3L new_net_719_v_fanout (
		.a(new_net_719),
		.b(new_net_1286),
		.c(new_net_287),
		.d(new_net_286)
	);

	spl2 new_net_5_v_fanout (
		.a(new_net_5),
		.b(new_net_725),
		.c(new_net_726)
	);

	spl3L new_net_9_v_fanout (
		.a(new_net_9),
		.b(new_net_597),
		.c(new_net_596),
		.d(new_net_727)
	);

	bfr new_net_1287_bfr_before (
		.din(new_net_1287),
		.dout(new_net_730)
	);

	bfr new_net_1288_bfr_before (
		.din(new_net_1288),
		.dout(new_net_1287)
	);

	bfr new_net_1289_bfr_before (
		.din(new_net_1289),
		.dout(new_net_1288)
	);

	bfr new_net_1290_bfr_before (
		.din(new_net_1290),
		.dout(new_net_1289)
	);

	bfr new_net_1291_bfr_before (
		.din(new_net_1291),
		.dout(new_net_309)
	);

	bfr new_net_1292_bfr_before (
		.din(new_net_1292),
		.dout(new_net_307)
	);

	spl4L new_net_4_v_fanout (
		.a(new_net_4),
		.b(new_net_305),
		.c(new_net_1290),
		.d(new_net_1291),
		.e(new_net_1292)
	);

	spl3L _0410__v_fanout (
		.a(_0410_),
		.b(new_net_576),
		.c(new_net_574),
		.d(new_net_575)
	);

	bfr new_net_1293_bfr_before (
		.din(new_net_1293),
		.dout(new_net_529)
	);

	bfr new_net_1294_bfr_before (
		.din(new_net_1294),
		.dout(new_net_532)
	);

	spl4L _0226__v_fanout (
		.a(_0226_),
		.b(new_net_530),
		.c(new_net_1293),
		.d(new_net_1294),
		.e(new_net_531)
	);

	bfr new_net_1295_bfr_before (
		.din(new_net_1295),
		.dout(new_net_521)
	);

	bfr new_net_1296_bfr_before (
		.din(new_net_1296),
		.dout(new_net_1295)
	);

	spl3L new_net_678_v_fanout (
		.a(new_net_678),
		.b(new_net_1296),
		.c(new_net_523),
		.d(new_net_522)
	);

	bfr new_net_1297_bfr_before (
		.din(new_net_1297),
		.dout(new_net_583)
	);

	bfr new_net_1298_bfr_before (
		.din(new_net_1298),
		.dout(new_net_1297)
	);

	spl3L new_net_688_v_fanout (
		.a(new_net_688),
		.b(new_net_582),
		.c(new_net_581),
		.d(new_net_1298)
	);

	spl2 new_net_3_v_fanout (
		.a(new_net_3),
		.b(new_net_731),
		.c(new_net_732)
	);

	spl2 new_net_8_v_fanout (
		.a(new_net_8),
		.b(new_net_734),
		.c(new_net_735)
	);

	bfr new_net_1299_bfr_before (
		.din(new_net_1299),
		.dout(new_net_624)
	);

	bfr new_net_1300_bfr_before (
		.din(new_net_1300),
		.dout(new_net_1299)
	);

	bfr new_net_1301_bfr_before (
		.din(new_net_1301),
		.dout(new_net_1300)
	);

	bfr new_net_1302_bfr_before (
		.din(new_net_1302),
		.dout(new_net_1301)
	);

	spl3L new_net_656_v_fanout (
		.a(new_net_656),
		.b(new_net_1302),
		.c(new_net_625),
		.d(new_net_626)
	);

	bfr new_net_1303_bfr_before (
		.din(new_net_1303),
		.dout(new_net_26)
	);

	bfr new_net_1304_bfr_before (
		.din(new_net_1304),
		.dout(new_net_1303)
	);

	bfr new_net_1305_bfr_before (
		.din(new_net_1305),
		.dout(new_net_1304)
	);

	bfr new_net_1306_bfr_before (
		.din(new_net_1306),
		.dout(new_net_1305)
	);

	spl3L new_net_660_v_fanout (
		.a(new_net_660),
		.b(new_net_1306),
		.c(new_net_25),
		.d(new_net_27)
	);

	spl3L new_net_7_v_fanout (
		.a(new_net_7),
		.b(new_net_434),
		.c(new_net_433),
		.d(new_net_736)
	);

	bfr new_net_1307_bfr_before (
		.din(new_net_1307),
		.dout(new_net_420)
	);

	bfr new_net_1308_bfr_before (
		.din(new_net_1308),
		.dout(new_net_1307)
	);

	spl3L new_net_638_v_fanout (
		.a(new_net_638),
		.b(new_net_418),
		.c(new_net_421),
		.d(new_net_1308)
	);

	spl3L _0411__v_fanout (
		.a(_0411_),
		.b(new_net_220),
		.c(new_net_219),
		.d(new_net_221)
	);

	bfr new_net_1309_bfr_before (
		.din(new_net_1309),
		.dout(new_net_333)
	);

	bfr new_net_1310_bfr_before (
		.din(new_net_1310),
		.dout(new_net_1309)
	);

	spl3L new_net_641_v_fanout (
		.a(new_net_641),
		.b(new_net_334),
		.c(new_net_330),
		.d(new_net_1310)
	);

	spl2 new_net_662_v_fanout (
		.a(new_net_662),
		.b(new_net_384),
		.c(new_net_385)
	);

	bfr new_net_1311_bfr_before (
		.din(new_net_1311),
		.dout(new_net_486)
	);

	spl3L new_net_640_v_fanout (
		.a(new_net_640),
		.b(new_net_482),
		.c(new_net_487),
		.d(new_net_1311)
	);

	spl2 _0234__v_fanout (
		.a(_0234_),
		.b(new_net_740),
		.c(new_net_739)
	);

	spl2 _0131__v_fanout (
		.a(_0131_),
		.b(new_net_374),
		.c(new_net_373)
	);

	spl3L new_net_717_v_fanout (
		.a(new_net_717),
		.b(new_net_87),
		.c(new_net_83),
		.d(new_net_84)
	);

	spl2 new_net_714_v_fanout (
		.a(new_net_714),
		.b(new_net_449),
		.c(new_net_448)
	);

	bfr new_net_1312_bfr_before (
		.din(new_net_1312),
		.dout(new_net_613)
	);

	bfr new_net_1313_bfr_before (
		.din(new_net_1313),
		.dout(new_net_616)
	);

	bfr new_net_1314_bfr_before (
		.din(new_net_1314),
		.dout(new_net_1313)
	);

	bfr new_net_1315_bfr_before (
		.din(new_net_1315),
		.dout(new_net_1314)
	);

	bfr new_net_1316_bfr_before (
		.din(new_net_1316),
		.dout(new_net_1315)
	);

	bfr new_net_1317_bfr_before (
		.din(new_net_1317),
		.dout(new_net_1316)
	);

	bfr new_net_1318_bfr_before (
		.din(new_net_1318),
		.dout(new_net_1317)
	);

	bfr new_net_1319_bfr_before (
		.din(new_net_1319),
		.dout(new_net_1318)
	);

	spl3L new_net_682_v_fanout (
		.a(new_net_682),
		.b(new_net_1319),
		.c(new_net_1312),
		.d(new_net_614)
	);

	spl2 _0271__v_fanout (
		.a(_0271_),
		.b(new_net_500),
		.c(new_net_499)
	);

	spl2 new_net_712_v_fanout (
		.a(new_net_712),
		.b(new_net_56),
		.c(new_net_58)
	);

	bfr new_net_1320_bfr_before (
		.din(new_net_1320),
		.dout(new_net_719)
	);

	spl2 new_net_6_v_fanout (
		.a(new_net_6),
		.b(new_net_1320),
		.c(new_net_285)
	);

	bfr new_net_1321_bfr_before (
		.din(new_net_1321),
		.dout(G2559)
	);

	bfr new_net_1322_bfr_before (
		.din(new_net_1322),
		.dout(new_net_1321)
	);

	bfr new_net_1323_bfr_before (
		.din(new_net_1323),
		.dout(new_net_1322)
	);

	bfr new_net_1324_bfr_before (
		.din(new_net_1324),
		.dout(new_net_1323)
	);

	bfr new_net_1325_bfr_before (
		.din(new_net_1325),
		.dout(new_net_1324)
	);

	bfr new_net_1326_bfr_before (
		.din(new_net_1326),
		.dout(new_net_1325)
	);

	bfr new_net_1327_bfr_before (
		.din(new_net_1327),
		.dout(new_net_1326)
	);

	bfr new_net_1328_bfr_before (
		.din(new_net_1328),
		.dout(new_net_1327)
	);

	bfr new_net_1329_bfr_before (
		.din(new_net_1329),
		.dout(new_net_1328)
	);

	bfr new_net_1330_bfr_before (
		.din(new_net_1330),
		.dout(new_net_1329)
	);

	bfr new_net_1331_bfr_before (
		.din(new_net_1331),
		.dout(new_net_1330)
	);

	bfr new_net_1332_bfr_before (
		.din(new_net_1332),
		.dout(new_net_1331)
	);

	bfr new_net_1333_bfr_before (
		.din(new_net_1333),
		.dout(new_net_1332)
	);

	bfr new_net_1334_bfr_before (
		.din(new_net_1334),
		.dout(new_net_1333)
	);

	bfr new_net_1335_bfr_before (
		.din(new_net_1335),
		.dout(new_net_1334)
	);

	bfr new_net_1336_bfr_before (
		.din(new_net_1336),
		.dout(new_net_1335)
	);

	bfr new_net_1337_bfr_before (
		.din(new_net_1337),
		.dout(new_net_1336)
	);

	bfr new_net_1338_bfr_before (
		.din(new_net_1338),
		.dout(new_net_1337)
	);

	bfr new_net_1339_bfr_before (
		.din(new_net_1339),
		.dout(new_net_1338)
	);

	bfr new_net_1340_bfr_before (
		.din(new_net_1340),
		.dout(new_net_1339)
	);

	spl3L new_net_715_v_fanout (
		.a(new_net_715),
		.b(new_net_1340),
		.c(new_net_255),
		.d(new_net_258)
	);

	bfr new_net_1341_bfr_before (
		.din(new_net_1341),
		.dout(new_net_364)
	);

	bfr new_net_1342_bfr_before (
		.din(new_net_1342),
		.dout(new_net_365)
	);

	spl4L new_net_671_v_fanout (
		.a(new_net_671),
		.b(new_net_368),
		.c(new_net_1341),
		.d(new_net_1342),
		.e(new_net_366)
	);

	bfr new_net_1343_bfr_before (
		.din(new_net_1343),
		.dout(new_net_681)
	);

	bfr new_net_1344_bfr_before (
		.din(new_net_1344),
		.dout(new_net_1343)
	);

	spl3L new_net_680_v_fanout (
		.a(new_net_680),
		.b(new_net_356),
		.c(new_net_1344),
		.d(new_net_357)
	);

	spl2 new_net_710_v_fanout (
		.a(new_net_710),
		.b(new_net_428),
		.c(new_net_427)
	);

	spl4L new_net_665_v_fanout (
		.a(new_net_665),
		.b(new_net_516),
		.c(new_net_503),
		.d(new_net_504),
		.e(new_net_517)
	);

	spl2 new_net_716_v_fanout (
		.a(new_net_716),
		.b(new_net_85),
		.c(new_net_86)
	);

	spl3L new_net_711_v_fanout (
		.a(new_net_711),
		.b(new_net_425),
		.c(new_net_424),
		.d(new_net_426)
	);

	spl3L new_net_713_v_fanout (
		.a(new_net_713),
		.b(new_net_54),
		.c(new_net_55),
		.d(new_net_57)
	);

	bfr new_net_1345_bfr_before (
		.din(new_net_1345),
		.dout(new_net_514)
	);

	spl4L new_net_664_v_fanout (
		.a(new_net_664),
		.b(new_net_512),
		.c(new_net_505),
		.d(new_net_1345),
		.e(new_net_515)
	);

	bfr new_net_1346_bfr_before (
		.din(new_net_1346),
		.dout(new_net_370)
	);

	bfr new_net_1347_bfr_before (
		.din(new_net_1347),
		.dout(new_net_1346)
	);

	bfr new_net_1348_bfr_before (
		.din(new_net_1348),
		.dout(new_net_1347)
	);

	bfr new_net_1349_bfr_before (
		.din(new_net_1349),
		.dout(new_net_1348)
	);

	bfr new_net_1350_bfr_before (
		.din(new_net_1350),
		.dout(new_net_1349)
	);

	bfr new_net_1351_bfr_before (
		.din(new_net_1351),
		.dout(new_net_1350)
	);

	bfr new_net_1352_bfr_before (
		.din(new_net_1352),
		.dout(new_net_1351)
	);

	bfr new_net_1353_bfr_before (
		.din(new_net_1353),
		.dout(new_net_1352)
	);

	bfr new_net_1354_bfr_before (
		.din(new_net_1354),
		.dout(new_net_1353)
	);

	bfr new_net_1355_bfr_before (
		.din(new_net_1355),
		.dout(new_net_1354)
	);

	bfr new_net_1356_bfr_before (
		.din(new_net_1356),
		.dout(new_net_1355)
	);

	bfr new_net_1357_bfr_before (
		.din(new_net_1357),
		.dout(new_net_1356)
	);

	bfr new_net_1358_bfr_before (
		.din(new_net_1358),
		.dout(new_net_363)
	);

	spl3L new_net_670_v_fanout (
		.a(new_net_670),
		.b(new_net_1358),
		.c(new_net_1357),
		.d(new_net_367)
	);

	spl2 _0200__v_fanout (
		.a(_0200_),
		.b(new_net_710),
		.c(new_net_711)
	);

	spl2 _0180__v_fanout (
		.a(_0180_),
		.b(new_net_313),
		.c(new_net_312)
	);

	spl2 _0170__v_fanout (
		.a(_0170_),
		.b(new_net_712),
		.c(new_net_713)
	);

	bfr new_net_1359_bfr_before (
		.din(new_net_1359),
		.dout(G2558)
	);

	bfr new_net_1360_bfr_before (
		.din(new_net_1360),
		.dout(new_net_1359)
	);

	bfr new_net_1361_bfr_before (
		.din(new_net_1361),
		.dout(new_net_1360)
	);

	bfr new_net_1362_bfr_before (
		.din(new_net_1362),
		.dout(new_net_1361)
	);

	bfr new_net_1363_bfr_before (
		.din(new_net_1363),
		.dout(new_net_1362)
	);

	bfr new_net_1364_bfr_before (
		.din(new_net_1364),
		.dout(new_net_1363)
	);

	bfr new_net_1365_bfr_before (
		.din(new_net_1365),
		.dout(new_net_1364)
	);

	bfr new_net_1366_bfr_before (
		.din(new_net_1366),
		.dout(new_net_1365)
	);

	bfr new_net_1367_bfr_before (
		.din(new_net_1367),
		.dout(new_net_1366)
	);

	bfr new_net_1368_bfr_before (
		.din(new_net_1368),
		.dout(new_net_1367)
	);

	bfr new_net_1369_bfr_before (
		.din(new_net_1369),
		.dout(new_net_1368)
	);

	bfr new_net_1370_bfr_before (
		.din(new_net_1370),
		.dout(new_net_1369)
	);

	bfr new_net_1371_bfr_before (
		.din(new_net_1371),
		.dout(new_net_1370)
	);

	bfr new_net_1372_bfr_before (
		.din(new_net_1372),
		.dout(new_net_1371)
	);

	bfr new_net_1373_bfr_before (
		.din(new_net_1373),
		.dout(new_net_1372)
	);

	bfr new_net_1374_bfr_before (
		.din(new_net_1374),
		.dout(new_net_1373)
	);

	bfr new_net_1375_bfr_before (
		.din(new_net_1375),
		.dout(new_net_1374)
	);

	bfr new_net_1376_bfr_before (
		.din(new_net_1376),
		.dout(new_net_1375)
	);

	bfr new_net_1377_bfr_before (
		.din(new_net_1377),
		.dout(new_net_1376)
	);

	bfr new_net_1378_bfr_before (
		.din(new_net_1378),
		.dout(new_net_1377)
	);

	bfr new_net_1379_bfr_before (
		.din(new_net_1379),
		.dout(new_net_1378)
	);

	bfr new_net_1380_bfr_before (
		.din(new_net_1380),
		.dout(new_net_467)
	);

	bfr new_net_1381_bfr_before (
		.din(new_net_1381),
		.dout(new_net_465)
	);

	spl4L new_net_0_v_fanout (
		.a(new_net_0),
		.b(new_net_1380),
		.c(new_net_1379),
		.d(new_net_466),
		.e(new_net_1381)
	);

	spl4L _0163__v_fanout (
		.a(_0163_),
		.b(new_net_452),
		.c(new_net_450),
		.d(new_net_451),
		.e(new_net_714)
	);

	spl2 _0105__v_fanout (
		.a(_0105_),
		.b(new_net_97),
		.c(new_net_96)
	);

	bfr new_net_1382_bfr_before (
		.din(new_net_1382),
		.dout(new_net_665)
	);

	spl3L new_net_663_v_fanout (
		.a(new_net_663),
		.b(new_net_513),
		.c(new_net_1382),
		.d(new_net_664)
	);

	spl3L _0187__v_fanout (
		.a(_0187_),
		.b(new_net_561),
		.c(new_net_560),
		.d(new_net_562)
	);

	spl3L new_net_2_v_fanout (
		.a(new_net_2),
		.b(new_net_257),
		.c(new_net_259),
		.d(new_net_715)
	);

	spl2 _0150__v_fanout (
		.a(_0150_),
		.b(new_net_716),
		.c(new_net_717)
	);

	bfr new_net_1383_bfr_before (
		.din(new_net_1383),
		.dout(new_net_718)
	);

	bfr new_net_1384_bfr_before (
		.din(new_net_1384),
		.dout(new_net_1383)
	);

	bfr new_net_1385_bfr_before (
		.din(new_net_1385),
		.dout(new_net_1384)
	);

	spl3L new_net_1_v_fanout (
		.a(new_net_1),
		.b(new_net_268),
		.c(new_net_269),
		.d(new_net_1385)
	);

	spl2 _0079__v_fanout (
		.a(_0079_),
		.b(new_net_459),
		.c(new_net_458)
	);

	bfr new_net_1386_bfr_before (
		.din(new_net_1386),
		.dout(new_net_141)
	);

	bfr new_net_1387_bfr_before (
		.din(new_net_1387),
		.dout(new_net_137)
	);

	spl4L new_net_674_v_fanout (
		.a(new_net_674),
		.b(new_net_1387),
		.c(new_net_1386),
		.d(new_net_133),
		.e(new_net_138)
	);

	bfr new_net_1388_bfr_after (
		.din(_0114_),
		.dout(new_net_1388)
	);

	spl2 _0114__v_fanout (
		.a(new_net_1388),
		.b(new_net_372),
		.c(new_net_371)
	);

	bfr new_net_1389_bfr_before (
		.din(new_net_1389),
		.dout(new_net_139)
	);

	spl4L new_net_673_v_fanout (
		.a(new_net_673),
		.b(new_net_1389),
		.c(new_net_132),
		.d(new_net_140),
		.e(new_net_144)
	);

	bfr new_net_1390_bfr_before (
		.din(new_net_1390),
		.dout(new_net_640)
	);

	bfr new_net_1391_bfr_before (
		.din(new_net_1391),
		.dout(new_net_1390)
	);

	spl3L new_net_639_v_fanout (
		.a(new_net_639),
		.b(new_net_488),
		.c(new_net_1391),
		.d(new_net_484)
	);

	spl2 _0125__v_fanout (
		.a(_0125_),
		.b(new_net_111),
		.c(new_net_110)
	);

	spl2 new_net_650_v_fanout (
		.a(new_net_650),
		.b(new_net_50),
		.c(new_net_49)
	);

	bfr new_net_1392_bfr_after (
		.din(_0140_),
		.dout(new_net_1392)
	);

	bfr new_net_1393_bfr_after (
		.din(new_net_1392),
		.dout(new_net_1393)
	);

	bfr new_net_1394_bfr_after (
		.din(new_net_1393),
		.dout(new_net_1394)
	);

	spl2 _0140__v_fanout (
		.a(new_net_1394),
		.b(new_net_380),
		.c(new_net_379)
	);

	bfr new_net_1395_bfr_after (
		.din(_0094_),
		.dout(new_net_1395)
	);

	bfr new_net_1396_bfr_after (
		.din(new_net_1395),
		.dout(new_net_1396)
	);

	bfr new_net_1397_bfr_after (
		.din(new_net_1396),
		.dout(new_net_1397)
	);

	spl2 _0094__v_fanout (
		.a(new_net_1397),
		.b(new_net_329),
		.c(new_net_328)
	);

	bfr new_net_1398_bfr_before (
		.din(new_net_1398),
		.dout(new_net_638)
	);

	bfr new_net_1399_bfr_before (
		.din(new_net_1399),
		.dout(new_net_1398)
	);

	spl3L new_net_637_v_fanout (
		.a(new_net_637),
		.b(new_net_422),
		.c(new_net_1399),
		.d(new_net_423)
	);

	bfr new_net_1400_bfr_before (
		.din(new_net_1400),
		.dout(new_net_662)
	);

	bfr new_net_1401_bfr_before (
		.din(new_net_1401),
		.dout(new_net_1400)
	);

	spl3L new_net_661_v_fanout (
		.a(new_net_661),
		.b(new_net_1401),
		.c(new_net_383),
		.d(new_net_382)
	);

	bfr new_net_1402_bfr_before (
		.din(new_net_1402),
		.dout(new_net_709)
	);

	bfr new_net_1403_bfr_before (
		.din(new_net_1403),
		.dout(new_net_1402)
	);

	bfr new_net_1404_bfr_before (
		.din(new_net_1404),
		.dout(new_net_1403)
	);

	spl2 new_net_11_v_fanout (
		.a(new_net_11),
		.b(new_net_299),
		.c(new_net_1404)
	);

	spl2 new_net_703_v_fanout (
		.a(new_net_703),
		.b(new_net_209),
		.c(new_net_208)
	);

	spl4L new_net_704_v_fanout (
		.a(new_net_704),
		.b(new_net_201),
		.c(new_net_200),
		.d(new_net_203),
		.e(new_net_204)
	);

	spl4L new_net_707_v_fanout (
		.a(new_net_707),
		.b(new_net_35),
		.c(new_net_33),
		.d(new_net_34),
		.e(new_net_36)
	);

	spl3L new_net_708_v_fanout (
		.a(new_net_708),
		.b(new_net_39),
		.c(new_net_37),
		.d(new_net_38)
	);

	bfr new_net_1405_bfr_after (
		.din(new_net_17),
		.dout(new_net_1405)
	);

	bfr new_net_1406_bfr_after (
		.din(new_net_1405),
		.dout(new_net_1406)
	);

	bfr new_net_1407_bfr_after (
		.din(new_net_1406),
		.dout(new_net_1407)
	);

	bfr new_net_1408_bfr_after (
		.din(new_net_1407),
		.dout(new_net_1408)
	);

	bfr new_net_1409_bfr_after (
		.din(new_net_1408),
		.dout(new_net_1409)
	);

	bfr new_net_1410_bfr_after (
		.din(new_net_1409),
		.dout(new_net_1410)
	);

	bfr new_net_1411_bfr_after (
		.din(new_net_1410),
		.dout(new_net_1411)
	);

	bfr new_net_1412_bfr_after (
		.din(new_net_1411),
		.dout(new_net_1412)
	);

	bfr new_net_1413_bfr_after (
		.din(new_net_1412),
		.dout(new_net_1413)
	);

	bfr new_net_1414_bfr_after (
		.din(new_net_1413),
		.dout(new_net_1414)
	);

	bfr new_net_1415_bfr_after (
		.din(new_net_1414),
		.dout(new_net_1415)
	);

	bfr new_net_1416_bfr_after (
		.din(new_net_1415),
		.dout(new_net_1416)
	);

	bfr new_net_1417_bfr_after (
		.din(new_net_1416),
		.dout(new_net_1417)
	);

	bfr new_net_1418_bfr_after (
		.din(new_net_1417),
		.dout(new_net_1418)
	);

	bfr new_net_1419_bfr_after (
		.din(new_net_1418),
		.dout(new_net_1419)
	);

	bfr new_net_1420_bfr_after (
		.din(new_net_1419),
		.dout(new_net_1420)
	);

	bfr new_net_1421_bfr_after (
		.din(new_net_1420),
		.dout(new_net_1421)
	);

	bfr new_net_1422_bfr_after (
		.din(new_net_1421),
		.dout(new_net_1422)
	);

	bfr new_net_1423_bfr_after (
		.din(new_net_1422),
		.dout(new_net_1423)
	);

	bfr new_net_1424_bfr_after (
		.din(new_net_1423),
		.dout(new_net_1424)
	);

	bfr new_net_1425_bfr_after (
		.din(new_net_1424),
		.dout(new_net_1425)
	);

	bfr new_net_1426_bfr_after (
		.din(new_net_1425),
		.dout(new_net_1426)
	);

	bfr new_net_1427_bfr_after (
		.din(new_net_1426),
		.dout(new_net_1427)
	);

	spl2 new_net_17_v_fanout (
		.a(new_net_1427),
		.b(G2555),
		.c(G2554)
	);

	spl4L new_net_705_v_fanout (
		.a(new_net_705),
		.b(new_net_205),
		.c(new_net_202),
		.d(new_net_207),
		.e(new_net_206)
	);

	spl2 new_net_706_v_fanout (
		.a(new_net_706),
		.b(new_net_41),
		.c(new_net_40)
	);

	spl3L _0028__v_fanout (
		.a(_0028_),
		.b(new_net_704),
		.c(new_net_705),
		.d(new_net_703)
	);

	spl2 _0099__v_fanout (
		.a(_0099_),
		.b(new_net_447),
		.c(new_net_446)
	);

	spl3L _0026__v_fanout (
		.a(_0026_),
		.b(new_net_706),
		.c(new_net_707),
		.d(new_net_708)
	);

	spl2 _0102__v_fanout (
		.a(_0102_),
		.b(new_net_263),
		.c(new_net_262)
	);

	spl3L new_net_693_v_fanout (
		.a(new_net_693),
		.b(new_net_124),
		.c(new_net_120),
		.d(new_net_123)
	);

	spl2 new_net_694_v_fanout (
		.a(new_net_694),
		.b(new_net_635),
		.c(new_net_634)
	);

	spl3L new_net_699_v_fanout (
		.a(new_net_699),
		.b(new_net_179),
		.c(new_net_176),
		.d(new_net_180)
	);

	bfr new_net_1428_bfr_after (
		.din(_0128_),
		.dout(new_net_1428)
	);

	bfr new_net_1429_bfr_after (
		.din(new_net_1428),
		.dout(new_net_1429)
	);

	bfr new_net_1430_bfr_after (
		.din(new_net_1429),
		.dout(new_net_1430)
	);

	spl2 _0128__v_fanout (
		.a(new_net_1430),
		.b(new_net_53),
		.c(new_net_52)
	);

	spl3L new_net_702_v_fanout (
		.a(new_net_702),
		.b(new_net_539),
		.c(new_net_536),
		.d(new_net_540)
	);

	spl2 _0073__v_fanout (
		.a(_0073_),
		.b(new_net_274),
		.c(new_net_273)
	);

	spl2 new_net_651_v_fanout (
		.a(new_net_651),
		.b(new_net_556),
		.c(new_net_557)
	);

	spl2 new_net_691_v_fanout (
		.a(new_net_691),
		.b(new_net_126),
		.c(new_net_125)
	);

	spl2 _0111__v_fanout (
		.a(_0111_),
		.b(new_net_162),
		.c(new_net_161)
	);

	spl4L new_net_653_v_fanout (
		.a(new_net_653),
		.b(new_net_551),
		.c(new_net_548),
		.d(new_net_554),
		.e(new_net_555)
	);

	bfr new_net_1431_bfr_after (
		.din(_0082_),
		.dout(new_net_1431)
	);

	bfr new_net_1432_bfr_after (
		.din(new_net_1431),
		.dout(new_net_1432)
	);

	bfr new_net_1433_bfr_after (
		.din(new_net_1432),
		.dout(new_net_1433)
	);

	spl2 _0082__v_fanout (
		.a(new_net_1433),
		.b(new_net_568),
		.c(new_net_567)
	);

	spl2 _0076__v_fanout (
		.a(_0076_),
		.b(new_net_351),
		.c(new_net_350)
	);

	spl2 _0134__v_fanout (
		.a(_0134_),
		.b(new_net_223),
		.c(new_net_222)
	);

	spl4L new_net_695_v_fanout (
		.a(new_net_695),
		.b(new_net_629),
		.c(new_net_636),
		.d(new_net_628),
		.e(new_net_632)
	);

	spl2 _0108__v_fanout (
		.a(_0108_),
		.b(new_net_109),
		.c(new_net_108)
	);

	spl3L new_net_696_v_fanout (
		.a(new_net_696),
		.b(new_net_633),
		.c(new_net_631),
		.d(new_net_630)
	);

	spl2 _0091__v_fanout (
		.a(_0091_),
		.b(new_net_186),
		.c(new_net_185)
	);

	spl4L new_net_701_v_fanout (
		.a(new_net_701),
		.b(new_net_538),
		.c(new_net_543),
		.d(new_net_537),
		.e(new_net_535)
	);

	spl2 _0119__v_fanout (
		.a(_0119_),
		.b(new_net_496),
		.c(new_net_495)
	);

	spl2 _0264__v_fanout (
		.a(_0264_),
		.b(new_net_327),
		.c(new_net_326)
	);

	spl2 _0088__v_fanout (
		.a(_0088_),
		.b(new_net_103),
		.c(new_net_102)
	);

	spl2 new_net_697_v_fanout (
		.a(new_net_697),
		.b(new_net_182),
		.c(new_net_181)
	);

	spl4L new_net_652_v_fanout (
		.a(new_net_652),
		.b(new_net_550),
		.c(new_net_546),
		.d(new_net_547),
		.e(new_net_549)
	);

	spl2 _0267__v_fanout (
		.a(_0267_),
		.b(new_net_390),
		.c(new_net_389)
	);

	spl4L new_net_698_v_fanout (
		.a(new_net_698),
		.b(new_net_175),
		.c(new_net_174),
		.d(new_net_177),
		.e(new_net_178)
	);

	spl2 _0137__v_fanout (
		.a(_0137_),
		.b(new_net_290),
		.c(new_net_289)
	);

	spl4L new_net_692_v_fanout (
		.a(new_net_692),
		.b(new_net_121),
		.c(new_net_118),
		.d(new_net_122),
		.e(new_net_119)
	);

	spl2 _0122__v_fanout (
		.a(_0122_),
		.b(new_net_490),
		.c(new_net_489)
	);

	spl2 new_net_700_v_fanout (
		.a(new_net_700),
		.b(new_net_542),
		.c(new_net_541)
	);

	spl2 new_net_642_v_fanout (
		.a(new_net_642),
		.b(new_net_405),
		.c(new_net_399)
	);

	spl3L _0005__v_fanout (
		.a(_0005_),
		.b(new_net_692),
		.c(new_net_691),
		.d(new_net_693)
	);

	spl4L new_net_646_v_fanout (
		.a(new_net_646),
		.b(new_net_403),
		.c(new_net_402),
		.d(new_net_391),
		.e(new_net_409)
	);

	spl2 _0097__v_fanout (
		.a(_0097_),
		.b(new_net_349),
		.c(new_net_348)
	);

	spl3L _0000__v_fanout (
		.a(_0000_),
		.b(new_net_694),
		.c(new_net_695),
		.d(new_net_696)
	);

	spl4L new_net_647_v_fanout (
		.a(new_net_647),
		.b(new_net_401),
		.c(new_net_393),
		.d(new_net_397),
		.e(new_net_395)
	);

	spl4L new_net_645_v_fanout (
		.a(new_net_645),
		.b(new_net_410),
		.c(new_net_406),
		.d(new_net_412),
		.e(new_net_394)
	);

	spl3L _0007__v_fanout (
		.a(_0007_),
		.b(new_net_698),
		.c(new_net_699),
		.d(new_net_697)
	);

	spl4L new_net_644_v_fanout (
		.a(new_net_644),
		.b(new_net_407),
		.c(new_net_398),
		.d(new_net_411),
		.e(new_net_408)
	);

	bfr new_net_1434_bfr_before (
		.din(new_net_1434),
		.dout(G2551)
	);

	bfr new_net_1435_bfr_before (
		.din(new_net_1435),
		.dout(new_net_1434)
	);

	bfr new_net_1436_bfr_before (
		.din(new_net_1436),
		.dout(new_net_1435)
	);

	bfr new_net_1437_bfr_before (
		.din(new_net_1437),
		.dout(new_net_1436)
	);

	bfr new_net_1438_bfr_before (
		.din(new_net_1438),
		.dout(new_net_1437)
	);

	bfr new_net_1439_bfr_before (
		.din(new_net_1439),
		.dout(new_net_1438)
	);

	bfr new_net_1440_bfr_before (
		.din(new_net_1440),
		.dout(new_net_1439)
	);

	bfr new_net_1441_bfr_before (
		.din(new_net_1441),
		.dout(new_net_1440)
	);

	bfr new_net_1442_bfr_before (
		.din(new_net_1442),
		.dout(new_net_1441)
	);

	bfr new_net_1443_bfr_before (
		.din(new_net_1443),
		.dout(new_net_1442)
	);

	bfr new_net_1444_bfr_before (
		.din(new_net_1444),
		.dout(new_net_1443)
	);

	bfr new_net_1445_bfr_before (
		.din(new_net_1445),
		.dout(new_net_1444)
	);

	bfr new_net_1446_bfr_before (
		.din(new_net_1446),
		.dout(new_net_1445)
	);

	bfr new_net_1447_bfr_before (
		.din(new_net_1447),
		.dout(new_net_1446)
	);

	bfr new_net_1448_bfr_before (
		.din(new_net_1448),
		.dout(new_net_1447)
	);

	bfr new_net_1449_bfr_before (
		.din(new_net_1449),
		.dout(new_net_1448)
	);

	bfr new_net_1450_bfr_before (
		.din(new_net_1450),
		.dout(new_net_1449)
	);

	bfr new_net_1451_bfr_before (
		.din(new_net_1451),
		.dout(new_net_1450)
	);

	bfr new_net_1452_bfr_before (
		.din(new_net_1452),
		.dout(new_net_1451)
	);

	bfr new_net_1453_bfr_before (
		.din(new_net_1453),
		.dout(new_net_1452)
	);

	bfr new_net_1454_bfr_before (
		.din(new_net_1454),
		.dout(new_net_1453)
	);

	bfr new_net_1455_bfr_before (
		.din(new_net_1455),
		.dout(new_net_1454)
	);

	bfr new_net_1456_bfr_before (
		.din(new_net_1456),
		.dout(new_net_1455)
	);

	bfr new_net_1457_bfr_before (
		.din(new_net_1457),
		.dout(new_net_1456)
	);

	bfr new_net_1458_bfr_before (
		.din(new_net_1458),
		.dout(new_net_1457)
	);

	bfr new_net_1459_bfr_before (
		.din(new_net_1459),
		.dout(new_net_1458)
	);

	spl3L new_net_10_v_fanout (
		.a(new_net_10),
		.b(new_net_590),
		.c(new_net_1459),
		.d(new_net_589)
	);

	spl3L new_net_655_v_fanout (
		.a(new_net_655),
		.b(new_net_652),
		.c(new_net_651),
		.d(new_net_552)
	);

	spl2 _0100__v_fanout (
		.a(_0100_),
		.b(new_net_620),
		.c(new_net_619)
	);

	spl4L new_net_643_v_fanout (
		.a(new_net_643),
		.b(new_net_392),
		.c(new_net_404),
		.d(new_net_400),
		.e(new_net_396)
	);

	spl3L _0002__v_fanout (
		.a(_0002_),
		.b(new_net_700),
		.c(new_net_701),
		.d(new_net_702)
	);

	spl2 new_net_654_v_fanout (
		.a(new_net_654),
		.b(new_net_553),
		.c(new_net_653)
	);

	spl4L new_net_649_v_fanout (
		.a(new_net_649),
		.b(new_net_645),
		.c(new_net_642),
		.d(new_net_644),
		.e(new_net_643)
	);

	spl4L new_net_677_v_fanout (
		.a(new_net_677),
		.b(new_net_143),
		.c(new_net_131),
		.d(new_net_134),
		.e(new_net_135)
	);

	bfr new_net_1460_bfr_before (
		.din(new_net_1460),
		.dout(new_net_674)
	);

	bfr new_net_1461_bfr_before (
		.din(new_net_1461),
		.dout(new_net_1460)
	);

	bfr new_net_1462_bfr_before (
		.din(new_net_1462),
		.dout(new_net_1461)
	);

	bfr new_net_1463_bfr_before (
		.din(new_net_1463),
		.dout(new_net_1462)
	);

	bfr new_net_1464_bfr_before (
		.din(new_net_1464),
		.dout(new_net_1463)
	);

	spl2 new_net_675_v_fanout (
		.a(new_net_675),
		.b(new_net_1464),
		.c(new_net_136)
	);

	spl2 new_net_666_v_fanout (
		.a(new_net_666),
		.b(new_net_518),
		.c(new_net_511)
	);

	bfr new_net_1465_bfr_before (
		.din(new_net_1465),
		.dout(new_net_673)
	);

	bfr new_net_1466_bfr_before (
		.din(new_net_1466),
		.dout(new_net_1465)
	);

	bfr new_net_1467_bfr_before (
		.din(new_net_1467),
		.dout(new_net_1466)
	);

	bfr new_net_1468_bfr_before (
		.din(new_net_1468),
		.dout(new_net_1467)
	);

	bfr new_net_1469_bfr_before (
		.din(new_net_1469),
		.dout(new_net_1468)
	);

	spl4L new_net_676_v_fanout (
		.a(new_net_676),
		.b(new_net_1469),
		.c(new_net_146),
		.d(new_net_145),
		.e(new_net_142)
	);

	spl2 new_net_648_v_fanout (
		.a(new_net_648),
		.b(new_net_646),
		.c(new_net_647)
	);

	spl4L new_net_668_v_fanout (
		.a(new_net_668),
		.b(new_net_509),
		.c(new_net_508),
		.d(new_net_501),
		.e(new_net_507)
	);

	bfr new_net_1470_bfr_before (
		.din(new_net_1470),
		.dout(new_net_663)
	);

	bfr new_net_1471_bfr_before (
		.din(new_net_1471),
		.dout(new_net_1470)
	);

	bfr new_net_1472_bfr_before (
		.din(new_net_1472),
		.dout(new_net_1471)
	);

	bfr new_net_1473_bfr_before (
		.din(new_net_1473),
		.dout(new_net_1472)
	);

	bfr new_net_1474_bfr_before (
		.din(new_net_1474),
		.dout(new_net_1473)
	);

	bfr new_net_1475_bfr_before (
		.din(new_net_1475),
		.dout(new_net_1474)
	);

	spl4L new_net_667_v_fanout (
		.a(new_net_667),
		.b(new_net_506),
		.c(new_net_502),
		.d(new_net_1475),
		.e(new_net_510)
	);

	bfr new_net_1476_bfr_after (
		.din(G119),
		.dout(new_net_1476)
	);

	bfr new_net_1477_bfr_after (
		.din(new_net_1476),
		.dout(new_net_1477)
	);

	bfr new_net_1478_bfr_before (
		.din(new_net_1478),
		.dout(new_net_469)
	);

	spl2 G119_v_fanout (
		.a(new_net_1477),
		.b(new_net_1478),
		.c(new_net_468)
	);

	spl2 G155_v_fanout (
		.a(G155),
		.b(new_net_414),
		.c(new_net_413)
	);

	bfr new_net_1479_bfr_before (
		.din(new_net_1479),
		.dout(new_net_637)
	);

	bfr new_net_1480_bfr_before (
		.din(new_net_1480),
		.dout(new_net_1479)
	);

	bfr new_net_1481_bfr_before (
		.din(new_net_1481),
		.dout(new_net_1480)
	);

	bfr new_net_1482_bfr_before (
		.din(new_net_1482),
		.dout(new_net_1481)
	);

	bfr new_net_1483_bfr_before (
		.din(new_net_1483),
		.dout(new_net_1482)
	);

	bfr new_net_1484_bfr_before (
		.din(new_net_1484),
		.dout(new_net_1483)
	);

	spl3L G136_v_fanout (
		.a(G136),
		.b(new_net_419),
		.c(new_net_417),
		.d(new_net_1484)
	);

	spl2 G148_v_fanout (
		.a(G148),
		.b(new_net_622),
		.c(new_net_621)
	);

	bfr new_net_1485_bfr_before (
		.din(new_net_1485),
		.dout(new_net_639)
	);

	bfr new_net_1486_bfr_before (
		.din(new_net_1486),
		.dout(new_net_1485)
	);

	bfr new_net_1487_bfr_before (
		.din(new_net_1487),
		.dout(new_net_1486)
	);

	bfr new_net_1488_bfr_before (
		.din(new_net_1488),
		.dout(new_net_1487)
	);

	bfr new_net_1489_bfr_before (
		.din(new_net_1489),
		.dout(new_net_1488)
	);

	bfr new_net_1490_bfr_before (
		.din(new_net_1490),
		.dout(new_net_1489)
	);

	bfr new_net_1491_bfr_before (
		.din(new_net_1491),
		.dout(new_net_1490)
	);

	spl3L G138_v_fanout (
		.a(G138),
		.b(new_net_483),
		.c(new_net_485),
		.d(new_net_1491)
	);

	bfr new_net_1492_bfr_before (
		.din(new_net_1492),
		.dout(G2539)
	);

	bfr new_net_1493_bfr_before (
		.din(new_net_1493),
		.dout(new_net_1492)
	);

	bfr new_net_1494_bfr_before (
		.din(new_net_1494),
		.dout(new_net_1493)
	);

	bfr new_net_1495_bfr_before (
		.din(new_net_1495),
		.dout(new_net_1494)
	);

	bfr new_net_1496_bfr_before (
		.din(new_net_1496),
		.dout(new_net_1495)
	);

	bfr new_net_1497_bfr_before (
		.din(new_net_1497),
		.dout(new_net_1496)
	);

	bfr new_net_1498_bfr_before (
		.din(new_net_1498),
		.dout(new_net_1497)
	);

	bfr new_net_1499_bfr_before (
		.din(new_net_1499),
		.dout(new_net_1498)
	);

	bfr new_net_1500_bfr_before (
		.din(new_net_1500),
		.dout(new_net_1499)
	);

	bfr new_net_1501_bfr_before (
		.din(new_net_1501),
		.dout(new_net_1500)
	);

	bfr new_net_1502_bfr_before (
		.din(new_net_1502),
		.dout(new_net_1501)
	);

	bfr new_net_1503_bfr_before (
		.din(new_net_1503),
		.dout(new_net_1502)
	);

	bfr new_net_1504_bfr_before (
		.din(new_net_1504),
		.dout(new_net_1503)
	);

	bfr new_net_1505_bfr_before (
		.din(new_net_1505),
		.dout(new_net_1504)
	);

	bfr new_net_1506_bfr_before (
		.din(new_net_1506),
		.dout(new_net_1505)
	);

	bfr new_net_1507_bfr_before (
		.din(new_net_1507),
		.dout(new_net_1506)
	);

	bfr new_net_1508_bfr_before (
		.din(new_net_1508),
		.dout(new_net_1507)
	);

	bfr new_net_1509_bfr_before (
		.din(new_net_1509),
		.dout(new_net_1508)
	);

	bfr new_net_1510_bfr_before (
		.din(new_net_1510),
		.dout(new_net_1509)
	);

	bfr new_net_1511_bfr_before (
		.din(new_net_1511),
		.dout(new_net_1510)
	);

	bfr new_net_1512_bfr_before (
		.din(new_net_1512),
		.dout(new_net_1511)
	);

	bfr new_net_1513_bfr_before (
		.din(new_net_1513),
		.dout(new_net_1512)
	);

	bfr new_net_1514_bfr_before (
		.din(new_net_1514),
		.dout(new_net_1513)
	);

	bfr new_net_1515_bfr_before (
		.din(new_net_1515),
		.dout(new_net_1514)
	);

	bfr new_net_1516_bfr_before (
		.din(new_net_1516),
		.dout(new_net_1515)
	);

	bfr new_net_1517_bfr_before (
		.din(new_net_1517),
		.dout(new_net_1516)
	);

	bfr new_net_1518_bfr_before (
		.din(new_net_1518),
		.dout(new_net_1517)
	);

	bfr new_net_1519_bfr_before (
		.din(new_net_1519),
		.dout(new_net_1518)
	);

	spl2 G32_v_fanout (
		.a(G32),
		.b(new_net_1519),
		.c(new_net_444)
	);

	bfr new_net_1520_bfr_before (
		.din(new_net_1520),
		.dout(G2540)
	);

	bfr new_net_1521_bfr_before (
		.din(new_net_1521),
		.dout(new_net_1520)
	);

	bfr new_net_1522_bfr_before (
		.din(new_net_1522),
		.dout(new_net_1521)
	);

	bfr new_net_1523_bfr_before (
		.din(new_net_1523),
		.dout(new_net_1522)
	);

	bfr new_net_1524_bfr_before (
		.din(new_net_1524),
		.dout(new_net_1523)
	);

	bfr new_net_1525_bfr_before (
		.din(new_net_1525),
		.dout(new_net_1524)
	);

	bfr new_net_1526_bfr_before (
		.din(new_net_1526),
		.dout(new_net_1525)
	);

	bfr new_net_1527_bfr_before (
		.din(new_net_1527),
		.dout(new_net_1526)
	);

	bfr new_net_1528_bfr_before (
		.din(new_net_1528),
		.dout(new_net_1527)
	);

	bfr new_net_1529_bfr_before (
		.din(new_net_1529),
		.dout(new_net_1528)
	);

	bfr new_net_1530_bfr_before (
		.din(new_net_1530),
		.dout(new_net_1529)
	);

	bfr new_net_1531_bfr_before (
		.din(new_net_1531),
		.dout(new_net_1530)
	);

	bfr new_net_1532_bfr_before (
		.din(new_net_1532),
		.dout(new_net_1531)
	);

	bfr new_net_1533_bfr_before (
		.din(new_net_1533),
		.dout(new_net_1532)
	);

	bfr new_net_1534_bfr_before (
		.din(new_net_1534),
		.dout(new_net_1533)
	);

	bfr new_net_1535_bfr_before (
		.din(new_net_1535),
		.dout(new_net_1534)
	);

	bfr new_net_1536_bfr_before (
		.din(new_net_1536),
		.dout(new_net_1535)
	);

	bfr new_net_1537_bfr_before (
		.din(new_net_1537),
		.dout(new_net_1536)
	);

	bfr new_net_1538_bfr_before (
		.din(new_net_1538),
		.dout(new_net_1537)
	);

	bfr new_net_1539_bfr_before (
		.din(new_net_1539),
		.dout(new_net_1538)
	);

	bfr new_net_1540_bfr_before (
		.din(new_net_1540),
		.dout(new_net_1539)
	);

	bfr new_net_1541_bfr_before (
		.din(new_net_1541),
		.dout(new_net_1540)
	);

	bfr new_net_1542_bfr_before (
		.din(new_net_1542),
		.dout(new_net_1541)
	);

	bfr new_net_1543_bfr_before (
		.din(new_net_1543),
		.dout(new_net_1542)
	);

	bfr new_net_1544_bfr_before (
		.din(new_net_1544),
		.dout(new_net_1543)
	);

	bfr new_net_1545_bfr_before (
		.din(new_net_1545),
		.dout(new_net_1544)
	);

	bfr new_net_1546_bfr_before (
		.din(new_net_1546),
		.dout(new_net_1545)
	);

	bfr new_net_1547_bfr_before (
		.din(new_net_1547),
		.dout(new_net_1546)
	);

	spl2 G106_v_fanout (
		.a(G106),
		.b(new_net_1547),
		.c(new_net_472)
	);

	bfr new_net_1548_bfr_before (
		.din(new_net_1548),
		.dout(G2542)
	);

	bfr new_net_1549_bfr_before (
		.din(new_net_1549),
		.dout(new_net_1548)
	);

	bfr new_net_1550_bfr_before (
		.din(new_net_1550),
		.dout(new_net_1549)
	);

	bfr new_net_1551_bfr_before (
		.din(new_net_1551),
		.dout(new_net_1550)
	);

	bfr new_net_1552_bfr_before (
		.din(new_net_1552),
		.dout(new_net_1551)
	);

	bfr new_net_1553_bfr_before (
		.din(new_net_1553),
		.dout(new_net_1552)
	);

	bfr new_net_1554_bfr_before (
		.din(new_net_1554),
		.dout(new_net_1553)
	);

	bfr new_net_1555_bfr_before (
		.din(new_net_1555),
		.dout(new_net_1554)
	);

	bfr new_net_1556_bfr_before (
		.din(new_net_1556),
		.dout(new_net_1555)
	);

	bfr new_net_1557_bfr_before (
		.din(new_net_1557),
		.dout(new_net_1556)
	);

	bfr new_net_1558_bfr_before (
		.din(new_net_1558),
		.dout(new_net_1557)
	);

	bfr new_net_1559_bfr_before (
		.din(new_net_1559),
		.dout(new_net_1558)
	);

	bfr new_net_1560_bfr_before (
		.din(new_net_1560),
		.dout(new_net_1559)
	);

	bfr new_net_1561_bfr_before (
		.din(new_net_1561),
		.dout(new_net_1560)
	);

	bfr new_net_1562_bfr_before (
		.din(new_net_1562),
		.dout(new_net_1561)
	);

	bfr new_net_1563_bfr_before (
		.din(new_net_1563),
		.dout(new_net_1562)
	);

	bfr new_net_1564_bfr_before (
		.din(new_net_1564),
		.dout(new_net_1563)
	);

	bfr new_net_1565_bfr_before (
		.din(new_net_1565),
		.dout(new_net_1564)
	);

	bfr new_net_1566_bfr_before (
		.din(new_net_1566),
		.dout(new_net_1565)
	);

	bfr new_net_1567_bfr_before (
		.din(new_net_1567),
		.dout(new_net_1566)
	);

	bfr new_net_1568_bfr_before (
		.din(new_net_1568),
		.dout(new_net_1567)
	);

	bfr new_net_1569_bfr_before (
		.din(new_net_1569),
		.dout(new_net_1568)
	);

	bfr new_net_1570_bfr_before (
		.din(new_net_1570),
		.dout(new_net_1569)
	);

	bfr new_net_1571_bfr_before (
		.din(new_net_1571),
		.dout(new_net_1570)
	);

	bfr new_net_1572_bfr_before (
		.din(new_net_1572),
		.dout(new_net_1571)
	);

	bfr new_net_1573_bfr_before (
		.din(new_net_1573),
		.dout(new_net_1572)
	);

	bfr new_net_1574_bfr_before (
		.din(new_net_1574),
		.dout(new_net_1573)
	);

	bfr new_net_1575_bfr_before (
		.din(new_net_1575),
		.dout(new_net_1574)
	);

	spl2 G76_v_fanout (
		.a(G76),
		.b(new_net_1575),
		.c(new_net_533)
	);

	bfr new_net_1576_bfr_before (
		.din(new_net_1576),
		.dout(G2545)
	);

	bfr new_net_1577_bfr_before (
		.din(new_net_1577),
		.dout(new_net_1576)
	);

	bfr new_net_1578_bfr_before (
		.din(new_net_1578),
		.dout(new_net_1577)
	);

	bfr new_net_1579_bfr_before (
		.din(new_net_1579),
		.dout(new_net_1578)
	);

	bfr new_net_1580_bfr_before (
		.din(new_net_1580),
		.dout(new_net_1579)
	);

	bfr new_net_1581_bfr_before (
		.din(new_net_1581),
		.dout(new_net_1580)
	);

	bfr new_net_1582_bfr_before (
		.din(new_net_1582),
		.dout(new_net_1581)
	);

	bfr new_net_1583_bfr_before (
		.din(new_net_1583),
		.dout(new_net_1582)
	);

	bfr new_net_1584_bfr_before (
		.din(new_net_1584),
		.dout(new_net_1583)
	);

	bfr new_net_1585_bfr_before (
		.din(new_net_1585),
		.dout(new_net_1584)
	);

	bfr new_net_1586_bfr_before (
		.din(new_net_1586),
		.dout(new_net_1585)
	);

	bfr new_net_1587_bfr_before (
		.din(new_net_1587),
		.dout(new_net_1586)
	);

	bfr new_net_1588_bfr_before (
		.din(new_net_1588),
		.dout(new_net_1587)
	);

	bfr new_net_1589_bfr_before (
		.din(new_net_1589),
		.dout(new_net_1588)
	);

	bfr new_net_1590_bfr_before (
		.din(new_net_1590),
		.dout(new_net_1589)
	);

	bfr new_net_1591_bfr_before (
		.din(new_net_1591),
		.dout(new_net_1590)
	);

	bfr new_net_1592_bfr_before (
		.din(new_net_1592),
		.dout(new_net_1591)
	);

	bfr new_net_1593_bfr_before (
		.din(new_net_1593),
		.dout(new_net_1592)
	);

	bfr new_net_1594_bfr_before (
		.din(new_net_1594),
		.dout(new_net_1593)
	);

	bfr new_net_1595_bfr_before (
		.din(new_net_1595),
		.dout(new_net_1594)
	);

	bfr new_net_1596_bfr_before (
		.din(new_net_1596),
		.dout(new_net_1595)
	);

	bfr new_net_1597_bfr_before (
		.din(new_net_1597),
		.dout(new_net_1596)
	);

	bfr new_net_1598_bfr_before (
		.din(new_net_1598),
		.dout(new_net_1597)
	);

	bfr new_net_1599_bfr_before (
		.din(new_net_1599),
		.dout(new_net_1598)
	);

	bfr new_net_1600_bfr_before (
		.din(new_net_1600),
		.dout(new_net_1599)
	);

	bfr new_net_1601_bfr_before (
		.din(new_net_1601),
		.dout(new_net_1600)
	);

	bfr new_net_1602_bfr_before (
		.din(new_net_1602),
		.dout(new_net_1601)
	);

	bfr new_net_1603_bfr_before (
		.din(new_net_1603),
		.dout(new_net_1602)
	);

	spl2 G43_v_fanout (
		.a(G43),
		.b(new_net_1603),
		.c(new_net_212)
	);

	bfr new_net_1604_bfr_before (
		.din(new_net_1604),
		.dout(new_net_641)
	);

	bfr new_net_1605_bfr_before (
		.din(new_net_1605),
		.dout(new_net_1604)
	);

	bfr new_net_1606_bfr_before (
		.din(new_net_1606),
		.dout(new_net_1605)
	);

	bfr new_net_1607_bfr_before (
		.din(new_net_1607),
		.dout(new_net_1606)
	);

	bfr new_net_1608_bfr_before (
		.din(new_net_1608),
		.dout(new_net_1607)
	);

	bfr new_net_1609_bfr_before (
		.din(new_net_1609),
		.dout(new_net_1608)
	);

	bfr new_net_1610_bfr_before (
		.din(new_net_1610),
		.dout(new_net_1609)
	);

	bfr new_net_1611_bfr_before (
		.din(new_net_1611),
		.dout(new_net_1610)
	);

	bfr new_net_1612_bfr_before (
		.din(new_net_1612),
		.dout(new_net_1611)
	);

	bfr new_net_1613_bfr_before (
		.din(new_net_1613),
		.dout(new_net_1612)
	);

	bfr new_net_1614_bfr_before (
		.din(new_net_1614),
		.dout(new_net_1613)
	);

	spl3L G133_v_fanout (
		.a(G133),
		.b(new_net_332),
		.c(new_net_331),
		.d(new_net_1614)
	);

	spl2 G117_v_fanout (
		.a(G117),
		.b(new_net_649),
		.c(new_net_648)
	);

	spl2 G152_v_fanout (
		.a(G152),
		.b(new_net_99),
		.c(new_net_98)
	);

	bfr new_net_1615_bfr_after (
		.din(G137),
		.dout(new_net_1615)
	);

	bfr new_net_1616_bfr_after (
		.din(new_net_1615),
		.dout(new_net_1616)
	);

	bfr new_net_1617_bfr_after (
		.din(new_net_1616),
		.dout(new_net_1617)
	);

	bfr new_net_1618_bfr_after (
		.din(new_net_1617),
		.dout(new_net_1618)
	);

	bfr new_net_1619_bfr_after (
		.din(new_net_1618),
		.dout(new_net_1619)
	);

	bfr new_net_1620_bfr_after (
		.din(new_net_1619),
		.dout(new_net_1620)
	);

	bfr new_net_1621_bfr_after (
		.din(new_net_1620),
		.dout(new_net_1621)
	);

	bfr new_net_1622_bfr_after (
		.din(new_net_1621),
		.dout(new_net_1622)
	);

	bfr new_net_1623_bfr_after (
		.din(new_net_1622),
		.dout(new_net_1623)
	);

	bfr new_net_1624_bfr_after (
		.din(new_net_1623),
		.dout(new_net_1624)
	);

	bfr new_net_1625_bfr_after (
		.din(new_net_1624),
		.dout(new_net_1625)
	);

	bfr new_net_1626_bfr_after (
		.din(new_net_1625),
		.dout(new_net_1626)
	);

	bfr new_net_1627_bfr_after (
		.din(new_net_1626),
		.dout(new_net_1627)
	);

	bfr new_net_1628_bfr_after (
		.din(new_net_1627),
		.dout(new_net_1628)
	);

	bfr new_net_1629_bfr_after (
		.din(new_net_1628),
		.dout(new_net_1629)
	);

	bfr new_net_1630_bfr_after (
		.din(new_net_1629),
		.dout(new_net_1630)
	);

	bfr new_net_1631_bfr_after (
		.din(new_net_1630),
		.dout(new_net_1631)
	);

	bfr new_net_1632_bfr_after (
		.din(new_net_1631),
		.dout(new_net_1632)
	);

	bfr new_net_1633_bfr_after (
		.din(new_net_1632),
		.dout(new_net_1633)
	);

	bfr new_net_1634_bfr_after (
		.din(new_net_1633),
		.dout(new_net_1634)
	);

	bfr new_net_1635_bfr_after (
		.din(new_net_1634),
		.dout(new_net_1635)
	);

	bfr new_net_1636_bfr_after (
		.din(new_net_1635),
		.dout(new_net_1636)
	);

	bfr new_net_1637_bfr_after (
		.din(new_net_1636),
		.dout(new_net_1637)
	);

	bfr new_net_1638_bfr_after (
		.din(new_net_1637),
		.dout(new_net_1638)
	);

	bfr new_net_1639_bfr_after (
		.din(new_net_1638),
		.dout(new_net_1639)
	);

	bfr new_net_1640_bfr_after (
		.din(new_net_1639),
		.dout(new_net_1640)
	);

	bfr new_net_1641_bfr_after (
		.din(new_net_1640),
		.dout(new_net_1641)
	);

	bfr new_net_1642_bfr_after (
		.din(new_net_1641),
		.dout(new_net_1642)
	);

	spl3L G137_v_fanout (
		.a(new_net_1642),
		.b(G2538),
		.c(G2536),
		.d(G2537)
	);

	bfr new_net_1643_bfr_before (
		.din(new_net_1643),
		.dout(new_net_67)
	);

	bfr new_net_1644_bfr_before (
		.din(new_net_1644),
		.dout(new_net_1643)
	);

	bfr new_net_1645_bfr_before (
		.din(new_net_1645),
		.dout(new_net_1644)
	);

	bfr new_net_1646_bfr_before (
		.din(new_net_1646),
		.dout(new_net_1645)
	);

	bfr new_net_1647_bfr_before (
		.din(new_net_1647),
		.dout(new_net_1646)
	);

	bfr new_net_1648_bfr_before (
		.din(new_net_1648),
		.dout(new_net_1647)
	);

	bfr new_net_1649_bfr_before (
		.din(new_net_1649),
		.dout(new_net_1648)
	);

	bfr new_net_1650_bfr_before (
		.din(new_net_1650),
		.dout(new_net_1649)
	);

	bfr new_net_1651_bfr_before (
		.din(new_net_1651),
		.dout(new_net_1650)
	);

	bfr new_net_1652_bfr_before (
		.din(new_net_1652),
		.dout(new_net_1651)
	);

	spl3L G144_v_fanout (
		.a(G144),
		.b(new_net_1652),
		.c(new_net_65),
		.d(new_net_66)
	);

	bfr new_net_1653_bfr_before (
		.din(new_net_1653),
		.dout(G2543)
	);

	bfr new_net_1654_bfr_before (
		.din(new_net_1654),
		.dout(new_net_1653)
	);

	bfr new_net_1655_bfr_before (
		.din(new_net_1655),
		.dout(new_net_1654)
	);

	bfr new_net_1656_bfr_before (
		.din(new_net_1656),
		.dout(new_net_1655)
	);

	bfr new_net_1657_bfr_before (
		.din(new_net_1657),
		.dout(new_net_1656)
	);

	bfr new_net_1658_bfr_before (
		.din(new_net_1658),
		.dout(new_net_1657)
	);

	bfr new_net_1659_bfr_before (
		.din(new_net_1659),
		.dout(new_net_1658)
	);

	bfr new_net_1660_bfr_before (
		.din(new_net_1660),
		.dout(new_net_1659)
	);

	bfr new_net_1661_bfr_before (
		.din(new_net_1661),
		.dout(new_net_1660)
	);

	bfr new_net_1662_bfr_before (
		.din(new_net_1662),
		.dout(new_net_1661)
	);

	bfr new_net_1663_bfr_before (
		.din(new_net_1663),
		.dout(new_net_1662)
	);

	bfr new_net_1664_bfr_before (
		.din(new_net_1664),
		.dout(new_net_1663)
	);

	bfr new_net_1665_bfr_before (
		.din(new_net_1665),
		.dout(new_net_1664)
	);

	bfr new_net_1666_bfr_before (
		.din(new_net_1666),
		.dout(new_net_1665)
	);

	bfr new_net_1667_bfr_before (
		.din(new_net_1667),
		.dout(new_net_1666)
	);

	bfr new_net_1668_bfr_before (
		.din(new_net_1668),
		.dout(new_net_1667)
	);

	bfr new_net_1669_bfr_before (
		.din(new_net_1669),
		.dout(new_net_1668)
	);

	bfr new_net_1670_bfr_before (
		.din(new_net_1670),
		.dout(new_net_1669)
	);

	bfr new_net_1671_bfr_before (
		.din(new_net_1671),
		.dout(new_net_1670)
	);

	bfr new_net_1672_bfr_before (
		.din(new_net_1672),
		.dout(new_net_1671)
	);

	bfr new_net_1673_bfr_before (
		.din(new_net_1673),
		.dout(new_net_1672)
	);

	bfr new_net_1674_bfr_before (
		.din(new_net_1674),
		.dout(new_net_1673)
	);

	bfr new_net_1675_bfr_before (
		.din(new_net_1675),
		.dout(new_net_1674)
	);

	bfr new_net_1676_bfr_before (
		.din(new_net_1676),
		.dout(new_net_1675)
	);

	bfr new_net_1677_bfr_before (
		.din(new_net_1677),
		.dout(new_net_1676)
	);

	bfr new_net_1678_bfr_before (
		.din(new_net_1678),
		.dout(new_net_1677)
	);

	bfr new_net_1679_bfr_before (
		.din(new_net_1679),
		.dout(new_net_1678)
	);

	bfr new_net_1680_bfr_before (
		.din(new_net_1680),
		.dout(new_net_1679)
	);

	spl2 G53_v_fanout (
		.a(G53),
		.b(new_net_1680),
		.c(new_net_277)
	);

	bfr new_net_1681_bfr_before (
		.din(new_net_1681),
		.dout(new_net_650)
	);

	bfr new_net_1682_bfr_before (
		.din(new_net_1682),
		.dout(new_net_1681)
	);

	bfr new_net_1683_bfr_before (
		.din(new_net_1683),
		.dout(new_net_1682)
	);

	bfr new_net_1684_bfr_before (
		.din(new_net_1684),
		.dout(new_net_1683)
	);

	bfr new_net_1685_bfr_before (
		.din(new_net_1685),
		.dout(new_net_1684)
	);

	bfr new_net_1686_bfr_before (
		.din(new_net_1686),
		.dout(new_net_1685)
	);

	bfr new_net_1687_bfr_before (
		.din(new_net_1687),
		.dout(new_net_1686)
	);

	spl3L G143_v_fanout (
		.a(G143),
		.b(new_net_1687),
		.c(new_net_48),
		.d(new_net_51)
	);

	bfr new_net_1688_bfr_after (
		.din(G29),
		.dout(new_net_1688)
	);

	bfr new_net_1689_bfr_after (
		.din(new_net_1688),
		.dout(new_net_1689)
	);

	bfr new_net_1690_bfr_after (
		.din(new_net_1689),
		.dout(new_net_1690)
	);

	bfr new_net_1691_bfr_after (
		.din(new_net_1690),
		.dout(new_net_1691)
	);

	bfr new_net_1692_bfr_after (
		.din(new_net_1691),
		.dout(new_net_1692)
	);

	bfr new_net_1693_bfr_after (
		.din(new_net_1692),
		.dout(new_net_1693)
	);

	bfr new_net_1694_bfr_after (
		.din(new_net_1693),
		.dout(new_net_1694)
	);

	bfr new_net_1695_bfr_after (
		.din(new_net_1694),
		.dout(new_net_1695)
	);

	bfr new_net_1696_bfr_after (
		.din(new_net_1695),
		.dout(new_net_1696)
	);

	bfr new_net_1697_bfr_after (
		.din(new_net_1696),
		.dout(new_net_1697)
	);

	bfr new_net_1698_bfr_after (
		.din(new_net_1697),
		.dout(new_net_1698)
	);

	bfr new_net_1699_bfr_after (
		.din(new_net_1698),
		.dout(new_net_1699)
	);

	bfr new_net_1700_bfr_after (
		.din(new_net_1699),
		.dout(new_net_1700)
	);

	bfr new_net_1701_bfr_after (
		.din(new_net_1700),
		.dout(new_net_1701)
	);

	bfr new_net_1702_bfr_after (
		.din(new_net_1701),
		.dout(new_net_1702)
	);

	bfr new_net_1703_bfr_after (
		.din(new_net_1702),
		.dout(new_net_1703)
	);

	bfr new_net_1704_bfr_after (
		.din(new_net_1703),
		.dout(new_net_1704)
	);

	bfr new_net_1705_bfr_after (
		.din(new_net_1704),
		.dout(new_net_1705)
	);

	bfr new_net_1706_bfr_before (
		.din(new_net_1706),
		.dout(new_net_325)
	);

	bfr new_net_1707_bfr_before (
		.din(new_net_1707),
		.dout(new_net_1706)
	);

	spl2 G29_v_fanout (
		.a(new_net_1705),
		.b(new_net_1707),
		.c(new_net_324)
	);

	spl2 G157_v_fanout (
		.a(G157),
		.b(new_net_471),
		.c(new_net_470)
	);

	bfr new_net_1708_bfr_after (
		.din(G120),
		.dout(new_net_1708)
	);

	spl2 G120_v_fanout (
		.a(new_net_1708),
		.b(new_net_654),
		.c(new_net_655)
	);

	spl2 G156_v_fanout (
		.a(G156),
		.b(new_net_443),
		.c(new_net_442)
	);

	spl2 G151_v_fanout (
		.a(G151),
		.b(new_net_292),
		.c(new_net_291)
	);

	bfr new_net_1709_bfr_before (
		.din(new_net_1709),
		.dout(new_net_656)
	);

	bfr new_net_1710_bfr_before (
		.din(new_net_1710),
		.dout(new_net_1709)
	);

	bfr new_net_1711_bfr_before (
		.din(new_net_1711),
		.dout(new_net_1710)
	);

	bfr new_net_1712_bfr_before (
		.din(new_net_1712),
		.dout(new_net_1711)
	);

	bfr new_net_1713_bfr_before (
		.din(new_net_1713),
		.dout(new_net_1712)
	);

	bfr new_net_1714_bfr_before (
		.din(new_net_1714),
		.dout(new_net_1713)
	);

	bfr new_net_1715_bfr_before (
		.din(new_net_1715),
		.dout(new_net_1714)
	);

	bfr new_net_1716_bfr_before (
		.din(new_net_1716),
		.dout(new_net_1715)
	);

	bfr new_net_1717_bfr_before (
		.din(new_net_1717),
		.dout(new_net_1716)
	);

	spl3L G141_v_fanout (
		.a(G141),
		.b(new_net_627),
		.c(new_net_623),
		.d(new_net_1717)
	);

	bfr new_net_1718_bfr_before (
		.din(new_net_1718),
		.dout(new_net_528)
	);

	bfr new_net_1719_bfr_before (
		.din(new_net_1719),
		.dout(new_net_1718)
	);

	bfr new_net_1720_bfr_before (
		.din(new_net_1720),
		.dout(new_net_1719)
	);

	bfr new_net_1721_bfr_before (
		.din(new_net_1721),
		.dout(new_net_1720)
	);

	bfr new_net_1722_bfr_before (
		.din(new_net_1722),
		.dout(new_net_1721)
	);

	bfr new_net_1723_bfr_before (
		.din(new_net_1723),
		.dout(new_net_1722)
	);

	bfr new_net_1724_bfr_before (
		.din(new_net_1724),
		.dout(new_net_1723)
	);

	bfr new_net_1725_bfr_before (
		.din(new_net_1725),
		.dout(new_net_1724)
	);

	bfr new_net_1726_bfr_before (
		.din(new_net_1726),
		.dout(new_net_1725)
	);

	bfr new_net_1727_bfr_before (
		.din(new_net_1727),
		.dout(new_net_1726)
	);

	spl3L G118_v_fanout (
		.a(G118),
		.b(new_net_527),
		.c(new_net_526),
		.d(new_net_1727)
	);

	bfr new_net_1728_bfr_before (
		.din(new_net_1728),
		.dout(new_net_657)
	);

	bfr new_net_1729_bfr_before (
		.din(new_net_1729),
		.dout(new_net_1728)
	);

	bfr new_net_1730_bfr_before (
		.din(new_net_1730),
		.dout(new_net_1729)
	);

	bfr new_net_1731_bfr_before (
		.din(new_net_1731),
		.dout(new_net_1730)
	);

	bfr new_net_1732_bfr_before (
		.din(new_net_1732),
		.dout(new_net_1731)
	);

	bfr new_net_1733_bfr_before (
		.din(new_net_1733),
		.dout(new_net_1732)
	);

	bfr new_net_1734_bfr_before (
		.din(new_net_1734),
		.dout(new_net_1733)
	);

	bfr new_net_1735_bfr_before (
		.din(new_net_1735),
		.dout(new_net_1734)
	);

	bfr new_net_1736_bfr_before (
		.din(new_net_1736),
		.dout(new_net_1735)
	);

	bfr new_net_1737_bfr_before (
		.din(new_net_1737),
		.dout(new_net_1736)
	);

	spl3L G128_v_fanout (
		.a(G128),
		.b(new_net_165),
		.c(new_net_163),
		.d(new_net_1737)
	);

	bfr new_net_1738_bfr_before (
		.din(new_net_1738),
		.dout(new_net_659)
	);

	bfr new_net_1739_bfr_before (
		.din(new_net_1739),
		.dout(new_net_1738)
	);

	bfr new_net_1740_bfr_before (
		.din(new_net_1740),
		.dout(new_net_1739)
	);

	bfr new_net_1741_bfr_before (
		.din(new_net_1741),
		.dout(new_net_1740)
	);

	bfr new_net_1742_bfr_before (
		.din(new_net_1742),
		.dout(new_net_1741)
	);

	bfr new_net_1743_bfr_before (
		.din(new_net_1743),
		.dout(new_net_1742)
	);

	bfr new_net_1744_bfr_before (
		.din(new_net_1744),
		.dout(new_net_1743)
	);

	bfr new_net_1745_bfr_before (
		.din(new_net_1745),
		.dout(new_net_1744)
	);

	bfr new_net_1746_bfr_before (
		.din(new_net_1746),
		.dout(new_net_1745)
	);

	bfr new_net_1747_bfr_before (
		.din(new_net_1747),
		.dout(new_net_1746)
	);

	bfr new_net_1748_bfr_before (
		.din(new_net_1748),
		.dout(new_net_1747)
	);

	bfr new_net_1749_bfr_before (
		.din(new_net_1749),
		.dout(new_net_1748)
	);

	spl3L G131_v_fanout (
		.a(G131),
		.b(new_net_438),
		.c(new_net_439),
		.d(new_net_1749)
	);

	bfr new_net_1750_bfr_before (
		.din(new_net_1750),
		.dout(new_net_660)
	);

	bfr new_net_1751_bfr_before (
		.din(new_net_1751),
		.dout(new_net_1750)
	);

	bfr new_net_1752_bfr_before (
		.din(new_net_1752),
		.dout(new_net_1751)
	);

	bfr new_net_1753_bfr_before (
		.din(new_net_1753),
		.dout(new_net_1752)
	);

	bfr new_net_1754_bfr_before (
		.din(new_net_1754),
		.dout(new_net_1753)
	);

	bfr new_net_1755_bfr_before (
		.din(new_net_1755),
		.dout(new_net_1754)
	);

	bfr new_net_1756_bfr_before (
		.din(new_net_1756),
		.dout(new_net_1755)
	);

	bfr new_net_1757_bfr_before (
		.din(new_net_1757),
		.dout(new_net_1756)
	);

	bfr new_net_1758_bfr_before (
		.din(new_net_1758),
		.dout(new_net_1757)
	);

	spl3L G142_v_fanout (
		.a(G142),
		.b(new_net_28),
		.c(new_net_24),
		.d(new_net_1758)
	);

	bfr new_net_1759_bfr_before (
		.din(new_net_1759),
		.dout(new_net_661)
	);

	bfr new_net_1760_bfr_before (
		.din(new_net_1760),
		.dout(new_net_1759)
	);

	bfr new_net_1761_bfr_before (
		.din(new_net_1761),
		.dout(new_net_1760)
	);

	bfr new_net_1762_bfr_before (
		.din(new_net_1762),
		.dout(new_net_1761)
	);

	bfr new_net_1763_bfr_before (
		.din(new_net_1763),
		.dout(new_net_1762)
	);

	bfr new_net_1764_bfr_before (
		.din(new_net_1764),
		.dout(new_net_1763)
	);

	bfr new_net_1765_bfr_before (
		.din(new_net_1765),
		.dout(new_net_1764)
	);

	spl3L G135_v_fanout (
		.a(G135),
		.b(new_net_386),
		.c(new_net_381),
		.d(new_net_1765)
	);

	spl3L G12_v_fanout (
		.a(G12),
		.b(new_net_668),
		.c(new_net_666),
		.d(new_net_667)
	);

	bfr new_net_1766_bfr_before (
		.din(new_net_1766),
		.dout(G2541)
	);

	bfr new_net_1767_bfr_before (
		.din(new_net_1767),
		.dout(new_net_1766)
	);

	bfr new_net_1768_bfr_before (
		.din(new_net_1768),
		.dout(new_net_1767)
	);

	bfr new_net_1769_bfr_before (
		.din(new_net_1769),
		.dout(new_net_1768)
	);

	bfr new_net_1770_bfr_before (
		.din(new_net_1770),
		.dout(new_net_1769)
	);

	bfr new_net_1771_bfr_before (
		.din(new_net_1771),
		.dout(new_net_1770)
	);

	bfr new_net_1772_bfr_before (
		.din(new_net_1772),
		.dout(new_net_1771)
	);

	bfr new_net_1773_bfr_before (
		.din(new_net_1773),
		.dout(new_net_1772)
	);

	bfr new_net_1774_bfr_before (
		.din(new_net_1774),
		.dout(new_net_1773)
	);

	bfr new_net_1775_bfr_before (
		.din(new_net_1775),
		.dout(new_net_1774)
	);

	bfr new_net_1776_bfr_before (
		.din(new_net_1776),
		.dout(new_net_1775)
	);

	bfr new_net_1777_bfr_before (
		.din(new_net_1777),
		.dout(new_net_1776)
	);

	bfr new_net_1778_bfr_before (
		.din(new_net_1778),
		.dout(new_net_1777)
	);

	bfr new_net_1779_bfr_before (
		.din(new_net_1779),
		.dout(new_net_1778)
	);

	bfr new_net_1780_bfr_before (
		.din(new_net_1780),
		.dout(new_net_1779)
	);

	bfr new_net_1781_bfr_before (
		.din(new_net_1781),
		.dout(new_net_1780)
	);

	bfr new_net_1782_bfr_before (
		.din(new_net_1782),
		.dout(new_net_1781)
	);

	bfr new_net_1783_bfr_before (
		.din(new_net_1783),
		.dout(new_net_1782)
	);

	bfr new_net_1784_bfr_before (
		.din(new_net_1784),
		.dout(new_net_1783)
	);

	bfr new_net_1785_bfr_before (
		.din(new_net_1785),
		.dout(new_net_1784)
	);

	bfr new_net_1786_bfr_before (
		.din(new_net_1786),
		.dout(new_net_1785)
	);

	bfr new_net_1787_bfr_before (
		.din(new_net_1787),
		.dout(new_net_1786)
	);

	bfr new_net_1788_bfr_before (
		.din(new_net_1788),
		.dout(new_net_1787)
	);

	bfr new_net_1789_bfr_before (
		.din(new_net_1789),
		.dout(new_net_1788)
	);

	bfr new_net_1790_bfr_before (
		.din(new_net_1790),
		.dout(new_net_1789)
	);

	bfr new_net_1791_bfr_before (
		.din(new_net_1791),
		.dout(new_net_1790)
	);

	bfr new_net_1792_bfr_before (
		.din(new_net_1792),
		.dout(new_net_1791)
	);

	bfr new_net_1793_bfr_before (
		.din(new_net_1793),
		.dout(new_net_1792)
	);

	spl2 G64_v_fanout (
		.a(G64),
		.b(new_net_1793),
		.c(new_net_198)
	);

	bfr new_net_1794_bfr_before (
		.din(new_net_1794),
		.dout(new_net_669)
	);

	bfr new_net_1795_bfr_before (
		.din(new_net_1795),
		.dout(new_net_1794)
	);

	bfr new_net_1796_bfr_before (
		.din(new_net_1796),
		.dout(new_net_1795)
	);

	bfr new_net_1797_bfr_before (
		.din(new_net_1797),
		.dout(new_net_1796)
	);

	bfr new_net_1798_bfr_before (
		.din(new_net_1798),
		.dout(new_net_1797)
	);

	bfr new_net_1799_bfr_before (
		.din(new_net_1799),
		.dout(new_net_1798)
	);

	bfr new_net_1800_bfr_before (
		.din(new_net_1800),
		.dout(new_net_1799)
	);

	bfr new_net_1801_bfr_before (
		.din(new_net_1801),
		.dout(new_net_1800)
	);

	bfr new_net_1802_bfr_before (
		.din(new_net_1802),
		.dout(new_net_1801)
	);

	bfr new_net_1803_bfr_before (
		.din(new_net_1803),
		.dout(new_net_1802)
	);

	spl3L G132_v_fanout (
		.a(G132),
		.b(new_net_302),
		.c(new_net_300),
		.d(new_net_1803)
	);

	bfr new_net_1804_bfr_before (
		.din(new_net_1804),
		.dout(new_net_671)
	);

	bfr new_net_1805_bfr_before (
		.din(new_net_1805),
		.dout(new_net_1804)
	);

	bfr new_net_1806_bfr_before (
		.din(new_net_1806),
		.dout(new_net_1805)
	);

	bfr new_net_1807_bfr_before (
		.din(new_net_1807),
		.dout(new_net_1806)
	);

	bfr new_net_1808_bfr_before (
		.din(new_net_1808),
		.dout(new_net_1807)
	);

	bfr new_net_1809_bfr_before (
		.din(new_net_1809),
		.dout(new_net_1808)
	);

	bfr new_net_1810_bfr_before (
		.din(new_net_1810),
		.dout(new_net_1809)
	);

	bfr new_net_1811_bfr_before (
		.din(new_net_1811),
		.dout(new_net_1810)
	);

	bfr new_net_1812_bfr_before (
		.din(new_net_1812),
		.dout(new_net_670)
	);

	bfr new_net_1813_bfr_before (
		.din(new_net_1813),
		.dout(new_net_1812)
	);

	bfr new_net_1814_bfr_before (
		.din(new_net_1814),
		.dout(new_net_1813)
	);

	bfr new_net_1815_bfr_before (
		.din(new_net_1815),
		.dout(new_net_1814)
	);

	bfr new_net_1816_bfr_before (
		.din(new_net_1816),
		.dout(new_net_1815)
	);

	bfr new_net_1817_bfr_before (
		.din(new_net_1817),
		.dout(new_net_1816)
	);

	bfr new_net_1818_bfr_before (
		.din(new_net_1818),
		.dout(new_net_1817)
	);

	bfr new_net_1819_bfr_before (
		.din(new_net_1819),
		.dout(new_net_1818)
	);

	spl3L G123_v_fanout (
		.a(G123),
		.b(new_net_1811),
		.c(new_net_369),
		.d(new_net_1819)
	);

	bfr new_net_1820_bfr_before (
		.din(new_net_1820),
		.dout(G2546)
	);

	bfr new_net_1821_bfr_before (
		.din(new_net_1821),
		.dout(new_net_1820)
	);

	bfr new_net_1822_bfr_before (
		.din(new_net_1822),
		.dout(new_net_1821)
	);

	bfr new_net_1823_bfr_before (
		.din(new_net_1823),
		.dout(new_net_1822)
	);

	bfr new_net_1824_bfr_before (
		.din(new_net_1824),
		.dout(new_net_1823)
	);

	bfr new_net_1825_bfr_before (
		.din(new_net_1825),
		.dout(new_net_1824)
	);

	bfr new_net_1826_bfr_before (
		.din(new_net_1826),
		.dout(new_net_1825)
	);

	bfr new_net_1827_bfr_before (
		.din(new_net_1827),
		.dout(new_net_1826)
	);

	bfr new_net_1828_bfr_before (
		.din(new_net_1828),
		.dout(new_net_1827)
	);

	bfr new_net_1829_bfr_before (
		.din(new_net_1829),
		.dout(new_net_1828)
	);

	bfr new_net_1830_bfr_before (
		.din(new_net_1830),
		.dout(new_net_1829)
	);

	bfr new_net_1831_bfr_before (
		.din(new_net_1831),
		.dout(new_net_1830)
	);

	bfr new_net_1832_bfr_before (
		.din(new_net_1832),
		.dout(new_net_1831)
	);

	bfr new_net_1833_bfr_before (
		.din(new_net_1833),
		.dout(new_net_1832)
	);

	bfr new_net_1834_bfr_before (
		.din(new_net_1834),
		.dout(new_net_1833)
	);

	bfr new_net_1835_bfr_before (
		.din(new_net_1835),
		.dout(new_net_1834)
	);

	bfr new_net_1836_bfr_before (
		.din(new_net_1836),
		.dout(new_net_1835)
	);

	bfr new_net_1837_bfr_before (
		.din(new_net_1837),
		.dout(new_net_1836)
	);

	bfr new_net_1838_bfr_before (
		.din(new_net_1838),
		.dout(new_net_1837)
	);

	bfr new_net_1839_bfr_before (
		.din(new_net_1839),
		.dout(new_net_1838)
	);

	bfr new_net_1840_bfr_before (
		.din(new_net_1840),
		.dout(new_net_1839)
	);

	bfr new_net_1841_bfr_before (
		.din(new_net_1841),
		.dout(new_net_1840)
	);

	bfr new_net_1842_bfr_before (
		.din(new_net_1842),
		.dout(new_net_1841)
	);

	bfr new_net_1843_bfr_before (
		.din(new_net_1843),
		.dout(new_net_1842)
	);

	bfr new_net_1844_bfr_before (
		.din(new_net_1844),
		.dout(new_net_1843)
	);

	bfr new_net_1845_bfr_before (
		.din(new_net_1845),
		.dout(new_net_1844)
	);

	bfr new_net_1846_bfr_before (
		.din(new_net_1846),
		.dout(new_net_1845)
	);

	bfr new_net_1847_bfr_before (
		.din(new_net_1847),
		.dout(new_net_1846)
	);

	spl2 G86_v_fanout (
		.a(G86),
		.b(new_net_1847),
		.c(new_net_335)
	);

	spl4L G146_v_fanout (
		.a(G146),
		.b(new_net_115),
		.c(new_net_114),
		.d(new_net_117),
		.e(new_net_116)
	);

	bfr new_net_1848_bfr_before (
		.din(new_net_1848),
		.dout(new_net_672)
	);

	bfr new_net_1849_bfr_before (
		.din(new_net_1849),
		.dout(new_net_1848)
	);

	bfr new_net_1850_bfr_before (
		.din(new_net_1850),
		.dout(new_net_1849)
	);

	bfr new_net_1851_bfr_before (
		.din(new_net_1851),
		.dout(new_net_1850)
	);

	bfr new_net_1852_bfr_before (
		.din(new_net_1852),
		.dout(new_net_1851)
	);

	bfr new_net_1853_bfr_before (
		.din(new_net_1853),
		.dout(new_net_1852)
	);

	bfr new_net_1854_bfr_before (
		.din(new_net_1854),
		.dout(new_net_1853)
	);

	bfr new_net_1855_bfr_before (
		.din(new_net_1855),
		.dout(new_net_1854)
	);

	bfr new_net_1856_bfr_before (
		.din(new_net_1856),
		.dout(new_net_1855)
	);

	bfr new_net_1857_bfr_before (
		.din(new_net_1857),
		.dout(new_net_1856)
	);

	bfr new_net_1858_bfr_before (
		.din(new_net_1858),
		.dout(new_net_1857)
	);

	bfr new_net_1859_bfr_before (
		.din(new_net_1859),
		.dout(new_net_1858)
	);

	bfr new_net_1860_bfr_before (
		.din(new_net_1860),
		.dout(new_net_1859)
	);

	bfr new_net_1861_bfr_before (
		.din(new_net_1861),
		.dout(new_net_1860)
	);

	bfr new_net_1862_bfr_before (
		.din(new_net_1862),
		.dout(new_net_1861)
	);

	bfr new_net_1863_bfr_before (
		.din(new_net_1863),
		.dout(new_net_1862)
	);

	bfr new_net_1864_bfr_before (
		.din(new_net_1864),
		.dout(new_net_1863)
	);

	bfr new_net_1865_bfr_before (
		.din(new_net_1865),
		.dout(new_net_1864)
	);

	bfr new_net_1866_bfr_before (
		.din(new_net_1866),
		.dout(new_net_1865)
	);

	bfr new_net_1867_bfr_before (
		.din(new_net_1867),
		.dout(new_net_1866)
	);

	bfr new_net_1868_bfr_before (
		.din(new_net_1868),
		.dout(new_net_1867)
	);

	bfr new_net_1869_bfr_before (
		.din(new_net_1869),
		.dout(new_net_1868)
	);

	bfr new_net_1870_bfr_before (
		.din(new_net_1870),
		.dout(new_net_1869)
	);

	bfr new_net_1871_bfr_before (
		.din(new_net_1871),
		.dout(new_net_1870)
	);

	bfr new_net_1872_bfr_before (
		.din(new_net_1872),
		.dout(new_net_1871)
	);

	bfr new_net_1873_bfr_before (
		.din(new_net_1873),
		.dout(new_net_1872)
	);

	bfr new_net_1874_bfr_before (
		.din(new_net_1874),
		.dout(new_net_1873)
	);

	spl2 G115_v_fanout (
		.a(G115),
		.b(new_net_1874),
		.c(new_net_347)
	);

	spl3L G23_v_fanout (
		.a(G23),
		.b(new_net_676),
		.c(new_net_677),
		.d(new_net_675)
	);

	bfr new_net_1875_bfr_after (
		.din(G124),
		.dout(new_net_1875)
	);

	bfr new_net_1876_bfr_after (
		.din(new_net_1875),
		.dout(new_net_1876)
	);

	bfr new_net_1877_bfr_after (
		.din(new_net_1876),
		.dout(new_net_1877)
	);

	bfr new_net_1878_bfr_after (
		.din(new_net_1877),
		.dout(new_net_1878)
	);

	bfr new_net_1879_bfr_after (
		.din(new_net_1878),
		.dout(new_net_1879)
	);

	bfr new_net_1880_bfr_after (
		.din(new_net_1879),
		.dout(new_net_1880)
	);

	bfr new_net_1881_bfr_after (
		.din(new_net_1880),
		.dout(new_net_1881)
	);

	bfr new_net_1882_bfr_after (
		.din(new_net_1881),
		.dout(new_net_1882)
	);

	bfr new_net_1883_bfr_after (
		.din(new_net_1882),
		.dout(new_net_1883)
	);

	bfr new_net_1884_bfr_after (
		.din(new_net_1883),
		.dout(new_net_1884)
	);

	bfr new_net_1885_bfr_after (
		.din(new_net_1884),
		.dout(new_net_1885)
	);

	bfr new_net_1886_bfr_after (
		.din(new_net_1885),
		.dout(new_net_1886)
	);

	bfr new_net_1887_bfr_after (
		.din(new_net_1886),
		.dout(new_net_1887)
	);

	bfr new_net_1888_bfr_after (
		.din(new_net_1887),
		.dout(new_net_1888)
	);

	bfr new_net_1889_bfr_after (
		.din(new_net_1888),
		.dout(new_net_1889)
	);

	bfr new_net_1890_bfr_after (
		.din(new_net_1889),
		.dout(new_net_1890)
	);

	bfr new_net_1891_bfr_after (
		.din(new_net_1890),
		.dout(new_net_1891)
	);

	bfr new_net_1892_bfr_after (
		.din(new_net_1891),
		.dout(new_net_1892)
	);

	bfr new_net_1893_bfr_after (
		.din(new_net_1892),
		.dout(new_net_1893)
	);

	bfr new_net_1894_bfr_after (
		.din(new_net_1893),
		.dout(new_net_1894)
	);

	bfr new_net_1895_bfr_after (
		.din(new_net_1894),
		.dout(new_net_1895)
	);

	bfr new_net_1896_bfr_after (
		.din(new_net_1895),
		.dout(new_net_1896)
	);

	bfr new_net_1897_bfr_after (
		.din(new_net_1896),
		.dout(new_net_1897)
	);

	bfr new_net_1898_bfr_after (
		.din(new_net_1897),
		.dout(new_net_1898)
	);

	bfr new_net_1899_bfr_after (
		.din(new_net_1898),
		.dout(new_net_1899)
	);

	bfr new_net_1900_bfr_after (
		.din(new_net_1899),
		.dout(new_net_1900)
	);

	bfr new_net_1901_bfr_after (
		.din(new_net_1900),
		.dout(new_net_1901)
	);

	bfr new_net_1902_bfr_after (
		.din(new_net_1901),
		.dout(new_net_1902)
	);

	spl2 G124_v_fanout (
		.a(new_net_1902),
		.b(G2535),
		.c(G2534)
	);

	spl2 G153_v_fanout (
		.a(G153),
		.b(new_net_342),
		.c(new_net_341)
	);

	bfr new_net_1903_bfr_before (
		.din(new_net_1903),
		.dout(new_net_678)
	);

	bfr new_net_1904_bfr_before (
		.din(new_net_1904),
		.dout(new_net_1903)
	);

	bfr new_net_1905_bfr_before (
		.din(new_net_1905),
		.dout(new_net_1904)
	);

	bfr new_net_1906_bfr_before (
		.din(new_net_1906),
		.dout(new_net_1905)
	);

	bfr new_net_1907_bfr_before (
		.din(new_net_1907),
		.dout(new_net_1906)
	);

	bfr new_net_1908_bfr_before (
		.din(new_net_1908),
		.dout(new_net_1907)
	);

	bfr new_net_1909_bfr_before (
		.din(new_net_1909),
		.dout(new_net_1908)
	);

	bfr new_net_1910_bfr_before (
		.din(new_net_1910),
		.dout(new_net_1909)
	);

	bfr new_net_1911_bfr_before (
		.din(new_net_1911),
		.dout(new_net_1910)
	);

	spl3L G139_v_fanout (
		.a(G139),
		.b(new_net_520),
		.c(new_net_519),
		.d(new_net_1911)
	);

	bfr new_net_1912_bfr_before (
		.din(new_net_1912),
		.dout(new_net_679)
	);

	bfr new_net_1913_bfr_before (
		.din(new_net_1913),
		.dout(new_net_1912)
	);

	bfr new_net_1914_bfr_before (
		.din(new_net_1914),
		.dout(new_net_1913)
	);

	bfr new_net_1915_bfr_before (
		.din(new_net_1915),
		.dout(new_net_1914)
	);

	bfr new_net_1916_bfr_before (
		.din(new_net_1916),
		.dout(new_net_1915)
	);

	bfr new_net_1917_bfr_before (
		.din(new_net_1917),
		.dout(new_net_1916)
	);

	bfr new_net_1918_bfr_before (
		.din(new_net_1918),
		.dout(new_net_1917)
	);

	bfr new_net_1919_bfr_before (
		.din(new_net_1919),
		.dout(new_net_1918)
	);

	bfr new_net_1920_bfr_before (
		.din(new_net_1920),
		.dout(new_net_1919)
	);

	bfr new_net_1921_bfr_before (
		.din(new_net_1921),
		.dout(new_net_1920)
	);

	bfr new_net_1922_bfr_before (
		.din(new_net_1922),
		.dout(new_net_1921)
	);

	bfr new_net_1923_bfr_before (
		.din(new_net_1923),
		.dout(new_net_1922)
	);

	spl3L G130_v_fanout (
		.a(G130),
		.b(new_net_281),
		.c(new_net_279),
		.d(new_net_1923)
	);

	spl2 G149_v_fanout (
		.a(G149),
		.b(new_net_233),
		.c(new_net_232)
	);

	bfr new_net_1924_bfr_before (
		.din(new_net_1924),
		.dout(new_net_680)
	);

	bfr new_net_1925_bfr_before (
		.din(new_net_1925),
		.dout(new_net_1924)
	);

	bfr new_net_1926_bfr_before (
		.din(new_net_1926),
		.dout(new_net_1925)
	);

	bfr new_net_1927_bfr_before (
		.din(new_net_1927),
		.dout(new_net_1926)
	);

	bfr new_net_1928_bfr_before (
		.din(new_net_1928),
		.dout(new_net_1927)
	);

	bfr new_net_1929_bfr_before (
		.din(new_net_1929),
		.dout(new_net_1928)
	);

	bfr new_net_1930_bfr_before (
		.din(new_net_1930),
		.dout(new_net_1929)
	);

	bfr new_net_1931_bfr_before (
		.din(new_net_1931),
		.dout(new_net_1930)
	);

	bfr new_net_1932_bfr_before (
		.din(new_net_1932),
		.dout(new_net_1931)
	);

	spl3L G134_v_fanout (
		.a(G134),
		.b(new_net_355),
		.c(new_net_352),
		.d(new_net_1932)
	);

	bfr new_net_1933_bfr_before (
		.din(new_net_1933),
		.dout(new_net_682)
	);

	bfr new_net_1934_bfr_before (
		.din(new_net_1934),
		.dout(new_net_1933)
	);

	bfr new_net_1935_bfr_before (
		.din(new_net_1935),
		.dout(new_net_1934)
	);

	bfr new_net_1936_bfr_before (
		.din(new_net_1936),
		.dout(new_net_1935)
	);

	bfr new_net_1937_bfr_before (
		.din(new_net_1937),
		.dout(new_net_1936)
	);

	bfr new_net_1938_bfr_before (
		.din(new_net_1938),
		.dout(new_net_1937)
	);

	bfr new_net_1939_bfr_before (
		.din(new_net_1939),
		.dout(new_net_1938)
	);

	bfr new_net_1940_bfr_before (
		.din(new_net_1940),
		.dout(new_net_1939)
	);

	spl2 G122_v_fanout (
		.a(G122),
		.b(new_net_615),
		.c(new_net_1940)
	);

	bfr new_net_1941_bfr_before (
		.din(new_net_1941),
		.dout(new_net_683)
	);

	bfr new_net_1942_bfr_before (
		.din(new_net_1942),
		.dout(new_net_1941)
	);

	bfr new_net_1943_bfr_before (
		.din(new_net_1943),
		.dout(new_net_1942)
	);

	bfr new_net_1944_bfr_before (
		.din(new_net_1944),
		.dout(new_net_1943)
	);

	bfr new_net_1945_bfr_before (
		.din(new_net_1945),
		.dout(new_net_1944)
	);

	bfr new_net_1946_bfr_before (
		.din(new_net_1946),
		.dout(new_net_1945)
	);

	bfr new_net_1947_bfr_before (
		.din(new_net_1947),
		.dout(new_net_1946)
	);

	bfr new_net_1948_bfr_before (
		.din(new_net_1948),
		.dout(new_net_1947)
	);

	bfr new_net_1949_bfr_before (
		.din(new_net_1949),
		.dout(new_net_1948)
	);

	bfr new_net_1950_bfr_before (
		.din(new_net_1950),
		.dout(new_net_1949)
	);

	spl3L G129_v_fanout (
		.a(G129),
		.b(new_net_218),
		.c(new_net_214),
		.d(new_net_1950)
	);

	spl4L G145_v_fanout (
		.a(G145),
		.b(new_net_160),
		.c(new_net_157),
		.d(new_net_159),
		.e(new_net_158)
	);

	spl2 G150_v_fanout (
		.a(G150),
		.b(new_net_265),
		.c(new_net_264)
	);

	bfr new_net_1951_bfr_after (
		.din(G8),
		.dout(new_net_1951)
	);

	bfr new_net_1952_bfr_after (
		.din(new_net_1951),
		.dout(new_net_1952)
	);

	bfr new_net_1953_bfr_after (
		.din(new_net_1952),
		.dout(new_net_1953)
	);

	bfr new_net_1954_bfr_after (
		.din(new_net_1953),
		.dout(new_net_1954)
	);

	bfr new_net_1955_bfr_after (
		.din(new_net_1954),
		.dout(new_net_1955)
	);

	bfr new_net_1956_bfr_after (
		.din(new_net_1955),
		.dout(new_net_1956)
	);

	bfr new_net_1957_bfr_after (
		.din(new_net_1956),
		.dout(new_net_1957)
	);

	bfr new_net_1958_bfr_after (
		.din(new_net_1957),
		.dout(new_net_1958)
	);

	bfr new_net_1959_bfr_after (
		.din(new_net_1958),
		.dout(new_net_1959)
	);

	bfr new_net_1960_bfr_after (
		.din(new_net_1959),
		.dout(new_net_1960)
	);

	bfr new_net_1961_bfr_before (
		.din(new_net_1961),
		.dout(new_net_685)
	);

	spl3L G8_v_fanout (
		.a(new_net_1960),
		.b(new_net_129),
		.c(new_net_1961),
		.d(new_net_128)
	);

	bfr new_net_1962_bfr_before (
		.din(new_net_1962),
		.dout(G2544)
	);

	bfr new_net_1963_bfr_before (
		.din(new_net_1963),
		.dout(new_net_1962)
	);

	bfr new_net_1964_bfr_before (
		.din(new_net_1964),
		.dout(new_net_1963)
	);

	bfr new_net_1965_bfr_before (
		.din(new_net_1965),
		.dout(new_net_1964)
	);

	bfr new_net_1966_bfr_before (
		.din(new_net_1966),
		.dout(new_net_1965)
	);

	bfr new_net_1967_bfr_before (
		.din(new_net_1967),
		.dout(new_net_1966)
	);

	bfr new_net_1968_bfr_before (
		.din(new_net_1968),
		.dout(new_net_1967)
	);

	bfr new_net_1969_bfr_before (
		.din(new_net_1969),
		.dout(new_net_1968)
	);

	bfr new_net_1970_bfr_before (
		.din(new_net_1970),
		.dout(new_net_1969)
	);

	bfr new_net_1971_bfr_before (
		.din(new_net_1971),
		.dout(new_net_1970)
	);

	bfr new_net_1972_bfr_before (
		.din(new_net_1972),
		.dout(new_net_1971)
	);

	bfr new_net_1973_bfr_before (
		.din(new_net_1973),
		.dout(new_net_1972)
	);

	bfr new_net_1974_bfr_before (
		.din(new_net_1974),
		.dout(new_net_1973)
	);

	bfr new_net_1975_bfr_before (
		.din(new_net_1975),
		.dout(new_net_1974)
	);

	bfr new_net_1976_bfr_before (
		.din(new_net_1976),
		.dout(new_net_1975)
	);

	bfr new_net_1977_bfr_before (
		.din(new_net_1977),
		.dout(new_net_1976)
	);

	bfr new_net_1978_bfr_before (
		.din(new_net_1978),
		.dout(new_net_1977)
	);

	bfr new_net_1979_bfr_before (
		.din(new_net_1979),
		.dout(new_net_1978)
	);

	bfr new_net_1980_bfr_before (
		.din(new_net_1980),
		.dout(new_net_1979)
	);

	bfr new_net_1981_bfr_before (
		.din(new_net_1981),
		.dout(new_net_1980)
	);

	bfr new_net_1982_bfr_before (
		.din(new_net_1982),
		.dout(new_net_1981)
	);

	bfr new_net_1983_bfr_before (
		.din(new_net_1983),
		.dout(new_net_1982)
	);

	bfr new_net_1984_bfr_before (
		.din(new_net_1984),
		.dout(new_net_1983)
	);

	bfr new_net_1985_bfr_before (
		.din(new_net_1985),
		.dout(new_net_1984)
	);

	bfr new_net_1986_bfr_before (
		.din(new_net_1986),
		.dout(new_net_1985)
	);

	bfr new_net_1987_bfr_before (
		.din(new_net_1987),
		.dout(new_net_1986)
	);

	bfr new_net_1988_bfr_before (
		.din(new_net_1988),
		.dout(new_net_1987)
	);

	bfr new_net_1989_bfr_before (
		.din(new_net_1989),
		.dout(new_net_1988)
	);

	spl2 G96_v_fanout (
		.a(G96),
		.b(new_net_1989),
		.c(new_net_31)
	);

	bfr new_net_1990_bfr_before (
		.din(new_net_1990),
		.dout(new_net_686)
	);

	bfr new_net_1991_bfr_before (
		.din(new_net_1991),
		.dout(new_net_1990)
	);

	bfr new_net_1992_bfr_before (
		.din(new_net_1992),
		.dout(new_net_1991)
	);

	bfr new_net_1993_bfr_before (
		.din(new_net_1993),
		.dout(new_net_1992)
	);

	bfr new_net_1994_bfr_before (
		.din(new_net_1994),
		.dout(new_net_1993)
	);

	bfr new_net_1995_bfr_before (
		.din(new_net_1995),
		.dout(new_net_1994)
	);

	bfr new_net_1996_bfr_before (
		.din(new_net_1996),
		.dout(new_net_1995)
	);

	bfr new_net_1997_bfr_before (
		.din(new_net_1997),
		.dout(new_net_1996)
	);

	bfr new_net_1998_bfr_before (
		.din(new_net_1998),
		.dout(new_net_1997)
	);

	bfr new_net_1999_bfr_before (
		.din(new_net_1999),
		.dout(new_net_1998)
	);

	bfr new_net_2000_bfr_before (
		.din(new_net_2000),
		.dout(new_net_1999)
	);

	spl3L G125_v_fanout (
		.a(G125),
		.b(new_net_72),
		.c(new_net_2000),
		.d(new_net_75)
	);

	bfr new_net_2001_bfr_before (
		.din(new_net_2001),
		.dout(new_net_688)
	);

	bfr new_net_2002_bfr_before (
		.din(new_net_2002),
		.dout(new_net_2001)
	);

	bfr new_net_2003_bfr_before (
		.din(new_net_2003),
		.dout(new_net_2002)
	);

	bfr new_net_2004_bfr_before (
		.din(new_net_2004),
		.dout(new_net_2003)
	);

	bfr new_net_2005_bfr_before (
		.din(new_net_2005),
		.dout(new_net_2004)
	);

	bfr new_net_2006_bfr_before (
		.din(new_net_2006),
		.dout(new_net_2005)
	);

	bfr new_net_2007_bfr_before (
		.din(new_net_2007),
		.dout(new_net_2006)
	);

	bfr new_net_2008_bfr_before (
		.din(new_net_2008),
		.dout(new_net_2007)
	);

	bfr new_net_2009_bfr_before (
		.din(new_net_2009),
		.dout(new_net_2008)
	);

	spl3L G140_v_fanout (
		.a(G140),
		.b(new_net_580),
		.c(new_net_579),
		.d(new_net_2009)
	);

	bfr new_net_2010_bfr_after (
		.din(G147),
		.dout(new_net_2010)
	);

	bfr new_net_2011_bfr_after (
		.din(new_net_2010),
		.dout(new_net_2011)
	);

	bfr new_net_2012_bfr_before (
		.din(new_net_2012),
		.dout(new_net_156)
	);

	spl2 G147_v_fanout (
		.a(new_net_2011),
		.b(new_net_2012),
		.c(new_net_155)
	);

	spl3L G121_v_fanout (
		.a(G121),
		.b(new_net_573),
		.c(new_net_571),
		.d(new_net_572)
	);

	spl2 G154_v_fanout (
		.a(G154),
		.b(new_net_378),
		.c(new_net_377)
	);

	bfr new_net_2013_bfr_before (
		.din(new_net_2013),
		.dout(new_net_689)
	);

	bfr new_net_2014_bfr_before (
		.din(new_net_2014),
		.dout(new_net_2013)
	);

	bfr new_net_2015_bfr_before (
		.din(new_net_2015),
		.dout(new_net_2014)
	);

	bfr new_net_2016_bfr_before (
		.din(new_net_2016),
		.dout(new_net_2015)
	);

	bfr new_net_2017_bfr_before (
		.din(new_net_2017),
		.dout(new_net_2016)
	);

	bfr new_net_2018_bfr_before (
		.din(new_net_2018),
		.dout(new_net_2017)
	);

	bfr new_net_2019_bfr_before (
		.din(new_net_2019),
		.dout(new_net_2018)
	);

	bfr new_net_2020_bfr_before (
		.din(new_net_2020),
		.dout(new_net_2019)
	);

	bfr new_net_2021_bfr_before (
		.din(new_net_2021),
		.dout(new_net_2020)
	);

	bfr new_net_2022_bfr_before (
		.din(new_net_2022),
		.dout(new_net_2021)
	);

	bfr new_net_2023_bfr_before (
		.din(new_net_2023),
		.dout(new_net_2022)
	);

	spl3L G126_v_fanout (
		.a(G126),
		.b(new_net_193),
		.c(new_net_2023),
		.d(new_net_195)
	);

	bfr new_net_2024_bfr_after (
		.din(new_net_954),
		.dout(new_net_2024)
	);

	bfr new_net_2025_bfr_after (
		.din(new_net_2024),
		.dout(new_net_2025)
	);

	bfr new_net_2026_bfr_after (
		.din(new_net_2025),
		.dout(new_net_2026)
	);

	bfr new_net_2027_bfr_after (
		.din(new_net_2026),
		.dout(new_net_2027)
	);

	bfr new_net_2028_bfr_after (
		.din(new_net_2027),
		.dout(new_net_2028)
	);

	bfr new_net_2029_bfr_after (
		.din(new_net_2028),
		.dout(new_net_2029)
	);

	bfr new_net_2030_bfr_after (
		.din(new_net_2029),
		.dout(new_net_2030)
	);

	bfr new_net_2031_bfr_after (
		.din(new_net_2030),
		.dout(new_net_2031)
	);

	bfr new_net_2032_bfr_after (
		.din(new_net_2031),
		.dout(new_net_2032)
	);

	bfr new_net_2033_bfr_after (
		.din(new_net_2032),
		.dout(new_net_2033)
	);

	bfr new_net_2034_bfr_after (
		.din(new_net_2033),
		.dout(new_net_2034)
	);

	bfr new_net_2035_bfr_after (
		.din(new_net_2034),
		.dout(new_net_2035)
	);

	bfr new_net_2036_bfr_after (
		.din(new_net_2035),
		.dout(new_net_2036)
	);

	bfr new_net_2037_bfr_after (
		.din(new_net_2036),
		.dout(new_net_2037)
	);

	bfr new_net_2038_bfr_after (
		.din(new_net_2037),
		.dout(new_net_2038)
	);

	bfr new_net_2039_bfr_after (
		.din(new_net_2038),
		.dout(new_net_2039)
	);

	bfr new_net_2040_bfr_after (
		.din(new_net_2039),
		.dout(new_net_2040)
	);

	bfr new_net_2041_bfr_after (
		.din(new_net_2040),
		.dout(new_net_2041)
	);

	bfr new_net_2042_bfr_after (
		.din(new_net_2041),
		.dout(new_net_2042)
	);

	bfr new_net_2043_bfr_after (
		.din(new_net_2042),
		.dout(new_net_2043)
	);

	bfr new_net_2044_bfr_after (
		.din(new_net_2043),
		.dout(new_net_2044)
	);

	bfr new_net_2045_bfr_after (
		.din(new_net_2044),
		.dout(new_net_2045)
	);

	bfr new_net_2046_bfr_after (
		.din(new_net_2045),
		.dout(new_net_2046)
	);

	bfr new_net_2047_bfr_after (
		.din(new_net_2046),
		.dout(new_net_2047)
	);

	bfr new_net_2048_bfr_after (
		.din(new_net_2047),
		.dout(new_net_2048)
	);

	bfr new_net_2049_bfr_after (
		.din(new_net_2048),
		.dout(new_net_2049)
	);

	bfr G2550_bfr_after (
		.din(new_net_2049),
		.dout(G2550)
	);

	bfr new_net_2050_bfr_after (
		.din(_0417_),
		.dout(new_net_2050)
	);

	bfr new_net_2051_bfr_after (
		.din(new_net_2050),
		.dout(new_net_2051)
	);

	bfr new_net_2052_bfr_after (
		.din(new_net_2051),
		.dout(new_net_2052)
	);

	bfr new_net_2053_bfr_after (
		.din(new_net_2052),
		.dout(new_net_2053)
	);

	bfr new_net_2054_bfr_after (
		.din(new_net_2053),
		.dout(new_net_2054)
	);

	bfr new_net_2055_bfr_after (
		.din(new_net_2054),
		.dout(new_net_2055)
	);

	bfr new_net_2056_bfr_after (
		.din(new_net_2055),
		.dout(new_net_2056)
	);

	bfr new_net_2057_bfr_after (
		.din(new_net_2056),
		.dout(new_net_2057)
	);

	bfr new_net_929_bfr_after (
		.din(new_net_2057),
		.dout(new_net_929)
	);

	bfr new_net_840_bfr_after (
		.din(_0227_),
		.dout(new_net_840)
	);

	bfr new_net_2058_bfr_after (
		.din(_0286_),
		.dout(new_net_2058)
	);

	bfr new_net_2059_bfr_after (
		.din(new_net_2058),
		.dout(new_net_2059)
	);

	bfr new_net_867_bfr_after (
		.din(new_net_2059),
		.dout(new_net_867)
	);

	bfr new_net_2060_bfr_after (
		.din(_0283_),
		.dout(new_net_2060)
	);

	bfr new_net_2061_bfr_after (
		.din(new_net_2060),
		.dout(new_net_2061)
	);

	bfr new_net_2062_bfr_after (
		.din(new_net_2061),
		.dout(new_net_2062)
	);

	bfr new_net_2063_bfr_after (
		.din(new_net_2062),
		.dout(new_net_2063)
	);

	bfr new_net_2064_bfr_after (
		.din(new_net_2063),
		.dout(new_net_2064)
	);

	bfr new_net_2065_bfr_after (
		.din(new_net_2064),
		.dout(new_net_2065)
	);

	bfr new_net_862_bfr_after (
		.din(new_net_2065),
		.dout(new_net_862)
	);

	bfr new_net_2066_bfr_after (
		.din(_0456_),
		.dout(new_net_2066)
	);

	bfr new_net_925_bfr_after (
		.din(new_net_2066),
		.dout(new_net_925)
	);

	bfr new_net_2067_bfr_after (
		.din(G16),
		.dout(new_net_2067)
	);

	bfr new_net_889_bfr_after (
		.din(new_net_2067),
		.dout(new_net_889)
	);

	bfr new_net_2068_bfr_after (
		.din(_0327_),
		.dout(new_net_2068)
	);

	bfr new_net_2069_bfr_after (
		.din(new_net_2068),
		.dout(new_net_2069)
	);

	bfr new_net_884_bfr_after (
		.din(new_net_2069),
		.dout(new_net_884)
	);

	bfr new_net_2070_bfr_after (
		.din(_0039_),
		.dout(new_net_2070)
	);

	bfr new_net_778_bfr_after (
		.din(new_net_2070),
		.dout(new_net_778)
	);

	bfr new_net_799_bfr_after (
		.din(_0064_),
		.dout(new_net_799)
	);

	bfr new_net_2071_bfr_after (
		.din(G94),
		.dout(new_net_2071)
	);

	bfr new_net_2072_bfr_after (
		.din(new_net_2071),
		.dout(new_net_2072)
	);

	bfr new_net_2073_bfr_after (
		.din(new_net_2072),
		.dout(new_net_2073)
	);

	bfr new_net_820_bfr_after (
		.din(new_net_2073),
		.dout(new_net_820)
	);

	bfr new_net_2074_bfr_after (
		.din(G110),
		.dout(new_net_2074)
	);

	bfr new_net_2075_bfr_after (
		.din(new_net_2074),
		.dout(new_net_2075)
	);

	bfr new_net_2076_bfr_after (
		.din(new_net_2075),
		.dout(new_net_2076)
	);

	bfr new_net_753_bfr_after (
		.din(new_net_2076),
		.dout(new_net_753)
	);

	bfr new_net_2077_bfr_after (
		.din(G78),
		.dout(new_net_2077)
	);

	bfr new_net_2078_bfr_after (
		.din(new_net_2077),
		.dout(new_net_2078)
	);

	bfr new_net_2079_bfr_after (
		.din(new_net_2078),
		.dout(new_net_2079)
	);

	bfr new_net_757_bfr_after (
		.din(new_net_2079),
		.dout(new_net_757)
	);

	bfr new_net_2080_bfr_after (
		.din(G67),
		.dout(new_net_2080)
	);

	bfr new_net_2081_bfr_after (
		.din(new_net_2080),
		.dout(new_net_2081)
	);

	bfr new_net_770_bfr_after (
		.din(new_net_2081),
		.dout(new_net_770)
	);

	bfr new_net_2082_bfr_after (
		.din(G39),
		.dout(new_net_2082)
	);

	bfr new_net_2083_bfr_after (
		.din(new_net_2082),
		.dout(new_net_2083)
	);

	bfr new_net_791_bfr_after (
		.din(new_net_2083),
		.dout(new_net_791)
	);

	bfr new_net_2084_bfr_after (
		.din(G103),
		.dout(new_net_2084)
	);

	bfr new_net_2085_bfr_after (
		.din(new_net_2084),
		.dout(new_net_2085)
	);

	bfr new_net_2086_bfr_after (
		.din(new_net_2085),
		.dout(new_net_2086)
	);

	bfr new_net_812_bfr_after (
		.din(new_net_2086),
		.dout(new_net_812)
	);

	bfr new_net_2087_bfr_after (
		.din(G102),
		.dout(new_net_2087)
	);

	bfr new_net_2088_bfr_after (
		.din(new_net_2087),
		.dout(new_net_2088)
	);

	bfr new_net_2089_bfr_after (
		.din(new_net_2088),
		.dout(new_net_2089)
	);

	bfr new_net_816_bfr_after (
		.din(new_net_2089),
		.dout(new_net_816)
	);

	bfr new_net_2090_bfr_after (
		.din(G68),
		.dout(new_net_2090)
	);

	bfr new_net_2091_bfr_after (
		.din(new_net_2090),
		.dout(new_net_2091)
	);

	bfr new_net_774_bfr_after (
		.din(new_net_2091),
		.dout(new_net_774)
	);

	bfr new_net_2092_bfr_after (
		.din(G75),
		.dout(new_net_2092)
	);

	bfr new_net_2093_bfr_after (
		.din(new_net_2092),
		.dout(new_net_2093)
	);

	bfr new_net_2094_bfr_after (
		.din(new_net_2093),
		.dout(new_net_2094)
	);

	bfr new_net_827_bfr_after (
		.din(new_net_2094),
		.dout(new_net_827)
	);

	bfr new_net_2095_bfr_after (
		.din(G61),
		.dout(new_net_2095)
	);

	bfr new_net_2096_bfr_after (
		.din(new_net_2095),
		.dout(new_net_2096)
	);

	bfr new_net_2097_bfr_after (
		.din(new_net_2096),
		.dout(new_net_2097)
	);

	bfr new_net_2098_bfr_after (
		.din(new_net_2097),
		.dout(new_net_2098)
	);

	bfr new_net_2099_bfr_after (
		.din(new_net_2098),
		.dout(new_net_2099)
	);

	bfr new_net_848_bfr_after (
		.din(new_net_2099),
		.dout(new_net_848)
	);

	bfr new_net_853_bfr_after (
		.din(G7),
		.dout(new_net_853)
	);

	bfr new_net_2100_bfr_after (
		.din(_0386_),
		.dout(new_net_2100)
	);

	bfr new_net_2101_bfr_after (
		.din(new_net_2100),
		.dout(new_net_2101)
	);

	bfr new_net_911_bfr_after (
		.din(new_net_2101),
		.dout(new_net_911)
	);

	bfr new_net_916_bfr_after (
		.din(_0330_),
		.dout(new_net_916)
	);

	bfr new_net_875_bfr_after (
		.din(_0309_),
		.dout(new_net_875)
	);

	bfr new_net_2102_bfr_after (
		.din(_0486_),
		.dout(new_net_2102)
	);

	bfr new_net_2103_bfr_after (
		.din(new_net_2102),
		.dout(new_net_2103)
	);

	bfr new_net_2104_bfr_after (
		.din(new_net_2103),
		.dout(new_net_2104)
	);

	bfr new_net_2105_bfr_after (
		.din(new_net_2104),
		.dout(new_net_2105)
	);

	bfr new_net_2106_bfr_after (
		.din(new_net_2105),
		.dout(new_net_2106)
	);

	bfr new_net_2107_bfr_after (
		.din(new_net_2106),
		.dout(new_net_2107)
	);

	bfr new_net_2108_bfr_after (
		.din(new_net_2107),
		.dout(new_net_2108)
	);

	bfr new_net_2109_bfr_after (
		.din(new_net_2108),
		.dout(new_net_2109)
	);

	bfr new_net_938_bfr_after (
		.din(new_net_2109),
		.dout(new_net_938)
	);

	bfr new_net_2110_bfr_after (
		.din(_0471_),
		.dout(new_net_2110)
	);

	bfr new_net_2111_bfr_after (
		.din(new_net_2110),
		.dout(new_net_2111)
	);

	bfr new_net_933_bfr_after (
		.din(new_net_2111),
		.dout(new_net_933)
	);

	bfr new_net_2112_bfr_after (
		.din(_0354_),
		.dout(new_net_2112)
	);

	bfr new_net_2113_bfr_after (
		.din(new_net_2112),
		.dout(new_net_2113)
	);

	bfr new_net_897_bfr_after (
		.din(new_net_2113),
		.dout(new_net_897)
	);

	bfr new_net_2114_bfr_after (
		.din(G100),
		.dout(new_net_2114)
	);

	bfr new_net_2115_bfr_after (
		.din(new_net_2114),
		.dout(new_net_2115)
	);

	bfr new_net_2116_bfr_after (
		.din(new_net_2115),
		.dout(new_net_2116)
	);

	bfr new_net_752_bfr_after (
		.din(new_net_2116),
		.dout(new_net_752)
	);

	bfr new_net_2117_bfr_after (
		.din(_0301_),
		.dout(new_net_2117)
	);

	bfr new_net_2118_bfr_after (
		.din(new_net_2117),
		.dout(new_net_2118)
	);

	bfr new_net_2119_bfr_after (
		.din(new_net_2118),
		.dout(new_net_2119)
	);

	bfr new_net_2120_bfr_after (
		.din(new_net_2119),
		.dout(new_net_2120)
	);

	bfr new_net_2121_bfr_after (
		.din(new_net_2120),
		.dout(new_net_2121)
	);

	bfr new_net_871_bfr_after (
		.din(new_net_2121),
		.dout(new_net_871)
	);

	bfr new_net_2122_bfr_after (
		.din(_0348_),
		.dout(new_net_2122)
	);

	bfr new_net_893_bfr_after (
		.din(new_net_2122),
		.dout(new_net_893)
	);

	bfr new_net_2123_bfr_after (
		.din(_0272_),
		.dout(new_net_2123)
	);

	bfr new_net_2124_bfr_after (
		.din(new_net_2123),
		.dout(new_net_2124)
	);

	bfr new_net_2125_bfr_after (
		.din(new_net_2124),
		.dout(new_net_2125)
	);

	bfr new_net_2126_bfr_after (
		.din(new_net_2125),
		.dout(new_net_2126)
	);

	bfr new_net_2127_bfr_after (
		.din(new_net_2126),
		.dout(new_net_2127)
	);

	bfr new_net_2128_bfr_after (
		.din(new_net_2127),
		.dout(new_net_2128)
	);

	bfr new_net_2129_bfr_after (
		.din(new_net_2128),
		.dout(new_net_2129)
	);

	bfr new_net_857_bfr_after (
		.din(new_net_2129),
		.dout(new_net_857)
	);

	bfr new_net_920_bfr_after (
		.din(_0434_),
		.dout(new_net_920)
	);

	bfr new_net_831_bfr_after (
		.din(_0207_),
		.dout(new_net_831)
	);

	bfr new_net_2130_bfr_after (
		.din(G11),
		.dout(new_net_2130)
	);

	bfr new_net_852_bfr_after (
		.din(new_net_2130),
		.dout(new_net_852)
	);

	bfr new_net_915_bfr_after (
		.din(_0350_),
		.dout(new_net_915)
	);

	bfr new_net_2131_bfr_after (
		.din(G44),
		.dout(new_net_2131)
	);

	bfr new_net_2132_bfr_after (
		.din(new_net_2131),
		.dout(new_net_2132)
	);

	bfr new_net_2133_bfr_after (
		.din(new_net_2132),
		.dout(new_net_2133)
	);

	bfr new_net_2134_bfr_after (
		.din(new_net_2133),
		.dout(new_net_2134)
	);

	bfr new_net_2135_bfr_after (
		.din(new_net_2134),
		.dout(new_net_2135)
	);

	bfr new_net_782_bfr_after (
		.din(new_net_2135),
		.dout(new_net_782)
	);

	bfr new_net_803_bfr_after (
		.din(_0098_),
		.dout(new_net_803)
	);

	bfr new_net_2136_bfr_after (
		.din(G101),
		.dout(new_net_2136)
	);

	bfr new_net_2137_bfr_after (
		.din(new_net_2136),
		.dout(new_net_2137)
	);

	bfr new_net_2138_bfr_after (
		.din(new_net_2137),
		.dout(new_net_2138)
	);

	bfr new_net_824_bfr_after (
		.din(new_net_2138),
		.dout(new_net_824)
	);

	bfr new_net_2139_bfr_after (
		.din(G66),
		.dout(new_net_2139)
	);

	bfr new_net_2140_bfr_after (
		.din(new_net_2139),
		.dout(new_net_2140)
	);

	bfr new_net_786_bfr_after (
		.din(new_net_2140),
		.dout(new_net_786)
	);

	bfr new_net_2141_bfr_after (
		.din(G77),
		.dout(new_net_2141)
	);

	bfr new_net_2142_bfr_after (
		.din(new_net_2141),
		.dout(new_net_2142)
	);

	bfr new_net_2143_bfr_after (
		.din(new_net_2142),
		.dout(new_net_2143)
	);

	bfr new_net_807_bfr_after (
		.din(new_net_2143),
		.dout(new_net_807)
	);

	bfr new_net_2144_bfr_after (
		.din(G99),
		.dout(new_net_2144)
	);

	bfr new_net_2145_bfr_after (
		.din(new_net_2144),
		.dout(new_net_2145)
	);

	bfr new_net_2146_bfr_after (
		.din(new_net_2145),
		.dout(new_net_2146)
	);

	bfr new_net_761_bfr_after (
		.din(new_net_2146),
		.dout(new_net_761)
	);

	bfr new_net_2147_bfr_after (
		.din(G47),
		.dout(new_net_2147)
	);

	bfr new_net_2148_bfr_after (
		.din(new_net_2147),
		.dout(new_net_2148)
	);

	bfr new_net_2149_bfr_after (
		.din(new_net_2148),
		.dout(new_net_2149)
	);

	bfr new_net_2150_bfr_after (
		.din(new_net_2149),
		.dout(new_net_2150)
	);

	bfr new_net_2151_bfr_after (
		.din(new_net_2150),
		.dout(new_net_2151)
	);

	bfr new_net_765_bfr_after (
		.din(new_net_2151),
		.dout(new_net_765)
	);

	bfr new_net_2152_bfr_after (
		.din(G60),
		.dout(new_net_2152)
	);

	bfr new_net_2153_bfr_after (
		.din(new_net_2152),
		.dout(new_net_2153)
	);

	bfr new_net_2154_bfr_after (
		.din(new_net_2153),
		.dout(new_net_2154)
	);

	bfr new_net_2155_bfr_after (
		.din(new_net_2154),
		.dout(new_net_2155)
	);

	bfr new_net_2156_bfr_after (
		.din(new_net_2155),
		.dout(new_net_2156)
	);

	bfr new_net_795_bfr_after (
		.din(new_net_2156),
		.dout(new_net_795)
	);

	bfr new_net_2157_bfr_after (
		.din(G85),
		.dout(new_net_2157)
	);

	bfr new_net_2158_bfr_after (
		.din(new_net_2157),
		.dout(new_net_2158)
	);

	bfr new_net_2159_bfr_after (
		.din(new_net_2158),
		.dout(new_net_2159)
	);

	bfr new_net_828_bfr_after (
		.din(new_net_2159),
		.dout(new_net_828)
	);

	bfr new_net_2160_bfr_after (
		.din(G72),
		.dout(new_net_2160)
	);

	bfr new_net_2161_bfr_after (
		.din(new_net_2160),
		.dout(new_net_2161)
	);

	bfr new_net_845_bfr_after (
		.din(new_net_2161),
		.dout(new_net_845)
	);

	bfr new_net_2162_bfr_after (
		.din(G4),
		.dout(new_net_2162)
	);

	bfr new_net_879_bfr_after (
		.din(new_net_2162),
		.dout(new_net_879)
	);

	bfr new_net_942_bfr_after (
		.din(_0495_),
		.dout(new_net_942)
	);

	bfr new_net_2163_bfr_after (
		.din(G114),
		.dout(new_net_2163)
	);

	bfr new_net_2164_bfr_after (
		.din(new_net_2163),
		.dout(new_net_2164)
	);

	bfr new_net_2165_bfr_after (
		.din(new_net_2164),
		.dout(new_net_2165)
	);

	bfr new_net_822_bfr_after (
		.din(new_net_2165),
		.dout(new_net_822)
	);

	bfr new_net_2166_bfr_after (
		.din(_0230_),
		.dout(new_net_2166)
	);

	bfr new_net_843_bfr_after (
		.din(new_net_2166),
		.dout(new_net_843)
	);

	bfr new_net_2167_bfr_after (
		.din(_0364_),
		.dout(new_net_2167)
	);

	bfr new_net_2168_bfr_after (
		.din(new_net_2167),
		.dout(new_net_2168)
	);

	bfr new_net_2169_bfr_after (
		.din(new_net_2168),
		.dout(new_net_2169)
	);

	bfr new_net_2170_bfr_after (
		.din(new_net_2169),
		.dout(new_net_2170)
	);

	bfr new_net_2171_bfr_after (
		.din(new_net_2170),
		.dout(new_net_2171)
	);

	bfr new_net_2172_bfr_after (
		.din(new_net_2171),
		.dout(new_net_2172)
	);

	bfr new_net_2173_bfr_after (
		.din(new_net_2172),
		.dout(new_net_2173)
	);

	bfr new_net_901_bfr_after (
		.din(new_net_2173),
		.dout(new_net_901)
	);

	bfr new_net_2174_bfr_after (
		.din(_0373_),
		.dout(new_net_2174)
	);

	bfr new_net_906_bfr_after (
		.din(new_net_2174),
		.dout(new_net_906)
	);

	bfr new_net_2175_bfr_after (
		.din(G80),
		.dout(new_net_2175)
	);

	bfr new_net_2176_bfr_after (
		.din(new_net_2175),
		.dout(new_net_2176)
	);

	bfr new_net_2177_bfr_after (
		.din(new_net_2176),
		.dout(new_net_2177)
	);

	bfr new_net_750_bfr_after (
		.din(new_net_2177),
		.dout(new_net_750)
	);

	bfr new_net_2178_bfr_after (
		.din(_0418_),
		.dout(new_net_2178)
	);

	bfr new_net_2179_bfr_after (
		.din(new_net_2178),
		.dout(new_net_2179)
	);

	bfr new_net_2180_bfr_after (
		.din(new_net_2179),
		.dout(new_net_2180)
	);

	bfr new_net_2181_bfr_after (
		.din(new_net_2180),
		.dout(new_net_2181)
	);

	bfr new_net_2182_bfr_after (
		.din(new_net_2181),
		.dout(new_net_2182)
	);

	bfr new_net_2183_bfr_after (
		.din(new_net_2182),
		.dout(new_net_2183)
	);

	bfr new_net_2184_bfr_after (
		.din(new_net_2183),
		.dout(new_net_2184)
	);

	bfr new_net_928_bfr_after (
		.din(new_net_2184),
		.dout(new_net_928)
	);

	bfr new_net_2185_bfr_after (
		.din(new_net_965),
		.dout(new_net_2185)
	);

	bfr new_net_2186_bfr_after (
		.din(new_net_2185),
		.dout(new_net_2186)
	);

	bfr new_net_2187_bfr_after (
		.din(new_net_2186),
		.dout(new_net_2187)
	);

	bfr new_net_2188_bfr_after (
		.din(new_net_2187),
		.dout(new_net_2188)
	);

	bfr new_net_2189_bfr_after (
		.din(new_net_2188),
		.dout(new_net_2189)
	);

	bfr new_net_2190_bfr_after (
		.din(new_net_2189),
		.dout(new_net_2190)
	);

	bfr new_net_2191_bfr_after (
		.din(new_net_2190),
		.dout(new_net_2191)
	);

	bfr new_net_2192_bfr_after (
		.din(new_net_2191),
		.dout(new_net_2192)
	);

	bfr new_net_2193_bfr_after (
		.din(new_net_2192),
		.dout(new_net_2193)
	);

	bfr new_net_2194_bfr_after (
		.din(new_net_2193),
		.dout(new_net_2194)
	);

	bfr new_net_2195_bfr_after (
		.din(new_net_2194),
		.dout(new_net_2195)
	);

	bfr new_net_2196_bfr_after (
		.din(new_net_2195),
		.dout(new_net_2196)
	);

	bfr new_net_2197_bfr_after (
		.din(new_net_2196),
		.dout(new_net_2197)
	);

	bfr new_net_2198_bfr_after (
		.din(new_net_2197),
		.dout(new_net_2198)
	);

	bfr new_net_2199_bfr_after (
		.din(new_net_2198),
		.dout(new_net_2199)
	);

	bfr new_net_2200_bfr_after (
		.din(new_net_2199),
		.dout(new_net_2200)
	);

	bfr new_net_2201_bfr_after (
		.din(new_net_2200),
		.dout(new_net_2201)
	);

	bfr new_net_2202_bfr_after (
		.din(new_net_2201),
		.dout(new_net_2202)
	);

	bfr new_net_2203_bfr_after (
		.din(new_net_2202),
		.dout(new_net_2203)
	);

	bfr new_net_2204_bfr_after (
		.din(new_net_2203),
		.dout(new_net_2204)
	);

	bfr new_net_2205_bfr_after (
		.din(new_net_2204),
		.dout(new_net_2205)
	);

	bfr new_net_2206_bfr_after (
		.din(new_net_2205),
		.dout(new_net_2206)
	);

	bfr new_net_2207_bfr_after (
		.din(new_net_2206),
		.dout(new_net_2207)
	);

	bfr new_net_2208_bfr_after (
		.din(new_net_2207),
		.dout(new_net_2208)
	);

	bfr G2547_bfr_after (
		.din(new_net_2208),
		.dout(G2547)
	);

	bfr new_net_2209_bfr_after (
		.din(_0291_),
		.dout(new_net_2209)
	);

	bfr new_net_2210_bfr_after (
		.din(new_net_2209),
		.dout(new_net_2210)
	);

	bfr new_net_2211_bfr_after (
		.din(new_net_2210),
		.dout(new_net_2211)
	);

	bfr new_net_2212_bfr_after (
		.din(new_net_2211),
		.dout(new_net_2212)
	);

	bfr new_net_2213_bfr_after (
		.din(new_net_2212),
		.dout(new_net_2213)
	);

	bfr new_net_2214_bfr_after (
		.din(new_net_2213),
		.dout(new_net_2214)
	);

	bfr new_net_2215_bfr_after (
		.din(new_net_2214),
		.dout(new_net_2215)
	);

	bfr new_net_2216_bfr_after (
		.din(new_net_2215),
		.dout(new_net_2216)
	);

	bfr new_net_866_bfr_after (
		.din(new_net_2216),
		.dout(new_net_866)
	);

	bfr new_net_2217_bfr_after (
		.din(G19),
		.dout(new_net_2217)
	);

	bfr new_net_861_bfr_after (
		.din(new_net_2217),
		.dout(new_net_861)
	);

	bfr new_net_924_bfr_after (
		.din(_0448_),
		.dout(new_net_924)
	);

	bfr new_net_2218_bfr_after (
		.din(_0331_),
		.dout(new_net_2218)
	);

	bfr new_net_2219_bfr_after (
		.din(new_net_2218),
		.dout(new_net_2219)
	);

	bfr new_net_2220_bfr_after (
		.din(new_net_2219),
		.dout(new_net_2220)
	);

	bfr new_net_2221_bfr_after (
		.din(new_net_2220),
		.dout(new_net_2221)
	);

	bfr new_net_2222_bfr_after (
		.din(new_net_2221),
		.dout(new_net_2222)
	);

	bfr new_net_888_bfr_after (
		.din(new_net_2222),
		.dout(new_net_888)
	);

	bfr new_net_2223_bfr_after (
		.din(_0322_),
		.dout(new_net_2223)
	);

	bfr new_net_2224_bfr_after (
		.din(new_net_2223),
		.dout(new_net_2224)
	);

	bfr new_net_2225_bfr_after (
		.din(new_net_2224),
		.dout(new_net_2225)
	);

	bfr new_net_2226_bfr_after (
		.din(new_net_2225),
		.dout(new_net_2226)
	);

	bfr new_net_2227_bfr_after (
		.din(new_net_2226),
		.dout(new_net_2227)
	);

	bfr new_net_883_bfr_after (
		.din(new_net_2227),
		.dout(new_net_883)
	);

	bfr new_net_2228_bfr_after (
		.din(G50),
		.dout(new_net_2228)
	);

	bfr new_net_2229_bfr_after (
		.din(new_net_2228),
		.dout(new_net_2229)
	);

	bfr new_net_2230_bfr_after (
		.din(new_net_2229),
		.dout(new_net_2230)
	);

	bfr new_net_2231_bfr_after (
		.din(new_net_2230),
		.dout(new_net_2231)
	);

	bfr new_net_2232_bfr_after (
		.din(new_net_2231),
		.dout(new_net_2232)
	);

	bfr new_net_847_bfr_after (
		.din(new_net_2232),
		.dout(new_net_847)
	);

	bfr new_net_910_bfr_after (
		.din(_0380_),
		.dout(new_net_910)
	);

	bfr new_net_2233_bfr_after (
		.din(_0371_),
		.dout(new_net_2233)
	);

	bfr new_net_2234_bfr_after (
		.din(new_net_2233),
		.dout(new_net_2234)
	);

	bfr new_net_905_bfr_after (
		.din(new_net_2234),
		.dout(new_net_905)
	);

	bfr new_net_2235_bfr_after (
		.din(G57),
		.dout(new_net_2235)
	);

	bfr new_net_2236_bfr_after (
		.din(new_net_2235),
		.dout(new_net_2236)
	);

	bfr new_net_2237_bfr_after (
		.din(new_net_2236),
		.dout(new_net_2237)
	);

	bfr new_net_2238_bfr_after (
		.din(new_net_2237),
		.dout(new_net_2238)
	);

	bfr new_net_2239_bfr_after (
		.din(new_net_2238),
		.dout(new_net_2239)
	);

	bfr new_net_777_bfr_after (
		.din(new_net_2239),
		.dout(new_net_777)
	);

	bfr new_net_2240_bfr_after (
		.din(G70),
		.dout(new_net_2240)
	);

	bfr new_net_2241_bfr_after (
		.din(new_net_2240),
		.dout(new_net_2241)
	);

	bfr new_net_798_bfr_after (
		.din(new_net_2241),
		.dout(new_net_798)
	);

	bfr new_net_2242_bfr_after (
		.din(G84),
		.dout(new_net_2242)
	);

	bfr new_net_2243_bfr_after (
		.din(new_net_2242),
		.dout(new_net_2243)
	);

	bfr new_net_2244_bfr_after (
		.din(new_net_2243),
		.dout(new_net_2244)
	);

	bfr new_net_819_bfr_after (
		.din(new_net_2244),
		.dout(new_net_819)
	);

	bfr new_net_2245_bfr_after (
		.din(G88),
		.dout(new_net_2245)
	);

	bfr new_net_2246_bfr_after (
		.din(new_net_2245),
		.dout(new_net_2246)
	);

	bfr new_net_2247_bfr_after (
		.din(new_net_2246),
		.dout(new_net_2247)
	);

	bfr new_net_756_bfr_after (
		.din(new_net_2247),
		.dout(new_net_756)
	);

	bfr new_net_2248_bfr_after (
		.din(G35),
		.dout(new_net_2248)
	);

	bfr new_net_2249_bfr_after (
		.din(new_net_2248),
		.dout(new_net_2249)
	);

	bfr new_net_769_bfr_after (
		.din(new_net_2249),
		.dout(new_net_769)
	);

	bfr new_net_2250_bfr_after (
		.din(_0053_),
		.dout(new_net_2250)
	);

	bfr new_net_790_bfr_after (
		.din(new_net_2250),
		.dout(new_net_790)
	);

	bfr new_net_2251_bfr_after (
		.din(G93),
		.dout(new_net_2251)
	);

	bfr new_net_2252_bfr_after (
		.din(new_net_2251),
		.dout(new_net_2252)
	);

	bfr new_net_2253_bfr_after (
		.din(new_net_2252),
		.dout(new_net_2253)
	);

	bfr new_net_811_bfr_after (
		.din(new_net_2253),
		.dout(new_net_811)
	);

	bfr new_net_2254_bfr_after (
		.din(G36),
		.dout(new_net_2254)
	);

	bfr new_net_2255_bfr_after (
		.din(new_net_2254),
		.dout(new_net_2255)
	);

	bfr new_net_773_bfr_after (
		.din(new_net_2255),
		.dout(new_net_773)
	);

	bfr new_net_2256_bfr_after (
		.din(G49),
		.dout(new_net_2256)
	);

	bfr new_net_2257_bfr_after (
		.din(new_net_2256),
		.dout(new_net_2257)
	);

	bfr new_net_2258_bfr_after (
		.din(new_net_2257),
		.dout(new_net_2258)
	);

	bfr new_net_2259_bfr_after (
		.din(new_net_2258),
		.dout(new_net_2259)
	);

	bfr new_net_2260_bfr_after (
		.din(new_net_2259),
		.dout(new_net_2260)
	);

	bfr new_net_794_bfr_after (
		.din(new_net_2260),
		.dout(new_net_794)
	);

	bfr new_net_2261_bfr_after (
		.din(G82),
		.dout(new_net_2261)
	);

	bfr new_net_2262_bfr_after (
		.din(new_net_2261),
		.dout(new_net_2262)
	);

	bfr new_net_2263_bfr_after (
		.din(new_net_2262),
		.dout(new_net_2263)
	);

	bfr new_net_815_bfr_after (
		.din(new_net_2263),
		.dout(new_net_815)
	);

	bfr new_net_2264_bfr_after (
		.din(_0306_),
		.dout(new_net_2264)
	);

	bfr new_net_2265_bfr_after (
		.din(new_net_2264),
		.dout(new_net_2265)
	);

	bfr new_net_2266_bfr_after (
		.din(new_net_2265),
		.dout(new_net_2266)
	);

	bfr new_net_2267_bfr_after (
		.din(new_net_2266),
		.dout(new_net_2267)
	);

	bfr new_net_2268_bfr_after (
		.din(new_net_2267),
		.dout(new_net_2268)
	);

	bfr new_net_874_bfr_after (
		.din(new_net_2268),
		.dout(new_net_874)
	);

	bfr new_net_2269_bfr_after (
		.din(_0468_),
		.dout(new_net_2269)
	);

	bfr new_net_2270_bfr_after (
		.din(new_net_2269),
		.dout(new_net_2270)
	);

	bfr new_net_932_bfr_after (
		.din(new_net_2270),
		.dout(new_net_932)
	);

	bfr new_net_937_bfr_after (
		.din(_0482_),
		.dout(new_net_937)
	);

	bfr new_net_2271_bfr_after (
		.din(_0351_),
		.dout(new_net_2271)
	);

	bfr new_net_2272_bfr_after (
		.din(new_net_2271),
		.dout(new_net_2272)
	);

	bfr new_net_2273_bfr_after (
		.din(new_net_2272),
		.dout(new_net_2273)
	);

	bfr new_net_2274_bfr_after (
		.din(new_net_2273),
		.dout(new_net_2274)
	);

	bfr new_net_2275_bfr_after (
		.din(new_net_2274),
		.dout(new_net_2275)
	);

	bfr new_net_896_bfr_after (
		.din(new_net_2275),
		.dout(new_net_896)
	);

	bfr new_net_2276_bfr_after (
		.din(G21),
		.dout(new_net_2276)
	);

	bfr new_net_870_bfr_after (
		.din(new_net_2276),
		.dout(new_net_870)
	);

	bfr new_net_2277_bfr_after (
		.din(1'b0),
		.dout(new_net_2277)
	);

	bfr new_net_2278_bfr_after (
		.din(new_net_2277),
		.dout(new_net_2278)
	);

	bfr new_net_2279_bfr_after (
		.din(new_net_2278),
		.dout(new_net_2279)
	);

	bfr new_net_2280_bfr_after (
		.din(new_net_2279),
		.dout(new_net_2280)
	);

	bfr new_net_2281_bfr_after (
		.din(new_net_2280),
		.dout(new_net_2281)
	);

	bfr new_net_2282_bfr_after (
		.din(new_net_2281),
		.dout(new_net_2282)
	);

	bfr new_net_2283_bfr_after (
		.din(new_net_2282),
		.dout(new_net_2283)
	);

	bfr new_net_2284_bfr_after (
		.din(new_net_2283),
		.dout(new_net_2284)
	);

	bfr new_net_2285_bfr_after (
		.din(new_net_2284),
		.dout(new_net_2285)
	);

	bfr new_net_2286_bfr_after (
		.din(new_net_2285),
		.dout(new_net_2286)
	);

	bfr new_net_2287_bfr_after (
		.din(new_net_2286),
		.dout(new_net_2287)
	);

	bfr new_net_2288_bfr_after (
		.din(new_net_2287),
		.dout(new_net_2288)
	);

	bfr new_net_2289_bfr_after (
		.din(new_net_2288),
		.dout(new_net_2289)
	);

	bfr new_net_2290_bfr_after (
		.din(new_net_2289),
		.dout(new_net_2290)
	);

	bfr new_net_2291_bfr_after (
		.din(new_net_2290),
		.dout(new_net_2291)
	);

	bfr new_net_2292_bfr_after (
		.din(new_net_2291),
		.dout(new_net_2292)
	);

	bfr new_net_2293_bfr_after (
		.din(new_net_2292),
		.dout(new_net_2293)
	);

	bfr new_net_2294_bfr_after (
		.din(new_net_2293),
		.dout(new_net_2294)
	);

	bfr new_net_2295_bfr_after (
		.din(new_net_2294),
		.dout(new_net_2295)
	);

	bfr new_net_2296_bfr_after (
		.din(new_net_2295),
		.dout(new_net_2296)
	);

	bfr new_net_2297_bfr_after (
		.din(new_net_2296),
		.dout(new_net_2297)
	);

	bfr new_net_2298_bfr_after (
		.din(new_net_2297),
		.dout(new_net_2298)
	);

	bfr new_net_2299_bfr_after (
		.din(new_net_2298),
		.dout(new_net_2299)
	);

	bfr new_net_2300_bfr_after (
		.din(new_net_2299),
		.dout(new_net_2300)
	);

	bfr new_net_2301_bfr_after (
		.din(new_net_2300),
		.dout(new_net_2301)
	);

	bfr new_net_2302_bfr_after (
		.din(new_net_2301),
		.dout(new_net_2302)
	);

	bfr new_net_2303_bfr_after (
		.din(new_net_2302),
		.dout(new_net_2303)
	);

	bfr new_net_2304_bfr_after (
		.din(new_net_2303),
		.dout(new_net_2304)
	);

	bfr G2592_bfr_after (
		.din(new_net_2304),
		.dout(G2592)
	);

	bfr new_net_834_bfr_after (
		.din(_0219_),
		.dout(new_net_834)
	);

	bfr new_net_2305_bfr_after (
		.din(G90),
		.dout(new_net_2305)
	);

	bfr new_net_2306_bfr_after (
		.din(new_net_2305),
		.dout(new_net_2306)
	);

	bfr new_net_2307_bfr_after (
		.din(new_net_2306),
		.dout(new_net_2307)
	);

	bfr new_net_751_bfr_after (
		.din(new_net_2307),
		.dout(new_net_751)
	);

	bfr new_net_2308_bfr_after (
		.din(_0343_),
		.dout(new_net_2308)
	);

	bfr new_net_2309_bfr_after (
		.din(new_net_2308),
		.dout(new_net_2309)
	);

	bfr new_net_2310_bfr_after (
		.din(new_net_2309),
		.dout(new_net_2310)
	);

	bfr new_net_2311_bfr_after (
		.din(new_net_2310),
		.dout(new_net_2311)
	);

	bfr new_net_2312_bfr_after (
		.din(new_net_2311),
		.dout(new_net_2312)
	);

	bfr new_net_2313_bfr_after (
		.din(new_net_2312),
		.dout(new_net_2313)
	);

	bfr new_net_892_bfr_after (
		.din(new_net_2313),
		.dout(new_net_892)
	);

	bfr new_net_2314_bfr_after (
		.din(new_net_950),
		.dout(new_net_2314)
	);

	bfr new_net_2315_bfr_after (
		.din(new_net_2314),
		.dout(new_net_2315)
	);

	bfr new_net_2316_bfr_after (
		.din(new_net_2315),
		.dout(new_net_2316)
	);

	bfr new_net_2317_bfr_after (
		.din(new_net_2316),
		.dout(new_net_2317)
	);

	bfr new_net_2318_bfr_after (
		.din(new_net_2317),
		.dout(new_net_2318)
	);

	bfr new_net_2319_bfr_after (
		.din(new_net_2318),
		.dout(new_net_2319)
	);

	bfr new_net_2320_bfr_after (
		.din(new_net_2319),
		.dout(new_net_2320)
	);

	bfr new_net_2321_bfr_after (
		.din(new_net_2320),
		.dout(new_net_2321)
	);

	bfr new_net_2322_bfr_after (
		.din(new_net_2321),
		.dout(new_net_2322)
	);

	bfr new_net_2323_bfr_after (
		.din(new_net_2322),
		.dout(new_net_2323)
	);

	bfr new_net_2324_bfr_after (
		.din(new_net_2323),
		.dout(new_net_2324)
	);

	bfr new_net_2325_bfr_after (
		.din(new_net_2324),
		.dout(new_net_2325)
	);

	bfr new_net_2326_bfr_after (
		.din(new_net_2325),
		.dout(new_net_2326)
	);

	bfr new_net_2327_bfr_after (
		.din(new_net_2326),
		.dout(new_net_2327)
	);

	bfr new_net_2328_bfr_after (
		.din(new_net_2327),
		.dout(new_net_2328)
	);

	bfr new_net_2329_bfr_after (
		.din(new_net_2328),
		.dout(new_net_2329)
	);

	bfr new_net_2330_bfr_after (
		.din(new_net_2329),
		.dout(new_net_2330)
	);

	bfr new_net_2331_bfr_after (
		.din(new_net_2330),
		.dout(new_net_2331)
	);

	bfr G2564_bfr_after (
		.din(new_net_2331),
		.dout(G2564)
	);

	bfr new_net_2332_bfr_after (
		.din(G30),
		.dout(new_net_2332)
	);

	bfr new_net_2333_bfr_after (
		.din(new_net_2332),
		.dout(new_net_2333)
	);

	bfr new_net_2334_bfr_after (
		.din(new_net_2333),
		.dout(new_net_2334)
	);

	bfr new_net_2335_bfr_after (
		.din(new_net_2334),
		.dout(new_net_2335)
	);

	bfr new_net_2336_bfr_after (
		.din(new_net_2335),
		.dout(new_net_2336)
	);

	bfr new_net_2337_bfr_after (
		.din(new_net_2336),
		.dout(new_net_2337)
	);

	bfr new_net_2338_bfr_after (
		.din(new_net_2337),
		.dout(new_net_2338)
	);

	bfr new_net_919_bfr_after (
		.din(new_net_2338),
		.dout(new_net_919)
	);

	bfr new_net_2339_bfr_after (
		.din(G105),
		.dout(new_net_2339)
	);

	bfr new_net_2340_bfr_after (
		.din(new_net_2339),
		.dout(new_net_2340)
	);

	bfr new_net_2341_bfr_after (
		.din(new_net_2340),
		.dout(new_net_2341)
	);

	bfr new_net_830_bfr_after (
		.din(new_net_2341),
		.dout(new_net_830)
	);

	bfr new_net_851_bfr_after (
		.din(G2),
		.dout(new_net_851)
	);

	bfr new_net_2342_bfr_after (
		.din(_0393_),
		.dout(new_net_2342)
	);

	bfr new_net_914_bfr_after (
		.din(new_net_2342),
		.dout(new_net_914)
	);

	bfr new_net_2343_bfr_after (
		.din(_0313_),
		.dout(new_net_2343)
	);

	bfr new_net_2344_bfr_after (
		.din(new_net_2343),
		.dout(new_net_2344)
	);

	bfr new_net_2345_bfr_after (
		.din(new_net_2344),
		.dout(new_net_2345)
	);

	bfr new_net_2346_bfr_after (
		.din(new_net_2345),
		.dout(new_net_2346)
	);

	bfr new_net_2347_bfr_after (
		.din(new_net_2346),
		.dout(new_net_2347)
	);

	bfr new_net_2348_bfr_after (
		.din(new_net_2347),
		.dout(new_net_2348)
	);

	bfr new_net_2349_bfr_after (
		.din(new_net_2348),
		.dout(new_net_2349)
	);

	bfr new_net_878_bfr_after (
		.din(new_net_2349),
		.dout(new_net_878)
	);

	bfr new_net_2350_bfr_after (
		.din(_0494_),
		.dout(new_net_2350)
	);

	bfr new_net_2351_bfr_after (
		.din(new_net_2350),
		.dout(new_net_2351)
	);

	bfr new_net_2352_bfr_after (
		.din(new_net_2351),
		.dout(new_net_2352)
	);

	bfr new_net_2353_bfr_after (
		.din(new_net_2352),
		.dout(new_net_2353)
	);

	bfr new_net_2354_bfr_after (
		.din(new_net_2353),
		.dout(new_net_2354)
	);

	bfr new_net_2355_bfr_after (
		.din(new_net_2354),
		.dout(new_net_2355)
	);

	bfr new_net_941_bfr_after (
		.din(new_net_2355),
		.dout(new_net_941)
	);

	bfr new_net_2356_bfr_after (
		.din(_0480_),
		.dout(new_net_2356)
	);

	bfr new_net_936_bfr_after (
		.din(new_net_2356),
		.dout(new_net_936)
	);

	bfr new_net_2357_bfr_after (
		.din(G34),
		.dout(new_net_2357)
	);

	bfr new_net_2358_bfr_after (
		.din(new_net_2357),
		.dout(new_net_2358)
	);

	bfr new_net_785_bfr_after (
		.din(new_net_2358),
		.dout(new_net_785)
	);

	bfr new_net_806_bfr_after (
		.din(_0141_),
		.dout(new_net_806)
	);

	bfr new_net_2359_bfr_after (
		.din(_0067_),
		.dout(new_net_2359)
	);

	bfr new_net_802_bfr_after (
		.din(new_net_2359),
		.dout(new_net_802)
	);

	bfr new_net_2360_bfr_after (
		.din(G81),
		.dout(new_net_2360)
	);

	bfr new_net_2361_bfr_after (
		.din(new_net_2360),
		.dout(new_net_2361)
	);

	bfr new_net_2362_bfr_after (
		.din(new_net_2361),
		.dout(new_net_2362)
	);

	bfr new_net_823_bfr_after (
		.din(new_net_2362),
		.dout(new_net_823)
	);

	bfr new_net_2363_bfr_after (
		.din(G55),
		.dout(new_net_2363)
	);

	bfr new_net_2364_bfr_after (
		.din(new_net_2363),
		.dout(new_net_2364)
	);

	bfr new_net_2365_bfr_after (
		.din(new_net_2364),
		.dout(new_net_2365)
	);

	bfr new_net_2366_bfr_after (
		.din(new_net_2365),
		.dout(new_net_2366)
	);

	bfr new_net_2367_bfr_after (
		.din(new_net_2366),
		.dout(new_net_2367)
	);

	bfr new_net_789_bfr_after (
		.din(new_net_2367),
		.dout(new_net_789)
	);

	bfr new_net_2368_bfr_after (
		.din(G87),
		.dout(new_net_2368)
	);

	bfr new_net_2369_bfr_after (
		.din(new_net_2368),
		.dout(new_net_2369)
	);

	bfr new_net_2370_bfr_after (
		.din(new_net_2369),
		.dout(new_net_2370)
	);

	bfr new_net_810_bfr_after (
		.din(new_net_2370),
		.dout(new_net_810)
	);

	bfr new_net_2371_bfr_after (
		.din(G89),
		.dout(new_net_2371)
	);

	bfr new_net_2372_bfr_after (
		.din(new_net_2371),
		.dout(new_net_2372)
	);

	bfr new_net_2373_bfr_after (
		.din(new_net_2372),
		.dout(new_net_2373)
	);

	bfr new_net_760_bfr_after (
		.din(new_net_2373),
		.dout(new_net_760)
	);

	bfr new_net_764_bfr_after (
		.din(_0022_),
		.dout(new_net_764)
	);

	bfr new_net_2374_bfr_after (
		.din(G56),
		.dout(new_net_2374)
	);

	bfr new_net_2375_bfr_after (
		.din(new_net_2374),
		.dout(new_net_2375)
	);

	bfr new_net_2376_bfr_after (
		.din(new_net_2375),
		.dout(new_net_2376)
	);

	bfr new_net_2377_bfr_after (
		.din(new_net_2376),
		.dout(new_net_2377)
	);

	bfr new_net_2378_bfr_after (
		.din(new_net_2377),
		.dout(new_net_2378)
	);

	bfr new_net_768_bfr_after (
		.din(new_net_2378),
		.dout(new_net_768)
	);

	bfr new_net_781_bfr_after (
		.din(_0043_),
		.dout(new_net_781)
	);

	bfr new_net_2379_bfr_after (
		.din(G6),
		.dout(new_net_2379)
	);

	bfr new_net_900_bfr_after (
		.din(new_net_2379),
		.dout(new_net_900)
	);

	bfr new_net_2380_bfr_after (
		.din(_0460_),
		.dout(new_net_2380)
	);

	bfr new_net_2381_bfr_after (
		.din(new_net_2380),
		.dout(new_net_2381)
	);

	bfr new_net_927_bfr_after (
		.din(new_net_2381),
		.dout(new_net_927)
	);

	bfr new_net_2382_bfr_after (
		.din(G31),
		.dout(new_net_2382)
	);

	bfr new_net_2383_bfr_after (
		.din(new_net_2382),
		.dout(new_net_2383)
	);

	bfr new_net_838_bfr_after (
		.din(new_net_2383),
		.dout(new_net_838)
	);

	bfr new_net_2384_bfr_after (
		.din(G15),
		.dout(new_net_2384)
	);

	bfr new_net_865_bfr_after (
		.din(new_net_2384),
		.dout(new_net_865)
	);

	bfr new_net_2385_bfr_after (
		.din(_0278_),
		.dout(new_net_2385)
	);

	bfr new_net_2386_bfr_after (
		.din(new_net_2385),
		.dout(new_net_2386)
	);

	bfr new_net_2387_bfr_after (
		.din(new_net_2386),
		.dout(new_net_2387)
	);

	bfr new_net_2388_bfr_after (
		.din(new_net_2387),
		.dout(new_net_2388)
	);

	bfr new_net_2389_bfr_after (
		.din(new_net_2388),
		.dout(new_net_2389)
	);

	bfr new_net_2390_bfr_after (
		.din(new_net_2389),
		.dout(new_net_2390)
	);

	bfr new_net_2391_bfr_after (
		.din(new_net_2390),
		.dout(new_net_2391)
	);

	bfr new_net_2392_bfr_after (
		.din(new_net_2391),
		.dout(new_net_2392)
	);

	bfr new_net_860_bfr_after (
		.din(new_net_2392),
		.dout(new_net_860)
	);

	bfr new_net_2393_bfr_after (
		.din(_0442_),
		.dout(new_net_2393)
	);

	bfr new_net_923_bfr_after (
		.din(new_net_2393),
		.dout(new_net_923)
	);

	bfr new_net_2394_bfr_after (
		.din(G24),
		.dout(new_net_2394)
	);

	bfr new_net_887_bfr_after (
		.din(new_net_2394),
		.dout(new_net_887)
	);

	bfr new_net_2395_bfr_after (
		.din(G26),
		.dout(new_net_2395)
	);

	bfr new_net_882_bfr_after (
		.din(new_net_2395),
		.dout(new_net_882)
	);

	bfr new_net_2396_bfr_after (
		.din(_0498_),
		.dout(new_net_2396)
	);

	bfr new_net_2397_bfr_after (
		.din(new_net_2396),
		.dout(new_net_2397)
	);

	bfr new_net_2398_bfr_after (
		.din(new_net_2397),
		.dout(new_net_2398)
	);

	bfr new_net_2399_bfr_after (
		.din(new_net_2398),
		.dout(new_net_2399)
	);

	bfr new_net_2400_bfr_after (
		.din(new_net_2399),
		.dout(new_net_2400)
	);

	bfr new_net_2401_bfr_after (
		.din(new_net_2400),
		.dout(new_net_2401)
	);

	bfr new_net_945_bfr_after (
		.din(new_net_2401),
		.dout(new_net_945)
	);

	bfr new_net_909_bfr_after (
		.din(_0382_),
		.dout(new_net_909)
	);

	bfr new_net_2402_bfr_after (
		.din(_0370_),
		.dout(new_net_2402)
	);

	bfr new_net_2403_bfr_after (
		.din(new_net_2402),
		.dout(new_net_2403)
	);

	bfr new_net_2404_bfr_after (
		.din(new_net_2403),
		.dout(new_net_2404)
	);

	bfr new_net_2405_bfr_after (
		.din(new_net_2404),
		.dout(new_net_2405)
	);

	bfr new_net_2406_bfr_after (
		.din(new_net_2405),
		.dout(new_net_2406)
	);

	bfr new_net_904_bfr_after (
		.din(new_net_2406),
		.dout(new_net_904)
	);

	bfr new_net_907_bfr_after (
		.din(_0376_),
		.dout(new_net_907)
	);

	bfr new_net_2407_bfr_after (
		.din(_0466_),
		.dout(new_net_2407)
	);

	bfr new_net_2408_bfr_after (
		.din(new_net_2407),
		.dout(new_net_2408)
	);

	bfr new_net_2409_bfr_after (
		.din(new_net_2408),
		.dout(new_net_2409)
	);

	bfr new_net_931_bfr_after (
		.din(new_net_2409),
		.dout(new_net_931)
	);

	bfr new_net_2410_bfr_after (
		.din(G104),
		.dout(new_net_2410)
	);

	bfr new_net_2411_bfr_after (
		.din(new_net_2410),
		.dout(new_net_2411)
	);

	bfr new_net_2412_bfr_after (
		.din(new_net_2411),
		.dout(new_net_2412)
	);

	bfr new_net_821_bfr_after (
		.din(new_net_2412),
		.dout(new_net_821)
	);

	bfr new_net_2413_bfr_after (
		.din(G52),
		.dout(new_net_2413)
	);

	bfr new_net_2414_bfr_after (
		.din(new_net_2413),
		.dout(new_net_2414)
	);

	bfr new_net_2415_bfr_after (
		.din(new_net_2414),
		.dout(new_net_2415)
	);

	bfr new_net_2416_bfr_after (
		.din(new_net_2415),
		.dout(new_net_2416)
	);

	bfr new_net_2417_bfr_after (
		.din(new_net_2416),
		.dout(new_net_2417)
	);

	bfr new_net_842_bfr_after (
		.din(new_net_2417),
		.dout(new_net_842)
	);

	bfr new_net_2418_bfr_after (
		.din(G98),
		.dout(new_net_2418)
	);

	bfr new_net_2419_bfr_after (
		.din(new_net_2418),
		.dout(new_net_2419)
	);

	bfr new_net_2420_bfr_after (
		.din(new_net_2419),
		.dout(new_net_2420)
	);

	bfr new_net_755_bfr_after (
		.din(new_net_2420),
		.dout(new_net_755)
	);

	bfr new_net_772_bfr_after (
		.din(_0035_),
		.dout(new_net_772)
	);

	bfr new_net_2421_bfr_after (
		.din(G38),
		.dout(new_net_2421)
	);

	bfr new_net_2422_bfr_after (
		.din(new_net_2421),
		.dout(new_net_2422)
	);

	bfr new_net_797_bfr_after (
		.din(new_net_2422),
		.dout(new_net_797)
	);

	bfr new_net_2423_bfr_after (
		.din(G92),
		.dout(new_net_2423)
	);

	bfr new_net_2424_bfr_after (
		.din(new_net_2423),
		.dout(new_net_2424)
	);

	bfr new_net_2425_bfr_after (
		.din(new_net_2424),
		.dout(new_net_2425)
	);

	bfr new_net_818_bfr_after (
		.din(new_net_2425),
		.dout(new_net_818)
	);

	bfr new_net_793_bfr_after (
		.din(_0057_),
		.dout(new_net_793)
	);

	bfr new_net_2426_bfr_after (
		.din(G83),
		.dout(new_net_2426)
	);

	bfr new_net_2427_bfr_after (
		.din(new_net_2426),
		.dout(new_net_2427)
	);

	bfr new_net_2428_bfr_after (
		.din(new_net_2427),
		.dout(new_net_2428)
	);

	bfr new_net_814_bfr_after (
		.din(new_net_2428),
		.dout(new_net_814)
	);

	bfr new_net_2429_bfr_after (
		.din(G46),
		.dout(new_net_2429)
	);

	bfr new_net_2430_bfr_after (
		.din(new_net_2429),
		.dout(new_net_2430)
	);

	bfr new_net_2431_bfr_after (
		.din(new_net_2430),
		.dout(new_net_2431)
	);

	bfr new_net_2432_bfr_after (
		.din(new_net_2431),
		.dout(new_net_2432)
	);

	bfr new_net_2433_bfr_after (
		.din(new_net_2432),
		.dout(new_net_2433)
	);

	bfr new_net_776_bfr_after (
		.din(new_net_2433),
		.dout(new_net_776)
	);

	bfr new_net_2434_bfr_after (
		.din(G51),
		.dout(new_net_2434)
	);

	bfr new_net_2435_bfr_after (
		.din(new_net_2434),
		.dout(new_net_2435)
	);

	bfr new_net_2436_bfr_after (
		.din(new_net_2435),
		.dout(new_net_2436)
	);

	bfr new_net_2437_bfr_after (
		.din(new_net_2436),
		.dout(new_net_2437)
	);

	bfr new_net_2438_bfr_after (
		.din(new_net_2437),
		.dout(new_net_2438)
	);

	bfr new_net_835_bfr_after (
		.din(new_net_2438),
		.dout(new_net_835)
	);

	bfr new_net_2439_bfr_after (
		.din(G63),
		.dout(new_net_2439)
	);

	bfr new_net_2440_bfr_after (
		.din(new_net_2439),
		.dout(new_net_2440)
	);

	bfr new_net_839_bfr_after (
		.din(new_net_2440),
		.dout(new_net_839)
	);

	bfr new_net_2441_bfr_after (
		.din(G28),
		.dout(new_net_2441)
	);

	bfr new_net_2442_bfr_after (
		.din(new_net_2441),
		.dout(new_net_2442)
	);

	bfr new_net_2443_bfr_after (
		.din(new_net_2442),
		.dout(new_net_2443)
	);

	bfr new_net_2444_bfr_after (
		.din(new_net_2443),
		.dout(new_net_2444)
	);

	bfr new_net_2445_bfr_after (
		.din(new_net_2444),
		.dout(new_net_2445)
	);

	bfr new_net_2446_bfr_after (
		.din(new_net_2445),
		.dout(new_net_2446)
	);

	bfr new_net_2447_bfr_after (
		.din(new_net_2446),
		.dout(new_net_2447)
	);

	bfr new_net_2448_bfr_after (
		.din(new_net_2447),
		.dout(new_net_2448)
	);

	bfr new_net_856_bfr_after (
		.din(new_net_2448),
		.dout(new_net_856)
	);

	bfr new_net_2449_bfr_after (
		.din(_0297_),
		.dout(new_net_2449)
	);

	bfr new_net_2450_bfr_after (
		.din(new_net_2449),
		.dout(new_net_2450)
	);

	bfr new_net_2451_bfr_after (
		.din(new_net_2450),
		.dout(new_net_2451)
	);

	bfr new_net_2452_bfr_after (
		.din(new_net_2451),
		.dout(new_net_2452)
	);

	bfr new_net_2453_bfr_after (
		.din(new_net_2452),
		.dout(new_net_2453)
	);

	bfr new_net_2454_bfr_after (
		.din(new_net_2453),
		.dout(new_net_2454)
	);

	bfr new_net_2455_bfr_after (
		.din(new_net_2454),
		.dout(new_net_2455)
	);

	bfr new_net_869_bfr_after (
		.din(new_net_2455),
		.dout(new_net_869)
	);

	bfr new_net_2456_bfr_after (
		.din(G25),
		.dout(new_net_2456)
	);

	bfr new_net_895_bfr_after (
		.din(new_net_2456),
		.dout(new_net_895)
	);

	bfr new_net_2457_bfr_after (
		.din(new_net_959),
		.dout(new_net_2457)
	);

	bfr new_net_2458_bfr_after (
		.din(new_net_2457),
		.dout(new_net_2458)
	);

	bfr new_net_2459_bfr_after (
		.din(new_net_2458),
		.dout(new_net_2459)
	);

	bfr new_net_2460_bfr_after (
		.din(new_net_2459),
		.dout(new_net_2460)
	);

	bfr new_net_2461_bfr_after (
		.din(new_net_2460),
		.dout(new_net_2461)
	);

	bfr new_net_2462_bfr_after (
		.din(new_net_2461),
		.dout(new_net_2462)
	);

	bfr new_net_2463_bfr_after (
		.din(new_net_2462),
		.dout(new_net_2463)
	);

	bfr new_net_2464_bfr_after (
		.din(new_net_2463),
		.dout(new_net_2464)
	);

	bfr new_net_2465_bfr_after (
		.din(new_net_2464),
		.dout(new_net_2465)
	);

	bfr G2586_bfr_after (
		.din(new_net_2465),
		.dout(G2586)
	);

	bfr new_net_2466_bfr_after (
		.din(G73),
		.dout(new_net_2466)
	);

	bfr new_net_2467_bfr_after (
		.din(new_net_2466),
		.dout(new_net_2467)
	);

	bfr new_net_833_bfr_after (
		.din(new_net_2467),
		.dout(new_net_833)
	);

	bfr new_net_2468_bfr_after (
		.din(new_net_948),
		.dout(new_net_2468)
	);

	bfr new_net_2469_bfr_after (
		.din(new_net_2468),
		.dout(new_net_2469)
	);

	bfr new_net_2470_bfr_after (
		.din(new_net_2469),
		.dout(new_net_2470)
	);

	bfr new_net_2471_bfr_after (
		.din(new_net_2470),
		.dout(new_net_2471)
	);

	bfr new_net_2472_bfr_after (
		.din(new_net_2471),
		.dout(new_net_2472)
	);

	bfr new_net_2473_bfr_after (
		.din(new_net_2472),
		.dout(new_net_2473)
	);

	bfr new_net_2474_bfr_after (
		.din(new_net_2473),
		.dout(new_net_2474)
	);

	bfr new_net_2475_bfr_after (
		.din(new_net_2474),
		.dout(new_net_2475)
	);

	bfr new_net_2476_bfr_after (
		.din(new_net_2475),
		.dout(new_net_2476)
	);

	bfr new_net_2477_bfr_after (
		.din(new_net_2476),
		.dout(new_net_2477)
	);

	bfr new_net_2478_bfr_after (
		.din(new_net_2477),
		.dout(new_net_2478)
	);

	bfr new_net_2479_bfr_after (
		.din(new_net_2478),
		.dout(new_net_2479)
	);

	bfr new_net_2480_bfr_after (
		.din(new_net_2479),
		.dout(new_net_2480)
	);

	bfr new_net_2481_bfr_after (
		.din(new_net_2480),
		.dout(new_net_2481)
	);

	bfr new_net_2482_bfr_after (
		.din(new_net_2481),
		.dout(new_net_2482)
	);

	bfr new_net_2483_bfr_after (
		.din(new_net_2482),
		.dout(new_net_2483)
	);

	bfr G2563_bfr_after (
		.din(new_net_2483),
		.dout(G2563)
	);

	bfr new_net_2484_bfr_after (
		.din(G20),
		.dout(new_net_2484)
	);

	bfr new_net_891_bfr_after (
		.din(new_net_2484),
		.dout(new_net_891)
	);

	bfr new_net_2485_bfr_after (
		.din(_0270_),
		.dout(new_net_2485)
	);

	bfr new_net_2486_bfr_after (
		.din(new_net_2485),
		.dout(new_net_2486)
	);

	bfr new_net_2487_bfr_after (
		.din(new_net_2486),
		.dout(new_net_2487)
	);

	bfr new_net_2488_bfr_after (
		.din(new_net_2487),
		.dout(new_net_2488)
	);

	bfr new_net_855_bfr_after (
		.din(new_net_2488),
		.dout(new_net_855)
	);

	bfr new_net_2489_bfr_after (
		.din(G127),
		.dout(new_net_2489)
	);

	bfr new_net_2490_bfr_after (
		.din(new_net_2489),
		.dout(new_net_2490)
	);

	bfr new_net_2491_bfr_after (
		.din(new_net_2490),
		.dout(new_net_2491)
	);

	bfr new_net_2492_bfr_after (
		.din(new_net_2491),
		.dout(new_net_2492)
	);

	bfr new_net_2493_bfr_after (
		.din(new_net_2492),
		.dout(new_net_2493)
	);

	bfr new_net_2494_bfr_after (
		.din(new_net_2493),
		.dout(new_net_2494)
	);

	bfr new_net_2495_bfr_after (
		.din(new_net_2494),
		.dout(new_net_2495)
	);

	bfr new_net_918_bfr_after (
		.din(new_net_2495),
		.dout(new_net_918)
	);

	bfr new_net_2496_bfr_after (
		.din(_0388_),
		.dout(new_net_2496)
	);

	bfr new_net_2497_bfr_after (
		.din(new_net_2496),
		.dout(new_net_2497)
	);

	bfr new_net_2498_bfr_after (
		.din(new_net_2497),
		.dout(new_net_2498)
	);

	bfr new_net_2499_bfr_after (
		.din(new_net_2498),
		.dout(new_net_2499)
	);

	bfr new_net_2500_bfr_after (
		.din(new_net_2499),
		.dout(new_net_2500)
	);

	bfr new_net_2501_bfr_after (
		.din(new_net_2500),
		.dout(new_net_2501)
	);

	bfr new_net_913_bfr_after (
		.din(new_net_2501),
		.dout(new_net_913)
	);

	bfr new_net_2502_bfr_after (
		.din(new_net_946),
		.dout(new_net_2502)
	);

	bfr new_net_2503_bfr_after (
		.din(new_net_2502),
		.dout(new_net_2503)
	);

	bfr new_net_2504_bfr_after (
		.din(new_net_2503),
		.dout(new_net_2504)
	);

	bfr new_net_2505_bfr_after (
		.din(new_net_2504),
		.dout(new_net_2505)
	);

	bfr new_net_2506_bfr_after (
		.din(new_net_2505),
		.dout(new_net_2506)
	);

	bfr new_net_2507_bfr_after (
		.din(new_net_2506),
		.dout(new_net_2507)
	);

	bfr new_net_2508_bfr_after (
		.din(new_net_2507),
		.dout(new_net_2508)
	);

	bfr new_net_2509_bfr_after (
		.din(new_net_2508),
		.dout(new_net_2509)
	);

	bfr new_net_2510_bfr_after (
		.din(new_net_2509),
		.dout(new_net_2510)
	);

	bfr new_net_2511_bfr_after (
		.din(new_net_2510),
		.dout(new_net_2511)
	);

	bfr new_net_2512_bfr_after (
		.din(new_net_2511),
		.dout(new_net_2512)
	);

	bfr new_net_2513_bfr_after (
		.din(new_net_2512),
		.dout(new_net_2513)
	);

	bfr new_net_2514_bfr_after (
		.din(new_net_2513),
		.dout(new_net_2514)
	);

	bfr new_net_2515_bfr_after (
		.din(new_net_2514),
		.dout(new_net_2515)
	);

	bfr new_net_2516_bfr_after (
		.din(new_net_2515),
		.dout(new_net_2516)
	);

	bfr new_net_2517_bfr_after (
		.din(new_net_2516),
		.dout(new_net_2517)
	);

	bfr new_net_2518_bfr_after (
		.din(new_net_2517),
		.dout(new_net_2518)
	);

	bfr new_net_2519_bfr_after (
		.din(new_net_2518),
		.dout(new_net_2519)
	);

	bfr G2565_bfr_after (
		.din(new_net_2519),
		.dout(G2565)
	);

	bfr new_net_2520_bfr_after (
		.din(new_net_961),
		.dout(new_net_2520)
	);

	bfr new_net_2521_bfr_after (
		.din(new_net_2520),
		.dout(new_net_2521)
	);

	bfr new_net_2522_bfr_after (
		.din(new_net_2521),
		.dout(new_net_2522)
	);

	bfr new_net_2523_bfr_after (
		.din(new_net_2522),
		.dout(new_net_2523)
	);

	bfr new_net_2524_bfr_after (
		.din(new_net_2523),
		.dout(new_net_2524)
	);

	bfr new_net_2525_bfr_after (
		.din(new_net_2524),
		.dout(new_net_2525)
	);

	bfr new_net_2526_bfr_after (
		.din(new_net_2525),
		.dout(new_net_2526)
	);

	bfr new_net_2527_bfr_after (
		.din(new_net_2526),
		.dout(new_net_2527)
	);

	bfr new_net_2528_bfr_after (
		.din(new_net_2527),
		.dout(new_net_2528)
	);

	bfr new_net_2529_bfr_after (
		.din(new_net_2528),
		.dout(new_net_2529)
	);

	bfr new_net_2530_bfr_after (
		.din(new_net_2529),
		.dout(new_net_2530)
	);

	bfr new_net_2531_bfr_after (
		.din(new_net_2530),
		.dout(new_net_2531)
	);

	bfr new_net_2532_bfr_after (
		.din(new_net_2531),
		.dout(new_net_2532)
	);

	bfr new_net_2533_bfr_after (
		.din(new_net_2532),
		.dout(new_net_2533)
	);

	bfr new_net_2534_bfr_after (
		.din(new_net_2533),
		.dout(new_net_2534)
	);

	bfr new_net_2535_bfr_after (
		.din(new_net_2534),
		.dout(new_net_2535)
	);

	bfr G2577_bfr_after (
		.din(new_net_2535),
		.dout(G2577)
	);

	bfr new_net_2536_bfr_after (
		.din(G14),
		.dout(new_net_2536)
	);

	bfr new_net_877_bfr_after (
		.din(new_net_2536),
		.dout(new_net_877)
	);

	bfr new_net_940_bfr_after (
		.din(_0492_),
		.dout(new_net_940)
	);

	bfr new_net_935_bfr_after (
		.din(_0478_),
		.dout(new_net_935)
	);

	bfr new_net_2537_bfr_after (
		.din(new_net_967),
		.dout(new_net_2537)
	);

	bfr new_net_2538_bfr_after (
		.din(new_net_2537),
		.dout(new_net_2538)
	);

	bfr new_net_2539_bfr_after (
		.din(new_net_2538),
		.dout(new_net_2539)
	);

	bfr new_net_2540_bfr_after (
		.din(new_net_2539),
		.dout(new_net_2540)
	);

	bfr new_net_2541_bfr_after (
		.din(new_net_2540),
		.dout(new_net_2541)
	);

	bfr new_net_2542_bfr_after (
		.din(new_net_2541),
		.dout(new_net_2542)
	);

	bfr new_net_2543_bfr_after (
		.din(new_net_2542),
		.dout(new_net_2543)
	);

	bfr new_net_2544_bfr_after (
		.din(new_net_2543),
		.dout(new_net_2544)
	);

	bfr new_net_2545_bfr_after (
		.din(new_net_2544),
		.dout(new_net_2545)
	);

	bfr new_net_2546_bfr_after (
		.din(new_net_2545),
		.dout(new_net_2546)
	);

	bfr new_net_2547_bfr_after (
		.din(new_net_2546),
		.dout(new_net_2547)
	);

	bfr new_net_2548_bfr_after (
		.din(new_net_2547),
		.dout(new_net_2548)
	);

	bfr new_net_2549_bfr_after (
		.din(new_net_2548),
		.dout(new_net_2549)
	);

	bfr new_net_2550_bfr_after (
		.din(new_net_2549),
		.dout(new_net_2550)
	);

	bfr new_net_2551_bfr_after (
		.din(new_net_2550),
		.dout(new_net_2551)
	);

	bfr new_net_2552_bfr_after (
		.din(new_net_2551),
		.dout(new_net_2552)
	);

	bfr new_net_2553_bfr_after (
		.din(new_net_2552),
		.dout(new_net_2553)
	);

	bfr new_net_2554_bfr_after (
		.din(new_net_2553),
		.dout(new_net_2554)
	);

	bfr new_net_2555_bfr_after (
		.din(new_net_2554),
		.dout(new_net_2555)
	);

	bfr new_net_2556_bfr_after (
		.din(new_net_2555),
		.dout(new_net_2556)
	);

	bfr new_net_2557_bfr_after (
		.din(new_net_2556),
		.dout(new_net_2557)
	);

	bfr new_net_2558_bfr_after (
		.din(new_net_2557),
		.dout(new_net_2558)
	);

	bfr new_net_2559_bfr_after (
		.din(new_net_2558),
		.dout(new_net_2559)
	);

	bfr new_net_2560_bfr_after (
		.din(new_net_2559),
		.dout(new_net_2560)
	);

	bfr G2553_bfr_after (
		.din(new_net_2560),
		.dout(G2553)
	);

	bfr new_net_2561_bfr_after (
		.din(_0358_),
		.dout(new_net_2561)
	);

	bfr new_net_2562_bfr_after (
		.din(new_net_2561),
		.dout(new_net_2562)
	);

	bfr new_net_2563_bfr_after (
		.din(new_net_2562),
		.dout(new_net_2563)
	);

	bfr new_net_2564_bfr_after (
		.din(new_net_2563),
		.dout(new_net_2564)
	);

	bfr new_net_2565_bfr_after (
		.din(new_net_2564),
		.dout(new_net_2565)
	);

	bfr new_net_2566_bfr_after (
		.din(new_net_2565),
		.dout(new_net_2566)
	);

	bfr new_net_2567_bfr_after (
		.din(new_net_2566),
		.dout(new_net_2567)
	);

	bfr new_net_2568_bfr_after (
		.din(new_net_2567),
		.dout(new_net_2568)
	);

	bfr new_net_899_bfr_after (
		.din(new_net_2568),
		.dout(new_net_899)
	);

	bfr new_net_2569_bfr_after (
		.din(G27),
		.dout(new_net_2569)
	);

	bfr new_net_873_bfr_after (
		.din(new_net_2569),
		.dout(new_net_873)
	);

	bfr new_net_2570_bfr_after (
		.din(G91),
		.dout(new_net_2570)
	);

	bfr new_net_2571_bfr_after (
		.din(new_net_2570),
		.dout(new_net_2571)
	);

	bfr new_net_2572_bfr_after (
		.din(new_net_2571),
		.dout(new_net_2572)
	);

	bfr new_net_826_bfr_after (
		.din(new_net_2572),
		.dout(new_net_826)
	);

	bfr new_net_2573_bfr_after (
		.din(_0046_),
		.dout(new_net_2573)
	);

	bfr new_net_784_bfr_after (
		.din(new_net_2573),
		.dout(new_net_784)
	);

	bfr new_net_2574_bfr_after (
		.din(G10),
		.dout(new_net_2574)
	);

	bfr new_net_2575_bfr_after (
		.din(new_net_2574),
		.dout(new_net_2575)
	);

	bfr new_net_2576_bfr_after (
		.din(new_net_2575),
		.dout(new_net_2576)
	);

	bfr new_net_2577_bfr_after (
		.din(new_net_2576),
		.dout(new_net_2577)
	);

	bfr new_net_2578_bfr_after (
		.din(new_net_2577),
		.dout(new_net_2578)
	);

	bfr new_net_2579_bfr_after (
		.din(new_net_2578),
		.dout(new_net_2579)
	);

	bfr new_net_2580_bfr_after (
		.din(new_net_2579),
		.dout(new_net_2580)
	);

	bfr new_net_2581_bfr_after (
		.din(new_net_2580),
		.dout(new_net_2581)
	);

	bfr new_net_2582_bfr_after (
		.din(new_net_2581),
		.dout(new_net_2582)
	);

	bfr new_net_2583_bfr_after (
		.din(new_net_2582),
		.dout(new_net_2583)
	);

	bfr new_net_805_bfr_after (
		.din(new_net_2583),
		.dout(new_net_805)
	);

	bfr new_net_2584_bfr_after (
		.din(G45),
		.dout(new_net_2584)
	);

	bfr new_net_2585_bfr_after (
		.din(new_net_2584),
		.dout(new_net_2585)
	);

	bfr new_net_2586_bfr_after (
		.din(new_net_2585),
		.dout(new_net_2586)
	);

	bfr new_net_2587_bfr_after (
		.din(new_net_2586),
		.dout(new_net_2587)
	);

	bfr new_net_2588_bfr_after (
		.din(new_net_2587),
		.dout(new_net_2588)
	);

	bfr new_net_788_bfr_after (
		.din(new_net_2588),
		.dout(new_net_788)
	);

	bfr new_net_2589_bfr_after (
		.din(G107),
		.dout(new_net_2589)
	);

	bfr new_net_2590_bfr_after (
		.din(new_net_2589),
		.dout(new_net_2590)
	);

	bfr new_net_2591_bfr_after (
		.din(new_net_2590),
		.dout(new_net_2591)
	);

	bfr new_net_809_bfr_after (
		.din(new_net_2591),
		.dout(new_net_809)
	);

	bfr new_net_2592_bfr_after (
		.din(G79),
		.dout(new_net_2592)
	);

	bfr new_net_2593_bfr_after (
		.din(new_net_2592),
		.dout(new_net_2593)
	);

	bfr new_net_2594_bfr_after (
		.din(new_net_2593),
		.dout(new_net_2594)
	);

	bfr new_net_759_bfr_after (
		.din(new_net_2594),
		.dout(new_net_759)
	);

	bfr new_net_2595_bfr_after (
		.din(_0025_),
		.dout(new_net_2595)
	);

	bfr new_net_767_bfr_after (
		.din(new_net_2595),
		.dout(new_net_767)
	);

	bfr new_net_2596_bfr_after (
		.din(G69),
		.dout(new_net_2596)
	);

	bfr new_net_2597_bfr_after (
		.din(new_net_2596),
		.dout(new_net_2597)
	);

	bfr new_net_763_bfr_after (
		.din(new_net_2597),
		.dout(new_net_763)
	);

	bfr new_net_2598_bfr_after (
		.din(G65),
		.dout(new_net_2598)
	);

	bfr new_net_2599_bfr_after (
		.din(new_net_2598),
		.dout(new_net_2599)
	);

	bfr new_net_780_bfr_after (
		.din(new_net_2599),
		.dout(new_net_780)
	);

	bfr new_net_2600_bfr_after (
		.din(G59),
		.dout(new_net_2600)
	);

	bfr new_net_2601_bfr_after (
		.din(new_net_2600),
		.dout(new_net_2601)
	);

	bfr new_net_2602_bfr_after (
		.din(new_net_2601),
		.dout(new_net_2602)
	);

	bfr new_net_2603_bfr_after (
		.din(new_net_2602),
		.dout(new_net_2603)
	);

	bfr new_net_2604_bfr_after (
		.din(new_net_2603),
		.dout(new_net_2604)
	);

	bfr new_net_801_bfr_after (
		.din(new_net_2604),
		.dout(new_net_801)
	);

	bfr new_net_2605_bfr_after (
		.din(_0222_),
		.dout(new_net_2605)
	);

	bfr new_net_837_bfr_after (
		.din(new_net_2605),
		.dout(new_net_837)
	);

	bfr new_net_2606_bfr_after (
		.din(_0287_),
		.dout(new_net_2606)
	);

	bfr new_net_2607_bfr_after (
		.din(new_net_2606),
		.dout(new_net_2607)
	);

	bfr new_net_2608_bfr_after (
		.din(new_net_2607),
		.dout(new_net_2608)
	);

	bfr new_net_2609_bfr_after (
		.din(new_net_2608),
		.dout(new_net_2609)
	);

	bfr new_net_2610_bfr_after (
		.din(new_net_2609),
		.dout(new_net_2610)
	);

	bfr new_net_2611_bfr_after (
		.din(new_net_2610),
		.dout(new_net_2611)
	);

	bfr new_net_2612_bfr_after (
		.din(new_net_2611),
		.dout(new_net_2612)
	);

	bfr new_net_2613_bfr_after (
		.din(new_net_2612),
		.dout(new_net_2613)
	);

	bfr new_net_864_bfr_after (
		.din(new_net_2613),
		.dout(new_net_864)
	);

	bfr new_net_859_bfr_after (
		.din(_0275_),
		.dout(new_net_859)
	);

	bfr new_net_2614_bfr_after (
		.din(_0422_),
		.dout(new_net_2614)
	);

	bfr new_net_2615_bfr_after (
		.din(new_net_2614),
		.dout(new_net_2615)
	);

	bfr new_net_922_bfr_after (
		.din(new_net_2615),
		.dout(new_net_922)
	);

	bfr new_net_886_bfr_after (
		.din(_0296_),
		.dout(new_net_886)
	);

	bfr new_net_881_bfr_after (
		.din(_0316_),
		.dout(new_net_881)
	);

	bfr new_net_2616_bfr_after (
		.din(_0496_),
		.dout(new_net_2616)
	);

	bfr new_net_2617_bfr_after (
		.din(new_net_2616),
		.dout(new_net_2617)
	);

	bfr new_net_2618_bfr_after (
		.din(new_net_2617),
		.dout(new_net_2618)
	);

	bfr new_net_2619_bfr_after (
		.din(new_net_2618),
		.dout(new_net_2619)
	);

	bfr new_net_2620_bfr_after (
		.din(new_net_2619),
		.dout(new_net_2620)
	);

	bfr new_net_2621_bfr_after (
		.din(new_net_2620),
		.dout(new_net_2621)
	);

	bfr new_net_2622_bfr_after (
		.din(new_net_2621),
		.dout(new_net_2622)
	);

	bfr new_net_2623_bfr_after (
		.din(new_net_2622),
		.dout(new_net_2623)
	);

	bfr new_net_944_bfr_after (
		.din(new_net_2623),
		.dout(new_net_944)
	);

	bfr new_net_2624_bfr_after (
		.din(_0378_),
		.dout(new_net_2624)
	);

	bfr new_net_908_bfr_after (
		.din(new_net_2624),
		.dout(new_net_908)
	);

	bfr new_net_2625_bfr_after (
		.din(G9),
		.dout(new_net_2625)
	);

	bfr new_net_2626_bfr_after (
		.din(new_net_2625),
		.dout(new_net_2626)
	);

	bfr new_net_903_bfr_after (
		.din(new_net_2626),
		.dout(new_net_903)
	);

	bfr new_net_2627_bfr_after (
		.din(_0414_),
		.dout(new_net_2627)
	);

	bfr new_net_2628_bfr_after (
		.din(new_net_2627),
		.dout(new_net_2628)
	);

	bfr new_net_2629_bfr_after (
		.din(new_net_2628),
		.dout(new_net_2629)
	);

	bfr new_net_2630_bfr_after (
		.din(new_net_2629),
		.dout(new_net_2630)
	);

	bfr new_net_2631_bfr_after (
		.din(new_net_2630),
		.dout(new_net_2631)
	);

	bfr new_net_2632_bfr_after (
		.din(new_net_2631),
		.dout(new_net_2632)
	);

	bfr new_net_2633_bfr_after (
		.din(new_net_2632),
		.dout(new_net_2633)
	);

	bfr new_net_2634_bfr_after (
		.din(new_net_2633),
		.dout(new_net_2634)
	);

	bfr new_net_2635_bfr_after (
		.din(new_net_2634),
		.dout(new_net_2635)
	);

	bfr new_net_930_bfr_after (
		.din(new_net_2635),
		.dout(new_net_930)
	);

	bfr new_net_2636_bfr_after (
		.din(new_net_963),
		.dout(new_net_2636)
	);

	bfr new_net_2637_bfr_after (
		.din(new_net_2636),
		.dout(new_net_2637)
	);

	bfr new_net_2638_bfr_after (
		.din(new_net_2637),
		.dout(new_net_2638)
	);

	bfr new_net_2639_bfr_after (
		.din(new_net_2638),
		.dout(new_net_2639)
	);

	bfr new_net_2640_bfr_after (
		.din(new_net_2639),
		.dout(new_net_2640)
	);

	bfr new_net_2641_bfr_after (
		.din(new_net_2640),
		.dout(new_net_2641)
	);

	bfr new_net_2642_bfr_after (
		.din(new_net_2641),
		.dout(new_net_2642)
	);

	bfr new_net_2643_bfr_after (
		.din(new_net_2642),
		.dout(new_net_2643)
	);

	bfr new_net_2644_bfr_after (
		.din(new_net_2643),
		.dout(new_net_2644)
	);

	bfr new_net_2645_bfr_after (
		.din(new_net_2644),
		.dout(new_net_2645)
	);

	bfr new_net_2646_bfr_after (
		.din(new_net_2645),
		.dout(new_net_2646)
	);

	bfr new_net_2647_bfr_after (
		.din(new_net_2646),
		.dout(new_net_2647)
	);

	bfr new_net_2648_bfr_after (
		.din(new_net_2647),
		.dout(new_net_2648)
	);

	bfr new_net_2649_bfr_after (
		.din(new_net_2648),
		.dout(new_net_2649)
	);

	bfr new_net_2650_bfr_after (
		.din(new_net_2649),
		.dout(new_net_2650)
	);

	bfr new_net_2651_bfr_after (
		.din(new_net_2650),
		.dout(new_net_2651)
	);

	bfr G2580_bfr_after (
		.din(new_net_2651),
		.dout(G2580)
	);

	bfr new_net_2652_bfr_after (
		.din(G42),
		.dout(new_net_2652)
	);

	bfr new_net_2653_bfr_after (
		.din(new_net_2652),
		.dout(new_net_2653)
	);

	bfr new_net_2654_bfr_after (
		.din(new_net_2653),
		.dout(new_net_2654)
	);

	bfr new_net_2655_bfr_after (
		.din(new_net_2654),
		.dout(new_net_2655)
	);

	bfr new_net_2656_bfr_after (
		.din(new_net_2655),
		.dout(new_net_2656)
	);

	bfr new_net_841_bfr_after (
		.din(new_net_2656),
		.dout(new_net_841)
	);

	bfr new_net_2657_bfr_after (
		.din(G5),
		.dout(new_net_2657)
	);

	bfr new_net_868_bfr_after (
		.din(new_net_2657),
		.dout(new_net_868)
	);

	bfr new_net_2658_bfr_after (
		.din(new_net_952),
		.dout(new_net_2658)
	);

	bfr new_net_2659_bfr_after (
		.din(new_net_2658),
		.dout(new_net_2659)
	);

	bfr new_net_2660_bfr_after (
		.din(new_net_2659),
		.dout(new_net_2660)
	);

	bfr new_net_2661_bfr_after (
		.din(new_net_2660),
		.dout(new_net_2661)
	);

	bfr new_net_2662_bfr_after (
		.din(new_net_2661),
		.dout(new_net_2662)
	);

	bfr new_net_2663_bfr_after (
		.din(new_net_2662),
		.dout(new_net_2663)
	);

	bfr new_net_2664_bfr_after (
		.din(new_net_2663),
		.dout(new_net_2664)
	);

	bfr new_net_2665_bfr_after (
		.din(new_net_2664),
		.dout(new_net_2665)
	);

	bfr new_net_2666_bfr_after (
		.din(new_net_2665),
		.dout(new_net_2666)
	);

	bfr new_net_2667_bfr_after (
		.din(new_net_2666),
		.dout(new_net_2667)
	);

	bfr new_net_2668_bfr_after (
		.din(new_net_2667),
		.dout(new_net_2668)
	);

	bfr new_net_2669_bfr_after (
		.din(new_net_2668),
		.dout(new_net_2669)
	);

	bfr new_net_2670_bfr_after (
		.din(new_net_2669),
		.dout(new_net_2670)
	);

	bfr new_net_2671_bfr_after (
		.din(new_net_2670),
		.dout(new_net_2671)
	);

	bfr new_net_2672_bfr_after (
		.din(new_net_2671),
		.dout(new_net_2672)
	);

	bfr new_net_2673_bfr_after (
		.din(new_net_2672),
		.dout(new_net_2673)
	);

	bfr new_net_2674_bfr_after (
		.din(new_net_2673),
		.dout(new_net_2674)
	);

	bfr new_net_2675_bfr_after (
		.din(new_net_2674),
		.dout(new_net_2675)
	);

	bfr new_net_2676_bfr_after (
		.din(new_net_2675),
		.dout(new_net_2676)
	);

	bfr new_net_2677_bfr_after (
		.din(new_net_2676),
		.dout(new_net_2677)
	);

	bfr new_net_2678_bfr_after (
		.din(new_net_2677),
		.dout(new_net_2678)
	);

	bfr new_net_2679_bfr_after (
		.din(new_net_2678),
		.dout(new_net_2679)
	);

	bfr new_net_2680_bfr_after (
		.din(new_net_2679),
		.dout(new_net_2680)
	);

	bfr new_net_2681_bfr_after (
		.din(new_net_2680),
		.dout(new_net_2681)
	);

	bfr new_net_2682_bfr_after (
		.din(new_net_2681),
		.dout(new_net_2682)
	);

	bfr G2548_bfr_after (
		.din(new_net_2682),
		.dout(G2548)
	);

	bfr new_net_2683_bfr_after (
		.din(G13),
		.dout(new_net_2683)
	);

	bfr new_net_863_bfr_after (
		.din(new_net_2683),
		.dout(new_net_863)
	);

	bfr new_net_2684_bfr_after (
		.din(_0458_),
		.dout(new_net_2684)
	);

	bfr new_net_2685_bfr_after (
		.din(new_net_2684),
		.dout(new_net_2685)
	);

	bfr new_net_926_bfr_after (
		.din(new_net_2685),
		.dout(new_net_926)
	);

	bfr new_net_2686_bfr_after (
		.din(G33),
		.dout(new_net_2686)
	);

	bfr new_net_2687_bfr_after (
		.din(new_net_2686),
		.dout(new_net_2687)
	);

	bfr new_net_779_bfr_after (
		.din(new_net_2687),
		.dout(new_net_779)
	);

	bfr new_net_2688_bfr_after (
		.din(G48),
		.dout(new_net_2688)
	);

	bfr new_net_2689_bfr_after (
		.din(new_net_2688),
		.dout(new_net_2689)
	);

	bfr new_net_2690_bfr_after (
		.din(new_net_2689),
		.dout(new_net_2690)
	);

	bfr new_net_2691_bfr_after (
		.din(new_net_2690),
		.dout(new_net_2691)
	);

	bfr new_net_2692_bfr_after (
		.din(new_net_2691),
		.dout(new_net_2692)
	);

	bfr new_net_800_bfr_after (
		.din(new_net_2692),
		.dout(new_net_800)
	);

	bfr new_net_2693_bfr_after (
		.din(G108),
		.dout(new_net_2693)
	);

	bfr new_net_2694_bfr_after (
		.din(new_net_2693),
		.dout(new_net_2694)
	);

	bfr new_net_2695_bfr_after (
		.din(new_net_2694),
		.dout(new_net_2695)
	);

	bfr new_net_754_bfr_after (
		.din(new_net_2695),
		.dout(new_net_754)
	);

	bfr new_net_2696_bfr_after (
		.din(G109),
		.dout(new_net_2696)
	);

	bfr new_net_2697_bfr_after (
		.din(new_net_2696),
		.dout(new_net_2697)
	);

	bfr new_net_2698_bfr_after (
		.din(new_net_2697),
		.dout(new_net_2698)
	);

	bfr new_net_758_bfr_after (
		.din(new_net_2698),
		.dout(new_net_758)
	);

	bfr new_net_771_bfr_after (
		.din(_0032_),
		.dout(new_net_771)
	);

	bfr new_net_2699_bfr_after (
		.din(G71),
		.dout(new_net_2699)
	);

	bfr new_net_2700_bfr_after (
		.din(new_net_2699),
		.dout(new_net_2700)
	);

	bfr new_net_792_bfr_after (
		.din(new_net_2700),
		.dout(new_net_792)
	);

	bfr new_net_2701_bfr_after (
		.din(G113),
		.dout(new_net_2701)
	);

	bfr new_net_2702_bfr_after (
		.din(new_net_2701),
		.dout(new_net_2702)
	);

	bfr new_net_2703_bfr_after (
		.din(new_net_2702),
		.dout(new_net_2703)
	);

	bfr new_net_813_bfr_after (
		.din(new_net_2703),
		.dout(new_net_813)
	);

	bfr new_net_775_bfr_after (
		.din(_0036_),
		.dout(new_net_775)
	);

	bfr new_net_2704_bfr_after (
		.din(_0060_),
		.dout(new_net_2704)
	);

	bfr new_net_796_bfr_after (
		.din(new_net_2704),
		.dout(new_net_796)
	);

	bfr new_net_2705_bfr_after (
		.din(G112),
		.dout(new_net_2705)
	);

	bfr new_net_2706_bfr_after (
		.din(new_net_2705),
		.dout(new_net_2706)
	);

	bfr new_net_2707_bfr_after (
		.din(new_net_2706),
		.dout(new_net_2707)
	);

	bfr new_net_817_bfr_after (
		.din(new_net_2707),
		.dout(new_net_817)
	);

	bfr new_net_2708_bfr_after (
		.din(G41),
		.dout(new_net_2708)
	);

	bfr new_net_2709_bfr_after (
		.din(new_net_2708),
		.dout(new_net_2709)
	);

	bfr new_net_832_bfr_after (
		.din(new_net_2709),
		.dout(new_net_832)
	);

	bfr new_net_2710_bfr_after (
		.din(_0337_),
		.dout(new_net_2710)
	);

	bfr new_net_2711_bfr_after (
		.din(new_net_2710),
		.dout(new_net_2711)
	);

	bfr new_net_2712_bfr_after (
		.din(new_net_2711),
		.dout(new_net_2712)
	);

	bfr new_net_2713_bfr_after (
		.din(new_net_2712),
		.dout(new_net_2713)
	);

	bfr new_net_2714_bfr_after (
		.din(new_net_2713),
		.dout(new_net_2714)
	);

	bfr new_net_2715_bfr_after (
		.din(new_net_2714),
		.dout(new_net_2715)
	);

	bfr new_net_2716_bfr_after (
		.din(new_net_2715),
		.dout(new_net_2716)
	);

	bfr new_net_2717_bfr_after (
		.din(new_net_2716),
		.dout(new_net_2717)
	);

	bfr new_net_890_bfr_after (
		.din(new_net_2717),
		.dout(new_net_890)
	);

	bfr new_net_854_bfr_after (
		.din(G116),
		.dout(new_net_854)
	);

	bfr new_net_2718_bfr_after (
		.din(_0398_),
		.dout(new_net_2718)
	);

	bfr new_net_2719_bfr_after (
		.din(new_net_2718),
		.dout(new_net_2719)
	);

	bfr new_net_2720_bfr_after (
		.din(new_net_2719),
		.dout(new_net_2720)
	);

	bfr new_net_2721_bfr_after (
		.din(new_net_2720),
		.dout(new_net_2721)
	);

	bfr new_net_2722_bfr_after (
		.din(new_net_2721),
		.dout(new_net_2722)
	);

	bfr new_net_2723_bfr_after (
		.din(new_net_2722),
		.dout(new_net_2723)
	);

	bfr new_net_2724_bfr_after (
		.din(new_net_2723),
		.dout(new_net_2724)
	);

	bfr new_net_2725_bfr_after (
		.din(new_net_2724),
		.dout(new_net_2725)
	);

	bfr new_net_2726_bfr_after (
		.din(new_net_2725),
		.dout(new_net_2726)
	);

	bfr new_net_2727_bfr_after (
		.din(new_net_2726),
		.dout(new_net_2727)
	);

	bfr new_net_2728_bfr_after (
		.din(new_net_2727),
		.dout(new_net_2728)
	);

	bfr new_net_917_bfr_after (
		.din(new_net_2728),
		.dout(new_net_917)
	);

	bfr new_net_2729_bfr_after (
		.din(_0244_),
		.dout(new_net_2729)
	);

	bfr new_net_849_bfr_after (
		.din(new_net_2729),
		.dout(new_net_849)
	);

	bfr new_net_2730_bfr_after (
		.din(G17),
		.dout(new_net_2730)
	);

	bfr new_net_912_bfr_after (
		.din(new_net_2730),
		.dout(new_net_912)
	);

	bfr new_net_876_bfr_after (
		.din(_0311_),
		.dout(new_net_876)
	);

	bfr new_net_2731_bfr_after (
		.din(_0491_),
		.dout(new_net_2731)
	);

	bfr new_net_2732_bfr_after (
		.din(new_net_2731),
		.dout(new_net_2732)
	);

	bfr new_net_2733_bfr_after (
		.din(new_net_2732),
		.dout(new_net_2733)
	);

	bfr new_net_2734_bfr_after (
		.din(new_net_2733),
		.dout(new_net_2734)
	);

	bfr new_net_2735_bfr_after (
		.din(new_net_2734),
		.dout(new_net_2735)
	);

	bfr new_net_2736_bfr_after (
		.din(new_net_2735),
		.dout(new_net_2736)
	);

	bfr new_net_2737_bfr_after (
		.din(new_net_2736),
		.dout(new_net_2737)
	);

	bfr new_net_2738_bfr_after (
		.din(new_net_2737),
		.dout(new_net_2738)
	);

	bfr new_net_939_bfr_after (
		.din(new_net_2738),
		.dout(new_net_939)
	);

	bfr new_net_934_bfr_after (
		.din(_0476_),
		.dout(new_net_934)
	);

	bfr new_net_2739_bfr_after (
		.din(new_net_957),
		.dout(new_net_2739)
	);

	bfr new_net_2740_bfr_after (
		.din(new_net_2739),
		.dout(new_net_2740)
	);

	bfr new_net_2741_bfr_after (
		.din(new_net_2740),
		.dout(new_net_2741)
	);

	bfr new_net_2742_bfr_after (
		.din(new_net_2741),
		.dout(new_net_2742)
	);

	bfr new_net_2743_bfr_after (
		.din(new_net_2742),
		.dout(new_net_2743)
	);

	bfr new_net_2744_bfr_after (
		.din(new_net_2743),
		.dout(new_net_2744)
	);

	bfr new_net_2745_bfr_after (
		.din(new_net_2744),
		.dout(new_net_2745)
	);

	bfr new_net_2746_bfr_after (
		.din(new_net_2745),
		.dout(new_net_2746)
	);

	bfr new_net_2747_bfr_after (
		.din(new_net_2746),
		.dout(new_net_2747)
	);

	bfr new_net_2748_bfr_after (
		.din(new_net_2747),
		.dout(new_net_2748)
	);

	bfr new_net_2749_bfr_after (
		.din(new_net_2748),
		.dout(new_net_2749)
	);

	bfr new_net_2750_bfr_after (
		.din(new_net_2749),
		.dout(new_net_2750)
	);

	bfr new_net_2751_bfr_after (
		.din(new_net_2750),
		.dout(new_net_2751)
	);

	bfr new_net_2752_bfr_after (
		.din(new_net_2751),
		.dout(new_net_2752)
	);

	bfr new_net_2753_bfr_after (
		.din(new_net_2752),
		.dout(new_net_2753)
	);

	bfr new_net_2754_bfr_after (
		.din(new_net_2753),
		.dout(new_net_2754)
	);

	bfr new_net_2755_bfr_after (
		.din(new_net_2754),
		.dout(new_net_2755)
	);

	bfr new_net_2756_bfr_after (
		.din(new_net_2755),
		.dout(new_net_2756)
	);

	bfr new_net_2757_bfr_after (
		.din(new_net_2756),
		.dout(new_net_2757)
	);

	bfr new_net_2758_bfr_after (
		.din(new_net_2757),
		.dout(new_net_2758)
	);

	bfr new_net_2759_bfr_after (
		.din(new_net_2758),
		.dout(new_net_2759)
	);

	bfr new_net_2760_bfr_after (
		.din(new_net_2759),
		.dout(new_net_2760)
	);

	bfr new_net_2761_bfr_after (
		.din(new_net_2760),
		.dout(new_net_2761)
	);

	bfr new_net_2762_bfr_after (
		.din(new_net_2761),
		.dout(new_net_2762)
	);

	bfr G2552_bfr_after (
		.din(new_net_2762),
		.dout(G2552)
	);

	bfr new_net_2763_bfr_after (
		.din(G18),
		.dout(new_net_2763)
	);

	bfr new_net_898_bfr_after (
		.din(new_net_2763),
		.dout(new_net_898)
	);

	bfr new_net_2764_bfr_after (
		.din(_0304_),
		.dout(new_net_2764)
	);

	bfr new_net_872_bfr_after (
		.din(new_net_2764),
		.dout(new_net_872)
	);

	bfr new_net_2765_bfr_after (
		.din(G62),
		.dout(new_net_2765)
	);

	bfr new_net_2766_bfr_after (
		.din(new_net_2765),
		.dout(new_net_2766)
	);

	bfr new_net_2767_bfr_after (
		.din(new_net_2766),
		.dout(new_net_2767)
	);

	bfr new_net_2768_bfr_after (
		.din(new_net_2767),
		.dout(new_net_2768)
	);

	bfr new_net_2769_bfr_after (
		.din(new_net_2768),
		.dout(new_net_2769)
	);

	bfr new_net_836_bfr_after (
		.din(new_net_2769),
		.dout(new_net_836)
	);

	bfr new_net_2770_bfr_after (
		.din(_0336_),
		.dout(new_net_2770)
	);

	bfr new_net_2771_bfr_after (
		.din(new_net_2770),
		.dout(new_net_2771)
	);

	bfr new_net_2772_bfr_after (
		.din(new_net_2771),
		.dout(new_net_2772)
	);

	bfr new_net_894_bfr_after (
		.din(new_net_2772),
		.dout(new_net_894)
	);

	bfr new_net_2773_bfr_after (
		.din(G54),
		.dout(new_net_2773)
	);

	bfr new_net_2774_bfr_after (
		.din(new_net_2773),
		.dout(new_net_2774)
	);

	bfr new_net_2775_bfr_after (
		.din(new_net_2774),
		.dout(new_net_2775)
	);

	bfr new_net_2776_bfr_after (
		.din(new_net_2775),
		.dout(new_net_2776)
	);

	bfr new_net_2777_bfr_after (
		.din(new_net_2776),
		.dout(new_net_2777)
	);

	bfr new_net_783_bfr_after (
		.din(new_net_2777),
		.dout(new_net_783)
	);

	bfr new_net_804_bfr_after (
		.din(_0101_),
		.dout(new_net_804)
	);

	bfr new_net_2778_bfr_after (
		.din(G111),
		.dout(new_net_2778)
	);

	bfr new_net_2779_bfr_after (
		.din(new_net_2778),
		.dout(new_net_2779)
	);

	bfr new_net_2780_bfr_after (
		.din(new_net_2779),
		.dout(new_net_2780)
	);

	bfr new_net_825_bfr_after (
		.din(new_net_2780),
		.dout(new_net_825)
	);

	bfr new_net_787_bfr_after (
		.din(_0050_),
		.dout(new_net_787)
	);

	bfr new_net_2781_bfr_after (
		.din(G97),
		.dout(new_net_2781)
	);

	bfr new_net_2782_bfr_after (
		.din(new_net_2781),
		.dout(new_net_2782)
	);

	bfr new_net_2783_bfr_after (
		.din(new_net_2782),
		.dout(new_net_2783)
	);

	bfr new_net_808_bfr_after (
		.din(new_net_2783),
		.dout(new_net_808)
	);

	bfr new_net_2784_bfr_after (
		.din(G37),
		.dout(new_net_2784)
	);

	bfr new_net_2785_bfr_after (
		.din(new_net_2784),
		.dout(new_net_2785)
	);

	bfr new_net_762_bfr_after (
		.din(new_net_2785),
		.dout(new_net_762)
	);

	bfr new_net_2786_bfr_after (
		.din(G58),
		.dout(new_net_2786)
	);

	bfr new_net_2787_bfr_after (
		.din(new_net_2786),
		.dout(new_net_2787)
	);

	bfr new_net_2788_bfr_after (
		.din(new_net_2787),
		.dout(new_net_2788)
	);

	bfr new_net_2789_bfr_after (
		.din(new_net_2788),
		.dout(new_net_2789)
	);

	bfr new_net_2790_bfr_after (
		.din(new_net_2789),
		.dout(new_net_2790)
	);

	bfr new_net_766_bfr_after (
		.din(new_net_2790),
		.dout(new_net_766)
	);

	bfr new_net_2791_bfr_after (
		.din(G95),
		.dout(new_net_2791)
	);

	bfr new_net_2792_bfr_after (
		.din(new_net_2791),
		.dout(new_net_2792)
	);

	bfr new_net_2793_bfr_after (
		.din(new_net_2792),
		.dout(new_net_2793)
	);

	bfr new_net_829_bfr_after (
		.din(new_net_2793),
		.dout(new_net_829)
	);

	bfr new_net_846_bfr_after (
		.din(_0241_),
		.dout(new_net_846)
	);

	bfr new_net_850_bfr_after (
		.din(_0258_),
		.dout(new_net_850)
	);

	bfr new_net_858_bfr_after (
		.din(_0274_),
		.dout(new_net_858)
	);

	bfr new_net_2794_bfr_after (
		.din(_0426_),
		.dout(new_net_2794)
	);

	bfr new_net_921_bfr_after (
		.din(new_net_2794),
		.dout(new_net_921)
	);

	bfr new_net_885_bfr_after (
		.din(_0312_),
		.dout(new_net_885)
	);

	bfr new_net_2795_bfr_after (
		.din(_0317_),
		.dout(new_net_2795)
	);

	bfr new_net_2796_bfr_after (
		.din(new_net_2795),
		.dout(new_net_2796)
	);

	bfr new_net_2797_bfr_after (
		.din(new_net_2796),
		.dout(new_net_2797)
	);

	bfr new_net_2798_bfr_after (
		.din(new_net_2797),
		.dout(new_net_2798)
	);

	bfr new_net_2799_bfr_after (
		.din(new_net_2798),
		.dout(new_net_2799)
	);

	bfr new_net_2800_bfr_after (
		.din(new_net_2799),
		.dout(new_net_2800)
	);

	bfr new_net_2801_bfr_after (
		.din(new_net_2800),
		.dout(new_net_2801)
	);

	bfr new_net_2802_bfr_after (
		.din(new_net_2801),
		.dout(new_net_2802)
	);

	bfr new_net_880_bfr_after (
		.din(new_net_2802),
		.dout(new_net_880)
	);

	bfr new_net_943_bfr_after (
		.din(G74),
		.dout(new_net_943)
	);

	bfr new_net_2803_bfr_after (
		.din(G40),
		.dout(new_net_2803)
	);

	bfr new_net_2804_bfr_after (
		.din(new_net_2803),
		.dout(new_net_2804)
	);

	bfr new_net_844_bfr_after (
		.din(new_net_2804),
		.dout(new_net_844)
	);

	bfr new_net_2805_bfr_after (
		.din(G22),
		.dout(new_net_2805)
	);

	bfr new_net_902_bfr_after (
		.din(new_net_2805),
		.dout(new_net_902)
	);

endmodule