module apc64bits(in, out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _apc32_1_apc16_1_adder1_lv1_a ;
  wire _apc32_1_apc16_1_adder1_lv1_b ;
  wire _apc32_1_apc16_1_adder1_lv1_cin ;
  wire _apc32_1_apc16_1_adder1_lv1_cout ;
  wire _apc32_1_apc16_1_adder1_lv1_d ;
  wire _apc32_1_apc16_1_adder1_lv1_m3_d ;
  wire _apc32_1_apc16_1_adder1_lv2_b ;
  wire _apc32_1_apc16_1_adder1_lv2_cin ;
  wire _apc32_1_apc16_1_adder1_lv2_cout ;
  wire _apc32_1_apc16_1_adder1_lv2_d ;
  wire _apc32_1_apc16_1_adder1_lv2_m3_d ;
  wire _apc32_1_apc16_1_adder2_lv1_a ;
  wire _apc32_1_apc16_1_adder2_lv1_b ;
  wire _apc32_1_apc16_1_adder2_lv1_cin ;
  wire _apc32_1_apc16_1_adder2_lv1_d ;
  wire _apc32_1_apc16_1_adder2_lv1_m3_d ;
  wire _apc32_1_apc16_1_adder2_lv2_cin ;
  wire _apc32_1_apc16_1_adder2_lv2_d ;
  wire _apc32_1_apc16_1_adder2_lv2_m3_d ;
  wire _apc32_1_apc16_1_half1_a ;
  wire _apc32_1_apc16_1_half1_cout ;
  wire _apc32_1_apc16_1_half1_s ;
  wire _apc32_1_apc16_1_half2_cout ;
  wire _apc32_1_apc16_1_half2_s ;
  wire _apc32_1_apc16_1_half3_cout ;
  wire _apc32_1_apc16_1_half3_s ;
  wire _apc32_1_apc16_2_adder1_lv1_a ;
  wire _apc32_1_apc16_2_adder1_lv1_b ;
  wire _apc32_1_apc16_2_adder1_lv1_cin ;
  wire _apc32_1_apc16_2_adder1_lv1_cout ;
  wire _apc32_1_apc16_2_adder1_lv1_d ;
  wire _apc32_1_apc16_2_adder1_lv1_m3_d ;
  wire _apc32_1_apc16_2_adder1_lv2_b ;
  wire _apc32_1_apc16_2_adder1_lv2_cin ;
  wire _apc32_1_apc16_2_adder1_lv2_cout ;
  wire _apc32_1_apc16_2_adder1_lv2_d ;
  wire _apc32_1_apc16_2_adder1_lv2_m3_d ;
  wire _apc32_1_apc16_2_adder2_lv1_a ;
  wire _apc32_1_apc16_2_adder2_lv1_b ;
  wire _apc32_1_apc16_2_adder2_lv1_cin ;
  wire _apc32_1_apc16_2_adder2_lv1_d ;
  wire _apc32_1_apc16_2_adder2_lv1_m3_d ;
  wire _apc32_1_apc16_2_adder2_lv2_cin ;
  wire _apc32_1_apc16_2_adder2_lv2_d ;
  wire _apc32_1_apc16_2_adder2_lv2_m3_d ;
  wire _apc32_1_apc16_2_half1_a ;
  wire _apc32_1_apc16_2_half1_cout ;
  wire _apc32_1_apc16_2_half1_s ;
  wire _apc32_1_apc16_2_half2_cout ;
  wire _apc32_1_apc16_2_half2_s ;
  wire _apc32_1_apc16_2_half3_cout ;
  wire _apc32_1_apc16_2_half3_s ;
  wire _apc32_1_out_0_;
  wire _apc32_1_out_1_;
  wire _apc32_1_out_2_;
  wire _apc32_1_out_3_;
  wire _apc32_1_out_4_;
  wire _apc32_1_out_5_;
  wire _apc32_2_apc16_1_adder1_lv1_a ;
  wire _apc32_2_apc16_1_adder1_lv1_b ;
  wire _apc32_2_apc16_1_adder1_lv1_cin ;
  wire _apc32_2_apc16_1_adder1_lv1_cout ;
  wire _apc32_2_apc16_1_adder1_lv1_d ;
  wire _apc32_2_apc16_1_adder1_lv1_m3_d ;
  wire _apc32_2_apc16_1_adder1_lv2_b ;
  wire _apc32_2_apc16_1_adder1_lv2_cin ;
  wire _apc32_2_apc16_1_adder1_lv2_cout ;
  wire _apc32_2_apc16_1_adder1_lv2_d ;
  wire _apc32_2_apc16_1_adder1_lv2_m3_d ;
  wire _apc32_2_apc16_1_adder2_lv1_a ;
  wire _apc32_2_apc16_1_adder2_lv1_b ;
  wire _apc32_2_apc16_1_adder2_lv1_cin ;
  wire _apc32_2_apc16_1_adder2_lv1_d ;
  wire _apc32_2_apc16_1_adder2_lv1_m3_d ;
  wire _apc32_2_apc16_1_adder2_lv2_cin ;
  wire _apc32_2_apc16_1_adder2_lv2_d ;
  wire _apc32_2_apc16_1_adder2_lv2_m3_d ;
  wire _apc32_2_apc16_1_half1_a ;
  wire _apc32_2_apc16_1_half1_cout ;
  wire _apc32_2_apc16_1_half1_s ;
  wire _apc32_2_apc16_1_half2_cout ;
  wire _apc32_2_apc16_1_half2_s ;
  wire _apc32_2_apc16_1_half3_cout ;
  wire _apc32_2_apc16_1_half3_s ;
  wire _apc32_2_apc16_2_adder1_lv1_a ;
  wire _apc32_2_apc16_2_adder1_lv1_b ;
  wire _apc32_2_apc16_2_adder1_lv1_cin ;
  wire _apc32_2_apc16_2_adder1_lv1_cout ;
  wire _apc32_2_apc16_2_adder1_lv1_d ;
  wire _apc32_2_apc16_2_adder1_lv1_m3_d ;
  wire _apc32_2_apc16_2_adder1_lv2_b ;
  wire _apc32_2_apc16_2_adder1_lv2_cin ;
  wire _apc32_2_apc16_2_adder1_lv2_cout ;
  wire _apc32_2_apc16_2_adder1_lv2_d ;
  wire _apc32_2_apc16_2_adder1_lv2_m3_d ;
  wire _apc32_2_apc16_2_adder2_lv1_a ;
  wire _apc32_2_apc16_2_adder2_lv1_b ;
  wire _apc32_2_apc16_2_adder2_lv1_cin ;
  wire _apc32_2_apc16_2_adder2_lv1_d ;
  wire _apc32_2_apc16_2_adder2_lv1_m3_d ;
  wire _apc32_2_apc16_2_adder2_lv2_cin ;
  wire _apc32_2_apc16_2_adder2_lv2_d ;
  wire _apc32_2_apc16_2_adder2_lv2_m3_d ;
  wire _apc32_2_apc16_2_half1_a ;
  wire _apc32_2_apc16_2_half1_cout ;
  wire _apc32_2_apc16_2_half1_s ;
  wire _apc32_2_apc16_2_half2_cout ;
  wire _apc32_2_apc16_2_half2_s ;
  wire _apc32_2_apc16_2_half3_cout ;
  wire _apc32_2_apc16_2_half3_s ;
  wire _apc32_2_out_0_;
  wire _apc32_2_out_1_;
  wire _apc32_2_out_2_;
  wire _apc32_2_out_3_;
  wire _apc32_2_out_4_;
  wire _apc32_2_out_5_;
  input in_0_;
  input in_1_;
  input in_2_;
  input in_3_;
  input in_4_;
  input in_5_;
  input in_6_;
  input in_7_;
  input in_8_;
  input in_9_;
  input in_10_;
  input in_11_;
  input in_12_;
  input in_13_;
  input in_14_;
  input in_15_;
  input in_16_;
  input in_17_;
  input in_18_;
  input in_19_;
  input in_20_;
  input in_21_;
  input in_22_;
  input in_23_;
  input in_24_;
  input in_25_;
  input in_26_;
  input in_27_;
  input in_28_;
  input in_29_;
  input in_30_;
  input in_31_;
  input in_32_;
  input in_33_;
  input in_34_;
  input in_35_;
  input in_36_;
  input in_37_;
  input in_38_;
  input in_39_;
  input in_40_;
  input in_41_;
  input in_42_;
  input in_43_;
  input in_44_;
  input in_45_;
  input in_46_;
  input in_47_;
  input in_48_;
  input in_49_;
  input in_50_;
  input in_51_;
  input in_52_;
  input in_53_;
  input in_54_;
  input in_55_;
  input in_56_;
  input in_57_;
  input in_58_;
  input in_59_;
  input in_60_;
  input in_61_;
  input in_62_;
  input in_63_;
  output out_0_;
  output out_1_;
  output out_2_;
  output out_3_;
  output out_4_;
  output out_5_;
  output out_6_;
  or_ii _093_ (
    .a(_apc32_2_out_0_),
    .b(_apc32_1_out_0_),
    .c(_000_)
  );
  or_ii _094_ (
    .a(_apc32_2_out_1_),
    .b(_apc32_1_out_1_),
    .c(_001_)
  );
  and_ii _095_ (
    .a(_apc32_2_out_1_),
    .b(_apc32_1_out_1_),
    .c(_002_)
  );
  and_bi _096_ (
    .a(_001_),
    .b(_002_),
    .c(_003_)
  );
  or_bi _097_ (
    .a(_000_),
    .b(_003_),
    .c(_004_)
  );
  and_bi _098_ (
    .a(_000_),
    .b(_003_),
    .c(_005_)
  );
  and_bi _099_ (
    .a(_004_),
    .b(_005_),
    .c(out_1_)
  );
  maj_bii _100_ (
    .a(_000_),
    .b(_apc32_2_out_1_),
    .c(_apc32_1_out_1_),
    .d(_006_)
  );
  or_ii _101_ (
    .a(_apc32_2_out_2_),
    .b(_apc32_1_out_2_),
    .c(_007_)
  );
  and_ii _102_ (
    .a(_apc32_2_out_2_),
    .b(_apc32_1_out_2_),
    .c(_008_)
  );
  and_bi _103_ (
    .a(_007_),
    .b(_008_),
    .c(_009_)
  );
  or_bi _104_ (
    .a(_006_),
    .b(_009_),
    .c(_010_)
  );
  and_bi _105_ (
    .a(_006_),
    .b(_009_),
    .c(_011_)
  );
  and_bi _106_ (
    .a(_010_),
    .b(_011_),
    .c(out_2_)
  );
  maj_bii _107_ (
    .a(_006_),
    .b(_apc32_2_out_2_),
    .c(_apc32_1_out_2_),
    .d(_012_)
  );
  or_ii _108_ (
    .a(_apc32_2_out_3_),
    .b(_apc32_1_out_3_),
    .c(_013_)
  );
  and_ii _109_ (
    .a(_apc32_2_out_3_),
    .b(_apc32_1_out_3_),
    .c(_014_)
  );
  and_bi _110_ (
    .a(_013_),
    .b(_014_),
    .c(_015_)
  );
  or_bi _111_ (
    .a(_012_),
    .b(_015_),
    .c(_016_)
  );
  and_bi _112_ (
    .a(_012_),
    .b(_015_),
    .c(_017_)
  );
  and_bi _113_ (
    .a(_016_),
    .b(_017_),
    .c(out_3_)
  );
  maj_bii _114_ (
    .a(_012_),
    .b(_apc32_2_out_3_),
    .c(_apc32_1_out_3_),
    .d(_018_)
  );
  or_ii _115_ (
    .a(_apc32_2_out_4_),
    .b(_apc32_1_out_4_),
    .c(_019_)
  );
  and_ii _116_ (
    .a(_apc32_2_out_4_),
    .b(_apc32_1_out_4_),
    .c(_020_)
  );
  and_bi _117_ (
    .a(_019_),
    .b(_020_),
    .c(_021_)
  );
  or_bi _118_ (
    .a(_018_),
    .b(_021_),
    .c(_022_)
  );
  and_bi _119_ (
    .a(_018_),
    .b(_021_),
    .c(_023_)
  );
  and_bi _120_ (
    .a(_022_),
    .b(_023_),
    .c(out_4_)
  );
  maj_bii _121_ (
    .a(_018_),
    .b(_apc32_2_out_4_),
    .c(_apc32_1_out_4_),
    .d(_024_)
  );
  or_ii _122_ (
    .a(_apc32_2_out_5_),
    .b(_apc32_1_out_5_),
    .c(_025_)
  );
  and_ii _123_ (
    .a(_apc32_2_out_5_),
    .b(_apc32_1_out_5_),
    .c(_026_)
  );
  and_bi _124_ (
    .a(_025_),
    .b(_026_),
    .c(_027_)
  );
  or_bi _125_ (
    .a(_024_),
    .b(_027_),
    .c(_028_)
  );
  and_bi _126_ (
    .a(_024_),
    .b(_027_),
    .c(_029_)
  );
  and_bi _127_ (
    .a(_028_),
    .b(_029_),
    .c(out_5_)
  );
  maj_bbi _128_ (
    .a(_apc32_2_out_5_),
    .b(_apc32_1_out_5_),
    .c(_024_),
    .d(out_6_)
  );
  and_ii _129_ (
    .a(_apc32_2_out_0_),
    .b(_apc32_1_out_0_),
    .c(_030_)
  );
  and_bi _130_ (
    .a(_000_),
    .b(_030_),
    .c(out_0_)
  );
  or_ii _131_ (
    .a(1'b0),
    .b(1'b0),
    .c(_031_)
  );
  or_ii _132_ (
    .a(_apc32_1_apc16_2_half1_s ),
    .b(_apc32_1_apc16_1_half1_s ),
    .c(_032_)
  );
  and_ii _133_ (
    .a(_apc32_1_apc16_2_half1_s ),
    .b(_apc32_1_apc16_1_half1_s ),
    .c(_033_)
  );
  and_bi _134_ (
    .a(_032_),
    .b(_033_),
    .c(_034_)
  );
  or_bi _135_ (
    .a(_031_),
    .b(_034_),
    .c(_035_)
  );
  and_bi _136_ (
    .a(_031_),
    .b(_034_),
    .c(_036_)
  );
  and_bi _137_ (
    .a(_035_),
    .b(_036_),
    .c(_apc32_1_out_1_)
  );
  maj_bii _138_ (
    .a(_031_),
    .b(_apc32_1_apc16_2_half1_s ),
    .c(_apc32_1_apc16_1_half1_s ),
    .d(_037_)
  );
  or_ii _139_ (
    .a(_apc32_1_apc16_2_half2_s ),
    .b(_apc32_1_apc16_1_half2_s ),
    .c(_038_)
  );
  and_ii _140_ (
    .a(_apc32_1_apc16_2_half2_s ),
    .b(_apc32_1_apc16_1_half2_s ),
    .c(_039_)
  );
  and_bi _141_ (
    .a(_038_),
    .b(_039_),
    .c(_040_)
  );
  or_bi _142_ (
    .a(_037_),
    .b(_040_),
    .c(_041_)
  );
  and_bi _143_ (
    .a(_037_),
    .b(_040_),
    .c(_042_)
  );
  and_bi _144_ (
    .a(_041_),
    .b(_042_),
    .c(_apc32_1_out_2_)
  );
  maj_bii _145_ (
    .a(_037_),
    .b(_apc32_1_apc16_2_half2_s ),
    .c(_apc32_1_apc16_1_half2_s ),
    .d(_043_)
  );
  or_ii _146_ (
    .a(_apc32_1_apc16_2_half3_s ),
    .b(_apc32_1_apc16_1_half3_s ),
    .c(_044_)
  );
  and_ii _147_ (
    .a(_apc32_1_apc16_2_half3_s ),
    .b(_apc32_1_apc16_1_half3_s ),
    .c(_045_)
  );
  and_bi _148_ (
    .a(_044_),
    .b(_045_),
    .c(_046_)
  );
  or_bi _149_ (
    .a(_043_),
    .b(_046_),
    .c(_047_)
  );
  and_bi _150_ (
    .a(_043_),
    .b(_046_),
    .c(_048_)
  );
  and_bi _151_ (
    .a(_047_),
    .b(_048_),
    .c(_apc32_1_out_3_)
  );
  maj_bii _152_ (
    .a(_043_),
    .b(_apc32_1_apc16_2_half3_s ),
    .c(_apc32_1_apc16_1_half3_s ),
    .d(_049_)
  );
  or_ii _153_ (
    .a(_apc32_1_apc16_2_half3_cout ),
    .b(_apc32_1_apc16_1_half3_cout ),
    .c(_050_)
  );
  and_ii _154_ (
    .a(_apc32_1_apc16_2_half3_cout ),
    .b(_apc32_1_apc16_1_half3_cout ),
    .c(_051_)
  );
  and_bi _155_ (
    .a(_050_),
    .b(_051_),
    .c(_052_)
  );
  or_bi _156_ (
    .a(_049_),
    .b(_052_),
    .c(_053_)
  );
  and_bi _157_ (
    .a(_049_),
    .b(_052_),
    .c(_054_)
  );
  and_bi _158_ (
    .a(_053_),
    .b(_054_),
    .c(_apc32_1_out_4_)
  );
  and_ii _159_ (
    .a(1'b0),
    .b(1'b0),
    .c(_055_)
  );
  and_bi _160_ (
    .a(_031_),
    .b(_055_),
    .c(_apc32_1_out_0_)
  );
  maj_bbi _161_ (
    .a(_apc32_1_apc16_2_half3_cout ),
    .b(_apc32_1_apc16_1_half3_cout ),
    .c(_049_),
    .d(_apc32_1_out_5_)
  );
  or_bb _162_ (
    .a(in_49_),
    .b(in_48_),
    .c(_apc32_1_apc16_1_adder1_lv1_a )
  );
  and_bb _163_ (
    .a(in_51_),
    .b(in_50_),
    .c(_apc32_1_apc16_1_adder1_lv1_b )
  );
  or_bb _164_ (
    .a(in_53_),
    .b(in_52_),
    .c(_apc32_1_apc16_1_adder1_lv1_cin )
  );
  and_bb _165_ (
    .a(in_55_),
    .b(in_54_),
    .c(_apc32_1_apc16_1_adder2_lv1_a )
  );
  or_bb _166_ (
    .a(in_57_),
    .b(in_56_),
    .c(_apc32_1_apc16_1_adder2_lv1_b )
  );
  and_bb _167_ (
    .a(in_59_),
    .b(in_58_),
    .c(_apc32_1_apc16_1_adder2_lv1_cin )
  );
  or_bb _168_ (
    .a(in_61_),
    .b(in_60_),
    .c(_apc32_1_apc16_1_adder2_lv2_cin )
  );
  and_bb _169_ (
    .a(in_63_),
    .b(in_62_),
    .c(_apc32_1_apc16_1_half1_a )
  );
  maj_bbb _170_ (
    .a(_apc32_1_apc16_1_adder1_lv1_cin ),
    .b(_apc32_1_apc16_1_adder1_lv1_b ),
    .c(_apc32_1_apc16_1_adder1_lv1_a ),
    .d(_apc32_1_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _171_ (
    .a(_apc32_1_apc16_1_adder1_lv1_b ),
    .b(_apc32_1_apc16_1_adder1_lv1_a ),
    .c(_apc32_1_apc16_1_adder1_lv1_cin ),
    .d(_apc32_1_apc16_1_adder1_lv1_d )
  );
  maj_bbi _172_ (
    .a(_apc32_1_apc16_1_adder1_lv1_d ),
    .b(_apc32_1_apc16_1_adder1_lv1_cin ),
    .c(_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc32_1_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _173_ (
    .a(_apc32_1_apc16_1_adder1_lv2_cin ),
    .b(_apc32_1_apc16_1_adder1_lv2_b ),
    .c(_apc32_1_apc16_1_adder1_lv1_cout ),
    .d(_apc32_1_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _174_ (
    .a(_apc32_1_apc16_1_adder1_lv2_b ),
    .b(_apc32_1_apc16_1_adder1_lv1_cout ),
    .c(_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc32_1_apc16_1_adder1_lv2_d )
  );
  maj_bbi _175_ (
    .a(_apc32_1_apc16_1_adder1_lv2_d ),
    .b(_apc32_1_apc16_1_adder1_lv2_cin ),
    .c(_apc32_1_apc16_1_adder1_lv2_cout ),
    .d(_apc32_1_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _176_ (
    .a(_apc32_1_apc16_1_adder2_lv1_cin ),
    .b(_apc32_1_apc16_1_adder2_lv1_b ),
    .c(_apc32_1_apc16_1_adder2_lv1_a ),
    .d(_apc32_1_apc16_1_adder1_lv2_b )
  );
  maj_bbi _177_ (
    .a(_apc32_1_apc16_1_adder2_lv1_b ),
    .b(_apc32_1_apc16_1_adder2_lv1_a ),
    .c(_apc32_1_apc16_1_adder2_lv1_cin ),
    .d(_apc32_1_apc16_1_adder2_lv1_d )
  );
  maj_bbi _178_ (
    .a(_apc32_1_apc16_1_adder2_lv1_d ),
    .b(_apc32_1_apc16_1_adder2_lv1_cin ),
    .c(_apc32_1_apc16_1_adder1_lv2_b ),
    .d(_apc32_1_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _179_ (
    .a(_apc32_1_apc16_1_adder2_lv2_cin ),
    .b(_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .c(_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .d(_apc32_1_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _180_ (
    .a(_apc32_1_apc16_1_adder2_lv1_m3_d ),
    .b(_apc32_1_apc16_1_adder1_lv1_m3_d ),
    .c(_apc32_1_apc16_1_adder2_lv2_cin ),
    .d(_apc32_1_apc16_1_adder2_lv2_d )
  );
  maj_bbi _181_ (
    .a(_apc32_1_apc16_1_adder2_lv2_d ),
    .b(_apc32_1_apc16_1_adder2_lv2_cin ),
    .c(_apc32_1_apc16_1_adder1_lv2_cin ),
    .d(_apc32_1_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _182_ (
    .a(_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc32_1_apc16_1_half1_a ),
    .c(_apc32_1_apc16_1_half1_cout )
  );
  or_bb _183_ (
    .a(_apc32_1_apc16_1_adder2_lv2_m3_d ),
    .b(_apc32_1_apc16_1_half1_a ),
    .c(_056_)
  );
  and_bi _184_ (
    .a(_056_),
    .b(_apc32_1_apc16_1_half1_cout ),
    .c(_apc32_1_apc16_1_half1_s )
  );
  and_bb _185_ (
    .a(_apc32_1_apc16_1_half1_cout ),
    .b(_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_apc32_1_apc16_1_half2_cout )
  );
  or_bb _186_ (
    .a(_apc32_1_apc16_1_half1_cout ),
    .b(_apc32_1_apc16_1_adder1_lv2_m3_d ),
    .c(_057_)
  );
  and_bi _187_ (
    .a(_057_),
    .b(_apc32_1_apc16_1_half2_cout ),
    .c(_apc32_1_apc16_1_half2_s )
  );
  and_bb _188_ (
    .a(_apc32_1_apc16_1_half2_cout ),
    .b(_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_apc32_1_apc16_1_half3_cout )
  );
  or_bb _189_ (
    .a(_apc32_1_apc16_1_half2_cout ),
    .b(_apc32_1_apc16_1_adder1_lv2_cout ),
    .c(_058_)
  );
  and_bi _190_ (
    .a(_058_),
    .b(_apc32_1_apc16_1_half3_cout ),
    .c(_apc32_1_apc16_1_half3_s )
  );
  or_bb _191_ (
    .a(in_33_),
    .b(in_32_),
    .c(_apc32_1_apc16_2_adder1_lv1_a )
  );
  and_bb _192_ (
    .a(in_35_),
    .b(in_34_),
    .c(_apc32_1_apc16_2_adder1_lv1_b )
  );
  or_bb _193_ (
    .a(in_37_),
    .b(in_36_),
    .c(_apc32_1_apc16_2_adder1_lv1_cin )
  );
  and_bb _194_ (
    .a(in_39_),
    .b(in_38_),
    .c(_apc32_1_apc16_2_adder2_lv1_a )
  );
  or_bb _195_ (
    .a(in_41_),
    .b(in_40_),
    .c(_apc32_1_apc16_2_adder2_lv1_b )
  );
  and_bb _196_ (
    .a(in_43_),
    .b(in_42_),
    .c(_apc32_1_apc16_2_adder2_lv1_cin )
  );
  or_bb _197_ (
    .a(in_45_),
    .b(in_44_),
    .c(_apc32_1_apc16_2_adder2_lv2_cin )
  );
  and_bb _198_ (
    .a(in_47_),
    .b(in_46_),
    .c(_apc32_1_apc16_2_half1_a )
  );
  maj_bbb _199_ (
    .a(_apc32_1_apc16_2_adder1_lv1_cin ),
    .b(_apc32_1_apc16_2_adder1_lv1_b ),
    .c(_apc32_1_apc16_2_adder1_lv1_a ),
    .d(_apc32_1_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _200_ (
    .a(_apc32_1_apc16_2_adder1_lv1_b ),
    .b(_apc32_1_apc16_2_adder1_lv1_a ),
    .c(_apc32_1_apc16_2_adder1_lv1_cin ),
    .d(_apc32_1_apc16_2_adder1_lv1_d )
  );
  maj_bbi _201_ (
    .a(_apc32_1_apc16_2_adder1_lv1_d ),
    .b(_apc32_1_apc16_2_adder1_lv1_cin ),
    .c(_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc32_1_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _202_ (
    .a(_apc32_1_apc16_2_adder1_lv2_cin ),
    .b(_apc32_1_apc16_2_adder1_lv2_b ),
    .c(_apc32_1_apc16_2_adder1_lv1_cout ),
    .d(_apc32_1_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _203_ (
    .a(_apc32_1_apc16_2_adder1_lv2_b ),
    .b(_apc32_1_apc16_2_adder1_lv1_cout ),
    .c(_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc32_1_apc16_2_adder1_lv2_d )
  );
  maj_bbi _204_ (
    .a(_apc32_1_apc16_2_adder1_lv2_d ),
    .b(_apc32_1_apc16_2_adder1_lv2_cin ),
    .c(_apc32_1_apc16_2_adder1_lv2_cout ),
    .d(_apc32_1_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _205_ (
    .a(_apc32_1_apc16_2_adder2_lv1_cin ),
    .b(_apc32_1_apc16_2_adder2_lv1_b ),
    .c(_apc32_1_apc16_2_adder2_lv1_a ),
    .d(_apc32_1_apc16_2_adder1_lv2_b )
  );
  maj_bbi _206_ (
    .a(_apc32_1_apc16_2_adder2_lv1_b ),
    .b(_apc32_1_apc16_2_adder2_lv1_a ),
    .c(_apc32_1_apc16_2_adder2_lv1_cin ),
    .d(_apc32_1_apc16_2_adder2_lv1_d )
  );
  maj_bbi _207_ (
    .a(_apc32_1_apc16_2_adder2_lv1_d ),
    .b(_apc32_1_apc16_2_adder2_lv1_cin ),
    .c(_apc32_1_apc16_2_adder1_lv2_b ),
    .d(_apc32_1_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _208_ (
    .a(_apc32_1_apc16_2_adder2_lv2_cin ),
    .b(_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .c(_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .d(_apc32_1_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _209_ (
    .a(_apc32_1_apc16_2_adder2_lv1_m3_d ),
    .b(_apc32_1_apc16_2_adder1_lv1_m3_d ),
    .c(_apc32_1_apc16_2_adder2_lv2_cin ),
    .d(_apc32_1_apc16_2_adder2_lv2_d )
  );
  maj_bbi _210_ (
    .a(_apc32_1_apc16_2_adder2_lv2_d ),
    .b(_apc32_1_apc16_2_adder2_lv2_cin ),
    .c(_apc32_1_apc16_2_adder1_lv2_cin ),
    .d(_apc32_1_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _211_ (
    .a(_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc32_1_apc16_2_half1_a ),
    .c(_apc32_1_apc16_2_half1_cout )
  );
  or_bb _212_ (
    .a(_apc32_1_apc16_2_adder2_lv2_m3_d ),
    .b(_apc32_1_apc16_2_half1_a ),
    .c(_059_)
  );
  and_bi _213_ (
    .a(_059_),
    .b(_apc32_1_apc16_2_half1_cout ),
    .c(_apc32_1_apc16_2_half1_s )
  );
  and_bb _214_ (
    .a(_apc32_1_apc16_2_half1_cout ),
    .b(_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_apc32_1_apc16_2_half2_cout )
  );
  or_bb _215_ (
    .a(_apc32_1_apc16_2_half1_cout ),
    .b(_apc32_1_apc16_2_adder1_lv2_m3_d ),
    .c(_060_)
  );
  and_bi _216_ (
    .a(_060_),
    .b(_apc32_1_apc16_2_half2_cout ),
    .c(_apc32_1_apc16_2_half2_s )
  );
  and_bb _217_ (
    .a(_apc32_1_apc16_2_half2_cout ),
    .b(_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_apc32_1_apc16_2_half3_cout )
  );
  or_bb _218_ (
    .a(_apc32_1_apc16_2_half2_cout ),
    .b(_apc32_1_apc16_2_adder1_lv2_cout ),
    .c(_061_)
  );
  and_bi _219_ (
    .a(_061_),
    .b(_apc32_1_apc16_2_half3_cout ),
    .c(_apc32_1_apc16_2_half3_s )
  );
  or_ii _220_ (
    .a(1'b0),
    .b(1'b0),
    .c(_062_)
  );
  or_ii _221_ (
    .a(_apc32_2_apc16_2_half1_s ),
    .b(_apc32_2_apc16_1_half1_s ),
    .c(_063_)
  );
  and_ii _222_ (
    .a(_apc32_2_apc16_2_half1_s ),
    .b(_apc32_2_apc16_1_half1_s ),
    .c(_064_)
  );
  and_bi _223_ (
    .a(_063_),
    .b(_064_),
    .c(_065_)
  );
  or_bi _224_ (
    .a(_062_),
    .b(_065_),
    .c(_066_)
  );
  and_bi _225_ (
    .a(_062_),
    .b(_065_),
    .c(_067_)
  );
  and_bi _226_ (
    .a(_066_),
    .b(_067_),
    .c(_apc32_2_out_1_)
  );
  maj_bii _227_ (
    .a(_062_),
    .b(_apc32_2_apc16_2_half1_s ),
    .c(_apc32_2_apc16_1_half1_s ),
    .d(_068_)
  );
  or_ii _228_ (
    .a(_apc32_2_apc16_2_half2_s ),
    .b(_apc32_2_apc16_1_half2_s ),
    .c(_069_)
  );
  and_ii _229_ (
    .a(_apc32_2_apc16_2_half2_s ),
    .b(_apc32_2_apc16_1_half2_s ),
    .c(_070_)
  );
  and_bi _230_ (
    .a(_069_),
    .b(_070_),
    .c(_071_)
  );
  or_bi _231_ (
    .a(_068_),
    .b(_071_),
    .c(_072_)
  );
  and_bi _232_ (
    .a(_068_),
    .b(_071_),
    .c(_073_)
  );
  and_bi _233_ (
    .a(_072_),
    .b(_073_),
    .c(_apc32_2_out_2_)
  );
  maj_bii _234_ (
    .a(_068_),
    .b(_apc32_2_apc16_2_half2_s ),
    .c(_apc32_2_apc16_1_half2_s ),
    .d(_074_)
  );
  or_ii _235_ (
    .a(_apc32_2_apc16_2_half3_s ),
    .b(_apc32_2_apc16_1_half3_s ),
    .c(_075_)
  );
  and_ii _236_ (
    .a(_apc32_2_apc16_2_half3_s ),
    .b(_apc32_2_apc16_1_half3_s ),
    .c(_076_)
  );
  and_bi _237_ (
    .a(_075_),
    .b(_076_),
    .c(_077_)
  );
  or_bi _238_ (
    .a(_074_),
    .b(_077_),
    .c(_078_)
  );
  and_bi _239_ (
    .a(_074_),
    .b(_077_),
    .c(_079_)
  );
  and_bi _240_ (
    .a(_078_),
    .b(_079_),
    .c(_apc32_2_out_3_)
  );
  maj_bii _241_ (
    .a(_074_),
    .b(_apc32_2_apc16_2_half3_s ),
    .c(_apc32_2_apc16_1_half3_s ),
    .d(_080_)
  );
  or_ii _242_ (
    .a(_apc32_2_apc16_2_half3_cout ),
    .b(_apc32_2_apc16_1_half3_cout ),
    .c(_081_)
  );
  and_ii _243_ (
    .a(_apc32_2_apc16_2_half3_cout ),
    .b(_apc32_2_apc16_1_half3_cout ),
    .c(_082_)
  );
  and_bi _244_ (
    .a(_081_),
    .b(_082_),
    .c(_083_)
  );
  or_bi _245_ (
    .a(_080_),
    .b(_083_),
    .c(_084_)
  );
  and_bi _246_ (
    .a(_080_),
    .b(_083_),
    .c(_085_)
  );
  and_bi _247_ (
    .a(_084_),
    .b(_085_),
    .c(_apc32_2_out_4_)
  );
  and_ii _248_ (
    .a(1'b0),
    .b(1'b0),
    .c(_086_)
  );
  and_bi _249_ (
    .a(_062_),
    .b(_086_),
    .c(_apc32_2_out_0_)
  );
  maj_bbi _250_ (
    .a(_apc32_2_apc16_2_half3_cout ),
    .b(_apc32_2_apc16_1_half3_cout ),
    .c(_080_),
    .d(_apc32_2_out_5_)
  );
  or_bb _251_ (
    .a(in_17_),
    .b(in_16_),
    .c(_apc32_2_apc16_1_adder1_lv1_a )
  );
  and_bb _252_ (
    .a(in_19_),
    .b(in_18_),
    .c(_apc32_2_apc16_1_adder1_lv1_b )
  );
  or_bb _253_ (
    .a(in_21_),
    .b(in_20_),
    .c(_apc32_2_apc16_1_adder1_lv1_cin )
  );
  and_bb _254_ (
    .a(in_23_),
    .b(in_22_),
    .c(_apc32_2_apc16_1_adder2_lv1_a )
  );
  or_bb _255_ (
    .a(in_25_),
    .b(in_24_),
    .c(_apc32_2_apc16_1_adder2_lv1_b )
  );
  and_bb _256_ (
    .a(in_27_),
    .b(in_26_),
    .c(_apc32_2_apc16_1_adder2_lv1_cin )
  );
  or_bb _257_ (
    .a(in_29_),
    .b(in_28_),
    .c(_apc32_2_apc16_1_adder2_lv2_cin )
  );
  and_bb _258_ (
    .a(in_31_),
    .b(in_30_),
    .c(_apc32_2_apc16_1_half1_a )
  );
  maj_bbb _259_ (
    .a(_apc32_2_apc16_1_adder1_lv1_cin ),
    .b(_apc32_2_apc16_1_adder1_lv1_b ),
    .c(_apc32_2_apc16_1_adder1_lv1_a ),
    .d(_apc32_2_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _260_ (
    .a(_apc32_2_apc16_1_adder1_lv1_b ),
    .b(_apc32_2_apc16_1_adder1_lv1_a ),
    .c(_apc32_2_apc16_1_adder1_lv1_cin ),
    .d(_apc32_2_apc16_1_adder1_lv1_d )
  );
  maj_bbi _261_ (
    .a(_apc32_2_apc16_1_adder1_lv1_d ),
    .b(_apc32_2_apc16_1_adder1_lv1_cin ),
    .c(_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc32_2_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _262_ (
    .a(_apc32_2_apc16_1_adder1_lv2_cin ),
    .b(_apc32_2_apc16_1_adder1_lv2_b ),
    .c(_apc32_2_apc16_1_adder1_lv1_cout ),
    .d(_apc32_2_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _263_ (
    .a(_apc32_2_apc16_1_adder1_lv2_b ),
    .b(_apc32_2_apc16_1_adder1_lv1_cout ),
    .c(_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc32_2_apc16_1_adder1_lv2_d )
  );
  maj_bbi _264_ (
    .a(_apc32_2_apc16_1_adder1_lv2_d ),
    .b(_apc32_2_apc16_1_adder1_lv2_cin ),
    .c(_apc32_2_apc16_1_adder1_lv2_cout ),
    .d(_apc32_2_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _265_ (
    .a(_apc32_2_apc16_1_adder2_lv1_cin ),
    .b(_apc32_2_apc16_1_adder2_lv1_b ),
    .c(_apc32_2_apc16_1_adder2_lv1_a ),
    .d(_apc32_2_apc16_1_adder1_lv2_b )
  );
  maj_bbi _266_ (
    .a(_apc32_2_apc16_1_adder2_lv1_b ),
    .b(_apc32_2_apc16_1_adder2_lv1_a ),
    .c(_apc32_2_apc16_1_adder2_lv1_cin ),
    .d(_apc32_2_apc16_1_adder2_lv1_d )
  );
  maj_bbi _267_ (
    .a(_apc32_2_apc16_1_adder2_lv1_d ),
    .b(_apc32_2_apc16_1_adder2_lv1_cin ),
    .c(_apc32_2_apc16_1_adder1_lv2_b ),
    .d(_apc32_2_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _268_ (
    .a(_apc32_2_apc16_1_adder2_lv2_cin ),
    .b(_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .c(_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .d(_apc32_2_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _269_ (
    .a(_apc32_2_apc16_1_adder2_lv1_m3_d ),
    .b(_apc32_2_apc16_1_adder1_lv1_m3_d ),
    .c(_apc32_2_apc16_1_adder2_lv2_cin ),
    .d(_apc32_2_apc16_1_adder2_lv2_d )
  );
  maj_bbi _270_ (
    .a(_apc32_2_apc16_1_adder2_lv2_d ),
    .b(_apc32_2_apc16_1_adder2_lv2_cin ),
    .c(_apc32_2_apc16_1_adder1_lv2_cin ),
    .d(_apc32_2_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _271_ (
    .a(_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc32_2_apc16_1_half1_a ),
    .c(_apc32_2_apc16_1_half1_cout )
  );
  or_bb _272_ (
    .a(_apc32_2_apc16_1_adder2_lv2_m3_d ),
    .b(_apc32_2_apc16_1_half1_a ),
    .c(_087_)
  );
  and_bi _273_ (
    .a(_087_),
    .b(_apc32_2_apc16_1_half1_cout ),
    .c(_apc32_2_apc16_1_half1_s )
  );
  and_bb _274_ (
    .a(_apc32_2_apc16_1_half1_cout ),
    .b(_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_apc32_2_apc16_1_half2_cout )
  );
  or_bb _275_ (
    .a(_apc32_2_apc16_1_half1_cout ),
    .b(_apc32_2_apc16_1_adder1_lv2_m3_d ),
    .c(_088_)
  );
  and_bi _276_ (
    .a(_088_),
    .b(_apc32_2_apc16_1_half2_cout ),
    .c(_apc32_2_apc16_1_half2_s )
  );
  and_bb _277_ (
    .a(_apc32_2_apc16_1_half2_cout ),
    .b(_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_apc32_2_apc16_1_half3_cout )
  );
  or_bb _278_ (
    .a(_apc32_2_apc16_1_half2_cout ),
    .b(_apc32_2_apc16_1_adder1_lv2_cout ),
    .c(_089_)
  );
  and_bi _279_ (
    .a(_089_),
    .b(_apc32_2_apc16_1_half3_cout ),
    .c(_apc32_2_apc16_1_half3_s )
  );
  or_bb _280_ (
    .a(in_1_),
    .b(in_0_),
    .c(_apc32_2_apc16_2_adder1_lv1_a )
  );
  and_bb _281_ (
    .a(in_3_),
    .b(in_2_),
    .c(_apc32_2_apc16_2_adder1_lv1_b )
  );
  or_bb _282_ (
    .a(in_5_),
    .b(in_4_),
    .c(_apc32_2_apc16_2_adder1_lv1_cin )
  );
  and_bb _283_ (
    .a(in_7_),
    .b(in_6_),
    .c(_apc32_2_apc16_2_adder2_lv1_a )
  );
  or_bb _284_ (
    .a(in_9_),
    .b(in_8_),
    .c(_apc32_2_apc16_2_adder2_lv1_b )
  );
  and_bb _285_ (
    .a(in_11_),
    .b(in_10_),
    .c(_apc32_2_apc16_2_adder2_lv1_cin )
  );
  or_bb _286_ (
    .a(in_13_),
    .b(in_12_),
    .c(_apc32_2_apc16_2_adder2_lv2_cin )
  );
  and_bb _287_ (
    .a(in_15_),
    .b(in_14_),
    .c(_apc32_2_apc16_2_half1_a )
  );
  maj_bbb _288_ (
    .a(_apc32_2_apc16_2_adder1_lv1_cin ),
    .b(_apc32_2_apc16_2_adder1_lv1_b ),
    .c(_apc32_2_apc16_2_adder1_lv1_a ),
    .d(_apc32_2_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _289_ (
    .a(_apc32_2_apc16_2_adder1_lv1_b ),
    .b(_apc32_2_apc16_2_adder1_lv1_a ),
    .c(_apc32_2_apc16_2_adder1_lv1_cin ),
    .d(_apc32_2_apc16_2_adder1_lv1_d )
  );
  maj_bbi _290_ (
    .a(_apc32_2_apc16_2_adder1_lv1_d ),
    .b(_apc32_2_apc16_2_adder1_lv1_cin ),
    .c(_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc32_2_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _291_ (
    .a(_apc32_2_apc16_2_adder1_lv2_cin ),
    .b(_apc32_2_apc16_2_adder1_lv2_b ),
    .c(_apc32_2_apc16_2_adder1_lv1_cout ),
    .d(_apc32_2_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _292_ (
    .a(_apc32_2_apc16_2_adder1_lv2_b ),
    .b(_apc32_2_apc16_2_adder1_lv1_cout ),
    .c(_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc32_2_apc16_2_adder1_lv2_d )
  );
  maj_bbi _293_ (
    .a(_apc32_2_apc16_2_adder1_lv2_d ),
    .b(_apc32_2_apc16_2_adder1_lv2_cin ),
    .c(_apc32_2_apc16_2_adder1_lv2_cout ),
    .d(_apc32_2_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _294_ (
    .a(_apc32_2_apc16_2_adder2_lv1_cin ),
    .b(_apc32_2_apc16_2_adder2_lv1_b ),
    .c(_apc32_2_apc16_2_adder2_lv1_a ),
    .d(_apc32_2_apc16_2_adder1_lv2_b )
  );
  maj_bbi _295_ (
    .a(_apc32_2_apc16_2_adder2_lv1_b ),
    .b(_apc32_2_apc16_2_adder2_lv1_a ),
    .c(_apc32_2_apc16_2_adder2_lv1_cin ),
    .d(_apc32_2_apc16_2_adder2_lv1_d )
  );
  maj_bbi _296_ (
    .a(_apc32_2_apc16_2_adder2_lv1_d ),
    .b(_apc32_2_apc16_2_adder2_lv1_cin ),
    .c(_apc32_2_apc16_2_adder1_lv2_b ),
    .d(_apc32_2_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _297_ (
    .a(_apc32_2_apc16_2_adder2_lv2_cin ),
    .b(_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .c(_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .d(_apc32_2_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _298_ (
    .a(_apc32_2_apc16_2_adder2_lv1_m3_d ),
    .b(_apc32_2_apc16_2_adder1_lv1_m3_d ),
    .c(_apc32_2_apc16_2_adder2_lv2_cin ),
    .d(_apc32_2_apc16_2_adder2_lv2_d )
  );
  maj_bbi _299_ (
    .a(_apc32_2_apc16_2_adder2_lv2_d ),
    .b(_apc32_2_apc16_2_adder2_lv2_cin ),
    .c(_apc32_2_apc16_2_adder1_lv2_cin ),
    .d(_apc32_2_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _300_ (
    .a(_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc32_2_apc16_2_half1_a ),
    .c(_apc32_2_apc16_2_half1_cout )
  );
  or_bb _301_ (
    .a(_apc32_2_apc16_2_adder2_lv2_m3_d ),
    .b(_apc32_2_apc16_2_half1_a ),
    .c(_090_)
  );
  and_bi _302_ (
    .a(_090_),
    .b(_apc32_2_apc16_2_half1_cout ),
    .c(_apc32_2_apc16_2_half1_s )
  );
  and_bb _303_ (
    .a(_apc32_2_apc16_2_half1_cout ),
    .b(_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_apc32_2_apc16_2_half2_cout )
  );
  or_bb _304_ (
    .a(_apc32_2_apc16_2_half1_cout ),
    .b(_apc32_2_apc16_2_adder1_lv2_m3_d ),
    .c(_091_)
  );
  and_bi _305_ (
    .a(_091_),
    .b(_apc32_2_apc16_2_half2_cout ),
    .c(_apc32_2_apc16_2_half2_s )
  );
  and_bb _306_ (
    .a(_apc32_2_apc16_2_half2_cout ),
    .b(_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_apc32_2_apc16_2_half3_cout )
  );
  or_bb _307_ (
    .a(_apc32_2_apc16_2_half2_cout ),
    .b(_apc32_2_apc16_2_adder1_lv2_cout ),
    .c(_092_)
  );
  and_bi _308_ (
    .a(_092_),
    .b(_apc32_2_apc16_2_half3_cout ),
    .c(_apc32_2_apc16_2_half3_s )
  );
endmodule
