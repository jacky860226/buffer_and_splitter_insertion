module c1355(G27,G41,G37,G21,G18,G24,G33,G30,G4,G3,G23,G39,G7,G1,G25,G19,G13,G17,G16,G22,G36,G6,G26,G31,G2,G12,G20,G29,G5,G28,G15,G9,G8,G14,G34,G10,G32,G35,G11,G38,G40);
    wire _090_;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_8;
    wire _255_;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_1647;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_739;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_24;
    wire _042_;
    wire _035_;
    wire _181_;
    wire new_Jinkela_wire_1479;
    wire _095_;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_870;
    wire _119_;
    wire _317_;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_1287;
    wire _054_;
    wire new_Jinkela_wire_775;
    wire _022_;
    wire _272_;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_254;
    wire _017_;
    wire _069_;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_1015;
    wire _316_;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_233;
    wire new_net_710;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_20;
    wire _012_;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_1408;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_612;
    wire _257_;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_366;
    wire _002_;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_1378;
    wire _268_;
    wire _282_;
    wire _217_;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_1518;
    wire _292_;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_1554;
    wire _333_;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_954;
    wire new_net_728;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_283;
    wire _123_;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_613;
    wire _320_;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_118;
    wire _122_;
    wire new_Jinkela_wire_1309;
    wire _187_;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_126;
    wire _089_;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_925;
    wire _267_;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_1069;
    wire _328_;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_66;
    wire _156_;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_930;
    wire new_Jinkela_wire_1;
    wire new_net_712;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_1281;
    wire _127_;
    wire new_Jinkela_wire_1530;
    wire _322_;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_1403;
    wire _212_;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_9;
    wire _053_;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_653;
    wire _068_;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_358;
    wire _265_;
    wire new_Jinkela_wire_457;
    wire _291_;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_251;
    wire _321_;
    wire _107_;
    wire _347_;
    wire _109_;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_553;
    wire new_net_708;
    wire new_Jinkela_wire_341;
    wire _007_;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_1137;
    wire _228_;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_786;
    wire _238_;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_79;
    wire new_net_694;
    wire _294_;
    wire _006_;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_950;
    wire new_net_722;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_415;
    wire _326_;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_528;
    wire _227_;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_87;
    wire _307_;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_437;
    wire _061_;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_1553;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_40;
    wire _281_;
    wire _205_;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_1108;
    wire _224_;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_830;
    wire _142_;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_1089;
    wire _311_;
    wire _164_;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_1145;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_857;
    wire _072_;
    wire new_Jinkela_wire_1191;
    wire _241_;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_371;
    wire _262_;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_1303;
    wire _044_;
    wire new_Jinkela_wire_150;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_1086;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_1512;
    wire _349_;
    wire _121_;
    wire new_Jinkela_wire_1617;
    wire _234_;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_1485;
    wire _008_;
    wire new_Jinkela_wire_311;
    wire _312_;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_1536;
    wire _271_;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_1569;
    wire _067_;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_851;
    wire _276_;
    wire _160_;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_797;
    wire _084_;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_310;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_1389;
    wire _278_;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_46;
    wire _049_;
    wire _085_;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_493;
    wire _159_;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_372;
    wire _210_;
    wire _232_;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_953;
    wire _176_;
    wire _339_;
    wire _093_;
    wire new_Jinkela_wire_552;
    wire _249_;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_748;
    wire new_net_686;
    wire new_Jinkela_wire_730;
    wire _298_;
    wire new_Jinkela_wire_891;
    wire _152_;
    wire new_Jinkela_wire_721;
    wire _088_;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_1324;
    wire _340_;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_1182;
    wire _200_;
    wire new_Jinkela_wire_859;
    wire _021_;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_107;
    wire _075_;
    wire _153_;
    wire _352_;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_1283;
    wire _080_;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_1169;
    wire _169_;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_401;
    wire _018_;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_1343;
    wire _237_;
    wire _043_;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_105;
    wire _304_;
    wire _259_;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_1239;
    wire _233_;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_1521;
    wire _225_;
    wire new_net_682;
    wire new_Jinkela_wire_1292;
    wire _261_;
    wire new_Jinkela_wire_1286;
    wire new_Jinkela_wire_113;
    wire _112_;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_559;
    wire _288_;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_687;
    wire _150_;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_266;
    wire _215_;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_1331;
    wire _342_;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_1093;
    wire _149_;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_1299;
    wire _223_;
    wire new_Jinkela_wire_1110;
    wire _062_;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_755;
    wire _036_;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_1082;
    wire _030_;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_1263;
    wire _229_;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_554;
    wire _277_;
    wire _325_;
    wire new_Jinkela_wire_649;
    wire _270_;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_999;
    wire _216_;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_1112;
    wire _258_;
    wire new_Jinkela_wire_783;
    wire _284_;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_742;
    wire _014_;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_1284;
    wire _243_;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_1078;
    wire _055_;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_111;
    wire _252_;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_766;
    wire _310_;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_438;
    wire _295_;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_1135;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_1151;
    wire _050_;
    wire new_Jinkela_wire_1092;
    wire _336_;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_605;
    wire _195_;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_1591;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_1097;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_836;
    wire _226_;
    wire new_Jinkela_wire_1398;
    wire _019_;
    wire new_Jinkela_wire_936;
    wire _148_;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_494;
    wire _344_;
    wire new_Jinkela_wire_458;
    wire _133_;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_430;
    wire new_net_702;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_781;
    wire _132_;
    wire new_Jinkela_wire_1063;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_904;
    wire _048_;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_39;
    wire _254_;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_1142;
    wire _345_;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_1450;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_326;
    wire _173_;
    wire new_Jinkela_wire_1635;
    wire _025_;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_1407;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_908;
    wire _015_;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_1440;
    wire _034_;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_623;
    wire _059_;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_1567;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_1276;
    wire _172_;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_1037;
    wire _263_;
    wire new_Jinkela_wire_396;
    wire _016_;
    wire new_Jinkela_wire_679;
    wire _219_;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_1475;
    wire _166_;
    wire new_Jinkela_wire_509;
    wire _011_;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_835;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_180;
    wire _086_;
    wire _091_;
    wire _031_;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_750;
    wire _060_;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_1421;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_1394;
    wire _182_;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_1186;
    wire _058_;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_608;
    wire _157_;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_1486;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_1141;
    wire _290_;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_1480;
    wire _028_;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_1194;
    wire _139_;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_1189;
    wire _247_;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_71;
    wire _197_;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_1252;
    wire _111_;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_1537;
    wire _300_;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_898;
    wire _348_;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_777;
    wire _202_;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_1630;
    wire _218_;
    wire _125_;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_1404;
    wire _302_;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_377;
    wire _114_;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_832;
    wire _190_;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_1562;
    wire new_net_692;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_435;
    wire _214_;
    wire _251_;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_1551;
    wire new_net_696;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_178;
    wire _242_;
    wire new_net_726;
    wire _178_;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_1358;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_1640;
    wire _355_;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_452;
    wire _032_;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_1114;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_133;
    wire _026_;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_1197;
    wire new_Jinkela_wire_55;
    wire _158_;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_1235;
    wire _128_;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_482;
    wire _273_;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_1397;
    wire _001_;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_1245;
    wire _033_;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_1636;
    wire _246_;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_597;
    wire _004_;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_1503;
    wire _180_;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_1495;
    wire _136_;
    wire new_Jinkela_wire_1159;
    wire _161_;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_1382;
    wire _013_;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_1393;
    wire _179_;
    wire new_Jinkela_wire_800;
    wire _305_;
    wire _131_;
    wire new_Jinkela_wire_84;
    wire _330_;
    wire _102_;
    wire new_Jinkela_wire_1014;
    wire _341_;
    wire new_Jinkela_wire_1452;
    wire _240_;
    wire _117_;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_895;
    wire _338_;
    wire _350_;
    wire _074_;
    wire _099_;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_1552;
    wire _235_;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_455;
    wire _335_;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_263;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_56;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_483;
    wire _083_;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_771;
    wire _155_;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_1073;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_929;
    wire _073_;
    wire new_Jinkela_wire_706;
    wire _253_;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_1002;
    wire _144_;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_1042;
    wire _005_;
    wire _289_;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_428;
    wire _076_;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_804;
    wire _285_;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_799;
    wire _275_;
    wire new_Jinkela_wire_200;
    wire _171_;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_1437;
    wire _167_;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_1380;
    wire _129_;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_1059;
    wire _287_;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_1184;
    wire _092_;
    wire new_Jinkela_wire_564;
    wire _313_;
    wire _301_;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_23;
    wire new_Jinkela_wire_1060;
    wire _115_;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_1514;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_1144;
    wire _087_;
    wire new_Jinkela_wire_1216;
    wire _244_;
    wire _329_;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_784;
    wire _020_;
    wire new_net_688;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_1101;
    wire _199_;
    wire _343_;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_279;
    wire _193_;
    wire new_Jinkela_wire_147;
    wire _207_;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_61;
    wire new_Jinkela_wire_669;
    wire _046_;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_1156;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_1412;
    wire _038_;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_1354;
    wire _296_;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_369;
    wire _078_;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_1103;
    wire _279_;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_1583;
    wire _185_;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_659;
    wire _047_;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_238;
    wire _239_;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_505;
    wire _071_;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_1326;
    wire new_Jinkela_wire_1055;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_591;
    wire _106_;
    wire _306_;
    wire new_net_716;
    wire _280_;
    wire new_Jinkela_wire_1212;
    wire _120_;
    wire new_Jinkela_wire_1381;
    wire _147_;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_557;
    wire _045_;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_232;
    wire _040_;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_210;
    wire _319_;
    wire new_Jinkela_wire_291;
    wire _094_;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_625;
    wire _145_;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_759;
    wire _297_;
    wire new_Jinkela_wire_850;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_1049;
    wire _209_;
    wire _256_;
    wire _337_;
    wire new_Jinkela_wire_516;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_420;
    wire _130_;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_293;
    wire _081_;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_914;
    wire _220_;
    wire new_Jinkela_wire_949;
    wire _351_;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_444;
    wire _357_;
    wire new_Jinkela_wire_1555;
    wire _327_;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_673;
    wire _332_;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_237;
    wire _211_;
    wire new_Jinkela_wire_1140;
    wire _027_;
    wire new_Jinkela_wire_1376;
    wire _113_;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_1258;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_566;
    wire _103_;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_565;
    wire _141_;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_1161;
    wire _334_;
    wire _168_;
    wire _000_;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_1224;
    wire _196_;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_4;
    wire _236_;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_468;
    wire _353_;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_972;
    wire _318_;
    wire _358_;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_1462;
    wire _293_;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_1166;
    wire _162_;
    wire new_Jinkela_wire_1298;
    wire _359_;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_1121;
    wire _077_;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_1545;
    wire _308_;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_294;
    wire _194_;
    wire _037_;
    wire new_net_724;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_933;
    wire new_net_706;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_1202;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_333;
    wire _009_;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_692;
    wire _175_;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_142;
    wire _303_;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_1445;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_1627;
    wire _070_;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_319;
    wire _116_;
    wire _143_;
    wire new_net_684;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_155;
    wire _137_;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_1050;
    wire _274_;
    wire new_net_718;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_578;
    wire _324_;
    wire new_Jinkela_wire_121;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_894;
    wire _221_;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_852;
    wire _192_;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_1294;
    wire new_net_700;
    wire _309_;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_638;
    wire _082_;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_1066;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_12;
    wire _188_;
    wire _023_;
    wire _346_;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_1105;
    wire _204_;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_1176;
    wire _191_;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_1234;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_1322;
    wire _134_;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_1361;
    wire _063_;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_346;
    wire _183_;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_1178;
    wire _051_;
    wire _138_;
    wire new_Jinkela_wire_876;
    wire _066_;
    wire _283_;
    wire _041_;
    wire _079_;
    wire new_Jinkela_wire_1626;
    wire _146_;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_1190;
    wire _186_;
    wire _024_;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_1200;
    wire new_net_704;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_1016;
    wire _189_;
    wire new_Jinkela_wire_137;
    wire _208_;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_1405;
    wire _331_;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_1341;
    wire _065_;
    wire new_net_690;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_806;
    wire _039_;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_1549;
    wire _096_;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_1266;
    wire _100_;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_149;
    wire _198_;
    wire _101_;
    wire new_Jinkela_wire_1315;
    wire new_Jinkela_wire_1233;
    wire _230_;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_314;
    wire _354_;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_701;
    wire _206_;
    wire _098_;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_1506;
    wire new_Jinkela_wire_1119;
    wire _105_;
    wire _118_;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_1612;
    wire new_net_720;
    wire _052_;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_241;
    wire _248_;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_751;
    wire _003_;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_1571;
    wire _104_;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_1040;
    wire _269_;
    wire new_Jinkela_wire_1111;
    wire _201_;
    wire new_Jinkela_wire_477;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_88;
    wire _126_;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_226;
    wire _124_;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_248;
    wire _108_;
    wire new_Jinkela_wire_480;
    wire _165_;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_1333;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_304;
    wire _203_;
    wire _213_;
    wire new_Jinkela_wire_1154;
    wire _010_;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_924;
    wire _177_;
    wire _029_;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_896;
    wire _151_;
    wire new_net_714;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_579;
    wire _097_;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_769;
    wire _163_;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_86;
    wire _231_;
    wire new_Jinkela_wire_1643;
    wire _170_;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_93;
    wire _286_;
    wire _140_;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_1262;
    wire _056_;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_720;
    wire _245_;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_1057;
    wire _356_;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_1439;
    wire _264_;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_966;
    wire _266_;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_1126;
    wire _315_;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_1011;
    wire _154_;
    wire new_Jinkela_wire_725;
    wire _110_;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_1436;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_1153;
    wire _174_;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_675;
    wire new_net_698;
    wire _314_;
    wire _323_;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_1307;
    wire _064_;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_1036;
    wire _222_;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_337;
    wire _260_;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_734;
    wire _184_;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_1420;
    wire _135_;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_952;
    wire _299_;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_956;
    wire _250_;
    wire new_Jinkela_wire_981;
    wire _057_;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_1391;
    input G27;
    input G41;
    input G37;
    input G21;
    input G18;
    input G24;
    input G33;
    input G30;
    input G4;
    input G3;
    input G23;
    input G39;
    input G7;
    input G1;
    input G25;
    input G19;
    input G13;
    input G17;
    input G16;
    input G22;
    input G36;
    input G6;
    input G26;
    input G31;
    input G2;
    input G12;
    input G20;
    input G29;
    input G5;
    input G28;
    input G15;
    input G9;
    input G8;
    input G14;
    input G34;
    input G10;
    input G32;
    input G35;
    input G11;
    input G38;
    input G40;
    output G1335;
    output G1336;
    output G1348;
    output G1324;
    output G1337;
    output G1350;
    output G1332;
    output G1326;
    output G1346;
    output G1344;
    output G1354;
    output G1341;
    output G1342;
    output G1347;
    output G1349;
    output G1328;
    output G1355;
    output G1327;
    output G1338;
    output G1334;
    output G1352;
    output G1331;
    output G1340;
    output G1343;
    output G1339;
    output G1329;
    output G1353;
    output G1330;
    output G1325;
    output G1351;
    output G1333;
    output G1345;

    and_bi _473_ (
        .a(new_Jinkela_wire_1251),
        .b(new_Jinkela_wire_1222),
        .c(_087_)
    );

    and_bi _474_ (
        .a(new_Jinkela_wire_1221),
        .b(new_Jinkela_wire_1252),
        .c(_088_)
    );

    or_bb _475_ (
        .a(_088_),
        .b(_087_),
        .c(_089_)
    );

    or_bi _476_ (
        .a(new_Jinkela_wire_341),
        .b(new_Jinkela_wire_48),
        .c(_090_)
    );

    and_bi _477_ (
        .a(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_46),
        .c(_091_)
    );

    or_bi _478_ (
        .a(_091_),
        .b(_090_),
        .c(_092_)
    );

    or_bb _479_ (
        .a(new_Jinkela_wire_437),
        .b(new_Jinkela_wire_730),
        .c(_093_)
    );

    and_bb _480_ (
        .a(new_Jinkela_wire_438),
        .b(new_Jinkela_wire_731),
        .c(_094_)
    );

    or_bi _481_ (
        .a(_094_),
        .b(_093_),
        .c(_095_)
    );

    or_bi _482_ (
        .a(new_Jinkela_wire_1349),
        .b(new_Jinkela_wire_1066),
        .c(_096_)
    );

    and_bi _483_ (
        .a(new_Jinkela_wire_1350),
        .b(new_Jinkela_wire_1067),
        .c(_097_)
    );

    and_bi _484_ (
        .a(_096_),
        .b(_097_),
        .c(_098_)
    );

    and_bi _485_ (
        .a(new_Jinkela_wire_1543),
        .b(new_Jinkela_wire_1630),
        .c(_099_)
    );

    and_bi _486_ (
        .a(new_Jinkela_wire_1631),
        .b(new_Jinkela_wire_1544),
        .c(_100_)
    );

    or_bb _487_ (
        .a(_100_),
        .b(_099_),
        .c(_101_)
    );

    or_bb _488_ (
        .a(new_Jinkela_wire_1521),
        .b(new_Jinkela_wire_1086),
        .c(_102_)
    );

    and_bb _489_ (
        .a(new_Jinkela_wire_1522),
        .b(new_Jinkela_wire_1087),
        .c(_103_)
    );

    and_bi _490_ (
        .a(_102_),
        .b(_103_),
        .c(_104_)
    );

    or_ii _491_ (
        .a(new_Jinkela_wire_1055),
        .b(new_Jinkela_wire_34),
        .c(_105_)
    );

    and_bi _492_ (
        .a(new_Jinkela_wire_1549),
        .b(new_Jinkela_wire_1291),
        .c(_106_)
    );

    and_bi _493_ (
        .a(new_Jinkela_wire_1294),
        .b(new_Jinkela_wire_1550),
        .c(_107_)
    );

    or_bb _494_ (
        .a(_107_),
        .b(_106_),
        .c(_108_)
    );

    or_bi _495_ (
        .a(new_Jinkela_wire_77),
        .b(new_Jinkela_wire_564),
        .c(_109_)
    );

    and_bi _496_ (
        .a(new_Jinkela_wire_76),
        .b(new_Jinkela_wire_565),
        .c(_110_)
    );

    or_bi _497_ (
        .a(_110_),
        .b(_109_),
        .c(_111_)
    );

    or_bb _498_ (
        .a(new_Jinkela_wire_498),
        .b(new_Jinkela_wire_142),
        .c(_112_)
    );

    and_bb _499_ (
        .a(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_141),
        .c(_113_)
    );

    or_bi _500_ (
        .a(_113_),
        .b(_112_),
        .c(_114_)
    );

    or_bi _501_ (
        .a(new_Jinkela_wire_1257),
        .b(new_Jinkela_wire_1271),
        .c(_115_)
    );

    and_bi _502_ (
        .a(new_Jinkela_wire_1258),
        .b(new_Jinkela_wire_1272),
        .c(_116_)
    );

    and_bi _503_ (
        .a(_115_),
        .b(_116_),
        .c(_117_)
    );

    and_bi _504_ (
        .a(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1072),
        .c(_118_)
    );

    and_bi _505_ (
        .a(new_Jinkela_wire_1070),
        .b(new_Jinkela_wire_1334),
        .c(_119_)
    );

    or_bb _506_ (
        .a(_119_),
        .b(_118_),
        .c(_120_)
    );

    or_bb _507_ (
        .a(new_Jinkela_wire_1396),
        .b(new_Jinkela_wire_1586),
        .c(_121_)
    );

    and_bb _508_ (
        .a(new_Jinkela_wire_1397),
        .b(new_Jinkela_wire_1587),
        .c(_122_)
    );

    or_bi _509_ (
        .a(new_Jinkela_wire_1084),
        .b(new_Jinkela_wire_1135),
        .c(_123_)
    );

    or_bb _510_ (
        .a(_123_),
        .b(new_Jinkela_wire_1556),
        .c(_124_)
    );

    and_bb _511_ (
        .a(new_Jinkela_wire_955),
        .b(new_Jinkela_wire_35),
        .c(_125_)
    );

    or_bb _512_ (
        .a(new_Jinkela_wire_145),
        .b(new_Jinkela_wire_728),
        .c(_126_)
    );

    and_bb _513_ (
        .a(new_Jinkela_wire_144),
        .b(new_Jinkela_wire_732),
        .c(_127_)
    );

    and_bi _514_ (
        .a(_126_),
        .b(_127_),
        .c(_128_)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_136),
        .c(new_Jinkela_wire_137),
        .b(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_686),
        .dout(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_180),
        .dout(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_155),
        .dout(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    spl2 new_Jinkela_splitter_78 (
        .a(G15),
        .c(new_Jinkela_wire_824),
        .b(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_244),
        .dout(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_210),
        .dout(new_Jinkela_wire_211)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_157),
        .dout(new_Jinkela_wire_158)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_158),
        .dout(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_211),
        .dout(new_Jinkela_wire_212)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_159),
        .dout(new_Jinkela_wire_160)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    spl2 new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_691),
        .c(new_Jinkela_wire_692),
        .b(new_Jinkela_wire_693)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_160),
        .dout(new_Jinkela_wire_161)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_764),
        .dout(new_Jinkela_wire_765)
    );

    spl3L new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_794),
        .d(new_Jinkela_wire_795),
        .c(new_Jinkela_wire_796),
        .b(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_161),
        .dout(new_Jinkela_wire_162)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_737),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_162),
        .dout(new_Jinkela_wire_163)
    );

    spl3L new_Jinkela_splitter_81 (
        .a(G9),
        .d(new_Jinkela_wire_856),
        .c(new_Jinkela_wire_857),
        .b(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_212),
        .dout(new_Jinkela_wire_213)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_163),
        .dout(new_Jinkela_wire_164)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_164),
        .dout(new_Jinkela_wire_165)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_765),
        .dout(new_Jinkela_wire_766)
    );

    spl2 new_Jinkela_splitter_30 (
        .a(G1),
        .c(new_Jinkela_wire_304),
        .b(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_238),
        .dout(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_739),
        .dout(new_Jinkela_wire_740)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_716),
        .dout(new_Jinkela_wire_717)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_166),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_213),
        .dout(new_Jinkela_wire_214)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_167),
        .dout(new_Jinkela_wire_168)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    spl2 new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_168),
        .c(new_Jinkela_wire_169),
        .b(new_Jinkela_wire_170)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    spl4L new_Jinkela_splitter_31 (
        .a(new_Jinkela_wire_306),
        .d(new_Jinkela_wire_307),
        .e(new_Jinkela_wire_308),
        .c(new_Jinkela_wire_309),
        .b(new_Jinkela_wire_310)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    spl4L new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_826),
        .d(new_Jinkela_wire_827),
        .e(new_Jinkela_wire_828),
        .c(new_Jinkela_wire_829),
        .b(new_Jinkela_wire_830)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_0),
        .dout(new_Jinkela_wire_1)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(G27),
        .c(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_2)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_721),
        .dout(new_Jinkela_wire_722)
    );

    spl3L new_Jinkela_splitter_33 (
        .a(G25),
        .d(new_Jinkela_wire_338),
        .c(new_Jinkela_wire_339),
        .b(new_Jinkela_wire_340)
    );

    spl2 new_Jinkela_splitter_3 (
        .a(G41),
        .c(new_Jinkela_wire_33),
        .b(new_Jinkela_wire_38)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_215),
        .dout(new_Jinkela_wire_216)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_722),
        .dout(new_Jinkela_wire_723)
    );

    spl4L new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_2),
        .d(new_Jinkela_wire_3),
        .e(new_Jinkela_wire_4),
        .c(new_Jinkela_wire_5),
        .b(new_Jinkela_wire_6)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_190),
        .dout(new_Jinkela_wire_191)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    spl4L new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_38),
        .d(new_Jinkela_wire_39),
        .e(new_Jinkela_wire_40),
        .c(new_Jinkela_wire_41),
        .b(new_Jinkela_wire_42)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_245),
        .dout(new_Jinkela_wire_246)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_191),
        .dout(new_Jinkela_wire_192)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_25 (
        .din(G37),
        .dout(new_Jinkela_wire_43)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_216),
        .dout(new_Jinkela_wire_217)
    );

    spl2 new_Jinkela_splitter_68 (
        .a(new_Jinkela_wire_724),
        .c(new_Jinkela_wire_725),
        .b(new_Jinkela_wire_726)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(G21),
        .c(new_Jinkela_wire_45),
        .b(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_192),
        .dout(new_Jinkela_wire_193)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    spl4L new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_33),
        .d(new_Jinkela_wire_34),
        .e(new_Jinkela_wire_35),
        .c(new_Jinkela_wire_36),
        .b(new_Jinkela_wire_37)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    spl2 new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_431),
        .c(new_Jinkela_wire_432),
        .b(new_Jinkela_wire_433)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_530),
        .dout(new_Jinkela_wire_531)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(new_Jinkela_wire_1650),
        .dout(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_451),
        .dout(new_Jinkela_wire_452)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(new_Jinkela_wire_1651),
        .c(new_Jinkela_wire_1652),
        .b(new_Jinkela_wire_1653)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_453),
        .dout(new_Jinkela_wire_454)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    spl2 new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_986),
        .c(new_Jinkela_wire_987),
        .b(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_454),
        .dout(new_Jinkela_wire_455)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_1030),
        .dout(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    spl2 new_Jinkela_splitter_101 (
        .a(_181_),
        .c(new_Jinkela_wire_1062),
        .b(new_Jinkela_wire_1063)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(_095_),
        .c(new_Jinkela_wire_1066),
        .b(new_Jinkela_wire_1067)
    );

    spl4L new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_532),
        .d(new_Jinkela_wire_533),
        .e(new_Jinkela_wire_534),
        .c(new_Jinkela_wire_535),
        .b(new_Jinkela_wire_536)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(G2),
        .c(new_Jinkela_wire_627),
        .b(new_Jinkela_wire_629)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(new_Jinkela_wire_1063),
        .c(new_Jinkela_wire_1064),
        .b(new_Jinkela_wire_1065)
    );

    spl2 new_Jinkela_splitter_104 (
        .a(_272_),
        .c(new_Jinkela_wire_1068),
        .b(new_Jinkela_wire_1069)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_1011),
        .dout(new_Jinkela_wire_1012)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(_292_),
        .c(new_Jinkela_wire_1079),
        .b(new_Jinkela_wire_1080)
    );

    spl2 new_Jinkela_splitter_57 (
        .a(G31),
        .c(new_Jinkela_wire_596),
        .b(new_Jinkela_wire_598)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_1013),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_463),
        .c(new_Jinkela_wire_464),
        .b(new_Jinkela_wire_465)
    );

    spl2 new_Jinkela_splitter_106 (
        .a(_316_),
        .c(new_Jinkela_wire_1074),
        .b(new_Jinkela_wire_1075)
    );

    spl4L new_Jinkela_splitter_105 (
        .a(_069_),
        .d(new_Jinkela_wire_1070),
        .e(new_Jinkela_wire_1071),
        .c(new_Jinkela_wire_1072),
        .b(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_483),
        .dout(new_Jinkela_wire_484)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_1016),
        .dout(new_Jinkela_wire_1017)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_484),
        .dout(new_Jinkela_wire_485)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1076),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    spl2 new_Jinkela_splitter_95 (
        .a(new_Jinkela_wire_1017),
        .c(new_Jinkela_wire_1018),
        .b(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_485),
        .dout(new_Jinkela_wire_486)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_598),
        .d(new_Jinkela_wire_599),
        .e(new_Jinkela_wire_600),
        .c(new_Jinkela_wire_601),
        .b(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_486),
        .dout(new_Jinkela_wire_487)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_net_710),
        .dout(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_net_728),
        .dout(new_Jinkela_wire_1081)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    spl3L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_566),
        .d(new_Jinkela_wire_567),
        .c(new_Jinkela_wire_568),
        .b(new_Jinkela_wire_569)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_488),
        .dout(new_Jinkela_wire_489)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1039),
        .dout(new_Jinkela_wire_1040)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    or_bb _683_ (
        .a(new_Jinkela_wire_1523),
        .b(new_Jinkela_wire_1243),
        .c(_281_)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_1345),
        .dout(new_Jinkela_wire_1346)
    );

    or_ii _684_ (
        .a(new_Jinkela_wire_1116),
        .b(new_Jinkela_wire_107),
        .c(_282_)
    );

    spl2 new_Jinkela_splitter_177 (
        .a(new_Jinkela_wire_1319),
        .c(new_Jinkela_wire_1320),
        .b(new_Jinkela_wire_1321)
    );

    and_ii _685_ (
        .a(new_Jinkela_wire_1117),
        .b(new_Jinkela_wire_106),
        .c(_283_)
    );

    spl2 new_Jinkela_splitter_178 (
        .a(new_Jinkela_wire_1321),
        .c(new_Jinkela_wire_1322),
        .b(new_Jinkela_wire_1323)
    );

    and_bi _686_ (
        .a(_282_),
        .b(_283_),
        .c(new_net_698)
    );

    or_bb _687_ (
        .a(new_Jinkela_wire_1525),
        .b(new_Jinkela_wire_1573),
        .c(_284_)
    );

    spl2 new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_1323),
        .c(new_Jinkela_wire_1324),
        .b(new_Jinkela_wire_1325)
    );

    or_ii _688_ (
        .a(new_Jinkela_wire_1208),
        .b(new_Jinkela_wire_465),
        .c(_285_)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_Jinkela_wire_1346),
        .dout(new_Jinkela_wire_1347)
    );

    and_ii _689_ (
        .a(new_Jinkela_wire_1209),
        .b(new_Jinkela_wire_464),
        .c(_286_)
    );

    bfr new_Jinkela_buffer_876 (
        .din(new_Jinkela_wire_1347),
        .dout(new_Jinkela_wire_1348)
    );

    and_bi _690_ (
        .a(_285_),
        .b(_286_),
        .c(new_net_724)
    );

    spl4L new_Jinkela_splitter_190 (
        .a(_343_),
        .d(new_Jinkela_wire_1358),
        .e(new_Jinkela_wire_1359),
        .c(new_Jinkela_wire_1360),
        .b(new_Jinkela_wire_1361)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_net_688),
        .dout(new_Jinkela_wire_1357)
    );

    or_bi _691_ (
        .a(new_Jinkela_wire_1120),
        .b(new_Jinkela_wire_1407),
        .c(_287_)
    );

    spl2 new_Jinkela_splitter_191 (
        .a(_207_),
        .c(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_1363)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1351),
        .dout(new_Jinkela_wire_1352)
    );

    or_bb _692_ (
        .a(new_Jinkela_wire_1348),
        .b(new_Jinkela_wire_1590),
        .c(_288_)
    );

    or_bb _693_ (
        .a(new_Jinkela_wire_1191),
        .b(new_Jinkela_wire_1510),
        .c(_289_)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1352),
        .dout(new_Jinkela_wire_1353)
    );

    and_bi _694_ (
        .a(new_Jinkela_wire_1341),
        .b(new_Jinkela_wire_496),
        .c(_290_)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(_038_),
        .c(new_Jinkela_wire_1368),
        .b(new_Jinkela_wire_1369)
    );

    and_bi _695_ (
        .a(new_Jinkela_wire_497),
        .b(new_Jinkela_wire_1342),
        .c(_291_)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1394),
        .dout(new_Jinkela_wire_1395)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1353),
        .dout(new_Jinkela_wire_1354)
    );

    or_bb _696_ (
        .a(_291_),
        .b(_290_),
        .c(new_net_696)
    );

    or_bb _697_ (
        .a(new_Jinkela_wire_1192),
        .b(new_Jinkela_wire_1537),
        .c(_292_)
    );

    spl2 new_Jinkela_splitter_189 (
        .a(new_Jinkela_wire_1354),
        .c(new_Jinkela_wire_1355),
        .b(new_Jinkela_wire_1356)
    );

    or_ii _698_ (
        .a(new_Jinkela_wire_1079),
        .b(new_Jinkela_wire_855),
        .c(_293_)
    );

    and_ii _699_ (
        .a(new_Jinkela_wire_1080),
        .b(new_Jinkela_wire_854),
        .c(_294_)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_1363),
        .dout(new_Jinkela_wire_1364)
    );

    and_bi _700_ (
        .a(_293_),
        .b(_294_),
        .c(new_net_716)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(_078_),
        .c(new_Jinkela_wire_1370),
        .b(new_Jinkela_wire_1371)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1364),
        .dout(new_Jinkela_wire_1365)
    );

    or_bi _701_ (
        .a(new_Jinkela_wire_1193),
        .b(new_Jinkela_wire_1320),
        .c(_295_)
    );

    spl4L new_Jinkela_splitter_194 (
        .a(_047_),
        .d(new_Jinkela_wire_1372),
        .e(new_Jinkela_wire_1373),
        .c(new_Jinkela_wire_1374),
        .b(new_Jinkela_wire_1375)
    );

    and_bi _702_ (
        .a(new_Jinkela_wire_1212),
        .b(new_Jinkela_wire_953),
        .c(_296_)
    );

    spl2 new_Jinkela_splitter_200 (
        .a(_319_),
        .c(new_Jinkela_wire_1398),
        .b(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1365),
        .dout(new_Jinkela_wire_1366)
    );

    and_bi _703_ (
        .a(new_Jinkela_wire_952),
        .b(new_Jinkela_wire_1213),
        .c(_297_)
    );

    spl2 new_Jinkela_splitter_197 (
        .a(_239_),
        .c(new_Jinkela_wire_1390),
        .b(new_Jinkela_wire_1391)
    );

    or_bb _704_ (
        .a(_297_),
        .b(_296_),
        .c(new_net_714)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1366),
        .dout(new_Jinkela_wire_1367)
    );

    or_bi _705_ (
        .a(new_Jinkela_wire_1190),
        .b(new_Jinkela_wire_1606),
        .c(_298_)
    );

    and_bi _706_ (
        .a(new_Jinkela_wire_1175),
        .b(new_Jinkela_wire_432),
        .c(_299_)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(_306_),
        .c(new_Jinkela_wire_1392),
        .b(new_Jinkela_wire_1393)
    );

    and_bi _707_ (
        .a(new_Jinkela_wire_433),
        .b(new_Jinkela_wire_1176),
        .c(_300_)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1376),
        .dout(new_Jinkela_wire_1377)
    );

    or_bb _708_ (
        .a(_300_),
        .b(_299_),
        .c(new_net_722)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_net_716),
        .dout(new_Jinkela_wire_1394)
    );

    or_bb _709_ (
        .a(new_Jinkela_wire_1592),
        .b(new_Jinkela_wire_1168),
        .c(_301_)
    );

    spl2 new_Jinkela_splitter_199 (
        .a(_120_),
        .c(new_Jinkela_wire_1396),
        .b(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    or_bi _710_ (
        .a(_301_),
        .b(new_Jinkela_wire_1414),
        .c(_302_)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1375),
        .dout(new_Jinkela_wire_1376)
    );

    or_bb _711_ (
        .a(new_Jinkela_wire_1268),
        .b(new_Jinkela_wire_1512),
        .c(_303_)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_1378),
        .dout(new_Jinkela_wire_1379)
    );

    or_ii _712_ (
        .a(new_Jinkela_wire_1443),
        .b(new_Jinkela_wire_692),
        .c(_304_)
    );

    and_ii _713_ (
        .a(new_Jinkela_wire_1444),
        .b(new_Jinkela_wire_693),
        .c(_305_)
    );

    and_bi _714_ (
        .a(_304_),
        .b(_305_),
        .c(new_net_718)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1379),
        .dout(new_Jinkela_wire_1380)
    );

    or_bb _715_ (
        .a(new_Jinkela_wire_1267),
        .b(new_Jinkela_wire_1539),
        .c(_306_)
    );

    bfr new_Jinkela_buffer_897 (
        .din(_209_),
        .dout(new_Jinkela_wire_1400)
    );

    or_ii _716_ (
        .a(new_Jinkela_wire_1392),
        .b(new_Jinkela_wire_1052),
        .c(_307_)
    );

    spl2 new_Jinkela_splitter_202 (
        .a(_081_),
        .c(new_Jinkela_wire_1404),
        .b(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    and_ii _717_ (
        .a(new_Jinkela_wire_1393),
        .b(new_Jinkela_wire_1053),
        .c(_308_)
    );

    and_bi _718_ (
        .a(_307_),
        .b(_308_),
        .c(new_net_704)
    );

    bfr new_Jinkela_buffer_898 (
        .din(_337_),
        .dout(new_Jinkela_wire_1401)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    or_bi _719_ (
        .a(new_Jinkela_wire_1269),
        .b(new_Jinkela_wire_1322),
        .c(_309_)
    );

    spl3L new_Jinkela_splitter_203 (
        .a(_220_),
        .d(new_Jinkela_wire_1406),
        .c(new_Jinkela_wire_1407),
        .b(new_Jinkela_wire_1408)
    );

    or_ii _720_ (
        .a(new_Jinkela_wire_1454),
        .b(new_Jinkela_wire_988),
        .c(_310_)
    );

    spl2 new_Jinkela_splitter_201 (
        .a(new_Jinkela_wire_1401),
        .c(new_Jinkela_wire_1402),
        .b(new_Jinkela_wire_1403)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    and_ii _721_ (
        .a(new_Jinkela_wire_1455),
        .b(new_Jinkela_wire_987),
        .c(_311_)
    );

    and_bi _722_ (
        .a(_310_),
        .b(_311_),
        .c(new_net_726)
    );

    spl3L new_Jinkela_splitter_195 (
        .a(new_Jinkela_wire_1383),
        .d(new_Jinkela_wire_1384),
        .c(new_Jinkela_wire_1385),
        .b(new_Jinkela_wire_1386)
    );

    or_bi _723_ (
        .a(new_Jinkela_wire_1270),
        .b(new_Jinkela_wire_1608),
        .c(_312_)
    );

    bfr new_Jinkela_buffer_905 (
        .din(_211_),
        .dout(new_Jinkela_wire_1415)
    );

    or_ii _724_ (
        .a(new_Jinkela_wire_1139),
        .b(new_Jinkela_wire_886),
        .c(_313_)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_193),
        .dout(new_Jinkela_wire_194)
    );

    or_bi _515_ (
        .a(new_Jinkela_wire_601),
        .b(new_Jinkela_wire_994),
        .c(_129_)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    and_bi _516_ (
        .a(new_Jinkela_wire_600),
        .b(new_Jinkela_wire_992),
        .c(_130_)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_194),
        .dout(new_Jinkela_wire_195)
    );

    or_bi _517_ (
        .a(_130_),
        .b(_129_),
        .c(_131_)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_246),
        .dout(new_Jinkela_wire_247)
    );

    or_bi _518_ (
        .a(new_Jinkela_wire_1299),
        .b(new_Jinkela_wire_1330),
        .c(_132_)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_195),
        .dout(new_Jinkela_wire_196)
    );

    and_bi _519_ (
        .a(new_Jinkela_wire_1300),
        .b(new_Jinkela_wire_1331),
        .c(_133_)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    and_bi _520_ (
        .a(_132_),
        .b(_133_),
        .c(_134_)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_196),
        .dout(new_Jinkela_wire_197)
    );

    or_bb _521_ (
        .a(new_Jinkela_wire_1469),
        .b(new_Jinkela_wire_1265),
        .c(_135_)
    );

    and_bb _522_ (
        .a(new_Jinkela_wire_1471),
        .b(new_Jinkela_wire_1266),
        .c(_136_)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_276),
        .dout(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_197),
        .dout(new_Jinkela_wire_198)
    );

    or_bi _523_ (
        .a(_136_),
        .b(_135_),
        .c(_137_)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    or_bb _524_ (
        .a(new_Jinkela_wire_792),
        .b(new_Jinkela_wire_338),
        .c(_138_)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    and_bb _525_ (
        .a(new_Jinkela_wire_793),
        .b(new_Jinkela_wire_339),
        .c(_139_)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_247),
        .dout(new_Jinkela_wire_248)
    );

    and_bi _526_ (
        .a(_138_),
        .b(_139_),
        .c(_140_)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_199),
        .dout(new_Jinkela_wire_200)
    );

    or_bi _527_ (
        .a(new_Jinkela_wire_3),
        .b(new_Jinkela_wire_567),
        .c(_141_)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    and_bi _528_ (
        .a(new_Jinkela_wire_4),
        .b(new_Jinkela_wire_568),
        .c(_142_)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    or_bi _529_ (
        .a(_142_),
        .b(_141_),
        .c(_143_)
    );

    spl3L new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_273),
        .d(new_Jinkela_wire_274),
        .c(new_Jinkela_wire_275),
        .b(new_Jinkela_wire_276)
    );

    or_bi _530_ (
        .a(new_Jinkela_wire_1626),
        .b(new_Jinkela_wire_1445),
        .c(_144_)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    and_bi _531_ (
        .a(new_Jinkela_wire_1627),
        .b(new_Jinkela_wire_1446),
        .c(_145_)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_221),
        .dout(new_Jinkela_wire_222)
    );

    and_bi _532_ (
        .a(_144_),
        .b(_145_),
        .c(_146_)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_202),
        .c(new_Jinkela_wire_203),
        .b(new_Jinkela_wire_204)
    );

    or_bb _533_ (
        .a(new_Jinkela_wire_923),
        .b(new_Jinkela_wire_630),
        .c(_147_)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_222),
        .dout(new_Jinkela_wire_223)
    );

    and_bb _534_ (
        .a(new_Jinkela_wire_926),
        .b(new_Jinkela_wire_628),
        .c(_148_)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_248),
        .dout(new_Jinkela_wire_249)
    );

    and_bi _535_ (
        .a(_147_),
        .b(_148_),
        .c(_149_)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    or_bi _536_ (
        .a(new_Jinkela_wire_534),
        .b(new_Jinkela_wire_957),
        .c(_150_)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    and_bi _537_ (
        .a(new_Jinkela_wire_535),
        .b(new_Jinkela_wire_959),
        .c(_151_)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    and_bi _538_ (
        .a(_150_),
        .b(_151_),
        .c(_152_)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    or_bi _539_ (
        .a(new_Jinkela_wire_1198),
        .b(new_Jinkela_wire_1177),
        .c(_153_)
    );

    and_bi _540_ (
        .a(new_Jinkela_wire_1199),
        .b(new_Jinkela_wire_1178),
        .c(_154_)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    or_bi _541_ (
        .a(_154_),
        .b(_153_),
        .c(_155_)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    or_bb _542_ (
        .a(new_Jinkela_wire_1339),
        .b(new_Jinkela_wire_1486),
        .c(_156_)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_226),
        .dout(new_Jinkela_wire_227)
    );

    and_bb _543_ (
        .a(new_Jinkela_wire_1340),
        .b(new_Jinkela_wire_1485),
        .c(_157_)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    and_bi _544_ (
        .a(_156_),
        .b(_157_),
        .c(_158_)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    and_bi _545_ (
        .a(new_Jinkela_wire_1297),
        .b(new_Jinkela_wire_1448),
        .c(_159_)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_251),
        .dout(new_Jinkela_wire_252)
    );

    and_bi _546_ (
        .a(new_Jinkela_wire_1449),
        .b(new_Jinkela_wire_1298),
        .c(_160_)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    or_bb _547_ (
        .a(_160_),
        .b(_159_),
        .c(_161_)
    );

    spl2 new_Jinkela_splitter_39 (
        .a(G13),
        .c(new_Jinkela_wire_402),
        .b(new_Jinkela_wire_404)
    );

    or_bi _548_ (
        .a(new_Jinkela_wire_1595),
        .b(new_Jinkela_wire_1309),
        .c(_162_)
    );

    spl3L new_Jinkela_splitter_36 (
        .a(G19),
        .d(new_Jinkela_wire_370),
        .c(new_Jinkela_wire_371),
        .b(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    or_ii _549_ (
        .a(new_Jinkela_wire_1021),
        .b(new_Jinkela_wire_39),
        .c(_163_)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    and_bi _550_ (
        .a(new_Jinkela_wire_1621),
        .b(new_Jinkela_wire_1361),
        .c(_164_)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    and_bi _551_ (
        .a(new_Jinkela_wire_1358),
        .b(new_Jinkela_wire_1622),
        .c(_165_)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_278),
        .dout(new_Jinkela_wire_279)
    );

    or_bb _552_ (
        .a(_165_),
        .b(_164_),
        .c(_166_)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_231),
        .dout(new_Jinkela_wire_232)
    );

    or_bi _553_ (
        .a(new_Jinkela_wire_828),
        .b(new_Jinkela_wire_1026),
        .c(_167_)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_253),
        .dout(new_Jinkela_wire_254)
    );

    and_bi _554_ (
        .a(new_Jinkela_wire_827),
        .b(new_Jinkela_wire_1025),
        .c(_168_)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_232),
        .dout(new_Jinkela_wire_233)
    );

    or_bi _555_ (
        .a(_168_),
        .b(_167_),
        .c(_169_)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_310),
        .dout(new_Jinkela_wire_311)
    );

    or_bb _556_ (
        .a(new_Jinkela_wire_206),
        .b(new_Jinkela_wire_271),
        .c(_170_)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    spl4L new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_890),
        .d(new_Jinkela_wire_891),
        .e(new_Jinkela_wire_892),
        .c(new_Jinkela_wire_893),
        .b(new_Jinkela_wire_894)
    );

    spl2 new_Jinkela_splitter_87 (
        .a(G14),
        .c(new_Jinkela_wire_922),
        .b(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_770),
        .dout(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    spl2 new_Jinkela_splitter_84 (
        .a(G8),
        .c(new_Jinkela_wire_888),
        .b(new_Jinkela_wire_890)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_773),
        .dout(new_Jinkela_wire_774)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_755),
        .c(new_Jinkela_wire_756),
        .b(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_830),
        .dout(new_Jinkela_wire_831)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_775),
        .dout(new_Jinkela_wire_776)
    );

    spl4L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_924),
        .d(new_Jinkela_wire_925),
        .e(new_Jinkela_wire_926),
        .c(new_Jinkela_wire_927),
        .b(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_776),
        .dout(new_Jinkela_wire_777)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_777),
        .dout(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_831),
        .dout(new_Jinkela_wire_832)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_778),
        .dout(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_803),
        .dout(new_Jinkela_wire_804)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_779),
        .dout(new_Jinkela_wire_780)
    );

    spl3L new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_858),
        .d(new_Jinkela_wire_859),
        .c(new_Jinkela_wire_860),
        .b(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_804),
        .dout(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_832),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1386),
        .dout(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_908 (
        .din(_334_),
        .dout(new_Jinkela_wire_1418)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(new_Jinkela_wire_1387),
        .c(new_Jinkela_wire_1388),
        .b(new_Jinkela_wire_1389)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(_236_),
        .c(new_Jinkela_wire_1424),
        .b(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1410),
        .dout(new_Jinkela_wire_1411)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(_358_),
        .c(new_Jinkela_wire_1426),
        .b(new_Jinkela_wire_1427)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1411),
        .dout(new_Jinkela_wire_1412)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1412),
        .dout(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1413),
        .dout(new_Jinkela_wire_1414)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(_162_),
        .c(new_Jinkela_wire_1428),
        .b(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_net_724),
        .dout(new_Jinkela_wire_1437)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(new_Jinkela_wire_1421),
        .c(new_Jinkela_wire_1422),
        .b(new_Jinkela_wire_1423)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(_175_),
        .c(new_Jinkela_wire_1441),
        .b(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_net_706),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(_303_),
        .c(new_Jinkela_wire_1443),
        .b(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1438),
        .dout(new_Jinkela_wire_1439)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_net_684),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1439),
        .dout(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(_143_),
        .c(new_Jinkela_wire_1445),
        .b(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1435),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_net_700),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_net_718),
        .dout(new_Jinkela_wire_1450)
    );

    spl2 new_Jinkela_splitter_211 (
        .a(_137_),
        .c(new_Jinkela_wire_1448),
        .b(new_Jinkela_wire_1449)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(_023_),
        .c(new_Jinkela_wire_1456),
        .b(new_Jinkela_wire_1457)
    );

    spl2 new_Jinkela_splitter_212 (
        .a(_192_),
        .c(new_Jinkela_wire_1451),
        .b(new_Jinkela_wire_1452)
    );

    spl2 new_Jinkela_splitter_213 (
        .a(_309_),
        .c(new_Jinkela_wire_1454),
        .b(new_Jinkela_wire_1455)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(_346_),
        .c(new_Jinkela_wire_1458),
        .b(new_Jinkela_wire_1459)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(_063_),
        .c(new_Jinkela_wire_1466),
        .b(new_Jinkela_wire_1467)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(_204_),
        .c(new_Jinkela_wire_1460),
        .b(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_489),
        .dout(new_Jinkela_wire_490)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1040),
        .dout(new_Jinkela_wire_1041)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_537),
        .dout(new_Jinkela_wire_538)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_490),
        .dout(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1041),
        .dout(new_Jinkela_wire_1042)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(_122_),
        .c(new_Jinkela_wire_1084),
        .b(new_Jinkela_wire_1085)
    );

    spl2 new_Jinkela_splitter_109 (
        .a(_089_),
        .c(new_Jinkela_wire_1086),
        .b(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1042),
        .dout(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_596),
        .dout(new_Jinkela_wire_597)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_492),
        .dout(new_Jinkela_wire_493)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_493),
        .dout(new_Jinkela_wire_494)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1044),
        .dout(new_Jinkela_wire_1045)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_494),
        .dout(new_Jinkela_wire_495)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1045),
        .dout(new_Jinkela_wire_1046)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_513),
        .dout(new_Jinkela_wire_514)
    );

    spl2 new_Jinkela_splitter_110 (
        .a(_328_),
        .c(new_Jinkela_wire_1088),
        .b(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1090),
        .dout(new_Jinkela_wire_1091)
    );

    spl2 new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_495),
        .c(new_Jinkela_wire_496),
        .b(new_Jinkela_wire_497)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1046),
        .dout(new_Jinkela_wire_1047)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_514),
        .dout(new_Jinkela_wire_515)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_net_712),
        .dout(new_Jinkela_wire_1090)
    );

    bfr new_Jinkela_buffer_801 (
        .din(_212_),
        .dout(new_Jinkela_wire_1095)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1047),
        .dout(new_Jinkela_wire_1048)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_539),
        .dout(new_Jinkela_wire_540)
    );

    spl2 new_Jinkela_splitter_111 (
        .a(_322_),
        .c(new_Jinkela_wire_1093),
        .b(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_515),
        .dout(new_Jinkela_wire_516)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1048),
        .dout(new_Jinkela_wire_1049)
    );

    spl4L new_Jinkela_splitter_113 (
        .a(_265_),
        .d(new_Jinkela_wire_1098),
        .e(new_Jinkela_wire_1099),
        .c(new_Jinkela_wire_1100),
        .b(new_Jinkela_wire_1101)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(G12),
        .c(new_Jinkela_wire_661),
        .b(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1049),
        .dout(new_Jinkela_wire_1050)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_540),
        .dout(new_Jinkela_wire_541)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1091),
        .dout(new_Jinkela_wire_1092)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1050),
        .dout(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(new_Jinkela_wire_1051),
        .c(new_Jinkela_wire_1052),
        .b(new_Jinkela_wire_1053)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_net_722),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_519),
        .dout(new_Jinkela_wire_520)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(_053_),
        .c(new_Jinkela_wire_1096),
        .b(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_net_708),
        .dout(new_Jinkela_wire_1102)
    );

    spl3L new_Jinkela_splitter_115 (
        .a(_228_),
        .d(new_Jinkela_wire_1107),
        .c(new_Jinkela_wire_1108),
        .b(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_520),
        .dout(new_Jinkela_wire_521)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(_007_),
        .c(new_Jinkela_wire_1105),
        .b(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_521),
        .dout(new_Jinkela_wire_522)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_522),
        .dout(new_Jinkela_wire_523)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_net_694),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_810 (
        .din(_227_),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_523),
        .dout(new_Jinkela_wire_524)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_663),
        .d(new_Jinkela_wire_664),
        .e(new_Jinkela_wire_665),
        .c(new_Jinkela_wire_666),
        .b(new_Jinkela_wire_667)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_524),
        .dout(new_Jinkela_wire_525)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(_281_),
        .c(new_Jinkela_wire_1116),
        .b(new_Jinkela_wire_1117)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_525),
        .c(new_Jinkela_wire_526),
        .b(new_Jinkela_wire_527)
    );

    spl2 new_Jinkela_splitter_117 (
        .a(_224_),
        .c(new_Jinkela_wire_1118),
        .b(new_Jinkela_wire_1119)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(new_Jinkela_wire_1119),
        .c(new_Jinkela_wire_1120),
        .b(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    spl2 new_Jinkela_splitter_119 (
        .a(_072_),
        .c(new_Jinkela_wire_1129),
        .b(new_Jinkela_wire_1130)
    );

    spl2 new_Jinkela_splitter_120 (
        .a(_044_),
        .c(new_Jinkela_wire_1131),
        .b(new_Jinkela_wire_1132)
    );

    spl4L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_629),
        .d(new_Jinkela_wire_630),
        .e(new_Jinkela_wire_631),
        .c(new_Jinkela_wire_632),
        .b(new_Jinkela_wire_633)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(_349_),
        .c(new_Jinkela_wire_1133),
        .b(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_546),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_233),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_254),
        .dout(new_Jinkela_wire_255)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_279),
        .dout(new_Jinkela_wire_280)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(new_Jinkela_wire_235),
        .c(new_Jinkela_wire_236),
        .b(new_Jinkela_wire_237)
    );

    spl3L new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_340),
        .d(new_Jinkela_wire_341),
        .c(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_255),
        .dout(new_Jinkela_wire_256)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_256),
        .dout(new_Jinkela_wire_257)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_280),
        .dout(new_Jinkela_wire_281)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_257),
        .dout(new_Jinkela_wire_258)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_258),
        .dout(new_Jinkela_wire_259)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_281),
        .dout(new_Jinkela_wire_282)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_259),
        .dout(new_Jinkela_wire_260)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_311),
        .dout(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_282),
        .dout(new_Jinkela_wire_283)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_343),
        .dout(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_283),
        .dout(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_263),
        .dout(new_Jinkela_wire_264)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    spl2 new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_266),
        .c(new_Jinkela_wire_267),
        .b(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_313),
        .dout(new_Jinkela_wire_314)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    spl3L new_Jinkela_splitter_42 (
        .a(G17),
        .d(new_Jinkela_wire_434),
        .c(new_Jinkela_wire_435),
        .b(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_314),
        .dout(new_Jinkela_wire_315)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_315),
        .dout(new_Jinkela_wire_316)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_290),
        .dout(new_Jinkela_wire_291)
    );

    spl4L new_Jinkela_splitter_40 (
        .a(new_Jinkela_wire_404),
        .d(new_Jinkela_wire_405),
        .e(new_Jinkela_wire_406),
        .c(new_Jinkela_wire_407),
        .b(new_Jinkela_wire_408)
    );

    spl3L new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_372),
        .d(new_Jinkela_wire_373),
        .c(new_Jinkela_wire_374),
        .b(new_Jinkela_wire_375)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_316),
        .dout(new_Jinkela_wire_317)
    );

    and_ii _725_ (
        .a(new_Jinkela_wire_1140),
        .b(new_Jinkela_wire_887),
        .c(_314_)
    );

    and_bi _726_ (
        .a(_313_),
        .b(_314_),
        .c(new_net_692)
    );

    or_bb _727_ (
        .a(new_Jinkela_wire_1128),
        .b(new_Jinkela_wire_1275),
        .c(_315_)
    );

    or_bb _728_ (
        .a(new_Jinkela_wire_1639),
        .b(new_Jinkela_wire_1515),
        .c(_316_)
    );

    or_ii _729_ (
        .a(new_Jinkela_wire_1074),
        .b(new_Jinkela_wire_920),
        .c(_317_)
    );

    and_ii _730_ (
        .a(new_Jinkela_wire_1075),
        .b(new_Jinkela_wire_921),
        .c(_318_)
    );

    and_bi _731_ (
        .a(_317_),
        .b(_318_),
        .c(G1331)
    );

    or_bb _732_ (
        .a(new_Jinkela_wire_1638),
        .b(new_Jinkela_wire_1542),
        .c(_319_)
    );

    or_ii _733_ (
        .a(new_Jinkela_wire_1398),
        .b(new_Jinkela_wire_302),
        .c(_320_)
    );

    and_ii _734_ (
        .a(new_Jinkela_wire_1399),
        .b(new_Jinkela_wire_303),
        .c(_321_)
    );

    and_bi _735_ (
        .a(_320_),
        .b(_321_),
        .c(G1330)
    );

    or_bi _736_ (
        .a(new_Jinkela_wire_1641),
        .b(new_Jinkela_wire_1325),
        .c(_322_)
    );

    or_ii _737_ (
        .a(new_Jinkela_wire_1093),
        .b(new_Jinkela_wire_562),
        .c(_323_)
    );

    and_ii _738_ (
        .a(new_Jinkela_wire_1094),
        .b(new_Jinkela_wire_563),
        .c(_324_)
    );

    and_bi _739_ (
        .a(_323_),
        .b(_324_),
        .c(G1329)
    );

    or_bi _740_ (
        .a(new_Jinkela_wire_1640),
        .b(new_Jinkela_wire_1610),
        .c(_325_)
    );

    or_ii _741_ (
        .a(new_Jinkela_wire_1202),
        .b(new_Jinkela_wire_790),
        .c(_326_)
    );

    and_ii _742_ (
        .a(new_Jinkela_wire_1203),
        .b(new_Jinkela_wire_791),
        .c(_327_)
    );

    and_bi _743_ (
        .a(_326_),
        .b(_327_),
        .c(G1328)
    );

    or_bb _744_ (
        .a(new_Jinkela_wire_1196),
        .b(new_Jinkela_wire_1514),
        .c(_328_)
    );

    or_ii _745_ (
        .a(new_Jinkela_wire_1088),
        .b(new_Jinkela_wire_203),
        .c(_329_)
    );

    and_ii _746_ (
        .a(new_Jinkela_wire_1089),
        .b(new_Jinkela_wire_204),
        .c(_330_)
    );

    and_bi _747_ (
        .a(_329_),
        .b(_330_),
        .c(G1327)
    );

    or_bb _748_ (
        .a(new_Jinkela_wire_1197),
        .b(new_Jinkela_wire_1541),
        .c(_331_)
    );

    or_ii _749_ (
        .a(new_Jinkela_wire_1516),
        .b(new_Jinkela_wire_236),
        .c(_332_)
    );

    and_ii _750_ (
        .a(new_Jinkela_wire_1517),
        .b(new_Jinkela_wire_237),
        .c(_333_)
    );

    and_bi _751_ (
        .a(_332_),
        .b(_333_),
        .c(G1326)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_785),
        .dout(new_Jinkela_wire_786)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_787),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_789),
        .c(new_Jinkela_wire_790),
        .b(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_835),
        .dout(new_Jinkela_wire_836)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_712 (
        .din(G34),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_836),
        .dout(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_837),
        .dout(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_888),
        .dout(new_Jinkela_wire_889)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_838),
        .dout(new_Jinkela_wire_839)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    spl2 new_Jinkela_splitter_90 (
        .a(G10),
        .c(new_Jinkela_wire_956),
        .b(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_840),
        .dout(new_Jinkela_wire_841)
    );

    spl2 new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_821),
        .c(new_Jinkela_wire_822),
        .b(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_841),
        .dout(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    and_bb _406_ (
        .a(new_Jinkela_wire_270),
        .b(new_Jinkela_wire_41),
        .c(_020_)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_842),
        .dout(new_Jinkela_wire_843)
    );

    and_bb _557_ (
        .a(new_Jinkela_wire_205),
        .b(new_Jinkela_wire_272),
        .c(_171_)
    );

    or_bi _558_ (
        .a(_171_),
        .b(_170_),
        .c(_172_)
    );

    or_bi _559_ (
        .a(new_Jinkela_wire_1185),
        .b(new_Jinkela_wire_1225),
        .c(_173_)
    );

    and_bi _560_ (
        .a(new_Jinkela_wire_1186),
        .b(new_Jinkela_wire_1226),
        .c(_174_)
    );

    and_bi _561_ (
        .a(_173_),
        .b(_174_),
        .c(_175_)
    );

    and_bi _562_ (
        .a(new_Jinkela_wire_1441),
        .b(new_Jinkela_wire_1488),
        .c(_176_)
    );

    and_bi _563_ (
        .a(new_Jinkela_wire_1487),
        .b(new_Jinkela_wire_1442),
        .c(_177_)
    );

    or_bb _564_ (
        .a(_177_),
        .b(_176_),
        .c(_178_)
    );

    or_bb _565_ (
        .a(new_Jinkela_wire_1285),
        .b(new_Jinkela_wire_1245),
        .c(_179_)
    );

    and_bb _566_ (
        .a(new_Jinkela_wire_1286),
        .b(new_Jinkela_wire_1246),
        .c(_180_)
    );

    or_bi _567_ (
        .a(new_Jinkela_wire_1305),
        .b(new_Jinkela_wire_1328),
        .c(_181_)
    );

    or_bb _568_ (
        .a(new_Jinkela_wire_1064),
        .b(new_Jinkela_wire_1428),
        .c(_182_)
    );

    or_bi _569_ (
        .a(new_Jinkela_wire_1308),
        .b(new_Jinkela_wire_1593),
        .c(_183_)
    );

    or_bb _570_ (
        .a(new_Jinkela_wire_1472),
        .b(new_Jinkela_wire_1065),
        .c(_184_)
    );

    and_bb _571_ (
        .a(new_Jinkela_wire_1646),
        .b(new_Jinkela_wire_1255),
        .c(_185_)
    );

    or_ii _572_ (
        .a(new_Jinkela_wire_529),
        .b(new_Jinkela_wire_37),
        .c(_186_)
    );

    and_bi _573_ (
        .a(new_Jinkela_wire_1493),
        .b(new_Jinkela_wire_1290),
        .c(_187_)
    );

    or_bi _385_ (
        .a(new_Jinkela_wire_860),
        .b(new_Jinkela_wire_309),
        .c(_359_)
    );

    and_bi _574_ (
        .a(new_Jinkela_wire_1289),
        .b(new_Jinkela_wire_1494),
        .c(_188_)
    );

    and_bi _363_ (
        .a(_335_),
        .b(_336_),
        .c(_337_)
    );

    or_bb _361_ (
        .a(new_Jinkela_wire_371),
        .b(new_Jinkela_wire_434),
        .c(_335_)
    );

    or_bb _575_ (
        .a(_188_),
        .b(_187_),
        .c(_189_)
    );

    and_bb _362_ (
        .a(new_Jinkela_wire_370),
        .b(new_Jinkela_wire_435),
        .c(_336_)
    );

    or_bi _576_ (
        .a(new_Jinkela_wire_176),
        .b(new_Jinkela_wire_665),
        .c(_190_)
    );

    and_bb _360_ (
        .a(new_Jinkela_wire_40),
        .b(new_Jinkela_wire_140),
        .c(_334_)
    );

    and_bi _577_ (
        .a(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_662),
        .c(_191_)
    );

    or_bi _364_ (
        .a(new_Jinkela_wire_79),
        .b(new_Jinkela_wire_698),
        .c(_338_)
    );

    or_bi _578_ (
        .a(_191_),
        .b(_190_),
        .c(_192_)
    );

    and_bi _368_ (
        .a(new_Jinkela_wire_1403),
        .b(new_Jinkela_wire_1180),
        .c(_342_)
    );

    or_bb _579_ (
        .a(new_Jinkela_wire_892),
        .b(new_Jinkela_wire_469),
        .c(_193_)
    );

    or_bi _367_ (
        .a(new_Jinkela_wire_1402),
        .b(new_Jinkela_wire_1179),
        .c(_341_)
    );

    and_bb _580_ (
        .a(new_Jinkela_wire_891),
        .b(new_Jinkela_wire_467),
        .c(_194_)
    );

    and_bi _365_ (
        .a(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_695),
        .c(_339_)
    );

    or_bi _581_ (
        .a(_194_),
        .b(_193_),
        .c(_195_)
    );

    and_bi _377_ (
        .a(new_Jinkela_wire_112),
        .b(new_Jinkela_wire_50),
        .c(_351_)
    );

    or_bi _582_ (
        .a(new_Jinkela_wire_1451),
        .b(new_Jinkela_wire_1216),
        .c(_196_)
    );

    or_bi _366_ (
        .a(_339_),
        .b(_338_),
        .c(_340_)
    );

    and_bi _369_ (
        .a(_341_),
        .b(_342_),
        .c(_343_)
    );

    and_bi _583_ (
        .a(new_Jinkela_wire_1452),
        .b(new_Jinkela_wire_1217),
        .c(_197_)
    );

    or_bb _370_ (
        .a(new_Jinkela_wire_1359),
        .b(new_Jinkela_wire_1422),
        .c(_344_)
    );

    and_bi _584_ (
        .a(_196_),
        .b(_197_),
        .c(_198_)
    );

    and_bb _371_ (
        .a(new_Jinkela_wire_1360),
        .b(new_Jinkela_wire_1423),
        .c(_345_)
    );

    and_bi _585_ (
        .a(new_Jinkela_wire_1519),
        .b(new_Jinkela_wire_1470),
        .c(_199_)
    );

    or_bi _372_ (
        .a(_345_),
        .b(_344_),
        .c(_346_)
    );

    and_bi _586_ (
        .a(new_Jinkela_wire_1468),
        .b(new_Jinkela_wire_1520),
        .c(_200_)
    );

    or_bb _373_ (
        .a(new_Jinkela_wire_241),
        .b(new_Jinkela_wire_502),
        .c(_347_)
    );

    or_bb _587_ (
        .a(_200_),
        .b(_199_),
        .c(_201_)
    );

    and_bb _374_ (
        .a(new_Jinkela_wire_239),
        .b(new_Jinkela_wire_501),
        .c(_348_)
    );

    or_bb _588_ (
        .a(new_Jinkela_wire_1576),
        .b(new_Jinkela_wire_1496),
        .c(_202_)
    );

    and_bi _375_ (
        .a(_347_),
        .b(_348_),
        .c(_349_)
    );

    and_bb _589_ (
        .a(new_Jinkela_wire_1577),
        .b(new_Jinkela_wire_1497),
        .c(_203_)
    );

    or_bi _376_ (
        .a(new_Jinkela_wire_113),
        .b(new_Jinkela_wire_49),
        .c(_350_)
    );

    or_bi _590_ (
        .a(new_Jinkela_wire_1588),
        .b(new_Jinkela_wire_1259),
        .c(_204_)
    );

    or_bb _591_ (
        .a(new_Jinkela_wire_1465),
        .b(_185_),
        .c(_205_)
    );

    or_bi _378_ (
        .a(_351_),
        .b(_350_),
        .c(_352_)
    );

    and_bi _592_ (
        .a(new_Jinkela_wire_1329),
        .b(new_Jinkela_wire_1306),
        .c(_206_)
    );

    or_bi _379_ (
        .a(new_Jinkela_wire_1133),
        .b(new_Jinkela_wire_1183),
        .c(_353_)
    );

    or_bb _593_ (
        .a(new_Jinkela_wire_1460),
        .b(new_Jinkela_wire_1527),
        .c(_207_)
    );

    and_bi _380_ (
        .a(new_Jinkela_wire_1134),
        .b(new_Jinkela_wire_1184),
        .c(_354_)
    );

    and_bi _594_ (
        .a(new_Jinkela_wire_1260),
        .b(new_Jinkela_wire_1589),
        .c(_208_)
    );

    and_bi _381_ (
        .a(_353_),
        .b(_354_),
        .c(_355_)
    );

    or_bb _595_ (
        .a(new_Jinkela_wire_1498),
        .b(new_Jinkela_wire_1062),
        .c(_209_)
    );

    or_bb _382_ (
        .a(new_Jinkela_wire_763),
        .b(new_Jinkela_wire_405),
        .c(_356_)
    );

    or_ii _596_ (
        .a(new_Jinkela_wire_1400),
        .b(new_Jinkela_wire_1362),
        .c(_210_)
    );

    and_bb _383_ (
        .a(new_Jinkela_wire_759),
        .b(new_Jinkela_wire_403),
        .c(_357_)
    );

    or_bb _597_ (
        .a(new_Jinkela_wire_1307),
        .b(new_Jinkela_wire_1594),
        .c(_211_)
    );

    and_bi _384_ (
        .a(_356_),
        .b(_357_),
        .c(_358_)
    );

    and_bi _598_ (
        .a(_210_),
        .b(new_Jinkela_wire_1417),
        .c(_212_)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    spl3L new_Jinkela_splitter_9 (
        .a(G18),
        .d(new_Jinkela_wire_76),
        .c(new_Jinkela_wire_77),
        .b(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    spl4L new_Jinkela_splitter_218 (
        .a(_134_),
        .d(new_Jinkela_wire_1468),
        .e(new_Jinkela_wire_1469),
        .c(new_Jinkela_wire_1470),
        .b(new_Jinkela_wire_1471)
    );

    spl2 new_Jinkela_splitter_221 (
        .a(_041_),
        .c(new_Jinkela_wire_1483),
        .b(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_43),
        .dout(new_Jinkela_wire_44)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(_066_),
        .c(new_Jinkela_wire_1481),
        .b(new_Jinkela_wire_1482)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(G24),
        .c(new_Jinkela_wire_108),
        .b(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    spl2 new_Jinkela_splitter_219 (
        .a(_183_),
        .c(new_Jinkela_wire_1472),
        .b(new_Jinkela_wire_1473)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_10),
        .dout(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    spl4L new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_47),
        .d(new_Jinkela_wire_48),
        .e(new_Jinkela_wire_49),
        .c(new_Jinkela_wire_50),
        .b(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_97 (
        .din(G33),
        .dout(new_Jinkela_wire_139)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1473),
        .dout(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1474),
        .dout(new_Jinkela_wire_1475)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    spl4L new_Jinkela_splitter_222 (
        .a(_146_),
        .d(new_Jinkela_wire_1485),
        .e(new_Jinkela_wire_1486),
        .c(new_Jinkela_wire_1487),
        .b(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_net_704),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1475),
        .dout(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    bfr new_Jinkela_buffer_937 (
        .din(_186_),
        .dout(new_Jinkela_wire_1489)
    );

    spl4L new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_110),
        .d(new_Jinkela_wire_111),
        .e(new_Jinkela_wire_112),
        .c(new_Jinkela_wire_113),
        .b(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1476),
        .dout(new_Jinkela_wire_1477)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(G4),
        .c(new_Jinkela_wire_171),
        .b(new_Jinkela_wire_173)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(_189_),
        .c(new_Jinkela_wire_1496),
        .b(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(_208_),
        .c(new_Jinkela_wire_1498),
        .b(new_Jinkela_wire_1499)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1479),
        .dout(new_Jinkela_wire_1480)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_18),
        .dout(new_Jinkela_wire_19)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_19),
        .dout(new_Jinkela_wire_20)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1491),
        .dout(new_Jinkela_wire_1492)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_108),
        .dout(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_20),
        .dout(new_Jinkela_wire_21)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(new_Jinkela_wire_1492),
        .c(new_Jinkela_wire_1493),
        .b(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(_101_),
        .c(new_Jinkela_wire_1521),
        .b(new_Jinkela_wire_1522)
    );

    spl2 new_Jinkela_splitter_230 (
        .a(_331_),
        .c(new_Jinkela_wire_1516),
        .b(new_Jinkela_wire_1517)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1499),
        .dout(new_Jinkela_wire_1500)
    );

    spl3L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_78),
        .d(new_Jinkela_wire_79),
        .c(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1500),
        .dout(new_Jinkela_wire_1501)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_55),
        .dout(new_Jinkela_wire_56)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1504),
        .dout(new_Jinkela_wire_1505)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    spl4L new_Jinkela_splitter_233 (
        .a(_230_),
        .d(new_Jinkela_wire_1523),
        .e(new_Jinkela_wire_1524),
        .c(new_Jinkela_wire_1525),
        .b(new_Jinkela_wire_1526)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_23),
        .dout(new_Jinkela_wire_24)
    );

    spl3L new_Jinkela_splitter_226 (
        .a(new_Jinkela_wire_1501),
        .d(new_Jinkela_wire_1502),
        .c(new_Jinkela_wire_1503),
        .b(new_Jinkela_wire_1504)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_net_690),
        .dout(new_Jinkela_wire_1518)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_24),
        .dout(new_Jinkela_wire_25)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(_198_),
        .c(new_Jinkela_wire_1519),
        .b(new_Jinkela_wire_1520)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_56),
        .dout(new_Jinkela_wire_57)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(_206_),
        .c(new_Jinkela_wire_1527),
        .b(new_Jinkela_wire_1528)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_25),
        .dout(new_Jinkela_wire_26)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1505),
        .dout(new_Jinkela_wire_1506)
    );

    spl3L new_Jinkela_splitter_15 (
        .a(G30),
        .d(new_Jinkela_wire_141),
        .c(new_Jinkela_wire_142),
        .b(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_958 (
        .din(_105_),
        .dout(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(_248_),
        .c(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1506),
        .dout(new_Jinkela_wire_1507)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1528),
        .dout(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    spl2 new_Jinkela_splitter_238 (
        .a(_098_),
        .c(new_Jinkela_wire_1543),
        .b(new_Jinkela_wire_1544)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_net_720),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_547),
        .dout(new_Jinkela_wire_548)
    );

    and_bi _386_ (
        .a(new_Jinkela_wire_859),
        .b(new_Jinkela_wire_307),
        .c(_000_)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_633),
        .dout(new_Jinkela_wire_634)
    );

    and_bi _387_ (
        .a(_359_),
        .b(_000_),
        .c(_001_)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    or_bi _388_ (
        .a(new_Jinkela_wire_1426),
        .b(new_Jinkela_wire_1301),
        .c(_002_)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_574),
        .dout(new_Jinkela_wire_575)
    );

    and_bi _389_ (
        .a(new_Jinkela_wire_1427),
        .b(new_Jinkela_wire_1302),
        .c(_003_)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    or_bi _390_ (
        .a(_003_),
        .b(_002_),
        .c(_004_)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    or_bb _391_ (
        .a(new_Jinkela_wire_1303),
        .b(new_Jinkela_wire_1288),
        .c(_005_)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    and_bb _392_ (
        .a(new_Jinkela_wire_1304),
        .b(new_Jinkela_wire_1287),
        .c(_006_)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    and_bi _393_ (
        .a(_005_),
        .b(_006_),
        .c(_007_)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_551),
        .dout(new_Jinkela_wire_552)
    );

    and_bi _394_ (
        .a(new_Jinkela_wire_1105),
        .b(new_Jinkela_wire_1458),
        .c(_008_)
    );

    spl2 new_Jinkela_splitter_66 (
        .a(G20),
        .c(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_696)
    );

    and_bi _395_ (
        .a(new_Jinkela_wire_1459),
        .b(new_Jinkela_wire_1106),
        .c(_009_)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    or_bb _396_ (
        .a(_009_),
        .b(_008_),
        .c(_010_)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    or_bb _397_ (
        .a(new_Jinkela_wire_209),
        .b(new_Jinkela_wire_175),
        .c(_011_)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    and_bb _398_ (
        .a(new_Jinkela_wire_208),
        .b(new_Jinkela_wire_174),
        .c(_012_)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    and_bi _399_ (
        .a(_011_),
        .b(_012_),
        .c(_013_)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    or_bi _400_ (
        .a(new_Jinkela_wire_631),
        .b(new_Jinkela_wire_305),
        .c(_014_)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    and_bi _401_ (
        .a(new_Jinkela_wire_632),
        .b(new_Jinkela_wire_308),
        .c(_015_)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_555),
        .dout(new_Jinkela_wire_556)
    );

    or_bi _402_ (
        .a(_015_),
        .b(_014_),
        .c(_016_)
    );

    or_bi _403_ (
        .a(new_Jinkela_wire_1326),
        .b(new_Jinkela_wire_1227),
        .c(_017_)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_627),
        .dout(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    and_bi _404_ (
        .a(new_Jinkela_wire_1327),
        .b(new_Jinkela_wire_1228),
        .c(_018_)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_578),
        .dout(new_Jinkela_wire_579)
    );

    and_bi _405_ (
        .a(_017_),
        .b(_018_),
        .c(_019_)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_557),
        .dout(new_Jinkela_wire_558)
    );

    or_bi _409_ (
        .a(_022_),
        .b(_021_),
        .c(_023_)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    or_bb _410_ (
        .a(new_Jinkela_wire_666),
        .b(new_Jinkela_wire_961),
        .c(_024_)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_558),
        .dout(new_Jinkela_wire_559)
    );

    and_bb _411_ (
        .a(new_Jinkela_wire_664),
        .b(new_Jinkela_wire_960),
        .c(_025_)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    and_bi _412_ (
        .a(_024_),
        .b(_025_),
        .c(_026_)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    or_bi _413_ (
        .a(new_Jinkela_wire_1022),
        .b(new_Jinkela_wire_856),
        .c(_027_)
    );

    and_bi _414_ (
        .a(new_Jinkela_wire_1023),
        .b(new_Jinkela_wire_857),
        .c(_028_)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    or_bi _415_ (
        .a(_028_),
        .b(_027_),
        .c(_029_)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    or_bi _416_ (
        .a(new_Jinkela_wire_1295),
        .b(new_Jinkela_wire_1613),
        .c(_030_)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_561),
        .c(new_Jinkela_wire_562),
        .b(new_Jinkela_wire_563)
    );

    and_bi _417_ (
        .a(new_Jinkela_wire_1296),
        .b(new_Jinkela_wire_1614),
        .c(_031_)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_581),
        .dout(new_Jinkela_wire_582)
    );

    and_bi _418_ (
        .a(_030_),
        .b(_031_),
        .c(_032_)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    or_bb _419_ (
        .a(new_Jinkela_wire_373),
        .b(new_Jinkela_wire_242),
        .c(_033_)
    );

    and_bb _420_ (
        .a(new_Jinkela_wire_374),
        .b(new_Jinkela_wire_243),
        .c(_034_)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    and_bi _421_ (
        .a(_033_),
        .b(_034_),
        .c(_035_)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    or_bi _422_ (
        .a(new_Jinkela_wire_597),
        .b(new_Jinkela_wire_5),
        .c(_036_)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    and_bi _423_ (
        .a(new_Jinkela_wire_599),
        .b(new_Jinkela_wire_1),
        .c(_037_)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_634),
        .dout(new_Jinkela_wire_635)
    );

    and_bi _424_ (
        .a(_036_),
        .b(_037_),
        .c(_038_)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_584),
        .dout(new_Jinkela_wire_585)
    );

    or_bi _425_ (
        .a(new_Jinkela_wire_1060),
        .b(new_Jinkela_wire_1368),
        .c(_039_)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    and_bi _426_ (
        .a(new_Jinkela_wire_1061),
        .b(new_Jinkela_wire_1369),
        .c(_040_)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    and_bi _427_ (
        .a(_039_),
        .b(_040_),
        .c(_041_)
    );

    spl4L new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_696),
        .d(new_Jinkela_wire_697),
        .e(new_Jinkela_wire_698),
        .c(new_Jinkela_wire_699),
        .b(new_Jinkela_wire_700)
    );

    or_bi _428_ (
        .a(new_Jinkela_wire_1292),
        .b(new_Jinkela_wire_1483),
        .c(_042_)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(G29),
        .c(new_Jinkela_wire_727),
        .b(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_586),
        .dout(new_Jinkela_wire_587)
    );

    and_bi _429_ (
        .a(new_Jinkela_wire_1293),
        .b(new_Jinkela_wire_1484),
        .c(_043_)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    and_bi _430_ (
        .a(_042_),
        .b(_043_),
        .c(_044_)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1122),
        .dout(new_Jinkela_wire_1123)
    );

    spl2 new_Jinkela_splitter_122 (
        .a(_121_),
        .c(new_Jinkela_wire_1135),
        .b(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1137),
        .dout(new_Jinkela_wire_1138)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1123),
        .dout(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_818 (
        .din(_234_),
        .dout(new_Jinkela_wire_1137)
    );

    spl4L new_Jinkela_splitter_124 (
        .a(_084_),
        .d(new_Jinkela_wire_1141),
        .e(new_Jinkela_wire_1142),
        .c(new_Jinkela_wire_1143),
        .b(new_Jinkela_wire_1144)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    spl2 new_Jinkela_splitter_123 (
        .a(_312_),
        .c(new_Jinkela_wire_1139),
        .b(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_1126),
        .dout(new_Jinkela_wire_1127)
    );

    spl2 new_Jinkela_splitter_127 (
        .a(_278_),
        .c(new_Jinkela_wire_1159),
        .b(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1127),
        .dout(new_Jinkela_wire_1128)
    );

    spl2 new_Jinkela_splitter_128 (
        .a(_085_),
        .c(new_Jinkela_wire_1161),
        .b(new_Jinkela_wire_1162)
    );

    spl2 new_Jinkela_splitter_130 (
        .a(_298_),
        .c(new_Jinkela_wire_1175),
        .b(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_1145),
        .dout(new_Jinkela_wire_1146)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_net_686),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_1146),
        .dout(new_Jinkela_wire_1147)
    );

    spl2 new_Jinkela_splitter_131 (
        .a(_152_),
        .c(new_Jinkela_wire_1177),
        .b(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1144),
        .dout(new_Jinkela_wire_1145)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_1147),
        .dout(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1172),
        .dout(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1163),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1148),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    spl2 new_Jinkela_splitter_133 (
        .a(_075_),
        .c(new_Jinkela_wire_1181),
        .b(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1164),
        .dout(new_Jinkela_wire_1165)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1173),
        .dout(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1151),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1165),
        .dout(new_Jinkela_wire_1166)
    );

    spl3L new_Jinkela_splitter_125 (
        .a(new_Jinkela_wire_1152),
        .d(new_Jinkela_wire_1153),
        .c(new_Jinkela_wire_1154),
        .b(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1155),
        .dout(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1166),
        .dout(new_Jinkela_wire_1167)
    );

    spl2 new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_1156),
        .c(new_Jinkela_wire_1157),
        .b(new_Jinkela_wire_1158)
    );

    spl2 new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_1167),
        .c(new_Jinkela_wire_1168),
        .b(new_Jinkela_wire_1169)
    );

    spl2 new_Jinkela_splitter_132 (
        .a(_340_),
        .c(new_Jinkela_wire_1179),
        .b(new_Jinkela_wire_1180)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1169),
        .dout(new_Jinkela_wire_1170)
    );

    spl2 new_Jinkela_splitter_134 (
        .a(_352_),
        .c(new_Jinkela_wire_1183),
        .b(new_Jinkela_wire_1184)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(_169_),
        .c(new_Jinkela_wire_1185),
        .b(new_Jinkela_wire_1186)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1170),
        .dout(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_net_682),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_843),
        .dout(new_Jinkela_wire_844)
    );

    or_bb _407_ (
        .a(new_Jinkela_wire_1355),
        .b(new_Jinkela_wire_1220),
        .c(_021_)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_317),
        .dout(new_Jinkela_wire_318)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_844),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    bfr new_Jinkela_buffer_644 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_845),
        .dout(new_Jinkela_wire_846)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_468),
        .d(new_Jinkela_wire_469),
        .e(new_Jinkela_wire_470),
        .c(new_Jinkela_wire_471),
        .b(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    spl2 new_Jinkela_splitter_93 (
        .a(G32),
        .c(new_Jinkela_wire_989),
        .b(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_318),
        .dout(new_Jinkela_wire_319)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_846),
        .dout(new_Jinkela_wire_847)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_319),
        .dout(new_Jinkela_wire_320)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_299),
        .dout(new_Jinkela_wire_300)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_320),
        .dout(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    spl2 new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_301),
        .c(new_Jinkela_wire_302),
        .b(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_321),
        .dout(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_871),
        .dout(new_Jinkela_wire_872)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_322),
        .dout(new_Jinkela_wire_323)
    );

    spl2 new_Jinkela_splitter_80 (
        .a(new_Jinkela_wire_853),
        .c(new_Jinkela_wire_854),
        .b(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_348),
        .dout(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_323),
        .dout(new_Jinkela_wire_324)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(G16),
        .c(new_Jinkela_wire_466),
        .b(new_Jinkela_wire_468)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_324),
        .dout(new_Jinkela_wire_325)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    spl4L new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_991),
        .d(new_Jinkela_wire_992),
        .e(new_Jinkela_wire_993),
        .c(new_Jinkela_wire_994),
        .b(new_Jinkela_wire_995)
    );

    spl4L new_Jinkela_splitter_91 (
        .a(new_Jinkela_wire_958),
        .d(new_Jinkela_wire_959),
        .e(new_Jinkela_wire_960),
        .c(new_Jinkela_wire_961),
        .b(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_325),
        .dout(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_326),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_350),
        .dout(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_876),
        .dout(new_Jinkela_wire_877)
    );

    spl3L new_Jinkela_splitter_48 (
        .a(G22),
        .d(new_Jinkela_wire_498),
        .c(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_500)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_877),
        .dout(new_Jinkela_wire_878)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_329),
        .dout(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_878),
        .dout(new_Jinkela_wire_879)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_879),
        .dout(new_Jinkela_wire_880)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_331),
        .dout(new_Jinkela_wire_332)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_58),
        .dout(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_588),
        .dout(new_Jinkela_wire_589)
    );

    spl2 new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_30),
        .c(new_Jinkela_wire_31),
        .b(new_Jinkela_wire_32)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_589),
        .dout(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_59),
        .dout(new_Jinkela_wire_60)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_590),
        .dout(new_Jinkela_wire_591)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_592),
        .dout(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    spl3L new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_143),
        .d(new_Jinkela_wire_144),
        .c(new_Jinkela_wire_145),
        .b(new_Jinkela_wire_146)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    spl2 new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_593),
        .c(new_Jinkela_wire_594),
        .b(new_Jinkela_wire_595)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_667),
        .dout(new_Jinkela_wire_668)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_694),
        .dout(new_Jinkela_wire_695)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_65),
        .dout(new_Jinkela_wire_66)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_87),
        .dout(new_Jinkela_wire_88)
    );

    spl2 new_Jinkela_splitter_72 (
        .a(G5),
        .c(new_Jinkela_wire_758),
        .b(new_Jinkela_wire_760)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_66),
        .dout(new_Jinkela_wire_67)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    spl3L new_Jinkela_splitter_21 (
        .a(G3),
        .d(new_Jinkela_wire_205),
        .c(new_Jinkela_wire_206),
        .b(new_Jinkela_wire_207)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_67),
        .dout(new_Jinkela_wire_68)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_88),
        .dout(new_Jinkela_wire_89)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_668),
        .dout(new_Jinkela_wire_669)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_617),
        .dout(new_Jinkela_wire_618)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_618),
        .dout(new_Jinkela_wire_619)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_70),
        .dout(new_Jinkela_wire_71)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_619),
        .dout(new_Jinkela_wire_620)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_146),
        .dout(new_Jinkela_wire_147)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_71),
        .dout(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_620),
        .dout(new_Jinkela_wire_621)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_669),
        .dout(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_621),
        .dout(new_Jinkela_wire_622)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_117),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    spl2 new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_73),
        .c(new_Jinkela_wire_74),
        .b(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_622),
        .dout(new_Jinkela_wire_623)
    );

    spl4L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_760),
        .d(new_Jinkela_wire_761),
        .e(new_Jinkela_wire_762),
        .c(new_Jinkela_wire_763),
        .b(new_Jinkela_wire_764)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_91),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_623),
        .dout(new_Jinkela_wire_624)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(new_Jinkela_wire_624),
        .c(new_Jinkela_wire_625),
        .b(new_Jinkela_wire_626)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_93),
        .dout(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    spl4L new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_173),
        .d(new_Jinkela_wire_174),
        .e(new_Jinkela_wire_175),
        .c(new_Jinkela_wire_176),
        .b(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_670),
        .dout(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_94),
        .dout(new_Jinkela_wire_95)
    );

    spl4L new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_729),
        .d(new_Jinkela_wire_730),
        .e(new_Jinkela_wire_731),
        .c(new_Jinkela_wire_732),
        .b(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_95),
        .dout(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    and_bi _599_ (
        .a(_205_),
        .b(new_Jinkela_wire_1095),
        .c(_213_)
    );

    or_bb _600_ (
        .a(new_Jinkela_wire_1591),
        .b(new_Jinkela_wire_1585),
        .c(_214_)
    );

    or_bb _601_ (
        .a(new_Jinkela_wire_1274),
        .b(new_Jinkela_wire_1171),
        .c(_215_)
    );

    or_bi _602_ (
        .a(new_Jinkela_wire_1195),
        .b(new_Jinkela_wire_1611),
        .c(_216_)
    );

    or_ii _603_ (
        .a(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_336),
        .c(_217_)
    );

    and_ii _604_ (
        .a(new_Jinkela_wire_1205),
        .b(new_Jinkela_wire_337),
        .c(_218_)
    );

    and_bi _605_ (
        .a(_217_),
        .b(_218_),
        .c(G1324)
    );

    and_bi _606_ (
        .a(new_Jinkela_wire_1136),
        .b(new_Jinkela_wire_1085),
        .c(_219_)
    );

    and_bi _607_ (
        .a(new_Jinkela_wire_1559),
        .b(new_Jinkela_wire_1229),
        .c(_220_)
    );

    and_bi _608_ (
        .a(new_Jinkela_wire_1579),
        .b(new_Jinkela_wire_1406),
        .c(_221_)
    );

    or_bb _609_ (
        .a(new_Jinkela_wire_1142),
        .b(new_Jinkela_wire_1374),
        .c(_222_)
    );

    or_bb _610_ (
        .a(new_Jinkela_wire_1645),
        .b(_221_),
        .c(_223_)
    );

    or_bi _611_ (
        .a(new_Jinkela_wire_1373),
        .b(new_Jinkela_wire_1143),
        .c(_224_)
    );

    or_ii _612_ (
        .a(new_Jinkela_wire_1118),
        .b(new_Jinkela_wire_1161),
        .c(_225_)
    );

    or_ii _613_ (
        .a(new_Jinkela_wire_1230),
        .b(new_Jinkela_wire_1558),
        .c(_226_)
    );

    and_bi _614_ (
        .a(_225_),
        .b(new_Jinkela_wire_1218),
        .c(_227_)
    );

    and_bi _615_ (
        .a(_223_),
        .b(new_Jinkela_wire_1115),
        .c(_228_)
    );

    or_bb _616_ (
        .a(new_Jinkela_wire_1108),
        .b(new_Jinkela_wire_1367),
        .c(_229_)
    );

    or_bb _617_ (
        .a(new_Jinkela_wire_1200),
        .b(new_Jinkela_wire_1480),
        .c(_230_)
    );

    or_bi _618_ (
        .a(new_Jinkela_wire_1524),
        .b(new_Jinkela_wire_1158),
        .c(_231_)
    );

    or_ii _619_ (
        .a(new_Jinkela_wire_1623),
        .b(new_Jinkela_wire_725),
        .c(_232_)
    );

    and_ii _620_ (
        .a(new_Jinkela_wire_1624),
        .b(new_Jinkela_wire_726),
        .c(_233_)
    );

    and_bi _621_ (
        .a(_232_),
        .b(_233_),
        .c(new_net_684)
    );

    or_bb _622_ (
        .a(new_Jinkela_wire_1503),
        .b(new_Jinkela_wire_1647),
        .c(_234_)
    );

    or_bb _623_ (
        .a(new_Jinkela_wire_1138),
        .b(new_Jinkela_wire_1107),
        .c(_235_)
    );

    or_bb _624_ (
        .a(new_Jinkela_wire_1336),
        .b(new_Jinkela_wire_1568),
        .c(_236_)
    );

    or_ii _625_ (
        .a(new_Jinkela_wire_1424),
        .b(new_Jinkela_wire_74),
        .c(_237_)
    );

    and_ii _626_ (
        .a(new_Jinkela_wire_1425),
        .b(new_Jinkela_wire_75),
        .c(_238_)
    );

    and_bi _627_ (
        .a(_237_),
        .b(_238_),
        .c(new_net_694)
    );

    or_bi _628_ (
        .a(new_Jinkela_wire_1194),
        .b(new_Jinkela_wire_1324),
        .c(_239_)
    );

    or_ii _629_ (
        .a(new_Jinkela_wire_1390),
        .b(new_Jinkela_wire_660),
        .c(_240_)
    );

    and_ii _630_ (
        .a(new_Jinkela_wire_1391),
        .b(new_Jinkela_wire_659),
        .c(_241_)
    );

    and_bi _631_ (
        .a(_240_),
        .b(_241_),
        .c(G1325)
    );

    or_bb _632_ (
        .a(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_1239),
        .c(_242_)
    );

    or_ii _633_ (
        .a(new_Jinkela_wire_1282),
        .b(new_Jinkela_wire_526),
        .c(_243_)
    );

    and_ii _634_ (
        .a(new_Jinkela_wire_1283),
        .b(new_Jinkela_wire_527),
        .c(_244_)
    );

    and_bi _635_ (
        .a(_243_),
        .b(_244_),
        .c(new_net_720)
    );

    or_bi _636_ (
        .a(new_Jinkela_wire_1335),
        .b(new_Jinkela_wire_1384),
        .c(_245_)
    );

    or_ii _637_ (
        .a(new_Jinkela_wire_1632),
        .b(new_Jinkela_wire_267),
        .c(_246_)
    );

    and_ii _638_ (
        .a(new_Jinkela_wire_1633),
        .b(new_Jinkela_wire_268),
        .c(_247_)
    );

    and_bi _639_ (
        .a(_246_),
        .b(_247_),
        .c(new_net_686)
    );

    or_bi _640_ (
        .a(new_Jinkela_wire_1338),
        .b(new_Jinkela_wire_1153),
        .c(_248_)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1545),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1529),
        .dout(new_Jinkela_wire_1530)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(new_Jinkela_wire_1509),
        .c(new_Jinkela_wire_1510),
        .b(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(new_Jinkela_wire_1511),
        .c(new_Jinkela_wire_1512),
        .b(new_Jinkela_wire_1513)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_354),
        .dout(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    spl2 new_Jinkela_splitter_241 (
        .a(_104_),
        .c(new_Jinkela_wire_1556),
        .b(new_Jinkela_wire_1557)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_335),
        .c(new_Jinkela_wire_336),
        .b(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    spl2 new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_1513),
        .c(new_Jinkela_wire_1514),
        .b(new_Jinkela_wire_1515)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1530),
        .dout(new_Jinkela_wire_1531)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1551),
        .dout(new_Jinkela_wire_1552)
    );

    spl3L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_436),
        .d(new_Jinkela_wire_437),
        .c(new_Jinkela_wire_438),
        .b(new_Jinkela_wire_439)
    );

    spl2 new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_885),
        .c(new_Jinkela_wire_886),
        .b(new_Jinkela_wire_887)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1531),
        .dout(new_Jinkela_wire_1532)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_762 (
        .din(G35),
        .dout(new_Jinkela_wire_1020)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_409),
        .dout(new_Jinkela_wire_410)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1532),
        .dout(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_381),
        .dout(new_Jinkela_wire_382)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1533),
        .dout(new_Jinkela_wire_1534)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(_108_),
        .c(new_Jinkela_wire_1586),
        .b(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_359),
        .dout(new_Jinkela_wire_360)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1552),
        .dout(new_Jinkela_wire_1553)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(new_Jinkela_wire_1548),
        .c(new_Jinkela_wire_1549),
        .b(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    spl2 new_Jinkela_splitter_247 (
        .a(new_Jinkela_wire_1578),
        .c(new_Jinkela_wire_1579),
        .b(new_Jinkela_wire_1580)
    );

    spl2 new_Jinkela_splitter_235 (
        .a(new_Jinkela_wire_1536),
        .c(new_Jinkela_wire_1537),
        .b(new_Jinkela_wire_1538)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    spl2 new_Jinkela_splitter_236 (
        .a(new_Jinkela_wire_1538),
        .c(new_Jinkela_wire_1539),
        .b(new_Jinkela_wire_1540)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_788 (
        .din(G38),
        .dout(new_Jinkela_wire_1054)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(new_Jinkela_wire_1540),
        .c(new_Jinkela_wire_1541),
        .b(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_363),
        .dout(new_Jinkela_wire_364)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1560),
        .dout(new_Jinkela_wire_1561)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    spl2 new_Jinkela_splitter_249 (
        .a(_203_),
        .c(new_Jinkela_wire_1588),
        .b(new_Jinkela_wire_1589)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(_269_),
        .c(new_Jinkela_wire_1574),
        .b(new_Jinkela_wire_1575)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_411),
        .dout(new_Jinkela_wire_412)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    bfr new_Jinkela_buffer_973 (
        .din(_124_),
        .dout(new_Jinkela_wire_1578)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_385),
        .dout(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(_201_),
        .c(new_Jinkela_wire_1576),
        .b(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_503),
        .dout(new_Jinkela_wire_504)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_937),
        .dout(new_Jinkela_wire_938)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    spl2 new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_367),
        .c(new_Jinkela_wire_368),
        .b(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_412),
        .dout(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    spl3L new_Jinkela_splitter_242 (
        .a(new_Jinkela_wire_1557),
        .d(new_Jinkela_wire_1558),
        .c(new_Jinkela_wire_1559),
        .b(new_Jinkela_wire_1560)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_386),
        .dout(new_Jinkela_wire_387)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    spl3L new_Jinkela_splitter_250 (
        .a(_213_),
        .d(new_Jinkela_wire_1590),
        .c(new_Jinkela_wire_1591),
        .b(new_Jinkela_wire_1592)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_387),
        .dout(new_Jinkela_wire_388)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    bfr new_Jinkela_buffer_988 (
        .din(_029_),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1564),
        .dout(new_Jinkela_wire_1565)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_388),
        .dout(new_Jinkela_wire_389)
    );

    spl3L new_Jinkela_splitter_96 (
        .a(G11),
        .d(new_Jinkela_wire_1022),
        .c(new_Jinkela_wire_1023),
        .b(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1565),
        .dout(new_Jinkela_wire_1566)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_413),
        .dout(new_Jinkela_wire_414)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_919),
        .c(new_Jinkela_wire_920),
        .b(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_971 (
        .din(new_Jinkela_wire_1566),
        .dout(new_Jinkela_wire_1567)
    );

    spl3L new_Jinkela_splitter_54 (
        .a(G26),
        .d(new_Jinkela_wire_564),
        .c(new_Jinkela_wire_565),
        .b(new_Jinkela_wire_566)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    spl4L new_Jinkela_splitter_251 (
        .a(_010_),
        .d(new_Jinkela_wire_1593),
        .e(new_Jinkela_wire_1594),
        .c(new_Jinkela_wire_1595),
        .b(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_390),
        .dout(new_Jinkela_wire_391)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1582),
        .dout(new_Jinkela_wire_1583)
    );

    spl3L new_Jinkela_splitter_243 (
        .a(new_Jinkela_wire_1567),
        .d(new_Jinkela_wire_1568),
        .c(new_Jinkela_wire_1569),
        .b(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    and_bi _431_ (
        .a(new_Jinkela_wire_1131),
        .b(new_Jinkela_wire_1456),
        .c(_045_)
    );

    and_bi _432_ (
        .a(new_Jinkela_wire_1457),
        .b(new_Jinkela_wire_1132),
        .c(_046_)
    );

    or_bb _433_ (
        .a(_046_),
        .b(_045_),
        .c(_047_)
    );

    or_bb _434_ (
        .a(new_Jinkela_wire_893),
        .b(new_Jinkela_wire_274),
        .c(_048_)
    );

    and_bb _435_ (
        .a(new_Jinkela_wire_889),
        .b(new_Jinkela_wire_275),
        .c(_049_)
    );

    and_bi _436_ (
        .a(_048_),
        .b(_049_),
        .c(_050_)
    );

    or_bi _437_ (
        .a(new_Jinkela_wire_761),
        .b(new_Jinkela_wire_533),
        .c(_051_)
    );

    and_bi _438_ (
        .a(new_Jinkela_wire_762),
        .b(new_Jinkela_wire_531),
        .c(_052_)
    );

    or_bi _439_ (
        .a(_052_),
        .b(_051_),
        .c(_053_)
    );

    or_bi _440_ (
        .a(new_Jinkela_wire_1214),
        .b(new_Jinkela_wire_1096),
        .c(_054_)
    );

    and_bi _441_ (
        .a(new_Jinkela_wire_1215),
        .b(new_Jinkela_wire_1097),
        .c(_055_)
    );

    and_bi _442_ (
        .a(_054_),
        .b(_055_),
        .c(_056_)
    );

    and_bb _443_ (
        .a(new_Jinkela_wire_1057),
        .b(new_Jinkela_wire_36),
        .c(_057_)
    );

    or_bb _444_ (
        .a(new_Jinkela_wire_1652),
        .b(new_Jinkela_wire_1629),
        .c(_058_)
    );

    and_bb _445_ (
        .a(new_Jinkela_wire_1653),
        .b(new_Jinkela_wire_1628),
        .c(_059_)
    );

    or_bi _446_ (
        .a(_059_),
        .b(_058_),
        .c(_060_)
    );

    or_bb _447_ (
        .a(new_Jinkela_wire_925),
        .b(new_Jinkela_wire_470),
        .c(_061_)
    );

    and_bb _448_ (
        .a(new_Jinkela_wire_927),
        .b(new_Jinkela_wire_471),
        .c(_062_)
    );

    and_bi _449_ (
        .a(_061_),
        .b(_062_),
        .c(_063_)
    );

    or_bi _450_ (
        .a(new_Jinkela_wire_825),
        .b(new_Jinkela_wire_407),
        .c(_064_)
    );

    and_bi _451_ (
        .a(new_Jinkela_wire_829),
        .b(new_Jinkela_wire_406),
        .c(_065_)
    );

    or_bi _452_ (
        .a(_065_),
        .b(_064_),
        .c(_066_)
    );

    or_bi _453_ (
        .a(new_Jinkela_wire_1466),
        .b(new_Jinkela_wire_1481),
        .c(_067_)
    );

    and_bi _454_ (
        .a(new_Jinkela_wire_1467),
        .b(new_Jinkela_wire_1482),
        .c(_068_)
    );

    and_bi _455_ (
        .a(_067_),
        .b(_068_),
        .c(_069_)
    );

    or_bb _456_ (
        .a(new_Jinkela_wire_109),
        .b(new_Jinkela_wire_699),
        .c(_070_)
    );

    and_bb _457_ (
        .a(new_Jinkela_wire_111),
        .b(new_Jinkela_wire_697),
        .c(_071_)
    );

    and_bi _458_ (
        .a(_070_),
        .b(_071_),
        .c(_072_)
    );

    or_bi _459_ (
        .a(new_Jinkela_wire_795),
        .b(new_Jinkela_wire_990),
        .c(_073_)
    );

    and_bi _460_ (
        .a(new_Jinkela_wire_796),
        .b(new_Jinkela_wire_993),
        .c(_074_)
    );

    and_bi _461_ (
        .a(_073_),
        .b(_074_),
        .c(_075_)
    );

    or_bi _462_ (
        .a(new_Jinkela_wire_1129),
        .b(new_Jinkela_wire_1181),
        .c(_076_)
    );

    and_bi _463_ (
        .a(new_Jinkela_wire_1130),
        .b(new_Jinkela_wire_1182),
        .c(_077_)
    );

    and_bi _464_ (
        .a(_076_),
        .b(_077_),
        .c(_078_)
    );

    or_bi _465_ (
        .a(new_Jinkela_wire_1071),
        .b(new_Jinkela_wire_1370),
        .c(_079_)
    );

    and_bi _466_ (
        .a(new_Jinkela_wire_1073),
        .b(new_Jinkela_wire_1371),
        .c(_080_)
    );

    and_bi _467_ (
        .a(_079_),
        .b(_080_),
        .c(_081_)
    );

    and_bi _468_ (
        .a(new_Jinkela_wire_1404),
        .b(new_Jinkela_wire_1253),
        .c(_082_)
    );

    and_bi _469_ (
        .a(new_Jinkela_wire_1254),
        .b(new_Jinkela_wire_1405),
        .c(_083_)
    );

    or_bb _470_ (
        .a(_083_),
        .b(_082_),
        .c(_084_)
    );

    or_bi _471_ (
        .a(new_Jinkela_wire_1141),
        .b(new_Jinkela_wire_1372),
        .c(_085_)
    );

    or_ii _472_ (
        .a(new_Jinkela_wire_44),
        .b(new_Jinkela_wire_42),
        .c(_086_)
    );

    and_bb _408_ (
        .a(new_Jinkela_wire_1356),
        .b(new_Jinkela_wire_1219),
        .c(_022_)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    spl4L new_Jinkela_splitter_137 (
        .a(_288_),
        .d(new_Jinkela_wire_1190),
        .e(new_Jinkela_wire_1191),
        .c(new_Jinkela_wire_1192),
        .b(new_Jinkela_wire_1193)
    );

    spl4L new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_240),
        .d(new_Jinkela_wire_241),
        .e(new_Jinkela_wire_242),
        .c(new_Jinkela_wire_243),
        .b(new_Jinkela_wire_244)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(_149_),
        .c(new_Jinkela_wire_1198),
        .b(new_Jinkela_wire_1199)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    spl2 new_Jinkela_splitter_136 (
        .a(_261_),
        .c(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    spl4L new_Jinkela_splitter_138 (
        .a(_215_),
        .d(new_Jinkela_wire_1194),
        .e(new_Jinkela_wire_1195),
        .c(new_Jinkela_wire_1196),
        .b(new_Jinkela_wire_1197)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(_229_),
        .c(new_Jinkela_wire_1200),
        .b(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_147),
        .dout(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    spl2 new_Jinkela_splitter_141 (
        .a(_325_),
        .c(new_Jinkela_wire_1202),
        .b(new_Jinkela_wire_1203)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    spl2 new_Jinkela_splitter_142 (
        .a(_216_),
        .c(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_1205)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(G23),
        .c(new_Jinkela_wire_238),
        .b(new_Jinkela_wire_240)
    );

    spl2 new_Jinkela_splitter_143 (
        .a(_258_),
        .c(new_Jinkela_wire_1206),
        .b(new_Jinkela_wire_1207)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(_295_),
        .c(new_Jinkela_wire_1212),
        .b(new_Jinkela_wire_1213)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_100),
        .dout(new_Jinkela_wire_101)
    );

    spl2 new_Jinkela_splitter_144 (
        .a(_284_),
        .c(new_Jinkela_wire_1208),
        .b(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(_252_),
        .c(new_Jinkela_wire_1210),
        .b(new_Jinkela_wire_1211)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_101),
        .dout(new_Jinkela_wire_102)
    );

    bfr new_Jinkela_buffer_840 (
        .din(_226_),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(_050_),
        .c(new_Jinkela_wire_1214),
        .b(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_102),
        .dout(new_Jinkela_wire_103)
    );

    spl2 new_Jinkela_splitter_148 (
        .a(_195_),
        .c(new_Jinkela_wire_1216),
        .b(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    spl2 new_Jinkela_splitter_151 (
        .a(_016_),
        .c(new_Jinkela_wire_1227),
        .b(new_Jinkela_wire_1228)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_net_702),
        .dout(new_Jinkela_wire_1223)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    spl4L new_Jinkela_splitter_149 (
        .a(_019_),
        .d(new_Jinkela_wire_1219),
        .e(new_Jinkela_wire_1220),
        .c(new_Jinkela_wire_1221),
        .b(new_Jinkela_wire_1222)
    );

    bfr new_Jinkela_buffer_195 (
        .din(G39),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    spl2 new_Jinkela_splitter_150 (
        .a(new_Jinkela_wire_1224),
        .c(new_Jinkela_wire_1225),
        .b(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_104),
        .dout(new_Jinkela_wire_105)
    );

    spl2 new_Jinkela_splitter_158 (
        .a(_182_),
        .c(new_Jinkela_wire_1255),
        .b(new_Jinkela_wire_1256)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_842 (
        .din(_172_),
        .dout(new_Jinkela_wire_1224)
    );

    spl3L new_Jinkela_splitter_152 (
        .a(_219_),
        .d(new_Jinkela_wire_1229),
        .c(new_Jinkela_wire_1230),
        .b(new_Jinkela_wire_1231)
    );

    spl2 new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_105),
        .c(new_Jinkela_wire_106),
        .b(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    spl2 new_Jinkela_splitter_155 (
        .a(_166_),
        .c(new_Jinkela_wire_1245),
        .b(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    spl2 new_Jinkela_splitter_160 (
        .a(_202_),
        .c(new_Jinkela_wire_1259),
        .b(new_Jinkela_wire_1260)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1247),
        .dout(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1232),
        .dout(new_Jinkela_wire_1233)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    spl2 new_Jinkela_splitter_157 (
        .a(_060_),
        .c(new_Jinkela_wire_1253),
        .b(new_Jinkela_wire_1254)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1233),
        .dout(new_Jinkela_wire_1234)
    );

    spl3L new_Jinkela_splitter_27 (
        .a(G7),
        .d(new_Jinkela_wire_271),
        .c(new_Jinkela_wire_272),
        .b(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1231),
        .dout(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1234),
        .dout(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1248),
        .dout(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_178),
        .dout(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_851 (
        .din(_086_),
        .dout(new_Jinkela_wire_1247)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1235),
        .dout(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    spl2 new_Jinkela_splitter_159 (
        .a(_111_),
        .c(new_Jinkela_wire_1257),
        .b(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1236),
        .dout(new_Jinkela_wire_1237)
    );

    spl3L new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_207),
        .d(new_Jinkela_wire_208),
        .c(new_Jinkela_wire_209),
        .b(new_Jinkela_wire_210)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_1237),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    spl3L new_Jinkela_splitter_153 (
        .a(new_Jinkela_wire_1238),
        .d(new_Jinkela_wire_1239),
        .c(new_Jinkela_wire_1240),
        .b(new_Jinkela_wire_1241)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_179),
        .dout(new_Jinkela_wire_180)
    );

    spl2 new_Jinkela_splitter_156 (
        .a(new_Jinkela_wire_1250),
        .c(new_Jinkela_wire_1251),
        .b(new_Jinkela_wire_1252)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1241),
        .dout(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_154),
        .dout(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_855 (
        .din(_125_),
        .dout(new_Jinkela_wire_1261)
    );

    spl4L new_Jinkela_splitter_162 (
        .a(_302_),
        .d(new_Jinkela_wire_1267),
        .e(new_Jinkela_wire_1268),
        .c(new_Jinkela_wire_1269),
        .b(new_Jinkela_wire_1270)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    spl2 new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_1242),
        .c(new_Jinkela_wire_1243),
        .b(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(_114_),
        .c(new_Jinkela_wire_1271),
        .b(new_Jinkela_wire_1272)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1261),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_net_692),
        .dout(new_Jinkela_wire_1273)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    spl2 new_Jinkela_splitter_166 (
        .a(_242_),
        .c(new_Jinkela_wire_1282),
        .b(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1280),
        .dout(new_Jinkela_wire_1281)
    );

    spl4L new_Jinkela_splitter_165 (
        .a(_251_),
        .d(new_Jinkela_wire_1276),
        .e(new_Jinkela_wire_1277),
        .c(new_Jinkela_wire_1278),
        .b(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(new_Jinkela_wire_1264),
        .c(new_Jinkela_wire_1265),
        .b(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_net_696),
        .dout(new_Jinkela_wire_1280)
    );

    spl3L new_Jinkela_splitter_75 (
        .a(G28),
        .d(new_Jinkela_wire_792),
        .c(new_Jinkela_wire_793),
        .b(new_Jinkela_wire_794)
    );

    spl2 new_Jinkela_splitter_164 (
        .a(_214_),
        .c(new_Jinkela_wire_1274),
        .b(new_Jinkela_wire_1275)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    spl2 new_Jinkela_splitter_171 (
        .a(_158_),
        .c(new_Jinkela_wire_1297),
        .b(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_net_726),
        .dout(new_Jinkela_wire_1284)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    spl4L new_Jinkela_splitter_168 (
        .a(_355_),
        .d(new_Jinkela_wire_1287),
        .e(new_Jinkela_wire_1288),
        .c(new_Jinkela_wire_1289),
        .b(new_Jinkela_wire_1290)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_702),
        .dout(new_Jinkela_wire_703)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(_178_),
        .c(new_Jinkela_wire_1285),
        .b(new_Jinkela_wire_1286)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    spl2 new_Jinkela_splitter_170 (
        .a(_026_),
        .c(new_Jinkela_wire_1295),
        .b(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    spl4L new_Jinkela_splitter_169 (
        .a(_032_),
        .d(new_Jinkela_wire_1291),
        .e(new_Jinkela_wire_1292),
        .c(new_Jinkela_wire_1293),
        .b(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    spl2 new_Jinkela_splitter_174 (
        .a(_004_),
        .c(new_Jinkela_wire_1303),
        .b(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_676),
        .dout(new_Jinkela_wire_677)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(_128_),
        .c(new_Jinkela_wire_1299),
        .b(new_Jinkela_wire_1300)
    );

    spl2 new_Jinkela_splitter_173 (
        .a(_001_),
        .c(new_Jinkela_wire_1301),
        .b(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    spl2 new_Jinkela_splitter_180 (
        .a(_013_),
        .c(new_Jinkela_wire_1326),
        .b(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(_180_),
        .c(new_Jinkela_wire_1305),
        .b(new_Jinkela_wire_1306)
    );

    spl4L new_Jinkela_splitter_184 (
        .a(_235_),
        .d(new_Jinkela_wire_1335),
        .e(new_Jinkela_wire_1336),
        .c(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_1338)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    spl4L new_Jinkela_splitter_176 (
        .a(_161_),
        .d(new_Jinkela_wire_1307),
        .e(new_Jinkela_wire_1308),
        .c(new_Jinkela_wire_1309),
        .b(new_Jinkela_wire_1310)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(_179_),
        .c(new_Jinkela_wire_1328),
        .b(new_Jinkela_wire_1329)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1310),
        .dout(new_Jinkela_wire_1311)
    );

    spl2 new_Jinkela_splitter_183 (
        .a(new_Jinkela_wire_1332),
        .c(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1334)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_658),
        .c(new_Jinkela_wire_659),
        .b(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_872 (
        .din(_117_),
        .dout(new_Jinkela_wire_1332)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_1311),
        .dout(new_Jinkela_wire_1312)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_704),
        .dout(new_Jinkela_wire_705)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(_131_),
        .c(new_Jinkela_wire_1330),
        .b(new_Jinkela_wire_1331)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_678),
        .dout(new_Jinkela_wire_679)
    );

    spl2 new_Jinkela_splitter_185 (
        .a(_155_),
        .c(new_Jinkela_wire_1339),
        .b(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1312),
        .dout(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1313),
        .dout(new_Jinkela_wire_1314)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_705),
        .dout(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1314),
        .dout(new_Jinkela_wire_1315)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_682),
        .dout(new_Jinkela_wire_683)
    );

    spl2 new_Jinkela_splitter_186 (
        .a(_289_),
        .c(new_Jinkela_wire_1341),
        .b(new_Jinkela_wire_1342)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1315),
        .dout(new_Jinkela_wire_1316)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_877 (
        .din(_020_),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1316),
        .dout(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    spl2 new_Jinkela_splitter_187 (
        .a(_275_),
        .c(new_Jinkela_wire_1343),
        .b(new_Jinkela_wire_1344)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_873 (
        .din(_287_),
        .dout(new_Jinkela_wire_1345)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1317),
        .dout(new_Jinkela_wire_1318)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    spl2 new_Jinkela_splitter_188 (
        .a(_092_),
        .c(new_Jinkela_wire_1349),
        .b(new_Jinkela_wire_1350)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1318),
        .dout(new_Jinkela_wire_1319)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_391),
        .dout(new_Jinkela_wire_392)
    );

    or_ii _641_ (
        .a(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_137),
        .c(_249_)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_441),
        .dout(new_Jinkela_wire_442)
    );

    and_ii _642_ (
        .a(new_Jinkela_wire_1555),
        .b(new_Jinkela_wire_138),
        .c(_250_)
    );

    bfr new_Jinkela_buffer_991 (
        .din(_163_),
        .dout(new_Jinkela_wire_1617)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_392),
        .dout(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1583),
        .dout(new_Jinkela_wire_1584)
    );

    and_bi _643_ (
        .a(_249_),
        .b(_250_),
        .c(new_net_712)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(new_Jinkela_wire_1571),
        .c(new_Jinkela_wire_1572),
        .b(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    or_bb _644_ (
        .a(new_Jinkela_wire_1201),
        .b(new_Jinkela_wire_1436),
        .c(_251_)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(new_Jinkela_wire_1612),
        .c(new_Jinkela_wire_1613),
        .b(new_Jinkela_wire_1614)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_393),
        .dout(new_Jinkela_wire_394)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1584),
        .dout(new_Jinkela_wire_1585)
    );

    or_bb _645_ (
        .a(new_Jinkela_wire_1277),
        .b(new_Jinkela_wire_1572),
        .c(_252_)
    );

    bfr new_Jinkela_buffer_390 (
        .din(G36),
        .dout(new_Jinkela_wire_528)
    );

    or_ii _646_ (
        .a(new_Jinkela_wire_1210),
        .b(new_Jinkela_wire_368),
        .c(_253_)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_394),
        .dout(new_Jinkela_wire_395)
    );

    and_ii _647_ (
        .a(new_Jinkela_wire_1211),
        .b(new_Jinkela_wire_369),
        .c(_254_)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_416),
        .dout(new_Jinkela_wire_417)
    );

    and_bi _648_ (
        .a(_253_),
        .b(_254_),
        .c(new_net_702)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    or_bb _649_ (
        .a(new_Jinkela_wire_1278),
        .b(new_Jinkela_wire_1244),
        .c(_255_)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(new_Jinkela_wire_1625),
        .c(new_Jinkela_wire_1626),
        .b(new_Jinkela_wire_1627)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_442),
        .dout(new_Jinkela_wire_443)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(_231_),
        .c(new_Jinkela_wire_1623),
        .b(new_Jinkela_wire_1624)
    );

    or_ii _650_ (
        .a(new_Jinkela_wire_1058),
        .b(new_Jinkela_wire_595),
        .c(_256_)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    and_ii _651_ (
        .a(new_Jinkela_wire_1059),
        .b(new_Jinkela_wire_594),
        .c(_257_)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1615),
        .dout(new_Jinkela_wire_1616)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_417),
        .dout(new_Jinkela_wire_418)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_net_714),
        .dout(new_Jinkela_wire_1615)
    );

    and_bi _652_ (
        .a(_256_),
        .b(_257_),
        .c(new_net_688)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    or_bi _653_ (
        .a(new_Jinkela_wire_1279),
        .b(new_Jinkela_wire_1388),
        .c(_258_)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_472),
        .dout(new_Jinkela_wire_473)
    );

    or_ii _654_ (
        .a(new_Jinkela_wire_1206),
        .b(new_Jinkela_wire_32),
        .c(_259_)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(G6),
        .c(new_Jinkela_wire_530),
        .b(new_Jinkela_wire_532)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1617),
        .dout(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    and_ii _655_ (
        .a(new_Jinkela_wire_1207),
        .b(new_Jinkela_wire_31),
        .c(_260_)
    );

    bfr new_Jinkela_buffer_995 (
        .din(_140_),
        .dout(new_Jinkela_wire_1625)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_418),
        .dout(new_Jinkela_wire_419)
    );

    and_bi _656_ (
        .a(_259_),
        .b(_260_),
        .c(new_net_700)
    );

    spl2 new_Jinkela_splitter_38 (
        .a(new_Jinkela_wire_399),
        .c(new_Jinkela_wire_400),
        .b(new_Jinkela_wire_401)
    );

    spl4L new_Jinkela_splitter_259 (
        .a(_056_),
        .d(new_Jinkela_wire_1628),
        .e(new_Jinkela_wire_1629),
        .c(new_Jinkela_wire_1630),
        .b(new_Jinkela_wire_1631)
    );

    or_bi _657_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_1157),
        .c(_261_)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1601),
        .dout(new_Jinkela_wire_1602)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_419),
        .dout(new_Jinkela_wire_420)
    );

    or_ii _658_ (
        .a(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_822),
        .c(_262_)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_443),
        .dout(new_Jinkela_wire_444)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1618),
        .dout(new_Jinkela_wire_1619)
    );

    and_ii _659_ (
        .a(new_Jinkela_wire_1189),
        .b(new_Jinkela_wire_823),
        .c(_263_)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    and_bi _660_ (
        .a(_262_),
        .b(_263_),
        .c(new_net_682)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_420),
        .dout(new_Jinkela_wire_421)
    );

    or_bb _661_ (
        .a(new_Jinkela_wire_1502),
        .b(new_Jinkela_wire_1256),
        .c(_264_)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_444),
        .dout(new_Jinkela_wire_445)
    );

    or_bb _662_ (
        .a(new_Jinkela_wire_1635),
        .b(new_Jinkela_wire_1109),
        .c(_265_)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(_245_),
        .c(new_Jinkela_wire_1632),
        .b(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_421),
        .dout(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1619),
        .dout(new_Jinkela_wire_1620)
    );

    or_bb _663_ (
        .a(new_Jinkela_wire_1099),
        .b(new_Jinkela_wire_1569),
        .c(_266_)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    and_bi _664_ (
        .a(new_Jinkela_wire_1636),
        .b(new_Jinkela_wire_756),
        .c(_267_)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_422),
        .dout(new_Jinkela_wire_423)
    );

    and_bi _665_ (
        .a(new_Jinkela_wire_757),
        .b(new_Jinkela_wire_1637),
        .c(_268_)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(new_Jinkela_wire_1605),
        .c(new_Jinkela_wire_1606),
        .b(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_445),
        .dout(new_Jinkela_wire_446)
    );

    or_bb _666_ (
        .a(_268_),
        .b(_267_),
        .c(new_net_728)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(new_Jinkela_wire_1607),
        .c(new_Jinkela_wire_1608),
        .b(new_Jinkela_wire_1609)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_423),
        .dout(new_Jinkela_wire_424)
    );

    or_bb _667_ (
        .a(new_Jinkela_wire_1098),
        .b(new_Jinkela_wire_1240),
        .c(_269_)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(new_Jinkela_wire_1620),
        .c(new_Jinkela_wire_1621),
        .b(new_Jinkela_wire_1622)
    );

    or_ii _668_ (
        .a(new_Jinkela_wire_1574),
        .b(new_Jinkela_wire_170),
        .c(_270_)
    );

    spl3L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_500),
        .d(new_Jinkela_wire_501),
        .c(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_503)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(new_Jinkela_wire_1609),
        .c(new_Jinkela_wire_1610),
        .b(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_424),
        .dout(new_Jinkela_wire_425)
    );

    and_ii _669_ (
        .a(new_Jinkela_wire_1575),
        .b(new_Jinkela_wire_169),
        .c(_271_)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_446),
        .dout(new_Jinkela_wire_447)
    );

    and_bi _670_ (
        .a(_270_),
        .b(_271_),
        .c(new_net_706)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_425),
        .dout(new_Jinkela_wire_426)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    or_bi _671_ (
        .a(new_Jinkela_wire_1100),
        .b(new_Jinkela_wire_1385),
        .c(_272_)
    );

    bfr new_Jinkela_buffer_996 (
        .din(_264_),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_474),
        .dout(new_Jinkela_wire_475)
    );

    or_ii _672_ (
        .a(new_Jinkela_wire_1068),
        .b(new_Jinkela_wire_626),
        .c(_273_)
    );

    spl4L new_Jinkela_splitter_262 (
        .a(_315_),
        .d(new_Jinkela_wire_1638),
        .e(new_Jinkela_wire_1639),
        .c(new_Jinkela_wire_1640),
        .b(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_426),
        .dout(new_Jinkela_wire_427)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(_266_),
        .c(new_Jinkela_wire_1636),
        .b(new_Jinkela_wire_1637)
    );

    and_ii _673_ (
        .a(new_Jinkela_wire_1069),
        .b(new_Jinkela_wire_625),
        .c(_274_)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(_184_),
        .c(new_Jinkela_wire_1646),
        .b(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_447),
        .dout(new_Jinkela_wire_448)
    );

    bfr new_Jinkela_buffer_999 (
        .din(_222_),
        .dout(new_Jinkela_wire_1643)
    );

    and_bi _674_ (
        .a(_273_),
        .b(_274_),
        .c(new_net_708)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_427),
        .dout(new_Jinkela_wire_428)
    );

    or_bi _675_ (
        .a(new_Jinkela_wire_1101),
        .b(new_Jinkela_wire_1154),
        .c(_275_)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_net_698),
        .dout(new_Jinkela_wire_1642)
    );

    and_bi _676_ (
        .a(new_Jinkela_wire_1343),
        .b(new_Jinkela_wire_1018),
        .c(_276_)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    and_bi _677_ (
        .a(new_Jinkela_wire_1019),
        .b(new_Jinkela_wire_1344),
        .c(_277_)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(_057_),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    or_bb _678_ (
        .a(_277_),
        .b(_276_),
        .c(new_net_710)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    or_bi _679_ (
        .a(new_Jinkela_wire_1526),
        .b(new_Jinkela_wire_1389),
        .c(_278_)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1644),
        .dout(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_475),
        .dout(new_Jinkela_wire_476)
    );

    or_ii _680_ (
        .a(new_Jinkela_wire_1159),
        .b(new_Jinkela_wire_400),
        .c(_279_)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_430),
        .dout(new_Jinkela_wire_431)
    );

    and_ii _681_ (
        .a(new_Jinkela_wire_1160),
        .b(new_Jinkela_wire_401),
        .c(_280_)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    and_bi _682_ (
        .a(_279_),
        .b(_280_),
        .c(new_net_690)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    spl3L new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_1024),
        .d(new_Jinkela_wire_1025),
        .c(new_Jinkela_wire_1026),
        .b(new_Jinkela_wire_1027)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_1054),
        .dout(new_Jinkela_wire_1055)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_969),
        .dout(new_Jinkela_wire_970)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_948),
        .dout(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    spl2 new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_951),
        .c(new_Jinkela_wire_952),
        .b(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_972),
        .dout(new_Jinkela_wire_973)
    );

    spl2 new_Jinkela_splitter_99 (
        .a(_255_),
        .c(new_Jinkela_wire_1058),
        .b(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_790 (
        .din(G40),
        .dout(new_Jinkela_wire_1056)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_976),
        .dout(new_Jinkela_wire_977)
    );

    spl2 new_Jinkela_splitter_100 (
        .a(_035_),
        .c(new_Jinkela_wire_1060),
        .b(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1056),
        .dout(new_Jinkela_wire_1057)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_980),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

endmodule
